library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(5119 downto 0);
    signal layer1_outputs : std_logic_vector(5119 downto 0);
    signal layer2_outputs : std_logic_vector(5119 downto 0);

begin

    layer0_outputs(0) <= not((inputs(223)) xor (inputs(222)));
    layer0_outputs(1) <= not((inputs(202)) and (inputs(79)));
    layer0_outputs(2) <= '1';
    layer0_outputs(3) <= (inputs(25)) xor (inputs(148));
    layer0_outputs(4) <= (inputs(156)) or (inputs(187));
    layer0_outputs(5) <= not((inputs(234)) xor (inputs(98)));
    layer0_outputs(6) <= (inputs(68)) or (inputs(238));
    layer0_outputs(7) <= '1';
    layer0_outputs(8) <= not(inputs(164));
    layer0_outputs(9) <= (inputs(50)) and not (inputs(109));
    layer0_outputs(10) <= (inputs(149)) or (inputs(151));
    layer0_outputs(11) <= (inputs(211)) or (inputs(83));
    layer0_outputs(12) <= (inputs(230)) or (inputs(138));
    layer0_outputs(13) <= not(inputs(122)) or (inputs(207));
    layer0_outputs(14) <= (inputs(23)) and not (inputs(16));
    layer0_outputs(15) <= inputs(40);
    layer0_outputs(16) <= not(inputs(115)) or (inputs(20));
    layer0_outputs(17) <= not((inputs(191)) xor (inputs(219)));
    layer0_outputs(18) <= (inputs(77)) xor (inputs(43));
    layer0_outputs(19) <= inputs(48);
    layer0_outputs(20) <= not(inputs(73));
    layer0_outputs(21) <= not(inputs(43)) or (inputs(145));
    layer0_outputs(22) <= '0';
    layer0_outputs(23) <= (inputs(75)) xor (inputs(92));
    layer0_outputs(24) <= '1';
    layer0_outputs(25) <= (inputs(67)) and not (inputs(143));
    layer0_outputs(26) <= (inputs(124)) and not (inputs(172));
    layer0_outputs(27) <= not(inputs(35));
    layer0_outputs(28) <= (inputs(108)) or (inputs(124));
    layer0_outputs(29) <= (inputs(188)) and not (inputs(0));
    layer0_outputs(30) <= not(inputs(155)) or (inputs(250));
    layer0_outputs(31) <= (inputs(84)) and (inputs(52));
    layer0_outputs(32) <= not((inputs(6)) or (inputs(93)));
    layer0_outputs(33) <= (inputs(219)) or (inputs(169));
    layer0_outputs(34) <= '1';
    layer0_outputs(35) <= '0';
    layer0_outputs(36) <= '0';
    layer0_outputs(37) <= not((inputs(5)) or (inputs(193)));
    layer0_outputs(38) <= '0';
    layer0_outputs(39) <= '0';
    layer0_outputs(40) <= not(inputs(185)) or (inputs(26));
    layer0_outputs(41) <= inputs(91);
    layer0_outputs(42) <= inputs(196);
    layer0_outputs(43) <= (inputs(120)) and not (inputs(31));
    layer0_outputs(44) <= not(inputs(165));
    layer0_outputs(45) <= not((inputs(221)) xor (inputs(57)));
    layer0_outputs(46) <= (inputs(154)) or (inputs(132));
    layer0_outputs(47) <= not(inputs(146)) or (inputs(248));
    layer0_outputs(48) <= not(inputs(77)) or (inputs(252));
    layer0_outputs(49) <= (inputs(14)) xor (inputs(57));
    layer0_outputs(50) <= (inputs(0)) and (inputs(171));
    layer0_outputs(51) <= inputs(151);
    layer0_outputs(52) <= (inputs(152)) and not (inputs(253));
    layer0_outputs(53) <= not((inputs(145)) xor (inputs(86)));
    layer0_outputs(54) <= not(inputs(170)) or (inputs(41));
    layer0_outputs(55) <= '0';
    layer0_outputs(56) <= not(inputs(0));
    layer0_outputs(57) <= '1';
    layer0_outputs(58) <= (inputs(23)) and not (inputs(139));
    layer0_outputs(59) <= not((inputs(167)) or (inputs(245)));
    layer0_outputs(60) <= not(inputs(219));
    layer0_outputs(61) <= (inputs(179)) and not (inputs(61));
    layer0_outputs(62) <= not((inputs(208)) or (inputs(224)));
    layer0_outputs(63) <= not(inputs(128));
    layer0_outputs(64) <= inputs(245);
    layer0_outputs(65) <= not((inputs(243)) xor (inputs(184)));
    layer0_outputs(66) <= inputs(80);
    layer0_outputs(67) <= not(inputs(125));
    layer0_outputs(68) <= not(inputs(208));
    layer0_outputs(69) <= (inputs(84)) and not (inputs(194));
    layer0_outputs(70) <= not(inputs(183)) or (inputs(7));
    layer0_outputs(71) <= '0';
    layer0_outputs(72) <= inputs(243);
    layer0_outputs(73) <= not(inputs(86));
    layer0_outputs(74) <= not((inputs(0)) or (inputs(52)));
    layer0_outputs(75) <= not(inputs(239)) or (inputs(11));
    layer0_outputs(76) <= inputs(204);
    layer0_outputs(77) <= (inputs(187)) or (inputs(71));
    layer0_outputs(78) <= (inputs(247)) xor (inputs(135));
    layer0_outputs(79) <= not(inputs(221)) or (inputs(145));
    layer0_outputs(80) <= not(inputs(20)) or (inputs(251));
    layer0_outputs(81) <= (inputs(62)) and not (inputs(138));
    layer0_outputs(82) <= (inputs(17)) xor (inputs(225));
    layer0_outputs(83) <= (inputs(176)) and (inputs(12));
    layer0_outputs(84) <= '0';
    layer0_outputs(85) <= not((inputs(156)) or (inputs(184)));
    layer0_outputs(86) <= not(inputs(201)) or (inputs(249));
    layer0_outputs(87) <= (inputs(149)) and not (inputs(8));
    layer0_outputs(88) <= not((inputs(201)) or (inputs(110)));
    layer0_outputs(89) <= '0';
    layer0_outputs(90) <= (inputs(33)) or (inputs(35));
    layer0_outputs(91) <= not(inputs(138)) or (inputs(78));
    layer0_outputs(92) <= inputs(201);
    layer0_outputs(93) <= inputs(127);
    layer0_outputs(94) <= (inputs(178)) and (inputs(246));
    layer0_outputs(95) <= (inputs(111)) and not (inputs(16));
    layer0_outputs(96) <= not((inputs(38)) or (inputs(186)));
    layer0_outputs(97) <= inputs(148);
    layer0_outputs(98) <= (inputs(30)) or (inputs(39));
    layer0_outputs(99) <= not((inputs(109)) xor (inputs(219)));
    layer0_outputs(100) <= (inputs(69)) and not (inputs(237));
    layer0_outputs(101) <= (inputs(168)) and (inputs(20));
    layer0_outputs(102) <= '1';
    layer0_outputs(103) <= inputs(25);
    layer0_outputs(104) <= not((inputs(12)) xor (inputs(202)));
    layer0_outputs(105) <= (inputs(221)) or (inputs(89));
    layer0_outputs(106) <= not(inputs(109));
    layer0_outputs(107) <= (inputs(200)) and not (inputs(205));
    layer0_outputs(108) <= not((inputs(114)) xor (inputs(224)));
    layer0_outputs(109) <= (inputs(162)) xor (inputs(213));
    layer0_outputs(110) <= not((inputs(108)) xor (inputs(92)));
    layer0_outputs(111) <= (inputs(83)) or (inputs(247));
    layer0_outputs(112) <= not(inputs(122));
    layer0_outputs(113) <= '1';
    layer0_outputs(114) <= not((inputs(62)) or (inputs(7)));
    layer0_outputs(115) <= (inputs(102)) and not (inputs(65));
    layer0_outputs(116) <= (inputs(7)) and (inputs(64));
    layer0_outputs(117) <= not(inputs(23));
    layer0_outputs(118) <= not(inputs(32)) or (inputs(169));
    layer0_outputs(119) <= inputs(65);
    layer0_outputs(120) <= (inputs(77)) and not (inputs(211));
    layer0_outputs(121) <= not(inputs(47));
    layer0_outputs(122) <= (inputs(216)) and not (inputs(35));
    layer0_outputs(123) <= (inputs(182)) and not (inputs(204));
    layer0_outputs(124) <= (inputs(140)) and not (inputs(26));
    layer0_outputs(125) <= not(inputs(241)) or (inputs(186));
    layer0_outputs(126) <= (inputs(170)) and not (inputs(185));
    layer0_outputs(127) <= not((inputs(197)) or (inputs(39)));
    layer0_outputs(128) <= not((inputs(218)) or (inputs(94)));
    layer0_outputs(129) <= (inputs(135)) xor (inputs(205));
    layer0_outputs(130) <= (inputs(221)) or (inputs(168));
    layer0_outputs(131) <= not(inputs(38));
    layer0_outputs(132) <= (inputs(163)) or (inputs(72));
    layer0_outputs(133) <= not(inputs(244));
    layer0_outputs(134) <= inputs(166);
    layer0_outputs(135) <= not((inputs(209)) xor (inputs(209)));
    layer0_outputs(136) <= not((inputs(32)) and (inputs(219)));
    layer0_outputs(137) <= not(inputs(56)) or (inputs(155));
    layer0_outputs(138) <= (inputs(212)) and not (inputs(173));
    layer0_outputs(139) <= inputs(165);
    layer0_outputs(140) <= inputs(176);
    layer0_outputs(141) <= not(inputs(53));
    layer0_outputs(142) <= (inputs(185)) and not (inputs(213));
    layer0_outputs(143) <= not((inputs(169)) xor (inputs(66)));
    layer0_outputs(144) <= not((inputs(205)) and (inputs(23)));
    layer0_outputs(145) <= '1';
    layer0_outputs(146) <= not(inputs(138));
    layer0_outputs(147) <= (inputs(62)) xor (inputs(29));
    layer0_outputs(148) <= (inputs(45)) xor (inputs(237));
    layer0_outputs(149) <= not(inputs(182));
    layer0_outputs(150) <= (inputs(107)) or (inputs(67));
    layer0_outputs(151) <= not((inputs(76)) or (inputs(58)));
    layer0_outputs(152) <= not((inputs(196)) or (inputs(173)));
    layer0_outputs(153) <= not(inputs(72));
    layer0_outputs(154) <= (inputs(199)) xor (inputs(241));
    layer0_outputs(155) <= inputs(199);
    layer0_outputs(156) <= not((inputs(68)) or (inputs(46)));
    layer0_outputs(157) <= not(inputs(89));
    layer0_outputs(158) <= (inputs(135)) and not (inputs(19));
    layer0_outputs(159) <= not(inputs(152));
    layer0_outputs(160) <= not((inputs(108)) or (inputs(14)));
    layer0_outputs(161) <= not((inputs(186)) xor (inputs(83)));
    layer0_outputs(162) <= inputs(77);
    layer0_outputs(163) <= inputs(72);
    layer0_outputs(164) <= not(inputs(59)) or (inputs(148));
    layer0_outputs(165) <= (inputs(146)) or (inputs(234));
    layer0_outputs(166) <= (inputs(31)) or (inputs(40));
    layer0_outputs(167) <= inputs(156);
    layer0_outputs(168) <= inputs(53);
    layer0_outputs(169) <= (inputs(88)) and not (inputs(0));
    layer0_outputs(170) <= '1';
    layer0_outputs(171) <= (inputs(191)) xor (inputs(140));
    layer0_outputs(172) <= not(inputs(214));
    layer0_outputs(173) <= inputs(101);
    layer0_outputs(174) <= (inputs(57)) or (inputs(117));
    layer0_outputs(175) <= inputs(111);
    layer0_outputs(176) <= (inputs(160)) xor (inputs(26));
    layer0_outputs(177) <= (inputs(31)) and (inputs(185));
    layer0_outputs(178) <= (inputs(1)) xor (inputs(121));
    layer0_outputs(179) <= inputs(5);
    layer0_outputs(180) <= inputs(26);
    layer0_outputs(181) <= not((inputs(32)) or (inputs(243)));
    layer0_outputs(182) <= not((inputs(0)) or (inputs(34)));
    layer0_outputs(183) <= (inputs(106)) or (inputs(165));
    layer0_outputs(184) <= not((inputs(1)) or (inputs(140)));
    layer0_outputs(185) <= inputs(104);
    layer0_outputs(186) <= not((inputs(182)) xor (inputs(97)));
    layer0_outputs(187) <= inputs(150);
    layer0_outputs(188) <= not(inputs(29)) or (inputs(131));
    layer0_outputs(189) <= inputs(231);
    layer0_outputs(190) <= not(inputs(181));
    layer0_outputs(191) <= (inputs(35)) xor (inputs(164));
    layer0_outputs(192) <= not((inputs(192)) and (inputs(249)));
    layer0_outputs(193) <= (inputs(15)) xor (inputs(6));
    layer0_outputs(194) <= not(inputs(116));
    layer0_outputs(195) <= inputs(214);
    layer0_outputs(196) <= (inputs(58)) and not (inputs(155));
    layer0_outputs(197) <= inputs(6);
    layer0_outputs(198) <= (inputs(76)) or (inputs(219));
    layer0_outputs(199) <= not(inputs(188));
    layer0_outputs(200) <= inputs(206);
    layer0_outputs(201) <= not(inputs(252)) or (inputs(48));
    layer0_outputs(202) <= (inputs(36)) or (inputs(195));
    layer0_outputs(203) <= (inputs(118)) and not (inputs(113));
    layer0_outputs(204) <= not(inputs(230)) or (inputs(119));
    layer0_outputs(205) <= not(inputs(103));
    layer0_outputs(206) <= inputs(62);
    layer0_outputs(207) <= (inputs(31)) xor (inputs(104));
    layer0_outputs(208) <= (inputs(20)) xor (inputs(57));
    layer0_outputs(209) <= (inputs(17)) and not (inputs(244));
    layer0_outputs(210) <= (inputs(64)) and not (inputs(239));
    layer0_outputs(211) <= (inputs(154)) or (inputs(21));
    layer0_outputs(212) <= not(inputs(116));
    layer0_outputs(213) <= inputs(4);
    layer0_outputs(214) <= '1';
    layer0_outputs(215) <= '1';
    layer0_outputs(216) <= (inputs(92)) and not (inputs(34));
    layer0_outputs(217) <= not(inputs(198)) or (inputs(49));
    layer0_outputs(218) <= inputs(18);
    layer0_outputs(219) <= (inputs(19)) or (inputs(201));
    layer0_outputs(220) <= not((inputs(47)) or (inputs(58)));
    layer0_outputs(221) <= inputs(2);
    layer0_outputs(222) <= (inputs(2)) and (inputs(47));
    layer0_outputs(223) <= (inputs(182)) xor (inputs(195));
    layer0_outputs(224) <= inputs(154);
    layer0_outputs(225) <= (inputs(210)) and not (inputs(146));
    layer0_outputs(226) <= (inputs(179)) and not (inputs(247));
    layer0_outputs(227) <= not((inputs(58)) or (inputs(59)));
    layer0_outputs(228) <= not((inputs(132)) or (inputs(190)));
    layer0_outputs(229) <= not((inputs(172)) xor (inputs(218)));
    layer0_outputs(230) <= '0';
    layer0_outputs(231) <= (inputs(166)) or (inputs(41));
    layer0_outputs(232) <= not(inputs(187));
    layer0_outputs(233) <= '0';
    layer0_outputs(234) <= (inputs(91)) or (inputs(154));
    layer0_outputs(235) <= inputs(211);
    layer0_outputs(236) <= (inputs(217)) and not (inputs(120));
    layer0_outputs(237) <= '0';
    layer0_outputs(238) <= not(inputs(67)) or (inputs(220));
    layer0_outputs(239) <= (inputs(202)) xor (inputs(103));
    layer0_outputs(240) <= (inputs(108)) xor (inputs(31));
    layer0_outputs(241) <= not(inputs(15)) or (inputs(143));
    layer0_outputs(242) <= not(inputs(45)) or (inputs(95));
    layer0_outputs(243) <= not(inputs(121));
    layer0_outputs(244) <= '1';
    layer0_outputs(245) <= '0';
    layer0_outputs(246) <= inputs(60);
    layer0_outputs(247) <= inputs(88);
    layer0_outputs(248) <= (inputs(111)) or (inputs(22));
    layer0_outputs(249) <= (inputs(248)) and not (inputs(253));
    layer0_outputs(250) <= not((inputs(73)) or (inputs(189)));
    layer0_outputs(251) <= '1';
    layer0_outputs(252) <= (inputs(73)) and (inputs(6));
    layer0_outputs(253) <= '0';
    layer0_outputs(254) <= not((inputs(167)) or (inputs(198)));
    layer0_outputs(255) <= inputs(102);
    layer0_outputs(256) <= (inputs(10)) or (inputs(49));
    layer0_outputs(257) <= not((inputs(121)) or (inputs(180)));
    layer0_outputs(258) <= not(inputs(120)) or (inputs(155));
    layer0_outputs(259) <= not(inputs(19));
    layer0_outputs(260) <= inputs(20);
    layer0_outputs(261) <= '1';
    layer0_outputs(262) <= not((inputs(102)) or (inputs(85)));
    layer0_outputs(263) <= (inputs(9)) or (inputs(85));
    layer0_outputs(264) <= not((inputs(184)) or (inputs(80)));
    layer0_outputs(265) <= not(inputs(224));
    layer0_outputs(266) <= not(inputs(76)) or (inputs(247));
    layer0_outputs(267) <= (inputs(243)) or (inputs(206));
    layer0_outputs(268) <= (inputs(205)) xor (inputs(133));
    layer0_outputs(269) <= not(inputs(5)) or (inputs(243));
    layer0_outputs(270) <= '1';
    layer0_outputs(271) <= not(inputs(182));
    layer0_outputs(272) <= (inputs(68)) or (inputs(191));
    layer0_outputs(273) <= (inputs(227)) or (inputs(128));
    layer0_outputs(274) <= '1';
    layer0_outputs(275) <= inputs(212);
    layer0_outputs(276) <= (inputs(119)) xor (inputs(8));
    layer0_outputs(277) <= not((inputs(65)) xor (inputs(252)));
    layer0_outputs(278) <= not(inputs(78)) or (inputs(145));
    layer0_outputs(279) <= (inputs(223)) xor (inputs(200));
    layer0_outputs(280) <= inputs(156);
    layer0_outputs(281) <= not((inputs(167)) or (inputs(142)));
    layer0_outputs(282) <= (inputs(118)) xor (inputs(202));
    layer0_outputs(283) <= (inputs(14)) or (inputs(113));
    layer0_outputs(284) <= not(inputs(159)) or (inputs(152));
    layer0_outputs(285) <= inputs(3);
    layer0_outputs(286) <= (inputs(121)) and not (inputs(228));
    layer0_outputs(287) <= not(inputs(148));
    layer0_outputs(288) <= inputs(243);
    layer0_outputs(289) <= not(inputs(96));
    layer0_outputs(290) <= not((inputs(52)) or (inputs(214)));
    layer0_outputs(291) <= inputs(196);
    layer0_outputs(292) <= not((inputs(90)) xor (inputs(47)));
    layer0_outputs(293) <= not((inputs(133)) xor (inputs(129)));
    layer0_outputs(294) <= (inputs(26)) or (inputs(133));
    layer0_outputs(295) <= not(inputs(140));
    layer0_outputs(296) <= '1';
    layer0_outputs(297) <= (inputs(63)) or (inputs(114));
    layer0_outputs(298) <= inputs(197);
    layer0_outputs(299) <= inputs(47);
    layer0_outputs(300) <= (inputs(228)) xor (inputs(70));
    layer0_outputs(301) <= (inputs(145)) and not (inputs(9));
    layer0_outputs(302) <= not(inputs(28)) or (inputs(38));
    layer0_outputs(303) <= (inputs(208)) xor (inputs(180));
    layer0_outputs(304) <= (inputs(164)) or (inputs(147));
    layer0_outputs(305) <= '0';
    layer0_outputs(306) <= (inputs(236)) or (inputs(81));
    layer0_outputs(307) <= not(inputs(148));
    layer0_outputs(308) <= not(inputs(192));
    layer0_outputs(309) <= '0';
    layer0_outputs(310) <= (inputs(162)) and not (inputs(24));
    layer0_outputs(311) <= (inputs(20)) or (inputs(21));
    layer0_outputs(312) <= not((inputs(150)) or (inputs(91)));
    layer0_outputs(313) <= not(inputs(204));
    layer0_outputs(314) <= not(inputs(105)) or (inputs(23));
    layer0_outputs(315) <= not(inputs(177));
    layer0_outputs(316) <= inputs(26);
    layer0_outputs(317) <= (inputs(16)) or (inputs(5));
    layer0_outputs(318) <= not((inputs(153)) and (inputs(229)));
    layer0_outputs(319) <= inputs(204);
    layer0_outputs(320) <= not(inputs(68));
    layer0_outputs(321) <= not(inputs(5)) or (inputs(88));
    layer0_outputs(322) <= (inputs(171)) xor (inputs(137));
    layer0_outputs(323) <= (inputs(195)) and not (inputs(240));
    layer0_outputs(324) <= (inputs(13)) or (inputs(145));
    layer0_outputs(325) <= not((inputs(51)) or (inputs(29)));
    layer0_outputs(326) <= inputs(148);
    layer0_outputs(327) <= not((inputs(10)) or (inputs(117)));
    layer0_outputs(328) <= not((inputs(174)) and (inputs(125)));
    layer0_outputs(329) <= (inputs(58)) or (inputs(156));
    layer0_outputs(330) <= (inputs(184)) or (inputs(158));
    layer0_outputs(331) <= (inputs(53)) or (inputs(203));
    layer0_outputs(332) <= inputs(152);
    layer0_outputs(333) <= not((inputs(154)) xor (inputs(235)));
    layer0_outputs(334) <= not((inputs(218)) and (inputs(225)));
    layer0_outputs(335) <= inputs(102);
    layer0_outputs(336) <= not((inputs(146)) xor (inputs(157)));
    layer0_outputs(337) <= not((inputs(123)) xor (inputs(143)));
    layer0_outputs(338) <= not(inputs(69)) or (inputs(115));
    layer0_outputs(339) <= not((inputs(115)) or (inputs(201)));
    layer0_outputs(340) <= not(inputs(15));
    layer0_outputs(341) <= not((inputs(219)) or (inputs(72)));
    layer0_outputs(342) <= not(inputs(0));
    layer0_outputs(343) <= inputs(55);
    layer0_outputs(344) <= inputs(133);
    layer0_outputs(345) <= not(inputs(83)) or (inputs(60));
    layer0_outputs(346) <= '0';
    layer0_outputs(347) <= not(inputs(174));
    layer0_outputs(348) <= (inputs(240)) xor (inputs(61));
    layer0_outputs(349) <= not(inputs(60));
    layer0_outputs(350) <= (inputs(117)) or (inputs(28));
    layer0_outputs(351) <= not((inputs(76)) or (inputs(122)));
    layer0_outputs(352) <= '1';
    layer0_outputs(353) <= not(inputs(118));
    layer0_outputs(354) <= not((inputs(162)) or (inputs(172)));
    layer0_outputs(355) <= (inputs(83)) and (inputs(37));
    layer0_outputs(356) <= not(inputs(241)) or (inputs(210));
    layer0_outputs(357) <= not(inputs(54)) or (inputs(44));
    layer0_outputs(358) <= not(inputs(182));
    layer0_outputs(359) <= not(inputs(19)) or (inputs(7));
    layer0_outputs(360) <= inputs(122);
    layer0_outputs(361) <= not(inputs(198)) or (inputs(53));
    layer0_outputs(362) <= (inputs(13)) and not (inputs(208));
    layer0_outputs(363) <= inputs(133);
    layer0_outputs(364) <= inputs(137);
    layer0_outputs(365) <= (inputs(135)) or (inputs(191));
    layer0_outputs(366) <= not((inputs(79)) xor (inputs(63)));
    layer0_outputs(367) <= (inputs(212)) xor (inputs(192));
    layer0_outputs(368) <= inputs(252);
    layer0_outputs(369) <= inputs(132);
    layer0_outputs(370) <= not(inputs(234));
    layer0_outputs(371) <= (inputs(160)) xor (inputs(47));
    layer0_outputs(372) <= not((inputs(132)) xor (inputs(222)));
    layer0_outputs(373) <= inputs(74);
    layer0_outputs(374) <= not(inputs(253)) or (inputs(26));
    layer0_outputs(375) <= not((inputs(171)) or (inputs(198)));
    layer0_outputs(376) <= '1';
    layer0_outputs(377) <= not((inputs(172)) or (inputs(116)));
    layer0_outputs(378) <= not((inputs(242)) xor (inputs(43)));
    layer0_outputs(379) <= not((inputs(155)) xor (inputs(31)));
    layer0_outputs(380) <= (inputs(74)) or (inputs(231));
    layer0_outputs(381) <= not(inputs(100)) or (inputs(33));
    layer0_outputs(382) <= (inputs(104)) or (inputs(255));
    layer0_outputs(383) <= (inputs(157)) and not (inputs(218));
    layer0_outputs(384) <= not((inputs(225)) xor (inputs(205)));
    layer0_outputs(385) <= not(inputs(166)) or (inputs(223));
    layer0_outputs(386) <= (inputs(92)) and not (inputs(237));
    layer0_outputs(387) <= not((inputs(87)) or (inputs(15)));
    layer0_outputs(388) <= inputs(135);
    layer0_outputs(389) <= not((inputs(156)) xor (inputs(207)));
    layer0_outputs(390) <= not(inputs(73)) or (inputs(26));
    layer0_outputs(391) <= not(inputs(89));
    layer0_outputs(392) <= (inputs(118)) and not (inputs(21));
    layer0_outputs(393) <= (inputs(54)) and not (inputs(45));
    layer0_outputs(394) <= inputs(45);
    layer0_outputs(395) <= (inputs(86)) xor (inputs(109));
    layer0_outputs(396) <= (inputs(255)) or (inputs(181));
    layer0_outputs(397) <= not((inputs(164)) xor (inputs(7)));
    layer0_outputs(398) <= (inputs(153)) and (inputs(203));
    layer0_outputs(399) <= not(inputs(127));
    layer0_outputs(400) <= '0';
    layer0_outputs(401) <= not(inputs(121)) or (inputs(163));
    layer0_outputs(402) <= not((inputs(234)) xor (inputs(222)));
    layer0_outputs(403) <= inputs(138);
    layer0_outputs(404) <= inputs(137);
    layer0_outputs(405) <= (inputs(210)) and not (inputs(83));
    layer0_outputs(406) <= not(inputs(229)) or (inputs(68));
    layer0_outputs(407) <= not(inputs(19));
    layer0_outputs(408) <= (inputs(125)) xor (inputs(70));
    layer0_outputs(409) <= '1';
    layer0_outputs(410) <= (inputs(188)) xor (inputs(140));
    layer0_outputs(411) <= not(inputs(70)) or (inputs(171));
    layer0_outputs(412) <= not((inputs(221)) or (inputs(117)));
    layer0_outputs(413) <= not((inputs(93)) xor (inputs(105)));
    layer0_outputs(414) <= not(inputs(213));
    layer0_outputs(415) <= '0';
    layer0_outputs(416) <= inputs(13);
    layer0_outputs(417) <= (inputs(179)) or (inputs(194));
    layer0_outputs(418) <= (inputs(100)) or (inputs(187));
    layer0_outputs(419) <= not(inputs(172));
    layer0_outputs(420) <= not((inputs(123)) xor (inputs(99)));
    layer0_outputs(421) <= (inputs(55)) and not (inputs(130));
    layer0_outputs(422) <= (inputs(187)) and not (inputs(23));
    layer0_outputs(423) <= (inputs(212)) and not (inputs(192));
    layer0_outputs(424) <= not((inputs(96)) or (inputs(69)));
    layer0_outputs(425) <= not((inputs(157)) and (inputs(18)));
    layer0_outputs(426) <= not(inputs(104)) or (inputs(129));
    layer0_outputs(427) <= (inputs(66)) xor (inputs(24));
    layer0_outputs(428) <= not((inputs(76)) or (inputs(93)));
    layer0_outputs(429) <= inputs(86);
    layer0_outputs(430) <= (inputs(74)) or (inputs(227));
    layer0_outputs(431) <= not(inputs(126)) or (inputs(237));
    layer0_outputs(432) <= not(inputs(153)) or (inputs(180));
    layer0_outputs(433) <= (inputs(206)) or (inputs(248));
    layer0_outputs(434) <= (inputs(57)) and (inputs(96));
    layer0_outputs(435) <= not((inputs(42)) or (inputs(83)));
    layer0_outputs(436) <= (inputs(43)) and not (inputs(116));
    layer0_outputs(437) <= not(inputs(16)) or (inputs(109));
    layer0_outputs(438) <= (inputs(251)) xor (inputs(214));
    layer0_outputs(439) <= (inputs(245)) xor (inputs(226));
    layer0_outputs(440) <= inputs(32);
    layer0_outputs(441) <= not(inputs(133)) or (inputs(11));
    layer0_outputs(442) <= not((inputs(168)) or (inputs(247)));
    layer0_outputs(443) <= not((inputs(50)) or (inputs(161)));
    layer0_outputs(444) <= (inputs(103)) and not (inputs(231));
    layer0_outputs(445) <= inputs(183);
    layer0_outputs(446) <= (inputs(62)) and not (inputs(20));
    layer0_outputs(447) <= not(inputs(69));
    layer0_outputs(448) <= not(inputs(11)) or (inputs(85));
    layer0_outputs(449) <= inputs(18);
    layer0_outputs(450) <= (inputs(109)) and (inputs(251));
    layer0_outputs(451) <= (inputs(49)) xor (inputs(122));
    layer0_outputs(452) <= (inputs(243)) and not (inputs(126));
    layer0_outputs(453) <= not((inputs(143)) xor (inputs(15)));
    layer0_outputs(454) <= not(inputs(1)) or (inputs(176));
    layer0_outputs(455) <= (inputs(230)) and not (inputs(38));
    layer0_outputs(456) <= inputs(109);
    layer0_outputs(457) <= inputs(237);
    layer0_outputs(458) <= (inputs(165)) and not (inputs(146));
    layer0_outputs(459) <= not((inputs(227)) or (inputs(78)));
    layer0_outputs(460) <= (inputs(215)) or (inputs(123));
    layer0_outputs(461) <= (inputs(206)) and not (inputs(97));
    layer0_outputs(462) <= not((inputs(216)) or (inputs(224)));
    layer0_outputs(463) <= '1';
    layer0_outputs(464) <= not((inputs(135)) or (inputs(43)));
    layer0_outputs(465) <= not(inputs(196)) or (inputs(251));
    layer0_outputs(466) <= not((inputs(88)) or (inputs(148)));
    layer0_outputs(467) <= (inputs(191)) or (inputs(160));
    layer0_outputs(468) <= not(inputs(187));
    layer0_outputs(469) <= (inputs(113)) and (inputs(151));
    layer0_outputs(470) <= '1';
    layer0_outputs(471) <= not(inputs(250));
    layer0_outputs(472) <= (inputs(158)) xor (inputs(91));
    layer0_outputs(473) <= (inputs(197)) and not (inputs(27));
    layer0_outputs(474) <= inputs(213);
    layer0_outputs(475) <= not(inputs(230)) or (inputs(42));
    layer0_outputs(476) <= (inputs(161)) and not (inputs(158));
    layer0_outputs(477) <= not((inputs(204)) or (inputs(150)));
    layer0_outputs(478) <= inputs(56);
    layer0_outputs(479) <= not(inputs(84)) or (inputs(202));
    layer0_outputs(480) <= inputs(187);
    layer0_outputs(481) <= (inputs(231)) and (inputs(69));
    layer0_outputs(482) <= not((inputs(153)) or (inputs(190)));
    layer0_outputs(483) <= not((inputs(157)) xor (inputs(238)));
    layer0_outputs(484) <= (inputs(19)) and (inputs(162));
    layer0_outputs(485) <= (inputs(83)) xor (inputs(224));
    layer0_outputs(486) <= not(inputs(120));
    layer0_outputs(487) <= (inputs(140)) and not (inputs(139));
    layer0_outputs(488) <= not((inputs(125)) or (inputs(86)));
    layer0_outputs(489) <= not(inputs(87)) or (inputs(157));
    layer0_outputs(490) <= not(inputs(227)) or (inputs(222));
    layer0_outputs(491) <= not((inputs(9)) or (inputs(137)));
    layer0_outputs(492) <= inputs(45);
    layer0_outputs(493) <= (inputs(158)) xor (inputs(233));
    layer0_outputs(494) <= inputs(149);
    layer0_outputs(495) <= inputs(125);
    layer0_outputs(496) <= (inputs(178)) and not (inputs(78));
    layer0_outputs(497) <= not(inputs(144)) or (inputs(6));
    layer0_outputs(498) <= (inputs(147)) and not (inputs(39));
    layer0_outputs(499) <= '1';
    layer0_outputs(500) <= not(inputs(196)) or (inputs(234));
    layer0_outputs(501) <= not((inputs(25)) xor (inputs(158)));
    layer0_outputs(502) <= (inputs(208)) and not (inputs(156));
    layer0_outputs(503) <= not((inputs(179)) or (inputs(158)));
    layer0_outputs(504) <= not(inputs(50)) or (inputs(90));
    layer0_outputs(505) <= not((inputs(106)) xor (inputs(12)));
    layer0_outputs(506) <= (inputs(225)) xor (inputs(187));
    layer0_outputs(507) <= inputs(54);
    layer0_outputs(508) <= not(inputs(206)) or (inputs(83));
    layer0_outputs(509) <= inputs(180);
    layer0_outputs(510) <= not((inputs(37)) and (inputs(13)));
    layer0_outputs(511) <= (inputs(3)) and not (inputs(33));
    layer0_outputs(512) <= (inputs(233)) and (inputs(98));
    layer0_outputs(513) <= (inputs(191)) xor (inputs(97));
    layer0_outputs(514) <= inputs(76);
    layer0_outputs(515) <= inputs(109);
    layer0_outputs(516) <= not((inputs(93)) or (inputs(8)));
    layer0_outputs(517) <= (inputs(52)) or (inputs(196));
    layer0_outputs(518) <= inputs(149);
    layer0_outputs(519) <= not(inputs(184)) or (inputs(6));
    layer0_outputs(520) <= (inputs(200)) and not (inputs(139));
    layer0_outputs(521) <= not(inputs(119)) or (inputs(105));
    layer0_outputs(522) <= (inputs(232)) and not (inputs(30));
    layer0_outputs(523) <= inputs(56);
    layer0_outputs(524) <= inputs(112);
    layer0_outputs(525) <= (inputs(252)) xor (inputs(251));
    layer0_outputs(526) <= '1';
    layer0_outputs(527) <= inputs(120);
    layer0_outputs(528) <= (inputs(14)) and (inputs(68));
    layer0_outputs(529) <= not((inputs(35)) xor (inputs(150)));
    layer0_outputs(530) <= (inputs(91)) xor (inputs(167));
    layer0_outputs(531) <= inputs(186);
    layer0_outputs(532) <= not((inputs(163)) or (inputs(109)));
    layer0_outputs(533) <= not((inputs(201)) or (inputs(240)));
    layer0_outputs(534) <= inputs(120);
    layer0_outputs(535) <= (inputs(110)) and (inputs(223));
    layer0_outputs(536) <= not((inputs(151)) or (inputs(194)));
    layer0_outputs(537) <= not(inputs(133));
    layer0_outputs(538) <= inputs(101);
    layer0_outputs(539) <= not(inputs(119));
    layer0_outputs(540) <= (inputs(21)) xor (inputs(248));
    layer0_outputs(541) <= not(inputs(78));
    layer0_outputs(542) <= '1';
    layer0_outputs(543) <= not((inputs(121)) and (inputs(208)));
    layer0_outputs(544) <= not(inputs(189)) or (inputs(79));
    layer0_outputs(545) <= (inputs(91)) and not (inputs(43));
    layer0_outputs(546) <= not(inputs(184));
    layer0_outputs(547) <= not(inputs(252));
    layer0_outputs(548) <= not((inputs(66)) or (inputs(87)));
    layer0_outputs(549) <= not((inputs(13)) xor (inputs(159)));
    layer0_outputs(550) <= not((inputs(201)) xor (inputs(141)));
    layer0_outputs(551) <= not((inputs(74)) or (inputs(76)));
    layer0_outputs(552) <= inputs(42);
    layer0_outputs(553) <= inputs(132);
    layer0_outputs(554) <= inputs(124);
    layer0_outputs(555) <= '1';
    layer0_outputs(556) <= not(inputs(223)) or (inputs(128));
    layer0_outputs(557) <= not(inputs(53)) or (inputs(46));
    layer0_outputs(558) <= inputs(182);
    layer0_outputs(559) <= (inputs(28)) and (inputs(43));
    layer0_outputs(560) <= '1';
    layer0_outputs(561) <= inputs(101);
    layer0_outputs(562) <= (inputs(141)) or (inputs(123));
    layer0_outputs(563) <= (inputs(87)) xor (inputs(39));
    layer0_outputs(564) <= not(inputs(3)) or (inputs(92));
    layer0_outputs(565) <= not((inputs(248)) or (inputs(127)));
    layer0_outputs(566) <= (inputs(180)) or (inputs(77));
    layer0_outputs(567) <= (inputs(68)) and not (inputs(167));
    layer0_outputs(568) <= inputs(213);
    layer0_outputs(569) <= not(inputs(53));
    layer0_outputs(570) <= '1';
    layer0_outputs(571) <= not((inputs(214)) or (inputs(80)));
    layer0_outputs(572) <= (inputs(45)) or (inputs(23));
    layer0_outputs(573) <= not(inputs(39)) or (inputs(235));
    layer0_outputs(574) <= inputs(61);
    layer0_outputs(575) <= not(inputs(217)) or (inputs(108));
    layer0_outputs(576) <= '0';
    layer0_outputs(577) <= inputs(56);
    layer0_outputs(578) <= (inputs(52)) or (inputs(35));
    layer0_outputs(579) <= not(inputs(240));
    layer0_outputs(580) <= not(inputs(121));
    layer0_outputs(581) <= inputs(195);
    layer0_outputs(582) <= not(inputs(148)) or (inputs(27));
    layer0_outputs(583) <= inputs(104);
    layer0_outputs(584) <= (inputs(155)) xor (inputs(160));
    layer0_outputs(585) <= (inputs(173)) xor (inputs(62));
    layer0_outputs(586) <= (inputs(121)) and not (inputs(219));
    layer0_outputs(587) <= not(inputs(49));
    layer0_outputs(588) <= not(inputs(84));
    layer0_outputs(589) <= (inputs(219)) or (inputs(17));
    layer0_outputs(590) <= '1';
    layer0_outputs(591) <= not((inputs(124)) or (inputs(194)));
    layer0_outputs(592) <= not(inputs(173));
    layer0_outputs(593) <= not(inputs(57)) or (inputs(61));
    layer0_outputs(594) <= not((inputs(89)) xor (inputs(15)));
    layer0_outputs(595) <= '0';
    layer0_outputs(596) <= not((inputs(74)) xor (inputs(6)));
    layer0_outputs(597) <= inputs(170);
    layer0_outputs(598) <= (inputs(196)) and not (inputs(91));
    layer0_outputs(599) <= not(inputs(104)) or (inputs(241));
    layer0_outputs(600) <= not(inputs(102)) or (inputs(6));
    layer0_outputs(601) <= not((inputs(174)) and (inputs(236)));
    layer0_outputs(602) <= (inputs(211)) and not (inputs(126));
    layer0_outputs(603) <= not((inputs(53)) or (inputs(61)));
    layer0_outputs(604) <= (inputs(31)) and (inputs(178));
    layer0_outputs(605) <= not((inputs(222)) or (inputs(7)));
    layer0_outputs(606) <= (inputs(247)) and (inputs(12));
    layer0_outputs(607) <= not((inputs(213)) xor (inputs(95)));
    layer0_outputs(608) <= not(inputs(230));
    layer0_outputs(609) <= not((inputs(10)) or (inputs(132)));
    layer0_outputs(610) <= not(inputs(163)) or (inputs(226));
    layer0_outputs(611) <= not((inputs(110)) or (inputs(214)));
    layer0_outputs(612) <= (inputs(5)) and not (inputs(66));
    layer0_outputs(613) <= (inputs(34)) xor (inputs(185));
    layer0_outputs(614) <= (inputs(206)) and not (inputs(176));
    layer0_outputs(615) <= (inputs(77)) and not (inputs(208));
    layer0_outputs(616) <= (inputs(151)) and not (inputs(81));
    layer0_outputs(617) <= (inputs(76)) and not (inputs(97));
    layer0_outputs(618) <= (inputs(242)) and (inputs(28));
    layer0_outputs(619) <= inputs(189);
    layer0_outputs(620) <= not(inputs(147));
    layer0_outputs(621) <= not((inputs(93)) or (inputs(91)));
    layer0_outputs(622) <= inputs(25);
    layer0_outputs(623) <= (inputs(68)) xor (inputs(41));
    layer0_outputs(624) <= (inputs(100)) and (inputs(99));
    layer0_outputs(625) <= not(inputs(131)) or (inputs(96));
    layer0_outputs(626) <= '0';
    layer0_outputs(627) <= not(inputs(51));
    layer0_outputs(628) <= (inputs(5)) and (inputs(156));
    layer0_outputs(629) <= not(inputs(158)) or (inputs(121));
    layer0_outputs(630) <= not(inputs(108));
    layer0_outputs(631) <= not((inputs(158)) or (inputs(228)));
    layer0_outputs(632) <= not((inputs(51)) xor (inputs(29)));
    layer0_outputs(633) <= '0';
    layer0_outputs(634) <= not(inputs(211)) or (inputs(49));
    layer0_outputs(635) <= not(inputs(122));
    layer0_outputs(636) <= not(inputs(38));
    layer0_outputs(637) <= not((inputs(39)) or (inputs(157)));
    layer0_outputs(638) <= not((inputs(156)) or (inputs(43)));
    layer0_outputs(639) <= not(inputs(106));
    layer0_outputs(640) <= not((inputs(11)) xor (inputs(187)));
    layer0_outputs(641) <= (inputs(121)) and not (inputs(41));
    layer0_outputs(642) <= not((inputs(176)) xor (inputs(148)));
    layer0_outputs(643) <= (inputs(29)) and not (inputs(75));
    layer0_outputs(644) <= not((inputs(93)) or (inputs(33)));
    layer0_outputs(645) <= not(inputs(118)) or (inputs(97));
    layer0_outputs(646) <= not(inputs(185)) or (inputs(0));
    layer0_outputs(647) <= inputs(228);
    layer0_outputs(648) <= (inputs(37)) or (inputs(103));
    layer0_outputs(649) <= not(inputs(177));
    layer0_outputs(650) <= (inputs(134)) or (inputs(234));
    layer0_outputs(651) <= not(inputs(85)) or (inputs(39));
    layer0_outputs(652) <= (inputs(111)) xor (inputs(137));
    layer0_outputs(653) <= '1';
    layer0_outputs(654) <= not((inputs(125)) and (inputs(159)));
    layer0_outputs(655) <= not(inputs(133));
    layer0_outputs(656) <= (inputs(57)) and not (inputs(140));
    layer0_outputs(657) <= (inputs(73)) or (inputs(176));
    layer0_outputs(658) <= not((inputs(252)) xor (inputs(172)));
    layer0_outputs(659) <= not(inputs(108));
    layer0_outputs(660) <= '0';
    layer0_outputs(661) <= not(inputs(187)) or (inputs(99));
    layer0_outputs(662) <= (inputs(184)) xor (inputs(82));
    layer0_outputs(663) <= inputs(56);
    layer0_outputs(664) <= inputs(138);
    layer0_outputs(665) <= not(inputs(223)) or (inputs(30));
    layer0_outputs(666) <= not(inputs(77)) or (inputs(65));
    layer0_outputs(667) <= inputs(36);
    layer0_outputs(668) <= (inputs(34)) or (inputs(171));
    layer0_outputs(669) <= not((inputs(186)) xor (inputs(8)));
    layer0_outputs(670) <= not((inputs(136)) or (inputs(39)));
    layer0_outputs(671) <= (inputs(203)) and (inputs(127));
    layer0_outputs(672) <= not((inputs(130)) or (inputs(149)));
    layer0_outputs(673) <= '0';
    layer0_outputs(674) <= not(inputs(30)) or (inputs(243));
    layer0_outputs(675) <= not(inputs(212));
    layer0_outputs(676) <= (inputs(179)) and not (inputs(131));
    layer0_outputs(677) <= inputs(236);
    layer0_outputs(678) <= not(inputs(35));
    layer0_outputs(679) <= (inputs(116)) or (inputs(76));
    layer0_outputs(680) <= not(inputs(49)) or (inputs(172));
    layer0_outputs(681) <= not(inputs(90));
    layer0_outputs(682) <= (inputs(121)) and not (inputs(122));
    layer0_outputs(683) <= inputs(125);
    layer0_outputs(684) <= not(inputs(68));
    layer0_outputs(685) <= (inputs(233)) and not (inputs(145));
    layer0_outputs(686) <= (inputs(137)) or (inputs(147));
    layer0_outputs(687) <= (inputs(48)) and not (inputs(76));
    layer0_outputs(688) <= not(inputs(55));
    layer0_outputs(689) <= not((inputs(24)) and (inputs(233)));
    layer0_outputs(690) <= not(inputs(1)) or (inputs(176));
    layer0_outputs(691) <= (inputs(193)) and not (inputs(48));
    layer0_outputs(692) <= not(inputs(184));
    layer0_outputs(693) <= (inputs(33)) or (inputs(236));
    layer0_outputs(694) <= not((inputs(89)) or (inputs(234)));
    layer0_outputs(695) <= (inputs(93)) and not (inputs(239));
    layer0_outputs(696) <= not((inputs(192)) and (inputs(130)));
    layer0_outputs(697) <= (inputs(181)) and (inputs(223));
    layer0_outputs(698) <= inputs(217);
    layer0_outputs(699) <= not(inputs(217)) or (inputs(123));
    layer0_outputs(700) <= not((inputs(108)) or (inputs(236)));
    layer0_outputs(701) <= inputs(55);
    layer0_outputs(702) <= '1';
    layer0_outputs(703) <= not(inputs(175));
    layer0_outputs(704) <= not(inputs(33)) or (inputs(90));
    layer0_outputs(705) <= not(inputs(251));
    layer0_outputs(706) <= not((inputs(175)) xor (inputs(65)));
    layer0_outputs(707) <= (inputs(139)) and not (inputs(51));
    layer0_outputs(708) <= not(inputs(55)) or (inputs(139));
    layer0_outputs(709) <= not(inputs(39));
    layer0_outputs(710) <= (inputs(78)) and not (inputs(60));
    layer0_outputs(711) <= not(inputs(25)) or (inputs(228));
    layer0_outputs(712) <= not((inputs(182)) xor (inputs(239)));
    layer0_outputs(713) <= not(inputs(57));
    layer0_outputs(714) <= not((inputs(204)) or (inputs(38)));
    layer0_outputs(715) <= not(inputs(104)) or (inputs(235));
    layer0_outputs(716) <= not((inputs(88)) xor (inputs(74)));
    layer0_outputs(717) <= (inputs(223)) and not (inputs(252));
    layer0_outputs(718) <= not((inputs(197)) or (inputs(215)));
    layer0_outputs(719) <= not((inputs(205)) or (inputs(54)));
    layer0_outputs(720) <= not((inputs(74)) and (inputs(217)));
    layer0_outputs(721) <= (inputs(8)) xor (inputs(69));
    layer0_outputs(722) <= (inputs(44)) and (inputs(247));
    layer0_outputs(723) <= inputs(180);
    layer0_outputs(724) <= (inputs(236)) xor (inputs(225));
    layer0_outputs(725) <= (inputs(45)) and (inputs(218));
    layer0_outputs(726) <= (inputs(152)) and not (inputs(7));
    layer0_outputs(727) <= inputs(133);
    layer0_outputs(728) <= (inputs(231)) and (inputs(213));
    layer0_outputs(729) <= not((inputs(13)) and (inputs(81)));
    layer0_outputs(730) <= '1';
    layer0_outputs(731) <= inputs(229);
    layer0_outputs(732) <= not((inputs(125)) or (inputs(72)));
    layer0_outputs(733) <= not(inputs(200)) or (inputs(128));
    layer0_outputs(734) <= (inputs(31)) xor (inputs(235));
    layer0_outputs(735) <= (inputs(123)) and not (inputs(161));
    layer0_outputs(736) <= inputs(132);
    layer0_outputs(737) <= (inputs(247)) and not (inputs(8));
    layer0_outputs(738) <= not((inputs(95)) or (inputs(62)));
    layer0_outputs(739) <= not(inputs(76)) or (inputs(145));
    layer0_outputs(740) <= not(inputs(203));
    layer0_outputs(741) <= not(inputs(181));
    layer0_outputs(742) <= '0';
    layer0_outputs(743) <= not(inputs(62));
    layer0_outputs(744) <= not((inputs(34)) or (inputs(42)));
    layer0_outputs(745) <= (inputs(68)) or (inputs(200));
    layer0_outputs(746) <= (inputs(249)) or (inputs(89));
    layer0_outputs(747) <= not((inputs(85)) or (inputs(12)));
    layer0_outputs(748) <= '0';
    layer0_outputs(749) <= not(inputs(72)) or (inputs(138));
    layer0_outputs(750) <= '1';
    layer0_outputs(751) <= (inputs(185)) or (inputs(60));
    layer0_outputs(752) <= (inputs(182)) xor (inputs(196));
    layer0_outputs(753) <= (inputs(55)) and not (inputs(210));
    layer0_outputs(754) <= (inputs(68)) and not (inputs(63));
    layer0_outputs(755) <= not((inputs(214)) or (inputs(125)));
    layer0_outputs(756) <= inputs(236);
    layer0_outputs(757) <= inputs(134);
    layer0_outputs(758) <= '1';
    layer0_outputs(759) <= not(inputs(105));
    layer0_outputs(760) <= (inputs(86)) and not (inputs(140));
    layer0_outputs(761) <= '0';
    layer0_outputs(762) <= not(inputs(215)) or (inputs(158));
    layer0_outputs(763) <= not((inputs(14)) and (inputs(32)));
    layer0_outputs(764) <= not((inputs(238)) and (inputs(18)));
    layer0_outputs(765) <= not(inputs(108)) or (inputs(205));
    layer0_outputs(766) <= (inputs(209)) or (inputs(113));
    layer0_outputs(767) <= not(inputs(186)) or (inputs(245));
    layer0_outputs(768) <= not(inputs(149)) or (inputs(114));
    layer0_outputs(769) <= not((inputs(170)) or (inputs(195)));
    layer0_outputs(770) <= not((inputs(250)) or (inputs(213)));
    layer0_outputs(771) <= (inputs(182)) and not (inputs(35));
    layer0_outputs(772) <= (inputs(42)) xor (inputs(187));
    layer0_outputs(773) <= inputs(179);
    layer0_outputs(774) <= not((inputs(250)) and (inputs(49)));
    layer0_outputs(775) <= not(inputs(206));
    layer0_outputs(776) <= inputs(56);
    layer0_outputs(777) <= (inputs(31)) or (inputs(58));
    layer0_outputs(778) <= not((inputs(31)) and (inputs(12)));
    layer0_outputs(779) <= not((inputs(176)) and (inputs(154)));
    layer0_outputs(780) <= (inputs(43)) and (inputs(8));
    layer0_outputs(781) <= (inputs(194)) or (inputs(70));
    layer0_outputs(782) <= (inputs(115)) or (inputs(19));
    layer0_outputs(783) <= not(inputs(175));
    layer0_outputs(784) <= not(inputs(202));
    layer0_outputs(785) <= not(inputs(168)) or (inputs(185));
    layer0_outputs(786) <= (inputs(80)) or (inputs(49));
    layer0_outputs(787) <= not(inputs(167));
    layer0_outputs(788) <= (inputs(243)) and not (inputs(44));
    layer0_outputs(789) <= (inputs(86)) and not (inputs(47));
    layer0_outputs(790) <= '1';
    layer0_outputs(791) <= not(inputs(152));
    layer0_outputs(792) <= not(inputs(102)) or (inputs(236));
    layer0_outputs(793) <= (inputs(23)) xor (inputs(49));
    layer0_outputs(794) <= not(inputs(143));
    layer0_outputs(795) <= not((inputs(156)) or (inputs(193)));
    layer0_outputs(796) <= not((inputs(142)) xor (inputs(8)));
    layer0_outputs(797) <= not(inputs(251)) or (inputs(34));
    layer0_outputs(798) <= not((inputs(200)) or (inputs(156)));
    layer0_outputs(799) <= not(inputs(180));
    layer0_outputs(800) <= not(inputs(158)) or (inputs(252));
    layer0_outputs(801) <= inputs(11);
    layer0_outputs(802) <= not((inputs(123)) xor (inputs(165)));
    layer0_outputs(803) <= (inputs(131)) or (inputs(164));
    layer0_outputs(804) <= (inputs(128)) and not (inputs(43));
    layer0_outputs(805) <= not((inputs(220)) or (inputs(80)));
    layer0_outputs(806) <= not(inputs(5)) or (inputs(104));
    layer0_outputs(807) <= (inputs(88)) xor (inputs(96));
    layer0_outputs(808) <= not((inputs(93)) or (inputs(119)));
    layer0_outputs(809) <= inputs(59);
    layer0_outputs(810) <= not((inputs(134)) xor (inputs(207)));
    layer0_outputs(811) <= not((inputs(41)) xor (inputs(219)));
    layer0_outputs(812) <= not((inputs(222)) and (inputs(191)));
    layer0_outputs(813) <= '1';
    layer0_outputs(814) <= (inputs(159)) and not (inputs(131));
    layer0_outputs(815) <= not((inputs(64)) or (inputs(171)));
    layer0_outputs(816) <= (inputs(135)) xor (inputs(105));
    layer0_outputs(817) <= inputs(214);
    layer0_outputs(818) <= (inputs(171)) and not (inputs(33));
    layer0_outputs(819) <= not(inputs(169));
    layer0_outputs(820) <= (inputs(113)) and not (inputs(60));
    layer0_outputs(821) <= inputs(36);
    layer0_outputs(822) <= not(inputs(80)) or (inputs(230));
    layer0_outputs(823) <= (inputs(150)) and not (inputs(175));
    layer0_outputs(824) <= not(inputs(139));
    layer0_outputs(825) <= (inputs(176)) xor (inputs(115));
    layer0_outputs(826) <= '0';
    layer0_outputs(827) <= inputs(23);
    layer0_outputs(828) <= inputs(203);
    layer0_outputs(829) <= not(inputs(201)) or (inputs(189));
    layer0_outputs(830) <= (inputs(32)) and not (inputs(154));
    layer0_outputs(831) <= (inputs(72)) and (inputs(7));
    layer0_outputs(832) <= not(inputs(50));
    layer0_outputs(833) <= not((inputs(64)) xor (inputs(123)));
    layer0_outputs(834) <= (inputs(135)) and not (inputs(104));
    layer0_outputs(835) <= (inputs(79)) xor (inputs(51));
    layer0_outputs(836) <= not(inputs(148)) or (inputs(186));
    layer0_outputs(837) <= (inputs(240)) and not (inputs(123));
    layer0_outputs(838) <= (inputs(30)) or (inputs(145));
    layer0_outputs(839) <= not(inputs(116));
    layer0_outputs(840) <= inputs(156);
    layer0_outputs(841) <= not(inputs(7));
    layer0_outputs(842) <= inputs(184);
    layer0_outputs(843) <= inputs(172);
    layer0_outputs(844) <= (inputs(38)) and (inputs(122));
    layer0_outputs(845) <= (inputs(73)) and not (inputs(141));
    layer0_outputs(846) <= (inputs(188)) or (inputs(60));
    layer0_outputs(847) <= not((inputs(220)) or (inputs(174)));
    layer0_outputs(848) <= not(inputs(205));
    layer0_outputs(849) <= not(inputs(126));
    layer0_outputs(850) <= not((inputs(190)) or (inputs(71)));
    layer0_outputs(851) <= (inputs(165)) or (inputs(67));
    layer0_outputs(852) <= not((inputs(242)) or (inputs(180)));
    layer0_outputs(853) <= (inputs(219)) or (inputs(116));
    layer0_outputs(854) <= inputs(224);
    layer0_outputs(855) <= not((inputs(189)) xor (inputs(179)));
    layer0_outputs(856) <= (inputs(73)) and not (inputs(24));
    layer0_outputs(857) <= not(inputs(214)) or (inputs(186));
    layer0_outputs(858) <= not((inputs(243)) or (inputs(155)));
    layer0_outputs(859) <= not(inputs(154));
    layer0_outputs(860) <= (inputs(59)) and (inputs(153));
    layer0_outputs(861) <= (inputs(241)) or (inputs(230));
    layer0_outputs(862) <= inputs(215);
    layer0_outputs(863) <= (inputs(252)) and (inputs(169));
    layer0_outputs(864) <= (inputs(90)) xor (inputs(35));
    layer0_outputs(865) <= '0';
    layer0_outputs(866) <= (inputs(208)) or (inputs(61));
    layer0_outputs(867) <= not(inputs(224));
    layer0_outputs(868) <= (inputs(221)) xor (inputs(109));
    layer0_outputs(869) <= not(inputs(179));
    layer0_outputs(870) <= not(inputs(78));
    layer0_outputs(871) <= (inputs(21)) or (inputs(207));
    layer0_outputs(872) <= not((inputs(25)) xor (inputs(178)));
    layer0_outputs(873) <= not(inputs(74));
    layer0_outputs(874) <= inputs(134);
    layer0_outputs(875) <= '0';
    layer0_outputs(876) <= inputs(21);
    layer0_outputs(877) <= (inputs(230)) and not (inputs(246));
    layer0_outputs(878) <= (inputs(52)) or (inputs(51));
    layer0_outputs(879) <= not((inputs(172)) and (inputs(188)));
    layer0_outputs(880) <= inputs(70);
    layer0_outputs(881) <= not(inputs(188)) or (inputs(253));
    layer0_outputs(882) <= '0';
    layer0_outputs(883) <= not((inputs(225)) or (inputs(164)));
    layer0_outputs(884) <= inputs(22);
    layer0_outputs(885) <= (inputs(123)) and not (inputs(211));
    layer0_outputs(886) <= not(inputs(54));
    layer0_outputs(887) <= (inputs(180)) xor (inputs(214));
    layer0_outputs(888) <= not((inputs(165)) or (inputs(39)));
    layer0_outputs(889) <= (inputs(199)) xor (inputs(4));
    layer0_outputs(890) <= not(inputs(148)) or (inputs(151));
    layer0_outputs(891) <= (inputs(156)) and not (inputs(208));
    layer0_outputs(892) <= not(inputs(90));
    layer0_outputs(893) <= (inputs(130)) or (inputs(99));
    layer0_outputs(894) <= (inputs(231)) or (inputs(139));
    layer0_outputs(895) <= inputs(57);
    layer0_outputs(896) <= (inputs(122)) and not (inputs(204));
    layer0_outputs(897) <= (inputs(13)) or (inputs(84));
    layer0_outputs(898) <= (inputs(121)) and not (inputs(49));
    layer0_outputs(899) <= not(inputs(169));
    layer0_outputs(900) <= inputs(211);
    layer0_outputs(901) <= not((inputs(194)) and (inputs(96)));
    layer0_outputs(902) <= (inputs(136)) or (inputs(133));
    layer0_outputs(903) <= (inputs(6)) and not (inputs(184));
    layer0_outputs(904) <= '1';
    layer0_outputs(905) <= not((inputs(208)) and (inputs(92)));
    layer0_outputs(906) <= inputs(76);
    layer0_outputs(907) <= not(inputs(119)) or (inputs(166));
    layer0_outputs(908) <= not(inputs(57));
    layer0_outputs(909) <= not((inputs(48)) xor (inputs(91)));
    layer0_outputs(910) <= not(inputs(98));
    layer0_outputs(911) <= not(inputs(181));
    layer0_outputs(912) <= inputs(73);
    layer0_outputs(913) <= not((inputs(55)) or (inputs(192)));
    layer0_outputs(914) <= not((inputs(132)) and (inputs(157)));
    layer0_outputs(915) <= inputs(200);
    layer0_outputs(916) <= inputs(135);
    layer0_outputs(917) <= inputs(89);
    layer0_outputs(918) <= not((inputs(178)) and (inputs(146)));
    layer0_outputs(919) <= (inputs(159)) and (inputs(18));
    layer0_outputs(920) <= inputs(75);
    layer0_outputs(921) <= '0';
    layer0_outputs(922) <= not(inputs(240)) or (inputs(52));
    layer0_outputs(923) <= '0';
    layer0_outputs(924) <= inputs(176);
    layer0_outputs(925) <= '0';
    layer0_outputs(926) <= not(inputs(85));
    layer0_outputs(927) <= (inputs(171)) or (inputs(198));
    layer0_outputs(928) <= (inputs(82)) and (inputs(240));
    layer0_outputs(929) <= not((inputs(189)) or (inputs(152)));
    layer0_outputs(930) <= '1';
    layer0_outputs(931) <= not(inputs(168));
    layer0_outputs(932) <= (inputs(27)) or (inputs(227));
    layer0_outputs(933) <= not(inputs(185)) or (inputs(83));
    layer0_outputs(934) <= not(inputs(112));
    layer0_outputs(935) <= (inputs(227)) xor (inputs(236));
    layer0_outputs(936) <= not(inputs(182)) or (inputs(213));
    layer0_outputs(937) <= not((inputs(66)) or (inputs(136)));
    layer0_outputs(938) <= not(inputs(67)) or (inputs(203));
    layer0_outputs(939) <= (inputs(212)) or (inputs(213));
    layer0_outputs(940) <= (inputs(90)) and not (inputs(38));
    layer0_outputs(941) <= (inputs(152)) and not (inputs(145));
    layer0_outputs(942) <= not((inputs(144)) xor (inputs(84)));
    layer0_outputs(943) <= not(inputs(73));
    layer0_outputs(944) <= not(inputs(36));
    layer0_outputs(945) <= not(inputs(237)) or (inputs(212));
    layer0_outputs(946) <= not(inputs(122)) or (inputs(16));
    layer0_outputs(947) <= not((inputs(209)) or (inputs(93)));
    layer0_outputs(948) <= '1';
    layer0_outputs(949) <= (inputs(231)) and not (inputs(161));
    layer0_outputs(950) <= (inputs(131)) xor (inputs(145));
    layer0_outputs(951) <= inputs(14);
    layer0_outputs(952) <= inputs(177);
    layer0_outputs(953) <= inputs(118);
    layer0_outputs(954) <= inputs(185);
    layer0_outputs(955) <= not(inputs(131));
    layer0_outputs(956) <= (inputs(184)) and not (inputs(66));
    layer0_outputs(957) <= (inputs(198)) and not (inputs(168));
    layer0_outputs(958) <= (inputs(214)) or (inputs(49));
    layer0_outputs(959) <= not((inputs(139)) xor (inputs(51)));
    layer0_outputs(960) <= not((inputs(211)) or (inputs(157)));
    layer0_outputs(961) <= (inputs(195)) or (inputs(146));
    layer0_outputs(962) <= not((inputs(21)) or (inputs(120)));
    layer0_outputs(963) <= inputs(167);
    layer0_outputs(964) <= not((inputs(255)) xor (inputs(233)));
    layer0_outputs(965) <= (inputs(107)) and not (inputs(21));
    layer0_outputs(966) <= not(inputs(36));
    layer0_outputs(967) <= not(inputs(64)) or (inputs(50));
    layer0_outputs(968) <= (inputs(216)) or (inputs(60));
    layer0_outputs(969) <= not((inputs(11)) and (inputs(21)));
    layer0_outputs(970) <= '0';
    layer0_outputs(971) <= not((inputs(169)) xor (inputs(129)));
    layer0_outputs(972) <= not(inputs(93)) or (inputs(156));
    layer0_outputs(973) <= inputs(233);
    layer0_outputs(974) <= inputs(16);
    layer0_outputs(975) <= '1';
    layer0_outputs(976) <= not(inputs(29));
    layer0_outputs(977) <= inputs(50);
    layer0_outputs(978) <= not(inputs(57));
    layer0_outputs(979) <= (inputs(245)) and not (inputs(78));
    layer0_outputs(980) <= not((inputs(241)) and (inputs(115)));
    layer0_outputs(981) <= not((inputs(215)) or (inputs(213)));
    layer0_outputs(982) <= not((inputs(223)) xor (inputs(154)));
    layer0_outputs(983) <= (inputs(193)) and not (inputs(44));
    layer0_outputs(984) <= not((inputs(151)) or (inputs(99)));
    layer0_outputs(985) <= not((inputs(193)) or (inputs(240)));
    layer0_outputs(986) <= (inputs(223)) xor (inputs(200));
    layer0_outputs(987) <= (inputs(15)) and not (inputs(92));
    layer0_outputs(988) <= (inputs(125)) or (inputs(63));
    layer0_outputs(989) <= (inputs(110)) and not (inputs(14));
    layer0_outputs(990) <= inputs(215);
    layer0_outputs(991) <= inputs(90);
    layer0_outputs(992) <= (inputs(85)) and not (inputs(224));
    layer0_outputs(993) <= (inputs(182)) or (inputs(178));
    layer0_outputs(994) <= (inputs(222)) and not (inputs(228));
    layer0_outputs(995) <= not(inputs(155));
    layer0_outputs(996) <= '0';
    layer0_outputs(997) <= not(inputs(32)) or (inputs(209));
    layer0_outputs(998) <= not(inputs(205));
    layer0_outputs(999) <= (inputs(55)) or (inputs(11));
    layer0_outputs(1000) <= (inputs(136)) and not (inputs(141));
    layer0_outputs(1001) <= not((inputs(33)) or (inputs(154)));
    layer0_outputs(1002) <= (inputs(153)) xor (inputs(49));
    layer0_outputs(1003) <= not(inputs(40)) or (inputs(32));
    layer0_outputs(1004) <= not((inputs(105)) xor (inputs(11)));
    layer0_outputs(1005) <= not(inputs(181));
    layer0_outputs(1006) <= (inputs(2)) and (inputs(40));
    layer0_outputs(1007) <= inputs(102);
    layer0_outputs(1008) <= (inputs(120)) and not (inputs(112));
    layer0_outputs(1009) <= not(inputs(4));
    layer0_outputs(1010) <= not(inputs(153));
    layer0_outputs(1011) <= not((inputs(1)) xor (inputs(127)));
    layer0_outputs(1012) <= '1';
    layer0_outputs(1013) <= inputs(56);
    layer0_outputs(1014) <= inputs(67);
    layer0_outputs(1015) <= not(inputs(215)) or (inputs(238));
    layer0_outputs(1016) <= not((inputs(32)) or (inputs(207)));
    layer0_outputs(1017) <= not((inputs(79)) xor (inputs(219)));
    layer0_outputs(1018) <= '1';
    layer0_outputs(1019) <= not(inputs(201)) or (inputs(86));
    layer0_outputs(1020) <= not((inputs(110)) or (inputs(93)));
    layer0_outputs(1021) <= not((inputs(232)) or (inputs(152)));
    layer0_outputs(1022) <= inputs(155);
    layer0_outputs(1023) <= not((inputs(123)) or (inputs(175)));
    layer0_outputs(1024) <= (inputs(202)) xor (inputs(109));
    layer0_outputs(1025) <= not(inputs(215)) or (inputs(14));
    layer0_outputs(1026) <= not(inputs(140));
    layer0_outputs(1027) <= not((inputs(128)) and (inputs(115)));
    layer0_outputs(1028) <= (inputs(62)) and not (inputs(111));
    layer0_outputs(1029) <= (inputs(102)) and not (inputs(51));
    layer0_outputs(1030) <= (inputs(250)) and not (inputs(189));
    layer0_outputs(1031) <= not(inputs(68)) or (inputs(190));
    layer0_outputs(1032) <= '0';
    layer0_outputs(1033) <= inputs(82);
    layer0_outputs(1034) <= '0';
    layer0_outputs(1035) <= not(inputs(231));
    layer0_outputs(1036) <= not(inputs(249)) or (inputs(101));
    layer0_outputs(1037) <= (inputs(204)) and (inputs(218));
    layer0_outputs(1038) <= (inputs(218)) and not (inputs(48));
    layer0_outputs(1039) <= not((inputs(248)) or (inputs(211)));
    layer0_outputs(1040) <= inputs(186);
    layer0_outputs(1041) <= '1';
    layer0_outputs(1042) <= not(inputs(141));
    layer0_outputs(1043) <= (inputs(128)) and not (inputs(112));
    layer0_outputs(1044) <= inputs(59);
    layer0_outputs(1045) <= (inputs(99)) and not (inputs(97));
    layer0_outputs(1046) <= (inputs(203)) xor (inputs(94));
    layer0_outputs(1047) <= inputs(133);
    layer0_outputs(1048) <= not((inputs(88)) xor (inputs(210)));
    layer0_outputs(1049) <= (inputs(71)) xor (inputs(79));
    layer0_outputs(1050) <= (inputs(35)) or (inputs(193));
    layer0_outputs(1051) <= inputs(71);
    layer0_outputs(1052) <= not(inputs(37)) or (inputs(19));
    layer0_outputs(1053) <= inputs(249);
    layer0_outputs(1054) <= not((inputs(101)) or (inputs(229)));
    layer0_outputs(1055) <= (inputs(51)) and (inputs(23));
    layer0_outputs(1056) <= (inputs(165)) or (inputs(126));
    layer0_outputs(1057) <= (inputs(5)) and not (inputs(218));
    layer0_outputs(1058) <= not(inputs(92)) or (inputs(37));
    layer0_outputs(1059) <= not(inputs(181));
    layer0_outputs(1060) <= inputs(214);
    layer0_outputs(1061) <= (inputs(193)) or (inputs(200));
    layer0_outputs(1062) <= not(inputs(107)) or (inputs(252));
    layer0_outputs(1063) <= inputs(218);
    layer0_outputs(1064) <= (inputs(157)) and not (inputs(233));
    layer0_outputs(1065) <= inputs(149);
    layer0_outputs(1066) <= (inputs(115)) and not (inputs(227));
    layer0_outputs(1067) <= '1';
    layer0_outputs(1068) <= (inputs(235)) or (inputs(202));
    layer0_outputs(1069) <= not((inputs(69)) or (inputs(104)));
    layer0_outputs(1070) <= inputs(240);
    layer0_outputs(1071) <= inputs(197);
    layer0_outputs(1072) <= inputs(183);
    layer0_outputs(1073) <= inputs(29);
    layer0_outputs(1074) <= not(inputs(139)) or (inputs(36));
    layer0_outputs(1075) <= '1';
    layer0_outputs(1076) <= not(inputs(82));
    layer0_outputs(1077) <= (inputs(163)) xor (inputs(51));
    layer0_outputs(1078) <= not(inputs(147));
    layer0_outputs(1079) <= (inputs(147)) or (inputs(171));
    layer0_outputs(1080) <= inputs(165);
    layer0_outputs(1081) <= (inputs(211)) or (inputs(82));
    layer0_outputs(1082) <= not((inputs(39)) xor (inputs(87)));
    layer0_outputs(1083) <= not((inputs(205)) or (inputs(228)));
    layer0_outputs(1084) <= not((inputs(225)) xor (inputs(81)));
    layer0_outputs(1085) <= inputs(182);
    layer0_outputs(1086) <= (inputs(149)) and not (inputs(47));
    layer0_outputs(1087) <= not((inputs(198)) or (inputs(89)));
    layer0_outputs(1088) <= (inputs(55)) and not (inputs(30));
    layer0_outputs(1089) <= not(inputs(112));
    layer0_outputs(1090) <= not((inputs(224)) xor (inputs(237)));
    layer0_outputs(1091) <= (inputs(21)) and not (inputs(47));
    layer0_outputs(1092) <= '1';
    layer0_outputs(1093) <= not((inputs(209)) xor (inputs(253)));
    layer0_outputs(1094) <= not(inputs(91)) or (inputs(144));
    layer0_outputs(1095) <= not(inputs(105));
    layer0_outputs(1096) <= not((inputs(243)) xor (inputs(147)));
    layer0_outputs(1097) <= not((inputs(226)) and (inputs(41)));
    layer0_outputs(1098) <= (inputs(218)) xor (inputs(74));
    layer0_outputs(1099) <= not(inputs(21));
    layer0_outputs(1100) <= not((inputs(105)) or (inputs(24)));
    layer0_outputs(1101) <= inputs(144);
    layer0_outputs(1102) <= (inputs(76)) or (inputs(54));
    layer0_outputs(1103) <= not((inputs(193)) or (inputs(32)));
    layer0_outputs(1104) <= not(inputs(106)) or (inputs(211));
    layer0_outputs(1105) <= '1';
    layer0_outputs(1106) <= (inputs(233)) and not (inputs(17));
    layer0_outputs(1107) <= not(inputs(161)) or (inputs(238));
    layer0_outputs(1108) <= not(inputs(196)) or (inputs(17));
    layer0_outputs(1109) <= not((inputs(116)) or (inputs(125)));
    layer0_outputs(1110) <= not((inputs(92)) or (inputs(4)));
    layer0_outputs(1111) <= inputs(132);
    layer0_outputs(1112) <= (inputs(140)) or (inputs(150));
    layer0_outputs(1113) <= (inputs(153)) xor (inputs(246));
    layer0_outputs(1114) <= (inputs(80)) or (inputs(182));
    layer0_outputs(1115) <= not(inputs(128)) or (inputs(49));
    layer0_outputs(1116) <= not((inputs(193)) or (inputs(76)));
    layer0_outputs(1117) <= not(inputs(138));
    layer0_outputs(1118) <= not(inputs(54));
    layer0_outputs(1119) <= inputs(37);
    layer0_outputs(1120) <= not(inputs(19)) or (inputs(159));
    layer0_outputs(1121) <= inputs(147);
    layer0_outputs(1122) <= (inputs(134)) and (inputs(12));
    layer0_outputs(1123) <= inputs(236);
    layer0_outputs(1124) <= (inputs(189)) or (inputs(88));
    layer0_outputs(1125) <= '0';
    layer0_outputs(1126) <= not((inputs(87)) xor (inputs(219)));
    layer0_outputs(1127) <= not((inputs(203)) or (inputs(230)));
    layer0_outputs(1128) <= '1';
    layer0_outputs(1129) <= not(inputs(117));
    layer0_outputs(1130) <= (inputs(121)) and not (inputs(96));
    layer0_outputs(1131) <= not(inputs(244)) or (inputs(254));
    layer0_outputs(1132) <= not(inputs(216));
    layer0_outputs(1133) <= (inputs(85)) or (inputs(179));
    layer0_outputs(1134) <= inputs(91);
    layer0_outputs(1135) <= not((inputs(4)) or (inputs(74)));
    layer0_outputs(1136) <= not((inputs(133)) or (inputs(173)));
    layer0_outputs(1137) <= not(inputs(154));
    layer0_outputs(1138) <= inputs(216);
    layer0_outputs(1139) <= not(inputs(58));
    layer0_outputs(1140) <= '1';
    layer0_outputs(1141) <= inputs(41);
    layer0_outputs(1142) <= not((inputs(115)) or (inputs(116)));
    layer0_outputs(1143) <= (inputs(129)) and not (inputs(231));
    layer0_outputs(1144) <= not(inputs(167));
    layer0_outputs(1145) <= not((inputs(133)) xor (inputs(80)));
    layer0_outputs(1146) <= not(inputs(7));
    layer0_outputs(1147) <= (inputs(127)) and not (inputs(48));
    layer0_outputs(1148) <= not(inputs(146)) or (inputs(246));
    layer0_outputs(1149) <= (inputs(10)) and not (inputs(181));
    layer0_outputs(1150) <= not((inputs(178)) or (inputs(34)));
    layer0_outputs(1151) <= not((inputs(94)) or (inputs(99)));
    layer0_outputs(1152) <= inputs(6);
    layer0_outputs(1153) <= not((inputs(4)) or (inputs(41)));
    layer0_outputs(1154) <= not(inputs(237)) or (inputs(48));
    layer0_outputs(1155) <= (inputs(243)) and not (inputs(110));
    layer0_outputs(1156) <= not((inputs(77)) xor (inputs(25)));
    layer0_outputs(1157) <= '1';
    layer0_outputs(1158) <= inputs(119);
    layer0_outputs(1159) <= (inputs(238)) and not (inputs(39));
    layer0_outputs(1160) <= not((inputs(50)) or (inputs(179)));
    layer0_outputs(1161) <= (inputs(202)) and not (inputs(225));
    layer0_outputs(1162) <= not(inputs(118)) or (inputs(67));
    layer0_outputs(1163) <= not(inputs(89));
    layer0_outputs(1164) <= (inputs(131)) or (inputs(60));
    layer0_outputs(1165) <= not(inputs(126)) or (inputs(244));
    layer0_outputs(1166) <= (inputs(118)) or (inputs(196));
    layer0_outputs(1167) <= not(inputs(78));
    layer0_outputs(1168) <= (inputs(41)) or (inputs(54));
    layer0_outputs(1169) <= (inputs(87)) and not (inputs(237));
    layer0_outputs(1170) <= not(inputs(248));
    layer0_outputs(1171) <= (inputs(188)) and not (inputs(150));
    layer0_outputs(1172) <= inputs(213);
    layer0_outputs(1173) <= not((inputs(163)) or (inputs(201)));
    layer0_outputs(1174) <= not((inputs(139)) or (inputs(132)));
    layer0_outputs(1175) <= (inputs(163)) and not (inputs(29));
    layer0_outputs(1176) <= not((inputs(22)) and (inputs(20)));
    layer0_outputs(1177) <= not(inputs(73)) or (inputs(31));
    layer0_outputs(1178) <= not((inputs(56)) xor (inputs(134)));
    layer0_outputs(1179) <= '0';
    layer0_outputs(1180) <= not((inputs(0)) or (inputs(235)));
    layer0_outputs(1181) <= (inputs(251)) xor (inputs(74));
    layer0_outputs(1182) <= inputs(38);
    layer0_outputs(1183) <= not(inputs(93));
    layer0_outputs(1184) <= not((inputs(182)) or (inputs(31)));
    layer0_outputs(1185) <= inputs(34);
    layer0_outputs(1186) <= (inputs(129)) or (inputs(190));
    layer0_outputs(1187) <= '1';
    layer0_outputs(1188) <= not((inputs(13)) and (inputs(224)));
    layer0_outputs(1189) <= (inputs(238)) or (inputs(233));
    layer0_outputs(1190) <= not(inputs(191));
    layer0_outputs(1191) <= not(inputs(126)) or (inputs(72));
    layer0_outputs(1192) <= not(inputs(152));
    layer0_outputs(1193) <= not(inputs(133)) or (inputs(67));
    layer0_outputs(1194) <= '0';
    layer0_outputs(1195) <= (inputs(50)) or (inputs(114));
    layer0_outputs(1196) <= not(inputs(245)) or (inputs(9));
    layer0_outputs(1197) <= not((inputs(87)) or (inputs(27)));
    layer0_outputs(1198) <= not((inputs(77)) or (inputs(113)));
    layer0_outputs(1199) <= not((inputs(41)) or (inputs(163)));
    layer0_outputs(1200) <= not((inputs(157)) xor (inputs(232)));
    layer0_outputs(1201) <= not((inputs(244)) xor (inputs(54)));
    layer0_outputs(1202) <= not(inputs(245)) or (inputs(151));
    layer0_outputs(1203) <= (inputs(40)) and not (inputs(161));
    layer0_outputs(1204) <= not((inputs(70)) xor (inputs(15)));
    layer0_outputs(1205) <= not(inputs(149)) or (inputs(30));
    layer0_outputs(1206) <= not((inputs(117)) xor (inputs(112)));
    layer0_outputs(1207) <= inputs(219);
    layer0_outputs(1208) <= not(inputs(172));
    layer0_outputs(1209) <= (inputs(36)) or (inputs(122));
    layer0_outputs(1210) <= not((inputs(245)) and (inputs(203)));
    layer0_outputs(1211) <= (inputs(227)) and not (inputs(13));
    layer0_outputs(1212) <= not(inputs(230));
    layer0_outputs(1213) <= not(inputs(117));
    layer0_outputs(1214) <= '1';
    layer0_outputs(1215) <= (inputs(155)) or (inputs(253));
    layer0_outputs(1216) <= (inputs(79)) or (inputs(229));
    layer0_outputs(1217) <= not(inputs(168)) or (inputs(140));
    layer0_outputs(1218) <= not((inputs(195)) xor (inputs(55)));
    layer0_outputs(1219) <= (inputs(65)) and not (inputs(44));
    layer0_outputs(1220) <= (inputs(70)) or (inputs(1));
    layer0_outputs(1221) <= (inputs(12)) and not (inputs(42));
    layer0_outputs(1222) <= (inputs(32)) and (inputs(24));
    layer0_outputs(1223) <= not(inputs(231)) or (inputs(174));
    layer0_outputs(1224) <= not(inputs(69)) or (inputs(145));
    layer0_outputs(1225) <= inputs(86);
    layer0_outputs(1226) <= (inputs(72)) and not (inputs(128));
    layer0_outputs(1227) <= not((inputs(174)) or (inputs(158)));
    layer0_outputs(1228) <= (inputs(219)) xor (inputs(139));
    layer0_outputs(1229) <= inputs(114);
    layer0_outputs(1230) <= '1';
    layer0_outputs(1231) <= (inputs(80)) or (inputs(126));
    layer0_outputs(1232) <= not(inputs(48));
    layer0_outputs(1233) <= (inputs(124)) or (inputs(42));
    layer0_outputs(1234) <= '1';
    layer0_outputs(1235) <= '1';
    layer0_outputs(1236) <= inputs(152);
    layer0_outputs(1237) <= inputs(75);
    layer0_outputs(1238) <= not((inputs(248)) and (inputs(110)));
    layer0_outputs(1239) <= (inputs(71)) or (inputs(180));
    layer0_outputs(1240) <= (inputs(134)) xor (inputs(246));
    layer0_outputs(1241) <= not((inputs(161)) xor (inputs(193)));
    layer0_outputs(1242) <= not(inputs(158)) or (inputs(45));
    layer0_outputs(1243) <= not((inputs(52)) or (inputs(176)));
    layer0_outputs(1244) <= (inputs(105)) or (inputs(99));
    layer0_outputs(1245) <= not((inputs(85)) xor (inputs(18)));
    layer0_outputs(1246) <= inputs(199);
    layer0_outputs(1247) <= (inputs(11)) and (inputs(211));
    layer0_outputs(1248) <= (inputs(23)) and not (inputs(133));
    layer0_outputs(1249) <= not(inputs(247));
    layer0_outputs(1250) <= inputs(89);
    layer0_outputs(1251) <= inputs(147);
    layer0_outputs(1252) <= not(inputs(23));
    layer0_outputs(1253) <= not((inputs(215)) or (inputs(109)));
    layer0_outputs(1254) <= (inputs(63)) and (inputs(80));
    layer0_outputs(1255) <= (inputs(14)) and not (inputs(176));
    layer0_outputs(1256) <= (inputs(141)) and not (inputs(21));
    layer0_outputs(1257) <= (inputs(42)) xor (inputs(47));
    layer0_outputs(1258) <= not((inputs(185)) and (inputs(237)));
    layer0_outputs(1259) <= (inputs(84)) or (inputs(58));
    layer0_outputs(1260) <= (inputs(149)) and not (inputs(75));
    layer0_outputs(1261) <= '0';
    layer0_outputs(1262) <= inputs(139);
    layer0_outputs(1263) <= not(inputs(245));
    layer0_outputs(1264) <= inputs(87);
    layer0_outputs(1265) <= (inputs(204)) and not (inputs(203));
    layer0_outputs(1266) <= not(inputs(149));
    layer0_outputs(1267) <= not(inputs(144));
    layer0_outputs(1268) <= not((inputs(177)) or (inputs(108)));
    layer0_outputs(1269) <= inputs(81);
    layer0_outputs(1270) <= not((inputs(22)) or (inputs(185)));
    layer0_outputs(1271) <= (inputs(137)) xor (inputs(226));
    layer0_outputs(1272) <= not(inputs(239)) or (inputs(37));
    layer0_outputs(1273) <= inputs(17);
    layer0_outputs(1274) <= not((inputs(89)) xor (inputs(215)));
    layer0_outputs(1275) <= not(inputs(234)) or (inputs(249));
    layer0_outputs(1276) <= not((inputs(146)) xor (inputs(69)));
    layer0_outputs(1277) <= inputs(188);
    layer0_outputs(1278) <= not((inputs(251)) xor (inputs(72)));
    layer0_outputs(1279) <= inputs(208);
    layer0_outputs(1280) <= not(inputs(52)) or (inputs(94));
    layer0_outputs(1281) <= not(inputs(49)) or (inputs(199));
    layer0_outputs(1282) <= (inputs(79)) and not (inputs(4));
    layer0_outputs(1283) <= (inputs(69)) and not (inputs(146));
    layer0_outputs(1284) <= not((inputs(255)) xor (inputs(205)));
    layer0_outputs(1285) <= inputs(137);
    layer0_outputs(1286) <= (inputs(225)) xor (inputs(40));
    layer0_outputs(1287) <= (inputs(220)) or (inputs(147));
    layer0_outputs(1288) <= (inputs(199)) or (inputs(211));
    layer0_outputs(1289) <= (inputs(85)) or (inputs(108));
    layer0_outputs(1290) <= inputs(22);
    layer0_outputs(1291) <= (inputs(23)) and not (inputs(13));
    layer0_outputs(1292) <= not(inputs(149));
    layer0_outputs(1293) <= not((inputs(224)) and (inputs(183)));
    layer0_outputs(1294) <= not(inputs(76)) or (inputs(9));
    layer0_outputs(1295) <= not(inputs(16));
    layer0_outputs(1296) <= (inputs(218)) or (inputs(28));
    layer0_outputs(1297) <= not(inputs(163));
    layer0_outputs(1298) <= (inputs(62)) and (inputs(138));
    layer0_outputs(1299) <= (inputs(45)) or (inputs(25));
    layer0_outputs(1300) <= not(inputs(75)) or (inputs(151));
    layer0_outputs(1301) <= inputs(218);
    layer0_outputs(1302) <= '1';
    layer0_outputs(1303) <= not(inputs(31));
    layer0_outputs(1304) <= not(inputs(174)) or (inputs(47));
    layer0_outputs(1305) <= not(inputs(223)) or (inputs(213));
    layer0_outputs(1306) <= '0';
    layer0_outputs(1307) <= '0';
    layer0_outputs(1308) <= (inputs(56)) xor (inputs(128));
    layer0_outputs(1309) <= not(inputs(183)) or (inputs(105));
    layer0_outputs(1310) <= not((inputs(26)) and (inputs(5)));
    layer0_outputs(1311) <= not(inputs(168));
    layer0_outputs(1312) <= not((inputs(17)) and (inputs(66)));
    layer0_outputs(1313) <= not((inputs(182)) xor (inputs(96)));
    layer0_outputs(1314) <= inputs(215);
    layer0_outputs(1315) <= not((inputs(96)) or (inputs(55)));
    layer0_outputs(1316) <= (inputs(227)) xor (inputs(29));
    layer0_outputs(1317) <= inputs(154);
    layer0_outputs(1318) <= (inputs(14)) xor (inputs(159));
    layer0_outputs(1319) <= not((inputs(83)) or (inputs(194)));
    layer0_outputs(1320) <= (inputs(135)) or (inputs(181));
    layer0_outputs(1321) <= (inputs(149)) or (inputs(157));
    layer0_outputs(1322) <= (inputs(174)) and not (inputs(77));
    layer0_outputs(1323) <= (inputs(85)) and not (inputs(33));
    layer0_outputs(1324) <= not(inputs(165));
    layer0_outputs(1325) <= not(inputs(111));
    layer0_outputs(1326) <= inputs(177);
    layer0_outputs(1327) <= not(inputs(14)) or (inputs(19));
    layer0_outputs(1328) <= not(inputs(230)) or (inputs(144));
    layer0_outputs(1329) <= inputs(172);
    layer0_outputs(1330) <= (inputs(23)) and not (inputs(10));
    layer0_outputs(1331) <= not((inputs(213)) or (inputs(55)));
    layer0_outputs(1332) <= not((inputs(158)) or (inputs(93)));
    layer0_outputs(1333) <= not(inputs(127)) or (inputs(235));
    layer0_outputs(1334) <= inputs(125);
    layer0_outputs(1335) <= '0';
    layer0_outputs(1336) <= not(inputs(216)) or (inputs(38));
    layer0_outputs(1337) <= not((inputs(237)) and (inputs(14)));
    layer0_outputs(1338) <= not(inputs(213)) or (inputs(91));
    layer0_outputs(1339) <= inputs(24);
    layer0_outputs(1340) <= not(inputs(124));
    layer0_outputs(1341) <= not((inputs(222)) and (inputs(142)));
    layer0_outputs(1342) <= (inputs(174)) or (inputs(185));
    layer0_outputs(1343) <= not(inputs(230));
    layer0_outputs(1344) <= inputs(181);
    layer0_outputs(1345) <= not(inputs(127));
    layer0_outputs(1346) <= not(inputs(26));
    layer0_outputs(1347) <= not(inputs(40));
    layer0_outputs(1348) <= (inputs(17)) xor (inputs(60));
    layer0_outputs(1349) <= '0';
    layer0_outputs(1350) <= '1';
    layer0_outputs(1351) <= '1';
    layer0_outputs(1352) <= not(inputs(45)) or (inputs(242));
    layer0_outputs(1353) <= not(inputs(184)) or (inputs(190));
    layer0_outputs(1354) <= '0';
    layer0_outputs(1355) <= not((inputs(220)) xor (inputs(18)));
    layer0_outputs(1356) <= (inputs(160)) xor (inputs(132));
    layer0_outputs(1357) <= not(inputs(126));
    layer0_outputs(1358) <= not((inputs(188)) xor (inputs(57)));
    layer0_outputs(1359) <= inputs(143);
    layer0_outputs(1360) <= '1';
    layer0_outputs(1361) <= not((inputs(162)) xor (inputs(109)));
    layer0_outputs(1362) <= inputs(175);
    layer0_outputs(1363) <= not(inputs(75)) or (inputs(223));
    layer0_outputs(1364) <= (inputs(158)) xor (inputs(33));
    layer0_outputs(1365) <= not(inputs(201)) or (inputs(219));
    layer0_outputs(1366) <= not(inputs(91)) or (inputs(219));
    layer0_outputs(1367) <= (inputs(157)) xor (inputs(126));
    layer0_outputs(1368) <= not(inputs(197));
    layer0_outputs(1369) <= inputs(65);
    layer0_outputs(1370) <= inputs(73);
    layer0_outputs(1371) <= (inputs(40)) and not (inputs(131));
    layer0_outputs(1372) <= not((inputs(10)) or (inputs(152)));
    layer0_outputs(1373) <= (inputs(37)) or (inputs(147));
    layer0_outputs(1374) <= (inputs(17)) or (inputs(117));
    layer0_outputs(1375) <= not(inputs(190)) or (inputs(164));
    layer0_outputs(1376) <= not((inputs(110)) or (inputs(163)));
    layer0_outputs(1377) <= not((inputs(10)) xor (inputs(193)));
    layer0_outputs(1378) <= (inputs(196)) and not (inputs(50));
    layer0_outputs(1379) <= '0';
    layer0_outputs(1380) <= '1';
    layer0_outputs(1381) <= not(inputs(24));
    layer0_outputs(1382) <= not(inputs(162));
    layer0_outputs(1383) <= not((inputs(175)) and (inputs(221)));
    layer0_outputs(1384) <= not(inputs(174));
    layer0_outputs(1385) <= inputs(61);
    layer0_outputs(1386) <= not((inputs(199)) or (inputs(234)));
    layer0_outputs(1387) <= not(inputs(198)) or (inputs(126));
    layer0_outputs(1388) <= not((inputs(244)) xor (inputs(141)));
    layer0_outputs(1389) <= '1';
    layer0_outputs(1390) <= not(inputs(246)) or (inputs(254));
    layer0_outputs(1391) <= inputs(216);
    layer0_outputs(1392) <= (inputs(95)) and not (inputs(190));
    layer0_outputs(1393) <= (inputs(212)) or (inputs(77));
    layer0_outputs(1394) <= not((inputs(53)) or (inputs(255)));
    layer0_outputs(1395) <= '1';
    layer0_outputs(1396) <= not(inputs(119)) or (inputs(174));
    layer0_outputs(1397) <= inputs(233);
    layer0_outputs(1398) <= (inputs(11)) xor (inputs(167));
    layer0_outputs(1399) <= (inputs(33)) and (inputs(212));
    layer0_outputs(1400) <= '1';
    layer0_outputs(1401) <= not(inputs(42));
    layer0_outputs(1402) <= not(inputs(84));
    layer0_outputs(1403) <= (inputs(167)) and not (inputs(76));
    layer0_outputs(1404) <= not(inputs(163)) or (inputs(206));
    layer0_outputs(1405) <= (inputs(203)) xor (inputs(81));
    layer0_outputs(1406) <= not(inputs(56));
    layer0_outputs(1407) <= not((inputs(137)) xor (inputs(50)));
    layer0_outputs(1408) <= (inputs(108)) or (inputs(194));
    layer0_outputs(1409) <= (inputs(191)) and not (inputs(29));
    layer0_outputs(1410) <= not(inputs(53));
    layer0_outputs(1411) <= not(inputs(12));
    layer0_outputs(1412) <= (inputs(183)) and not (inputs(85));
    layer0_outputs(1413) <= not(inputs(121));
    layer0_outputs(1414) <= not((inputs(203)) or (inputs(195)));
    layer0_outputs(1415) <= not(inputs(193));
    layer0_outputs(1416) <= not(inputs(153));
    layer0_outputs(1417) <= not((inputs(55)) and (inputs(42)));
    layer0_outputs(1418) <= not(inputs(9));
    layer0_outputs(1419) <= (inputs(3)) and (inputs(62));
    layer0_outputs(1420) <= (inputs(56)) and not (inputs(246));
    layer0_outputs(1421) <= (inputs(192)) or (inputs(21));
    layer0_outputs(1422) <= (inputs(234)) and not (inputs(203));
    layer0_outputs(1423) <= (inputs(15)) or (inputs(161));
    layer0_outputs(1424) <= (inputs(76)) and not (inputs(250));
    layer0_outputs(1425) <= '0';
    layer0_outputs(1426) <= not(inputs(187));
    layer0_outputs(1427) <= not((inputs(181)) xor (inputs(110)));
    layer0_outputs(1428) <= not(inputs(5));
    layer0_outputs(1429) <= not(inputs(134)) or (inputs(104));
    layer0_outputs(1430) <= not((inputs(86)) xor (inputs(7)));
    layer0_outputs(1431) <= not(inputs(103));
    layer0_outputs(1432) <= (inputs(52)) or (inputs(17));
    layer0_outputs(1433) <= not((inputs(63)) xor (inputs(134)));
    layer0_outputs(1434) <= not(inputs(29)) or (inputs(80));
    layer0_outputs(1435) <= not((inputs(20)) or (inputs(167)));
    layer0_outputs(1436) <= not(inputs(37)) or (inputs(18));
    layer0_outputs(1437) <= inputs(245);
    layer0_outputs(1438) <= not((inputs(223)) xor (inputs(125)));
    layer0_outputs(1439) <= inputs(153);
    layer0_outputs(1440) <= not((inputs(254)) or (inputs(41)));
    layer0_outputs(1441) <= not(inputs(164)) or (inputs(66));
    layer0_outputs(1442) <= not(inputs(242)) or (inputs(212));
    layer0_outputs(1443) <= not(inputs(86)) or (inputs(164));
    layer0_outputs(1444) <= (inputs(150)) and not (inputs(235));
    layer0_outputs(1445) <= (inputs(61)) and not (inputs(52));
    layer0_outputs(1446) <= not(inputs(134)) or (inputs(47));
    layer0_outputs(1447) <= inputs(61);
    layer0_outputs(1448) <= inputs(182);
    layer0_outputs(1449) <= (inputs(213)) and not (inputs(138));
    layer0_outputs(1450) <= (inputs(205)) and not (inputs(184));
    layer0_outputs(1451) <= (inputs(31)) and not (inputs(37));
    layer0_outputs(1452) <= inputs(3);
    layer0_outputs(1453) <= not(inputs(61)) or (inputs(176));
    layer0_outputs(1454) <= (inputs(121)) xor (inputs(147));
    layer0_outputs(1455) <= (inputs(160)) or (inputs(189));
    layer0_outputs(1456) <= inputs(46);
    layer0_outputs(1457) <= not((inputs(114)) and (inputs(194)));
    layer0_outputs(1458) <= not((inputs(4)) or (inputs(133)));
    layer0_outputs(1459) <= not(inputs(15)) or (inputs(135));
    layer0_outputs(1460) <= (inputs(33)) or (inputs(125));
    layer0_outputs(1461) <= not((inputs(92)) or (inputs(199)));
    layer0_outputs(1462) <= not((inputs(57)) or (inputs(251)));
    layer0_outputs(1463) <= not(inputs(124));
    layer0_outputs(1464) <= '0';
    layer0_outputs(1465) <= (inputs(38)) or (inputs(139));
    layer0_outputs(1466) <= (inputs(240)) and (inputs(43));
    layer0_outputs(1467) <= '1';
    layer0_outputs(1468) <= not((inputs(46)) xor (inputs(217)));
    layer0_outputs(1469) <= (inputs(124)) and not (inputs(67));
    layer0_outputs(1470) <= not(inputs(33));
    layer0_outputs(1471) <= (inputs(1)) or (inputs(101));
    layer0_outputs(1472) <= not((inputs(211)) and (inputs(131)));
    layer0_outputs(1473) <= not(inputs(38)) or (inputs(17));
    layer0_outputs(1474) <= inputs(26);
    layer0_outputs(1475) <= inputs(148);
    layer0_outputs(1476) <= not(inputs(93));
    layer0_outputs(1477) <= '1';
    layer0_outputs(1478) <= not(inputs(68));
    layer0_outputs(1479) <= inputs(244);
    layer0_outputs(1480) <= (inputs(40)) and not (inputs(160));
    layer0_outputs(1481) <= not(inputs(120)) or (inputs(48));
    layer0_outputs(1482) <= not((inputs(22)) or (inputs(241)));
    layer0_outputs(1483) <= (inputs(73)) or (inputs(197));
    layer0_outputs(1484) <= inputs(89);
    layer0_outputs(1485) <= not((inputs(51)) and (inputs(167)));
    layer0_outputs(1486) <= '0';
    layer0_outputs(1487) <= not(inputs(5)) or (inputs(226));
    layer0_outputs(1488) <= '0';
    layer0_outputs(1489) <= (inputs(66)) and (inputs(172));
    layer0_outputs(1490) <= not((inputs(70)) and (inputs(97)));
    layer0_outputs(1491) <= not((inputs(22)) or (inputs(170)));
    layer0_outputs(1492) <= (inputs(151)) and not (inputs(237));
    layer0_outputs(1493) <= not((inputs(131)) or (inputs(124)));
    layer0_outputs(1494) <= (inputs(28)) or (inputs(212));
    layer0_outputs(1495) <= not(inputs(57));
    layer0_outputs(1496) <= not(inputs(183)) or (inputs(4));
    layer0_outputs(1497) <= (inputs(208)) or (inputs(8));
    layer0_outputs(1498) <= not(inputs(197)) or (inputs(142));
    layer0_outputs(1499) <= (inputs(92)) or (inputs(198));
    layer0_outputs(1500) <= (inputs(242)) or (inputs(112));
    layer0_outputs(1501) <= not(inputs(122)) or (inputs(33));
    layer0_outputs(1502) <= (inputs(233)) and not (inputs(25));
    layer0_outputs(1503) <= inputs(155);
    layer0_outputs(1504) <= not(inputs(72));
    layer0_outputs(1505) <= (inputs(254)) or (inputs(228));
    layer0_outputs(1506) <= '0';
    layer0_outputs(1507) <= inputs(52);
    layer0_outputs(1508) <= not((inputs(218)) and (inputs(41)));
    layer0_outputs(1509) <= (inputs(3)) and not (inputs(39));
    layer0_outputs(1510) <= (inputs(125)) and not (inputs(151));
    layer0_outputs(1511) <= (inputs(224)) xor (inputs(215));
    layer0_outputs(1512) <= (inputs(2)) and not (inputs(43));
    layer0_outputs(1513) <= inputs(133);
    layer0_outputs(1514) <= not((inputs(65)) or (inputs(68)));
    layer0_outputs(1515) <= '0';
    layer0_outputs(1516) <= (inputs(125)) xor (inputs(18));
    layer0_outputs(1517) <= inputs(0);
    layer0_outputs(1518) <= not(inputs(118)) or (inputs(67));
    layer0_outputs(1519) <= '1';
    layer0_outputs(1520) <= not(inputs(122));
    layer0_outputs(1521) <= not((inputs(205)) xor (inputs(7)));
    layer0_outputs(1522) <= (inputs(175)) and not (inputs(95));
    layer0_outputs(1523) <= (inputs(183)) and not (inputs(242));
    layer0_outputs(1524) <= '1';
    layer0_outputs(1525) <= inputs(48);
    layer0_outputs(1526) <= not(inputs(196));
    layer0_outputs(1527) <= not(inputs(153));
    layer0_outputs(1528) <= inputs(141);
    layer0_outputs(1529) <= (inputs(234)) and not (inputs(50));
    layer0_outputs(1530) <= not((inputs(176)) xor (inputs(167)));
    layer0_outputs(1531) <= '0';
    layer0_outputs(1532) <= not(inputs(174)) or (inputs(211));
    layer0_outputs(1533) <= inputs(136);
    layer0_outputs(1534) <= not((inputs(13)) or (inputs(196)));
    layer0_outputs(1535) <= not(inputs(152));
    layer0_outputs(1536) <= (inputs(144)) and (inputs(251));
    layer0_outputs(1537) <= not(inputs(108)) or (inputs(14));
    layer0_outputs(1538) <= inputs(164);
    layer0_outputs(1539) <= not(inputs(187)) or (inputs(192));
    layer0_outputs(1540) <= inputs(89);
    layer0_outputs(1541) <= (inputs(37)) and not (inputs(179));
    layer0_outputs(1542) <= not((inputs(160)) or (inputs(3)));
    layer0_outputs(1543) <= not((inputs(61)) xor (inputs(24)));
    layer0_outputs(1544) <= not(inputs(88)) or (inputs(90));
    layer0_outputs(1545) <= not(inputs(74));
    layer0_outputs(1546) <= not(inputs(123));
    layer0_outputs(1547) <= (inputs(204)) and (inputs(162));
    layer0_outputs(1548) <= not(inputs(163)) or (inputs(154));
    layer0_outputs(1549) <= (inputs(136)) and not (inputs(177));
    layer0_outputs(1550) <= not(inputs(228));
    layer0_outputs(1551) <= not(inputs(85)) or (inputs(205));
    layer0_outputs(1552) <= inputs(131);
    layer0_outputs(1553) <= not((inputs(74)) xor (inputs(58)));
    layer0_outputs(1554) <= not(inputs(191));
    layer0_outputs(1555) <= not(inputs(117));
    layer0_outputs(1556) <= not(inputs(90));
    layer0_outputs(1557) <= (inputs(55)) and not (inputs(102));
    layer0_outputs(1558) <= not(inputs(213)) or (inputs(206));
    layer0_outputs(1559) <= not((inputs(156)) xor (inputs(50)));
    layer0_outputs(1560) <= not((inputs(147)) or (inputs(124)));
    layer0_outputs(1561) <= not(inputs(120)) or (inputs(2));
    layer0_outputs(1562) <= not(inputs(14));
    layer0_outputs(1563) <= not((inputs(22)) and (inputs(179)));
    layer0_outputs(1564) <= (inputs(140)) and not (inputs(224));
    layer0_outputs(1565) <= not((inputs(208)) or (inputs(21)));
    layer0_outputs(1566) <= (inputs(28)) or (inputs(130));
    layer0_outputs(1567) <= (inputs(168)) xor (inputs(32));
    layer0_outputs(1568) <= not(inputs(35)) or (inputs(72));
    layer0_outputs(1569) <= not(inputs(211));
    layer0_outputs(1570) <= not((inputs(26)) or (inputs(21)));
    layer0_outputs(1571) <= not(inputs(56));
    layer0_outputs(1572) <= '1';
    layer0_outputs(1573) <= inputs(191);
    layer0_outputs(1574) <= not((inputs(175)) or (inputs(138)));
    layer0_outputs(1575) <= inputs(36);
    layer0_outputs(1576) <= not(inputs(116));
    layer0_outputs(1577) <= not(inputs(107)) or (inputs(51));
    layer0_outputs(1578) <= inputs(60);
    layer0_outputs(1579) <= (inputs(192)) and not (inputs(7));
    layer0_outputs(1580) <= (inputs(86)) and not (inputs(178));
    layer0_outputs(1581) <= (inputs(28)) and not (inputs(3));
    layer0_outputs(1582) <= (inputs(53)) or (inputs(38));
    layer0_outputs(1583) <= (inputs(107)) and not (inputs(209));
    layer0_outputs(1584) <= (inputs(9)) and (inputs(144));
    layer0_outputs(1585) <= (inputs(221)) xor (inputs(158));
    layer0_outputs(1586) <= not((inputs(220)) or (inputs(153)));
    layer0_outputs(1587) <= '1';
    layer0_outputs(1588) <= (inputs(255)) and not (inputs(241));
    layer0_outputs(1589) <= (inputs(253)) or (inputs(205));
    layer0_outputs(1590) <= not(inputs(11));
    layer0_outputs(1591) <= not(inputs(117)) or (inputs(64));
    layer0_outputs(1592) <= not((inputs(227)) xor (inputs(240)));
    layer0_outputs(1593) <= (inputs(142)) xor (inputs(176));
    layer0_outputs(1594) <= (inputs(147)) xor (inputs(8));
    layer0_outputs(1595) <= (inputs(92)) and (inputs(36));
    layer0_outputs(1596) <= '1';
    layer0_outputs(1597) <= not(inputs(133));
    layer0_outputs(1598) <= not((inputs(108)) or (inputs(85)));
    layer0_outputs(1599) <= not((inputs(120)) or (inputs(120)));
    layer0_outputs(1600) <= (inputs(134)) or (inputs(117));
    layer0_outputs(1601) <= not((inputs(249)) or (inputs(13)));
    layer0_outputs(1602) <= inputs(202);
    layer0_outputs(1603) <= not(inputs(173)) or (inputs(107));
    layer0_outputs(1604) <= not((inputs(66)) and (inputs(209)));
    layer0_outputs(1605) <= inputs(77);
    layer0_outputs(1606) <= (inputs(77)) or (inputs(108));
    layer0_outputs(1607) <= not((inputs(47)) and (inputs(16)));
    layer0_outputs(1608) <= not(inputs(186));
    layer0_outputs(1609) <= not(inputs(79)) or (inputs(31));
    layer0_outputs(1610) <= not((inputs(43)) or (inputs(248)));
    layer0_outputs(1611) <= not(inputs(135)) or (inputs(86));
    layer0_outputs(1612) <= not((inputs(230)) or (inputs(94)));
    layer0_outputs(1613) <= not(inputs(190));
    layer0_outputs(1614) <= (inputs(186)) and not (inputs(46));
    layer0_outputs(1615) <= (inputs(160)) and not (inputs(31));
    layer0_outputs(1616) <= inputs(98);
    layer0_outputs(1617) <= (inputs(111)) or (inputs(162));
    layer0_outputs(1618) <= (inputs(44)) and (inputs(176));
    layer0_outputs(1619) <= inputs(140);
    layer0_outputs(1620) <= not(inputs(135));
    layer0_outputs(1621) <= not(inputs(18)) or (inputs(195));
    layer0_outputs(1622) <= (inputs(148)) and not (inputs(109));
    layer0_outputs(1623) <= not(inputs(117));
    layer0_outputs(1624) <= not(inputs(48)) or (inputs(230));
    layer0_outputs(1625) <= (inputs(172)) xor (inputs(177));
    layer0_outputs(1626) <= inputs(58);
    layer0_outputs(1627) <= not(inputs(107)) or (inputs(23));
    layer0_outputs(1628) <= not(inputs(180));
    layer0_outputs(1629) <= (inputs(248)) xor (inputs(140));
    layer0_outputs(1630) <= '1';
    layer0_outputs(1631) <= not((inputs(202)) xor (inputs(171)));
    layer0_outputs(1632) <= (inputs(161)) or (inputs(103));
    layer0_outputs(1633) <= not(inputs(12));
    layer0_outputs(1634) <= not(inputs(229));
    layer0_outputs(1635) <= not((inputs(146)) xor (inputs(215)));
    layer0_outputs(1636) <= '0';
    layer0_outputs(1637) <= (inputs(101)) and not (inputs(35));
    layer0_outputs(1638) <= (inputs(73)) or (inputs(94));
    layer0_outputs(1639) <= (inputs(145)) and not (inputs(141));
    layer0_outputs(1640) <= not((inputs(42)) or (inputs(70)));
    layer0_outputs(1641) <= inputs(202);
    layer0_outputs(1642) <= (inputs(93)) or (inputs(101));
    layer0_outputs(1643) <= not((inputs(248)) xor (inputs(241)));
    layer0_outputs(1644) <= inputs(36);
    layer0_outputs(1645) <= (inputs(119)) and not (inputs(189));
    layer0_outputs(1646) <= not((inputs(195)) or (inputs(94)));
    layer0_outputs(1647) <= (inputs(187)) and (inputs(207));
    layer0_outputs(1648) <= not((inputs(210)) and (inputs(223)));
    layer0_outputs(1649) <= not((inputs(99)) and (inputs(227)));
    layer0_outputs(1650) <= not((inputs(109)) or (inputs(201)));
    layer0_outputs(1651) <= not((inputs(63)) or (inputs(92)));
    layer0_outputs(1652) <= (inputs(80)) or (inputs(47));
    layer0_outputs(1653) <= not((inputs(41)) and (inputs(74)));
    layer0_outputs(1654) <= not(inputs(45));
    layer0_outputs(1655) <= (inputs(8)) and (inputs(236));
    layer0_outputs(1656) <= '1';
    layer0_outputs(1657) <= not(inputs(142)) or (inputs(82));
    layer0_outputs(1658) <= not((inputs(54)) or (inputs(53)));
    layer0_outputs(1659) <= not((inputs(180)) xor (inputs(191)));
    layer0_outputs(1660) <= not(inputs(171));
    layer0_outputs(1661) <= (inputs(103)) or (inputs(179));
    layer0_outputs(1662) <= '1';
    layer0_outputs(1663) <= (inputs(177)) or (inputs(193));
    layer0_outputs(1664) <= not(inputs(169)) or (inputs(168));
    layer0_outputs(1665) <= inputs(236);
    layer0_outputs(1666) <= not((inputs(14)) or (inputs(216)));
    layer0_outputs(1667) <= not(inputs(151));
    layer0_outputs(1668) <= not((inputs(84)) or (inputs(208)));
    layer0_outputs(1669) <= '0';
    layer0_outputs(1670) <= (inputs(166)) xor (inputs(189));
    layer0_outputs(1671) <= (inputs(189)) and (inputs(64));
    layer0_outputs(1672) <= not(inputs(242));
    layer0_outputs(1673) <= inputs(215);
    layer0_outputs(1674) <= not(inputs(12));
    layer0_outputs(1675) <= not((inputs(201)) or (inputs(78)));
    layer0_outputs(1676) <= not((inputs(134)) xor (inputs(30)));
    layer0_outputs(1677) <= inputs(205);
    layer0_outputs(1678) <= (inputs(195)) xor (inputs(227));
    layer0_outputs(1679) <= not(inputs(82));
    layer0_outputs(1680) <= (inputs(213)) or (inputs(68));
    layer0_outputs(1681) <= not(inputs(170));
    layer0_outputs(1682) <= '0';
    layer0_outputs(1683) <= not(inputs(155)) or (inputs(99));
    layer0_outputs(1684) <= (inputs(91)) and not (inputs(146));
    layer0_outputs(1685) <= (inputs(9)) and (inputs(34));
    layer0_outputs(1686) <= not(inputs(54)) or (inputs(25));
    layer0_outputs(1687) <= not((inputs(86)) or (inputs(104)));
    layer0_outputs(1688) <= not(inputs(22));
    layer0_outputs(1689) <= (inputs(243)) or (inputs(217));
    layer0_outputs(1690) <= not(inputs(122)) or (inputs(0));
    layer0_outputs(1691) <= (inputs(59)) and not (inputs(128));
    layer0_outputs(1692) <= not(inputs(91));
    layer0_outputs(1693) <= not((inputs(244)) xor (inputs(79)));
    layer0_outputs(1694) <= (inputs(235)) and not (inputs(17));
    layer0_outputs(1695) <= inputs(133);
    layer0_outputs(1696) <= (inputs(178)) or (inputs(59));
    layer0_outputs(1697) <= (inputs(227)) and (inputs(7));
    layer0_outputs(1698) <= not((inputs(115)) xor (inputs(33)));
    layer0_outputs(1699) <= inputs(18);
    layer0_outputs(1700) <= (inputs(208)) and (inputs(17));
    layer0_outputs(1701) <= not(inputs(196)) or (inputs(232));
    layer0_outputs(1702) <= (inputs(166)) and not (inputs(235));
    layer0_outputs(1703) <= (inputs(101)) and not (inputs(88));
    layer0_outputs(1704) <= not((inputs(137)) or (inputs(234)));
    layer0_outputs(1705) <= not(inputs(179));
    layer0_outputs(1706) <= not(inputs(170)) or (inputs(110));
    layer0_outputs(1707) <= (inputs(221)) and (inputs(56));
    layer0_outputs(1708) <= (inputs(55)) and not (inputs(44));
    layer0_outputs(1709) <= not(inputs(125));
    layer0_outputs(1710) <= not(inputs(135)) or (inputs(113));
    layer0_outputs(1711) <= (inputs(35)) or (inputs(97));
    layer0_outputs(1712) <= not((inputs(177)) xor (inputs(212)));
    layer0_outputs(1713) <= inputs(198);
    layer0_outputs(1714) <= not(inputs(84)) or (inputs(97));
    layer0_outputs(1715) <= (inputs(137)) or (inputs(46));
    layer0_outputs(1716) <= not(inputs(134)) or (inputs(102));
    layer0_outputs(1717) <= (inputs(35)) or (inputs(243));
    layer0_outputs(1718) <= not((inputs(225)) xor (inputs(230)));
    layer0_outputs(1719) <= (inputs(217)) and not (inputs(10));
    layer0_outputs(1720) <= not(inputs(101));
    layer0_outputs(1721) <= not(inputs(25));
    layer0_outputs(1722) <= not(inputs(102)) or (inputs(178));
    layer0_outputs(1723) <= '1';
    layer0_outputs(1724) <= (inputs(69)) or (inputs(242));
    layer0_outputs(1725) <= '0';
    layer0_outputs(1726) <= not((inputs(57)) or (inputs(127)));
    layer0_outputs(1727) <= not(inputs(9));
    layer0_outputs(1728) <= (inputs(230)) xor (inputs(124));
    layer0_outputs(1729) <= (inputs(193)) xor (inputs(166));
    layer0_outputs(1730) <= (inputs(4)) and (inputs(244));
    layer0_outputs(1731) <= (inputs(58)) and not (inputs(132));
    layer0_outputs(1732) <= inputs(148);
    layer0_outputs(1733) <= inputs(140);
    layer0_outputs(1734) <= '1';
    layer0_outputs(1735) <= inputs(41);
    layer0_outputs(1736) <= inputs(38);
    layer0_outputs(1737) <= inputs(100);
    layer0_outputs(1738) <= not(inputs(184));
    layer0_outputs(1739) <= (inputs(113)) and not (inputs(16));
    layer0_outputs(1740) <= not(inputs(188));
    layer0_outputs(1741) <= (inputs(86)) and not (inputs(50));
    layer0_outputs(1742) <= (inputs(88)) and not (inputs(182));
    layer0_outputs(1743) <= (inputs(82)) or (inputs(153));
    layer0_outputs(1744) <= '0';
    layer0_outputs(1745) <= inputs(207);
    layer0_outputs(1746) <= (inputs(93)) or (inputs(85));
    layer0_outputs(1747) <= not((inputs(109)) xor (inputs(158)));
    layer0_outputs(1748) <= not(inputs(77));
    layer0_outputs(1749) <= not((inputs(53)) or (inputs(148)));
    layer0_outputs(1750) <= not(inputs(205));
    layer0_outputs(1751) <= '1';
    layer0_outputs(1752) <= inputs(99);
    layer0_outputs(1753) <= (inputs(3)) xor (inputs(238));
    layer0_outputs(1754) <= not((inputs(183)) or (inputs(28)));
    layer0_outputs(1755) <= not((inputs(56)) and (inputs(57)));
    layer0_outputs(1756) <= (inputs(194)) and not (inputs(235));
    layer0_outputs(1757) <= (inputs(34)) or (inputs(108));
    layer0_outputs(1758) <= inputs(249);
    layer0_outputs(1759) <= inputs(234);
    layer0_outputs(1760) <= not((inputs(149)) or (inputs(22)));
    layer0_outputs(1761) <= inputs(52);
    layer0_outputs(1762) <= (inputs(189)) or (inputs(201));
    layer0_outputs(1763) <= '1';
    layer0_outputs(1764) <= '1';
    layer0_outputs(1765) <= not((inputs(170)) or (inputs(117)));
    layer0_outputs(1766) <= not(inputs(248)) or (inputs(79));
    layer0_outputs(1767) <= (inputs(3)) and not (inputs(53));
    layer0_outputs(1768) <= not((inputs(13)) xor (inputs(65)));
    layer0_outputs(1769) <= (inputs(86)) or (inputs(110));
    layer0_outputs(1770) <= not(inputs(131));
    layer0_outputs(1771) <= not((inputs(236)) and (inputs(206)));
    layer0_outputs(1772) <= not(inputs(186));
    layer0_outputs(1773) <= not(inputs(157));
    layer0_outputs(1774) <= not((inputs(142)) and (inputs(173)));
    layer0_outputs(1775) <= not(inputs(102));
    layer0_outputs(1776) <= not((inputs(203)) or (inputs(202)));
    layer0_outputs(1777) <= not(inputs(27));
    layer0_outputs(1778) <= (inputs(157)) or (inputs(165));
    layer0_outputs(1779) <= (inputs(208)) and (inputs(96));
    layer0_outputs(1780) <= (inputs(237)) or (inputs(233));
    layer0_outputs(1781) <= (inputs(29)) and (inputs(62));
    layer0_outputs(1782) <= (inputs(119)) and not (inputs(191));
    layer0_outputs(1783) <= not((inputs(219)) xor (inputs(250)));
    layer0_outputs(1784) <= (inputs(213)) xor (inputs(95));
    layer0_outputs(1785) <= inputs(205);
    layer0_outputs(1786) <= not(inputs(239));
    layer0_outputs(1787) <= (inputs(36)) and not (inputs(233));
    layer0_outputs(1788) <= (inputs(90)) or (inputs(220));
    layer0_outputs(1789) <= (inputs(144)) and not (inputs(149));
    layer0_outputs(1790) <= inputs(119);
    layer0_outputs(1791) <= not(inputs(179)) or (inputs(17));
    layer0_outputs(1792) <= not(inputs(80));
    layer0_outputs(1793) <= not(inputs(124));
    layer0_outputs(1794) <= (inputs(212)) and not (inputs(244));
    layer0_outputs(1795) <= (inputs(15)) xor (inputs(240));
    layer0_outputs(1796) <= (inputs(26)) or (inputs(184));
    layer0_outputs(1797) <= not(inputs(102)) or (inputs(75));
    layer0_outputs(1798) <= not(inputs(8)) or (inputs(211));
    layer0_outputs(1799) <= not(inputs(250));
    layer0_outputs(1800) <= not((inputs(239)) and (inputs(7)));
    layer0_outputs(1801) <= not((inputs(244)) xor (inputs(78)));
    layer0_outputs(1802) <= (inputs(112)) and (inputs(170));
    layer0_outputs(1803) <= (inputs(97)) and (inputs(188));
    layer0_outputs(1804) <= (inputs(20)) or (inputs(167));
    layer0_outputs(1805) <= (inputs(186)) or (inputs(26));
    layer0_outputs(1806) <= (inputs(173)) or (inputs(71));
    layer0_outputs(1807) <= not((inputs(85)) or (inputs(220)));
    layer0_outputs(1808) <= (inputs(68)) or (inputs(40));
    layer0_outputs(1809) <= (inputs(141)) and not (inputs(64));
    layer0_outputs(1810) <= not(inputs(113)) or (inputs(194));
    layer0_outputs(1811) <= '0';
    layer0_outputs(1812) <= inputs(135);
    layer0_outputs(1813) <= not(inputs(205));
    layer0_outputs(1814) <= not((inputs(216)) or (inputs(88)));
    layer0_outputs(1815) <= not(inputs(203));
    layer0_outputs(1816) <= (inputs(253)) and not (inputs(7));
    layer0_outputs(1817) <= (inputs(74)) xor (inputs(196));
    layer0_outputs(1818) <= not((inputs(235)) xor (inputs(214)));
    layer0_outputs(1819) <= not((inputs(63)) or (inputs(207)));
    layer0_outputs(1820) <= not(inputs(149)) or (inputs(69));
    layer0_outputs(1821) <= (inputs(219)) xor (inputs(238));
    layer0_outputs(1822) <= (inputs(121)) or (inputs(220));
    layer0_outputs(1823) <= not(inputs(136));
    layer0_outputs(1824) <= (inputs(79)) and (inputs(99));
    layer0_outputs(1825) <= not((inputs(146)) xor (inputs(9)));
    layer0_outputs(1826) <= not((inputs(28)) and (inputs(128)));
    layer0_outputs(1827) <= not((inputs(137)) or (inputs(206)));
    layer0_outputs(1828) <= not((inputs(25)) or (inputs(167)));
    layer0_outputs(1829) <= not(inputs(12));
    layer0_outputs(1830) <= (inputs(49)) and not (inputs(65));
    layer0_outputs(1831) <= not(inputs(230));
    layer0_outputs(1832) <= not(inputs(45)) or (inputs(13));
    layer0_outputs(1833) <= inputs(94);
    layer0_outputs(1834) <= not((inputs(251)) and (inputs(242)));
    layer0_outputs(1835) <= not((inputs(228)) xor (inputs(242)));
    layer0_outputs(1836) <= inputs(28);
    layer0_outputs(1837) <= not(inputs(177));
    layer0_outputs(1838) <= (inputs(235)) and not (inputs(41));
    layer0_outputs(1839) <= not(inputs(204)) or (inputs(236));
    layer0_outputs(1840) <= (inputs(170)) xor (inputs(155));
    layer0_outputs(1841) <= '1';
    layer0_outputs(1842) <= (inputs(26)) and (inputs(25));
    layer0_outputs(1843) <= not((inputs(126)) or (inputs(106)));
    layer0_outputs(1844) <= (inputs(58)) xor (inputs(47));
    layer0_outputs(1845) <= inputs(46);
    layer0_outputs(1846) <= (inputs(40)) or (inputs(156));
    layer0_outputs(1847) <= not((inputs(197)) or (inputs(162)));
    layer0_outputs(1848) <= not((inputs(189)) or (inputs(239)));
    layer0_outputs(1849) <= not((inputs(113)) and (inputs(252)));
    layer0_outputs(1850) <= (inputs(72)) and not (inputs(254));
    layer0_outputs(1851) <= not((inputs(104)) xor (inputs(72)));
    layer0_outputs(1852) <= inputs(188);
    layer0_outputs(1853) <= not(inputs(198)) or (inputs(240));
    layer0_outputs(1854) <= inputs(36);
    layer0_outputs(1855) <= inputs(13);
    layer0_outputs(1856) <= (inputs(235)) and (inputs(128));
    layer0_outputs(1857) <= '1';
    layer0_outputs(1858) <= inputs(105);
    layer0_outputs(1859) <= not((inputs(13)) or (inputs(135)));
    layer0_outputs(1860) <= (inputs(156)) and not (inputs(110));
    layer0_outputs(1861) <= inputs(71);
    layer0_outputs(1862) <= not((inputs(72)) xor (inputs(14)));
    layer0_outputs(1863) <= not((inputs(228)) or (inputs(90)));
    layer0_outputs(1864) <= (inputs(77)) and not (inputs(2));
    layer0_outputs(1865) <= (inputs(239)) and not (inputs(1));
    layer0_outputs(1866) <= (inputs(119)) or (inputs(253));
    layer0_outputs(1867) <= (inputs(113)) xor (inputs(127));
    layer0_outputs(1868) <= inputs(139);
    layer0_outputs(1869) <= (inputs(254)) and (inputs(215));
    layer0_outputs(1870) <= not(inputs(114)) or (inputs(245));
    layer0_outputs(1871) <= (inputs(133)) or (inputs(158));
    layer0_outputs(1872) <= not((inputs(33)) xor (inputs(212)));
    layer0_outputs(1873) <= not((inputs(142)) xor (inputs(198)));
    layer0_outputs(1874) <= (inputs(147)) and not (inputs(220));
    layer0_outputs(1875) <= not((inputs(242)) and (inputs(10)));
    layer0_outputs(1876) <= (inputs(7)) and not (inputs(246));
    layer0_outputs(1877) <= not(inputs(189));
    layer0_outputs(1878) <= not((inputs(102)) or (inputs(236)));
    layer0_outputs(1879) <= inputs(101);
    layer0_outputs(1880) <= inputs(249);
    layer0_outputs(1881) <= (inputs(82)) or (inputs(184));
    layer0_outputs(1882) <= (inputs(98)) xor (inputs(177));
    layer0_outputs(1883) <= (inputs(137)) or (inputs(82));
    layer0_outputs(1884) <= not((inputs(228)) and (inputs(141)));
    layer0_outputs(1885) <= not((inputs(144)) xor (inputs(4)));
    layer0_outputs(1886) <= (inputs(171)) and (inputs(171));
    layer0_outputs(1887) <= inputs(117);
    layer0_outputs(1888) <= not(inputs(71)) or (inputs(186));
    layer0_outputs(1889) <= inputs(69);
    layer0_outputs(1890) <= inputs(63);
    layer0_outputs(1891) <= not(inputs(123)) or (inputs(67));
    layer0_outputs(1892) <= not((inputs(95)) and (inputs(180)));
    layer0_outputs(1893) <= (inputs(11)) xor (inputs(179));
    layer0_outputs(1894) <= not((inputs(141)) and (inputs(229)));
    layer0_outputs(1895) <= inputs(118);
    layer0_outputs(1896) <= not((inputs(181)) xor (inputs(211)));
    layer0_outputs(1897) <= not(inputs(125)) or (inputs(67));
    layer0_outputs(1898) <= not(inputs(105));
    layer0_outputs(1899) <= (inputs(85)) or (inputs(100));
    layer0_outputs(1900) <= not((inputs(95)) xor (inputs(187)));
    layer0_outputs(1901) <= (inputs(21)) and not (inputs(162));
    layer0_outputs(1902) <= not(inputs(16));
    layer0_outputs(1903) <= not((inputs(137)) or (inputs(232)));
    layer0_outputs(1904) <= not((inputs(26)) xor (inputs(87)));
    layer0_outputs(1905) <= inputs(87);
    layer0_outputs(1906) <= not(inputs(139));
    layer0_outputs(1907) <= inputs(227);
    layer0_outputs(1908) <= not(inputs(225)) or (inputs(52));
    layer0_outputs(1909) <= (inputs(70)) and (inputs(87));
    layer0_outputs(1910) <= (inputs(101)) and not (inputs(83));
    layer0_outputs(1911) <= not(inputs(127));
    layer0_outputs(1912) <= '0';
    layer0_outputs(1913) <= (inputs(48)) and not (inputs(92));
    layer0_outputs(1914) <= inputs(236);
    layer0_outputs(1915) <= not(inputs(30));
    layer0_outputs(1916) <= (inputs(220)) or (inputs(79));
    layer0_outputs(1917) <= inputs(238);
    layer0_outputs(1918) <= (inputs(129)) xor (inputs(232));
    layer0_outputs(1919) <= not(inputs(68));
    layer0_outputs(1920) <= not(inputs(165)) or (inputs(63));
    layer0_outputs(1921) <= (inputs(189)) and not (inputs(27));
    layer0_outputs(1922) <= (inputs(125)) or (inputs(100));
    layer0_outputs(1923) <= not(inputs(159)) or (inputs(194));
    layer0_outputs(1924) <= not(inputs(16));
    layer0_outputs(1925) <= (inputs(81)) or (inputs(189));
    layer0_outputs(1926) <= not(inputs(94)) or (inputs(19));
    layer0_outputs(1927) <= inputs(242);
    layer0_outputs(1928) <= not(inputs(117));
    layer0_outputs(1929) <= (inputs(190)) and not (inputs(129));
    layer0_outputs(1930) <= (inputs(44)) and not (inputs(161));
    layer0_outputs(1931) <= (inputs(9)) and not (inputs(72));
    layer0_outputs(1932) <= inputs(254);
    layer0_outputs(1933) <= not((inputs(38)) xor (inputs(59)));
    layer0_outputs(1934) <= (inputs(128)) xor (inputs(148));
    layer0_outputs(1935) <= (inputs(27)) and not (inputs(229));
    layer0_outputs(1936) <= (inputs(217)) or (inputs(38));
    layer0_outputs(1937) <= not((inputs(59)) or (inputs(11)));
    layer0_outputs(1938) <= inputs(101);
    layer0_outputs(1939) <= (inputs(124)) and not (inputs(225));
    layer0_outputs(1940) <= (inputs(107)) and not (inputs(35));
    layer0_outputs(1941) <= (inputs(182)) or (inputs(185));
    layer0_outputs(1942) <= inputs(251);
    layer0_outputs(1943) <= (inputs(167)) or (inputs(159));
    layer0_outputs(1944) <= (inputs(75)) and not (inputs(29));
    layer0_outputs(1945) <= not(inputs(125));
    layer0_outputs(1946) <= not((inputs(40)) xor (inputs(35)));
    layer0_outputs(1947) <= (inputs(103)) and not (inputs(233));
    layer0_outputs(1948) <= not(inputs(175)) or (inputs(227));
    layer0_outputs(1949) <= inputs(163);
    layer0_outputs(1950) <= '1';
    layer0_outputs(1951) <= not((inputs(16)) and (inputs(138)));
    layer0_outputs(1952) <= not((inputs(233)) xor (inputs(195)));
    layer0_outputs(1953) <= inputs(236);
    layer0_outputs(1954) <= (inputs(6)) and (inputs(17));
    layer0_outputs(1955) <= not(inputs(34));
    layer0_outputs(1956) <= (inputs(35)) and not (inputs(1));
    layer0_outputs(1957) <= (inputs(253)) and not (inputs(24));
    layer0_outputs(1958) <= not((inputs(178)) or (inputs(26)));
    layer0_outputs(1959) <= (inputs(227)) or (inputs(87));
    layer0_outputs(1960) <= (inputs(204)) and (inputs(62));
    layer0_outputs(1961) <= not(inputs(120)) or (inputs(24));
    layer0_outputs(1962) <= not(inputs(152));
    layer0_outputs(1963) <= not((inputs(149)) xor (inputs(164)));
    layer0_outputs(1964) <= (inputs(45)) and not (inputs(6));
    layer0_outputs(1965) <= not(inputs(210)) or (inputs(246));
    layer0_outputs(1966) <= not(inputs(251));
    layer0_outputs(1967) <= not(inputs(42));
    layer0_outputs(1968) <= '1';
    layer0_outputs(1969) <= inputs(245);
    layer0_outputs(1970) <= not(inputs(63));
    layer0_outputs(1971) <= not((inputs(24)) or (inputs(172)));
    layer0_outputs(1972) <= not((inputs(139)) or (inputs(171)));
    layer0_outputs(1973) <= not(inputs(221)) or (inputs(7));
    layer0_outputs(1974) <= not((inputs(248)) or (inputs(108)));
    layer0_outputs(1975) <= '0';
    layer0_outputs(1976) <= not(inputs(141));
    layer0_outputs(1977) <= not((inputs(205)) and (inputs(236)));
    layer0_outputs(1978) <= not(inputs(180));
    layer0_outputs(1979) <= not(inputs(75));
    layer0_outputs(1980) <= not(inputs(42)) or (inputs(203));
    layer0_outputs(1981) <= (inputs(235)) and not (inputs(40));
    layer0_outputs(1982) <= (inputs(25)) or (inputs(39));
    layer0_outputs(1983) <= not(inputs(145)) or (inputs(68));
    layer0_outputs(1984) <= not(inputs(180));
    layer0_outputs(1985) <= (inputs(39)) and not (inputs(129));
    layer0_outputs(1986) <= not(inputs(247)) or (inputs(1));
    layer0_outputs(1987) <= not((inputs(137)) xor (inputs(34)));
    layer0_outputs(1988) <= (inputs(145)) and not (inputs(64));
    layer0_outputs(1989) <= (inputs(152)) and not (inputs(88));
    layer0_outputs(1990) <= not((inputs(27)) or (inputs(172)));
    layer0_outputs(1991) <= inputs(68);
    layer0_outputs(1992) <= inputs(189);
    layer0_outputs(1993) <= (inputs(105)) and not (inputs(20));
    layer0_outputs(1994) <= not((inputs(190)) xor (inputs(180)));
    layer0_outputs(1995) <= (inputs(49)) and not (inputs(177));
    layer0_outputs(1996) <= inputs(74);
    layer0_outputs(1997) <= inputs(105);
    layer0_outputs(1998) <= not(inputs(20)) or (inputs(115));
    layer0_outputs(1999) <= not((inputs(174)) xor (inputs(92)));
    layer0_outputs(2000) <= (inputs(87)) or (inputs(103));
    layer0_outputs(2001) <= not((inputs(245)) xor (inputs(15)));
    layer0_outputs(2002) <= inputs(21);
    layer0_outputs(2003) <= (inputs(56)) and not (inputs(139));
    layer0_outputs(2004) <= not((inputs(104)) xor (inputs(96)));
    layer0_outputs(2005) <= inputs(100);
    layer0_outputs(2006) <= inputs(214);
    layer0_outputs(2007) <= '1';
    layer0_outputs(2008) <= not(inputs(53)) or (inputs(122));
    layer0_outputs(2009) <= not(inputs(99));
    layer0_outputs(2010) <= (inputs(201)) and not (inputs(242));
    layer0_outputs(2011) <= (inputs(118)) and not (inputs(114));
    layer0_outputs(2012) <= '0';
    layer0_outputs(2013) <= not(inputs(233));
    layer0_outputs(2014) <= not((inputs(157)) or (inputs(223)));
    layer0_outputs(2015) <= not(inputs(145));
    layer0_outputs(2016) <= not((inputs(252)) and (inputs(226)));
    layer0_outputs(2017) <= inputs(57);
    layer0_outputs(2018) <= not((inputs(119)) or (inputs(64)));
    layer0_outputs(2019) <= inputs(86);
    layer0_outputs(2020) <= inputs(104);
    layer0_outputs(2021) <= not(inputs(183));
    layer0_outputs(2022) <= (inputs(90)) and not (inputs(39));
    layer0_outputs(2023) <= not((inputs(142)) or (inputs(39)));
    layer0_outputs(2024) <= not((inputs(182)) or (inputs(25)));
    layer0_outputs(2025) <= inputs(76);
    layer0_outputs(2026) <= not((inputs(75)) xor (inputs(67)));
    layer0_outputs(2027) <= inputs(170);
    layer0_outputs(2028) <= (inputs(173)) and (inputs(62));
    layer0_outputs(2029) <= not((inputs(114)) xor (inputs(243)));
    layer0_outputs(2030) <= not(inputs(215));
    layer0_outputs(2031) <= inputs(243);
    layer0_outputs(2032) <= not(inputs(143)) or (inputs(226));
    layer0_outputs(2033) <= not(inputs(119));
    layer0_outputs(2034) <= not((inputs(59)) xor (inputs(203)));
    layer0_outputs(2035) <= not(inputs(150));
    layer0_outputs(2036) <= not((inputs(40)) and (inputs(114)));
    layer0_outputs(2037) <= (inputs(232)) and not (inputs(240));
    layer0_outputs(2038) <= not((inputs(227)) xor (inputs(155)));
    layer0_outputs(2039) <= inputs(108);
    layer0_outputs(2040) <= (inputs(221)) xor (inputs(111));
    layer0_outputs(2041) <= (inputs(179)) and not (inputs(233));
    layer0_outputs(2042) <= not((inputs(241)) xor (inputs(210)));
    layer0_outputs(2043) <= not((inputs(0)) or (inputs(152)));
    layer0_outputs(2044) <= not(inputs(3)) or (inputs(222));
    layer0_outputs(2045) <= (inputs(194)) and (inputs(161));
    layer0_outputs(2046) <= inputs(116);
    layer0_outputs(2047) <= not((inputs(44)) xor (inputs(113)));
    layer0_outputs(2048) <= not(inputs(233));
    layer0_outputs(2049) <= inputs(126);
    layer0_outputs(2050) <= not((inputs(140)) or (inputs(53)));
    layer0_outputs(2051) <= (inputs(27)) and not (inputs(220));
    layer0_outputs(2052) <= not((inputs(174)) and (inputs(59)));
    layer0_outputs(2053) <= not(inputs(158));
    layer0_outputs(2054) <= not(inputs(89));
    layer0_outputs(2055) <= inputs(75);
    layer0_outputs(2056) <= not(inputs(60));
    layer0_outputs(2057) <= (inputs(72)) and not (inputs(229));
    layer0_outputs(2058) <= not(inputs(142)) or (inputs(71));
    layer0_outputs(2059) <= (inputs(118)) or (inputs(80));
    layer0_outputs(2060) <= '0';
    layer0_outputs(2061) <= (inputs(238)) and not (inputs(251));
    layer0_outputs(2062) <= not(inputs(109));
    layer0_outputs(2063) <= not((inputs(237)) and (inputs(16)));
    layer0_outputs(2064) <= inputs(26);
    layer0_outputs(2065) <= (inputs(228)) or (inputs(8));
    layer0_outputs(2066) <= not((inputs(47)) xor (inputs(141)));
    layer0_outputs(2067) <= (inputs(52)) or (inputs(194));
    layer0_outputs(2068) <= inputs(19);
    layer0_outputs(2069) <= (inputs(33)) xor (inputs(176));
    layer0_outputs(2070) <= '1';
    layer0_outputs(2071) <= inputs(65);
    layer0_outputs(2072) <= not(inputs(98)) or (inputs(198));
    layer0_outputs(2073) <= inputs(4);
    layer0_outputs(2074) <= not((inputs(226)) and (inputs(221)));
    layer0_outputs(2075) <= (inputs(135)) or (inputs(27));
    layer0_outputs(2076) <= '0';
    layer0_outputs(2077) <= not((inputs(221)) or (inputs(32)));
    layer0_outputs(2078) <= not(inputs(87));
    layer0_outputs(2079) <= not((inputs(6)) and (inputs(145)));
    layer0_outputs(2080) <= not((inputs(171)) or (inputs(197)));
    layer0_outputs(2081) <= (inputs(77)) and (inputs(170));
    layer0_outputs(2082) <= (inputs(166)) xor (inputs(5));
    layer0_outputs(2083) <= (inputs(228)) and not (inputs(78));
    layer0_outputs(2084) <= not((inputs(250)) xor (inputs(191)));
    layer0_outputs(2085) <= inputs(137);
    layer0_outputs(2086) <= '1';
    layer0_outputs(2087) <= not((inputs(252)) and (inputs(20)));
    layer0_outputs(2088) <= (inputs(231)) and not (inputs(47));
    layer0_outputs(2089) <= (inputs(85)) or (inputs(84));
    layer0_outputs(2090) <= (inputs(244)) and not (inputs(102));
    layer0_outputs(2091) <= not(inputs(181));
    layer0_outputs(2092) <= (inputs(107)) and not (inputs(194));
    layer0_outputs(2093) <= not((inputs(38)) or (inputs(203)));
    layer0_outputs(2094) <= not(inputs(193));
    layer0_outputs(2095) <= not(inputs(125));
    layer0_outputs(2096) <= (inputs(142)) or (inputs(235));
    layer0_outputs(2097) <= (inputs(0)) or (inputs(99));
    layer0_outputs(2098) <= not((inputs(36)) or (inputs(239)));
    layer0_outputs(2099) <= (inputs(118)) and not (inputs(175));
    layer0_outputs(2100) <= (inputs(237)) and (inputs(114));
    layer0_outputs(2101) <= (inputs(190)) and not (inputs(221));
    layer0_outputs(2102) <= (inputs(37)) or (inputs(180));
    layer0_outputs(2103) <= not((inputs(155)) xor (inputs(36)));
    layer0_outputs(2104) <= (inputs(90)) or (inputs(107));
    layer0_outputs(2105) <= not((inputs(0)) or (inputs(239)));
    layer0_outputs(2106) <= (inputs(94)) or (inputs(215));
    layer0_outputs(2107) <= not(inputs(186)) or (inputs(195));
    layer0_outputs(2108) <= not((inputs(92)) xor (inputs(186)));
    layer0_outputs(2109) <= inputs(135);
    layer0_outputs(2110) <= not((inputs(61)) or (inputs(149)));
    layer0_outputs(2111) <= inputs(88);
    layer0_outputs(2112) <= not((inputs(136)) xor (inputs(155)));
    layer0_outputs(2113) <= not(inputs(107)) or (inputs(163));
    layer0_outputs(2114) <= not(inputs(113)) or (inputs(179));
    layer0_outputs(2115) <= not((inputs(139)) xor (inputs(28)));
    layer0_outputs(2116) <= inputs(70);
    layer0_outputs(2117) <= not((inputs(51)) or (inputs(154)));
    layer0_outputs(2118) <= (inputs(28)) xor (inputs(48));
    layer0_outputs(2119) <= (inputs(146)) and not (inputs(221));
    layer0_outputs(2120) <= not((inputs(3)) or (inputs(181)));
    layer0_outputs(2121) <= not((inputs(75)) xor (inputs(90)));
    layer0_outputs(2122) <= not((inputs(11)) or (inputs(250)));
    layer0_outputs(2123) <= not((inputs(50)) or (inputs(168)));
    layer0_outputs(2124) <= not(inputs(82));
    layer0_outputs(2125) <= (inputs(199)) and (inputs(32));
    layer0_outputs(2126) <= not((inputs(206)) or (inputs(39)));
    layer0_outputs(2127) <= not(inputs(231)) or (inputs(24));
    layer0_outputs(2128) <= (inputs(87)) and not (inputs(230));
    layer0_outputs(2129) <= (inputs(234)) and not (inputs(2));
    layer0_outputs(2130) <= not(inputs(73));
    layer0_outputs(2131) <= (inputs(150)) xor (inputs(156));
    layer0_outputs(2132) <= inputs(255);
    layer0_outputs(2133) <= not((inputs(44)) or (inputs(172)));
    layer0_outputs(2134) <= (inputs(171)) and not (inputs(218));
    layer0_outputs(2135) <= not(inputs(187));
    layer0_outputs(2136) <= (inputs(234)) and not (inputs(111));
    layer0_outputs(2137) <= inputs(214);
    layer0_outputs(2138) <= not((inputs(144)) xor (inputs(249)));
    layer0_outputs(2139) <= not((inputs(249)) xor (inputs(70)));
    layer0_outputs(2140) <= inputs(171);
    layer0_outputs(2141) <= (inputs(232)) and not (inputs(81));
    layer0_outputs(2142) <= not((inputs(83)) or (inputs(246)));
    layer0_outputs(2143) <= (inputs(144)) and (inputs(65));
    layer0_outputs(2144) <= not((inputs(128)) or (inputs(230)));
    layer0_outputs(2145) <= not(inputs(157)) or (inputs(213));
    layer0_outputs(2146) <= '1';
    layer0_outputs(2147) <= '0';
    layer0_outputs(2148) <= not(inputs(207)) or (inputs(71));
    layer0_outputs(2149) <= (inputs(179)) and not (inputs(201));
    layer0_outputs(2150) <= (inputs(57)) or (inputs(117));
    layer0_outputs(2151) <= (inputs(165)) and not (inputs(209));
    layer0_outputs(2152) <= '1';
    layer0_outputs(2153) <= inputs(131);
    layer0_outputs(2154) <= not((inputs(44)) or (inputs(133)));
    layer0_outputs(2155) <= (inputs(241)) and (inputs(216));
    layer0_outputs(2156) <= inputs(211);
    layer0_outputs(2157) <= not((inputs(181)) xor (inputs(111)));
    layer0_outputs(2158) <= (inputs(21)) or (inputs(56));
    layer0_outputs(2159) <= not((inputs(155)) and (inputs(60)));
    layer0_outputs(2160) <= (inputs(152)) and not (inputs(22));
    layer0_outputs(2161) <= not(inputs(107));
    layer0_outputs(2162) <= not((inputs(92)) xor (inputs(161)));
    layer0_outputs(2163) <= (inputs(189)) xor (inputs(29));
    layer0_outputs(2164) <= (inputs(127)) or (inputs(170));
    layer0_outputs(2165) <= not(inputs(54)) or (inputs(127));
    layer0_outputs(2166) <= inputs(230);
    layer0_outputs(2167) <= not(inputs(101));
    layer0_outputs(2168) <= (inputs(21)) and (inputs(169));
    layer0_outputs(2169) <= inputs(36);
    layer0_outputs(2170) <= (inputs(236)) or (inputs(237));
    layer0_outputs(2171) <= not(inputs(120)) or (inputs(125));
    layer0_outputs(2172) <= '0';
    layer0_outputs(2173) <= (inputs(69)) xor (inputs(202));
    layer0_outputs(2174) <= (inputs(28)) or (inputs(48));
    layer0_outputs(2175) <= (inputs(181)) or (inputs(119));
    layer0_outputs(2176) <= (inputs(15)) or (inputs(79));
    layer0_outputs(2177) <= (inputs(185)) and not (inputs(84));
    layer0_outputs(2178) <= not((inputs(87)) xor (inputs(189)));
    layer0_outputs(2179) <= '0';
    layer0_outputs(2180) <= (inputs(46)) or (inputs(223));
    layer0_outputs(2181) <= inputs(92);
    layer0_outputs(2182) <= not((inputs(80)) and (inputs(112)));
    layer0_outputs(2183) <= inputs(147);
    layer0_outputs(2184) <= not(inputs(51)) or (inputs(150));
    layer0_outputs(2185) <= not(inputs(102));
    layer0_outputs(2186) <= not(inputs(72)) or (inputs(147));
    layer0_outputs(2187) <= (inputs(153)) and not (inputs(212));
    layer0_outputs(2188) <= not((inputs(148)) or (inputs(11)));
    layer0_outputs(2189) <= (inputs(18)) or (inputs(71));
    layer0_outputs(2190) <= '1';
    layer0_outputs(2191) <= not((inputs(53)) or (inputs(61)));
    layer0_outputs(2192) <= not(inputs(137));
    layer0_outputs(2193) <= not(inputs(95)) or (inputs(128));
    layer0_outputs(2194) <= (inputs(40)) or (inputs(49));
    layer0_outputs(2195) <= (inputs(16)) or (inputs(155));
    layer0_outputs(2196) <= inputs(100);
    layer0_outputs(2197) <= not((inputs(7)) xor (inputs(248)));
    layer0_outputs(2198) <= '1';
    layer0_outputs(2199) <= inputs(100);
    layer0_outputs(2200) <= inputs(135);
    layer0_outputs(2201) <= inputs(77);
    layer0_outputs(2202) <= not(inputs(176)) or (inputs(19));
    layer0_outputs(2203) <= not((inputs(52)) or (inputs(203)));
    layer0_outputs(2204) <= inputs(39);
    layer0_outputs(2205) <= inputs(183);
    layer0_outputs(2206) <= '0';
    layer0_outputs(2207) <= '1';
    layer0_outputs(2208) <= not((inputs(230)) or (inputs(154)));
    layer0_outputs(2209) <= inputs(172);
    layer0_outputs(2210) <= '1';
    layer0_outputs(2211) <= (inputs(20)) xor (inputs(167));
    layer0_outputs(2212) <= inputs(101);
    layer0_outputs(2213) <= inputs(151);
    layer0_outputs(2214) <= not((inputs(212)) or (inputs(103)));
    layer0_outputs(2215) <= inputs(183);
    layer0_outputs(2216) <= (inputs(76)) and not (inputs(192));
    layer0_outputs(2217) <= (inputs(98)) or (inputs(64));
    layer0_outputs(2218) <= inputs(20);
    layer0_outputs(2219) <= (inputs(53)) and not (inputs(3));
    layer0_outputs(2220) <= (inputs(34)) xor (inputs(230));
    layer0_outputs(2221) <= (inputs(45)) and not (inputs(50));
    layer0_outputs(2222) <= (inputs(51)) xor (inputs(41));
    layer0_outputs(2223) <= not(inputs(170)) or (inputs(155));
    layer0_outputs(2224) <= not((inputs(140)) or (inputs(139)));
    layer0_outputs(2225) <= (inputs(139)) xor (inputs(120));
    layer0_outputs(2226) <= not((inputs(136)) and (inputs(139)));
    layer0_outputs(2227) <= not((inputs(2)) xor (inputs(214)));
    layer0_outputs(2228) <= not(inputs(51));
    layer0_outputs(2229) <= (inputs(151)) or (inputs(13));
    layer0_outputs(2230) <= not(inputs(102));
    layer0_outputs(2231) <= (inputs(168)) and not (inputs(227));
    layer0_outputs(2232) <= (inputs(133)) or (inputs(180));
    layer0_outputs(2233) <= (inputs(140)) and not (inputs(237));
    layer0_outputs(2234) <= (inputs(97)) or (inputs(144));
    layer0_outputs(2235) <= (inputs(163)) and not (inputs(249));
    layer0_outputs(2236) <= not((inputs(40)) or (inputs(173)));
    layer0_outputs(2237) <= not((inputs(229)) or (inputs(170)));
    layer0_outputs(2238) <= inputs(13);
    layer0_outputs(2239) <= not((inputs(46)) or (inputs(166)));
    layer0_outputs(2240) <= (inputs(141)) and not (inputs(144));
    layer0_outputs(2241) <= (inputs(242)) or (inputs(201));
    layer0_outputs(2242) <= (inputs(196)) and (inputs(236));
    layer0_outputs(2243) <= '1';
    layer0_outputs(2244) <= not((inputs(80)) and (inputs(229)));
    layer0_outputs(2245) <= not((inputs(181)) or (inputs(20)));
    layer0_outputs(2246) <= inputs(50);
    layer0_outputs(2247) <= not(inputs(46)) or (inputs(207));
    layer0_outputs(2248) <= inputs(164);
    layer0_outputs(2249) <= not(inputs(180));
    layer0_outputs(2250) <= not(inputs(238));
    layer0_outputs(2251) <= not(inputs(86)) or (inputs(27));
    layer0_outputs(2252) <= (inputs(63)) and not (inputs(218));
    layer0_outputs(2253) <= not(inputs(120));
    layer0_outputs(2254) <= (inputs(22)) and not (inputs(82));
    layer0_outputs(2255) <= (inputs(59)) or (inputs(214));
    layer0_outputs(2256) <= not((inputs(80)) or (inputs(121)));
    layer0_outputs(2257) <= not(inputs(53)) or (inputs(208));
    layer0_outputs(2258) <= (inputs(112)) or (inputs(166));
    layer0_outputs(2259) <= not(inputs(196));
    layer0_outputs(2260) <= (inputs(48)) or (inputs(56));
    layer0_outputs(2261) <= inputs(214);
    layer0_outputs(2262) <= not(inputs(87));
    layer0_outputs(2263) <= not((inputs(138)) or (inputs(231)));
    layer0_outputs(2264) <= not((inputs(44)) and (inputs(26)));
    layer0_outputs(2265) <= not(inputs(222)) or (inputs(146));
    layer0_outputs(2266) <= not(inputs(165));
    layer0_outputs(2267) <= not(inputs(37));
    layer0_outputs(2268) <= inputs(237);
    layer0_outputs(2269) <= not(inputs(151));
    layer0_outputs(2270) <= not(inputs(150)) or (inputs(27));
    layer0_outputs(2271) <= not(inputs(245)) or (inputs(33));
    layer0_outputs(2272) <= inputs(172);
    layer0_outputs(2273) <= (inputs(118)) and (inputs(82));
    layer0_outputs(2274) <= (inputs(186)) or (inputs(170));
    layer0_outputs(2275) <= (inputs(172)) and not (inputs(15));
    layer0_outputs(2276) <= inputs(100);
    layer0_outputs(2277) <= inputs(59);
    layer0_outputs(2278) <= (inputs(228)) or (inputs(81));
    layer0_outputs(2279) <= not(inputs(95)) or (inputs(202));
    layer0_outputs(2280) <= (inputs(17)) and not (inputs(248));
    layer0_outputs(2281) <= not(inputs(126));
    layer0_outputs(2282) <= (inputs(224)) or (inputs(63));
    layer0_outputs(2283) <= not((inputs(50)) xor (inputs(45)));
    layer0_outputs(2284) <= inputs(113);
    layer0_outputs(2285) <= (inputs(128)) and (inputs(7));
    layer0_outputs(2286) <= not((inputs(124)) or (inputs(167)));
    layer0_outputs(2287) <= not((inputs(171)) or (inputs(188)));
    layer0_outputs(2288) <= not((inputs(124)) or (inputs(42)));
    layer0_outputs(2289) <= (inputs(82)) and not (inputs(126));
    layer0_outputs(2290) <= (inputs(39)) or (inputs(59));
    layer0_outputs(2291) <= not(inputs(205)) or (inputs(249));
    layer0_outputs(2292) <= not(inputs(186)) or (inputs(99));
    layer0_outputs(2293) <= inputs(101);
    layer0_outputs(2294) <= not(inputs(169));
    layer0_outputs(2295) <= (inputs(45)) and not (inputs(248));
    layer0_outputs(2296) <= (inputs(158)) and (inputs(41));
    layer0_outputs(2297) <= inputs(9);
    layer0_outputs(2298) <= not((inputs(128)) xor (inputs(217)));
    layer0_outputs(2299) <= not(inputs(67)) or (inputs(111));
    layer0_outputs(2300) <= not(inputs(2)) or (inputs(102));
    layer0_outputs(2301) <= not((inputs(93)) xor (inputs(168)));
    layer0_outputs(2302) <= not(inputs(62)) or (inputs(28));
    layer0_outputs(2303) <= not(inputs(96));
    layer0_outputs(2304) <= not(inputs(16));
    layer0_outputs(2305) <= not(inputs(106)) or (inputs(78));
    layer0_outputs(2306) <= (inputs(8)) or (inputs(24));
    layer0_outputs(2307) <= (inputs(206)) or (inputs(20));
    layer0_outputs(2308) <= not(inputs(65));
    layer0_outputs(2309) <= inputs(100);
    layer0_outputs(2310) <= not(inputs(79));
    layer0_outputs(2311) <= (inputs(136)) or (inputs(137));
    layer0_outputs(2312) <= not(inputs(246)) or (inputs(193));
    layer0_outputs(2313) <= '0';
    layer0_outputs(2314) <= not((inputs(7)) or (inputs(194)));
    layer0_outputs(2315) <= (inputs(85)) xor (inputs(51));
    layer0_outputs(2316) <= not(inputs(167)) or (inputs(12));
    layer0_outputs(2317) <= (inputs(198)) or (inputs(97));
    layer0_outputs(2318) <= not(inputs(219));
    layer0_outputs(2319) <= inputs(136);
    layer0_outputs(2320) <= not(inputs(240)) or (inputs(190));
    layer0_outputs(2321) <= not((inputs(135)) xor (inputs(29)));
    layer0_outputs(2322) <= not(inputs(201)) or (inputs(69));
    layer0_outputs(2323) <= (inputs(15)) or (inputs(124));
    layer0_outputs(2324) <= not((inputs(4)) or (inputs(241)));
    layer0_outputs(2325) <= (inputs(224)) and (inputs(220));
    layer0_outputs(2326) <= '1';
    layer0_outputs(2327) <= not(inputs(147));
    layer0_outputs(2328) <= (inputs(159)) xor (inputs(247));
    layer0_outputs(2329) <= (inputs(93)) xor (inputs(82));
    layer0_outputs(2330) <= (inputs(127)) xor (inputs(31));
    layer0_outputs(2331) <= not((inputs(165)) or (inputs(206)));
    layer0_outputs(2332) <= not((inputs(145)) or (inputs(200)));
    layer0_outputs(2333) <= not(inputs(74)) or (inputs(128));
    layer0_outputs(2334) <= not((inputs(250)) and (inputs(5)));
    layer0_outputs(2335) <= (inputs(54)) and not (inputs(228));
    layer0_outputs(2336) <= (inputs(218)) or (inputs(98));
    layer0_outputs(2337) <= (inputs(19)) xor (inputs(17));
    layer0_outputs(2338) <= inputs(151);
    layer0_outputs(2339) <= not(inputs(209)) or (inputs(190));
    layer0_outputs(2340) <= not(inputs(139));
    layer0_outputs(2341) <= (inputs(81)) xor (inputs(185));
    layer0_outputs(2342) <= inputs(228);
    layer0_outputs(2343) <= (inputs(88)) and not (inputs(162));
    layer0_outputs(2344) <= not((inputs(86)) or (inputs(159)));
    layer0_outputs(2345) <= not(inputs(76));
    layer0_outputs(2346) <= (inputs(214)) or (inputs(205));
    layer0_outputs(2347) <= not(inputs(115));
    layer0_outputs(2348) <= not(inputs(53));
    layer0_outputs(2349) <= (inputs(35)) and (inputs(193));
    layer0_outputs(2350) <= not((inputs(188)) or (inputs(190)));
    layer0_outputs(2351) <= not((inputs(35)) or (inputs(221)));
    layer0_outputs(2352) <= inputs(150);
    layer0_outputs(2353) <= not(inputs(239)) or (inputs(96));
    layer0_outputs(2354) <= not(inputs(81)) or (inputs(217));
    layer0_outputs(2355) <= not((inputs(220)) xor (inputs(11)));
    layer0_outputs(2356) <= not(inputs(29)) or (inputs(84));
    layer0_outputs(2357) <= not(inputs(76)) or (inputs(92));
    layer0_outputs(2358) <= not(inputs(207));
    layer0_outputs(2359) <= not(inputs(113));
    layer0_outputs(2360) <= not((inputs(86)) xor (inputs(204)));
    layer0_outputs(2361) <= (inputs(89)) and not (inputs(168));
    layer0_outputs(2362) <= not(inputs(148));
    layer0_outputs(2363) <= not((inputs(185)) or (inputs(14)));
    layer0_outputs(2364) <= not(inputs(52));
    layer0_outputs(2365) <= inputs(23);
    layer0_outputs(2366) <= not(inputs(83)) or (inputs(176));
    layer0_outputs(2367) <= (inputs(120)) and not (inputs(174));
    layer0_outputs(2368) <= not((inputs(118)) and (inputs(136)));
    layer0_outputs(2369) <= (inputs(49)) or (inputs(122));
    layer0_outputs(2370) <= inputs(150);
    layer0_outputs(2371) <= not((inputs(167)) xor (inputs(159)));
    layer0_outputs(2372) <= inputs(51);
    layer0_outputs(2373) <= not((inputs(48)) xor (inputs(69)));
    layer0_outputs(2374) <= not((inputs(80)) or (inputs(200)));
    layer0_outputs(2375) <= not(inputs(102)) or (inputs(188));
    layer0_outputs(2376) <= not((inputs(77)) or (inputs(111)));
    layer0_outputs(2377) <= inputs(180);
    layer0_outputs(2378) <= not((inputs(151)) or (inputs(6)));
    layer0_outputs(2379) <= '1';
    layer0_outputs(2380) <= '1';
    layer0_outputs(2381) <= (inputs(209)) or (inputs(67));
    layer0_outputs(2382) <= (inputs(176)) xor (inputs(173));
    layer0_outputs(2383) <= not(inputs(107));
    layer0_outputs(2384) <= not(inputs(3)) or (inputs(95));
    layer0_outputs(2385) <= not((inputs(47)) and (inputs(15)));
    layer0_outputs(2386) <= not((inputs(247)) or (inputs(105)));
    layer0_outputs(2387) <= inputs(99);
    layer0_outputs(2388) <= not(inputs(44));
    layer0_outputs(2389) <= not(inputs(195));
    layer0_outputs(2390) <= (inputs(239)) or (inputs(81));
    layer0_outputs(2391) <= (inputs(51)) and (inputs(60));
    layer0_outputs(2392) <= (inputs(114)) xor (inputs(231));
    layer0_outputs(2393) <= (inputs(107)) xor (inputs(142));
    layer0_outputs(2394) <= inputs(216);
    layer0_outputs(2395) <= (inputs(59)) and not (inputs(152));
    layer0_outputs(2396) <= not(inputs(40));
    layer0_outputs(2397) <= (inputs(52)) and not (inputs(220));
    layer0_outputs(2398) <= not((inputs(60)) and (inputs(209)));
    layer0_outputs(2399) <= (inputs(134)) or (inputs(15));
    layer0_outputs(2400) <= '1';
    layer0_outputs(2401) <= (inputs(117)) or (inputs(16));
    layer0_outputs(2402) <= (inputs(240)) and (inputs(230));
    layer0_outputs(2403) <= '1';
    layer0_outputs(2404) <= not((inputs(114)) or (inputs(237)));
    layer0_outputs(2405) <= (inputs(130)) or (inputs(240));
    layer0_outputs(2406) <= inputs(247);
    layer0_outputs(2407) <= (inputs(212)) or (inputs(232));
    layer0_outputs(2408) <= (inputs(159)) or (inputs(166));
    layer0_outputs(2409) <= not(inputs(125));
    layer0_outputs(2410) <= (inputs(128)) xor (inputs(182));
    layer0_outputs(2411) <= not(inputs(199));
    layer0_outputs(2412) <= not((inputs(88)) xor (inputs(216)));
    layer0_outputs(2413) <= (inputs(3)) and not (inputs(178));
    layer0_outputs(2414) <= not((inputs(231)) or (inputs(246)));
    layer0_outputs(2415) <= (inputs(162)) and (inputs(129));
    layer0_outputs(2416) <= not(inputs(144));
    layer0_outputs(2417) <= '0';
    layer0_outputs(2418) <= not((inputs(218)) xor (inputs(186)));
    layer0_outputs(2419) <= not((inputs(163)) or (inputs(113)));
    layer0_outputs(2420) <= inputs(3);
    layer0_outputs(2421) <= (inputs(203)) and (inputs(117));
    layer0_outputs(2422) <= not((inputs(134)) or (inputs(112)));
    layer0_outputs(2423) <= (inputs(129)) or (inputs(49));
    layer0_outputs(2424) <= '0';
    layer0_outputs(2425) <= not((inputs(121)) or (inputs(108)));
    layer0_outputs(2426) <= (inputs(226)) xor (inputs(243));
    layer0_outputs(2427) <= (inputs(57)) and not (inputs(170));
    layer0_outputs(2428) <= (inputs(192)) xor (inputs(106));
    layer0_outputs(2429) <= (inputs(7)) xor (inputs(63));
    layer0_outputs(2430) <= not(inputs(183)) or (inputs(78));
    layer0_outputs(2431) <= not(inputs(58));
    layer0_outputs(2432) <= (inputs(79)) and (inputs(211));
    layer0_outputs(2433) <= (inputs(20)) or (inputs(234));
    layer0_outputs(2434) <= '0';
    layer0_outputs(2435) <= (inputs(47)) and not (inputs(252));
    layer0_outputs(2436) <= not((inputs(82)) or (inputs(254)));
    layer0_outputs(2437) <= (inputs(34)) and not (inputs(102));
    layer0_outputs(2438) <= (inputs(2)) or (inputs(37));
    layer0_outputs(2439) <= not((inputs(238)) and (inputs(114)));
    layer0_outputs(2440) <= not((inputs(8)) and (inputs(183)));
    layer0_outputs(2441) <= not(inputs(71)) or (inputs(25));
    layer0_outputs(2442) <= not(inputs(102));
    layer0_outputs(2443) <= '0';
    layer0_outputs(2444) <= inputs(230);
    layer0_outputs(2445) <= (inputs(138)) or (inputs(226));
    layer0_outputs(2446) <= inputs(85);
    layer0_outputs(2447) <= not(inputs(78));
    layer0_outputs(2448) <= (inputs(4)) and not (inputs(197));
    layer0_outputs(2449) <= (inputs(30)) and not (inputs(126));
    layer0_outputs(2450) <= not(inputs(200));
    layer0_outputs(2451) <= (inputs(180)) or (inputs(186));
    layer0_outputs(2452) <= inputs(215);
    layer0_outputs(2453) <= (inputs(95)) and not (inputs(36));
    layer0_outputs(2454) <= not(inputs(65));
    layer0_outputs(2455) <= (inputs(149)) xor (inputs(172));
    layer0_outputs(2456) <= (inputs(180)) and not (inputs(28));
    layer0_outputs(2457) <= not(inputs(60));
    layer0_outputs(2458) <= not(inputs(76));
    layer0_outputs(2459) <= inputs(196);
    layer0_outputs(2460) <= not(inputs(94));
    layer0_outputs(2461) <= inputs(168);
    layer0_outputs(2462) <= (inputs(147)) or (inputs(65));
    layer0_outputs(2463) <= not((inputs(189)) or (inputs(255)));
    layer0_outputs(2464) <= (inputs(206)) or (inputs(180));
    layer0_outputs(2465) <= (inputs(235)) and (inputs(225));
    layer0_outputs(2466) <= (inputs(48)) and not (inputs(26));
    layer0_outputs(2467) <= not((inputs(73)) or (inputs(23)));
    layer0_outputs(2468) <= not((inputs(111)) and (inputs(246)));
    layer0_outputs(2469) <= '1';
    layer0_outputs(2470) <= '1';
    layer0_outputs(2471) <= not(inputs(90));
    layer0_outputs(2472) <= (inputs(245)) xor (inputs(85));
    layer0_outputs(2473) <= not((inputs(91)) xor (inputs(159)));
    layer0_outputs(2474) <= inputs(157);
    layer0_outputs(2475) <= not(inputs(234)) or (inputs(27));
    layer0_outputs(2476) <= not(inputs(165)) or (inputs(230));
    layer0_outputs(2477) <= '0';
    layer0_outputs(2478) <= not(inputs(93)) or (inputs(109));
    layer0_outputs(2479) <= inputs(166);
    layer0_outputs(2480) <= '0';
    layer0_outputs(2481) <= not(inputs(237));
    layer0_outputs(2482) <= (inputs(236)) and (inputs(4));
    layer0_outputs(2483) <= '1';
    layer0_outputs(2484) <= '1';
    layer0_outputs(2485) <= not(inputs(239)) or (inputs(3));
    layer0_outputs(2486) <= (inputs(56)) xor (inputs(244));
    layer0_outputs(2487) <= not((inputs(20)) xor (inputs(158)));
    layer0_outputs(2488) <= not((inputs(10)) or (inputs(52)));
    layer0_outputs(2489) <= (inputs(62)) or (inputs(93));
    layer0_outputs(2490) <= inputs(42);
    layer0_outputs(2491) <= '0';
    layer0_outputs(2492) <= not(inputs(151)) or (inputs(252));
    layer0_outputs(2493) <= (inputs(192)) or (inputs(86));
    layer0_outputs(2494) <= inputs(248);
    layer0_outputs(2495) <= not(inputs(107)) or (inputs(45));
    layer0_outputs(2496) <= inputs(163);
    layer0_outputs(2497) <= not(inputs(136));
    layer0_outputs(2498) <= not((inputs(10)) and (inputs(244)));
    layer0_outputs(2499) <= not(inputs(241));
    layer0_outputs(2500) <= (inputs(144)) or (inputs(102));
    layer0_outputs(2501) <= (inputs(178)) and not (inputs(245));
    layer0_outputs(2502) <= not((inputs(151)) xor (inputs(237)));
    layer0_outputs(2503) <= not(inputs(207)) or (inputs(1));
    layer0_outputs(2504) <= not((inputs(171)) or (inputs(207)));
    layer0_outputs(2505) <= (inputs(242)) and not (inputs(225));
    layer0_outputs(2506) <= '0';
    layer0_outputs(2507) <= not(inputs(117));
    layer0_outputs(2508) <= (inputs(162)) or (inputs(89));
    layer0_outputs(2509) <= (inputs(130)) and (inputs(194));
    layer0_outputs(2510) <= inputs(239);
    layer0_outputs(2511) <= (inputs(253)) and (inputs(209));
    layer0_outputs(2512) <= (inputs(135)) or (inputs(152));
    layer0_outputs(2513) <= not((inputs(133)) or (inputs(4)));
    layer0_outputs(2514) <= (inputs(102)) and not (inputs(226));
    layer0_outputs(2515) <= '0';
    layer0_outputs(2516) <= not(inputs(103)) or (inputs(177));
    layer0_outputs(2517) <= '1';
    layer0_outputs(2518) <= inputs(179);
    layer0_outputs(2519) <= not((inputs(126)) or (inputs(124)));
    layer0_outputs(2520) <= (inputs(110)) and not (inputs(53));
    layer0_outputs(2521) <= (inputs(252)) xor (inputs(229));
    layer0_outputs(2522) <= (inputs(235)) and not (inputs(61));
    layer0_outputs(2523) <= not(inputs(103));
    layer0_outputs(2524) <= (inputs(209)) or (inputs(71));
    layer0_outputs(2525) <= not(inputs(108));
    layer0_outputs(2526) <= '0';
    layer0_outputs(2527) <= '1';
    layer0_outputs(2528) <= (inputs(40)) or (inputs(52));
    layer0_outputs(2529) <= not(inputs(216)) or (inputs(146));
    layer0_outputs(2530) <= inputs(206);
    layer0_outputs(2531) <= (inputs(242)) and (inputs(69));
    layer0_outputs(2532) <= not(inputs(184));
    layer0_outputs(2533) <= not((inputs(142)) xor (inputs(98)));
    layer0_outputs(2534) <= '1';
    layer0_outputs(2535) <= (inputs(27)) xor (inputs(70));
    layer0_outputs(2536) <= (inputs(176)) and (inputs(88));
    layer0_outputs(2537) <= not(inputs(135)) or (inputs(248));
    layer0_outputs(2538) <= not(inputs(152)) or (inputs(161));
    layer0_outputs(2539) <= not(inputs(182));
    layer0_outputs(2540) <= not((inputs(180)) xor (inputs(131)));
    layer0_outputs(2541) <= not(inputs(153));
    layer0_outputs(2542) <= not(inputs(168)) or (inputs(1));
    layer0_outputs(2543) <= (inputs(10)) and not (inputs(231));
    layer0_outputs(2544) <= (inputs(112)) and (inputs(51));
    layer0_outputs(2545) <= not(inputs(27));
    layer0_outputs(2546) <= (inputs(47)) and (inputs(28));
    layer0_outputs(2547) <= not(inputs(252)) or (inputs(242));
    layer0_outputs(2548) <= not(inputs(175)) or (inputs(130));
    layer0_outputs(2549) <= not((inputs(253)) xor (inputs(157)));
    layer0_outputs(2550) <= not((inputs(228)) and (inputs(211)));
    layer0_outputs(2551) <= not(inputs(94));
    layer0_outputs(2552) <= inputs(216);
    layer0_outputs(2553) <= (inputs(3)) and not (inputs(133));
    layer0_outputs(2554) <= (inputs(168)) and not (inputs(193));
    layer0_outputs(2555) <= not(inputs(124)) or (inputs(130));
    layer0_outputs(2556) <= '0';
    layer0_outputs(2557) <= inputs(90);
    layer0_outputs(2558) <= not(inputs(60));
    layer0_outputs(2559) <= not(inputs(200));
    layer0_outputs(2560) <= '1';
    layer0_outputs(2561) <= (inputs(235)) and not (inputs(194));
    layer0_outputs(2562) <= not((inputs(216)) xor (inputs(161)));
    layer0_outputs(2563) <= not((inputs(53)) xor (inputs(249)));
    layer0_outputs(2564) <= '0';
    layer0_outputs(2565) <= not((inputs(44)) and (inputs(190)));
    layer0_outputs(2566) <= '1';
    layer0_outputs(2567) <= not(inputs(120));
    layer0_outputs(2568) <= inputs(252);
    layer0_outputs(2569) <= '0';
    layer0_outputs(2570) <= not(inputs(210)) or (inputs(140));
    layer0_outputs(2571) <= '0';
    layer0_outputs(2572) <= not(inputs(83));
    layer0_outputs(2573) <= not(inputs(206));
    layer0_outputs(2574) <= inputs(91);
    layer0_outputs(2575) <= (inputs(255)) xor (inputs(155));
    layer0_outputs(2576) <= (inputs(175)) xor (inputs(91));
    layer0_outputs(2577) <= not(inputs(121));
    layer0_outputs(2578) <= not(inputs(149));
    layer0_outputs(2579) <= (inputs(0)) and not (inputs(113));
    layer0_outputs(2580) <= not((inputs(253)) or (inputs(39)));
    layer0_outputs(2581) <= (inputs(213)) or (inputs(96));
    layer0_outputs(2582) <= not(inputs(168));
    layer0_outputs(2583) <= (inputs(149)) and not (inputs(163));
    layer0_outputs(2584) <= inputs(200);
    layer0_outputs(2585) <= (inputs(218)) xor (inputs(248));
    layer0_outputs(2586) <= not(inputs(107));
    layer0_outputs(2587) <= not(inputs(125)) or (inputs(2));
    layer0_outputs(2588) <= inputs(123);
    layer0_outputs(2589) <= not((inputs(107)) and (inputs(96)));
    layer0_outputs(2590) <= not((inputs(41)) and (inputs(174)));
    layer0_outputs(2591) <= not(inputs(7));
    layer0_outputs(2592) <= inputs(3);
    layer0_outputs(2593) <= not((inputs(227)) and (inputs(63)));
    layer0_outputs(2594) <= not((inputs(108)) or (inputs(27)));
    layer0_outputs(2595) <= not(inputs(110));
    layer0_outputs(2596) <= (inputs(80)) and not (inputs(93));
    layer0_outputs(2597) <= not((inputs(146)) or (inputs(186)));
    layer0_outputs(2598) <= (inputs(182)) or (inputs(81));
    layer0_outputs(2599) <= (inputs(87)) and not (inputs(105));
    layer0_outputs(2600) <= not(inputs(126)) or (inputs(64));
    layer0_outputs(2601) <= not((inputs(62)) or (inputs(180)));
    layer0_outputs(2602) <= '0';
    layer0_outputs(2603) <= '1';
    layer0_outputs(2604) <= not((inputs(57)) xor (inputs(82)));
    layer0_outputs(2605) <= (inputs(241)) xor (inputs(9));
    layer0_outputs(2606) <= not(inputs(133));
    layer0_outputs(2607) <= not((inputs(130)) or (inputs(235)));
    layer0_outputs(2608) <= not(inputs(156)) or (inputs(79));
    layer0_outputs(2609) <= (inputs(191)) xor (inputs(80));
    layer0_outputs(2610) <= not((inputs(100)) or (inputs(61)));
    layer0_outputs(2611) <= inputs(217);
    layer0_outputs(2612) <= not(inputs(135));
    layer0_outputs(2613) <= not((inputs(109)) xor (inputs(10)));
    layer0_outputs(2614) <= not(inputs(149));
    layer0_outputs(2615) <= not((inputs(43)) or (inputs(220)));
    layer0_outputs(2616) <= (inputs(163)) and not (inputs(111));
    layer0_outputs(2617) <= not(inputs(15));
    layer0_outputs(2618) <= (inputs(195)) xor (inputs(8));
    layer0_outputs(2619) <= not((inputs(80)) or (inputs(112)));
    layer0_outputs(2620) <= (inputs(17)) and not (inputs(48));
    layer0_outputs(2621) <= not(inputs(188));
    layer0_outputs(2622) <= not(inputs(210));
    layer0_outputs(2623) <= inputs(246);
    layer0_outputs(2624) <= (inputs(98)) xor (inputs(9));
    layer0_outputs(2625) <= not((inputs(30)) or (inputs(202)));
    layer0_outputs(2626) <= (inputs(131)) and not (inputs(62));
    layer0_outputs(2627) <= (inputs(16)) or (inputs(125));
    layer0_outputs(2628) <= not(inputs(25));
    layer0_outputs(2629) <= not((inputs(200)) or (inputs(96)));
    layer0_outputs(2630) <= inputs(106);
    layer0_outputs(2631) <= not((inputs(144)) and (inputs(251)));
    layer0_outputs(2632) <= not((inputs(118)) or (inputs(230)));
    layer0_outputs(2633) <= not(inputs(139));
    layer0_outputs(2634) <= (inputs(226)) and not (inputs(10));
    layer0_outputs(2635) <= (inputs(113)) xor (inputs(1));
    layer0_outputs(2636) <= (inputs(242)) or (inputs(250));
    layer0_outputs(2637) <= not(inputs(133));
    layer0_outputs(2638) <= (inputs(115)) and not (inputs(62));
    layer0_outputs(2639) <= not(inputs(182));
    layer0_outputs(2640) <= (inputs(170)) or (inputs(141));
    layer0_outputs(2641) <= not(inputs(105)) or (inputs(191));
    layer0_outputs(2642) <= (inputs(173)) or (inputs(38));
    layer0_outputs(2643) <= not((inputs(253)) or (inputs(16)));
    layer0_outputs(2644) <= not(inputs(45)) or (inputs(207));
    layer0_outputs(2645) <= not((inputs(26)) xor (inputs(182)));
    layer0_outputs(2646) <= (inputs(193)) xor (inputs(230));
    layer0_outputs(2647) <= (inputs(162)) or (inputs(66));
    layer0_outputs(2648) <= not(inputs(106)) or (inputs(129));
    layer0_outputs(2649) <= not(inputs(182));
    layer0_outputs(2650) <= not(inputs(110)) or (inputs(192));
    layer0_outputs(2651) <= '1';
    layer0_outputs(2652) <= (inputs(23)) and (inputs(28));
    layer0_outputs(2653) <= (inputs(12)) or (inputs(116));
    layer0_outputs(2654) <= inputs(52);
    layer0_outputs(2655) <= (inputs(6)) xor (inputs(155));
    layer0_outputs(2656) <= '1';
    layer0_outputs(2657) <= (inputs(217)) xor (inputs(110));
    layer0_outputs(2658) <= inputs(181);
    layer0_outputs(2659) <= (inputs(118)) or (inputs(209));
    layer0_outputs(2660) <= inputs(34);
    layer0_outputs(2661) <= (inputs(164)) and not (inputs(131));
    layer0_outputs(2662) <= not((inputs(227)) and (inputs(115)));
    layer0_outputs(2663) <= not((inputs(235)) and (inputs(25)));
    layer0_outputs(2664) <= inputs(241);
    layer0_outputs(2665) <= not(inputs(172));
    layer0_outputs(2666) <= inputs(216);
    layer0_outputs(2667) <= not(inputs(85)) or (inputs(209));
    layer0_outputs(2668) <= inputs(167);
    layer0_outputs(2669) <= (inputs(186)) or (inputs(225));
    layer0_outputs(2670) <= not(inputs(105)) or (inputs(244));
    layer0_outputs(2671) <= not(inputs(7)) or (inputs(21));
    layer0_outputs(2672) <= inputs(65);
    layer0_outputs(2673) <= not(inputs(210)) or (inputs(130));
    layer0_outputs(2674) <= (inputs(183)) or (inputs(178));
    layer0_outputs(2675) <= not(inputs(150));
    layer0_outputs(2676) <= not(inputs(209));
    layer0_outputs(2677) <= (inputs(199)) and not (inputs(160));
    layer0_outputs(2678) <= not(inputs(36)) or (inputs(84));
    layer0_outputs(2679) <= not(inputs(183)) or (inputs(253));
    layer0_outputs(2680) <= (inputs(90)) and not (inputs(133));
    layer0_outputs(2681) <= not(inputs(89)) or (inputs(22));
    layer0_outputs(2682) <= not(inputs(70));
    layer0_outputs(2683) <= inputs(197);
    layer0_outputs(2684) <= not((inputs(84)) or (inputs(197)));
    layer0_outputs(2685) <= inputs(185);
    layer0_outputs(2686) <= not(inputs(59)) or (inputs(191));
    layer0_outputs(2687) <= not((inputs(67)) or (inputs(105)));
    layer0_outputs(2688) <= (inputs(214)) or (inputs(130));
    layer0_outputs(2689) <= inputs(119);
    layer0_outputs(2690) <= not((inputs(70)) and (inputs(127)));
    layer0_outputs(2691) <= not(inputs(177));
    layer0_outputs(2692) <= not(inputs(106));
    layer0_outputs(2693) <= (inputs(244)) and not (inputs(173));
    layer0_outputs(2694) <= (inputs(127)) or (inputs(115));
    layer0_outputs(2695) <= not((inputs(195)) or (inputs(178)));
    layer0_outputs(2696) <= not(inputs(187)) or (inputs(84));
    layer0_outputs(2697) <= not(inputs(144));
    layer0_outputs(2698) <= not((inputs(200)) or (inputs(144)));
    layer0_outputs(2699) <= not(inputs(142));
    layer0_outputs(2700) <= inputs(238);
    layer0_outputs(2701) <= not(inputs(122));
    layer0_outputs(2702) <= inputs(152);
    layer0_outputs(2703) <= not(inputs(69));
    layer0_outputs(2704) <= (inputs(18)) and not (inputs(161));
    layer0_outputs(2705) <= (inputs(218)) xor (inputs(146));
    layer0_outputs(2706) <= not(inputs(151));
    layer0_outputs(2707) <= (inputs(156)) and not (inputs(160));
    layer0_outputs(2708) <= (inputs(167)) or (inputs(224));
    layer0_outputs(2709) <= (inputs(217)) and not (inputs(44));
    layer0_outputs(2710) <= not((inputs(35)) or (inputs(57)));
    layer0_outputs(2711) <= not((inputs(116)) or (inputs(25)));
    layer0_outputs(2712) <= (inputs(177)) and not (inputs(221));
    layer0_outputs(2713) <= (inputs(254)) or (inputs(103));
    layer0_outputs(2714) <= (inputs(94)) and not (inputs(16));
    layer0_outputs(2715) <= not(inputs(101));
    layer0_outputs(2716) <= (inputs(249)) and (inputs(109));
    layer0_outputs(2717) <= not(inputs(223));
    layer0_outputs(2718) <= (inputs(232)) and not (inputs(160));
    layer0_outputs(2719) <= (inputs(243)) xor (inputs(149));
    layer0_outputs(2720) <= not(inputs(134));
    layer0_outputs(2721) <= not((inputs(210)) and (inputs(11)));
    layer0_outputs(2722) <= not((inputs(130)) xor (inputs(46)));
    layer0_outputs(2723) <= not(inputs(174)) or (inputs(79));
    layer0_outputs(2724) <= not(inputs(110)) or (inputs(239));
    layer0_outputs(2725) <= inputs(238);
    layer0_outputs(2726) <= (inputs(132)) or (inputs(162));
    layer0_outputs(2727) <= '0';
    layer0_outputs(2728) <= not((inputs(221)) or (inputs(238)));
    layer0_outputs(2729) <= not((inputs(37)) or (inputs(151)));
    layer0_outputs(2730) <= not((inputs(173)) or (inputs(6)));
    layer0_outputs(2731) <= '0';
    layer0_outputs(2732) <= not((inputs(222)) xor (inputs(134)));
    layer0_outputs(2733) <= '0';
    layer0_outputs(2734) <= not((inputs(192)) or (inputs(238)));
    layer0_outputs(2735) <= not((inputs(176)) xor (inputs(36)));
    layer0_outputs(2736) <= not(inputs(133)) or (inputs(81));
    layer0_outputs(2737) <= '0';
    layer0_outputs(2738) <= '1';
    layer0_outputs(2739) <= (inputs(79)) xor (inputs(12));
    layer0_outputs(2740) <= not(inputs(117));
    layer0_outputs(2741) <= '1';
    layer0_outputs(2742) <= not(inputs(239)) or (inputs(77));
    layer0_outputs(2743) <= (inputs(190)) or (inputs(153));
    layer0_outputs(2744) <= not(inputs(126));
    layer0_outputs(2745) <= not(inputs(231));
    layer0_outputs(2746) <= not(inputs(184));
    layer0_outputs(2747) <= inputs(179);
    layer0_outputs(2748) <= not(inputs(19));
    layer0_outputs(2749) <= not(inputs(191)) or (inputs(136));
    layer0_outputs(2750) <= not(inputs(0));
    layer0_outputs(2751) <= inputs(168);
    layer0_outputs(2752) <= not(inputs(101));
    layer0_outputs(2753) <= (inputs(97)) and (inputs(33));
    layer0_outputs(2754) <= '0';
    layer0_outputs(2755) <= (inputs(241)) or (inputs(50));
    layer0_outputs(2756) <= not((inputs(107)) and (inputs(77)));
    layer0_outputs(2757) <= inputs(88);
    layer0_outputs(2758) <= inputs(177);
    layer0_outputs(2759) <= (inputs(209)) and not (inputs(117));
    layer0_outputs(2760) <= (inputs(107)) or (inputs(163));
    layer0_outputs(2761) <= (inputs(23)) or (inputs(140));
    layer0_outputs(2762) <= (inputs(108)) and not (inputs(204));
    layer0_outputs(2763) <= not(inputs(223));
    layer0_outputs(2764) <= (inputs(91)) or (inputs(67));
    layer0_outputs(2765) <= '0';
    layer0_outputs(2766) <= not(inputs(196));
    layer0_outputs(2767) <= not(inputs(188));
    layer0_outputs(2768) <= (inputs(221)) and not (inputs(119));
    layer0_outputs(2769) <= not(inputs(72)) or (inputs(191));
    layer0_outputs(2770) <= (inputs(185)) or (inputs(22));
    layer0_outputs(2771) <= (inputs(154)) and not (inputs(41));
    layer0_outputs(2772) <= inputs(66);
    layer0_outputs(2773) <= (inputs(73)) or (inputs(99));
    layer0_outputs(2774) <= not((inputs(92)) xor (inputs(110)));
    layer0_outputs(2775) <= (inputs(164)) and not (inputs(136));
    layer0_outputs(2776) <= not(inputs(23));
    layer0_outputs(2777) <= (inputs(117)) and not (inputs(206));
    layer0_outputs(2778) <= '1';
    layer0_outputs(2779) <= (inputs(200)) and not (inputs(210));
    layer0_outputs(2780) <= inputs(132);
    layer0_outputs(2781) <= inputs(22);
    layer0_outputs(2782) <= (inputs(248)) or (inputs(172));
    layer0_outputs(2783) <= not((inputs(101)) xor (inputs(80)));
    layer0_outputs(2784) <= '0';
    layer0_outputs(2785) <= inputs(164);
    layer0_outputs(2786) <= (inputs(224)) and (inputs(179));
    layer0_outputs(2787) <= not((inputs(120)) or (inputs(161)));
    layer0_outputs(2788) <= (inputs(47)) and not (inputs(83));
    layer0_outputs(2789) <= '1';
    layer0_outputs(2790) <= (inputs(78)) and (inputs(246));
    layer0_outputs(2791) <= not(inputs(132)) or (inputs(229));
    layer0_outputs(2792) <= not(inputs(133)) or (inputs(62));
    layer0_outputs(2793) <= not((inputs(211)) or (inputs(77)));
    layer0_outputs(2794) <= inputs(106);
    layer0_outputs(2795) <= not((inputs(95)) or (inputs(255)));
    layer0_outputs(2796) <= (inputs(172)) and not (inputs(15));
    layer0_outputs(2797) <= (inputs(80)) or (inputs(252));
    layer0_outputs(2798) <= (inputs(96)) xor (inputs(58));
    layer0_outputs(2799) <= (inputs(152)) and not (inputs(171));
    layer0_outputs(2800) <= not(inputs(101));
    layer0_outputs(2801) <= not((inputs(200)) or (inputs(194)));
    layer0_outputs(2802) <= not(inputs(189));
    layer0_outputs(2803) <= '1';
    layer0_outputs(2804) <= not(inputs(216)) or (inputs(194));
    layer0_outputs(2805) <= (inputs(210)) and not (inputs(38));
    layer0_outputs(2806) <= '0';
    layer0_outputs(2807) <= not(inputs(125));
    layer0_outputs(2808) <= not((inputs(227)) or (inputs(50)));
    layer0_outputs(2809) <= not(inputs(235)) or (inputs(238));
    layer0_outputs(2810) <= not(inputs(62));
    layer0_outputs(2811) <= not((inputs(214)) or (inputs(180)));
    layer0_outputs(2812) <= inputs(195);
    layer0_outputs(2813) <= not(inputs(186)) or (inputs(124));
    layer0_outputs(2814) <= (inputs(229)) or (inputs(89));
    layer0_outputs(2815) <= not((inputs(0)) or (inputs(205)));
    layer0_outputs(2816) <= not((inputs(229)) or (inputs(101)));
    layer0_outputs(2817) <= (inputs(160)) and not (inputs(65));
    layer0_outputs(2818) <= (inputs(233)) or (inputs(162));
    layer0_outputs(2819) <= (inputs(193)) xor (inputs(72));
    layer0_outputs(2820) <= not(inputs(172)) or (inputs(6));
    layer0_outputs(2821) <= (inputs(35)) or (inputs(81));
    layer0_outputs(2822) <= (inputs(188)) or (inputs(75));
    layer0_outputs(2823) <= not((inputs(95)) and (inputs(5)));
    layer0_outputs(2824) <= not(inputs(120));
    layer0_outputs(2825) <= not(inputs(245)) or (inputs(63));
    layer0_outputs(2826) <= not((inputs(97)) and (inputs(226)));
    layer0_outputs(2827) <= not(inputs(204));
    layer0_outputs(2828) <= (inputs(18)) and not (inputs(223));
    layer0_outputs(2829) <= not(inputs(250)) or (inputs(250));
    layer0_outputs(2830) <= not(inputs(40));
    layer0_outputs(2831) <= not((inputs(235)) or (inputs(205)));
    layer0_outputs(2832) <= not(inputs(91)) or (inputs(140));
    layer0_outputs(2833) <= (inputs(123)) and not (inputs(0));
    layer0_outputs(2834) <= not(inputs(21));
    layer0_outputs(2835) <= '0';
    layer0_outputs(2836) <= (inputs(14)) and not (inputs(162));
    layer0_outputs(2837) <= (inputs(96)) and not (inputs(173));
    layer0_outputs(2838) <= not(inputs(168));
    layer0_outputs(2839) <= not((inputs(81)) or (inputs(126)));
    layer0_outputs(2840) <= (inputs(199)) and not (inputs(53));
    layer0_outputs(2841) <= inputs(55);
    layer0_outputs(2842) <= inputs(140);
    layer0_outputs(2843) <= not(inputs(147));
    layer0_outputs(2844) <= not(inputs(55));
    layer0_outputs(2845) <= not(inputs(8)) or (inputs(37));
    layer0_outputs(2846) <= not((inputs(255)) or (inputs(1)));
    layer0_outputs(2847) <= (inputs(12)) and not (inputs(106));
    layer0_outputs(2848) <= '0';
    layer0_outputs(2849) <= not((inputs(35)) and (inputs(253)));
    layer0_outputs(2850) <= (inputs(205)) or (inputs(211));
    layer0_outputs(2851) <= (inputs(99)) xor (inputs(210));
    layer0_outputs(2852) <= not(inputs(100)) or (inputs(156));
    layer0_outputs(2853) <= '0';
    layer0_outputs(2854) <= (inputs(10)) xor (inputs(118));
    layer0_outputs(2855) <= not((inputs(224)) or (inputs(163)));
    layer0_outputs(2856) <= not(inputs(166)) or (inputs(163));
    layer0_outputs(2857) <= inputs(94);
    layer0_outputs(2858) <= not((inputs(237)) or (inputs(122)));
    layer0_outputs(2859) <= not(inputs(150)) or (inputs(8));
    layer0_outputs(2860) <= not((inputs(149)) and (inputs(239)));
    layer0_outputs(2861) <= not((inputs(105)) and (inputs(44)));
    layer0_outputs(2862) <= (inputs(51)) and not (inputs(175));
    layer0_outputs(2863) <= not(inputs(114));
    layer0_outputs(2864) <= (inputs(72)) or (inputs(73));
    layer0_outputs(2865) <= not(inputs(153));
    layer0_outputs(2866) <= not(inputs(218));
    layer0_outputs(2867) <= '0';
    layer0_outputs(2868) <= not(inputs(99));
    layer0_outputs(2869) <= not(inputs(21)) or (inputs(80));
    layer0_outputs(2870) <= (inputs(90)) xor (inputs(33));
    layer0_outputs(2871) <= not(inputs(206)) or (inputs(4));
    layer0_outputs(2872) <= not(inputs(112));
    layer0_outputs(2873) <= not((inputs(4)) or (inputs(162)));
    layer0_outputs(2874) <= (inputs(68)) and not (inputs(131));
    layer0_outputs(2875) <= not(inputs(17));
    layer0_outputs(2876) <= not((inputs(226)) xor (inputs(132)));
    layer0_outputs(2877) <= '1';
    layer0_outputs(2878) <= not(inputs(92));
    layer0_outputs(2879) <= '0';
    layer0_outputs(2880) <= inputs(162);
    layer0_outputs(2881) <= (inputs(229)) or (inputs(251));
    layer0_outputs(2882) <= not((inputs(252)) or (inputs(203)));
    layer0_outputs(2883) <= not(inputs(58)) or (inputs(134));
    layer0_outputs(2884) <= not(inputs(89));
    layer0_outputs(2885) <= not((inputs(175)) or (inputs(77)));
    layer0_outputs(2886) <= not((inputs(112)) and (inputs(142)));
    layer0_outputs(2887) <= not(inputs(100)) or (inputs(144));
    layer0_outputs(2888) <= not((inputs(53)) or (inputs(204)));
    layer0_outputs(2889) <= not(inputs(43)) or (inputs(255));
    layer0_outputs(2890) <= not(inputs(78));
    layer0_outputs(2891) <= not(inputs(160)) or (inputs(207));
    layer0_outputs(2892) <= not(inputs(57)) or (inputs(238));
    layer0_outputs(2893) <= (inputs(153)) and not (inputs(66));
    layer0_outputs(2894) <= (inputs(94)) and not (inputs(27));
    layer0_outputs(2895) <= inputs(134);
    layer0_outputs(2896) <= not(inputs(131));
    layer0_outputs(2897) <= inputs(88);
    layer0_outputs(2898) <= (inputs(0)) and not (inputs(126));
    layer0_outputs(2899) <= not((inputs(143)) or (inputs(90)));
    layer0_outputs(2900) <= not((inputs(128)) or (inputs(202)));
    layer0_outputs(2901) <= not(inputs(99)) or (inputs(214));
    layer0_outputs(2902) <= '0';
    layer0_outputs(2903) <= not((inputs(162)) or (inputs(187)));
    layer0_outputs(2904) <= not(inputs(141));
    layer0_outputs(2905) <= (inputs(228)) xor (inputs(200));
    layer0_outputs(2906) <= (inputs(120)) and not (inputs(70));
    layer0_outputs(2907) <= not(inputs(132)) or (inputs(245));
    layer0_outputs(2908) <= not(inputs(87));
    layer0_outputs(2909) <= inputs(148);
    layer0_outputs(2910) <= (inputs(125)) or (inputs(184));
    layer0_outputs(2911) <= (inputs(128)) and not (inputs(159));
    layer0_outputs(2912) <= (inputs(231)) and not (inputs(217));
    layer0_outputs(2913) <= inputs(11);
    layer0_outputs(2914) <= not(inputs(180)) or (inputs(221));
    layer0_outputs(2915) <= (inputs(164)) xor (inputs(144));
    layer0_outputs(2916) <= not(inputs(136)) or (inputs(57));
    layer0_outputs(2917) <= not((inputs(241)) or (inputs(154)));
    layer0_outputs(2918) <= inputs(54);
    layer0_outputs(2919) <= (inputs(137)) or (inputs(138));
    layer0_outputs(2920) <= inputs(107);
    layer0_outputs(2921) <= (inputs(238)) or (inputs(143));
    layer0_outputs(2922) <= not(inputs(151)) or (inputs(94));
    layer0_outputs(2923) <= (inputs(7)) or (inputs(53));
    layer0_outputs(2924) <= not(inputs(119));
    layer0_outputs(2925) <= not((inputs(243)) and (inputs(225)));
    layer0_outputs(2926) <= not(inputs(249));
    layer0_outputs(2927) <= (inputs(171)) or (inputs(155));
    layer0_outputs(2928) <= (inputs(241)) and not (inputs(28));
    layer0_outputs(2929) <= not(inputs(136)) or (inputs(228));
    layer0_outputs(2930) <= (inputs(222)) xor (inputs(25));
    layer0_outputs(2931) <= '0';
    layer0_outputs(2932) <= inputs(78);
    layer0_outputs(2933) <= inputs(207);
    layer0_outputs(2934) <= inputs(61);
    layer0_outputs(2935) <= not(inputs(38));
    layer0_outputs(2936) <= not((inputs(82)) or (inputs(195)));
    layer0_outputs(2937) <= (inputs(56)) and not (inputs(219));
    layer0_outputs(2938) <= (inputs(195)) or (inputs(145));
    layer0_outputs(2939) <= not((inputs(75)) or (inputs(111)));
    layer0_outputs(2940) <= inputs(232);
    layer0_outputs(2941) <= inputs(67);
    layer0_outputs(2942) <= '1';
    layer0_outputs(2943) <= (inputs(251)) or (inputs(89));
    layer0_outputs(2944) <= not(inputs(54)) or (inputs(60));
    layer0_outputs(2945) <= inputs(26);
    layer0_outputs(2946) <= inputs(80);
    layer0_outputs(2947) <= (inputs(66)) and not (inputs(238));
    layer0_outputs(2948) <= not((inputs(188)) or (inputs(173)));
    layer0_outputs(2949) <= not((inputs(16)) or (inputs(153)));
    layer0_outputs(2950) <= inputs(214);
    layer0_outputs(2951) <= (inputs(250)) and not (inputs(74));
    layer0_outputs(2952) <= not((inputs(123)) and (inputs(37)));
    layer0_outputs(2953) <= not((inputs(242)) xor (inputs(127)));
    layer0_outputs(2954) <= not(inputs(83));
    layer0_outputs(2955) <= not(inputs(16));
    layer0_outputs(2956) <= not(inputs(177));
    layer0_outputs(2957) <= inputs(35);
    layer0_outputs(2958) <= (inputs(13)) and not (inputs(80));
    layer0_outputs(2959) <= not(inputs(102));
    layer0_outputs(2960) <= inputs(231);
    layer0_outputs(2961) <= not((inputs(132)) xor (inputs(251)));
    layer0_outputs(2962) <= (inputs(29)) xor (inputs(201));
    layer0_outputs(2963) <= (inputs(178)) and (inputs(53));
    layer0_outputs(2964) <= (inputs(2)) xor (inputs(34));
    layer0_outputs(2965) <= not(inputs(219));
    layer0_outputs(2966) <= not((inputs(232)) or (inputs(223)));
    layer0_outputs(2967) <= (inputs(0)) and (inputs(163));
    layer0_outputs(2968) <= not((inputs(56)) or (inputs(112)));
    layer0_outputs(2969) <= (inputs(73)) and not (inputs(14));
    layer0_outputs(2970) <= inputs(60);
    layer0_outputs(2971) <= (inputs(64)) and not (inputs(229));
    layer0_outputs(2972) <= (inputs(106)) or (inputs(158));
    layer0_outputs(2973) <= not(inputs(128)) or (inputs(157));
    layer0_outputs(2974) <= (inputs(211)) or (inputs(78));
    layer0_outputs(2975) <= not((inputs(246)) or (inputs(90)));
    layer0_outputs(2976) <= not(inputs(71));
    layer0_outputs(2977) <= inputs(85);
    layer0_outputs(2978) <= not(inputs(116));
    layer0_outputs(2979) <= not((inputs(141)) or (inputs(64)));
    layer0_outputs(2980) <= not(inputs(164)) or (inputs(250));
    layer0_outputs(2981) <= not(inputs(125)) or (inputs(206));
    layer0_outputs(2982) <= (inputs(186)) and not (inputs(42));
    layer0_outputs(2983) <= inputs(56);
    layer0_outputs(2984) <= (inputs(50)) or (inputs(120));
    layer0_outputs(2985) <= not((inputs(127)) xor (inputs(56)));
    layer0_outputs(2986) <= (inputs(164)) xor (inputs(149));
    layer0_outputs(2987) <= not(inputs(104)) or (inputs(148));
    layer0_outputs(2988) <= inputs(152);
    layer0_outputs(2989) <= not(inputs(58));
    layer0_outputs(2990) <= (inputs(194)) or (inputs(89));
    layer0_outputs(2991) <= (inputs(102)) or (inputs(29));
    layer0_outputs(2992) <= not(inputs(160));
    layer0_outputs(2993) <= (inputs(163)) and not (inputs(165));
    layer0_outputs(2994) <= not(inputs(111)) or (inputs(50));
    layer0_outputs(2995) <= (inputs(141)) xor (inputs(61));
    layer0_outputs(2996) <= not(inputs(168)) or (inputs(234));
    layer0_outputs(2997) <= '1';
    layer0_outputs(2998) <= (inputs(71)) and not (inputs(192));
    layer0_outputs(2999) <= not(inputs(97));
    layer0_outputs(3000) <= not(inputs(121)) or (inputs(92));
    layer0_outputs(3001) <= not(inputs(67));
    layer0_outputs(3002) <= (inputs(118)) and not (inputs(65));
    layer0_outputs(3003) <= '1';
    layer0_outputs(3004) <= (inputs(225)) and (inputs(254));
    layer0_outputs(3005) <= not(inputs(136));
    layer0_outputs(3006) <= not(inputs(174)) or (inputs(59));
    layer0_outputs(3007) <= (inputs(16)) and (inputs(207));
    layer0_outputs(3008) <= '0';
    layer0_outputs(3009) <= not(inputs(125));
    layer0_outputs(3010) <= not(inputs(17)) or (inputs(127));
    layer0_outputs(3011) <= (inputs(141)) and (inputs(1));
    layer0_outputs(3012) <= (inputs(140)) and not (inputs(242));
    layer0_outputs(3013) <= not(inputs(25));
    layer0_outputs(3014) <= (inputs(56)) or (inputs(39));
    layer0_outputs(3015) <= (inputs(196)) or (inputs(189));
    layer0_outputs(3016) <= not((inputs(82)) or (inputs(172)));
    layer0_outputs(3017) <= (inputs(222)) or (inputs(196));
    layer0_outputs(3018) <= (inputs(248)) or (inputs(81));
    layer0_outputs(3019) <= not(inputs(141));
    layer0_outputs(3020) <= (inputs(164)) or (inputs(248));
    layer0_outputs(3021) <= '0';
    layer0_outputs(3022) <= (inputs(18)) and (inputs(29));
    layer0_outputs(3023) <= not((inputs(58)) or (inputs(55)));
    layer0_outputs(3024) <= not((inputs(205)) or (inputs(192)));
    layer0_outputs(3025) <= (inputs(126)) xor (inputs(124));
    layer0_outputs(3026) <= (inputs(202)) or (inputs(24));
    layer0_outputs(3027) <= not(inputs(119)) or (inputs(157));
    layer0_outputs(3028) <= not(inputs(42)) or (inputs(55));
    layer0_outputs(3029) <= '0';
    layer0_outputs(3030) <= inputs(190);
    layer0_outputs(3031) <= '0';
    layer0_outputs(3032) <= not((inputs(134)) or (inputs(108)));
    layer0_outputs(3033) <= inputs(90);
    layer0_outputs(3034) <= (inputs(88)) and not (inputs(70));
    layer0_outputs(3035) <= (inputs(22)) and (inputs(56));
    layer0_outputs(3036) <= (inputs(109)) and not (inputs(42));
    layer0_outputs(3037) <= (inputs(171)) and not (inputs(97));
    layer0_outputs(3038) <= not(inputs(152));
    layer0_outputs(3039) <= not((inputs(236)) or (inputs(138)));
    layer0_outputs(3040) <= not((inputs(27)) or (inputs(197)));
    layer0_outputs(3041) <= (inputs(197)) and not (inputs(239));
    layer0_outputs(3042) <= (inputs(146)) and not (inputs(98));
    layer0_outputs(3043) <= not(inputs(180)) or (inputs(12));
    layer0_outputs(3044) <= not(inputs(151)) or (inputs(169));
    layer0_outputs(3045) <= (inputs(232)) or (inputs(102));
    layer0_outputs(3046) <= not(inputs(36)) or (inputs(144));
    layer0_outputs(3047) <= not((inputs(50)) or (inputs(120)));
    layer0_outputs(3048) <= (inputs(200)) and not (inputs(220));
    layer0_outputs(3049) <= (inputs(124)) xor (inputs(220));
    layer0_outputs(3050) <= (inputs(54)) and not (inputs(48));
    layer0_outputs(3051) <= not((inputs(91)) or (inputs(106)));
    layer0_outputs(3052) <= (inputs(246)) and not (inputs(60));
    layer0_outputs(3053) <= not((inputs(151)) and (inputs(150)));
    layer0_outputs(3054) <= (inputs(82)) and not (inputs(228));
    layer0_outputs(3055) <= not(inputs(87)) or (inputs(221));
    layer0_outputs(3056) <= (inputs(207)) xor (inputs(115));
    layer0_outputs(3057) <= inputs(172);
    layer0_outputs(3058) <= not((inputs(13)) or (inputs(205)));
    layer0_outputs(3059) <= (inputs(185)) and not (inputs(220));
    layer0_outputs(3060) <= not((inputs(198)) or (inputs(222)));
    layer0_outputs(3061) <= (inputs(162)) xor (inputs(51));
    layer0_outputs(3062) <= inputs(171);
    layer0_outputs(3063) <= not(inputs(105));
    layer0_outputs(3064) <= not((inputs(176)) and (inputs(228)));
    layer0_outputs(3065) <= not(inputs(40)) or (inputs(208));
    layer0_outputs(3066) <= (inputs(240)) and not (inputs(71));
    layer0_outputs(3067) <= inputs(36);
    layer0_outputs(3068) <= not((inputs(1)) or (inputs(227)));
    layer0_outputs(3069) <= not((inputs(205)) or (inputs(189)));
    layer0_outputs(3070) <= not(inputs(112));
    layer0_outputs(3071) <= not(inputs(58));
    layer0_outputs(3072) <= (inputs(118)) and not (inputs(179));
    layer0_outputs(3073) <= not((inputs(87)) or (inputs(226)));
    layer0_outputs(3074) <= (inputs(3)) xor (inputs(101));
    layer0_outputs(3075) <= inputs(177);
    layer0_outputs(3076) <= not(inputs(116));
    layer0_outputs(3077) <= (inputs(80)) or (inputs(182));
    layer0_outputs(3078) <= not((inputs(110)) or (inputs(96)));
    layer0_outputs(3079) <= (inputs(48)) and (inputs(190));
    layer0_outputs(3080) <= not((inputs(12)) xor (inputs(85)));
    layer0_outputs(3081) <= (inputs(117)) and not (inputs(82));
    layer0_outputs(3082) <= not((inputs(130)) xor (inputs(36)));
    layer0_outputs(3083) <= (inputs(237)) or (inputs(11));
    layer0_outputs(3084) <= (inputs(170)) and not (inputs(135));
    layer0_outputs(3085) <= not(inputs(124)) or (inputs(3));
    layer0_outputs(3086) <= (inputs(172)) or (inputs(177));
    layer0_outputs(3087) <= not(inputs(89));
    layer0_outputs(3088) <= not((inputs(120)) or (inputs(244)));
    layer0_outputs(3089) <= not(inputs(139));
    layer0_outputs(3090) <= not((inputs(97)) xor (inputs(100)));
    layer0_outputs(3091) <= inputs(195);
    layer0_outputs(3092) <= (inputs(69)) and (inputs(216));
    layer0_outputs(3093) <= (inputs(169)) and not (inputs(23));
    layer0_outputs(3094) <= inputs(10);
    layer0_outputs(3095) <= (inputs(44)) and not (inputs(113));
    layer0_outputs(3096) <= not((inputs(223)) and (inputs(168)));
    layer0_outputs(3097) <= '0';
    layer0_outputs(3098) <= not((inputs(41)) or (inputs(55)));
    layer0_outputs(3099) <= (inputs(87)) and not (inputs(159));
    layer0_outputs(3100) <= (inputs(225)) and not (inputs(131));
    layer0_outputs(3101) <= (inputs(109)) xor (inputs(8));
    layer0_outputs(3102) <= (inputs(84)) and not (inputs(63));
    layer0_outputs(3103) <= not((inputs(20)) xor (inputs(121)));
    layer0_outputs(3104) <= '0';
    layer0_outputs(3105) <= (inputs(66)) and (inputs(98));
    layer0_outputs(3106) <= (inputs(132)) and not (inputs(78));
    layer0_outputs(3107) <= (inputs(84)) and not (inputs(5));
    layer0_outputs(3108) <= not(inputs(38));
    layer0_outputs(3109) <= not(inputs(242)) or (inputs(237));
    layer0_outputs(3110) <= not(inputs(24)) or (inputs(114));
    layer0_outputs(3111) <= (inputs(97)) xor (inputs(229));
    layer0_outputs(3112) <= not((inputs(192)) or (inputs(42)));
    layer0_outputs(3113) <= (inputs(119)) or (inputs(39));
    layer0_outputs(3114) <= not((inputs(225)) or (inputs(101)));
    layer0_outputs(3115) <= (inputs(87)) and not (inputs(68));
    layer0_outputs(3116) <= inputs(144);
    layer0_outputs(3117) <= not(inputs(187)) or (inputs(204));
    layer0_outputs(3118) <= not(inputs(55));
    layer0_outputs(3119) <= not(inputs(249)) or (inputs(245));
    layer0_outputs(3120) <= inputs(219);
    layer0_outputs(3121) <= not(inputs(114));
    layer0_outputs(3122) <= inputs(228);
    layer0_outputs(3123) <= not((inputs(54)) or (inputs(82)));
    layer0_outputs(3124) <= inputs(86);
    layer0_outputs(3125) <= not(inputs(232)) or (inputs(196));
    layer0_outputs(3126) <= not(inputs(235));
    layer0_outputs(3127) <= (inputs(151)) and not (inputs(31));
    layer0_outputs(3128) <= not((inputs(11)) or (inputs(244)));
    layer0_outputs(3129) <= not(inputs(156)) or (inputs(111));
    layer0_outputs(3130) <= (inputs(143)) xor (inputs(71));
    layer0_outputs(3131) <= (inputs(125)) or (inputs(4));
    layer0_outputs(3132) <= (inputs(117)) xor (inputs(100));
    layer0_outputs(3133) <= not(inputs(171)) or (inputs(161));
    layer0_outputs(3134) <= not((inputs(210)) or (inputs(28)));
    layer0_outputs(3135) <= not(inputs(184)) or (inputs(58));
    layer0_outputs(3136) <= (inputs(92)) xor (inputs(253));
    layer0_outputs(3137) <= (inputs(22)) xor (inputs(237));
    layer0_outputs(3138) <= not(inputs(18));
    layer0_outputs(3139) <= not(inputs(218)) or (inputs(255));
    layer0_outputs(3140) <= (inputs(193)) or (inputs(155));
    layer0_outputs(3141) <= not(inputs(249));
    layer0_outputs(3142) <= inputs(26);
    layer0_outputs(3143) <= not(inputs(156)) or (inputs(231));
    layer0_outputs(3144) <= not((inputs(124)) or (inputs(122)));
    layer0_outputs(3145) <= inputs(91);
    layer0_outputs(3146) <= inputs(214);
    layer0_outputs(3147) <= (inputs(79)) and not (inputs(130));
    layer0_outputs(3148) <= inputs(166);
    layer0_outputs(3149) <= inputs(140);
    layer0_outputs(3150) <= not((inputs(108)) xor (inputs(112)));
    layer0_outputs(3151) <= inputs(196);
    layer0_outputs(3152) <= inputs(254);
    layer0_outputs(3153) <= not(inputs(127)) or (inputs(1));
    layer0_outputs(3154) <= (inputs(222)) xor (inputs(28));
    layer0_outputs(3155) <= not((inputs(110)) and (inputs(175)));
    layer0_outputs(3156) <= not(inputs(140)) or (inputs(208));
    layer0_outputs(3157) <= inputs(116);
    layer0_outputs(3158) <= not(inputs(146)) or (inputs(15));
    layer0_outputs(3159) <= inputs(229);
    layer0_outputs(3160) <= (inputs(194)) or (inputs(64));
    layer0_outputs(3161) <= not(inputs(74));
    layer0_outputs(3162) <= '1';
    layer0_outputs(3163) <= not((inputs(39)) xor (inputs(87)));
    layer0_outputs(3164) <= (inputs(151)) xor (inputs(112));
    layer0_outputs(3165) <= not((inputs(73)) or (inputs(25)));
    layer0_outputs(3166) <= (inputs(241)) or (inputs(68));
    layer0_outputs(3167) <= not(inputs(13));
    layer0_outputs(3168) <= (inputs(123)) or (inputs(189));
    layer0_outputs(3169) <= (inputs(32)) and not (inputs(117));
    layer0_outputs(3170) <= not((inputs(207)) or (inputs(226)));
    layer0_outputs(3171) <= inputs(150);
    layer0_outputs(3172) <= (inputs(173)) and not (inputs(11));
    layer0_outputs(3173) <= inputs(72);
    layer0_outputs(3174) <= (inputs(128)) or (inputs(119));
    layer0_outputs(3175) <= (inputs(155)) and not (inputs(174));
    layer0_outputs(3176) <= not((inputs(41)) or (inputs(46)));
    layer0_outputs(3177) <= not(inputs(136));
    layer0_outputs(3178) <= not(inputs(232));
    layer0_outputs(3179) <= (inputs(94)) and not (inputs(160));
    layer0_outputs(3180) <= (inputs(3)) and not (inputs(236));
    layer0_outputs(3181) <= inputs(179);
    layer0_outputs(3182) <= '1';
    layer0_outputs(3183) <= inputs(65);
    layer0_outputs(3184) <= inputs(104);
    layer0_outputs(3185) <= not(inputs(207));
    layer0_outputs(3186) <= (inputs(215)) or (inputs(95));
    layer0_outputs(3187) <= '1';
    layer0_outputs(3188) <= not((inputs(189)) or (inputs(166)));
    layer0_outputs(3189) <= inputs(30);
    layer0_outputs(3190) <= not(inputs(89)) or (inputs(158));
    layer0_outputs(3191) <= not(inputs(183));
    layer0_outputs(3192) <= not(inputs(222)) or (inputs(204));
    layer0_outputs(3193) <= inputs(156);
    layer0_outputs(3194) <= not(inputs(52));
    layer0_outputs(3195) <= (inputs(118)) or (inputs(143));
    layer0_outputs(3196) <= not((inputs(153)) or (inputs(240)));
    layer0_outputs(3197) <= not((inputs(233)) xor (inputs(78)));
    layer0_outputs(3198) <= '1';
    layer0_outputs(3199) <= not((inputs(6)) or (inputs(83)));
    layer0_outputs(3200) <= (inputs(148)) and (inputs(0));
    layer0_outputs(3201) <= not((inputs(37)) xor (inputs(148)));
    layer0_outputs(3202) <= (inputs(120)) xor (inputs(46));
    layer0_outputs(3203) <= (inputs(92)) or (inputs(93));
    layer0_outputs(3204) <= not((inputs(146)) xor (inputs(254)));
    layer0_outputs(3205) <= inputs(110);
    layer0_outputs(3206) <= inputs(58);
    layer0_outputs(3207) <= (inputs(190)) or (inputs(168));
    layer0_outputs(3208) <= not(inputs(130)) or (inputs(95));
    layer0_outputs(3209) <= not(inputs(120));
    layer0_outputs(3210) <= (inputs(44)) and (inputs(32));
    layer0_outputs(3211) <= not(inputs(103)) or (inputs(107));
    layer0_outputs(3212) <= not(inputs(222));
    layer0_outputs(3213) <= not((inputs(19)) and (inputs(16)));
    layer0_outputs(3214) <= (inputs(66)) and (inputs(144));
    layer0_outputs(3215) <= not((inputs(57)) or (inputs(229)));
    layer0_outputs(3216) <= not(inputs(153));
    layer0_outputs(3217) <= not(inputs(153)) or (inputs(246));
    layer0_outputs(3218) <= inputs(149);
    layer0_outputs(3219) <= not(inputs(136));
    layer0_outputs(3220) <= inputs(197);
    layer0_outputs(3221) <= not(inputs(85));
    layer0_outputs(3222) <= not((inputs(34)) or (inputs(73)));
    layer0_outputs(3223) <= (inputs(59)) or (inputs(37));
    layer0_outputs(3224) <= (inputs(86)) xor (inputs(192));
    layer0_outputs(3225) <= inputs(190);
    layer0_outputs(3226) <= not(inputs(217));
    layer0_outputs(3227) <= '1';
    layer0_outputs(3228) <= inputs(54);
    layer0_outputs(3229) <= not(inputs(237));
    layer0_outputs(3230) <= (inputs(183)) xor (inputs(249));
    layer0_outputs(3231) <= (inputs(205)) or (inputs(104));
    layer0_outputs(3232) <= '0';
    layer0_outputs(3233) <= (inputs(125)) or (inputs(173));
    layer0_outputs(3234) <= inputs(61);
    layer0_outputs(3235) <= (inputs(217)) and not (inputs(29));
    layer0_outputs(3236) <= not(inputs(229)) or (inputs(66));
    layer0_outputs(3237) <= (inputs(19)) and not (inputs(115));
    layer0_outputs(3238) <= (inputs(4)) or (inputs(183));
    layer0_outputs(3239) <= not(inputs(225));
    layer0_outputs(3240) <= (inputs(100)) or (inputs(54));
    layer0_outputs(3241) <= not((inputs(166)) or (inputs(209)));
    layer0_outputs(3242) <= not((inputs(185)) or (inputs(55)));
    layer0_outputs(3243) <= not(inputs(72)) or (inputs(32));
    layer0_outputs(3244) <= not(inputs(44));
    layer0_outputs(3245) <= not((inputs(21)) or (inputs(200)));
    layer0_outputs(3246) <= (inputs(95)) xor (inputs(3));
    layer0_outputs(3247) <= (inputs(0)) or (inputs(93));
    layer0_outputs(3248) <= not(inputs(37));
    layer0_outputs(3249) <= not((inputs(178)) xor (inputs(8)));
    layer0_outputs(3250) <= (inputs(232)) and (inputs(139));
    layer0_outputs(3251) <= (inputs(170)) or (inputs(248));
    layer0_outputs(3252) <= (inputs(152)) and not (inputs(162));
    layer0_outputs(3253) <= (inputs(153)) and not (inputs(83));
    layer0_outputs(3254) <= not((inputs(244)) xor (inputs(78)));
    layer0_outputs(3255) <= not(inputs(72));
    layer0_outputs(3256) <= (inputs(44)) or (inputs(28));
    layer0_outputs(3257) <= (inputs(100)) or (inputs(230));
    layer0_outputs(3258) <= (inputs(200)) or (inputs(113));
    layer0_outputs(3259) <= not((inputs(125)) or (inputs(146)));
    layer0_outputs(3260) <= '0';
    layer0_outputs(3261) <= (inputs(154)) and not (inputs(22));
    layer0_outputs(3262) <= not(inputs(210));
    layer0_outputs(3263) <= not(inputs(55)) or (inputs(191));
    layer0_outputs(3264) <= (inputs(173)) and (inputs(224));
    layer0_outputs(3265) <= not(inputs(150));
    layer0_outputs(3266) <= (inputs(107)) or (inputs(175));
    layer0_outputs(3267) <= not(inputs(236));
    layer0_outputs(3268) <= not((inputs(128)) and (inputs(110)));
    layer0_outputs(3269) <= not((inputs(198)) or (inputs(36)));
    layer0_outputs(3270) <= not(inputs(67));
    layer0_outputs(3271) <= not(inputs(117));
    layer0_outputs(3272) <= (inputs(103)) xor (inputs(22));
    layer0_outputs(3273) <= not(inputs(167));
    layer0_outputs(3274) <= (inputs(186)) and not (inputs(89));
    layer0_outputs(3275) <= not(inputs(80));
    layer0_outputs(3276) <= (inputs(129)) xor (inputs(225));
    layer0_outputs(3277) <= (inputs(187)) and not (inputs(75));
    layer0_outputs(3278) <= (inputs(215)) or (inputs(232));
    layer0_outputs(3279) <= (inputs(165)) and not (inputs(5));
    layer0_outputs(3280) <= (inputs(110)) and (inputs(229));
    layer0_outputs(3281) <= not(inputs(154));
    layer0_outputs(3282) <= not(inputs(104)) or (inputs(208));
    layer0_outputs(3283) <= (inputs(164)) and not (inputs(25));
    layer0_outputs(3284) <= (inputs(107)) and (inputs(20));
    layer0_outputs(3285) <= not(inputs(152)) or (inputs(42));
    layer0_outputs(3286) <= (inputs(173)) and not (inputs(206));
    layer0_outputs(3287) <= not(inputs(40));
    layer0_outputs(3288) <= not((inputs(174)) or (inputs(26)));
    layer0_outputs(3289) <= (inputs(240)) and not (inputs(254));
    layer0_outputs(3290) <= (inputs(49)) xor (inputs(166));
    layer0_outputs(3291) <= '1';
    layer0_outputs(3292) <= '0';
    layer0_outputs(3293) <= not(inputs(82)) or (inputs(143));
    layer0_outputs(3294) <= not((inputs(246)) and (inputs(2)));
    layer0_outputs(3295) <= (inputs(161)) and not (inputs(45));
    layer0_outputs(3296) <= not((inputs(181)) xor (inputs(35)));
    layer0_outputs(3297) <= not(inputs(240)) or (inputs(46));
    layer0_outputs(3298) <= (inputs(190)) xor (inputs(123));
    layer0_outputs(3299) <= not(inputs(97));
    layer0_outputs(3300) <= inputs(37);
    layer0_outputs(3301) <= not(inputs(141)) or (inputs(205));
    layer0_outputs(3302) <= (inputs(65)) and not (inputs(62));
    layer0_outputs(3303) <= '1';
    layer0_outputs(3304) <= not(inputs(87)) or (inputs(168));
    layer0_outputs(3305) <= (inputs(31)) or (inputs(181));
    layer0_outputs(3306) <= (inputs(163)) or (inputs(83));
    layer0_outputs(3307) <= not(inputs(77)) or (inputs(127));
    layer0_outputs(3308) <= (inputs(129)) xor (inputs(105));
    layer0_outputs(3309) <= inputs(96);
    layer0_outputs(3310) <= (inputs(233)) or (inputs(91));
    layer0_outputs(3311) <= (inputs(154)) or (inputs(229));
    layer0_outputs(3312) <= '0';
    layer0_outputs(3313) <= not(inputs(124));
    layer0_outputs(3314) <= (inputs(217)) or (inputs(197));
    layer0_outputs(3315) <= not(inputs(78));
    layer0_outputs(3316) <= not(inputs(218));
    layer0_outputs(3317) <= (inputs(194)) or (inputs(162));
    layer0_outputs(3318) <= (inputs(81)) or (inputs(216));
    layer0_outputs(3319) <= inputs(118);
    layer0_outputs(3320) <= inputs(175);
    layer0_outputs(3321) <= (inputs(60)) and not (inputs(5));
    layer0_outputs(3322) <= (inputs(93)) and (inputs(27));
    layer0_outputs(3323) <= (inputs(106)) xor (inputs(14));
    layer0_outputs(3324) <= (inputs(0)) or (inputs(197));
    layer0_outputs(3325) <= '0';
    layer0_outputs(3326) <= inputs(76);
    layer0_outputs(3327) <= (inputs(3)) and not (inputs(165));
    layer0_outputs(3328) <= (inputs(254)) or (inputs(26));
    layer0_outputs(3329) <= '0';
    layer0_outputs(3330) <= (inputs(186)) or (inputs(229));
    layer0_outputs(3331) <= not((inputs(203)) or (inputs(119)));
    layer0_outputs(3332) <= not(inputs(108));
    layer0_outputs(3333) <= (inputs(86)) and not (inputs(111));
    layer0_outputs(3334) <= '1';
    layer0_outputs(3335) <= (inputs(212)) xor (inputs(224));
    layer0_outputs(3336) <= not((inputs(17)) and (inputs(112)));
    layer0_outputs(3337) <= '0';
    layer0_outputs(3338) <= (inputs(16)) and not (inputs(219));
    layer0_outputs(3339) <= not((inputs(241)) xor (inputs(101)));
    layer0_outputs(3340) <= (inputs(184)) or (inputs(75));
    layer0_outputs(3341) <= inputs(165);
    layer0_outputs(3342) <= not(inputs(149));
    layer0_outputs(3343) <= not(inputs(104));
    layer0_outputs(3344) <= (inputs(52)) xor (inputs(84));
    layer0_outputs(3345) <= not(inputs(77)) or (inputs(250));
    layer0_outputs(3346) <= '0';
    layer0_outputs(3347) <= not(inputs(71));
    layer0_outputs(3348) <= (inputs(139)) and not (inputs(50));
    layer0_outputs(3349) <= not(inputs(232));
    layer0_outputs(3350) <= inputs(58);
    layer0_outputs(3351) <= (inputs(173)) and not (inputs(111));
    layer0_outputs(3352) <= '0';
    layer0_outputs(3353) <= (inputs(230)) and not (inputs(78));
    layer0_outputs(3354) <= (inputs(227)) or (inputs(192));
    layer0_outputs(3355) <= not(inputs(107));
    layer0_outputs(3356) <= '0';
    layer0_outputs(3357) <= not((inputs(59)) or (inputs(77)));
    layer0_outputs(3358) <= (inputs(245)) and (inputs(50));
    layer0_outputs(3359) <= not((inputs(48)) xor (inputs(180)));
    layer0_outputs(3360) <= (inputs(59)) xor (inputs(192));
    layer0_outputs(3361) <= not((inputs(20)) and (inputs(197)));
    layer0_outputs(3362) <= not(inputs(220)) or (inputs(34));
    layer0_outputs(3363) <= not((inputs(165)) or (inputs(236)));
    layer0_outputs(3364) <= not((inputs(75)) xor (inputs(209)));
    layer0_outputs(3365) <= not(inputs(12));
    layer0_outputs(3366) <= not(inputs(226));
    layer0_outputs(3367) <= inputs(97);
    layer0_outputs(3368) <= (inputs(141)) xor (inputs(50));
    layer0_outputs(3369) <= (inputs(193)) or (inputs(225));
    layer0_outputs(3370) <= (inputs(49)) or (inputs(58));
    layer0_outputs(3371) <= (inputs(132)) or (inputs(251));
    layer0_outputs(3372) <= not((inputs(112)) or (inputs(160)));
    layer0_outputs(3373) <= (inputs(177)) or (inputs(43));
    layer0_outputs(3374) <= (inputs(85)) xor (inputs(11));
    layer0_outputs(3375) <= (inputs(204)) and (inputs(109));
    layer0_outputs(3376) <= not((inputs(18)) xor (inputs(221)));
    layer0_outputs(3377) <= not(inputs(12));
    layer0_outputs(3378) <= not(inputs(100));
    layer0_outputs(3379) <= not(inputs(77));
    layer0_outputs(3380) <= inputs(213);
    layer0_outputs(3381) <= (inputs(82)) or (inputs(61));
    layer0_outputs(3382) <= (inputs(142)) and not (inputs(170));
    layer0_outputs(3383) <= (inputs(160)) xor (inputs(109));
    layer0_outputs(3384) <= inputs(17);
    layer0_outputs(3385) <= inputs(122);
    layer0_outputs(3386) <= not((inputs(42)) xor (inputs(72)));
    layer0_outputs(3387) <= (inputs(158)) and (inputs(167));
    layer0_outputs(3388) <= not(inputs(35)) or (inputs(24));
    layer0_outputs(3389) <= (inputs(156)) or (inputs(196));
    layer0_outputs(3390) <= (inputs(156)) and not (inputs(73));
    layer0_outputs(3391) <= '1';
    layer0_outputs(3392) <= inputs(61);
    layer0_outputs(3393) <= (inputs(249)) or (inputs(233));
    layer0_outputs(3394) <= (inputs(171)) or (inputs(60));
    layer0_outputs(3395) <= inputs(146);
    layer0_outputs(3396) <= not(inputs(103)) or (inputs(113));
    layer0_outputs(3397) <= (inputs(27)) xor (inputs(162));
    layer0_outputs(3398) <= not(inputs(154));
    layer0_outputs(3399) <= not((inputs(214)) xor (inputs(112)));
    layer0_outputs(3400) <= not((inputs(40)) or (inputs(142)));
    layer0_outputs(3401) <= (inputs(24)) and (inputs(223));
    layer0_outputs(3402) <= not(inputs(117));
    layer0_outputs(3403) <= (inputs(66)) or (inputs(191));
    layer0_outputs(3404) <= (inputs(19)) and not (inputs(248));
    layer0_outputs(3405) <= not((inputs(97)) or (inputs(184)));
    layer0_outputs(3406) <= (inputs(202)) and not (inputs(130));
    layer0_outputs(3407) <= not(inputs(85));
    layer0_outputs(3408) <= not((inputs(175)) or (inputs(247)));
    layer0_outputs(3409) <= inputs(66);
    layer0_outputs(3410) <= not((inputs(234)) or (inputs(228)));
    layer0_outputs(3411) <= (inputs(69)) and (inputs(17));
    layer0_outputs(3412) <= not(inputs(106)) or (inputs(230));
    layer0_outputs(3413) <= not((inputs(30)) or (inputs(166)));
    layer0_outputs(3414) <= not(inputs(44)) or (inputs(249));
    layer0_outputs(3415) <= not((inputs(232)) or (inputs(21)));
    layer0_outputs(3416) <= not(inputs(106));
    layer0_outputs(3417) <= not((inputs(24)) or (inputs(63)));
    layer0_outputs(3418) <= not((inputs(150)) or (inputs(115)));
    layer0_outputs(3419) <= (inputs(123)) and (inputs(163));
    layer0_outputs(3420) <= (inputs(167)) and not (inputs(130));
    layer0_outputs(3421) <= (inputs(140)) or (inputs(133));
    layer0_outputs(3422) <= inputs(160);
    layer0_outputs(3423) <= not((inputs(32)) or (inputs(89)));
    layer0_outputs(3424) <= not(inputs(31));
    layer0_outputs(3425) <= (inputs(173)) xor (inputs(222));
    layer0_outputs(3426) <= not((inputs(24)) or (inputs(142)));
    layer0_outputs(3427) <= '1';
    layer0_outputs(3428) <= not(inputs(121)) or (inputs(203));
    layer0_outputs(3429) <= not(inputs(240)) or (inputs(69));
    layer0_outputs(3430) <= not(inputs(197));
    layer0_outputs(3431) <= not((inputs(115)) xor (inputs(84)));
    layer0_outputs(3432) <= (inputs(168)) or (inputs(20));
    layer0_outputs(3433) <= not(inputs(100));
    layer0_outputs(3434) <= not((inputs(211)) or (inputs(125)));
    layer0_outputs(3435) <= not((inputs(147)) xor (inputs(139)));
    layer0_outputs(3436) <= not((inputs(8)) xor (inputs(163)));
    layer0_outputs(3437) <= (inputs(12)) or (inputs(56));
    layer0_outputs(3438) <= (inputs(45)) or (inputs(162));
    layer0_outputs(3439) <= (inputs(56)) and not (inputs(5));
    layer0_outputs(3440) <= (inputs(159)) and not (inputs(245));
    layer0_outputs(3441) <= not(inputs(57));
    layer0_outputs(3442) <= not(inputs(55)) or (inputs(117));
    layer0_outputs(3443) <= '1';
    layer0_outputs(3444) <= (inputs(160)) or (inputs(106));
    layer0_outputs(3445) <= (inputs(248)) or (inputs(105));
    layer0_outputs(3446) <= (inputs(180)) or (inputs(186));
    layer0_outputs(3447) <= not((inputs(43)) or (inputs(81)));
    layer0_outputs(3448) <= not((inputs(210)) and (inputs(64)));
    layer0_outputs(3449) <= (inputs(100)) and not (inputs(177));
    layer0_outputs(3450) <= not((inputs(250)) or (inputs(242)));
    layer0_outputs(3451) <= inputs(115);
    layer0_outputs(3452) <= not(inputs(150)) or (inputs(207));
    layer0_outputs(3453) <= inputs(116);
    layer0_outputs(3454) <= not(inputs(10));
    layer0_outputs(3455) <= (inputs(110)) and not (inputs(236));
    layer0_outputs(3456) <= '1';
    layer0_outputs(3457) <= not((inputs(47)) xor (inputs(129)));
    layer0_outputs(3458) <= not(inputs(159)) or (inputs(50));
    layer0_outputs(3459) <= not((inputs(55)) or (inputs(172)));
    layer0_outputs(3460) <= (inputs(221)) and not (inputs(147));
    layer0_outputs(3461) <= not(inputs(195));
    layer0_outputs(3462) <= (inputs(18)) and (inputs(6));
    layer0_outputs(3463) <= '0';
    layer0_outputs(3464) <= (inputs(26)) or (inputs(121));
    layer0_outputs(3465) <= not((inputs(181)) or (inputs(59)));
    layer0_outputs(3466) <= not((inputs(151)) or (inputs(135)));
    layer0_outputs(3467) <= not(inputs(26));
    layer0_outputs(3468) <= (inputs(132)) and not (inputs(169));
    layer0_outputs(3469) <= (inputs(10)) and not (inputs(202));
    layer0_outputs(3470) <= (inputs(159)) and not (inputs(199));
    layer0_outputs(3471) <= not(inputs(107)) or (inputs(98));
    layer0_outputs(3472) <= not(inputs(152));
    layer0_outputs(3473) <= not((inputs(233)) xor (inputs(63)));
    layer0_outputs(3474) <= (inputs(107)) and not (inputs(2));
    layer0_outputs(3475) <= (inputs(148)) and not (inputs(48));
    layer0_outputs(3476) <= not(inputs(149));
    layer0_outputs(3477) <= '0';
    layer0_outputs(3478) <= not((inputs(105)) or (inputs(241)));
    layer0_outputs(3479) <= '0';
    layer0_outputs(3480) <= not((inputs(173)) and (inputs(159)));
    layer0_outputs(3481) <= not(inputs(174)) or (inputs(222));
    layer0_outputs(3482) <= not((inputs(98)) or (inputs(31)));
    layer0_outputs(3483) <= '0';
    layer0_outputs(3484) <= (inputs(168)) xor (inputs(175));
    layer0_outputs(3485) <= (inputs(129)) and not (inputs(50));
    layer0_outputs(3486) <= (inputs(151)) xor (inputs(62));
    layer0_outputs(3487) <= inputs(245);
    layer0_outputs(3488) <= (inputs(216)) and not (inputs(206));
    layer0_outputs(3489) <= not((inputs(91)) and (inputs(62)));
    layer0_outputs(3490) <= (inputs(126)) or (inputs(73));
    layer0_outputs(3491) <= not((inputs(131)) xor (inputs(122)));
    layer0_outputs(3492) <= '0';
    layer0_outputs(3493) <= not(inputs(212));
    layer0_outputs(3494) <= not((inputs(25)) xor (inputs(156)));
    layer0_outputs(3495) <= '1';
    layer0_outputs(3496) <= not(inputs(18)) or (inputs(211));
    layer0_outputs(3497) <= (inputs(117)) or (inputs(221));
    layer0_outputs(3498) <= '0';
    layer0_outputs(3499) <= not(inputs(247)) or (inputs(91));
    layer0_outputs(3500) <= inputs(140);
    layer0_outputs(3501) <= not(inputs(86)) or (inputs(187));
    layer0_outputs(3502) <= not((inputs(235)) xor (inputs(12)));
    layer0_outputs(3503) <= (inputs(109)) xor (inputs(79));
    layer0_outputs(3504) <= inputs(15);
    layer0_outputs(3505) <= '0';
    layer0_outputs(3506) <= (inputs(30)) xor (inputs(123));
    layer0_outputs(3507) <= not(inputs(65));
    layer0_outputs(3508) <= '1';
    layer0_outputs(3509) <= not(inputs(58));
    layer0_outputs(3510) <= not(inputs(152)) or (inputs(180));
    layer0_outputs(3511) <= not(inputs(38)) or (inputs(145));
    layer0_outputs(3512) <= not((inputs(99)) or (inputs(64)));
    layer0_outputs(3513) <= (inputs(239)) or (inputs(234));
    layer0_outputs(3514) <= inputs(237);
    layer0_outputs(3515) <= not((inputs(250)) and (inputs(70)));
    layer0_outputs(3516) <= not(inputs(153));
    layer0_outputs(3517) <= (inputs(118)) and not (inputs(2));
    layer0_outputs(3518) <= (inputs(156)) xor (inputs(18));
    layer0_outputs(3519) <= (inputs(13)) and not (inputs(44));
    layer0_outputs(3520) <= (inputs(240)) or (inputs(246));
    layer0_outputs(3521) <= (inputs(5)) or (inputs(220));
    layer0_outputs(3522) <= inputs(118);
    layer0_outputs(3523) <= inputs(184);
    layer0_outputs(3524) <= not((inputs(253)) or (inputs(97)));
    layer0_outputs(3525) <= (inputs(80)) or (inputs(94));
    layer0_outputs(3526) <= inputs(147);
    layer0_outputs(3527) <= not((inputs(189)) xor (inputs(157)));
    layer0_outputs(3528) <= (inputs(202)) and not (inputs(192));
    layer0_outputs(3529) <= (inputs(46)) xor (inputs(83));
    layer0_outputs(3530) <= not((inputs(11)) or (inputs(252)));
    layer0_outputs(3531) <= not(inputs(101)) or (inputs(217));
    layer0_outputs(3532) <= not((inputs(141)) or (inputs(65)));
    layer0_outputs(3533) <= not(inputs(38));
    layer0_outputs(3534) <= (inputs(109)) xor (inputs(65));
    layer0_outputs(3535) <= (inputs(35)) and not (inputs(239));
    layer0_outputs(3536) <= not(inputs(98)) or (inputs(8));
    layer0_outputs(3537) <= not((inputs(187)) or (inputs(27)));
    layer0_outputs(3538) <= not((inputs(177)) xor (inputs(104)));
    layer0_outputs(3539) <= not((inputs(17)) xor (inputs(103)));
    layer0_outputs(3540) <= (inputs(199)) and not (inputs(30));
    layer0_outputs(3541) <= not(inputs(135));
    layer0_outputs(3542) <= (inputs(134)) and not (inputs(240));
    layer0_outputs(3543) <= not((inputs(220)) or (inputs(99)));
    layer0_outputs(3544) <= '0';
    layer0_outputs(3545) <= (inputs(2)) or (inputs(165));
    layer0_outputs(3546) <= (inputs(137)) and not (inputs(193));
    layer0_outputs(3547) <= (inputs(137)) xor (inputs(53));
    layer0_outputs(3548) <= inputs(197);
    layer0_outputs(3549) <= not((inputs(8)) xor (inputs(49)));
    layer0_outputs(3550) <= inputs(245);
    layer0_outputs(3551) <= '1';
    layer0_outputs(3552) <= inputs(120);
    layer0_outputs(3553) <= '0';
    layer0_outputs(3554) <= not((inputs(76)) or (inputs(164)));
    layer0_outputs(3555) <= inputs(132);
    layer0_outputs(3556) <= (inputs(10)) and not (inputs(238));
    layer0_outputs(3557) <= inputs(107);
    layer0_outputs(3558) <= not(inputs(231));
    layer0_outputs(3559) <= '0';
    layer0_outputs(3560) <= not(inputs(103)) or (inputs(81));
    layer0_outputs(3561) <= not(inputs(153));
    layer0_outputs(3562) <= (inputs(157)) xor (inputs(196));
    layer0_outputs(3563) <= inputs(202);
    layer0_outputs(3564) <= (inputs(41)) and not (inputs(77));
    layer0_outputs(3565) <= not(inputs(228)) or (inputs(94));
    layer0_outputs(3566) <= (inputs(188)) or (inputs(92));
    layer0_outputs(3567) <= inputs(174);
    layer0_outputs(3568) <= inputs(196);
    layer0_outputs(3569) <= (inputs(251)) xor (inputs(22));
    layer0_outputs(3570) <= '1';
    layer0_outputs(3571) <= not(inputs(242)) or (inputs(80));
    layer0_outputs(3572) <= not(inputs(106)) or (inputs(174));
    layer0_outputs(3573) <= not(inputs(199));
    layer0_outputs(3574) <= (inputs(226)) and not (inputs(56));
    layer0_outputs(3575) <= not((inputs(45)) xor (inputs(206)));
    layer0_outputs(3576) <= not(inputs(127));
    layer0_outputs(3577) <= not(inputs(105)) or (inputs(119));
    layer0_outputs(3578) <= not(inputs(162));
    layer0_outputs(3579) <= not(inputs(129)) or (inputs(136));
    layer0_outputs(3580) <= inputs(106);
    layer0_outputs(3581) <= not((inputs(234)) or (inputs(116)));
    layer0_outputs(3582) <= '1';
    layer0_outputs(3583) <= not(inputs(190)) or (inputs(209));
    layer0_outputs(3584) <= not(inputs(243));
    layer0_outputs(3585) <= not(inputs(73)) or (inputs(81));
    layer0_outputs(3586) <= not(inputs(165)) or (inputs(94));
    layer0_outputs(3587) <= inputs(136);
    layer0_outputs(3588) <= inputs(102);
    layer0_outputs(3589) <= (inputs(30)) or (inputs(249));
    layer0_outputs(3590) <= (inputs(32)) or (inputs(232));
    layer0_outputs(3591) <= inputs(133);
    layer0_outputs(3592) <= not(inputs(241));
    layer0_outputs(3593) <= (inputs(68)) and (inputs(59));
    layer0_outputs(3594) <= (inputs(81)) and (inputs(38));
    layer0_outputs(3595) <= not(inputs(138)) or (inputs(39));
    layer0_outputs(3596) <= not(inputs(2)) or (inputs(75));
    layer0_outputs(3597) <= not(inputs(102));
    layer0_outputs(3598) <= not(inputs(190));
    layer0_outputs(3599) <= (inputs(231)) xor (inputs(226));
    layer0_outputs(3600) <= inputs(71);
    layer0_outputs(3601) <= inputs(142);
    layer0_outputs(3602) <= not(inputs(98));
    layer0_outputs(3603) <= (inputs(54)) and (inputs(183));
    layer0_outputs(3604) <= inputs(215);
    layer0_outputs(3605) <= (inputs(141)) and not (inputs(145));
    layer0_outputs(3606) <= inputs(33);
    layer0_outputs(3607) <= not(inputs(59)) or (inputs(145));
    layer0_outputs(3608) <= '1';
    layer0_outputs(3609) <= not((inputs(249)) xor (inputs(206)));
    layer0_outputs(3610) <= (inputs(60)) or (inputs(145));
    layer0_outputs(3611) <= (inputs(37)) or (inputs(68));
    layer0_outputs(3612) <= not(inputs(0));
    layer0_outputs(3613) <= (inputs(104)) and not (inputs(203));
    layer0_outputs(3614) <= (inputs(206)) and not (inputs(195));
    layer0_outputs(3615) <= (inputs(204)) xor (inputs(166));
    layer0_outputs(3616) <= not(inputs(102));
    layer0_outputs(3617) <= not(inputs(153)) or (inputs(184));
    layer0_outputs(3618) <= inputs(85);
    layer0_outputs(3619) <= '1';
    layer0_outputs(3620) <= not(inputs(90));
    layer0_outputs(3621) <= '0';
    layer0_outputs(3622) <= inputs(19);
    layer0_outputs(3623) <= not((inputs(232)) xor (inputs(15)));
    layer0_outputs(3624) <= not((inputs(189)) xor (inputs(120)));
    layer0_outputs(3625) <= (inputs(161)) and (inputs(207));
    layer0_outputs(3626) <= not(inputs(22));
    layer0_outputs(3627) <= not(inputs(119));
    layer0_outputs(3628) <= (inputs(146)) and not (inputs(250));
    layer0_outputs(3629) <= (inputs(83)) and not (inputs(113));
    layer0_outputs(3630) <= not(inputs(56)) or (inputs(143));
    layer0_outputs(3631) <= (inputs(183)) and not (inputs(196));
    layer0_outputs(3632) <= not((inputs(26)) or (inputs(167)));
    layer0_outputs(3633) <= not(inputs(199));
    layer0_outputs(3634) <= inputs(198);
    layer0_outputs(3635) <= not(inputs(14)) or (inputs(14));
    layer0_outputs(3636) <= not(inputs(129));
    layer0_outputs(3637) <= not(inputs(249)) or (inputs(54));
    layer0_outputs(3638) <= not(inputs(46));
    layer0_outputs(3639) <= (inputs(179)) or (inputs(148));
    layer0_outputs(3640) <= not(inputs(85));
    layer0_outputs(3641) <= (inputs(94)) and not (inputs(0));
    layer0_outputs(3642) <= not((inputs(251)) xor (inputs(105)));
    layer0_outputs(3643) <= not(inputs(233)) or (inputs(142));
    layer0_outputs(3644) <= not(inputs(164));
    layer0_outputs(3645) <= (inputs(11)) xor (inputs(40));
    layer0_outputs(3646) <= (inputs(15)) xor (inputs(128));
    layer0_outputs(3647) <= inputs(3);
    layer0_outputs(3648) <= not(inputs(35));
    layer0_outputs(3649) <= (inputs(5)) and (inputs(194));
    layer0_outputs(3650) <= (inputs(135)) and not (inputs(55));
    layer0_outputs(3651) <= (inputs(125)) or (inputs(20));
    layer0_outputs(3652) <= not(inputs(175));
    layer0_outputs(3653) <= not((inputs(174)) or (inputs(143)));
    layer0_outputs(3654) <= not(inputs(182)) or (inputs(94));
    layer0_outputs(3655) <= not((inputs(142)) or (inputs(141)));
    layer0_outputs(3656) <= not(inputs(152)) or (inputs(242));
    layer0_outputs(3657) <= '0';
    layer0_outputs(3658) <= inputs(150);
    layer0_outputs(3659) <= (inputs(137)) or (inputs(23));
    layer0_outputs(3660) <= '0';
    layer0_outputs(3661) <= not((inputs(2)) or (inputs(178)));
    layer0_outputs(3662) <= (inputs(167)) and not (inputs(107));
    layer0_outputs(3663) <= not((inputs(176)) xor (inputs(122)));
    layer0_outputs(3664) <= '1';
    layer0_outputs(3665) <= not((inputs(217)) or (inputs(195)));
    layer0_outputs(3666) <= inputs(105);
    layer0_outputs(3667) <= not(inputs(18));
    layer0_outputs(3668) <= (inputs(126)) or (inputs(21));
    layer0_outputs(3669) <= not((inputs(6)) or (inputs(152)));
    layer0_outputs(3670) <= not((inputs(229)) xor (inputs(224)));
    layer0_outputs(3671) <= not(inputs(62)) or (inputs(76));
    layer0_outputs(3672) <= not(inputs(234)) or (inputs(98));
    layer0_outputs(3673) <= (inputs(141)) or (inputs(223));
    layer0_outputs(3674) <= not((inputs(203)) or (inputs(221)));
    layer0_outputs(3675) <= not((inputs(20)) or (inputs(165)));
    layer0_outputs(3676) <= not(inputs(199)) or (inputs(12));
    layer0_outputs(3677) <= (inputs(52)) xor (inputs(77));
    layer0_outputs(3678) <= '1';
    layer0_outputs(3679) <= not(inputs(250)) or (inputs(66));
    layer0_outputs(3680) <= not(inputs(108));
    layer0_outputs(3681) <= inputs(36);
    layer0_outputs(3682) <= not((inputs(84)) xor (inputs(54)));
    layer0_outputs(3683) <= (inputs(220)) and not (inputs(67));
    layer0_outputs(3684) <= not((inputs(160)) xor (inputs(71)));
    layer0_outputs(3685) <= inputs(44);
    layer0_outputs(3686) <= inputs(221);
    layer0_outputs(3687) <= (inputs(199)) xor (inputs(32));
    layer0_outputs(3688) <= (inputs(215)) xor (inputs(161));
    layer0_outputs(3689) <= not((inputs(138)) or (inputs(244)));
    layer0_outputs(3690) <= not(inputs(247));
    layer0_outputs(3691) <= not(inputs(41));
    layer0_outputs(3692) <= not((inputs(43)) or (inputs(254)));
    layer0_outputs(3693) <= (inputs(73)) xor (inputs(76));
    layer0_outputs(3694) <= not(inputs(61)) or (inputs(18));
    layer0_outputs(3695) <= not((inputs(39)) xor (inputs(2)));
    layer0_outputs(3696) <= not((inputs(224)) and (inputs(204)));
    layer0_outputs(3697) <= (inputs(136)) or (inputs(229));
    layer0_outputs(3698) <= inputs(138);
    layer0_outputs(3699) <= not(inputs(86));
    layer0_outputs(3700) <= not(inputs(103)) or (inputs(170));
    layer0_outputs(3701) <= not(inputs(169));
    layer0_outputs(3702) <= (inputs(145)) or (inputs(18));
    layer0_outputs(3703) <= inputs(124);
    layer0_outputs(3704) <= (inputs(26)) xor (inputs(246));
    layer0_outputs(3705) <= (inputs(95)) and not (inputs(13));
    layer0_outputs(3706) <= not(inputs(73)) or (inputs(77));
    layer0_outputs(3707) <= (inputs(83)) or (inputs(123));
    layer0_outputs(3708) <= not((inputs(167)) or (inputs(126)));
    layer0_outputs(3709) <= inputs(139);
    layer0_outputs(3710) <= inputs(91);
    layer0_outputs(3711) <= (inputs(185)) and not (inputs(18));
    layer0_outputs(3712) <= not(inputs(212));
    layer0_outputs(3713) <= (inputs(89)) and not (inputs(109));
    layer0_outputs(3714) <= inputs(191);
    layer0_outputs(3715) <= inputs(132);
    layer0_outputs(3716) <= (inputs(130)) and (inputs(223));
    layer0_outputs(3717) <= not((inputs(47)) or (inputs(103)));
    layer0_outputs(3718) <= inputs(91);
    layer0_outputs(3719) <= not(inputs(167)) or (inputs(60));
    layer0_outputs(3720) <= (inputs(137)) xor (inputs(12));
    layer0_outputs(3721) <= not(inputs(215)) or (inputs(184));
    layer0_outputs(3722) <= not((inputs(239)) or (inputs(138)));
    layer0_outputs(3723) <= (inputs(252)) or (inputs(118));
    layer0_outputs(3724) <= not((inputs(31)) or (inputs(233)));
    layer0_outputs(3725) <= not(inputs(24));
    layer0_outputs(3726) <= not((inputs(73)) xor (inputs(57)));
    layer0_outputs(3727) <= not((inputs(40)) or (inputs(165)));
    layer0_outputs(3728) <= not((inputs(7)) or (inputs(174)));
    layer0_outputs(3729) <= not(inputs(181));
    layer0_outputs(3730) <= (inputs(71)) xor (inputs(226));
    layer0_outputs(3731) <= '0';
    layer0_outputs(3732) <= inputs(20);
    layer0_outputs(3733) <= not((inputs(125)) and (inputs(226)));
    layer0_outputs(3734) <= (inputs(46)) or (inputs(7));
    layer0_outputs(3735) <= (inputs(48)) xor (inputs(192));
    layer0_outputs(3736) <= not(inputs(182));
    layer0_outputs(3737) <= not((inputs(185)) or (inputs(211)));
    layer0_outputs(3738) <= not(inputs(195));
    layer0_outputs(3739) <= not((inputs(106)) or (inputs(251)));
    layer0_outputs(3740) <= (inputs(141)) or (inputs(139));
    layer0_outputs(3741) <= not(inputs(66));
    layer0_outputs(3742) <= (inputs(204)) or (inputs(63));
    layer0_outputs(3743) <= (inputs(62)) and not (inputs(145));
    layer0_outputs(3744) <= (inputs(29)) and (inputs(215));
    layer0_outputs(3745) <= not((inputs(33)) and (inputs(165)));
    layer0_outputs(3746) <= not(inputs(93));
    layer0_outputs(3747) <= not((inputs(225)) and (inputs(208)));
    layer0_outputs(3748) <= inputs(57);
    layer0_outputs(3749) <= not((inputs(151)) or (inputs(128)));
    layer0_outputs(3750) <= not((inputs(71)) and (inputs(217)));
    layer0_outputs(3751) <= not(inputs(18)) or (inputs(21));
    layer0_outputs(3752) <= (inputs(224)) and not (inputs(135));
    layer0_outputs(3753) <= inputs(124);
    layer0_outputs(3754) <= inputs(57);
    layer0_outputs(3755) <= (inputs(44)) or (inputs(182));
    layer0_outputs(3756) <= '0';
    layer0_outputs(3757) <= inputs(58);
    layer0_outputs(3758) <= (inputs(211)) and not (inputs(247));
    layer0_outputs(3759) <= not(inputs(24)) or (inputs(49));
    layer0_outputs(3760) <= not((inputs(185)) or (inputs(174)));
    layer0_outputs(3761) <= not((inputs(94)) or (inputs(225)));
    layer0_outputs(3762) <= (inputs(74)) or (inputs(70));
    layer0_outputs(3763) <= inputs(71);
    layer0_outputs(3764) <= not((inputs(246)) or (inputs(35)));
    layer0_outputs(3765) <= (inputs(140)) and not (inputs(43));
    layer0_outputs(3766) <= (inputs(29)) and not (inputs(238));
    layer0_outputs(3767) <= not(inputs(50));
    layer0_outputs(3768) <= not((inputs(31)) and (inputs(7)));
    layer0_outputs(3769) <= (inputs(209)) or (inputs(41));
    layer0_outputs(3770) <= not(inputs(222)) or (inputs(37));
    layer0_outputs(3771) <= '0';
    layer0_outputs(3772) <= not(inputs(158));
    layer0_outputs(3773) <= not(inputs(203));
    layer0_outputs(3774) <= not(inputs(244)) or (inputs(110));
    layer0_outputs(3775) <= inputs(235);
    layer0_outputs(3776) <= (inputs(105)) and (inputs(6));
    layer0_outputs(3777) <= (inputs(239)) or (inputs(123));
    layer0_outputs(3778) <= inputs(221);
    layer0_outputs(3779) <= (inputs(1)) and (inputs(77));
    layer0_outputs(3780) <= not((inputs(179)) or (inputs(25)));
    layer0_outputs(3781) <= inputs(149);
    layer0_outputs(3782) <= '0';
    layer0_outputs(3783) <= not(inputs(164));
    layer0_outputs(3784) <= not(inputs(70)) or (inputs(143));
    layer0_outputs(3785) <= inputs(27);
    layer0_outputs(3786) <= not((inputs(207)) or (inputs(15)));
    layer0_outputs(3787) <= not(inputs(58));
    layer0_outputs(3788) <= not((inputs(99)) or (inputs(231)));
    layer0_outputs(3789) <= (inputs(75)) or (inputs(64));
    layer0_outputs(3790) <= not((inputs(195)) or (inputs(217)));
    layer0_outputs(3791) <= (inputs(240)) and not (inputs(154));
    layer0_outputs(3792) <= not(inputs(189));
    layer0_outputs(3793) <= inputs(121);
    layer0_outputs(3794) <= not(inputs(64)) or (inputs(211));
    layer0_outputs(3795) <= '0';
    layer0_outputs(3796) <= not(inputs(156)) or (inputs(59));
    layer0_outputs(3797) <= (inputs(82)) or (inputs(38));
    layer0_outputs(3798) <= not(inputs(106));
    layer0_outputs(3799) <= not(inputs(71)) or (inputs(179));
    layer0_outputs(3800) <= not(inputs(149)) or (inputs(84));
    layer0_outputs(3801) <= (inputs(154)) or (inputs(16));
    layer0_outputs(3802) <= inputs(126);
    layer0_outputs(3803) <= not(inputs(228)) or (inputs(35));
    layer0_outputs(3804) <= (inputs(230)) and (inputs(190));
    layer0_outputs(3805) <= inputs(141);
    layer0_outputs(3806) <= inputs(169);
    layer0_outputs(3807) <= (inputs(238)) xor (inputs(117));
    layer0_outputs(3808) <= not(inputs(181)) or (inputs(123));
    layer0_outputs(3809) <= (inputs(18)) or (inputs(90));
    layer0_outputs(3810) <= not((inputs(114)) or (inputs(39)));
    layer0_outputs(3811) <= inputs(179);
    layer0_outputs(3812) <= (inputs(97)) and not (inputs(55));
    layer0_outputs(3813) <= inputs(133);
    layer0_outputs(3814) <= (inputs(99)) and not (inputs(222));
    layer0_outputs(3815) <= inputs(197);
    layer0_outputs(3816) <= (inputs(244)) or (inputs(30));
    layer0_outputs(3817) <= not((inputs(228)) or (inputs(81)));
    layer0_outputs(3818) <= not((inputs(164)) or (inputs(134)));
    layer0_outputs(3819) <= not(inputs(94));
    layer0_outputs(3820) <= (inputs(108)) and not (inputs(30));
    layer0_outputs(3821) <= not(inputs(166));
    layer0_outputs(3822) <= inputs(110);
    layer0_outputs(3823) <= '0';
    layer0_outputs(3824) <= (inputs(26)) and not (inputs(250));
    layer0_outputs(3825) <= not((inputs(51)) or (inputs(239)));
    layer0_outputs(3826) <= not((inputs(20)) or (inputs(64)));
    layer0_outputs(3827) <= inputs(75);
    layer0_outputs(3828) <= not(inputs(166));
    layer0_outputs(3829) <= not((inputs(88)) xor (inputs(212)));
    layer0_outputs(3830) <= (inputs(213)) or (inputs(188));
    layer0_outputs(3831) <= not(inputs(218));
    layer0_outputs(3832) <= (inputs(150)) or (inputs(39));
    layer0_outputs(3833) <= '1';
    layer0_outputs(3834) <= (inputs(11)) and not (inputs(210));
    layer0_outputs(3835) <= not(inputs(103));
    layer0_outputs(3836) <= not(inputs(131)) or (inputs(46));
    layer0_outputs(3837) <= (inputs(247)) or (inputs(195));
    layer0_outputs(3838) <= not(inputs(12)) or (inputs(212));
    layer0_outputs(3839) <= inputs(107);
    layer0_outputs(3840) <= not(inputs(79)) or (inputs(30));
    layer0_outputs(3841) <= not((inputs(38)) or (inputs(235)));
    layer0_outputs(3842) <= inputs(26);
    layer0_outputs(3843) <= (inputs(218)) and not (inputs(59));
    layer0_outputs(3844) <= not((inputs(124)) or (inputs(178)));
    layer0_outputs(3845) <= inputs(160);
    layer0_outputs(3846) <= not((inputs(95)) or (inputs(9)));
    layer0_outputs(3847) <= not(inputs(28));
    layer0_outputs(3848) <= not(inputs(141));
    layer0_outputs(3849) <= (inputs(45)) or (inputs(138));
    layer0_outputs(3850) <= '0';
    layer0_outputs(3851) <= not(inputs(116)) or (inputs(210));
    layer0_outputs(3852) <= not((inputs(101)) or (inputs(12)));
    layer0_outputs(3853) <= (inputs(250)) and not (inputs(52));
    layer0_outputs(3854) <= not(inputs(41));
    layer0_outputs(3855) <= (inputs(103)) or (inputs(64));
    layer0_outputs(3856) <= (inputs(150)) xor (inputs(193));
    layer0_outputs(3857) <= not(inputs(86));
    layer0_outputs(3858) <= inputs(183);
    layer0_outputs(3859) <= (inputs(202)) and not (inputs(114));
    layer0_outputs(3860) <= not((inputs(88)) and (inputs(176)));
    layer0_outputs(3861) <= not((inputs(101)) xor (inputs(96)));
    layer0_outputs(3862) <= (inputs(88)) xor (inputs(253));
    layer0_outputs(3863) <= (inputs(16)) and not (inputs(199));
    layer0_outputs(3864) <= (inputs(77)) xor (inputs(208));
    layer0_outputs(3865) <= not(inputs(224));
    layer0_outputs(3866) <= not((inputs(201)) xor (inputs(65)));
    layer0_outputs(3867) <= (inputs(71)) or (inputs(78));
    layer0_outputs(3868) <= not(inputs(192));
    layer0_outputs(3869) <= inputs(98);
    layer0_outputs(3870) <= inputs(138);
    layer0_outputs(3871) <= not(inputs(202)) or (inputs(24));
    layer0_outputs(3872) <= not(inputs(135));
    layer0_outputs(3873) <= not((inputs(192)) xor (inputs(153)));
    layer0_outputs(3874) <= not((inputs(117)) and (inputs(137)));
    layer0_outputs(3875) <= not((inputs(75)) or (inputs(84)));
    layer0_outputs(3876) <= not(inputs(63));
    layer0_outputs(3877) <= (inputs(201)) and not (inputs(250));
    layer0_outputs(3878) <= (inputs(116)) or (inputs(121));
    layer0_outputs(3879) <= inputs(40);
    layer0_outputs(3880) <= not(inputs(80));
    layer0_outputs(3881) <= (inputs(215)) and not (inputs(52));
    layer0_outputs(3882) <= (inputs(249)) and not (inputs(24));
    layer0_outputs(3883) <= not(inputs(216));
    layer0_outputs(3884) <= (inputs(127)) and (inputs(253));
    layer0_outputs(3885) <= not(inputs(135));
    layer0_outputs(3886) <= (inputs(100)) and not (inputs(205));
    layer0_outputs(3887) <= not((inputs(162)) or (inputs(84)));
    layer0_outputs(3888) <= not((inputs(78)) or (inputs(96)));
    layer0_outputs(3889) <= not(inputs(200)) or (inputs(225));
    layer0_outputs(3890) <= not(inputs(68));
    layer0_outputs(3891) <= (inputs(251)) or (inputs(23));
    layer0_outputs(3892) <= '1';
    layer0_outputs(3893) <= inputs(150);
    layer0_outputs(3894) <= inputs(134);
    layer0_outputs(3895) <= not((inputs(103)) and (inputs(242)));
    layer0_outputs(3896) <= not(inputs(234));
    layer0_outputs(3897) <= not((inputs(23)) or (inputs(74)));
    layer0_outputs(3898) <= not((inputs(97)) xor (inputs(134)));
    layer0_outputs(3899) <= not((inputs(110)) xor (inputs(110)));
    layer0_outputs(3900) <= (inputs(14)) and not (inputs(91));
    layer0_outputs(3901) <= not((inputs(51)) xor (inputs(228)));
    layer0_outputs(3902) <= not(inputs(160)) or (inputs(13));
    layer0_outputs(3903) <= (inputs(239)) or (inputs(145));
    layer0_outputs(3904) <= (inputs(216)) and (inputs(104));
    layer0_outputs(3905) <= (inputs(10)) and not (inputs(45));
    layer0_outputs(3906) <= not(inputs(23));
    layer0_outputs(3907) <= (inputs(48)) or (inputs(115));
    layer0_outputs(3908) <= (inputs(178)) or (inputs(180));
    layer0_outputs(3909) <= not(inputs(221));
    layer0_outputs(3910) <= '0';
    layer0_outputs(3911) <= (inputs(116)) and not (inputs(235));
    layer0_outputs(3912) <= not((inputs(243)) xor (inputs(176)));
    layer0_outputs(3913) <= (inputs(196)) or (inputs(178));
    layer0_outputs(3914) <= (inputs(101)) and not (inputs(156));
    layer0_outputs(3915) <= '0';
    layer0_outputs(3916) <= (inputs(1)) and not (inputs(216));
    layer0_outputs(3917) <= '0';
    layer0_outputs(3918) <= not(inputs(54)) or (inputs(149));
    layer0_outputs(3919) <= not(inputs(59)) or (inputs(146));
    layer0_outputs(3920) <= (inputs(35)) xor (inputs(209));
    layer0_outputs(3921) <= not((inputs(217)) xor (inputs(232)));
    layer0_outputs(3922) <= not((inputs(224)) or (inputs(222)));
    layer0_outputs(3923) <= (inputs(253)) or (inputs(30));
    layer0_outputs(3924) <= (inputs(197)) or (inputs(74));
    layer0_outputs(3925) <= not(inputs(56));
    layer0_outputs(3926) <= not((inputs(169)) or (inputs(228)));
    layer0_outputs(3927) <= inputs(161);
    layer0_outputs(3928) <= (inputs(189)) or (inputs(195));
    layer0_outputs(3929) <= (inputs(2)) xor (inputs(197));
    layer0_outputs(3930) <= not(inputs(96)) or (inputs(24));
    layer0_outputs(3931) <= not(inputs(216));
    layer0_outputs(3932) <= not(inputs(218)) or (inputs(243));
    layer0_outputs(3933) <= not((inputs(228)) or (inputs(233)));
    layer0_outputs(3934) <= not((inputs(236)) or (inputs(198)));
    layer0_outputs(3935) <= inputs(29);
    layer0_outputs(3936) <= (inputs(28)) or (inputs(175));
    layer0_outputs(3937) <= not((inputs(74)) or (inputs(202)));
    layer0_outputs(3938) <= (inputs(161)) xor (inputs(229));
    layer0_outputs(3939) <= not((inputs(140)) or (inputs(139)));
    layer0_outputs(3940) <= not(inputs(200));
    layer0_outputs(3941) <= not(inputs(19));
    layer0_outputs(3942) <= not(inputs(98));
    layer0_outputs(3943) <= inputs(16);
    layer0_outputs(3944) <= not((inputs(60)) and (inputs(177)));
    layer0_outputs(3945) <= not(inputs(186)) or (inputs(37));
    layer0_outputs(3946) <= inputs(183);
    layer0_outputs(3947) <= (inputs(36)) or (inputs(227));
    layer0_outputs(3948) <= not(inputs(54));
    layer0_outputs(3949) <= not(inputs(181)) or (inputs(232));
    layer0_outputs(3950) <= (inputs(210)) xor (inputs(247));
    layer0_outputs(3951) <= (inputs(50)) and not (inputs(85));
    layer0_outputs(3952) <= not(inputs(38));
    layer0_outputs(3953) <= not(inputs(89));
    layer0_outputs(3954) <= not(inputs(137)) or (inputs(98));
    layer0_outputs(3955) <= (inputs(122)) and not (inputs(212));
    layer0_outputs(3956) <= '1';
    layer0_outputs(3957) <= not(inputs(107));
    layer0_outputs(3958) <= inputs(88);
    layer0_outputs(3959) <= not((inputs(159)) xor (inputs(212)));
    layer0_outputs(3960) <= (inputs(67)) xor (inputs(61));
    layer0_outputs(3961) <= (inputs(149)) and not (inputs(14));
    layer0_outputs(3962) <= not(inputs(149)) or (inputs(4));
    layer0_outputs(3963) <= (inputs(82)) or (inputs(4));
    layer0_outputs(3964) <= not((inputs(196)) or (inputs(160)));
    layer0_outputs(3965) <= (inputs(203)) and not (inputs(243));
    layer0_outputs(3966) <= inputs(139);
    layer0_outputs(3967) <= inputs(169);
    layer0_outputs(3968) <= inputs(106);
    layer0_outputs(3969) <= inputs(91);
    layer0_outputs(3970) <= inputs(65);
    layer0_outputs(3971) <= not(inputs(225)) or (inputs(54));
    layer0_outputs(3972) <= (inputs(179)) and not (inputs(43));
    layer0_outputs(3973) <= not((inputs(212)) or (inputs(178)));
    layer0_outputs(3974) <= not((inputs(52)) or (inputs(76)));
    layer0_outputs(3975) <= (inputs(204)) xor (inputs(55));
    layer0_outputs(3976) <= not((inputs(148)) or (inputs(142)));
    layer0_outputs(3977) <= not((inputs(11)) xor (inputs(184)));
    layer0_outputs(3978) <= (inputs(171)) or (inputs(195));
    layer0_outputs(3979) <= not((inputs(5)) xor (inputs(137)));
    layer0_outputs(3980) <= not(inputs(37)) or (inputs(44));
    layer0_outputs(3981) <= not(inputs(248));
    layer0_outputs(3982) <= not(inputs(255)) or (inputs(242));
    layer0_outputs(3983) <= '0';
    layer0_outputs(3984) <= not(inputs(86)) or (inputs(177));
    layer0_outputs(3985) <= (inputs(2)) and not (inputs(57));
    layer0_outputs(3986) <= (inputs(86)) or (inputs(85));
    layer0_outputs(3987) <= not(inputs(108)) or (inputs(210));
    layer0_outputs(3988) <= not((inputs(94)) or (inputs(240)));
    layer0_outputs(3989) <= not((inputs(53)) and (inputs(145)));
    layer0_outputs(3990) <= (inputs(164)) xor (inputs(166));
    layer0_outputs(3991) <= inputs(45);
    layer0_outputs(3992) <= (inputs(48)) and not (inputs(79));
    layer0_outputs(3993) <= (inputs(153)) and (inputs(84));
    layer0_outputs(3994) <= not((inputs(179)) or (inputs(54)));
    layer0_outputs(3995) <= not((inputs(255)) xor (inputs(107)));
    layer0_outputs(3996) <= '0';
    layer0_outputs(3997) <= (inputs(27)) or (inputs(213));
    layer0_outputs(3998) <= not(inputs(188));
    layer0_outputs(3999) <= not((inputs(142)) or (inputs(46)));
    layer0_outputs(4000) <= (inputs(136)) xor (inputs(41));
    layer0_outputs(4001) <= (inputs(82)) xor (inputs(95));
    layer0_outputs(4002) <= (inputs(11)) and not (inputs(97));
    layer0_outputs(4003) <= not(inputs(150));
    layer0_outputs(4004) <= (inputs(150)) and (inputs(95));
    layer0_outputs(4005) <= (inputs(27)) or (inputs(11));
    layer0_outputs(4006) <= not(inputs(190));
    layer0_outputs(4007) <= not(inputs(186)) or (inputs(165));
    layer0_outputs(4008) <= not((inputs(79)) and (inputs(24)));
    layer0_outputs(4009) <= not((inputs(6)) and (inputs(58)));
    layer0_outputs(4010) <= (inputs(48)) or (inputs(135));
    layer0_outputs(4011) <= (inputs(118)) or (inputs(241));
    layer0_outputs(4012) <= not(inputs(130)) or (inputs(19));
    layer0_outputs(4013) <= not((inputs(137)) or (inputs(168)));
    layer0_outputs(4014) <= (inputs(229)) and not (inputs(2));
    layer0_outputs(4015) <= '0';
    layer0_outputs(4016) <= '1';
    layer0_outputs(4017) <= (inputs(75)) and (inputs(200));
    layer0_outputs(4018) <= not((inputs(228)) xor (inputs(195)));
    layer0_outputs(4019) <= (inputs(64)) and not (inputs(204));
    layer0_outputs(4020) <= not((inputs(98)) xor (inputs(105)));
    layer0_outputs(4021) <= inputs(249);
    layer0_outputs(4022) <= not((inputs(192)) and (inputs(255)));
    layer0_outputs(4023) <= (inputs(73)) and not (inputs(181));
    layer0_outputs(4024) <= not((inputs(58)) and (inputs(51)));
    layer0_outputs(4025) <= (inputs(205)) and not (inputs(255));
    layer0_outputs(4026) <= not(inputs(19)) or (inputs(188));
    layer0_outputs(4027) <= (inputs(62)) and not (inputs(233));
    layer0_outputs(4028) <= (inputs(75)) xor (inputs(212));
    layer0_outputs(4029) <= inputs(197);
    layer0_outputs(4030) <= '1';
    layer0_outputs(4031) <= inputs(135);
    layer0_outputs(4032) <= not((inputs(192)) xor (inputs(149)));
    layer0_outputs(4033) <= (inputs(163)) and not (inputs(28));
    layer0_outputs(4034) <= not((inputs(14)) xor (inputs(88)));
    layer0_outputs(4035) <= not((inputs(8)) or (inputs(22)));
    layer0_outputs(4036) <= not((inputs(211)) or (inputs(166)));
    layer0_outputs(4037) <= not((inputs(168)) xor (inputs(62)));
    layer0_outputs(4038) <= inputs(79);
    layer0_outputs(4039) <= (inputs(74)) and (inputs(214));
    layer0_outputs(4040) <= (inputs(37)) and not (inputs(234));
    layer0_outputs(4041) <= (inputs(250)) and (inputs(70));
    layer0_outputs(4042) <= (inputs(103)) and not (inputs(242));
    layer0_outputs(4043) <= (inputs(138)) or (inputs(62));
    layer0_outputs(4044) <= (inputs(78)) or (inputs(222));
    layer0_outputs(4045) <= inputs(94);
    layer0_outputs(4046) <= (inputs(63)) and not (inputs(1));
    layer0_outputs(4047) <= not(inputs(55));
    layer0_outputs(4048) <= '0';
    layer0_outputs(4049) <= '0';
    layer0_outputs(4050) <= not((inputs(72)) xor (inputs(56)));
    layer0_outputs(4051) <= not((inputs(69)) xor (inputs(0)));
    layer0_outputs(4052) <= not((inputs(6)) and (inputs(79)));
    layer0_outputs(4053) <= not(inputs(181));
    layer0_outputs(4054) <= '0';
    layer0_outputs(4055) <= not(inputs(245));
    layer0_outputs(4056) <= not((inputs(219)) or (inputs(5)));
    layer0_outputs(4057) <= (inputs(192)) or (inputs(231));
    layer0_outputs(4058) <= not(inputs(151)) or (inputs(223));
    layer0_outputs(4059) <= not(inputs(16)) or (inputs(0));
    layer0_outputs(4060) <= inputs(214);
    layer0_outputs(4061) <= '1';
    layer0_outputs(4062) <= not(inputs(223)) or (inputs(52));
    layer0_outputs(4063) <= not(inputs(237));
    layer0_outputs(4064) <= (inputs(4)) or (inputs(20));
    layer0_outputs(4065) <= (inputs(34)) and not (inputs(224));
    layer0_outputs(4066) <= not((inputs(116)) and (inputs(116)));
    layer0_outputs(4067) <= '1';
    layer0_outputs(4068) <= '0';
    layer0_outputs(4069) <= not((inputs(112)) xor (inputs(29)));
    layer0_outputs(4070) <= (inputs(252)) and not (inputs(217));
    layer0_outputs(4071) <= inputs(137);
    layer0_outputs(4072) <= (inputs(36)) xor (inputs(120));
    layer0_outputs(4073) <= '0';
    layer0_outputs(4074) <= not((inputs(131)) or (inputs(171)));
    layer0_outputs(4075) <= '0';
    layer0_outputs(4076) <= not((inputs(188)) or (inputs(194)));
    layer0_outputs(4077) <= (inputs(234)) and not (inputs(232));
    layer0_outputs(4078) <= '1';
    layer0_outputs(4079) <= (inputs(22)) and (inputs(26));
    layer0_outputs(4080) <= (inputs(181)) xor (inputs(14));
    layer0_outputs(4081) <= (inputs(76)) or (inputs(187));
    layer0_outputs(4082) <= not(inputs(239));
    layer0_outputs(4083) <= (inputs(42)) xor (inputs(44));
    layer0_outputs(4084) <= (inputs(46)) and not (inputs(17));
    layer0_outputs(4085) <= not((inputs(147)) and (inputs(249)));
    layer0_outputs(4086) <= inputs(225);
    layer0_outputs(4087) <= not(inputs(28));
    layer0_outputs(4088) <= not(inputs(241));
    layer0_outputs(4089) <= '0';
    layer0_outputs(4090) <= not((inputs(43)) and (inputs(246)));
    layer0_outputs(4091) <= not(inputs(41)) or (inputs(229));
    layer0_outputs(4092) <= not(inputs(200));
    layer0_outputs(4093) <= '0';
    layer0_outputs(4094) <= not(inputs(120));
    layer0_outputs(4095) <= not((inputs(194)) and (inputs(34)));
    layer0_outputs(4096) <= not((inputs(88)) xor (inputs(120)));
    layer0_outputs(4097) <= '1';
    layer0_outputs(4098) <= (inputs(159)) xor (inputs(218));
    layer0_outputs(4099) <= not(inputs(104)) or (inputs(47));
    layer0_outputs(4100) <= not(inputs(20));
    layer0_outputs(4101) <= not(inputs(137));
    layer0_outputs(4102) <= (inputs(214)) xor (inputs(96));
    layer0_outputs(4103) <= not(inputs(191));
    layer0_outputs(4104) <= not(inputs(184)) or (inputs(48));
    layer0_outputs(4105) <= (inputs(52)) and not (inputs(11));
    layer0_outputs(4106) <= not(inputs(212));
    layer0_outputs(4107) <= not(inputs(94)) or (inputs(87));
    layer0_outputs(4108) <= (inputs(235)) and not (inputs(192));
    layer0_outputs(4109) <= (inputs(74)) and not (inputs(175));
    layer0_outputs(4110) <= (inputs(116)) and not (inputs(103));
    layer0_outputs(4111) <= not((inputs(249)) and (inputs(66)));
    layer0_outputs(4112) <= not(inputs(120));
    layer0_outputs(4113) <= not((inputs(83)) or (inputs(70)));
    layer0_outputs(4114) <= not(inputs(187)) or (inputs(234));
    layer0_outputs(4115) <= (inputs(220)) and (inputs(212));
    layer0_outputs(4116) <= (inputs(232)) xor (inputs(34));
    layer0_outputs(4117) <= not((inputs(84)) or (inputs(20)));
    layer0_outputs(4118) <= not(inputs(42));
    layer0_outputs(4119) <= not((inputs(113)) xor (inputs(83)));
    layer0_outputs(4120) <= (inputs(73)) xor (inputs(254));
    layer0_outputs(4121) <= inputs(178);
    layer0_outputs(4122) <= '0';
    layer0_outputs(4123) <= not((inputs(216)) and (inputs(254)));
    layer0_outputs(4124) <= (inputs(149)) and not (inputs(24));
    layer0_outputs(4125) <= (inputs(33)) or (inputs(9));
    layer0_outputs(4126) <= not(inputs(140));
    layer0_outputs(4127) <= (inputs(246)) and (inputs(159));
    layer0_outputs(4128) <= not((inputs(49)) xor (inputs(199)));
    layer0_outputs(4129) <= (inputs(11)) or (inputs(118));
    layer0_outputs(4130) <= not((inputs(171)) or (inputs(224)));
    layer0_outputs(4131) <= '0';
    layer0_outputs(4132) <= not(inputs(220));
    layer0_outputs(4133) <= inputs(187);
    layer0_outputs(4134) <= (inputs(144)) and not (inputs(123));
    layer0_outputs(4135) <= inputs(137);
    layer0_outputs(4136) <= not(inputs(176)) or (inputs(32));
    layer0_outputs(4137) <= not(inputs(191)) or (inputs(247));
    layer0_outputs(4138) <= not((inputs(188)) or (inputs(56)));
    layer0_outputs(4139) <= not((inputs(139)) and (inputs(143)));
    layer0_outputs(4140) <= not((inputs(4)) and (inputs(70)));
    layer0_outputs(4141) <= not(inputs(124)) or (inputs(145));
    layer0_outputs(4142) <= not(inputs(224));
    layer0_outputs(4143) <= inputs(198);
    layer0_outputs(4144) <= not(inputs(104));
    layer0_outputs(4145) <= (inputs(233)) and not (inputs(42));
    layer0_outputs(4146) <= not(inputs(110)) or (inputs(41));
    layer0_outputs(4147) <= not(inputs(212));
    layer0_outputs(4148) <= (inputs(186)) and not (inputs(238));
    layer0_outputs(4149) <= not((inputs(209)) or (inputs(34)));
    layer0_outputs(4150) <= '1';
    layer0_outputs(4151) <= not(inputs(134));
    layer0_outputs(4152) <= (inputs(124)) and not (inputs(204));
    layer0_outputs(4153) <= (inputs(92)) xor (inputs(37));
    layer0_outputs(4154) <= (inputs(98)) or (inputs(86));
    layer0_outputs(4155) <= (inputs(219)) or (inputs(136));
    layer0_outputs(4156) <= not((inputs(206)) xor (inputs(22)));
    layer0_outputs(4157) <= (inputs(0)) and not (inputs(191));
    layer0_outputs(4158) <= '0';
    layer0_outputs(4159) <= inputs(98);
    layer0_outputs(4160) <= not(inputs(175));
    layer0_outputs(4161) <= not((inputs(51)) or (inputs(40)));
    layer0_outputs(4162) <= not((inputs(248)) or (inputs(129)));
    layer0_outputs(4163) <= not((inputs(214)) or (inputs(99)));
    layer0_outputs(4164) <= '1';
    layer0_outputs(4165) <= not(inputs(123));
    layer0_outputs(4166) <= not(inputs(4));
    layer0_outputs(4167) <= not((inputs(177)) xor (inputs(32)));
    layer0_outputs(4168) <= (inputs(177)) and (inputs(119));
    layer0_outputs(4169) <= (inputs(70)) and (inputs(255));
    layer0_outputs(4170) <= not(inputs(87));
    layer0_outputs(4171) <= not((inputs(118)) xor (inputs(96)));
    layer0_outputs(4172) <= (inputs(162)) or (inputs(27));
    layer0_outputs(4173) <= not(inputs(46)) or (inputs(29));
    layer0_outputs(4174) <= not(inputs(157));
    layer0_outputs(4175) <= not(inputs(235)) or (inputs(217));
    layer0_outputs(4176) <= not(inputs(160)) or (inputs(107));
    layer0_outputs(4177) <= '0';
    layer0_outputs(4178) <= not(inputs(142)) or (inputs(114));
    layer0_outputs(4179) <= (inputs(231)) and not (inputs(93));
    layer0_outputs(4180) <= (inputs(112)) and not (inputs(29));
    layer0_outputs(4181) <= (inputs(227)) and not (inputs(202));
    layer0_outputs(4182) <= inputs(174);
    layer0_outputs(4183) <= inputs(167);
    layer0_outputs(4184) <= (inputs(138)) or (inputs(254));
    layer0_outputs(4185) <= '1';
    layer0_outputs(4186) <= not((inputs(67)) and (inputs(12)));
    layer0_outputs(4187) <= (inputs(209)) and (inputs(132));
    layer0_outputs(4188) <= '1';
    layer0_outputs(4189) <= '0';
    layer0_outputs(4190) <= not(inputs(121)) or (inputs(33));
    layer0_outputs(4191) <= not(inputs(71)) or (inputs(178));
    layer0_outputs(4192) <= (inputs(170)) or (inputs(165));
    layer0_outputs(4193) <= not((inputs(247)) xor (inputs(233)));
    layer0_outputs(4194) <= (inputs(154)) and not (inputs(251));
    layer0_outputs(4195) <= '0';
    layer0_outputs(4196) <= (inputs(244)) and not (inputs(36));
    layer0_outputs(4197) <= (inputs(169)) and (inputs(100));
    layer0_outputs(4198) <= not(inputs(166)) or (inputs(237));
    layer0_outputs(4199) <= not(inputs(205)) or (inputs(250));
    layer0_outputs(4200) <= inputs(127);
    layer0_outputs(4201) <= (inputs(215)) or (inputs(204));
    layer0_outputs(4202) <= (inputs(116)) or (inputs(239));
    layer0_outputs(4203) <= '1';
    layer0_outputs(4204) <= (inputs(212)) xor (inputs(177));
    layer0_outputs(4205) <= not((inputs(157)) xor (inputs(245)));
    layer0_outputs(4206) <= (inputs(115)) xor (inputs(2));
    layer0_outputs(4207) <= not((inputs(0)) and (inputs(184)));
    layer0_outputs(4208) <= '1';
    layer0_outputs(4209) <= not((inputs(124)) or (inputs(250)));
    layer0_outputs(4210) <= '0';
    layer0_outputs(4211) <= not((inputs(100)) or (inputs(104)));
    layer0_outputs(4212) <= (inputs(94)) or (inputs(48));
    layer0_outputs(4213) <= not((inputs(160)) and (inputs(201)));
    layer0_outputs(4214) <= not(inputs(148));
    layer0_outputs(4215) <= not(inputs(131)) or (inputs(235));
    layer0_outputs(4216) <= (inputs(70)) or (inputs(240));
    layer0_outputs(4217) <= inputs(140);
    layer0_outputs(4218) <= not(inputs(11));
    layer0_outputs(4219) <= not((inputs(30)) xor (inputs(205)));
    layer0_outputs(4220) <= (inputs(21)) and not (inputs(225));
    layer0_outputs(4221) <= (inputs(9)) and not (inputs(198));
    layer0_outputs(4222) <= not((inputs(253)) or (inputs(193)));
    layer0_outputs(4223) <= not((inputs(1)) and (inputs(213)));
    layer0_outputs(4224) <= not(inputs(116));
    layer0_outputs(4225) <= (inputs(25)) or (inputs(236));
    layer0_outputs(4226) <= inputs(27);
    layer0_outputs(4227) <= not(inputs(134)) or (inputs(35));
    layer0_outputs(4228) <= inputs(119);
    layer0_outputs(4229) <= not(inputs(37));
    layer0_outputs(4230) <= not((inputs(81)) xor (inputs(199)));
    layer0_outputs(4231) <= (inputs(48)) or (inputs(244));
    layer0_outputs(4232) <= (inputs(44)) xor (inputs(118));
    layer0_outputs(4233) <= not((inputs(213)) or (inputs(105)));
    layer0_outputs(4234) <= not((inputs(115)) xor (inputs(143)));
    layer0_outputs(4235) <= not(inputs(131)) or (inputs(27));
    layer0_outputs(4236) <= (inputs(137)) or (inputs(166));
    layer0_outputs(4237) <= (inputs(34)) xor (inputs(29));
    layer0_outputs(4238) <= not(inputs(166)) or (inputs(233));
    layer0_outputs(4239) <= (inputs(173)) or (inputs(81));
    layer0_outputs(4240) <= (inputs(106)) and not (inputs(236));
    layer0_outputs(4241) <= not((inputs(49)) and (inputs(130)));
    layer0_outputs(4242) <= not(inputs(90));
    layer0_outputs(4243) <= (inputs(218)) or (inputs(200));
    layer0_outputs(4244) <= not(inputs(74)) or (inputs(36));
    layer0_outputs(4245) <= not((inputs(221)) and (inputs(212)));
    layer0_outputs(4246) <= (inputs(22)) and not (inputs(211));
    layer0_outputs(4247) <= not((inputs(200)) or (inputs(177)));
    layer0_outputs(4248) <= not((inputs(103)) and (inputs(199)));
    layer0_outputs(4249) <= (inputs(121)) and (inputs(241));
    layer0_outputs(4250) <= (inputs(204)) and not (inputs(226));
    layer0_outputs(4251) <= not((inputs(115)) xor (inputs(65)));
    layer0_outputs(4252) <= not(inputs(125));
    layer0_outputs(4253) <= inputs(247);
    layer0_outputs(4254) <= (inputs(117)) xor (inputs(161));
    layer0_outputs(4255) <= (inputs(186)) or (inputs(169));
    layer0_outputs(4256) <= not((inputs(228)) or (inputs(198)));
    layer0_outputs(4257) <= (inputs(42)) and not (inputs(189));
    layer0_outputs(4258) <= not(inputs(220)) or (inputs(103));
    layer0_outputs(4259) <= not(inputs(123)) or (inputs(53));
    layer0_outputs(4260) <= not(inputs(64));
    layer0_outputs(4261) <= (inputs(225)) and (inputs(92));
    layer0_outputs(4262) <= (inputs(175)) and not (inputs(94));
    layer0_outputs(4263) <= '0';
    layer0_outputs(4264) <= (inputs(6)) xor (inputs(54));
    layer0_outputs(4265) <= not(inputs(193)) or (inputs(145));
    layer0_outputs(4266) <= (inputs(79)) and not (inputs(6));
    layer0_outputs(4267) <= (inputs(6)) and not (inputs(13));
    layer0_outputs(4268) <= (inputs(113)) or (inputs(216));
    layer0_outputs(4269) <= not(inputs(150));
    layer0_outputs(4270) <= not(inputs(100));
    layer0_outputs(4271) <= not((inputs(128)) xor (inputs(27)));
    layer0_outputs(4272) <= (inputs(25)) xor (inputs(43));
    layer0_outputs(4273) <= not((inputs(132)) or (inputs(97)));
    layer0_outputs(4274) <= (inputs(58)) xor (inputs(157));
    layer0_outputs(4275) <= not(inputs(167));
    layer0_outputs(4276) <= (inputs(40)) or (inputs(178));
    layer0_outputs(4277) <= inputs(199);
    layer0_outputs(4278) <= not(inputs(56)) or (inputs(210));
    layer0_outputs(4279) <= not((inputs(67)) and (inputs(145)));
    layer0_outputs(4280) <= (inputs(162)) and (inputs(212));
    layer0_outputs(4281) <= not(inputs(112)) or (inputs(107));
    layer0_outputs(4282) <= not((inputs(3)) and (inputs(61)));
    layer0_outputs(4283) <= not((inputs(114)) or (inputs(88)));
    layer0_outputs(4284) <= '1';
    layer0_outputs(4285) <= not((inputs(119)) or (inputs(39)));
    layer0_outputs(4286) <= '1';
    layer0_outputs(4287) <= not((inputs(168)) and (inputs(52)));
    layer0_outputs(4288) <= not(inputs(213));
    layer0_outputs(4289) <= not((inputs(110)) xor (inputs(120)));
    layer0_outputs(4290) <= not((inputs(233)) xor (inputs(25)));
    layer0_outputs(4291) <= (inputs(200)) or (inputs(255));
    layer0_outputs(4292) <= inputs(166);
    layer0_outputs(4293) <= (inputs(108)) or (inputs(171));
    layer0_outputs(4294) <= inputs(77);
    layer0_outputs(4295) <= not((inputs(215)) xor (inputs(192)));
    layer0_outputs(4296) <= (inputs(90)) xor (inputs(239));
    layer0_outputs(4297) <= '1';
    layer0_outputs(4298) <= '1';
    layer0_outputs(4299) <= not(inputs(137)) or (inputs(174));
    layer0_outputs(4300) <= inputs(221);
    layer0_outputs(4301) <= inputs(203);
    layer0_outputs(4302) <= '1';
    layer0_outputs(4303) <= not(inputs(253)) or (inputs(49));
    layer0_outputs(4304) <= (inputs(167)) or (inputs(53));
    layer0_outputs(4305) <= not(inputs(75));
    layer0_outputs(4306) <= (inputs(36)) xor (inputs(9));
    layer0_outputs(4307) <= inputs(169);
    layer0_outputs(4308) <= not(inputs(163)) or (inputs(1));
    layer0_outputs(4309) <= (inputs(104)) or (inputs(213));
    layer0_outputs(4310) <= not((inputs(231)) or (inputs(235)));
    layer0_outputs(4311) <= (inputs(157)) or (inputs(126));
    layer0_outputs(4312) <= inputs(167);
    layer0_outputs(4313) <= not(inputs(139)) or (inputs(76));
    layer0_outputs(4314) <= not((inputs(173)) or (inputs(100)));
    layer0_outputs(4315) <= (inputs(46)) and not (inputs(51));
    layer0_outputs(4316) <= inputs(165);
    layer0_outputs(4317) <= (inputs(76)) xor (inputs(45));
    layer0_outputs(4318) <= not((inputs(149)) or (inputs(44)));
    layer0_outputs(4319) <= not(inputs(134)) or (inputs(30));
    layer0_outputs(4320) <= not((inputs(208)) or (inputs(124)));
    layer0_outputs(4321) <= not(inputs(249));
    layer0_outputs(4322) <= not(inputs(246)) or (inputs(35));
    layer0_outputs(4323) <= inputs(84);
    layer0_outputs(4324) <= '1';
    layer0_outputs(4325) <= not(inputs(165));
    layer0_outputs(4326) <= not(inputs(24)) or (inputs(213));
    layer0_outputs(4327) <= not(inputs(76));
    layer0_outputs(4328) <= not((inputs(51)) xor (inputs(19)));
    layer0_outputs(4329) <= not((inputs(129)) xor (inputs(87)));
    layer0_outputs(4330) <= (inputs(134)) and (inputs(159));
    layer0_outputs(4331) <= (inputs(14)) and (inputs(150));
    layer0_outputs(4332) <= not(inputs(25));
    layer0_outputs(4333) <= (inputs(10)) xor (inputs(199));
    layer0_outputs(4334) <= not((inputs(188)) or (inputs(58)));
    layer0_outputs(4335) <= (inputs(130)) xor (inputs(102));
    layer0_outputs(4336) <= not((inputs(132)) or (inputs(223)));
    layer0_outputs(4337) <= not((inputs(13)) or (inputs(17)));
    layer0_outputs(4338) <= inputs(25);
    layer0_outputs(4339) <= not((inputs(187)) or (inputs(139)));
    layer0_outputs(4340) <= not(inputs(104));
    layer0_outputs(4341) <= (inputs(31)) xor (inputs(37));
    layer0_outputs(4342) <= (inputs(66)) xor (inputs(63));
    layer0_outputs(4343) <= '1';
    layer0_outputs(4344) <= not((inputs(36)) and (inputs(3)));
    layer0_outputs(4345) <= not((inputs(183)) or (inputs(94)));
    layer0_outputs(4346) <= not(inputs(145)) or (inputs(178));
    layer0_outputs(4347) <= not(inputs(127)) or (inputs(171));
    layer0_outputs(4348) <= '0';
    layer0_outputs(4349) <= not(inputs(112)) or (inputs(80));
    layer0_outputs(4350) <= not(inputs(109)) or (inputs(162));
    layer0_outputs(4351) <= (inputs(133)) and not (inputs(34));
    layer0_outputs(4352) <= '0';
    layer0_outputs(4353) <= '0';
    layer0_outputs(4354) <= not(inputs(115));
    layer0_outputs(4355) <= not(inputs(148));
    layer0_outputs(4356) <= (inputs(193)) or (inputs(198));
    layer0_outputs(4357) <= (inputs(207)) and not (inputs(254));
    layer0_outputs(4358) <= not((inputs(220)) xor (inputs(43)));
    layer0_outputs(4359) <= (inputs(102)) and not (inputs(21));
    layer0_outputs(4360) <= not((inputs(17)) and (inputs(187)));
    layer0_outputs(4361) <= (inputs(52)) and not (inputs(6));
    layer0_outputs(4362) <= (inputs(228)) or (inputs(86));
    layer0_outputs(4363) <= (inputs(122)) and not (inputs(81));
    layer0_outputs(4364) <= inputs(169);
    layer0_outputs(4365) <= not((inputs(221)) and (inputs(111)));
    layer0_outputs(4366) <= inputs(218);
    layer0_outputs(4367) <= (inputs(73)) xor (inputs(93));
    layer0_outputs(4368) <= (inputs(87)) and not (inputs(39));
    layer0_outputs(4369) <= not((inputs(240)) or (inputs(213)));
    layer0_outputs(4370) <= not(inputs(194));
    layer0_outputs(4371) <= not((inputs(212)) and (inputs(30)));
    layer0_outputs(4372) <= '1';
    layer0_outputs(4373) <= (inputs(29)) and (inputs(37));
    layer0_outputs(4374) <= (inputs(69)) and (inputs(153));
    layer0_outputs(4375) <= '0';
    layer0_outputs(4376) <= (inputs(149)) or (inputs(129));
    layer0_outputs(4377) <= not(inputs(208));
    layer0_outputs(4378) <= not((inputs(61)) and (inputs(206)));
    layer0_outputs(4379) <= (inputs(82)) or (inputs(234));
    layer0_outputs(4380) <= (inputs(115)) xor (inputs(241));
    layer0_outputs(4381) <= (inputs(249)) and not (inputs(26));
    layer0_outputs(4382) <= not((inputs(54)) or (inputs(157)));
    layer0_outputs(4383) <= (inputs(68)) xor (inputs(122));
    layer0_outputs(4384) <= not((inputs(194)) or (inputs(204)));
    layer0_outputs(4385) <= not((inputs(127)) xor (inputs(119)));
    layer0_outputs(4386) <= not((inputs(174)) and (inputs(63)));
    layer0_outputs(4387) <= not((inputs(113)) or (inputs(84)));
    layer0_outputs(4388) <= not((inputs(250)) or (inputs(248)));
    layer0_outputs(4389) <= '1';
    layer0_outputs(4390) <= (inputs(89)) or (inputs(233));
    layer0_outputs(4391) <= (inputs(188)) and not (inputs(127));
    layer0_outputs(4392) <= '1';
    layer0_outputs(4393) <= not(inputs(142));
    layer0_outputs(4394) <= not(inputs(50)) or (inputs(1));
    layer0_outputs(4395) <= (inputs(142)) xor (inputs(250));
    layer0_outputs(4396) <= (inputs(248)) or (inputs(89));
    layer0_outputs(4397) <= not(inputs(1));
    layer0_outputs(4398) <= not((inputs(96)) or (inputs(59)));
    layer0_outputs(4399) <= (inputs(253)) and not (inputs(213));
    layer0_outputs(4400) <= not((inputs(73)) or (inputs(220)));
    layer0_outputs(4401) <= not(inputs(74));
    layer0_outputs(4402) <= inputs(64);
    layer0_outputs(4403) <= not(inputs(106));
    layer0_outputs(4404) <= not(inputs(151));
    layer0_outputs(4405) <= (inputs(108)) or (inputs(14));
    layer0_outputs(4406) <= not(inputs(88));
    layer0_outputs(4407) <= not((inputs(208)) or (inputs(10)));
    layer0_outputs(4408) <= inputs(124);
    layer0_outputs(4409) <= (inputs(85)) and not (inputs(177));
    layer0_outputs(4410) <= (inputs(156)) or (inputs(169));
    layer0_outputs(4411) <= (inputs(113)) and not (inputs(148));
    layer0_outputs(4412) <= not((inputs(55)) xor (inputs(133)));
    layer0_outputs(4413) <= not(inputs(170));
    layer0_outputs(4414) <= not(inputs(76)) or (inputs(193));
    layer0_outputs(4415) <= (inputs(218)) xor (inputs(147));
    layer0_outputs(4416) <= '1';
    layer0_outputs(4417) <= not(inputs(119)) or (inputs(9));
    layer0_outputs(4418) <= (inputs(201)) and not (inputs(95));
    layer0_outputs(4419) <= (inputs(82)) or (inputs(231));
    layer0_outputs(4420) <= (inputs(59)) and not (inputs(3));
    layer0_outputs(4421) <= '0';
    layer0_outputs(4422) <= not(inputs(216)) or (inputs(249));
    layer0_outputs(4423) <= not((inputs(213)) xor (inputs(206)));
    layer0_outputs(4424) <= not(inputs(40));
    layer0_outputs(4425) <= (inputs(164)) and not (inputs(124));
    layer0_outputs(4426) <= (inputs(167)) xor (inputs(33));
    layer0_outputs(4427) <= inputs(186);
    layer0_outputs(4428) <= inputs(83);
    layer0_outputs(4429) <= not((inputs(81)) or (inputs(147)));
    layer0_outputs(4430) <= (inputs(106)) and not (inputs(201));
    layer0_outputs(4431) <= inputs(213);
    layer0_outputs(4432) <= not(inputs(123));
    layer0_outputs(4433) <= not(inputs(179)) or (inputs(241));
    layer0_outputs(4434) <= '1';
    layer0_outputs(4435) <= inputs(138);
    layer0_outputs(4436) <= (inputs(45)) or (inputs(11));
    layer0_outputs(4437) <= (inputs(89)) and (inputs(187));
    layer0_outputs(4438) <= not((inputs(239)) or (inputs(182)));
    layer0_outputs(4439) <= '0';
    layer0_outputs(4440) <= '0';
    layer0_outputs(4441) <= (inputs(62)) and not (inputs(13));
    layer0_outputs(4442) <= not(inputs(116));
    layer0_outputs(4443) <= not((inputs(70)) xor (inputs(87)));
    layer0_outputs(4444) <= not((inputs(220)) and (inputs(146)));
    layer0_outputs(4445) <= not((inputs(161)) or (inputs(176)));
    layer0_outputs(4446) <= (inputs(190)) or (inputs(198));
    layer0_outputs(4447) <= inputs(5);
    layer0_outputs(4448) <= not((inputs(69)) and (inputs(9)));
    layer0_outputs(4449) <= inputs(248);
    layer0_outputs(4450) <= (inputs(88)) or (inputs(234));
    layer0_outputs(4451) <= not(inputs(51)) or (inputs(1));
    layer0_outputs(4452) <= inputs(136);
    layer0_outputs(4453) <= (inputs(193)) and not (inputs(14));
    layer0_outputs(4454) <= not((inputs(157)) or (inputs(148)));
    layer0_outputs(4455) <= inputs(167);
    layer0_outputs(4456) <= (inputs(49)) and not (inputs(2));
    layer0_outputs(4457) <= inputs(3);
    layer0_outputs(4458) <= not(inputs(113));
    layer0_outputs(4459) <= not((inputs(14)) xor (inputs(115)));
    layer0_outputs(4460) <= inputs(42);
    layer0_outputs(4461) <= not(inputs(173));
    layer0_outputs(4462) <= not(inputs(46)) or (inputs(79));
    layer0_outputs(4463) <= (inputs(57)) xor (inputs(204));
    layer0_outputs(4464) <= (inputs(247)) or (inputs(71));
    layer0_outputs(4465) <= inputs(119);
    layer0_outputs(4466) <= (inputs(157)) xor (inputs(37));
    layer0_outputs(4467) <= not(inputs(114));
    layer0_outputs(4468) <= inputs(89);
    layer0_outputs(4469) <= not((inputs(5)) and (inputs(177)));
    layer0_outputs(4470) <= (inputs(109)) xor (inputs(242));
    layer0_outputs(4471) <= (inputs(31)) or (inputs(219));
    layer0_outputs(4472) <= (inputs(14)) or (inputs(172));
    layer0_outputs(4473) <= (inputs(206)) xor (inputs(30));
    layer0_outputs(4474) <= '0';
    layer0_outputs(4475) <= (inputs(121)) or (inputs(86));
    layer0_outputs(4476) <= not((inputs(96)) xor (inputs(81)));
    layer0_outputs(4477) <= not((inputs(62)) and (inputs(3)));
    layer0_outputs(4478) <= not((inputs(18)) or (inputs(254)));
    layer0_outputs(4479) <= inputs(58);
    layer0_outputs(4480) <= not(inputs(116));
    layer0_outputs(4481) <= (inputs(46)) or (inputs(117));
    layer0_outputs(4482) <= not(inputs(57)) or (inputs(141));
    layer0_outputs(4483) <= '0';
    layer0_outputs(4484) <= not((inputs(193)) xor (inputs(196)));
    layer0_outputs(4485) <= inputs(1);
    layer0_outputs(4486) <= (inputs(251)) and not (inputs(20));
    layer0_outputs(4487) <= inputs(180);
    layer0_outputs(4488) <= not(inputs(133));
    layer0_outputs(4489) <= (inputs(223)) and not (inputs(0));
    layer0_outputs(4490) <= '0';
    layer0_outputs(4491) <= not(inputs(143));
    layer0_outputs(4492) <= not((inputs(67)) xor (inputs(142)));
    layer0_outputs(4493) <= (inputs(223)) or (inputs(197));
    layer0_outputs(4494) <= not(inputs(128));
    layer0_outputs(4495) <= (inputs(5)) and not (inputs(158));
    layer0_outputs(4496) <= inputs(153);
    layer0_outputs(4497) <= not((inputs(100)) or (inputs(248)));
    layer0_outputs(4498) <= not((inputs(109)) or (inputs(255)));
    layer0_outputs(4499) <= not(inputs(190));
    layer0_outputs(4500) <= not(inputs(3));
    layer0_outputs(4501) <= inputs(118);
    layer0_outputs(4502) <= '1';
    layer0_outputs(4503) <= inputs(229);
    layer0_outputs(4504) <= '0';
    layer0_outputs(4505) <= '0';
    layer0_outputs(4506) <= not(inputs(241));
    layer0_outputs(4507) <= not((inputs(9)) or (inputs(228)));
    layer0_outputs(4508) <= (inputs(131)) or (inputs(124));
    layer0_outputs(4509) <= not(inputs(38));
    layer0_outputs(4510) <= not((inputs(254)) and (inputs(210)));
    layer0_outputs(4511) <= not(inputs(158));
    layer0_outputs(4512) <= inputs(102);
    layer0_outputs(4513) <= not(inputs(228));
    layer0_outputs(4514) <= not((inputs(233)) or (inputs(190)));
    layer0_outputs(4515) <= (inputs(48)) or (inputs(152));
    layer0_outputs(4516) <= (inputs(134)) and not (inputs(93));
    layer0_outputs(4517) <= '1';
    layer0_outputs(4518) <= not(inputs(153)) or (inputs(208));
    layer0_outputs(4519) <= not((inputs(111)) or (inputs(218)));
    layer0_outputs(4520) <= not((inputs(8)) xor (inputs(193)));
    layer0_outputs(4521) <= not(inputs(198));
    layer0_outputs(4522) <= (inputs(244)) and not (inputs(71));
    layer0_outputs(4523) <= (inputs(118)) xor (inputs(172));
    layer0_outputs(4524) <= not((inputs(104)) or (inputs(83)));
    layer0_outputs(4525) <= not(inputs(57));
    layer0_outputs(4526) <= not((inputs(98)) and (inputs(126)));
    layer0_outputs(4527) <= '0';
    layer0_outputs(4528) <= inputs(34);
    layer0_outputs(4529) <= '0';
    layer0_outputs(4530) <= not(inputs(152));
    layer0_outputs(4531) <= (inputs(95)) and not (inputs(16));
    layer0_outputs(4532) <= not(inputs(151)) or (inputs(144));
    layer0_outputs(4533) <= not((inputs(44)) and (inputs(25)));
    layer0_outputs(4534) <= not(inputs(97));
    layer0_outputs(4535) <= not((inputs(247)) or (inputs(55)));
    layer0_outputs(4536) <= not(inputs(215)) or (inputs(67));
    layer0_outputs(4537) <= '0';
    layer0_outputs(4538) <= (inputs(156)) or (inputs(154));
    layer0_outputs(4539) <= (inputs(40)) xor (inputs(55));
    layer0_outputs(4540) <= not((inputs(163)) or (inputs(148)));
    layer0_outputs(4541) <= (inputs(254)) or (inputs(76));
    layer0_outputs(4542) <= (inputs(124)) and not (inputs(72));
    layer0_outputs(4543) <= not((inputs(182)) or (inputs(21)));
    layer0_outputs(4544) <= (inputs(106)) or (inputs(116));
    layer0_outputs(4545) <= '1';
    layer0_outputs(4546) <= (inputs(236)) and not (inputs(118));
    layer0_outputs(4547) <= not((inputs(161)) or (inputs(137)));
    layer0_outputs(4548) <= not(inputs(92));
    layer0_outputs(4549) <= not((inputs(10)) or (inputs(89)));
    layer0_outputs(4550) <= inputs(94);
    layer0_outputs(4551) <= (inputs(12)) and (inputs(99));
    layer0_outputs(4552) <= '1';
    layer0_outputs(4553) <= not(inputs(24));
    layer0_outputs(4554) <= inputs(231);
    layer0_outputs(4555) <= (inputs(42)) and not (inputs(99));
    layer0_outputs(4556) <= not(inputs(50)) or (inputs(32));
    layer0_outputs(4557) <= (inputs(16)) and not (inputs(161));
    layer0_outputs(4558) <= (inputs(159)) xor (inputs(92));
    layer0_outputs(4559) <= not(inputs(9));
    layer0_outputs(4560) <= (inputs(120)) or (inputs(51));
    layer0_outputs(4561) <= inputs(179);
    layer0_outputs(4562) <= not(inputs(150));
    layer0_outputs(4563) <= not(inputs(58));
    layer0_outputs(4564) <= (inputs(15)) and not (inputs(228));
    layer0_outputs(4565) <= inputs(77);
    layer0_outputs(4566) <= (inputs(102)) and not (inputs(142));
    layer0_outputs(4567) <= inputs(66);
    layer0_outputs(4568) <= not((inputs(155)) and (inputs(242)));
    layer0_outputs(4569) <= (inputs(107)) or (inputs(235));
    layer0_outputs(4570) <= (inputs(202)) or (inputs(159));
    layer0_outputs(4571) <= (inputs(90)) and (inputs(171));
    layer0_outputs(4572) <= '0';
    layer0_outputs(4573) <= (inputs(212)) xor (inputs(181));
    layer0_outputs(4574) <= (inputs(37)) and not (inputs(4));
    layer0_outputs(4575) <= (inputs(92)) xor (inputs(108));
    layer0_outputs(4576) <= (inputs(203)) or (inputs(209));
    layer0_outputs(4577) <= (inputs(121)) xor (inputs(63));
    layer0_outputs(4578) <= not(inputs(92)) or (inputs(17));
    layer0_outputs(4579) <= (inputs(39)) and not (inputs(1));
    layer0_outputs(4580) <= not(inputs(148));
    layer0_outputs(4581) <= (inputs(111)) xor (inputs(207));
    layer0_outputs(4582) <= '0';
    layer0_outputs(4583) <= not(inputs(115));
    layer0_outputs(4584) <= inputs(224);
    layer0_outputs(4585) <= not((inputs(158)) and (inputs(197)));
    layer0_outputs(4586) <= '1';
    layer0_outputs(4587) <= (inputs(30)) or (inputs(37));
    layer0_outputs(4588) <= not(inputs(22)) or (inputs(207));
    layer0_outputs(4589) <= not((inputs(3)) and (inputs(233)));
    layer0_outputs(4590) <= inputs(104);
    layer0_outputs(4591) <= not((inputs(19)) and (inputs(254)));
    layer0_outputs(4592) <= not(inputs(165)) or (inputs(232));
    layer0_outputs(4593) <= (inputs(140)) xor (inputs(8));
    layer0_outputs(4594) <= (inputs(134)) or (inputs(122));
    layer0_outputs(4595) <= not((inputs(127)) or (inputs(231)));
    layer0_outputs(4596) <= (inputs(151)) and not (inputs(51));
    layer0_outputs(4597) <= not((inputs(208)) and (inputs(26)));
    layer0_outputs(4598) <= not((inputs(175)) or (inputs(40)));
    layer0_outputs(4599) <= not((inputs(131)) xor (inputs(168)));
    layer0_outputs(4600) <= not((inputs(198)) or (inputs(227)));
    layer0_outputs(4601) <= (inputs(23)) or (inputs(182));
    layer0_outputs(4602) <= (inputs(180)) and not (inputs(4));
    layer0_outputs(4603) <= inputs(156);
    layer0_outputs(4604) <= '1';
    layer0_outputs(4605) <= (inputs(115)) xor (inputs(65));
    layer0_outputs(4606) <= not((inputs(246)) and (inputs(145)));
    layer0_outputs(4607) <= not(inputs(254)) or (inputs(36));
    layer0_outputs(4608) <= inputs(11);
    layer0_outputs(4609) <= (inputs(235)) or (inputs(162));
    layer0_outputs(4610) <= (inputs(30)) and not (inputs(19));
    layer0_outputs(4611) <= not(inputs(170)) or (inputs(235));
    layer0_outputs(4612) <= (inputs(148)) or (inputs(202));
    layer0_outputs(4613) <= not(inputs(39));
    layer0_outputs(4614) <= inputs(104);
    layer0_outputs(4615) <= (inputs(247)) and not (inputs(124));
    layer0_outputs(4616) <= '1';
    layer0_outputs(4617) <= '1';
    layer0_outputs(4618) <= inputs(60);
    layer0_outputs(4619) <= (inputs(139)) or (inputs(61));
    layer0_outputs(4620) <= not(inputs(244));
    layer0_outputs(4621) <= inputs(118);
    layer0_outputs(4622) <= (inputs(244)) xor (inputs(109));
    layer0_outputs(4623) <= not((inputs(235)) xor (inputs(237)));
    layer0_outputs(4624) <= (inputs(75)) xor (inputs(178));
    layer0_outputs(4625) <= not((inputs(98)) xor (inputs(162)));
    layer0_outputs(4626) <= not((inputs(165)) or (inputs(27)));
    layer0_outputs(4627) <= '1';
    layer0_outputs(4628) <= (inputs(102)) and not (inputs(184));
    layer0_outputs(4629) <= not(inputs(154)) or (inputs(128));
    layer0_outputs(4630) <= not(inputs(70));
    layer0_outputs(4631) <= '0';
    layer0_outputs(4632) <= not((inputs(166)) or (inputs(189)));
    layer0_outputs(4633) <= not(inputs(181));
    layer0_outputs(4634) <= not(inputs(179)) or (inputs(243));
    layer0_outputs(4635) <= (inputs(238)) xor (inputs(227));
    layer0_outputs(4636) <= not((inputs(113)) and (inputs(227)));
    layer0_outputs(4637) <= not(inputs(24));
    layer0_outputs(4638) <= inputs(183);
    layer0_outputs(4639) <= not((inputs(129)) xor (inputs(207)));
    layer0_outputs(4640) <= (inputs(232)) and not (inputs(169));
    layer0_outputs(4641) <= inputs(81);
    layer0_outputs(4642) <= not((inputs(159)) and (inputs(45)));
    layer0_outputs(4643) <= (inputs(59)) and not (inputs(28));
    layer0_outputs(4644) <= not(inputs(109)) or (inputs(9));
    layer0_outputs(4645) <= (inputs(174)) or (inputs(142));
    layer0_outputs(4646) <= '0';
    layer0_outputs(4647) <= (inputs(219)) and (inputs(198));
    layer0_outputs(4648) <= (inputs(193)) and not (inputs(58));
    layer0_outputs(4649) <= (inputs(200)) and not (inputs(157));
    layer0_outputs(4650) <= '0';
    layer0_outputs(4651) <= (inputs(53)) and not (inputs(166));
    layer0_outputs(4652) <= not((inputs(96)) and (inputs(128)));
    layer0_outputs(4653) <= not(inputs(160)) or (inputs(2));
    layer0_outputs(4654) <= (inputs(45)) or (inputs(132));
    layer0_outputs(4655) <= (inputs(46)) and not (inputs(27));
    layer0_outputs(4656) <= inputs(83);
    layer0_outputs(4657) <= not(inputs(104)) or (inputs(163));
    layer0_outputs(4658) <= inputs(222);
    layer0_outputs(4659) <= (inputs(243)) or (inputs(64));
    layer0_outputs(4660) <= not(inputs(63)) or (inputs(2));
    layer0_outputs(4661) <= inputs(120);
    layer0_outputs(4662) <= inputs(178);
    layer0_outputs(4663) <= (inputs(46)) xor (inputs(43));
    layer0_outputs(4664) <= (inputs(90)) and not (inputs(20));
    layer0_outputs(4665) <= (inputs(71)) and not (inputs(0));
    layer0_outputs(4666) <= not(inputs(217));
    layer0_outputs(4667) <= '1';
    layer0_outputs(4668) <= inputs(151);
    layer0_outputs(4669) <= not(inputs(54));
    layer0_outputs(4670) <= not(inputs(109)) or (inputs(165));
    layer0_outputs(4671) <= (inputs(202)) or (inputs(226));
    layer0_outputs(4672) <= not(inputs(166));
    layer0_outputs(4673) <= not((inputs(56)) or (inputs(17)));
    layer0_outputs(4674) <= inputs(163);
    layer0_outputs(4675) <= not(inputs(229)) or (inputs(67));
    layer0_outputs(4676) <= inputs(136);
    layer0_outputs(4677) <= not((inputs(160)) or (inputs(120)));
    layer0_outputs(4678) <= not(inputs(45));
    layer0_outputs(4679) <= '1';
    layer0_outputs(4680) <= inputs(168);
    layer0_outputs(4681) <= (inputs(74)) or (inputs(130));
    layer0_outputs(4682) <= not((inputs(67)) and (inputs(202)));
    layer0_outputs(4683) <= not((inputs(122)) xor (inputs(113)));
    layer0_outputs(4684) <= (inputs(199)) or (inputs(172));
    layer0_outputs(4685) <= inputs(238);
    layer0_outputs(4686) <= not(inputs(218));
    layer0_outputs(4687) <= not(inputs(236)) or (inputs(179));
    layer0_outputs(4688) <= not(inputs(230)) or (inputs(23));
    layer0_outputs(4689) <= inputs(73);
    layer0_outputs(4690) <= (inputs(7)) and (inputs(168));
    layer0_outputs(4691) <= inputs(169);
    layer0_outputs(4692) <= not((inputs(42)) xor (inputs(38)));
    layer0_outputs(4693) <= not((inputs(31)) xor (inputs(197)));
    layer0_outputs(4694) <= not(inputs(39)) or (inputs(140));
    layer0_outputs(4695) <= '1';
    layer0_outputs(4696) <= not(inputs(87));
    layer0_outputs(4697) <= not(inputs(71)) or (inputs(216));
    layer0_outputs(4698) <= not(inputs(41)) or (inputs(61));
    layer0_outputs(4699) <= (inputs(29)) or (inputs(61));
    layer0_outputs(4700) <= not(inputs(122)) or (inputs(82));
    layer0_outputs(4701) <= (inputs(166)) and not (inputs(103));
    layer0_outputs(4702) <= not(inputs(72));
    layer0_outputs(4703) <= not(inputs(153)) or (inputs(113));
    layer0_outputs(4704) <= '1';
    layer0_outputs(4705) <= (inputs(6)) xor (inputs(69));
    layer0_outputs(4706) <= not(inputs(144)) or (inputs(229));
    layer0_outputs(4707) <= (inputs(47)) xor (inputs(239));
    layer0_outputs(4708) <= not((inputs(0)) and (inputs(106)));
    layer0_outputs(4709) <= inputs(86);
    layer0_outputs(4710) <= not(inputs(237));
    layer0_outputs(4711) <= not(inputs(83)) or (inputs(10));
    layer0_outputs(4712) <= inputs(14);
    layer0_outputs(4713) <= (inputs(164)) and not (inputs(67));
    layer0_outputs(4714) <= not((inputs(131)) or (inputs(142)));
    layer0_outputs(4715) <= not(inputs(155)) or (inputs(61));
    layer0_outputs(4716) <= inputs(184);
    layer0_outputs(4717) <= (inputs(254)) xor (inputs(12));
    layer0_outputs(4718) <= inputs(98);
    layer0_outputs(4719) <= (inputs(129)) and not (inputs(24));
    layer0_outputs(4720) <= (inputs(24)) xor (inputs(159));
    layer0_outputs(4721) <= not((inputs(244)) or (inputs(227)));
    layer0_outputs(4722) <= not((inputs(24)) xor (inputs(220)));
    layer0_outputs(4723) <= not(inputs(30));
    layer0_outputs(4724) <= not((inputs(162)) or (inputs(28)));
    layer0_outputs(4725) <= '1';
    layer0_outputs(4726) <= not((inputs(97)) xor (inputs(62)));
    layer0_outputs(4727) <= inputs(121);
    layer0_outputs(4728) <= (inputs(85)) or (inputs(134));
    layer0_outputs(4729) <= not((inputs(14)) and (inputs(126)));
    layer0_outputs(4730) <= not(inputs(174));
    layer0_outputs(4731) <= not(inputs(114)) or (inputs(252));
    layer0_outputs(4732) <= (inputs(173)) and not (inputs(30));
    layer0_outputs(4733) <= '1';
    layer0_outputs(4734) <= not(inputs(158));
    layer0_outputs(4735) <= (inputs(223)) xor (inputs(19));
    layer0_outputs(4736) <= (inputs(111)) and (inputs(234));
    layer0_outputs(4737) <= not((inputs(220)) or (inputs(53)));
    layer0_outputs(4738) <= not((inputs(168)) or (inputs(41)));
    layer0_outputs(4739) <= (inputs(78)) or (inputs(222));
    layer0_outputs(4740) <= (inputs(203)) xor (inputs(157));
    layer0_outputs(4741) <= inputs(152);
    layer0_outputs(4742) <= not(inputs(42));
    layer0_outputs(4743) <= not(inputs(252)) or (inputs(132));
    layer0_outputs(4744) <= not((inputs(158)) or (inputs(138)));
    layer0_outputs(4745) <= not(inputs(185));
    layer0_outputs(4746) <= not(inputs(148));
    layer0_outputs(4747) <= (inputs(132)) xor (inputs(91));
    layer0_outputs(4748) <= not(inputs(101)) or (inputs(197));
    layer0_outputs(4749) <= not(inputs(243));
    layer0_outputs(4750) <= '1';
    layer0_outputs(4751) <= not((inputs(183)) and (inputs(194)));
    layer0_outputs(4752) <= (inputs(232)) and not (inputs(77));
    layer0_outputs(4753) <= not(inputs(117));
    layer0_outputs(4754) <= (inputs(59)) and not (inputs(227));
    layer0_outputs(4755) <= inputs(196);
    layer0_outputs(4756) <= inputs(181);
    layer0_outputs(4757) <= not(inputs(150)) or (inputs(35));
    layer0_outputs(4758) <= (inputs(162)) or (inputs(231));
    layer0_outputs(4759) <= not((inputs(41)) or (inputs(66)));
    layer0_outputs(4760) <= not((inputs(158)) xor (inputs(221)));
    layer0_outputs(4761) <= not(inputs(61));
    layer0_outputs(4762) <= inputs(131);
    layer0_outputs(4763) <= inputs(118);
    layer0_outputs(4764) <= (inputs(253)) and not (inputs(252));
    layer0_outputs(4765) <= (inputs(197)) and not (inputs(165));
    layer0_outputs(4766) <= not((inputs(244)) or (inputs(81)));
    layer0_outputs(4767) <= '1';
    layer0_outputs(4768) <= not(inputs(53));
    layer0_outputs(4769) <= (inputs(162)) or (inputs(165));
    layer0_outputs(4770) <= not(inputs(28)) or (inputs(4));
    layer0_outputs(4771) <= not(inputs(47)) or (inputs(175));
    layer0_outputs(4772) <= inputs(118);
    layer0_outputs(4773) <= '1';
    layer0_outputs(4774) <= not((inputs(8)) xor (inputs(150)));
    layer0_outputs(4775) <= not(inputs(178)) or (inputs(130));
    layer0_outputs(4776) <= (inputs(122)) or (inputs(126));
    layer0_outputs(4777) <= not(inputs(45)) or (inputs(134));
    layer0_outputs(4778) <= (inputs(22)) and not (inputs(66));
    layer0_outputs(4779) <= not(inputs(180));
    layer0_outputs(4780) <= (inputs(185)) and not (inputs(16));
    layer0_outputs(4781) <= (inputs(21)) or (inputs(8));
    layer0_outputs(4782) <= not(inputs(73)) or (inputs(20));
    layer0_outputs(4783) <= (inputs(232)) xor (inputs(253));
    layer0_outputs(4784) <= (inputs(95)) xor (inputs(179));
    layer0_outputs(4785) <= inputs(56);
    layer0_outputs(4786) <= (inputs(191)) and not (inputs(60));
    layer0_outputs(4787) <= not((inputs(204)) or (inputs(90)));
    layer0_outputs(4788) <= not(inputs(134)) or (inputs(245));
    layer0_outputs(4789) <= not((inputs(49)) or (inputs(145)));
    layer0_outputs(4790) <= not((inputs(229)) xor (inputs(214)));
    layer0_outputs(4791) <= inputs(153);
    layer0_outputs(4792) <= '0';
    layer0_outputs(4793) <= (inputs(223)) and not (inputs(108));
    layer0_outputs(4794) <= '1';
    layer0_outputs(4795) <= (inputs(15)) xor (inputs(226));
    layer0_outputs(4796) <= not((inputs(33)) xor (inputs(43)));
    layer0_outputs(4797) <= (inputs(166)) or (inputs(19));
    layer0_outputs(4798) <= not(inputs(165));
    layer0_outputs(4799) <= not(inputs(143)) or (inputs(63));
    layer0_outputs(4800) <= inputs(197);
    layer0_outputs(4801) <= not(inputs(90));
    layer0_outputs(4802) <= inputs(191);
    layer0_outputs(4803) <= (inputs(89)) or (inputs(151));
    layer0_outputs(4804) <= not(inputs(33)) or (inputs(246));
    layer0_outputs(4805) <= not((inputs(229)) or (inputs(167)));
    layer0_outputs(4806) <= not(inputs(100));
    layer0_outputs(4807) <= inputs(216);
    layer0_outputs(4808) <= (inputs(184)) xor (inputs(43));
    layer0_outputs(4809) <= not((inputs(89)) and (inputs(255)));
    layer0_outputs(4810) <= not(inputs(21));
    layer0_outputs(4811) <= (inputs(134)) or (inputs(126));
    layer0_outputs(4812) <= not((inputs(249)) and (inputs(231)));
    layer0_outputs(4813) <= '1';
    layer0_outputs(4814) <= not(inputs(185)) or (inputs(59));
    layer0_outputs(4815) <= '1';
    layer0_outputs(4816) <= (inputs(59)) xor (inputs(146));
    layer0_outputs(4817) <= not((inputs(224)) or (inputs(33)));
    layer0_outputs(4818) <= (inputs(198)) xor (inputs(144));
    layer0_outputs(4819) <= not(inputs(205));
    layer0_outputs(4820) <= (inputs(198)) xor (inputs(110));
    layer0_outputs(4821) <= '1';
    layer0_outputs(4822) <= '1';
    layer0_outputs(4823) <= not(inputs(172));
    layer0_outputs(4824) <= '1';
    layer0_outputs(4825) <= not(inputs(81));
    layer0_outputs(4826) <= (inputs(168)) xor (inputs(59));
    layer0_outputs(4827) <= not(inputs(228));
    layer0_outputs(4828) <= (inputs(18)) and not (inputs(188));
    layer0_outputs(4829) <= (inputs(238)) and (inputs(114));
    layer0_outputs(4830) <= not(inputs(73)) or (inputs(43));
    layer0_outputs(4831) <= (inputs(155)) xor (inputs(118));
    layer0_outputs(4832) <= '0';
    layer0_outputs(4833) <= (inputs(207)) xor (inputs(215));
    layer0_outputs(4834) <= (inputs(57)) and not (inputs(103));
    layer0_outputs(4835) <= not((inputs(190)) or (inputs(63)));
    layer0_outputs(4836) <= not((inputs(201)) and (inputs(43)));
    layer0_outputs(4837) <= not((inputs(217)) or (inputs(143)));
    layer0_outputs(4838) <= inputs(88);
    layer0_outputs(4839) <= inputs(33);
    layer0_outputs(4840) <= not((inputs(59)) and (inputs(249)));
    layer0_outputs(4841) <= not(inputs(120));
    layer0_outputs(4842) <= not(inputs(101));
    layer0_outputs(4843) <= not(inputs(167));
    layer0_outputs(4844) <= (inputs(178)) or (inputs(241));
    layer0_outputs(4845) <= (inputs(19)) or (inputs(104));
    layer0_outputs(4846) <= not((inputs(21)) xor (inputs(95)));
    layer0_outputs(4847) <= not(inputs(90)) or (inputs(218));
    layer0_outputs(4848) <= (inputs(36)) and not (inputs(203));
    layer0_outputs(4849) <= (inputs(113)) or (inputs(84));
    layer0_outputs(4850) <= (inputs(238)) or (inputs(69));
    layer0_outputs(4851) <= not(inputs(220));
    layer0_outputs(4852) <= not((inputs(110)) or (inputs(201)));
    layer0_outputs(4853) <= not((inputs(184)) and (inputs(207)));
    layer0_outputs(4854) <= '1';
    layer0_outputs(4855) <= not(inputs(105)) or (inputs(7));
    layer0_outputs(4856) <= not(inputs(123));
    layer0_outputs(4857) <= (inputs(88)) and (inputs(114));
    layer0_outputs(4858) <= not((inputs(236)) or (inputs(212)));
    layer0_outputs(4859) <= not((inputs(96)) or (inputs(105)));
    layer0_outputs(4860) <= (inputs(121)) xor (inputs(9));
    layer0_outputs(4861) <= not(inputs(141)) or (inputs(23));
    layer0_outputs(4862) <= not((inputs(219)) or (inputs(132)));
    layer0_outputs(4863) <= not((inputs(232)) or (inputs(94)));
    layer0_outputs(4864) <= inputs(111);
    layer0_outputs(4865) <= not((inputs(20)) and (inputs(198)));
    layer0_outputs(4866) <= (inputs(24)) xor (inputs(2));
    layer0_outputs(4867) <= not((inputs(65)) and (inputs(233)));
    layer0_outputs(4868) <= inputs(147);
    layer0_outputs(4869) <= not(inputs(127));
    layer0_outputs(4870) <= '1';
    layer0_outputs(4871) <= not(inputs(86));
    layer0_outputs(4872) <= (inputs(185)) and (inputs(244));
    layer0_outputs(4873) <= not(inputs(202));
    layer0_outputs(4874) <= (inputs(13)) xor (inputs(130));
    layer0_outputs(4875) <= not(inputs(105));
    layer0_outputs(4876) <= inputs(188);
    layer0_outputs(4877) <= (inputs(201)) and not (inputs(194));
    layer0_outputs(4878) <= not((inputs(79)) and (inputs(195)));
    layer0_outputs(4879) <= not(inputs(236));
    layer0_outputs(4880) <= not((inputs(112)) and (inputs(245)));
    layer0_outputs(4881) <= (inputs(200)) and not (inputs(17));
    layer0_outputs(4882) <= '0';
    layer0_outputs(4883) <= '0';
    layer0_outputs(4884) <= not(inputs(234)) or (inputs(37));
    layer0_outputs(4885) <= (inputs(82)) and not (inputs(142));
    layer0_outputs(4886) <= not((inputs(144)) or (inputs(104)));
    layer0_outputs(4887) <= not((inputs(230)) xor (inputs(114)));
    layer0_outputs(4888) <= not((inputs(64)) or (inputs(19)));
    layer0_outputs(4889) <= (inputs(41)) and not (inputs(84));
    layer0_outputs(4890) <= (inputs(72)) and not (inputs(23));
    layer0_outputs(4891) <= not((inputs(74)) or (inputs(214)));
    layer0_outputs(4892) <= (inputs(71)) and (inputs(201));
    layer0_outputs(4893) <= not((inputs(9)) xor (inputs(103)));
    layer0_outputs(4894) <= (inputs(247)) and not (inputs(198));
    layer0_outputs(4895) <= not((inputs(145)) or (inputs(177)));
    layer0_outputs(4896) <= not((inputs(66)) and (inputs(58)));
    layer0_outputs(4897) <= inputs(71);
    layer0_outputs(4898) <= not(inputs(53)) or (inputs(207));
    layer0_outputs(4899) <= (inputs(36)) and not (inputs(40));
    layer0_outputs(4900) <= not((inputs(1)) or (inputs(254)));
    layer0_outputs(4901) <= not(inputs(115)) or (inputs(46));
    layer0_outputs(4902) <= '1';
    layer0_outputs(4903) <= not((inputs(143)) and (inputs(216)));
    layer0_outputs(4904) <= not(inputs(37));
    layer0_outputs(4905) <= (inputs(254)) or (inputs(103));
    layer0_outputs(4906) <= inputs(75);
    layer0_outputs(4907) <= inputs(88);
    layer0_outputs(4908) <= not((inputs(54)) or (inputs(127)));
    layer0_outputs(4909) <= not((inputs(164)) xor (inputs(6)));
    layer0_outputs(4910) <= not(inputs(56)) or (inputs(188));
    layer0_outputs(4911) <= not((inputs(54)) or (inputs(104)));
    layer0_outputs(4912) <= inputs(152);
    layer0_outputs(4913) <= inputs(254);
    layer0_outputs(4914) <= not((inputs(45)) and (inputs(171)));
    layer0_outputs(4915) <= (inputs(129)) xor (inputs(168));
    layer0_outputs(4916) <= (inputs(7)) or (inputs(179));
    layer0_outputs(4917) <= not(inputs(13)) or (inputs(66));
    layer0_outputs(4918) <= not((inputs(240)) or (inputs(141)));
    layer0_outputs(4919) <= not(inputs(122));
    layer0_outputs(4920) <= '0';
    layer0_outputs(4921) <= (inputs(78)) xor (inputs(119));
    layer0_outputs(4922) <= (inputs(164)) and not (inputs(244));
    layer0_outputs(4923) <= (inputs(202)) and not (inputs(62));
    layer0_outputs(4924) <= '1';
    layer0_outputs(4925) <= inputs(61);
    layer0_outputs(4926) <= inputs(225);
    layer0_outputs(4927) <= '0';
    layer0_outputs(4928) <= (inputs(38)) xor (inputs(196));
    layer0_outputs(4929) <= '0';
    layer0_outputs(4930) <= (inputs(40)) or (inputs(38));
    layer0_outputs(4931) <= '0';
    layer0_outputs(4932) <= inputs(155);
    layer0_outputs(4933) <= not(inputs(253)) or (inputs(185));
    layer0_outputs(4934) <= not(inputs(183)) or (inputs(59));
    layer0_outputs(4935) <= (inputs(54)) and not (inputs(159));
    layer0_outputs(4936) <= not((inputs(39)) xor (inputs(141)));
    layer0_outputs(4937) <= not(inputs(15));
    layer0_outputs(4938) <= not((inputs(98)) or (inputs(83)));
    layer0_outputs(4939) <= not((inputs(88)) or (inputs(250)));
    layer0_outputs(4940) <= (inputs(129)) and (inputs(215));
    layer0_outputs(4941) <= inputs(198);
    layer0_outputs(4942) <= not((inputs(189)) or (inputs(216)));
    layer0_outputs(4943) <= not((inputs(70)) or (inputs(231)));
    layer0_outputs(4944) <= (inputs(220)) and not (inputs(36));
    layer0_outputs(4945) <= (inputs(59)) and (inputs(64));
    layer0_outputs(4946) <= (inputs(79)) or (inputs(236));
    layer0_outputs(4947) <= not(inputs(246)) or (inputs(5));
    layer0_outputs(4948) <= (inputs(54)) xor (inputs(103));
    layer0_outputs(4949) <= not(inputs(213)) or (inputs(96));
    layer0_outputs(4950) <= (inputs(111)) or (inputs(38));
    layer0_outputs(4951) <= not((inputs(177)) or (inputs(107)));
    layer0_outputs(4952) <= not(inputs(215)) or (inputs(202));
    layer0_outputs(4953) <= not(inputs(41));
    layer0_outputs(4954) <= inputs(94);
    layer0_outputs(4955) <= inputs(143);
    layer0_outputs(4956) <= inputs(15);
    layer0_outputs(4957) <= inputs(72);
    layer0_outputs(4958) <= inputs(22);
    layer0_outputs(4959) <= not(inputs(30)) or (inputs(140));
    layer0_outputs(4960) <= (inputs(102)) and not (inputs(251));
    layer0_outputs(4961) <= inputs(108);
    layer0_outputs(4962) <= not((inputs(153)) xor (inputs(1)));
    layer0_outputs(4963) <= not(inputs(158));
    layer0_outputs(4964) <= not((inputs(44)) or (inputs(238)));
    layer0_outputs(4965) <= not(inputs(100));
    layer0_outputs(4966) <= not(inputs(106)) or (inputs(34));
    layer0_outputs(4967) <= not(inputs(121));
    layer0_outputs(4968) <= not(inputs(59));
    layer0_outputs(4969) <= not((inputs(248)) or (inputs(191)));
    layer0_outputs(4970) <= not(inputs(116));
    layer0_outputs(4971) <= inputs(224);
    layer0_outputs(4972) <= not((inputs(36)) xor (inputs(163)));
    layer0_outputs(4973) <= not(inputs(67)) or (inputs(26));
    layer0_outputs(4974) <= not(inputs(43)) or (inputs(70));
    layer0_outputs(4975) <= (inputs(140)) and not (inputs(52));
    layer0_outputs(4976) <= inputs(130);
    layer0_outputs(4977) <= not(inputs(207)) or (inputs(114));
    layer0_outputs(4978) <= not((inputs(38)) or (inputs(17)));
    layer0_outputs(4979) <= (inputs(26)) and not (inputs(222));
    layer0_outputs(4980) <= not(inputs(85)) or (inputs(182));
    layer0_outputs(4981) <= not((inputs(77)) or (inputs(43)));
    layer0_outputs(4982) <= not(inputs(214));
    layer0_outputs(4983) <= not((inputs(197)) or (inputs(220)));
    layer0_outputs(4984) <= inputs(159);
    layer0_outputs(4985) <= '0';
    layer0_outputs(4986) <= not(inputs(42));
    layer0_outputs(4987) <= '1';
    layer0_outputs(4988) <= inputs(118);
    layer0_outputs(4989) <= not(inputs(119)) or (inputs(67));
    layer0_outputs(4990) <= not(inputs(141)) or (inputs(46));
    layer0_outputs(4991) <= (inputs(24)) or (inputs(165));
    layer0_outputs(4992) <= not(inputs(130)) or (inputs(18));
    layer0_outputs(4993) <= inputs(66);
    layer0_outputs(4994) <= not(inputs(142)) or (inputs(113));
    layer0_outputs(4995) <= inputs(44);
    layer0_outputs(4996) <= (inputs(1)) and not (inputs(140));
    layer0_outputs(4997) <= (inputs(105)) or (inputs(69));
    layer0_outputs(4998) <= inputs(144);
    layer0_outputs(4999) <= (inputs(55)) and not (inputs(49));
    layer0_outputs(5000) <= '1';
    layer0_outputs(5001) <= inputs(151);
    layer0_outputs(5002) <= not(inputs(250));
    layer0_outputs(5003) <= not(inputs(136));
    layer0_outputs(5004) <= not(inputs(147));
    layer0_outputs(5005) <= (inputs(49)) and not (inputs(185));
    layer0_outputs(5006) <= not(inputs(221)) or (inputs(133));
    layer0_outputs(5007) <= not(inputs(237));
    layer0_outputs(5008) <= inputs(153);
    layer0_outputs(5009) <= (inputs(120)) and (inputs(183));
    layer0_outputs(5010) <= not((inputs(127)) xor (inputs(206)));
    layer0_outputs(5011) <= not(inputs(12)) or (inputs(77));
    layer0_outputs(5012) <= not(inputs(159)) or (inputs(44));
    layer0_outputs(5013) <= not(inputs(134)) or (inputs(10));
    layer0_outputs(5014) <= not((inputs(46)) and (inputs(145)));
    layer0_outputs(5015) <= not((inputs(96)) xor (inputs(230)));
    layer0_outputs(5016) <= inputs(178);
    layer0_outputs(5017) <= not((inputs(180)) or (inputs(51)));
    layer0_outputs(5018) <= (inputs(207)) or (inputs(243));
    layer0_outputs(5019) <= not(inputs(216));
    layer0_outputs(5020) <= (inputs(25)) and not (inputs(193));
    layer0_outputs(5021) <= (inputs(216)) or (inputs(110));
    layer0_outputs(5022) <= (inputs(94)) or (inputs(38));
    layer0_outputs(5023) <= not(inputs(226)) or (inputs(66));
    layer0_outputs(5024) <= inputs(164);
    layer0_outputs(5025) <= not((inputs(70)) or (inputs(220)));
    layer0_outputs(5026) <= inputs(190);
    layer0_outputs(5027) <= not((inputs(199)) and (inputs(112)));
    layer0_outputs(5028) <= not(inputs(118)) or (inputs(233));
    layer0_outputs(5029) <= inputs(22);
    layer0_outputs(5030) <= not((inputs(131)) or (inputs(155)));
    layer0_outputs(5031) <= inputs(136);
    layer0_outputs(5032) <= '1';
    layer0_outputs(5033) <= not(inputs(143)) or (inputs(127));
    layer0_outputs(5034) <= (inputs(119)) or (inputs(255));
    layer0_outputs(5035) <= not(inputs(189));
    layer0_outputs(5036) <= (inputs(151)) and (inputs(214));
    layer0_outputs(5037) <= (inputs(5)) or (inputs(36));
    layer0_outputs(5038) <= not((inputs(34)) or (inputs(32)));
    layer0_outputs(5039) <= '1';
    layer0_outputs(5040) <= not((inputs(76)) and (inputs(211)));
    layer0_outputs(5041) <= not(inputs(207)) or (inputs(227));
    layer0_outputs(5042) <= not(inputs(138)) or (inputs(188));
    layer0_outputs(5043) <= not(inputs(181));
    layer0_outputs(5044) <= not(inputs(81));
    layer0_outputs(5045) <= (inputs(69)) xor (inputs(154));
    layer0_outputs(5046) <= not(inputs(172));
    layer0_outputs(5047) <= inputs(170);
    layer0_outputs(5048) <= (inputs(122)) xor (inputs(97));
    layer0_outputs(5049) <= inputs(26);
    layer0_outputs(5050) <= not((inputs(54)) or (inputs(170)));
    layer0_outputs(5051) <= not(inputs(242));
    layer0_outputs(5052) <= not((inputs(103)) xor (inputs(116)));
    layer0_outputs(5053) <= (inputs(187)) and not (inputs(131));
    layer0_outputs(5054) <= not(inputs(245));
    layer0_outputs(5055) <= (inputs(164)) and not (inputs(161));
    layer0_outputs(5056) <= not(inputs(216));
    layer0_outputs(5057) <= (inputs(28)) and not (inputs(175));
    layer0_outputs(5058) <= (inputs(166)) or (inputs(166));
    layer0_outputs(5059) <= (inputs(198)) and not (inputs(49));
    layer0_outputs(5060) <= (inputs(49)) and (inputs(247));
    layer0_outputs(5061) <= (inputs(101)) and not (inputs(175));
    layer0_outputs(5062) <= inputs(105);
    layer0_outputs(5063) <= not(inputs(104)) or (inputs(115));
    layer0_outputs(5064) <= inputs(138);
    layer0_outputs(5065) <= not(inputs(74)) or (inputs(255));
    layer0_outputs(5066) <= (inputs(214)) and (inputs(206));
    layer0_outputs(5067) <= inputs(23);
    layer0_outputs(5068) <= (inputs(70)) and not (inputs(25));
    layer0_outputs(5069) <= '1';
    layer0_outputs(5070) <= not((inputs(255)) or (inputs(216)));
    layer0_outputs(5071) <= (inputs(166)) and not (inputs(115));
    layer0_outputs(5072) <= (inputs(53)) and not (inputs(236));
    layer0_outputs(5073) <= '0';
    layer0_outputs(5074) <= '0';
    layer0_outputs(5075) <= not((inputs(129)) xor (inputs(90)));
    layer0_outputs(5076) <= not((inputs(83)) xor (inputs(143)));
    layer0_outputs(5077) <= (inputs(231)) or (inputs(75));
    layer0_outputs(5078) <= (inputs(156)) and not (inputs(65));
    layer0_outputs(5079) <= not(inputs(119)) or (inputs(158));
    layer0_outputs(5080) <= (inputs(176)) and not (inputs(190));
    layer0_outputs(5081) <= '1';
    layer0_outputs(5082) <= not(inputs(193));
    layer0_outputs(5083) <= not((inputs(227)) xor (inputs(178)));
    layer0_outputs(5084) <= not((inputs(255)) or (inputs(150)));
    layer0_outputs(5085) <= '0';
    layer0_outputs(5086) <= inputs(234);
    layer0_outputs(5087) <= '1';
    layer0_outputs(5088) <= not(inputs(174)) or (inputs(143));
    layer0_outputs(5089) <= not(inputs(1));
    layer0_outputs(5090) <= '1';
    layer0_outputs(5091) <= not(inputs(62));
    layer0_outputs(5092) <= not(inputs(191)) or (inputs(69));
    layer0_outputs(5093) <= (inputs(174)) and not (inputs(131));
    layer0_outputs(5094) <= not(inputs(95)) or (inputs(96));
    layer0_outputs(5095) <= inputs(40);
    layer0_outputs(5096) <= not((inputs(164)) xor (inputs(63)));
    layer0_outputs(5097) <= not(inputs(132));
    layer0_outputs(5098) <= not(inputs(26));
    layer0_outputs(5099) <= (inputs(159)) and not (inputs(244));
    layer0_outputs(5100) <= not((inputs(189)) xor (inputs(129)));
    layer0_outputs(5101) <= (inputs(187)) xor (inputs(97));
    layer0_outputs(5102) <= inputs(150);
    layer0_outputs(5103) <= inputs(234);
    layer0_outputs(5104) <= not((inputs(74)) xor (inputs(98)));
    layer0_outputs(5105) <= (inputs(127)) and not (inputs(227));
    layer0_outputs(5106) <= not(inputs(87)) or (inputs(224));
    layer0_outputs(5107) <= not(inputs(127));
    layer0_outputs(5108) <= inputs(92);
    layer0_outputs(5109) <= (inputs(10)) and not (inputs(87));
    layer0_outputs(5110) <= inputs(113);
    layer0_outputs(5111) <= (inputs(225)) and (inputs(62));
    layer0_outputs(5112) <= (inputs(230)) xor (inputs(108));
    layer0_outputs(5113) <= not(inputs(135));
    layer0_outputs(5114) <= inputs(120);
    layer0_outputs(5115) <= (inputs(99)) and (inputs(128));
    layer0_outputs(5116) <= (inputs(136)) and not (inputs(43));
    layer0_outputs(5117) <= not(inputs(175)) or (inputs(129));
    layer0_outputs(5118) <= not((inputs(108)) or (inputs(132)));
    layer0_outputs(5119) <= not((inputs(142)) xor (inputs(187)));
    layer1_outputs(0) <= (layer0_outputs(2850)) or (layer0_outputs(1993));
    layer1_outputs(1) <= (layer0_outputs(2438)) xor (layer0_outputs(317));
    layer1_outputs(2) <= not(layer0_outputs(5058));
    layer1_outputs(3) <= (layer0_outputs(2787)) and (layer0_outputs(2481));
    layer1_outputs(4) <= not((layer0_outputs(1935)) or (layer0_outputs(3628)));
    layer1_outputs(5) <= layer0_outputs(1583);
    layer1_outputs(6) <= (layer0_outputs(1117)) or (layer0_outputs(1988));
    layer1_outputs(7) <= not(layer0_outputs(3902));
    layer1_outputs(8) <= (layer0_outputs(480)) and not (layer0_outputs(98));
    layer1_outputs(9) <= not(layer0_outputs(1435)) or (layer0_outputs(2329));
    layer1_outputs(10) <= not(layer0_outputs(2093));
    layer1_outputs(11) <= (layer0_outputs(2648)) xor (layer0_outputs(631));
    layer1_outputs(12) <= not(layer0_outputs(589));
    layer1_outputs(13) <= (layer0_outputs(2928)) and not (layer0_outputs(5041));
    layer1_outputs(14) <= layer0_outputs(4744);
    layer1_outputs(15) <= layer0_outputs(4536);
    layer1_outputs(16) <= layer0_outputs(4171);
    layer1_outputs(17) <= not(layer0_outputs(3913));
    layer1_outputs(18) <= layer0_outputs(4628);
    layer1_outputs(19) <= (layer0_outputs(226)) and not (layer0_outputs(3657));
    layer1_outputs(20) <= not(layer0_outputs(1362));
    layer1_outputs(21) <= not((layer0_outputs(4956)) and (layer0_outputs(781)));
    layer1_outputs(22) <= not((layer0_outputs(4449)) xor (layer0_outputs(90)));
    layer1_outputs(23) <= (layer0_outputs(4373)) and (layer0_outputs(2894));
    layer1_outputs(24) <= not(layer0_outputs(1165)) or (layer0_outputs(1653));
    layer1_outputs(25) <= (layer0_outputs(803)) or (layer0_outputs(1626));
    layer1_outputs(26) <= (layer0_outputs(2552)) or (layer0_outputs(2828));
    layer1_outputs(27) <= layer0_outputs(1317);
    layer1_outputs(28) <= (layer0_outputs(4081)) and not (layer0_outputs(3383));
    layer1_outputs(29) <= layer0_outputs(2736);
    layer1_outputs(30) <= (layer0_outputs(1737)) or (layer0_outputs(1491));
    layer1_outputs(31) <= not(layer0_outputs(1672)) or (layer0_outputs(3761));
    layer1_outputs(32) <= layer0_outputs(3263);
    layer1_outputs(33) <= not(layer0_outputs(3026));
    layer1_outputs(34) <= layer0_outputs(3495);
    layer1_outputs(35) <= not(layer0_outputs(2689));
    layer1_outputs(36) <= not(layer0_outputs(2848));
    layer1_outputs(37) <= not((layer0_outputs(532)) xor (layer0_outputs(3800)));
    layer1_outputs(38) <= not(layer0_outputs(4210)) or (layer0_outputs(1865));
    layer1_outputs(39) <= not((layer0_outputs(4749)) xor (layer0_outputs(3270)));
    layer1_outputs(40) <= layer0_outputs(1372);
    layer1_outputs(41) <= layer0_outputs(4010);
    layer1_outputs(42) <= (layer0_outputs(151)) xor (layer0_outputs(4498));
    layer1_outputs(43) <= (layer0_outputs(2766)) and (layer0_outputs(4577));
    layer1_outputs(44) <= (layer0_outputs(3789)) and not (layer0_outputs(1295));
    layer1_outputs(45) <= not(layer0_outputs(3046));
    layer1_outputs(46) <= (layer0_outputs(1948)) or (layer0_outputs(697));
    layer1_outputs(47) <= layer0_outputs(1299);
    layer1_outputs(48) <= not((layer0_outputs(3590)) and (layer0_outputs(2553)));
    layer1_outputs(49) <= not(layer0_outputs(303)) or (layer0_outputs(985));
    layer1_outputs(50) <= not((layer0_outputs(2314)) xor (layer0_outputs(1958)));
    layer1_outputs(51) <= (layer0_outputs(1230)) or (layer0_outputs(2882));
    layer1_outputs(52) <= not(layer0_outputs(1887));
    layer1_outputs(53) <= (layer0_outputs(4120)) and not (layer0_outputs(200));
    layer1_outputs(54) <= (layer0_outputs(1430)) and not (layer0_outputs(5063));
    layer1_outputs(55) <= layer0_outputs(1604);
    layer1_outputs(56) <= not((layer0_outputs(1302)) or (layer0_outputs(1723)));
    layer1_outputs(57) <= not(layer0_outputs(3752)) or (layer0_outputs(4024));
    layer1_outputs(58) <= not(layer0_outputs(3172)) or (layer0_outputs(3617));
    layer1_outputs(59) <= not(layer0_outputs(598)) or (layer0_outputs(4379));
    layer1_outputs(60) <= not(layer0_outputs(822)) or (layer0_outputs(4382));
    layer1_outputs(61) <= (layer0_outputs(1708)) or (layer0_outputs(2000));
    layer1_outputs(62) <= not(layer0_outputs(4891));
    layer1_outputs(63) <= not(layer0_outputs(4213)) or (layer0_outputs(747));
    layer1_outputs(64) <= (layer0_outputs(3489)) or (layer0_outputs(1723));
    layer1_outputs(65) <= (layer0_outputs(2307)) and not (layer0_outputs(2053));
    layer1_outputs(66) <= not((layer0_outputs(2168)) and (layer0_outputs(1700)));
    layer1_outputs(67) <= layer0_outputs(2008);
    layer1_outputs(68) <= not((layer0_outputs(1123)) xor (layer0_outputs(2541)));
    layer1_outputs(69) <= not(layer0_outputs(1797));
    layer1_outputs(70) <= not((layer0_outputs(600)) and (layer0_outputs(4722)));
    layer1_outputs(71) <= (layer0_outputs(3818)) and not (layer0_outputs(4721));
    layer1_outputs(72) <= '1';
    layer1_outputs(73) <= (layer0_outputs(1647)) or (layer0_outputs(4713));
    layer1_outputs(74) <= not(layer0_outputs(3373));
    layer1_outputs(75) <= not(layer0_outputs(766));
    layer1_outputs(76) <= not((layer0_outputs(4819)) or (layer0_outputs(4100)));
    layer1_outputs(77) <= (layer0_outputs(2377)) and not (layer0_outputs(2967));
    layer1_outputs(78) <= not(layer0_outputs(878));
    layer1_outputs(79) <= not((layer0_outputs(1442)) xor (layer0_outputs(3331)));
    layer1_outputs(80) <= not((layer0_outputs(491)) or (layer0_outputs(1228)));
    layer1_outputs(81) <= (layer0_outputs(741)) and not (layer0_outputs(4293));
    layer1_outputs(82) <= (layer0_outputs(2879)) or (layer0_outputs(1035));
    layer1_outputs(83) <= not((layer0_outputs(3540)) xor (layer0_outputs(1952)));
    layer1_outputs(84) <= not(layer0_outputs(1240)) or (layer0_outputs(3203));
    layer1_outputs(85) <= not(layer0_outputs(1782));
    layer1_outputs(86) <= not(layer0_outputs(5040)) or (layer0_outputs(1863));
    layer1_outputs(87) <= layer0_outputs(777);
    layer1_outputs(88) <= '1';
    layer1_outputs(89) <= not((layer0_outputs(3147)) and (layer0_outputs(667)));
    layer1_outputs(90) <= not((layer0_outputs(385)) xor (layer0_outputs(737)));
    layer1_outputs(91) <= (layer0_outputs(3705)) and not (layer0_outputs(120));
    layer1_outputs(92) <= layer0_outputs(3632);
    layer1_outputs(93) <= not(layer0_outputs(4346)) or (layer0_outputs(3302));
    layer1_outputs(94) <= layer0_outputs(4254);
    layer1_outputs(95) <= layer0_outputs(2175);
    layer1_outputs(96) <= not((layer0_outputs(4811)) or (layer0_outputs(4045)));
    layer1_outputs(97) <= layer0_outputs(3655);
    layer1_outputs(98) <= layer0_outputs(4007);
    layer1_outputs(99) <= layer0_outputs(2183);
    layer1_outputs(100) <= not(layer0_outputs(2274));
    layer1_outputs(101) <= not(layer0_outputs(2027));
    layer1_outputs(102) <= not(layer0_outputs(1380));
    layer1_outputs(103) <= layer0_outputs(533);
    layer1_outputs(104) <= not(layer0_outputs(503));
    layer1_outputs(105) <= (layer0_outputs(3471)) and (layer0_outputs(718));
    layer1_outputs(106) <= (layer0_outputs(347)) and (layer0_outputs(204));
    layer1_outputs(107) <= layer0_outputs(2038);
    layer1_outputs(108) <= layer0_outputs(4128);
    layer1_outputs(109) <= not(layer0_outputs(1621));
    layer1_outputs(110) <= (layer0_outputs(2866)) and not (layer0_outputs(3452));
    layer1_outputs(111) <= not((layer0_outputs(4791)) and (layer0_outputs(3405)));
    layer1_outputs(112) <= not((layer0_outputs(1434)) and (layer0_outputs(1530)));
    layer1_outputs(113) <= (layer0_outputs(573)) and not (layer0_outputs(1290));
    layer1_outputs(114) <= not(layer0_outputs(1721)) or (layer0_outputs(1533));
    layer1_outputs(115) <= not(layer0_outputs(1624));
    layer1_outputs(116) <= layer0_outputs(686);
    layer1_outputs(117) <= (layer0_outputs(162)) xor (layer0_outputs(1275));
    layer1_outputs(118) <= layer0_outputs(4684);
    layer1_outputs(119) <= not(layer0_outputs(3909)) or (layer0_outputs(3965));
    layer1_outputs(120) <= not(layer0_outputs(3254)) or (layer0_outputs(3231));
    layer1_outputs(121) <= not((layer0_outputs(3460)) or (layer0_outputs(4933)));
    layer1_outputs(122) <= layer0_outputs(1673);
    layer1_outputs(123) <= not(layer0_outputs(2467));
    layer1_outputs(124) <= not((layer0_outputs(2091)) or (layer0_outputs(2694)));
    layer1_outputs(125) <= not((layer0_outputs(1804)) and (layer0_outputs(3667)));
    layer1_outputs(126) <= (layer0_outputs(2771)) and not (layer0_outputs(1056));
    layer1_outputs(127) <= not(layer0_outputs(1878));
    layer1_outputs(128) <= (layer0_outputs(4454)) and not (layer0_outputs(1889));
    layer1_outputs(129) <= not(layer0_outputs(271));
    layer1_outputs(130) <= not((layer0_outputs(2099)) and (layer0_outputs(5002)));
    layer1_outputs(131) <= not(layer0_outputs(2389)) or (layer0_outputs(1840));
    layer1_outputs(132) <= layer0_outputs(2784);
    layer1_outputs(133) <= not(layer0_outputs(887));
    layer1_outputs(134) <= (layer0_outputs(4690)) and not (layer0_outputs(1103));
    layer1_outputs(135) <= (layer0_outputs(3157)) and not (layer0_outputs(688));
    layer1_outputs(136) <= not((layer0_outputs(5044)) xor (layer0_outputs(4629)));
    layer1_outputs(137) <= not((layer0_outputs(377)) and (layer0_outputs(3495)));
    layer1_outputs(138) <= not(layer0_outputs(632)) or (layer0_outputs(212));
    layer1_outputs(139) <= (layer0_outputs(1136)) and not (layer0_outputs(1062));
    layer1_outputs(140) <= not(layer0_outputs(315)) or (layer0_outputs(3837));
    layer1_outputs(141) <= '0';
    layer1_outputs(142) <= layer0_outputs(4182);
    layer1_outputs(143) <= not(layer0_outputs(2876));
    layer1_outputs(144) <= not(layer0_outputs(1870));
    layer1_outputs(145) <= not((layer0_outputs(1377)) xor (layer0_outputs(1039)));
    layer1_outputs(146) <= layer0_outputs(326);
    layer1_outputs(147) <= (layer0_outputs(287)) and not (layer0_outputs(4083));
    layer1_outputs(148) <= layer0_outputs(4958);
    layer1_outputs(149) <= layer0_outputs(982);
    layer1_outputs(150) <= (layer0_outputs(4688)) and not (layer0_outputs(4590));
    layer1_outputs(151) <= layer0_outputs(1574);
    layer1_outputs(152) <= not(layer0_outputs(800));
    layer1_outputs(153) <= not(layer0_outputs(711)) or (layer0_outputs(4222));
    layer1_outputs(154) <= not(layer0_outputs(5113));
    layer1_outputs(155) <= not(layer0_outputs(41));
    layer1_outputs(156) <= not(layer0_outputs(3484));
    layer1_outputs(157) <= not(layer0_outputs(826));
    layer1_outputs(158) <= not(layer0_outputs(1405)) or (layer0_outputs(707));
    layer1_outputs(159) <= not((layer0_outputs(2029)) xor (layer0_outputs(4106)));
    layer1_outputs(160) <= not(layer0_outputs(1101)) or (layer0_outputs(2935));
    layer1_outputs(161) <= not(layer0_outputs(1945)) or (layer0_outputs(3421));
    layer1_outputs(162) <= not((layer0_outputs(2891)) xor (layer0_outputs(2445)));
    layer1_outputs(163) <= not((layer0_outputs(5090)) and (layer0_outputs(1081)));
    layer1_outputs(164) <= not((layer0_outputs(3939)) or (layer0_outputs(2526)));
    layer1_outputs(165) <= not(layer0_outputs(4942)) or (layer0_outputs(345));
    layer1_outputs(166) <= not(layer0_outputs(2321));
    layer1_outputs(167) <= not(layer0_outputs(2068));
    layer1_outputs(168) <= not((layer0_outputs(1267)) or (layer0_outputs(437)));
    layer1_outputs(169) <= not(layer0_outputs(4220));
    layer1_outputs(170) <= layer0_outputs(2807);
    layer1_outputs(171) <= '1';
    layer1_outputs(172) <= not((layer0_outputs(1769)) or (layer0_outputs(695)));
    layer1_outputs(173) <= not(layer0_outputs(2684));
    layer1_outputs(174) <= not(layer0_outputs(704)) or (layer0_outputs(1048));
    layer1_outputs(175) <= not(layer0_outputs(3697)) or (layer0_outputs(4967));
    layer1_outputs(176) <= (layer0_outputs(1628)) and (layer0_outputs(5007));
    layer1_outputs(177) <= not(layer0_outputs(4538));
    layer1_outputs(178) <= not(layer0_outputs(678));
    layer1_outputs(179) <= layer0_outputs(1895);
    layer1_outputs(180) <= not(layer0_outputs(720)) or (layer0_outputs(946));
    layer1_outputs(181) <= (layer0_outputs(3071)) and (layer0_outputs(666));
    layer1_outputs(182) <= (layer0_outputs(750)) or (layer0_outputs(3366));
    layer1_outputs(183) <= not(layer0_outputs(1609)) or (layer0_outputs(2482));
    layer1_outputs(184) <= (layer0_outputs(807)) or (layer0_outputs(975));
    layer1_outputs(185) <= not(layer0_outputs(2964)) or (layer0_outputs(3294));
    layer1_outputs(186) <= not(layer0_outputs(3859));
    layer1_outputs(187) <= (layer0_outputs(1427)) and (layer0_outputs(2427));
    layer1_outputs(188) <= not(layer0_outputs(2695)) or (layer0_outputs(4664));
    layer1_outputs(189) <= (layer0_outputs(2215)) xor (layer0_outputs(3759));
    layer1_outputs(190) <= layer0_outputs(1689);
    layer1_outputs(191) <= (layer0_outputs(4666)) and not (layer0_outputs(2394));
    layer1_outputs(192) <= (layer0_outputs(4992)) and not (layer0_outputs(3076));
    layer1_outputs(193) <= '1';
    layer1_outputs(194) <= (layer0_outputs(2643)) and not (layer0_outputs(4179));
    layer1_outputs(195) <= not((layer0_outputs(5104)) and (layer0_outputs(1877)));
    layer1_outputs(196) <= not((layer0_outputs(4167)) xor (layer0_outputs(3228)));
    layer1_outputs(197) <= (layer0_outputs(2231)) and not (layer0_outputs(1833));
    layer1_outputs(198) <= not((layer0_outputs(2478)) xor (layer0_outputs(3392)));
    layer1_outputs(199) <= (layer0_outputs(3320)) or (layer0_outputs(2020));
    layer1_outputs(200) <= (layer0_outputs(4599)) and (layer0_outputs(802));
    layer1_outputs(201) <= '1';
    layer1_outputs(202) <= not((layer0_outputs(608)) and (layer0_outputs(964)));
    layer1_outputs(203) <= not(layer0_outputs(582));
    layer1_outputs(204) <= not(layer0_outputs(2346));
    layer1_outputs(205) <= (layer0_outputs(4378)) and not (layer0_outputs(959));
    layer1_outputs(206) <= (layer0_outputs(951)) or (layer0_outputs(5052));
    layer1_outputs(207) <= layer0_outputs(1371);
    layer1_outputs(208) <= layer0_outputs(1513);
    layer1_outputs(209) <= '1';
    layer1_outputs(210) <= (layer0_outputs(172)) and (layer0_outputs(4879));
    layer1_outputs(211) <= not(layer0_outputs(485));
    layer1_outputs(212) <= not((layer0_outputs(2437)) xor (layer0_outputs(4131)));
    layer1_outputs(213) <= not(layer0_outputs(2495));
    layer1_outputs(214) <= not((layer0_outputs(2557)) or (layer0_outputs(3613)));
    layer1_outputs(215) <= (layer0_outputs(2252)) and not (layer0_outputs(638));
    layer1_outputs(216) <= (layer0_outputs(4004)) xor (layer0_outputs(1049));
    layer1_outputs(217) <= not((layer0_outputs(3123)) and (layer0_outputs(3738)));
    layer1_outputs(218) <= not(layer0_outputs(1948)) or (layer0_outputs(509));
    layer1_outputs(219) <= layer0_outputs(5031);
    layer1_outputs(220) <= '0';
    layer1_outputs(221) <= not((layer0_outputs(4939)) and (layer0_outputs(1569)));
    layer1_outputs(222) <= not(layer0_outputs(1593)) or (layer0_outputs(2931));
    layer1_outputs(223) <= (layer0_outputs(857)) and not (layer0_outputs(2943));
    layer1_outputs(224) <= (layer0_outputs(3474)) and not (layer0_outputs(2795));
    layer1_outputs(225) <= layer0_outputs(4186);
    layer1_outputs(226) <= not(layer0_outputs(808));
    layer1_outputs(227) <= not((layer0_outputs(47)) xor (layer0_outputs(3869)));
    layer1_outputs(228) <= not((layer0_outputs(839)) xor (layer0_outputs(766)));
    layer1_outputs(229) <= '1';
    layer1_outputs(230) <= not(layer0_outputs(297));
    layer1_outputs(231) <= not(layer0_outputs(1949));
    layer1_outputs(232) <= (layer0_outputs(1827)) and not (layer0_outputs(3107));
    layer1_outputs(233) <= not((layer0_outputs(1084)) or (layer0_outputs(1200)));
    layer1_outputs(234) <= layer0_outputs(4532);
    layer1_outputs(235) <= (layer0_outputs(4955)) and (layer0_outputs(2818));
    layer1_outputs(236) <= (layer0_outputs(2458)) and (layer0_outputs(3246));
    layer1_outputs(237) <= not(layer0_outputs(3388)) or (layer0_outputs(1079));
    layer1_outputs(238) <= (layer0_outputs(3251)) xor (layer0_outputs(342));
    layer1_outputs(239) <= layer0_outputs(3099);
    layer1_outputs(240) <= not(layer0_outputs(390));
    layer1_outputs(241) <= not(layer0_outputs(5047));
    layer1_outputs(242) <= (layer0_outputs(3406)) or (layer0_outputs(246));
    layer1_outputs(243) <= (layer0_outputs(385)) xor (layer0_outputs(1033));
    layer1_outputs(244) <= (layer0_outputs(4678)) xor (layer0_outputs(369));
    layer1_outputs(245) <= '0';
    layer1_outputs(246) <= (layer0_outputs(4758)) or (layer0_outputs(4342));
    layer1_outputs(247) <= not(layer0_outputs(954));
    layer1_outputs(248) <= (layer0_outputs(516)) and not (layer0_outputs(2777));
    layer1_outputs(249) <= not(layer0_outputs(575));
    layer1_outputs(250) <= layer0_outputs(203);
    layer1_outputs(251) <= not(layer0_outputs(143));
    layer1_outputs(252) <= not((layer0_outputs(2911)) and (layer0_outputs(1504)));
    layer1_outputs(253) <= layer0_outputs(2173);
    layer1_outputs(254) <= not(layer0_outputs(1285)) or (layer0_outputs(248));
    layer1_outputs(255) <= not(layer0_outputs(2644));
    layer1_outputs(256) <= not(layer0_outputs(980)) or (layer0_outputs(4406));
    layer1_outputs(257) <= layer0_outputs(3547);
    layer1_outputs(258) <= (layer0_outputs(1392)) or (layer0_outputs(2888));
    layer1_outputs(259) <= not(layer0_outputs(1561));
    layer1_outputs(260) <= (layer0_outputs(653)) and not (layer0_outputs(4734));
    layer1_outputs(261) <= layer0_outputs(4075);
    layer1_outputs(262) <= not((layer0_outputs(4105)) or (layer0_outputs(2706)));
    layer1_outputs(263) <= (layer0_outputs(2511)) and not (layer0_outputs(1829));
    layer1_outputs(264) <= not(layer0_outputs(709)) or (layer0_outputs(3698));
    layer1_outputs(265) <= not((layer0_outputs(881)) and (layer0_outputs(3773)));
    layer1_outputs(266) <= '1';
    layer1_outputs(267) <= layer0_outputs(3669);
    layer1_outputs(268) <= (layer0_outputs(452)) or (layer0_outputs(4068));
    layer1_outputs(269) <= (layer0_outputs(2896)) and (layer0_outputs(3754));
    layer1_outputs(270) <= not(layer0_outputs(1746));
    layer1_outputs(271) <= not(layer0_outputs(1823)) or (layer0_outputs(2845));
    layer1_outputs(272) <= (layer0_outputs(73)) and not (layer0_outputs(536));
    layer1_outputs(273) <= not((layer0_outputs(4823)) and (layer0_outputs(4306)));
    layer1_outputs(274) <= (layer0_outputs(588)) or (layer0_outputs(2455));
    layer1_outputs(275) <= not(layer0_outputs(2834)) or (layer0_outputs(1765));
    layer1_outputs(276) <= not(layer0_outputs(3122));
    layer1_outputs(277) <= (layer0_outputs(2711)) and not (layer0_outputs(2328));
    layer1_outputs(278) <= not(layer0_outputs(4726)) or (layer0_outputs(2858));
    layer1_outputs(279) <= not(layer0_outputs(4540));
    layer1_outputs(280) <= (layer0_outputs(3969)) or (layer0_outputs(3529));
    layer1_outputs(281) <= not((layer0_outputs(2322)) and (layer0_outputs(4598)));
    layer1_outputs(282) <= not(layer0_outputs(4460));
    layer1_outputs(283) <= not(layer0_outputs(2167));
    layer1_outputs(284) <= not(layer0_outputs(3041)) or (layer0_outputs(1993));
    layer1_outputs(285) <= '0';
    layer1_outputs(286) <= (layer0_outputs(3864)) xor (layer0_outputs(1730));
    layer1_outputs(287) <= layer0_outputs(62);
    layer1_outputs(288) <= not((layer0_outputs(851)) or (layer0_outputs(4576)));
    layer1_outputs(289) <= not((layer0_outputs(2204)) xor (layer0_outputs(5107)));
    layer1_outputs(290) <= layer0_outputs(459);
    layer1_outputs(291) <= not(layer0_outputs(304));
    layer1_outputs(292) <= (layer0_outputs(3269)) and not (layer0_outputs(4442));
    layer1_outputs(293) <= not((layer0_outputs(1330)) and (layer0_outputs(5074)));
    layer1_outputs(294) <= not(layer0_outputs(4572)) or (layer0_outputs(4489));
    layer1_outputs(295) <= not(layer0_outputs(3600));
    layer1_outputs(296) <= not(layer0_outputs(3979)) or (layer0_outputs(1549));
    layer1_outputs(297) <= not((layer0_outputs(4000)) and (layer0_outputs(3016)));
    layer1_outputs(298) <= (layer0_outputs(4452)) or (layer0_outputs(3825));
    layer1_outputs(299) <= not((layer0_outputs(4354)) or (layer0_outputs(1343)));
    layer1_outputs(300) <= not(layer0_outputs(2308)) or (layer0_outputs(4701));
    layer1_outputs(301) <= (layer0_outputs(3395)) and not (layer0_outputs(3388));
    layer1_outputs(302) <= layer0_outputs(3829);
    layer1_outputs(303) <= (layer0_outputs(1764)) and not (layer0_outputs(3208));
    layer1_outputs(304) <= (layer0_outputs(3778)) xor (layer0_outputs(1472));
    layer1_outputs(305) <= layer0_outputs(887);
    layer1_outputs(306) <= layer0_outputs(1722);
    layer1_outputs(307) <= not(layer0_outputs(1002));
    layer1_outputs(308) <= not((layer0_outputs(1097)) and (layer0_outputs(2838)));
    layer1_outputs(309) <= not(layer0_outputs(410)) or (layer0_outputs(362));
    layer1_outputs(310) <= layer0_outputs(343);
    layer1_outputs(311) <= '0';
    layer1_outputs(312) <= (layer0_outputs(2126)) and not (layer0_outputs(3603));
    layer1_outputs(313) <= '1';
    layer1_outputs(314) <= not(layer0_outputs(2446));
    layer1_outputs(315) <= (layer0_outputs(1548)) or (layer0_outputs(2205));
    layer1_outputs(316) <= not(layer0_outputs(2117)) or (layer0_outputs(1775));
    layer1_outputs(317) <= (layer0_outputs(4144)) and not (layer0_outputs(129));
    layer1_outputs(318) <= not(layer0_outputs(3361)) or (layer0_outputs(2839));
    layer1_outputs(319) <= (layer0_outputs(4946)) and not (layer0_outputs(1718));
    layer1_outputs(320) <= not((layer0_outputs(2441)) and (layer0_outputs(4862)));
    layer1_outputs(321) <= (layer0_outputs(1575)) and (layer0_outputs(665));
    layer1_outputs(322) <= not(layer0_outputs(148));
    layer1_outputs(323) <= (layer0_outputs(500)) or (layer0_outputs(3419));
    layer1_outputs(324) <= layer0_outputs(1142);
    layer1_outputs(325) <= layer0_outputs(353);
    layer1_outputs(326) <= not((layer0_outputs(2568)) and (layer0_outputs(3085)));
    layer1_outputs(327) <= layer0_outputs(4884);
    layer1_outputs(328) <= layer0_outputs(2720);
    layer1_outputs(329) <= layer0_outputs(444);
    layer1_outputs(330) <= not(layer0_outputs(2154));
    layer1_outputs(331) <= (layer0_outputs(4545)) and not (layer0_outputs(2893));
    layer1_outputs(332) <= (layer0_outputs(1046)) or (layer0_outputs(5077));
    layer1_outputs(333) <= layer0_outputs(1171);
    layer1_outputs(334) <= (layer0_outputs(1960)) and not (layer0_outputs(4824));
    layer1_outputs(335) <= not((layer0_outputs(1535)) xor (layer0_outputs(3417)));
    layer1_outputs(336) <= not(layer0_outputs(1766)) or (layer0_outputs(2851));
    layer1_outputs(337) <= '0';
    layer1_outputs(338) <= not(layer0_outputs(4755));
    layer1_outputs(339) <= not(layer0_outputs(1340)) or (layer0_outputs(673));
    layer1_outputs(340) <= layer0_outputs(2929);
    layer1_outputs(341) <= (layer0_outputs(625)) and (layer0_outputs(4748));
    layer1_outputs(342) <= not((layer0_outputs(2856)) and (layer0_outputs(3110)));
    layer1_outputs(343) <= not((layer0_outputs(4327)) and (layer0_outputs(4273)));
    layer1_outputs(344) <= '0';
    layer1_outputs(345) <= not((layer0_outputs(5071)) and (layer0_outputs(2852)));
    layer1_outputs(346) <= not(layer0_outputs(196));
    layer1_outputs(347) <= (layer0_outputs(706)) and (layer0_outputs(2497));
    layer1_outputs(348) <= not((layer0_outputs(3546)) and (layer0_outputs(4196)));
    layer1_outputs(349) <= not(layer0_outputs(942)) or (layer0_outputs(1257));
    layer1_outputs(350) <= layer0_outputs(3283);
    layer1_outputs(351) <= not((layer0_outputs(338)) xor (layer0_outputs(1401)));
    layer1_outputs(352) <= layer0_outputs(2229);
    layer1_outputs(353) <= not(layer0_outputs(4042));
    layer1_outputs(354) <= (layer0_outputs(2750)) and (layer0_outputs(3390));
    layer1_outputs(355) <= not(layer0_outputs(3638));
    layer1_outputs(356) <= (layer0_outputs(3583)) and not (layer0_outputs(471));
    layer1_outputs(357) <= layer0_outputs(1268);
    layer1_outputs(358) <= '0';
    layer1_outputs(359) <= not(layer0_outputs(4662));
    layer1_outputs(360) <= (layer0_outputs(3119)) and not (layer0_outputs(4763));
    layer1_outputs(361) <= not((layer0_outputs(2093)) xor (layer0_outputs(4371)));
    layer1_outputs(362) <= (layer0_outputs(1039)) or (layer0_outputs(1230));
    layer1_outputs(363) <= not(layer0_outputs(1003));
    layer1_outputs(364) <= '1';
    layer1_outputs(365) <= not(layer0_outputs(2227)) or (layer0_outputs(1982));
    layer1_outputs(366) <= '1';
    layer1_outputs(367) <= not(layer0_outputs(3039));
    layer1_outputs(368) <= not((layer0_outputs(1949)) or (layer0_outputs(3423)));
    layer1_outputs(369) <= not((layer0_outputs(1912)) and (layer0_outputs(4940)));
    layer1_outputs(370) <= not(layer0_outputs(3715));
    layer1_outputs(371) <= '1';
    layer1_outputs(372) <= (layer0_outputs(662)) and not (layer0_outputs(3120));
    layer1_outputs(373) <= not((layer0_outputs(4116)) xor (layer0_outputs(2405)));
    layer1_outputs(374) <= (layer0_outputs(4883)) xor (layer0_outputs(2783));
    layer1_outputs(375) <= not(layer0_outputs(1579));
    layer1_outputs(376) <= layer0_outputs(4700);
    layer1_outputs(377) <= layer0_outputs(4508);
    layer1_outputs(378) <= not(layer0_outputs(1703));
    layer1_outputs(379) <= not(layer0_outputs(1015));
    layer1_outputs(380) <= not((layer0_outputs(191)) and (layer0_outputs(4551)));
    layer1_outputs(381) <= not(layer0_outputs(2832)) or (layer0_outputs(5036));
    layer1_outputs(382) <= not((layer0_outputs(4741)) and (layer0_outputs(4736)));
    layer1_outputs(383) <= (layer0_outputs(33)) and not (layer0_outputs(2317));
    layer1_outputs(384) <= not((layer0_outputs(5032)) and (layer0_outputs(2781)));
    layer1_outputs(385) <= (layer0_outputs(1514)) and not (layer0_outputs(4333));
    layer1_outputs(386) <= not(layer0_outputs(1873));
    layer1_outputs(387) <= not(layer0_outputs(1448));
    layer1_outputs(388) <= layer0_outputs(4905);
    layer1_outputs(389) <= (layer0_outputs(4609)) and not (layer0_outputs(4234));
    layer1_outputs(390) <= (layer0_outputs(3091)) and not (layer0_outputs(2659));
    layer1_outputs(391) <= (layer0_outputs(5048)) and not (layer0_outputs(1080));
    layer1_outputs(392) <= not(layer0_outputs(4873)) or (layer0_outputs(1099));
    layer1_outputs(393) <= not(layer0_outputs(3465)) or (layer0_outputs(3611));
    layer1_outputs(394) <= (layer0_outputs(5034)) and not (layer0_outputs(3966));
    layer1_outputs(395) <= not(layer0_outputs(715));
    layer1_outputs(396) <= layer0_outputs(4258);
    layer1_outputs(397) <= layer0_outputs(3849);
    layer1_outputs(398) <= (layer0_outputs(2942)) and not (layer0_outputs(2142));
    layer1_outputs(399) <= not((layer0_outputs(2468)) and (layer0_outputs(3755)));
    layer1_outputs(400) <= (layer0_outputs(993)) xor (layer0_outputs(3296));
    layer1_outputs(401) <= not(layer0_outputs(938)) or (layer0_outputs(1716));
    layer1_outputs(402) <= not((layer0_outputs(2366)) and (layer0_outputs(1369)));
    layer1_outputs(403) <= not(layer0_outputs(3513));
    layer1_outputs(404) <= not((layer0_outputs(3194)) and (layer0_outputs(2710)));
    layer1_outputs(405) <= not(layer0_outputs(289));
    layer1_outputs(406) <= not((layer0_outputs(406)) and (layer0_outputs(1999)));
    layer1_outputs(407) <= (layer0_outputs(3908)) or (layer0_outputs(4418));
    layer1_outputs(408) <= (layer0_outputs(3524)) and not (layer0_outputs(2688));
    layer1_outputs(409) <= layer0_outputs(2524);
    layer1_outputs(410) <= not(layer0_outputs(1973)) or (layer0_outputs(990));
    layer1_outputs(411) <= not((layer0_outputs(1034)) and (layer0_outputs(3882)));
    layer1_outputs(412) <= not(layer0_outputs(5086));
    layer1_outputs(413) <= not(layer0_outputs(111)) or (layer0_outputs(4264));
    layer1_outputs(414) <= not((layer0_outputs(2542)) or (layer0_outputs(208)));
    layer1_outputs(415) <= not(layer0_outputs(3307)) or (layer0_outputs(2992));
    layer1_outputs(416) <= not((layer0_outputs(842)) xor (layer0_outputs(2974)));
    layer1_outputs(417) <= layer0_outputs(2925);
    layer1_outputs(418) <= not(layer0_outputs(4201));
    layer1_outputs(419) <= not(layer0_outputs(2975));
    layer1_outputs(420) <= (layer0_outputs(1207)) or (layer0_outputs(553));
    layer1_outputs(421) <= not(layer0_outputs(636)) or (layer0_outputs(408));
    layer1_outputs(422) <= not(layer0_outputs(2121)) or (layer0_outputs(4719));
    layer1_outputs(423) <= not((layer0_outputs(4077)) and (layer0_outputs(1273)));
    layer1_outputs(424) <= not((layer0_outputs(233)) or (layer0_outputs(2046)));
    layer1_outputs(425) <= not(layer0_outputs(3180));
    layer1_outputs(426) <= not((layer0_outputs(4067)) and (layer0_outputs(3355)));
    layer1_outputs(427) <= '0';
    layer1_outputs(428) <= not((layer0_outputs(2853)) xor (layer0_outputs(705)));
    layer1_outputs(429) <= (layer0_outputs(545)) and not (layer0_outputs(2340));
    layer1_outputs(430) <= not(layer0_outputs(4276));
    layer1_outputs(431) <= (layer0_outputs(4902)) or (layer0_outputs(4364));
    layer1_outputs(432) <= (layer0_outputs(4053)) and not (layer0_outputs(3815));
    layer1_outputs(433) <= not((layer0_outputs(4005)) or (layer0_outputs(3552)));
    layer1_outputs(434) <= not(layer0_outputs(1548));
    layer1_outputs(435) <= not(layer0_outputs(2298));
    layer1_outputs(436) <= layer0_outputs(3807);
    layer1_outputs(437) <= not(layer0_outputs(563)) or (layer0_outputs(3586));
    layer1_outputs(438) <= (layer0_outputs(2061)) xor (layer0_outputs(638));
    layer1_outputs(439) <= not((layer0_outputs(4806)) and (layer0_outputs(2800)));
    layer1_outputs(440) <= (layer0_outputs(1168)) or (layer0_outputs(3917));
    layer1_outputs(441) <= not(layer0_outputs(3542)) or (layer0_outputs(4882));
    layer1_outputs(442) <= not(layer0_outputs(3202));
    layer1_outputs(443) <= layer0_outputs(3195);
    layer1_outputs(444) <= (layer0_outputs(4686)) xor (layer0_outputs(2448));
    layer1_outputs(445) <= not(layer0_outputs(3649));
    layer1_outputs(446) <= layer0_outputs(226);
    layer1_outputs(447) <= layer0_outputs(563);
    layer1_outputs(448) <= not(layer0_outputs(2402));
    layer1_outputs(449) <= layer0_outputs(2517);
    layer1_outputs(450) <= not((layer0_outputs(2556)) xor (layer0_outputs(1962)));
    layer1_outputs(451) <= not(layer0_outputs(1755));
    layer1_outputs(452) <= not(layer0_outputs(4405));
    layer1_outputs(453) <= layer0_outputs(1627);
    layer1_outputs(454) <= (layer0_outputs(4547)) or (layer0_outputs(1541));
    layer1_outputs(455) <= layer0_outputs(1356);
    layer1_outputs(456) <= not((layer0_outputs(273)) or (layer0_outputs(1313)));
    layer1_outputs(457) <= layer0_outputs(3718);
    layer1_outputs(458) <= not(layer0_outputs(3020));
    layer1_outputs(459) <= not((layer0_outputs(3204)) xor (layer0_outputs(3995)));
    layer1_outputs(460) <= not(layer0_outputs(1690));
    layer1_outputs(461) <= '1';
    layer1_outputs(462) <= not((layer0_outputs(3962)) or (layer0_outputs(3997)));
    layer1_outputs(463) <= layer0_outputs(1933);
    layer1_outputs(464) <= (layer0_outputs(1456)) xor (layer0_outputs(1994));
    layer1_outputs(465) <= not(layer0_outputs(464)) or (layer0_outputs(3686));
    layer1_outputs(466) <= layer0_outputs(262);
    layer1_outputs(467) <= not(layer0_outputs(3942)) or (layer0_outputs(466));
    layer1_outputs(468) <= (layer0_outputs(3002)) and (layer0_outputs(2717));
    layer1_outputs(469) <= not(layer0_outputs(3363));
    layer1_outputs(470) <= not(layer0_outputs(5062));
    layer1_outputs(471) <= not((layer0_outputs(888)) and (layer0_outputs(1190)));
    layer1_outputs(472) <= not((layer0_outputs(114)) xor (layer0_outputs(1507)));
    layer1_outputs(473) <= layer0_outputs(1783);
    layer1_outputs(474) <= not(layer0_outputs(2570)) or (layer0_outputs(441));
    layer1_outputs(475) <= (layer0_outputs(655)) xor (layer0_outputs(3930));
    layer1_outputs(476) <= (layer0_outputs(3048)) and (layer0_outputs(2463));
    layer1_outputs(477) <= (layer0_outputs(731)) and not (layer0_outputs(3896));
    layer1_outputs(478) <= (layer0_outputs(1520)) xor (layer0_outputs(3067));
    layer1_outputs(479) <= layer0_outputs(282);
    layer1_outputs(480) <= layer0_outputs(361);
    layer1_outputs(481) <= not((layer0_outputs(4785)) xor (layer0_outputs(3816)));
    layer1_outputs(482) <= layer0_outputs(3047);
    layer1_outputs(483) <= (layer0_outputs(4966)) and not (layer0_outputs(4718));
    layer1_outputs(484) <= not(layer0_outputs(1742));
    layer1_outputs(485) <= (layer0_outputs(139)) or (layer0_outputs(4555));
    layer1_outputs(486) <= layer0_outputs(1796);
    layer1_outputs(487) <= not((layer0_outputs(1019)) or (layer0_outputs(4317)));
    layer1_outputs(488) <= (layer0_outputs(4557)) or (layer0_outputs(3677));
    layer1_outputs(489) <= not((layer0_outputs(1234)) xor (layer0_outputs(1816)));
    layer1_outputs(490) <= not((layer0_outputs(3149)) and (layer0_outputs(1894)));
    layer1_outputs(491) <= layer0_outputs(3420);
    layer1_outputs(492) <= (layer0_outputs(2920)) and not (layer0_outputs(4951));
    layer1_outputs(493) <= not(layer0_outputs(668));
    layer1_outputs(494) <= not((layer0_outputs(3288)) and (layer0_outputs(3736)));
    layer1_outputs(495) <= not(layer0_outputs(4165));
    layer1_outputs(496) <= not((layer0_outputs(975)) or (layer0_outputs(3745)));
    layer1_outputs(497) <= (layer0_outputs(196)) or (layer0_outputs(3102));
    layer1_outputs(498) <= not(layer0_outputs(712));
    layer1_outputs(499) <= (layer0_outputs(4405)) xor (layer0_outputs(4969));
    layer1_outputs(500) <= not((layer0_outputs(3874)) and (layer0_outputs(3683)));
    layer1_outputs(501) <= (layer0_outputs(3950)) and not (layer0_outputs(2466));
    layer1_outputs(502) <= not((layer0_outputs(3961)) or (layer0_outputs(2630)));
    layer1_outputs(503) <= layer0_outputs(1129);
    layer1_outputs(504) <= not((layer0_outputs(1758)) or (layer0_outputs(2515)));
    layer1_outputs(505) <= (layer0_outputs(3858)) and (layer0_outputs(5098));
    layer1_outputs(506) <= (layer0_outputs(107)) or (layer0_outputs(2290));
    layer1_outputs(507) <= not(layer0_outputs(1478));
    layer1_outputs(508) <= not((layer0_outputs(2187)) and (layer0_outputs(2007)));
    layer1_outputs(509) <= not(layer0_outputs(2047));
    layer1_outputs(510) <= '0';
    layer1_outputs(511) <= not((layer0_outputs(173)) or (layer0_outputs(4027)));
    layer1_outputs(512) <= layer0_outputs(1804);
    layer1_outputs(513) <= not((layer0_outputs(4950)) or (layer0_outputs(329)));
    layer1_outputs(514) <= (layer0_outputs(3814)) and not (layer0_outputs(4321));
    layer1_outputs(515) <= (layer0_outputs(2825)) and (layer0_outputs(5065));
    layer1_outputs(516) <= (layer0_outputs(2937)) and not (layer0_outputs(1479));
    layer1_outputs(517) <= (layer0_outputs(4560)) or (layer0_outputs(3593));
    layer1_outputs(518) <= (layer0_outputs(3806)) and not (layer0_outputs(4889));
    layer1_outputs(519) <= (layer0_outputs(253)) or (layer0_outputs(2393));
    layer1_outputs(520) <= not(layer0_outputs(3849));
    layer1_outputs(521) <= (layer0_outputs(1459)) or (layer0_outputs(3577));
    layer1_outputs(522) <= not(layer0_outputs(4114)) or (layer0_outputs(2895));
    layer1_outputs(523) <= layer0_outputs(3015);
    layer1_outputs(524) <= not((layer0_outputs(2337)) and (layer0_outputs(1652)));
    layer1_outputs(525) <= not(layer0_outputs(243)) or (layer0_outputs(4479));
    layer1_outputs(526) <= (layer0_outputs(42)) or (layer0_outputs(4753));
    layer1_outputs(527) <= not(layer0_outputs(2823)) or (layer0_outputs(2814));
    layer1_outputs(528) <= not((layer0_outputs(4298)) and (layer0_outputs(4535)));
    layer1_outputs(529) <= not(layer0_outputs(752)) or (layer0_outputs(1767));
    layer1_outputs(530) <= '0';
    layer1_outputs(531) <= layer0_outputs(3151);
    layer1_outputs(532) <= '0';
    layer1_outputs(533) <= '0';
    layer1_outputs(534) <= not((layer0_outputs(3464)) or (layer0_outputs(1339)));
    layer1_outputs(535) <= not(layer0_outputs(3945)) or (layer0_outputs(3726));
    layer1_outputs(536) <= not((layer0_outputs(641)) xor (layer0_outputs(3460)));
    layer1_outputs(537) <= (layer0_outputs(1514)) xor (layer0_outputs(4123));
    layer1_outputs(538) <= not(layer0_outputs(4561)) or (layer0_outputs(614));
    layer1_outputs(539) <= (layer0_outputs(2966)) xor (layer0_outputs(4620));
    layer1_outputs(540) <= layer0_outputs(266);
    layer1_outputs(541) <= not((layer0_outputs(1871)) or (layer0_outputs(496)));
    layer1_outputs(542) <= not(layer0_outputs(2115)) or (layer0_outputs(2704));
    layer1_outputs(543) <= not(layer0_outputs(2134)) or (layer0_outputs(3143));
    layer1_outputs(544) <= not(layer0_outputs(2055)) or (layer0_outputs(3422));
    layer1_outputs(545) <= (layer0_outputs(61)) and not (layer0_outputs(2746));
    layer1_outputs(546) <= not((layer0_outputs(4828)) xor (layer0_outputs(4034)));
    layer1_outputs(547) <= (layer0_outputs(2860)) xor (layer0_outputs(3219));
    layer1_outputs(548) <= layer0_outputs(152);
    layer1_outputs(549) <= '0';
    layer1_outputs(550) <= (layer0_outputs(873)) and not (layer0_outputs(75));
    layer1_outputs(551) <= (layer0_outputs(4215)) and not (layer0_outputs(3545));
    layer1_outputs(552) <= (layer0_outputs(1353)) and (layer0_outputs(4411));
    layer1_outputs(553) <= layer0_outputs(3085);
    layer1_outputs(554) <= not((layer0_outputs(1589)) or (layer0_outputs(3926)));
    layer1_outputs(555) <= (layer0_outputs(1947)) and not (layer0_outputs(3354));
    layer1_outputs(556) <= not(layer0_outputs(2459)) or (layer0_outputs(1761));
    layer1_outputs(557) <= not((layer0_outputs(4734)) and (layer0_outputs(390)));
    layer1_outputs(558) <= not(layer0_outputs(3238));
    layer1_outputs(559) <= not(layer0_outputs(4337)) or (layer0_outputs(475));
    layer1_outputs(560) <= layer0_outputs(2822);
    layer1_outputs(561) <= (layer0_outputs(4908)) and not (layer0_outputs(4307));
    layer1_outputs(562) <= not((layer0_outputs(2304)) xor (layer0_outputs(4412)));
    layer1_outputs(563) <= (layer0_outputs(4480)) and (layer0_outputs(599));
    layer1_outputs(564) <= not(layer0_outputs(3936)) or (layer0_outputs(3211));
    layer1_outputs(565) <= not(layer0_outputs(3506)) or (layer0_outputs(4217));
    layer1_outputs(566) <= not(layer0_outputs(3751));
    layer1_outputs(567) <= (layer0_outputs(351)) and (layer0_outputs(2816));
    layer1_outputs(568) <= not(layer0_outputs(3858));
    layer1_outputs(569) <= (layer0_outputs(4957)) and not (layer0_outputs(4453));
    layer1_outputs(570) <= layer0_outputs(1085);
    layer1_outputs(571) <= layer0_outputs(902);
    layer1_outputs(572) <= not((layer0_outputs(5088)) xor (layer0_outputs(4084)));
    layer1_outputs(573) <= layer0_outputs(4038);
    layer1_outputs(574) <= layer0_outputs(3149);
    layer1_outputs(575) <= not(layer0_outputs(4765));
    layer1_outputs(576) <= not((layer0_outputs(3706)) or (layer0_outputs(4011)));
    layer1_outputs(577) <= (layer0_outputs(359)) and (layer0_outputs(964));
    layer1_outputs(578) <= not((layer0_outputs(1058)) xor (layer0_outputs(1624)));
    layer1_outputs(579) <= not((layer0_outputs(4532)) and (layer0_outputs(1768)));
    layer1_outputs(580) <= (layer0_outputs(3677)) xor (layer0_outputs(1672));
    layer1_outputs(581) <= layer0_outputs(3305);
    layer1_outputs(582) <= not((layer0_outputs(989)) and (layer0_outputs(484)));
    layer1_outputs(583) <= (layer0_outputs(362)) or (layer0_outputs(2275));
    layer1_outputs(584) <= (layer0_outputs(610)) and (layer0_outputs(3379));
    layer1_outputs(585) <= layer0_outputs(3469);
    layer1_outputs(586) <= '1';
    layer1_outputs(587) <= layer0_outputs(5059);
    layer1_outputs(588) <= not(layer0_outputs(775)) or (layer0_outputs(2708));
    layer1_outputs(589) <= layer0_outputs(1080);
    layer1_outputs(590) <= layer0_outputs(2216);
    layer1_outputs(591) <= not((layer0_outputs(1468)) xor (layer0_outputs(3714)));
    layer1_outputs(592) <= not(layer0_outputs(1888)) or (layer0_outputs(4149));
    layer1_outputs(593) <= (layer0_outputs(2303)) and not (layer0_outputs(1590));
    layer1_outputs(594) <= (layer0_outputs(5019)) xor (layer0_outputs(4347));
    layer1_outputs(595) <= (layer0_outputs(2592)) and (layer0_outputs(780));
    layer1_outputs(596) <= layer0_outputs(4239);
    layer1_outputs(597) <= '0';
    layer1_outputs(598) <= not((layer0_outputs(3608)) and (layer0_outputs(2393)));
    layer1_outputs(599) <= (layer0_outputs(3834)) and not (layer0_outputs(4068));
    layer1_outputs(600) <= not((layer0_outputs(2101)) xor (layer0_outputs(1828)));
    layer1_outputs(601) <= not(layer0_outputs(354));
    layer1_outputs(602) <= not((layer0_outputs(1709)) and (layer0_outputs(295)));
    layer1_outputs(603) <= not(layer0_outputs(44));
    layer1_outputs(604) <= not(layer0_outputs(4959)) or (layer0_outputs(2361));
    layer1_outputs(605) <= not(layer0_outputs(4963)) or (layer0_outputs(1113));
    layer1_outputs(606) <= not((layer0_outputs(674)) and (layer0_outputs(3663)));
    layer1_outputs(607) <= not(layer0_outputs(2921));
    layer1_outputs(608) <= not(layer0_outputs(4605));
    layer1_outputs(609) <= layer0_outputs(4696);
    layer1_outputs(610) <= layer0_outputs(3857);
    layer1_outputs(611) <= not(layer0_outputs(1197));
    layer1_outputs(612) <= not(layer0_outputs(403)) or (layer0_outputs(2017));
    layer1_outputs(613) <= (layer0_outputs(4618)) or (layer0_outputs(1010));
    layer1_outputs(614) <= '0';
    layer1_outputs(615) <= not((layer0_outputs(4921)) or (layer0_outputs(2076)));
    layer1_outputs(616) <= '1';
    layer1_outputs(617) <= layer0_outputs(3762);
    layer1_outputs(618) <= layer0_outputs(1266);
    layer1_outputs(619) <= not(layer0_outputs(452));
    layer1_outputs(620) <= (layer0_outputs(161)) and not (layer0_outputs(2533));
    layer1_outputs(621) <= layer0_outputs(834);
    layer1_outputs(622) <= (layer0_outputs(399)) and not (layer0_outputs(3193));
    layer1_outputs(623) <= (layer0_outputs(4648)) and not (layer0_outputs(3399));
    layer1_outputs(624) <= (layer0_outputs(3776)) and (layer0_outputs(5096));
    layer1_outputs(625) <= (layer0_outputs(651)) and (layer0_outputs(3888));
    layer1_outputs(626) <= not(layer0_outputs(953));
    layer1_outputs(627) <= layer0_outputs(2639);
    layer1_outputs(628) <= (layer0_outputs(4716)) and (layer0_outputs(2622));
    layer1_outputs(629) <= (layer0_outputs(3518)) or (layer0_outputs(5065));
    layer1_outputs(630) <= layer0_outputs(4871);
    layer1_outputs(631) <= not((layer0_outputs(4039)) or (layer0_outputs(1308)));
    layer1_outputs(632) <= (layer0_outputs(158)) and not (layer0_outputs(2081));
    layer1_outputs(633) <= (layer0_outputs(5080)) and (layer0_outputs(1693));
    layer1_outputs(634) <= not(layer0_outputs(4835));
    layer1_outputs(635) <= not(layer0_outputs(973));
    layer1_outputs(636) <= not(layer0_outputs(2032));
    layer1_outputs(637) <= not((layer0_outputs(3217)) and (layer0_outputs(4451)));
    layer1_outputs(638) <= layer0_outputs(3461);
    layer1_outputs(639) <= layer0_outputs(1879);
    layer1_outputs(640) <= not(layer0_outputs(2914));
    layer1_outputs(641) <= (layer0_outputs(2487)) and (layer0_outputs(3055));
    layer1_outputs(642) <= layer0_outputs(1077);
    layer1_outputs(643) <= layer0_outputs(4954);
    layer1_outputs(644) <= not(layer0_outputs(1247));
    layer1_outputs(645) <= (layer0_outputs(2112)) and (layer0_outputs(5014));
    layer1_outputs(646) <= not(layer0_outputs(4356));
    layer1_outputs(647) <= layer0_outputs(4376);
    layer1_outputs(648) <= not((layer0_outputs(1986)) xor (layer0_outputs(4668)));
    layer1_outputs(649) <= '0';
    layer1_outputs(650) <= not((layer0_outputs(4246)) xor (layer0_outputs(2881)));
    layer1_outputs(651) <= '1';
    layer1_outputs(652) <= (layer0_outputs(628)) and (layer0_outputs(84));
    layer1_outputs(653) <= not((layer0_outputs(484)) or (layer0_outputs(2808)));
    layer1_outputs(654) <= layer0_outputs(2881);
    layer1_outputs(655) <= layer0_outputs(2874);
    layer1_outputs(656) <= not(layer0_outputs(4990)) or (layer0_outputs(1060));
    layer1_outputs(657) <= (layer0_outputs(3641)) and (layer0_outputs(4847));
    layer1_outputs(658) <= (layer0_outputs(1565)) xor (layer0_outputs(4239));
    layer1_outputs(659) <= not((layer0_outputs(770)) and (layer0_outputs(1598)));
    layer1_outputs(660) <= not(layer0_outputs(4151)) or (layer0_outputs(1774));
    layer1_outputs(661) <= not((layer0_outputs(4320)) xor (layer0_outputs(5089)));
    layer1_outputs(662) <= not((layer0_outputs(2695)) xor (layer0_outputs(4065)));
    layer1_outputs(663) <= (layer0_outputs(994)) or (layer0_outputs(2235));
    layer1_outputs(664) <= '1';
    layer1_outputs(665) <= layer0_outputs(2626);
    layer1_outputs(666) <= layer0_outputs(4982);
    layer1_outputs(667) <= (layer0_outputs(1494)) and not (layer0_outputs(2147));
    layer1_outputs(668) <= (layer0_outputs(386)) and not (layer0_outputs(1684));
    layer1_outputs(669) <= not((layer0_outputs(781)) xor (layer0_outputs(275)));
    layer1_outputs(670) <= not(layer0_outputs(1552)) or (layer0_outputs(4933));
    layer1_outputs(671) <= not((layer0_outputs(2515)) and (layer0_outputs(4093)));
    layer1_outputs(672) <= (layer0_outputs(2408)) or (layer0_outputs(3223));
    layer1_outputs(673) <= not(layer0_outputs(2981));
    layer1_outputs(674) <= not(layer0_outputs(3001));
    layer1_outputs(675) <= not(layer0_outputs(3702)) or (layer0_outputs(1984));
    layer1_outputs(676) <= not((layer0_outputs(1505)) or (layer0_outputs(555)));
    layer1_outputs(677) <= layer0_outputs(1367);
    layer1_outputs(678) <= '0';
    layer1_outputs(679) <= not((layer0_outputs(2727)) xor (layer0_outputs(3239)));
    layer1_outputs(680) <= (layer0_outputs(787)) and not (layer0_outputs(2995));
    layer1_outputs(681) <= (layer0_outputs(519)) xor (layer0_outputs(5006));
    layer1_outputs(682) <= (layer0_outputs(608)) and not (layer0_outputs(4014));
    layer1_outputs(683) <= not(layer0_outputs(1458));
    layer1_outputs(684) <= '1';
    layer1_outputs(685) <= (layer0_outputs(1921)) and (layer0_outputs(17));
    layer1_outputs(686) <= layer0_outputs(2089);
    layer1_outputs(687) <= not(layer0_outputs(1866));
    layer1_outputs(688) <= not(layer0_outputs(4090));
    layer1_outputs(689) <= not(layer0_outputs(2054));
    layer1_outputs(690) <= not((layer0_outputs(4768)) and (layer0_outputs(1406)));
    layer1_outputs(691) <= '0';
    layer1_outputs(692) <= not(layer0_outputs(2332));
    layer1_outputs(693) <= (layer0_outputs(4909)) and not (layer0_outputs(515));
    layer1_outputs(694) <= not(layer0_outputs(3374)) or (layer0_outputs(840));
    layer1_outputs(695) <= not((layer0_outputs(1633)) xor (layer0_outputs(79)));
    layer1_outputs(696) <= '1';
    layer1_outputs(697) <= not(layer0_outputs(4837));
    layer1_outputs(698) <= (layer0_outputs(449)) and not (layer0_outputs(3747));
    layer1_outputs(699) <= (layer0_outputs(4873)) and not (layer0_outputs(3132));
    layer1_outputs(700) <= layer0_outputs(4007);
    layer1_outputs(701) <= not((layer0_outputs(907)) and (layer0_outputs(2732)));
    layer1_outputs(702) <= (layer0_outputs(1339)) and (layer0_outputs(3282));
    layer1_outputs(703) <= layer0_outputs(3979);
    layer1_outputs(704) <= layer0_outputs(4156);
    layer1_outputs(705) <= not(layer0_outputs(1780));
    layer1_outputs(706) <= (layer0_outputs(2409)) and not (layer0_outputs(3002));
    layer1_outputs(707) <= not(layer0_outputs(3273));
    layer1_outputs(708) <= not((layer0_outputs(3230)) xor (layer0_outputs(617)));
    layer1_outputs(709) <= layer0_outputs(679);
    layer1_outputs(710) <= not(layer0_outputs(142));
    layer1_outputs(711) <= not(layer0_outputs(4972));
    layer1_outputs(712) <= not((layer0_outputs(1398)) or (layer0_outputs(3681)));
    layer1_outputs(713) <= (layer0_outputs(104)) xor (layer0_outputs(868));
    layer1_outputs(714) <= (layer0_outputs(3929)) and (layer0_outputs(4731));
    layer1_outputs(715) <= layer0_outputs(546);
    layer1_outputs(716) <= layer0_outputs(2787);
    layer1_outputs(717) <= (layer0_outputs(745)) and not (layer0_outputs(4630));
    layer1_outputs(718) <= layer0_outputs(4272);
    layer1_outputs(719) <= layer0_outputs(1900);
    layer1_outputs(720) <= not(layer0_outputs(2078));
    layer1_outputs(721) <= not(layer0_outputs(1890)) or (layer0_outputs(901));
    layer1_outputs(722) <= (layer0_outputs(4343)) and not (layer0_outputs(3802));
    layer1_outputs(723) <= not((layer0_outputs(1417)) or (layer0_outputs(5039)));
    layer1_outputs(724) <= not((layer0_outputs(4026)) and (layer0_outputs(3771)));
    layer1_outputs(725) <= not((layer0_outputs(4428)) or (layer0_outputs(1629)));
    layer1_outputs(726) <= not(layer0_outputs(2428)) or (layer0_outputs(1601));
    layer1_outputs(727) <= not(layer0_outputs(3626));
    layer1_outputs(728) <= not(layer0_outputs(1215)) or (layer0_outputs(2734));
    layer1_outputs(729) <= not(layer0_outputs(1623)) or (layer0_outputs(4391));
    layer1_outputs(730) <= (layer0_outputs(1960)) and not (layer0_outputs(3410));
    layer1_outputs(731) <= not(layer0_outputs(3710));
    layer1_outputs(732) <= (layer0_outputs(3501)) and (layer0_outputs(4808));
    layer1_outputs(733) <= layer0_outputs(2976);
    layer1_outputs(734) <= not(layer0_outputs(3411));
    layer1_outputs(735) <= layer0_outputs(2256);
    layer1_outputs(736) <= not(layer0_outputs(2518)) or (layer0_outputs(3732));
    layer1_outputs(737) <= not(layer0_outputs(1100));
    layer1_outputs(738) <= not((layer0_outputs(2072)) and (layer0_outputs(2286)));
    layer1_outputs(739) <= (layer0_outputs(86)) and not (layer0_outputs(813));
    layer1_outputs(740) <= not((layer0_outputs(954)) or (layer0_outputs(1585)));
    layer1_outputs(741) <= not((layer0_outputs(4018)) and (layer0_outputs(2088)));
    layer1_outputs(742) <= '0';
    layer1_outputs(743) <= layer0_outputs(3148);
    layer1_outputs(744) <= not(layer0_outputs(1894)) or (layer0_outputs(3700));
    layer1_outputs(745) <= (layer0_outputs(3949)) or (layer0_outputs(382));
    layer1_outputs(746) <= (layer0_outputs(3653)) xor (layer0_outputs(652));
    layer1_outputs(747) <= not(layer0_outputs(4774)) or (layer0_outputs(3685));
    layer1_outputs(748) <= (layer0_outputs(3109)) xor (layer0_outputs(632));
    layer1_outputs(749) <= layer0_outputs(263);
    layer1_outputs(750) <= (layer0_outputs(2712)) xor (layer0_outputs(3289));
    layer1_outputs(751) <= not(layer0_outputs(4986)) or (layer0_outputs(240));
    layer1_outputs(752) <= not(layer0_outputs(4674));
    layer1_outputs(753) <= not((layer0_outputs(3708)) xor (layer0_outputs(4600)));
    layer1_outputs(754) <= layer0_outputs(2552);
    layer1_outputs(755) <= (layer0_outputs(3425)) and not (layer0_outputs(3131));
    layer1_outputs(756) <= '0';
    layer1_outputs(757) <= '1';
    layer1_outputs(758) <= '0';
    layer1_outputs(759) <= not((layer0_outputs(1031)) or (layer0_outputs(910)));
    layer1_outputs(760) <= (layer0_outputs(3537)) and (layer0_outputs(4069));
    layer1_outputs(761) <= '1';
    layer1_outputs(762) <= not(layer0_outputs(558));
    layer1_outputs(763) <= (layer0_outputs(4657)) and (layer0_outputs(2459));
    layer1_outputs(764) <= layer0_outputs(3949);
    layer1_outputs(765) <= not((layer0_outputs(526)) or (layer0_outputs(2936)));
    layer1_outputs(766) <= not(layer0_outputs(2790)) or (layer0_outputs(4845));
    layer1_outputs(767) <= not((layer0_outputs(5070)) and (layer0_outputs(2886)));
    layer1_outputs(768) <= '0';
    layer1_outputs(769) <= (layer0_outputs(4202)) and (layer0_outputs(4642));
    layer1_outputs(770) <= (layer0_outputs(945)) xor (layer0_outputs(20));
    layer1_outputs(771) <= (layer0_outputs(1656)) and (layer0_outputs(1785));
    layer1_outputs(772) <= not((layer0_outputs(448)) or (layer0_outputs(4289)));
    layer1_outputs(773) <= (layer0_outputs(2883)) and (layer0_outputs(1711));
    layer1_outputs(774) <= not((layer0_outputs(4107)) or (layer0_outputs(4230)));
    layer1_outputs(775) <= (layer0_outputs(2635)) or (layer0_outputs(370));
    layer1_outputs(776) <= not(layer0_outputs(900)) or (layer0_outputs(1397));
    layer1_outputs(777) <= (layer0_outputs(4253)) or (layer0_outputs(4796));
    layer1_outputs(778) <= (layer0_outputs(2139)) xor (layer0_outputs(719));
    layer1_outputs(779) <= layer0_outputs(2967);
    layer1_outputs(780) <= (layer0_outputs(1897)) and not (layer0_outputs(3673));
    layer1_outputs(781) <= (layer0_outputs(3433)) or (layer0_outputs(3252));
    layer1_outputs(782) <= (layer0_outputs(4222)) and (layer0_outputs(3973));
    layer1_outputs(783) <= (layer0_outputs(1363)) and (layer0_outputs(1085));
    layer1_outputs(784) <= layer0_outputs(3304);
    layer1_outputs(785) <= not(layer0_outputs(4900));
    layer1_outputs(786) <= (layer0_outputs(3672)) or (layer0_outputs(479));
    layer1_outputs(787) <= not(layer0_outputs(4680)) or (layer0_outputs(3935));
    layer1_outputs(788) <= layer0_outputs(4952);
    layer1_outputs(789) <= not(layer0_outputs(53)) or (layer0_outputs(4747));
    layer1_outputs(790) <= (layer0_outputs(4621)) and (layer0_outputs(2697));
    layer1_outputs(791) <= not(layer0_outputs(2440)) or (layer0_outputs(1502));
    layer1_outputs(792) <= (layer0_outputs(4500)) and (layer0_outputs(2395));
    layer1_outputs(793) <= layer0_outputs(48);
    layer1_outputs(794) <= layer0_outputs(1015);
    layer1_outputs(795) <= not(layer0_outputs(447)) or (layer0_outputs(3151));
    layer1_outputs(796) <= layer0_outputs(2476);
    layer1_outputs(797) <= (layer0_outputs(276)) or (layer0_outputs(4318));
    layer1_outputs(798) <= layer0_outputs(1863);
    layer1_outputs(799) <= not(layer0_outputs(4396));
    layer1_outputs(800) <= not(layer0_outputs(3353));
    layer1_outputs(801) <= '1';
    layer1_outputs(802) <= layer0_outputs(4044);
    layer1_outputs(803) <= (layer0_outputs(135)) and not (layer0_outputs(5093));
    layer1_outputs(804) <= not(layer0_outputs(1138));
    layer1_outputs(805) <= (layer0_outputs(2060)) xor (layer0_outputs(527));
    layer1_outputs(806) <= not(layer0_outputs(4974)) or (layer0_outputs(2927));
    layer1_outputs(807) <= layer0_outputs(3357);
    layer1_outputs(808) <= not((layer0_outputs(935)) xor (layer0_outputs(1440)));
    layer1_outputs(809) <= (layer0_outputs(5004)) xor (layer0_outputs(1869));
    layer1_outputs(810) <= layer0_outputs(1729);
    layer1_outputs(811) <= not(layer0_outputs(898)) or (layer0_outputs(3684));
    layer1_outputs(812) <= '0';
    layer1_outputs(813) <= (layer0_outputs(3111)) or (layer0_outputs(5036));
    layer1_outputs(814) <= (layer0_outputs(4855)) and not (layer0_outputs(2803));
    layer1_outputs(815) <= not((layer0_outputs(3021)) and (layer0_outputs(1218)));
    layer1_outputs(816) <= not((layer0_outputs(4248)) xor (layer0_outputs(1087)));
    layer1_outputs(817) <= layer0_outputs(1324);
    layer1_outputs(818) <= layer0_outputs(3444);
    layer1_outputs(819) <= not((layer0_outputs(4237)) or (layer0_outputs(5055)));
    layer1_outputs(820) <= not((layer0_outputs(329)) or (layer0_outputs(3781)));
    layer1_outputs(821) <= layer0_outputs(3216);
    layer1_outputs(822) <= not(layer0_outputs(1527)) or (layer0_outputs(4153));
    layer1_outputs(823) <= (layer0_outputs(4110)) or (layer0_outputs(1946));
    layer1_outputs(824) <= not(layer0_outputs(921)) or (layer0_outputs(125));
    layer1_outputs(825) <= not((layer0_outputs(4388)) or (layer0_outputs(3017)));
    layer1_outputs(826) <= not((layer0_outputs(2404)) and (layer0_outputs(442)));
    layer1_outputs(827) <= not(layer0_outputs(4530));
    layer1_outputs(828) <= not(layer0_outputs(2090)) or (layer0_outputs(4681));
    layer1_outputs(829) <= not((layer0_outputs(4529)) or (layer0_outputs(637)));
    layer1_outputs(830) <= not(layer0_outputs(1431)) or (layer0_outputs(4988));
    layer1_outputs(831) <= not(layer0_outputs(314));
    layer1_outputs(832) <= not(layer0_outputs(3657));
    layer1_outputs(833) <= not(layer0_outputs(2649)) or (layer0_outputs(3180));
    layer1_outputs(834) <= layer0_outputs(3648);
    layer1_outputs(835) <= not(layer0_outputs(1938));
    layer1_outputs(836) <= layer0_outputs(4615);
    layer1_outputs(837) <= layer0_outputs(426);
    layer1_outputs(838) <= (layer0_outputs(2416)) and not (layer0_outputs(1045));
    layer1_outputs(839) <= not(layer0_outputs(1574));
    layer1_outputs(840) <= not((layer0_outputs(1349)) and (layer0_outputs(336)));
    layer1_outputs(841) <= not((layer0_outputs(372)) xor (layer0_outputs(3391)));
    layer1_outputs(842) <= (layer0_outputs(2985)) and not (layer0_outputs(3873));
    layer1_outputs(843) <= not((layer0_outputs(15)) and (layer0_outputs(162)));
    layer1_outputs(844) <= not(layer0_outputs(3737)) or (layer0_outputs(4654));
    layer1_outputs(845) <= layer0_outputs(1327);
    layer1_outputs(846) <= '0';
    layer1_outputs(847) <= (layer0_outputs(4507)) and not (layer0_outputs(389));
    layer1_outputs(848) <= (layer0_outputs(2470)) and not (layer0_outputs(224));
    layer1_outputs(849) <= not(layer0_outputs(866));
    layer1_outputs(850) <= (layer0_outputs(1725)) and not (layer0_outputs(1602));
    layer1_outputs(851) <= layer0_outputs(1455);
    layer1_outputs(852) <= layer0_outputs(2962);
    layer1_outputs(853) <= (layer0_outputs(4041)) and not (layer0_outputs(1590));
    layer1_outputs(854) <= not(layer0_outputs(1498));
    layer1_outputs(855) <= not((layer0_outputs(3468)) or (layer0_outputs(4512)));
    layer1_outputs(856) <= not(layer0_outputs(1463)) or (layer0_outputs(5003));
    layer1_outputs(857) <= layer0_outputs(1706);
    layer1_outputs(858) <= not(layer0_outputs(3719));
    layer1_outputs(859) <= layer0_outputs(4350);
    layer1_outputs(860) <= not((layer0_outputs(2700)) xor (layer0_outputs(5071)));
    layer1_outputs(861) <= (layer0_outputs(566)) and (layer0_outputs(4281));
    layer1_outputs(862) <= (layer0_outputs(3892)) and not (layer0_outputs(2220));
    layer1_outputs(863) <= layer0_outputs(3743);
    layer1_outputs(864) <= layer0_outputs(2512);
    layer1_outputs(865) <= not(layer0_outputs(1363)) or (layer0_outputs(1353));
    layer1_outputs(866) <= (layer0_outputs(4612)) and not (layer0_outputs(1957));
    layer1_outputs(867) <= not(layer0_outputs(1213));
    layer1_outputs(868) <= layer0_outputs(3875);
    layer1_outputs(869) <= (layer0_outputs(4564)) or (layer0_outputs(4833));
    layer1_outputs(870) <= (layer0_outputs(2118)) xor (layer0_outputs(3018));
    layer1_outputs(871) <= not(layer0_outputs(4907));
    layer1_outputs(872) <= not(layer0_outputs(3314));
    layer1_outputs(873) <= not((layer0_outputs(4397)) xor (layer0_outputs(2903)));
    layer1_outputs(874) <= not((layer0_outputs(4631)) or (layer0_outputs(4187)));
    layer1_outputs(875) <= not(layer0_outputs(3639)) or (layer0_outputs(2861));
    layer1_outputs(876) <= not((layer0_outputs(488)) or (layer0_outputs(1385)));
    layer1_outputs(877) <= layer0_outputs(3242);
    layer1_outputs(878) <= (layer0_outputs(3960)) xor (layer0_outputs(5072));
    layer1_outputs(879) <= not((layer0_outputs(541)) and (layer0_outputs(2419)));
    layer1_outputs(880) <= not(layer0_outputs(370));
    layer1_outputs(881) <= not(layer0_outputs(5049));
    layer1_outputs(882) <= (layer0_outputs(1294)) xor (layer0_outputs(106));
    layer1_outputs(883) <= not((layer0_outputs(2125)) and (layer0_outputs(4015)));
    layer1_outputs(884) <= layer0_outputs(1153);
    layer1_outputs(885) <= not(layer0_outputs(3680));
    layer1_outputs(886) <= not(layer0_outputs(3142));
    layer1_outputs(887) <= (layer0_outputs(435)) and not (layer0_outputs(1792));
    layer1_outputs(888) <= not(layer0_outputs(719));
    layer1_outputs(889) <= (layer0_outputs(1427)) and (layer0_outputs(3569));
    layer1_outputs(890) <= not(layer0_outputs(2878)) or (layer0_outputs(1893));
    layer1_outputs(891) <= (layer0_outputs(3621)) and not (layer0_outputs(779));
    layer1_outputs(892) <= not(layer0_outputs(2429)) or (layer0_outputs(4964));
    layer1_outputs(893) <= (layer0_outputs(520)) and (layer0_outputs(1107));
    layer1_outputs(894) <= (layer0_outputs(2268)) and not (layer0_outputs(2931));
    layer1_outputs(895) <= (layer0_outputs(2663)) or (layer0_outputs(4118));
    layer1_outputs(896) <= (layer0_outputs(4245)) and (layer0_outputs(195));
    layer1_outputs(897) <= not(layer0_outputs(4310)) or (layer0_outputs(3135));
    layer1_outputs(898) <= '0';
    layer1_outputs(899) <= (layer0_outputs(4651)) or (layer0_outputs(455));
    layer1_outputs(900) <= not(layer0_outputs(4779)) or (layer0_outputs(1856));
    layer1_outputs(901) <= not(layer0_outputs(4359));
    layer1_outputs(902) <= not((layer0_outputs(4831)) xor (layer0_outputs(207)));
    layer1_outputs(903) <= layer0_outputs(263);
    layer1_outputs(904) <= layer0_outputs(4242);
    layer1_outputs(905) <= layer0_outputs(1822);
    layer1_outputs(906) <= (layer0_outputs(3731)) or (layer0_outputs(2073));
    layer1_outputs(907) <= not((layer0_outputs(2781)) or (layer0_outputs(562)));
    layer1_outputs(908) <= layer0_outputs(2865);
    layer1_outputs(909) <= (layer0_outputs(802)) and not (layer0_outputs(3157));
    layer1_outputs(910) <= (layer0_outputs(197)) xor (layer0_outputs(3652));
    layer1_outputs(911) <= not((layer0_outputs(3608)) and (layer0_outputs(2562)));
    layer1_outputs(912) <= layer0_outputs(1167);
    layer1_outputs(913) <= layer0_outputs(1126);
    layer1_outputs(914) <= (layer0_outputs(4490)) xor (layer0_outputs(5069));
    layer1_outputs(915) <= not((layer0_outputs(1428)) xor (layer0_outputs(1943)));
    layer1_outputs(916) <= not(layer0_outputs(1556));
    layer1_outputs(917) <= not(layer0_outputs(1237)) or (layer0_outputs(180));
    layer1_outputs(918) <= layer0_outputs(1632);
    layer1_outputs(919) <= layer0_outputs(529);
    layer1_outputs(920) <= (layer0_outputs(3282)) xor (layer0_outputs(4490));
    layer1_outputs(921) <= (layer0_outputs(2802)) and not (layer0_outputs(2539));
    layer1_outputs(922) <= layer0_outputs(466);
    layer1_outputs(923) <= not((layer0_outputs(3101)) xor (layer0_outputs(2360)));
    layer1_outputs(924) <= layer0_outputs(3072);
    layer1_outputs(925) <= (layer0_outputs(3534)) xor (layer0_outputs(2158));
    layer1_outputs(926) <= layer0_outputs(1347);
    layer1_outputs(927) <= (layer0_outputs(1553)) and (layer0_outputs(3538));
    layer1_outputs(928) <= '1';
    layer1_outputs(929) <= (layer0_outputs(4281)) and (layer0_outputs(1289));
    layer1_outputs(930) <= not(layer0_outputs(525));
    layer1_outputs(931) <= (layer0_outputs(2384)) and not (layer0_outputs(2236));
    layer1_outputs(932) <= not((layer0_outputs(3442)) or (layer0_outputs(2046)));
    layer1_outputs(933) <= not(layer0_outputs(2234)) or (layer0_outputs(251));
    layer1_outputs(934) <= '0';
    layer1_outputs(935) <= not((layer0_outputs(269)) and (layer0_outputs(2895)));
    layer1_outputs(936) <= '1';
    layer1_outputs(937) <= not((layer0_outputs(2877)) xor (layer0_outputs(2418)));
    layer1_outputs(938) <= (layer0_outputs(5054)) and not (layer0_outputs(2214));
    layer1_outputs(939) <= not(layer0_outputs(2111));
    layer1_outputs(940) <= (layer0_outputs(1110)) or (layer0_outputs(4528));
    layer1_outputs(941) <= layer0_outputs(2883);
    layer1_outputs(942) <= (layer0_outputs(4783)) xor (layer0_outputs(4899));
    layer1_outputs(943) <= not(layer0_outputs(421));
    layer1_outputs(944) <= layer0_outputs(1704);
    layer1_outputs(945) <= not((layer0_outputs(2792)) or (layer0_outputs(3000)));
    layer1_outputs(946) <= not(layer0_outputs(4782));
    layer1_outputs(947) <= layer0_outputs(3640);
    layer1_outputs(948) <= layer0_outputs(2064);
    layer1_outputs(949) <= layer0_outputs(4431);
    layer1_outputs(950) <= not(layer0_outputs(669)) or (layer0_outputs(3455));
    layer1_outputs(951) <= not((layer0_outputs(2397)) or (layer0_outputs(4784)));
    layer1_outputs(952) <= (layer0_outputs(4632)) and not (layer0_outputs(2940));
    layer1_outputs(953) <= (layer0_outputs(605)) xor (layer0_outputs(1715));
    layer1_outputs(954) <= (layer0_outputs(2512)) xor (layer0_outputs(508));
    layer1_outputs(955) <= (layer0_outputs(1024)) or (layer0_outputs(2938));
    layer1_outputs(956) <= (layer0_outputs(4001)) and (layer0_outputs(2607));
    layer1_outputs(957) <= not(layer0_outputs(1903)) or (layer0_outputs(371));
    layer1_outputs(958) <= not(layer0_outputs(947));
    layer1_outputs(959) <= '0';
    layer1_outputs(960) <= layer0_outputs(916);
    layer1_outputs(961) <= layer0_outputs(4603);
    layer1_outputs(962) <= layer0_outputs(2338);
    layer1_outputs(963) <= not(layer0_outputs(4535));
    layer1_outputs(964) <= layer0_outputs(4101);
    layer1_outputs(965) <= not(layer0_outputs(3642)) or (layer0_outputs(1496));
    layer1_outputs(966) <= (layer0_outputs(4691)) and not (layer0_outputs(1111));
    layer1_outputs(967) <= not(layer0_outputs(4672));
    layer1_outputs(968) <= (layer0_outputs(564)) or (layer0_outputs(3424));
    layer1_outputs(969) <= layer0_outputs(3076);
    layer1_outputs(970) <= layer0_outputs(2773);
    layer1_outputs(971) <= not(layer0_outputs(1837));
    layer1_outputs(972) <= not(layer0_outputs(3669));
    layer1_outputs(973) <= layer0_outputs(2583);
    layer1_outputs(974) <= not((layer0_outputs(717)) and (layer0_outputs(5073)));
    layer1_outputs(975) <= not(layer0_outputs(2990)) or (layer0_outputs(4194));
    layer1_outputs(976) <= (layer0_outputs(773)) xor (layer0_outputs(867));
    layer1_outputs(977) <= not((layer0_outputs(1922)) or (layer0_outputs(1930)));
    layer1_outputs(978) <= layer0_outputs(3950);
    layer1_outputs(979) <= not(layer0_outputs(976));
    layer1_outputs(980) <= not(layer0_outputs(1253));
    layer1_outputs(981) <= (layer0_outputs(2129)) or (layer0_outputs(1304));
    layer1_outputs(982) <= (layer0_outputs(1023)) and not (layer0_outputs(4201));
    layer1_outputs(983) <= (layer0_outputs(1395)) or (layer0_outputs(374));
    layer1_outputs(984) <= (layer0_outputs(52)) xor (layer0_outputs(5010));
    layer1_outputs(985) <= not((layer0_outputs(1473)) xor (layer0_outputs(4663)));
    layer1_outputs(986) <= not((layer0_outputs(854)) and (layer0_outputs(1138)));
    layer1_outputs(987) <= not(layer0_outputs(2412));
    layer1_outputs(988) <= (layer0_outputs(4702)) and not (layer0_outputs(4457));
    layer1_outputs(989) <= not(layer0_outputs(4498)) or (layer0_outputs(1320));
    layer1_outputs(990) <= (layer0_outputs(3883)) and not (layer0_outputs(11));
    layer1_outputs(991) <= (layer0_outputs(4415)) and (layer0_outputs(173));
    layer1_outputs(992) <= '0';
    layer1_outputs(993) <= not((layer0_outputs(4910)) and (layer0_outputs(86)));
    layer1_outputs(994) <= (layer0_outputs(322)) and (layer0_outputs(4466));
    layer1_outputs(995) <= not((layer0_outputs(3171)) xor (layer0_outputs(4733)));
    layer1_outputs(996) <= not((layer0_outputs(3154)) xor (layer0_outputs(508)));
    layer1_outputs(997) <= layer0_outputs(5001);
    layer1_outputs(998) <= (layer0_outputs(48)) and not (layer0_outputs(3870));
    layer1_outputs(999) <= not(layer0_outputs(600));
    layer1_outputs(1000) <= (layer0_outputs(4509)) and not (layer0_outputs(3672));
    layer1_outputs(1001) <= not(layer0_outputs(2980));
    layer1_outputs(1002) <= (layer0_outputs(5015)) and not (layer0_outputs(2667));
    layer1_outputs(1003) <= not(layer0_outputs(1296));
    layer1_outputs(1004) <= not(layer0_outputs(4028));
    layer1_outputs(1005) <= '0';
    layer1_outputs(1006) <= (layer0_outputs(2589)) and not (layer0_outputs(4754));
    layer1_outputs(1007) <= (layer0_outputs(2050)) or (layer0_outputs(101));
    layer1_outputs(1008) <= not(layer0_outputs(2542)) or (layer0_outputs(1405));
    layer1_outputs(1009) <= (layer0_outputs(1593)) xor (layer0_outputs(594));
    layer1_outputs(1010) <= (layer0_outputs(3341)) or (layer0_outputs(5053));
    layer1_outputs(1011) <= (layer0_outputs(3597)) and (layer0_outputs(4952));
    layer1_outputs(1012) <= not((layer0_outputs(2963)) and (layer0_outputs(4255)));
    layer1_outputs(1013) <= not(layer0_outputs(155));
    layer1_outputs(1014) <= not((layer0_outputs(4331)) and (layer0_outputs(1625)));
    layer1_outputs(1015) <= (layer0_outputs(2999)) xor (layer0_outputs(929));
    layer1_outputs(1016) <= not(layer0_outputs(4760)) or (layer0_outputs(2428));
    layer1_outputs(1017) <= layer0_outputs(346);
    layer1_outputs(1018) <= not(layer0_outputs(909));
    layer1_outputs(1019) <= layer0_outputs(4632);
    layer1_outputs(1020) <= '0';
    layer1_outputs(1021) <= not((layer0_outputs(4794)) or (layer0_outputs(706)));
    layer1_outputs(1022) <= not(layer0_outputs(1431)) or (layer0_outputs(4180));
    layer1_outputs(1023) <= not(layer0_outputs(1227));
    layer1_outputs(1024) <= layer0_outputs(2067);
    layer1_outputs(1025) <= (layer0_outputs(4216)) and not (layer0_outputs(2640));
    layer1_outputs(1026) <= not(layer0_outputs(3421)) or (layer0_outputs(4437));
    layer1_outputs(1027) <= (layer0_outputs(4748)) and not (layer0_outputs(1000));
    layer1_outputs(1028) <= (layer0_outputs(4009)) and not (layer0_outputs(1209));
    layer1_outputs(1029) <= not(layer0_outputs(2715));
    layer1_outputs(1030) <= layer0_outputs(486);
    layer1_outputs(1031) <= not(layer0_outputs(4492));
    layer1_outputs(1032) <= (layer0_outputs(2453)) or (layer0_outputs(1678));
    layer1_outputs(1033) <= (layer0_outputs(4991)) and not (layer0_outputs(4646));
    layer1_outputs(1034) <= (layer0_outputs(3077)) and not (layer0_outputs(3413));
    layer1_outputs(1035) <= not(layer0_outputs(917));
    layer1_outputs(1036) <= '1';
    layer1_outputs(1037) <= not(layer0_outputs(1365)) or (layer0_outputs(1061));
    layer1_outputs(1038) <= (layer0_outputs(3087)) or (layer0_outputs(3057));
    layer1_outputs(1039) <= not((layer0_outputs(34)) xor (layer0_outputs(384)));
    layer1_outputs(1040) <= not(layer0_outputs(2832));
    layer1_outputs(1041) <= not((layer0_outputs(769)) and (layer0_outputs(4973)));
    layer1_outputs(1042) <= layer0_outputs(3088);
    layer1_outputs(1043) <= layer0_outputs(4816);
    layer1_outputs(1044) <= (layer0_outputs(784)) and not (layer0_outputs(1112));
    layer1_outputs(1045) <= layer0_outputs(5064);
    layer1_outputs(1046) <= layer0_outputs(4431);
    layer1_outputs(1047) <= not(layer0_outputs(4917)) or (layer0_outputs(2697));
    layer1_outputs(1048) <= not((layer0_outputs(4158)) xor (layer0_outputs(4063)));
    layer1_outputs(1049) <= (layer0_outputs(725)) xor (layer0_outputs(394));
    layer1_outputs(1050) <= not(layer0_outputs(1643));
    layer1_outputs(1051) <= not(layer0_outputs(3309));
    layer1_outputs(1052) <= (layer0_outputs(2536)) and not (layer0_outputs(1819));
    layer1_outputs(1053) <= not(layer0_outputs(259)) or (layer0_outputs(888));
    layer1_outputs(1054) <= not(layer0_outputs(341));
    layer1_outputs(1055) <= (layer0_outputs(1534)) and (layer0_outputs(1276));
    layer1_outputs(1056) <= not(layer0_outputs(1020));
    layer1_outputs(1057) <= layer0_outputs(2104);
    layer1_outputs(1058) <= not((layer0_outputs(3516)) or (layer0_outputs(846)));
    layer1_outputs(1059) <= (layer0_outputs(4932)) xor (layer0_outputs(2122));
    layer1_outputs(1060) <= not(layer0_outputs(1546));
    layer1_outputs(1061) <= not(layer0_outputs(2690));
    layer1_outputs(1062) <= not(layer0_outputs(3836));
    layer1_outputs(1063) <= layer0_outputs(883);
    layer1_outputs(1064) <= not(layer0_outputs(1838)) or (layer0_outputs(3682));
    layer1_outputs(1065) <= not(layer0_outputs(4647)) or (layer0_outputs(1166));
    layer1_outputs(1066) <= not((layer0_outputs(3853)) and (layer0_outputs(2287)));
    layer1_outputs(1067) <= (layer0_outputs(949)) xor (layer0_outputs(3769));
    layer1_outputs(1068) <= layer0_outputs(3666);
    layer1_outputs(1069) <= not(layer0_outputs(751));
    layer1_outputs(1070) <= (layer0_outputs(3078)) xor (layer0_outputs(1082));
    layer1_outputs(1071) <= not((layer0_outputs(2474)) or (layer0_outputs(4788)));
    layer1_outputs(1072) <= layer0_outputs(2259);
    layer1_outputs(1073) <= not((layer0_outputs(1821)) or (layer0_outputs(3735)));
    layer1_outputs(1074) <= (layer0_outputs(1523)) and not (layer0_outputs(3494));
    layer1_outputs(1075) <= not(layer0_outputs(2627)) or (layer0_outputs(1884));
    layer1_outputs(1076) <= (layer0_outputs(2271)) and (layer0_outputs(3599));
    layer1_outputs(1077) <= not(layer0_outputs(957));
    layer1_outputs(1078) <= not((layer0_outputs(3393)) or (layer0_outputs(2175)));
    layer1_outputs(1079) <= not(layer0_outputs(4036)) or (layer0_outputs(3017));
    layer1_outputs(1080) <= '1';
    layer1_outputs(1081) <= not((layer0_outputs(2567)) or (layer0_outputs(366)));
    layer1_outputs(1082) <= not((layer0_outputs(1303)) or (layer0_outputs(1486)));
    layer1_outputs(1083) <= not(layer0_outputs(3412));
    layer1_outputs(1084) <= layer0_outputs(4665);
    layer1_outputs(1085) <= layer0_outputs(3418);
    layer1_outputs(1086) <= not(layer0_outputs(4772)) or (layer0_outputs(3377));
    layer1_outputs(1087) <= (layer0_outputs(1178)) and not (layer0_outputs(2149));
    layer1_outputs(1088) <= not((layer0_outputs(718)) or (layer0_outputs(4663)));
    layer1_outputs(1089) <= (layer0_outputs(2462)) or (layer0_outputs(5068));
    layer1_outputs(1090) <= not((layer0_outputs(4372)) or (layer0_outputs(1759)));
    layer1_outputs(1091) <= not((layer0_outputs(1090)) xor (layer0_outputs(773)));
    layer1_outputs(1092) <= not(layer0_outputs(363));
    layer1_outputs(1093) <= (layer0_outputs(1801)) and not (layer0_outputs(360));
    layer1_outputs(1094) <= not((layer0_outputs(623)) or (layer0_outputs(552)));
    layer1_outputs(1095) <= (layer0_outputs(683)) or (layer0_outputs(2751));
    layer1_outputs(1096) <= not(layer0_outputs(1250));
    layer1_outputs(1097) <= (layer0_outputs(3774)) and not (layer0_outputs(962));
    layer1_outputs(1098) <= not(layer0_outputs(562));
    layer1_outputs(1099) <= not((layer0_outputs(1578)) xor (layer0_outputs(312)));
    layer1_outputs(1100) <= not(layer0_outputs(3924));
    layer1_outputs(1101) <= (layer0_outputs(354)) xor (layer0_outputs(4077));
    layer1_outputs(1102) <= (layer0_outputs(1845)) xor (layer0_outputs(3596));
    layer1_outputs(1103) <= (layer0_outputs(4677)) and not (layer0_outputs(1505));
    layer1_outputs(1104) <= layer0_outputs(4018);
    layer1_outputs(1105) <= (layer0_outputs(4623)) and not (layer0_outputs(4691));
    layer1_outputs(1106) <= not(layer0_outputs(436));
    layer1_outputs(1107) <= not(layer0_outputs(5004));
    layer1_outputs(1108) <= (layer0_outputs(2369)) and (layer0_outputs(221));
    layer1_outputs(1109) <= (layer0_outputs(259)) and not (layer0_outputs(3437));
    layer1_outputs(1110) <= (layer0_outputs(268)) and (layer0_outputs(1712));
    layer1_outputs(1111) <= layer0_outputs(2292);
    layer1_outputs(1112) <= (layer0_outputs(4529)) or (layer0_outputs(2615));
    layer1_outputs(1113) <= layer0_outputs(4803);
    layer1_outputs(1114) <= (layer0_outputs(4145)) or (layer0_outputs(1826));
    layer1_outputs(1115) <= layer0_outputs(607);
    layer1_outputs(1116) <= (layer0_outputs(1956)) or (layer0_outputs(3371));
    layer1_outputs(1117) <= (layer0_outputs(924)) or (layer0_outputs(2776));
    layer1_outputs(1118) <= (layer0_outputs(3674)) and (layer0_outputs(4217));
    layer1_outputs(1119) <= layer0_outputs(2041);
    layer1_outputs(1120) <= not((layer0_outputs(4407)) xor (layer0_outputs(311)));
    layer1_outputs(1121) <= not((layer0_outputs(3919)) and (layer0_outputs(99)));
    layer1_outputs(1122) <= (layer0_outputs(4298)) and not (layer0_outputs(1600));
    layer1_outputs(1123) <= (layer0_outputs(3997)) and (layer0_outputs(3696));
    layer1_outputs(1124) <= not((layer0_outputs(3651)) or (layer0_outputs(2854)));
    layer1_outputs(1125) <= (layer0_outputs(2885)) and (layer0_outputs(4205));
    layer1_outputs(1126) <= not(layer0_outputs(4003)) or (layer0_outputs(200));
    layer1_outputs(1127) <= not((layer0_outputs(2944)) xor (layer0_outputs(2382)));
    layer1_outputs(1128) <= (layer0_outputs(3129)) xor (layer0_outputs(2189));
    layer1_outputs(1129) <= not(layer0_outputs(2206)) or (layer0_outputs(2610));
    layer1_outputs(1130) <= layer0_outputs(3748);
    layer1_outputs(1131) <= (layer0_outputs(1665)) or (layer0_outputs(3453));
    layer1_outputs(1132) <= '1';
    layer1_outputs(1133) <= (layer0_outputs(4052)) xor (layer0_outputs(2886));
    layer1_outputs(1134) <= not(layer0_outputs(2208));
    layer1_outputs(1135) <= not(layer0_outputs(1714)) or (layer0_outputs(4747));
    layer1_outputs(1136) <= not((layer0_outputs(4357)) and (layer0_outputs(4584)));
    layer1_outputs(1137) <= layer0_outputs(3957);
    layer1_outputs(1138) <= layer0_outputs(3168);
    layer1_outputs(1139) <= (layer0_outputs(4563)) and (layer0_outputs(4390));
    layer1_outputs(1140) <= layer0_outputs(5114);
    layer1_outputs(1141) <= not(layer0_outputs(4830)) or (layer0_outputs(1122));
    layer1_outputs(1142) <= (layer0_outputs(3917)) xor (layer0_outputs(908));
    layer1_outputs(1143) <= (layer0_outputs(3160)) xor (layer0_outputs(1954));
    layer1_outputs(1144) <= layer0_outputs(4111);
    layer1_outputs(1145) <= (layer0_outputs(1224)) and not (layer0_outputs(4573));
    layer1_outputs(1146) <= not(layer0_outputs(3450));
    layer1_outputs(1147) <= (layer0_outputs(1917)) or (layer0_outputs(4826));
    layer1_outputs(1148) <= not(layer0_outputs(981));
    layer1_outputs(1149) <= not(layer0_outputs(2987)) or (layer0_outputs(5109));
    layer1_outputs(1150) <= layer0_outputs(2396);
    layer1_outputs(1151) <= (layer0_outputs(3624)) xor (layer0_outputs(836));
    layer1_outputs(1152) <= not((layer0_outputs(2518)) and (layer0_outputs(3605)));
    layer1_outputs(1153) <= not((layer0_outputs(3766)) or (layer0_outputs(3830)));
    layer1_outputs(1154) <= layer0_outputs(3855);
    layer1_outputs(1155) <= (layer0_outputs(2120)) and not (layer0_outputs(5020));
    layer1_outputs(1156) <= layer0_outputs(4779);
    layer1_outputs(1157) <= layer0_outputs(2658);
    layer1_outputs(1158) <= not(layer0_outputs(2640));
    layer1_outputs(1159) <= layer0_outputs(1388);
    layer1_outputs(1160) <= not(layer0_outputs(1718)) or (layer0_outputs(1218));
    layer1_outputs(1161) <= (layer0_outputs(2963)) xor (layer0_outputs(150));
    layer1_outputs(1162) <= not((layer0_outputs(391)) and (layer0_outputs(3404)));
    layer1_outputs(1163) <= not(layer0_outputs(3739)) or (layer0_outputs(2141));
    layer1_outputs(1164) <= not(layer0_outputs(1321));
    layer1_outputs(1165) <= (layer0_outputs(4087)) xor (layer0_outputs(2213));
    layer1_outputs(1166) <= '1';
    layer1_outputs(1167) <= not(layer0_outputs(986)) or (layer0_outputs(1259));
    layer1_outputs(1168) <= not((layer0_outputs(4319)) or (layer0_outputs(939)));
    layer1_outputs(1169) <= '0';
    layer1_outputs(1170) <= (layer0_outputs(841)) and not (layer0_outputs(2508));
    layer1_outputs(1171) <= not((layer0_outputs(2863)) and (layer0_outputs(3780)));
    layer1_outputs(1172) <= layer0_outputs(2844);
    layer1_outputs(1173) <= '0';
    layer1_outputs(1174) <= (layer0_outputs(3409)) or (layer0_outputs(4170));
    layer1_outputs(1175) <= not((layer0_outputs(3082)) and (layer0_outputs(2188)));
    layer1_outputs(1176) <= layer0_outputs(1918);
    layer1_outputs(1177) <= not(layer0_outputs(1426)) or (layer0_outputs(701));
    layer1_outputs(1178) <= not(layer0_outputs(3654));
    layer1_outputs(1179) <= not(layer0_outputs(4887)) or (layer0_outputs(1133));
    layer1_outputs(1180) <= (layer0_outputs(4055)) and (layer0_outputs(205));
    layer1_outputs(1181) <= not(layer0_outputs(4807));
    layer1_outputs(1182) <= (layer0_outputs(1925)) or (layer0_outputs(1756));
    layer1_outputs(1183) <= layer0_outputs(2191);
    layer1_outputs(1184) <= (layer0_outputs(809)) or (layer0_outputs(2425));
    layer1_outputs(1185) <= (layer0_outputs(2412)) and (layer0_outputs(402));
    layer1_outputs(1186) <= (layer0_outputs(3332)) and (layer0_outputs(2192));
    layer1_outputs(1187) <= (layer0_outputs(1529)) and not (layer0_outputs(2234));
    layer1_outputs(1188) <= not(layer0_outputs(2646));
    layer1_outputs(1189) <= '1';
    layer1_outputs(1190) <= (layer0_outputs(53)) and (layer0_outputs(337));
    layer1_outputs(1191) <= not(layer0_outputs(4426)) or (layer0_outputs(5103));
    layer1_outputs(1192) <= not((layer0_outputs(3679)) or (layer0_outputs(288)));
    layer1_outputs(1193) <= not(layer0_outputs(2724));
    layer1_outputs(1194) <= not(layer0_outputs(1794));
    layer1_outputs(1195) <= not((layer0_outputs(189)) or (layer0_outputs(1264)));
    layer1_outputs(1196) <= not(layer0_outputs(1111)) or (layer0_outputs(310));
    layer1_outputs(1197) <= not((layer0_outputs(267)) xor (layer0_outputs(1821)));
    layer1_outputs(1198) <= not(layer0_outputs(2401));
    layer1_outputs(1199) <= layer0_outputs(2520);
    layer1_outputs(1200) <= layer0_outputs(795);
    layer1_outputs(1201) <= layer0_outputs(1473);
    layer1_outputs(1202) <= not((layer0_outputs(3101)) or (layer0_outputs(2099)));
    layer1_outputs(1203) <= not((layer0_outputs(2662)) and (layer0_outputs(4342)));
    layer1_outputs(1204) <= not(layer0_outputs(2440)) or (layer0_outputs(3971));
    layer1_outputs(1205) <= (layer0_outputs(5001)) and not (layer0_outputs(4422));
    layer1_outputs(1206) <= layer0_outputs(1463);
    layer1_outputs(1207) <= (layer0_outputs(550)) and not (layer0_outputs(846));
    layer1_outputs(1208) <= (layer0_outputs(1147)) and not (layer0_outputs(3403));
    layer1_outputs(1209) <= not(layer0_outputs(3252));
    layer1_outputs(1210) <= (layer0_outputs(4046)) and (layer0_outputs(245));
    layer1_outputs(1211) <= '1';
    layer1_outputs(1212) <= (layer0_outputs(3121)) or (layer0_outputs(3600));
    layer1_outputs(1213) <= (layer0_outputs(2882)) xor (layer0_outputs(584));
    layer1_outputs(1214) <= not((layer0_outputs(4578)) or (layer0_outputs(1464)));
    layer1_outputs(1215) <= (layer0_outputs(3585)) xor (layer0_outputs(3414));
    layer1_outputs(1216) <= layer0_outputs(2319);
    layer1_outputs(1217) <= not((layer0_outputs(1747)) xor (layer0_outputs(3928)));
    layer1_outputs(1218) <= layer0_outputs(1413);
    layer1_outputs(1219) <= layer0_outputs(4160);
    layer1_outputs(1220) <= '0';
    layer1_outputs(1221) <= not((layer0_outputs(2470)) and (layer0_outputs(3347)));
    layer1_outputs(1222) <= (layer0_outputs(108)) and not (layer0_outputs(1958));
    layer1_outputs(1223) <= not((layer0_outputs(4710)) and (layer0_outputs(4611)));
    layer1_outputs(1224) <= (layer0_outputs(2298)) or (layer0_outputs(3734));
    layer1_outputs(1225) <= not(layer0_outputs(2083)) or (layer0_outputs(22));
    layer1_outputs(1226) <= layer0_outputs(523);
    layer1_outputs(1227) <= not((layer0_outputs(2380)) or (layer0_outputs(3883)));
    layer1_outputs(1228) <= not(layer0_outputs(4909));
    layer1_outputs(1229) <= layer0_outputs(517);
    layer1_outputs(1230) <= not(layer0_outputs(2024)) or (layer0_outputs(3561));
    layer1_outputs(1231) <= not(layer0_outputs(3040)) or (layer0_outputs(3258));
    layer1_outputs(1232) <= (layer0_outputs(1551)) or (layer0_outputs(871));
    layer1_outputs(1233) <= not((layer0_outputs(2015)) xor (layer0_outputs(3768)));
    layer1_outputs(1234) <= (layer0_outputs(2097)) and (layer0_outputs(1000));
    layer1_outputs(1235) <= (layer0_outputs(3709)) and not (layer0_outputs(1226));
    layer1_outputs(1236) <= not(layer0_outputs(3350));
    layer1_outputs(1237) <= (layer0_outputs(2436)) and not (layer0_outputs(3435));
    layer1_outputs(1238) <= (layer0_outputs(2633)) and (layer0_outputs(1242));
    layer1_outputs(1239) <= not(layer0_outputs(890)) or (layer0_outputs(2725));
    layer1_outputs(1240) <= (layer0_outputs(3212)) xor (layer0_outputs(4981));
    layer1_outputs(1241) <= (layer0_outputs(3010)) xor (layer0_outputs(4249));
    layer1_outputs(1242) <= not((layer0_outputs(398)) or (layer0_outputs(4738)));
    layer1_outputs(1243) <= layer0_outputs(1424);
    layer1_outputs(1244) <= not(layer0_outputs(4449));
    layer1_outputs(1245) <= not(layer0_outputs(1793)) or (layer0_outputs(3937));
    layer1_outputs(1246) <= '0';
    layer1_outputs(1247) <= layer0_outputs(5101);
    layer1_outputs(1248) <= not(layer0_outputs(4581));
    layer1_outputs(1249) <= not(layer0_outputs(4528)) or (layer0_outputs(1312));
    layer1_outputs(1250) <= not(layer0_outputs(990)) or (layer0_outputs(2862));
    layer1_outputs(1251) <= not(layer0_outputs(799));
    layer1_outputs(1252) <= (layer0_outputs(2344)) and not (layer0_outputs(5063));
    layer1_outputs(1253) <= layer0_outputs(581);
    layer1_outputs(1254) <= not(layer0_outputs(1888));
    layer1_outputs(1255) <= not(layer0_outputs(2830));
    layer1_outputs(1256) <= layer0_outputs(2604);
    layer1_outputs(1257) <= (layer0_outputs(2738)) and not (layer0_outputs(3908));
    layer1_outputs(1258) <= not(layer0_outputs(4451));
    layer1_outputs(1259) <= (layer0_outputs(3013)) or (layer0_outputs(121));
    layer1_outputs(1260) <= (layer0_outputs(3555)) or (layer0_outputs(4566));
    layer1_outputs(1261) <= layer0_outputs(577);
    layer1_outputs(1262) <= not(layer0_outputs(2970));
    layer1_outputs(1263) <= (layer0_outputs(1433)) and (layer0_outputs(2972));
    layer1_outputs(1264) <= not((layer0_outputs(29)) or (layer0_outputs(2769)));
    layer1_outputs(1265) <= not((layer0_outputs(3312)) xor (layer0_outputs(1866)));
    layer1_outputs(1266) <= not(layer0_outputs(2646));
    layer1_outputs(1267) <= not((layer0_outputs(4415)) xor (layer0_outputs(3800)));
    layer1_outputs(1268) <= not(layer0_outputs(323)) or (layer0_outputs(4889));
    layer1_outputs(1269) <= layer0_outputs(2052);
    layer1_outputs(1270) <= not((layer0_outputs(771)) or (layer0_outputs(2572)));
    layer1_outputs(1271) <= not(layer0_outputs(648));
    layer1_outputs(1272) <= layer0_outputs(4238);
    layer1_outputs(1273) <= not(layer0_outputs(792));
    layer1_outputs(1274) <= layer0_outputs(3086);
    layer1_outputs(1275) <= not(layer0_outputs(332)) or (layer0_outputs(4886));
    layer1_outputs(1276) <= not(layer0_outputs(4638)) or (layer0_outputs(949));
    layer1_outputs(1277) <= (layer0_outputs(4771)) and (layer0_outputs(2410));
    layer1_outputs(1278) <= not(layer0_outputs(60));
    layer1_outputs(1279) <= layer0_outputs(4435);
    layer1_outputs(1280) <= not(layer0_outputs(2728)) or (layer0_outputs(2800));
    layer1_outputs(1281) <= '1';
    layer1_outputs(1282) <= not(layer0_outputs(4113));
    layer1_outputs(1283) <= layer0_outputs(2101);
    layer1_outputs(1284) <= not((layer0_outputs(2950)) or (layer0_outputs(3656)));
    layer1_outputs(1285) <= not(layer0_outputs(1222));
    layer1_outputs(1286) <= layer0_outputs(4948);
    layer1_outputs(1287) <= layer0_outputs(4791);
    layer1_outputs(1288) <= layer0_outputs(4740);
    layer1_outputs(1289) <= (layer0_outputs(4424)) xor (layer0_outputs(1584));
    layer1_outputs(1290) <= not(layer0_outputs(3367)) or (layer0_outputs(3507));
    layer1_outputs(1291) <= not(layer0_outputs(365));
    layer1_outputs(1292) <= layer0_outputs(3728);
    layer1_outputs(1293) <= not(layer0_outputs(2063)) or (layer0_outputs(4124));
    layer1_outputs(1294) <= (layer0_outputs(3538)) and not (layer0_outputs(2444));
    layer1_outputs(1295) <= not(layer0_outputs(2172)) or (layer0_outputs(2354));
    layer1_outputs(1296) <= not(layer0_outputs(4066));
    layer1_outputs(1297) <= (layer0_outputs(2885)) and not (layer0_outputs(216));
    layer1_outputs(1298) <= (layer0_outputs(3106)) or (layer0_outputs(2051));
    layer1_outputs(1299) <= not((layer0_outputs(1269)) or (layer0_outputs(4031)));
    layer1_outputs(1300) <= (layer0_outputs(2987)) xor (layer0_outputs(4218));
    layer1_outputs(1301) <= not(layer0_outputs(4601));
    layer1_outputs(1302) <= not(layer0_outputs(612));
    layer1_outputs(1303) <= (layer0_outputs(4286)) and (layer0_outputs(1752));
    layer1_outputs(1304) <= not((layer0_outputs(4991)) or (layer0_outputs(4352)));
    layer1_outputs(1305) <= not((layer0_outputs(2930)) xor (layer0_outputs(1992)));
    layer1_outputs(1306) <= layer0_outputs(4403);
    layer1_outputs(1307) <= layer0_outputs(4177);
    layer1_outputs(1308) <= not((layer0_outputs(3259)) xor (layer0_outputs(745)));
    layer1_outputs(1309) <= not((layer0_outputs(4845)) or (layer0_outputs(1575)));
    layer1_outputs(1310) <= not(layer0_outputs(3914)) or (layer0_outputs(4930));
    layer1_outputs(1311) <= layer0_outputs(2686);
    layer1_outputs(1312) <= not(layer0_outputs(1839)) or (layer0_outputs(2604));
    layer1_outputs(1313) <= not(layer0_outputs(2406));
    layer1_outputs(1314) <= not(layer0_outputs(2292)) or (layer0_outputs(3397));
    layer1_outputs(1315) <= layer0_outputs(1871);
    layer1_outputs(1316) <= '1';
    layer1_outputs(1317) <= not((layer0_outputs(4585)) and (layer0_outputs(1869)));
    layer1_outputs(1318) <= (layer0_outputs(4299)) and (layer0_outputs(1386));
    layer1_outputs(1319) <= (layer0_outputs(3272)) and not (layer0_outputs(4568));
    layer1_outputs(1320) <= '0';
    layer1_outputs(1321) <= layer0_outputs(4901);
    layer1_outputs(1322) <= (layer0_outputs(4801)) and (layer0_outputs(694));
    layer1_outputs(1323) <= '1';
    layer1_outputs(1324) <= (layer0_outputs(3386)) xor (layer0_outputs(3846));
    layer1_outputs(1325) <= not((layer0_outputs(2107)) or (layer0_outputs(4616)));
    layer1_outputs(1326) <= not(layer0_outputs(891));
    layer1_outputs(1327) <= not((layer0_outputs(3550)) or (layer0_outputs(12)));
    layer1_outputs(1328) <= not(layer0_outputs(1189)) or (layer0_outputs(1852));
    layer1_outputs(1329) <= (layer0_outputs(3348)) or (layer0_outputs(1786));
    layer1_outputs(1330) <= layer0_outputs(1817);
    layer1_outputs(1331) <= '1';
    layer1_outputs(1332) <= not(layer0_outputs(3256)) or (layer0_outputs(194));
    layer1_outputs(1333) <= (layer0_outputs(3218)) and not (layer0_outputs(93));
    layer1_outputs(1334) <= (layer0_outputs(2567)) and not (layer0_outputs(3028));
    layer1_outputs(1335) <= not(layer0_outputs(3315)) or (layer0_outputs(567));
    layer1_outputs(1336) <= not(layer0_outputs(4817)) or (layer0_outputs(1154));
    layer1_outputs(1337) <= not(layer0_outputs(1311));
    layer1_outputs(1338) <= not(layer0_outputs(3627)) or (layer0_outputs(4575));
    layer1_outputs(1339) <= not(layer0_outputs(3808)) or (layer0_outputs(3074));
    layer1_outputs(1340) <= '1';
    layer1_outputs(1341) <= layer0_outputs(2943);
    layer1_outputs(1342) <= not(layer0_outputs(2770)) or (layer0_outputs(4191));
    layer1_outputs(1343) <= not(layer0_outputs(2081)) or (layer0_outputs(1596));
    layer1_outputs(1344) <= layer0_outputs(3209);
    layer1_outputs(1345) <= layer0_outputs(3432);
    layer1_outputs(1346) <= not(layer0_outputs(1330));
    layer1_outputs(1347) <= (layer0_outputs(3746)) and not (layer0_outputs(2812));
    layer1_outputs(1348) <= (layer0_outputs(1554)) and not (layer0_outputs(1716));
    layer1_outputs(1349) <= layer0_outputs(2287);
    layer1_outputs(1350) <= (layer0_outputs(806)) or (layer0_outputs(703));
    layer1_outputs(1351) <= (layer0_outputs(2628)) or (layer0_outputs(711));
    layer1_outputs(1352) <= layer0_outputs(1454);
    layer1_outputs(1353) <= (layer0_outputs(445)) or (layer0_outputs(3572));
    layer1_outputs(1354) <= (layer0_outputs(686)) and not (layer0_outputs(5038));
    layer1_outputs(1355) <= '1';
    layer1_outputs(1356) <= not(layer0_outputs(4437)) or (layer0_outputs(1885));
    layer1_outputs(1357) <= not(layer0_outputs(4075));
    layer1_outputs(1358) <= layer0_outputs(1773);
    layer1_outputs(1359) <= (layer0_outputs(2140)) and not (layer0_outputs(467));
    layer1_outputs(1360) <= (layer0_outputs(56)) and not (layer0_outputs(3121));
    layer1_outputs(1361) <= not((layer0_outputs(4412)) and (layer0_outputs(3226)));
    layer1_outputs(1362) <= (layer0_outputs(3658)) xor (layer0_outputs(1260));
    layer1_outputs(1363) <= not(layer0_outputs(4479));
    layer1_outputs(1364) <= (layer0_outputs(1057)) xor (layer0_outputs(1586));
    layer1_outputs(1365) <= (layer0_outputs(91)) and not (layer0_outputs(3678));
    layer1_outputs(1366) <= not(layer0_outputs(4146)) or (layer0_outputs(1048));
    layer1_outputs(1367) <= not(layer0_outputs(1420));
    layer1_outputs(1368) <= (layer0_outputs(1465)) xor (layer0_outputs(2326));
    layer1_outputs(1369) <= not((layer0_outputs(3780)) and (layer0_outputs(3459)));
    layer1_outputs(1370) <= (layer0_outputs(1766)) and not (layer0_outputs(4021));
    layer1_outputs(1371) <= not((layer0_outputs(4669)) or (layer0_outputs(3986)));
    layer1_outputs(1372) <= (layer0_outputs(4094)) xor (layer0_outputs(4854));
    layer1_outputs(1373) <= '1';
    layer1_outputs(1374) <= not(layer0_outputs(4944));
    layer1_outputs(1375) <= not(layer0_outputs(46)) or (layer0_outputs(3130));
    layer1_outputs(1376) <= not(layer0_outputs(381));
    layer1_outputs(1377) <= (layer0_outputs(1975)) and not (layer0_outputs(3794));
    layer1_outputs(1378) <= not(layer0_outputs(3878));
    layer1_outputs(1379) <= layer0_outputs(4355);
    layer1_outputs(1380) <= (layer0_outputs(4308)) and not (layer0_outputs(3437));
    layer1_outputs(1381) <= (layer0_outputs(3649)) and not (layer0_outputs(1333));
    layer1_outputs(1382) <= (layer0_outputs(3293)) and (layer0_outputs(4235));
    layer1_outputs(1383) <= (layer0_outputs(2964)) and (layer0_outputs(3008));
    layer1_outputs(1384) <= (layer0_outputs(2628)) and not (layer0_outputs(3722));
    layer1_outputs(1385) <= (layer0_outputs(3362)) and not (layer0_outputs(2884));
    layer1_outputs(1386) <= not(layer0_outputs(4223)) or (layer0_outputs(3089));
    layer1_outputs(1387) <= not(layer0_outputs(783)) or (layer0_outputs(3882));
    layer1_outputs(1388) <= not(layer0_outputs(2786)) or (layer0_outputs(1345));
    layer1_outputs(1389) <= not(layer0_outputs(4692));
    layer1_outputs(1390) <= layer0_outputs(4374);
    layer1_outputs(1391) <= (layer0_outputs(3443)) and not (layer0_outputs(4695));
    layer1_outputs(1392) <= not(layer0_outputs(2928));
    layer1_outputs(1393) <= '1';
    layer1_outputs(1394) <= not((layer0_outputs(601)) xor (layer0_outputs(1990)));
    layer1_outputs(1395) <= '1';
    layer1_outputs(1396) <= not((layer0_outputs(2741)) or (layer0_outputs(4125)));
    layer1_outputs(1397) <= (layer0_outputs(103)) and not (layer0_outputs(2718));
    layer1_outputs(1398) <= layer0_outputs(2579);
    layer1_outputs(1399) <= layer0_outputs(1217);
    layer1_outputs(1400) <= (layer0_outputs(2339)) or (layer0_outputs(1154));
    layer1_outputs(1401) <= (layer0_outputs(1977)) or (layer0_outputs(2320));
    layer1_outputs(1402) <= not(layer0_outputs(2756)) or (layer0_outputs(2961));
    layer1_outputs(1403) <= '1';
    layer1_outputs(1404) <= layer0_outputs(4491);
    layer1_outputs(1405) <= not((layer0_outputs(181)) or (layer0_outputs(2869)));
    layer1_outputs(1406) <= (layer0_outputs(4687)) and not (layer0_outputs(4108));
    layer1_outputs(1407) <= (layer0_outputs(4265)) and not (layer0_outputs(1483));
    layer1_outputs(1408) <= not(layer0_outputs(2896));
    layer1_outputs(1409) <= (layer0_outputs(4194)) xor (layer0_outputs(4320));
    layer1_outputs(1410) <= '0';
    layer1_outputs(1411) <= layer0_outputs(3633);
    layer1_outputs(1412) <= not(layer0_outputs(2551));
    layer1_outputs(1413) <= '1';
    layer1_outputs(1414) <= not(layer0_outputs(1260)) or (layer0_outputs(1909));
    layer1_outputs(1415) <= not(layer0_outputs(602)) or (layer0_outputs(418));
    layer1_outputs(1416) <= not((layer0_outputs(1534)) xor (layer0_outputs(4937)));
    layer1_outputs(1417) <= layer0_outputs(732);
    layer1_outputs(1418) <= '1';
    layer1_outputs(1419) <= not(layer0_outputs(664));
    layer1_outputs(1420) <= (layer0_outputs(4712)) and (layer0_outputs(5005));
    layer1_outputs(1421) <= not((layer0_outputs(2620)) and (layer0_outputs(2395)));
    layer1_outputs(1422) <= not((layer0_outputs(4332)) xor (layer0_outputs(1921)));
    layer1_outputs(1423) <= not(layer0_outputs(870));
    layer1_outputs(1424) <= not(layer0_outputs(4154));
    layer1_outputs(1425) <= not((layer0_outputs(4275)) or (layer0_outputs(2473)));
    layer1_outputs(1426) <= '1';
    layer1_outputs(1427) <= layer0_outputs(4621);
    layer1_outputs(1428) <= (layer0_outputs(3532)) and not (layer0_outputs(4569));
    layer1_outputs(1429) <= layer0_outputs(364);
    layer1_outputs(1430) <= (layer0_outputs(3065)) or (layer0_outputs(3207));
    layer1_outputs(1431) <= not(layer0_outputs(970)) or (layer0_outputs(1945));
    layer1_outputs(1432) <= not(layer0_outputs(3589));
    layer1_outputs(1433) <= not(layer0_outputs(2456));
    layer1_outputs(1434) <= (layer0_outputs(2642)) and not (layer0_outputs(428));
    layer1_outputs(1435) <= not(layer0_outputs(1229));
    layer1_outputs(1436) <= not(layer0_outputs(3854)) or (layer0_outputs(1459));
    layer1_outputs(1437) <= (layer0_outputs(1974)) and (layer0_outputs(4695));
    layer1_outputs(1438) <= layer0_outputs(3645);
    layer1_outputs(1439) <= (layer0_outputs(2626)) and not (layer0_outputs(2277));
    layer1_outputs(1440) <= not(layer0_outputs(4330)) or (layer0_outputs(431));
    layer1_outputs(1441) <= (layer0_outputs(1209)) or (layer0_outputs(3951));
    layer1_outputs(1442) <= not((layer0_outputs(2248)) and (layer0_outputs(3794)));
    layer1_outputs(1443) <= layer0_outputs(4579);
    layer1_outputs(1444) <= '1';
    layer1_outputs(1445) <= not((layer0_outputs(1417)) and (layer0_outputs(2011)));
    layer1_outputs(1446) <= layer0_outputs(2990);
    layer1_outputs(1447) <= layer0_outputs(190);
    layer1_outputs(1448) <= layer0_outputs(1936);
    layer1_outputs(1449) <= not(layer0_outputs(2702));
    layer1_outputs(1450) <= layer0_outputs(806);
    layer1_outputs(1451) <= not(layer0_outputs(516));
    layer1_outputs(1452) <= not((layer0_outputs(5109)) xor (layer0_outputs(4602)));
    layer1_outputs(1453) <= not((layer0_outputs(1988)) and (layer0_outputs(1083)));
    layer1_outputs(1454) <= not(layer0_outputs(3159));
    layer1_outputs(1455) <= (layer0_outputs(4352)) and (layer0_outputs(3382));
    layer1_outputs(1456) <= '0';
    layer1_outputs(1457) <= layer0_outputs(1364);
    layer1_outputs(1458) <= not((layer0_outputs(642)) and (layer0_outputs(3351)));
    layer1_outputs(1459) <= '0';
    layer1_outputs(1460) <= layer0_outputs(3707);
    layer1_outputs(1461) <= not(layer0_outputs(2538));
    layer1_outputs(1462) <= layer0_outputs(2806);
    layer1_outputs(1463) <= not((layer0_outputs(829)) or (layer0_outputs(2129)));
    layer1_outputs(1464) <= not(layer0_outputs(3069)) or (layer0_outputs(1881));
    layer1_outputs(1465) <= (layer0_outputs(113)) and not (layer0_outputs(4047));
    layer1_outputs(1466) <= not((layer0_outputs(823)) or (layer0_outputs(117)));
    layer1_outputs(1467) <= (layer0_outputs(2796)) or (layer0_outputs(1289));
    layer1_outputs(1468) <= not((layer0_outputs(167)) or (layer0_outputs(2661)));
    layer1_outputs(1469) <= not((layer0_outputs(141)) or (layer0_outputs(3203)));
    layer1_outputs(1470) <= not(layer0_outputs(457));
    layer1_outputs(1471) <= not(layer0_outputs(5077));
    layer1_outputs(1472) <= (layer0_outputs(222)) and (layer0_outputs(588));
    layer1_outputs(1473) <= layer0_outputs(1602);
    layer1_outputs(1474) <= layer0_outputs(1448);
    layer1_outputs(1475) <= not(layer0_outputs(455));
    layer1_outputs(1476) <= not(layer0_outputs(3627));
    layer1_outputs(1477) <= layer0_outputs(3265);
    layer1_outputs(1478) <= not(layer0_outputs(2971)) or (layer0_outputs(1337));
    layer1_outputs(1479) <= (layer0_outputs(714)) and not (layer0_outputs(3022));
    layer1_outputs(1480) <= not(layer0_outputs(1675));
    layer1_outputs(1481) <= (layer0_outputs(4200)) or (layer0_outputs(4029));
    layer1_outputs(1482) <= not(layer0_outputs(2407));
    layer1_outputs(1483) <= not((layer0_outputs(3038)) and (layer0_outputs(2514)));
    layer1_outputs(1484) <= layer0_outputs(149);
    layer1_outputs(1485) <= not(layer0_outputs(2385));
    layer1_outputs(1486) <= not((layer0_outputs(1135)) and (layer0_outputs(1725)));
    layer1_outputs(1487) <= not(layer0_outputs(4935));
    layer1_outputs(1488) <= not((layer0_outputs(1326)) xor (layer0_outputs(2444)));
    layer1_outputs(1489) <= layer0_outputs(2307);
    layer1_outputs(1490) <= layer0_outputs(2546);
    layer1_outputs(1491) <= not(layer0_outputs(184)) or (layer0_outputs(412));
    layer1_outputs(1492) <= not(layer0_outputs(652));
    layer1_outputs(1493) <= (layer0_outputs(2447)) and (layer0_outputs(1941));
    layer1_outputs(1494) <= (layer0_outputs(214)) and (layer0_outputs(4264));
    layer1_outputs(1495) <= not((layer0_outputs(1373)) xor (layer0_outputs(286)));
    layer1_outputs(1496) <= (layer0_outputs(1738)) or (layer0_outputs(4576));
    layer1_outputs(1497) <= not(layer0_outputs(174));
    layer1_outputs(1498) <= (layer0_outputs(4766)) and not (layer0_outputs(5013));
    layer1_outputs(1499) <= not((layer0_outputs(4050)) and (layer0_outputs(3543)));
    layer1_outputs(1500) <= '0';
    layer1_outputs(1501) <= (layer0_outputs(4443)) and (layer0_outputs(4595));
    layer1_outputs(1502) <= layer0_outputs(1204);
    layer1_outputs(1503) <= not(layer0_outputs(172));
    layer1_outputs(1504) <= (layer0_outputs(2351)) and not (layer0_outputs(2683));
    layer1_outputs(1505) <= (layer0_outputs(493)) and (layer0_outputs(1983));
    layer1_outputs(1506) <= (layer0_outputs(2560)) and not (layer0_outputs(3025));
    layer1_outputs(1507) <= not(layer0_outputs(418));
    layer1_outputs(1508) <= not(layer0_outputs(335)) or (layer0_outputs(1040));
    layer1_outputs(1509) <= (layer0_outputs(2758)) and (layer0_outputs(4971));
    layer1_outputs(1510) <= (layer0_outputs(4429)) and not (layer0_outputs(3921));
    layer1_outputs(1511) <= layer0_outputs(25);
    layer1_outputs(1512) <= (layer0_outputs(5085)) and (layer0_outputs(2913));
    layer1_outputs(1513) <= not((layer0_outputs(109)) and (layer0_outputs(443)));
    layer1_outputs(1514) <= (layer0_outputs(2745)) and not (layer0_outputs(4985));
    layer1_outputs(1515) <= layer0_outputs(1181);
    layer1_outputs(1516) <= (layer0_outputs(822)) and not (layer0_outputs(3604));
    layer1_outputs(1517) <= (layer0_outputs(4072)) and not (layer0_outputs(3920));
    layer1_outputs(1518) <= (layer0_outputs(2545)) and not (layer0_outputs(4772));
    layer1_outputs(1519) <= not(layer0_outputs(1192));
    layer1_outputs(1520) <= not((layer0_outputs(4787)) and (layer0_outputs(842)));
    layer1_outputs(1521) <= (layer0_outputs(4823)) and (layer0_outputs(4943));
    layer1_outputs(1522) <= not(layer0_outputs(4481));
    layer1_outputs(1523) <= not((layer0_outputs(4171)) and (layer0_outputs(1722)));
    layer1_outputs(1524) <= (layer0_outputs(4550)) and not (layer0_outputs(3372));
    layer1_outputs(1525) <= (layer0_outputs(794)) and not (layer0_outputs(2102));
    layer1_outputs(1526) <= (layer0_outputs(311)) and not (layer0_outputs(3137));
    layer1_outputs(1527) <= layer0_outputs(2158);
    layer1_outputs(1528) <= layer0_outputs(3614);
    layer1_outputs(1529) <= layer0_outputs(3769);
    layer1_outputs(1530) <= not(layer0_outputs(795)) or (layer0_outputs(4631));
    layer1_outputs(1531) <= '0';
    layer1_outputs(1532) <= not(layer0_outputs(4216)) or (layer0_outputs(3027));
    layer1_outputs(1533) <= not((layer0_outputs(2314)) and (layer0_outputs(1233)));
    layer1_outputs(1534) <= layer0_outputs(4207);
    layer1_outputs(1535) <= not(layer0_outputs(3894));
    layer1_outputs(1536) <= (layer0_outputs(3765)) and not (layer0_outputs(2220));
    layer1_outputs(1537) <= (layer0_outputs(859)) and not (layer0_outputs(2666));
    layer1_outputs(1538) <= layer0_outputs(4676);
    layer1_outputs(1539) <= not((layer0_outputs(1159)) xor (layer0_outputs(918)));
    layer1_outputs(1540) <= (layer0_outputs(1932)) and (layer0_outputs(2588));
    layer1_outputs(1541) <= not(layer0_outputs(1979)) or (layer0_outputs(2156));
    layer1_outputs(1542) <= not(layer0_outputs(4746));
    layer1_outputs(1543) <= not(layer0_outputs(2813));
    layer1_outputs(1544) <= not((layer0_outputs(998)) and (layer0_outputs(3728)));
    layer1_outputs(1545) <= not(layer0_outputs(4404));
    layer1_outputs(1546) <= (layer0_outputs(919)) or (layer0_outputs(3798));
    layer1_outputs(1547) <= not(layer0_outputs(506)) or (layer0_outputs(2701));
    layer1_outputs(1548) <= layer0_outputs(223);
    layer1_outputs(1549) <= not(layer0_outputs(3754));
    layer1_outputs(1550) <= (layer0_outputs(3344)) xor (layer0_outputs(491));
    layer1_outputs(1551) <= layer0_outputs(359);
    layer1_outputs(1552) <= not(layer0_outputs(4515));
    layer1_outputs(1553) <= layer0_outputs(586);
    layer1_outputs(1554) <= (layer0_outputs(3170)) and not (layer0_outputs(3310));
    layer1_outputs(1555) <= not(layer0_outputs(1136));
    layer1_outputs(1556) <= layer0_outputs(1389);
    layer1_outputs(1557) <= (layer0_outputs(4404)) and not (layer0_outputs(2421));
    layer1_outputs(1558) <= layer0_outputs(1658);
    layer1_outputs(1559) <= layer0_outputs(3324);
    layer1_outputs(1560) <= layer0_outputs(432);
    layer1_outputs(1561) <= not((layer0_outputs(171)) xor (layer0_outputs(4495)));
    layer1_outputs(1562) <= not(layer0_outputs(3134)) or (layer0_outputs(10));
    layer1_outputs(1563) <= not(layer0_outputs(5017));
    layer1_outputs(1564) <= layer0_outputs(1842);
    layer1_outputs(1565) <= layer0_outputs(4758);
    layer1_outputs(1566) <= not(layer0_outputs(1357)) or (layer0_outputs(1939));
    layer1_outputs(1567) <= layer0_outputs(1184);
    layer1_outputs(1568) <= not(layer0_outputs(2172)) or (layer0_outputs(1810));
    layer1_outputs(1569) <= layer0_outputs(651);
    layer1_outputs(1570) <= not(layer0_outputs(3050));
    layer1_outputs(1571) <= not(layer0_outputs(4430)) or (layer0_outputs(1091));
    layer1_outputs(1572) <= not(layer0_outputs(1926)) or (layer0_outputs(896));
    layer1_outputs(1573) <= (layer0_outputs(144)) xor (layer0_outputs(1717));
    layer1_outputs(1574) <= not((layer0_outputs(4815)) and (layer0_outputs(2372)));
    layer1_outputs(1575) <= not((layer0_outputs(4028)) xor (layer0_outputs(1369)));
    layer1_outputs(1576) <= layer0_outputs(3789);
    layer1_outputs(1577) <= layer0_outputs(3926);
    layer1_outputs(1578) <= (layer0_outputs(1364)) xor (layer0_outputs(3164));
    layer1_outputs(1579) <= (layer0_outputs(2902)) and not (layer0_outputs(4407));
    layer1_outputs(1580) <= not((layer0_outputs(4661)) or (layer0_outputs(4324)));
    layer1_outputs(1581) <= not(layer0_outputs(1493)) or (layer0_outputs(1086));
    layer1_outputs(1582) <= (layer0_outputs(2114)) and not (layer0_outputs(194));
    layer1_outputs(1583) <= (layer0_outputs(1070)) xor (layer0_outputs(1815));
    layer1_outputs(1584) <= (layer0_outputs(1801)) xor (layer0_outputs(1066));
    layer1_outputs(1585) <= layer0_outputs(4305);
    layer1_outputs(1586) <= (layer0_outputs(3039)) xor (layer0_outputs(3140));
    layer1_outputs(1587) <= layer0_outputs(3423);
    layer1_outputs(1588) <= not((layer0_outputs(2059)) or (layer0_outputs(3152)));
    layer1_outputs(1589) <= not((layer0_outputs(3673)) xor (layer0_outputs(1977)));
    layer1_outputs(1590) <= (layer0_outputs(3916)) or (layer0_outputs(4102));
    layer1_outputs(1591) <= (layer0_outputs(4563)) and (layer0_outputs(1282));
    layer1_outputs(1592) <= not(layer0_outputs(4701));
    layer1_outputs(1593) <= layer0_outputs(1329);
    layer1_outputs(1594) <= not(layer0_outputs(518));
    layer1_outputs(1595) <= not(layer0_outputs(1226));
    layer1_outputs(1596) <= not(layer0_outputs(4714));
    layer1_outputs(1597) <= layer0_outputs(960);
    layer1_outputs(1598) <= not(layer0_outputs(3215));
    layer1_outputs(1599) <= not(layer0_outputs(1555));
    layer1_outputs(1600) <= (layer0_outputs(2673)) and not (layer0_outputs(247));
    layer1_outputs(1601) <= layer0_outputs(1743);
    layer1_outputs(1602) <= '1';
    layer1_outputs(1603) <= '1';
    layer1_outputs(1604) <= (layer0_outputs(3953)) and (layer0_outputs(5048));
    layer1_outputs(1605) <= not((layer0_outputs(3742)) xor (layer0_outputs(3922)));
    layer1_outputs(1606) <= not((layer0_outputs(1661)) or (layer0_outputs(112)));
    layer1_outputs(1607) <= '1';
    layer1_outputs(1608) <= (layer0_outputs(2569)) and not (layer0_outputs(2431));
    layer1_outputs(1609) <= not((layer0_outputs(2146)) or (layer0_outputs(4840)));
    layer1_outputs(1610) <= not(layer0_outputs(3543)) or (layer0_outputs(59));
    layer1_outputs(1611) <= layer0_outputs(3713);
    layer1_outputs(1612) <= '0';
    layer1_outputs(1613) <= layer0_outputs(2186);
    layer1_outputs(1614) <= not(layer0_outputs(2450));
    layer1_outputs(1615) <= (layer0_outputs(3775)) xor (layer0_outputs(3910));
    layer1_outputs(1616) <= not(layer0_outputs(1278));
    layer1_outputs(1617) <= layer0_outputs(1886);
    layer1_outputs(1618) <= layer0_outputs(138);
    layer1_outputs(1619) <= not(layer0_outputs(258));
    layer1_outputs(1620) <= not((layer0_outputs(3339)) and (layer0_outputs(3694)));
    layer1_outputs(1621) <= not(layer0_outputs(475)) or (layer0_outputs(646));
    layer1_outputs(1622) <= '0';
    layer1_outputs(1623) <= (layer0_outputs(1271)) and not (layer0_outputs(3220));
    layer1_outputs(1624) <= (layer0_outputs(647)) and not (layer0_outputs(376));
    layer1_outputs(1625) <= layer0_outputs(4385);
    layer1_outputs(1626) <= layer0_outputs(3987);
    layer1_outputs(1627) <= (layer0_outputs(3595)) and not (layer0_outputs(835));
    layer1_outputs(1628) <= not(layer0_outputs(3884)) or (layer0_outputs(2714));
    layer1_outputs(1629) <= layer0_outputs(4468);
    layer1_outputs(1630) <= (layer0_outputs(1685)) or (layer0_outputs(2343));
    layer1_outputs(1631) <= not(layer0_outputs(3877));
    layer1_outputs(1632) <= layer0_outputs(2774);
    layer1_outputs(1633) <= not((layer0_outputs(2977)) xor (layer0_outputs(3073)));
    layer1_outputs(1634) <= (layer0_outputs(2624)) and not (layer0_outputs(2636));
    layer1_outputs(1635) <= (layer0_outputs(2619)) and (layer0_outputs(1883));
    layer1_outputs(1636) <= not(layer0_outputs(3582));
    layer1_outputs(1637) <= not(layer0_outputs(122));
    layer1_outputs(1638) <= not(layer0_outputs(2436));
    layer1_outputs(1639) <= '1';
    layer1_outputs(1640) <= not(layer0_outputs(349));
    layer1_outputs(1641) <= not(layer0_outputs(894));
    layer1_outputs(1642) <= not((layer0_outputs(2888)) and (layer0_outputs(573)));
    layer1_outputs(1643) <= (layer0_outputs(3918)) and (layer0_outputs(3956));
    layer1_outputs(1644) <= (layer0_outputs(5008)) and (layer0_outputs(2698));
    layer1_outputs(1645) <= layer0_outputs(1535);
    layer1_outputs(1646) <= (layer0_outputs(2908)) or (layer0_outputs(932));
    layer1_outputs(1647) <= layer0_outputs(2743);
    layer1_outputs(1648) <= (layer0_outputs(1942)) and not (layer0_outputs(3163));
    layer1_outputs(1649) <= layer0_outputs(1831);
    layer1_outputs(1650) <= layer0_outputs(3005);
    layer1_outputs(1651) <= (layer0_outputs(146)) and (layer0_outputs(2316));
    layer1_outputs(1652) <= not(layer0_outputs(4466));
    layer1_outputs(1653) <= layer0_outputs(3165);
    layer1_outputs(1654) <= (layer0_outputs(2162)) and not (layer0_outputs(4709));
    layer1_outputs(1655) <= not((layer0_outputs(1738)) and (layer0_outputs(5091)));
    layer1_outputs(1656) <= not(layer0_outputs(3491)) or (layer0_outputs(3328));
    layer1_outputs(1657) <= not(layer0_outputs(981));
    layer1_outputs(1658) <= not(layer0_outputs(4074));
    layer1_outputs(1659) <= not(layer0_outputs(4295));
    layer1_outputs(1660) <= (layer0_outputs(4146)) xor (layer0_outputs(4335));
    layer1_outputs(1661) <= layer0_outputs(1790);
    layer1_outputs(1662) <= not(layer0_outputs(2696)) or (layer0_outputs(1474));
    layer1_outputs(1663) <= (layer0_outputs(3183)) and not (layer0_outputs(3636));
    layer1_outputs(1664) <= not((layer0_outputs(3086)) or (layer0_outputs(2358)));
    layer1_outputs(1665) <= not((layer0_outputs(1762)) or (layer0_outputs(87)));
    layer1_outputs(1666) <= not((layer0_outputs(3462)) and (layer0_outputs(3492)));
    layer1_outputs(1667) <= (layer0_outputs(3973)) and (layer0_outputs(18));
    layer1_outputs(1668) <= not(layer0_outputs(4027));
    layer1_outputs(1669) <= not(layer0_outputs(4610));
    layer1_outputs(1670) <= not(layer0_outputs(1925)) or (layer0_outputs(4375));
    layer1_outputs(1671) <= (layer0_outputs(1185)) and (layer0_outputs(5066));
    layer1_outputs(1672) <= layer0_outputs(537);
    layer1_outputs(1673) <= layer0_outputs(2634);
    layer1_outputs(1674) <= not(layer0_outputs(987));
    layer1_outputs(1675) <= (layer0_outputs(4777)) and not (layer0_outputs(809));
    layer1_outputs(1676) <= (layer0_outputs(2465)) and (layer0_outputs(710));
    layer1_outputs(1677) <= layer0_outputs(4566);
    layer1_outputs(1678) <= layer0_outputs(2614);
    layer1_outputs(1679) <= not(layer0_outputs(1178)) or (layer0_outputs(4115));
    layer1_outputs(1680) <= (layer0_outputs(963)) and (layer0_outputs(2682));
    layer1_outputs(1681) <= layer0_outputs(2039);
    layer1_outputs(1682) <= (layer0_outputs(2439)) and not (layer0_outputs(2613));
    layer1_outputs(1683) <= not((layer0_outputs(845)) xor (layer0_outputs(2104)));
    layer1_outputs(1684) <= not(layer0_outputs(2944));
    layer1_outputs(1685) <= not(layer0_outputs(2174));
    layer1_outputs(1686) <= not(layer0_outputs(1445));
    layer1_outputs(1687) <= (layer0_outputs(2742)) and not (layer0_outputs(3247));
    layer1_outputs(1688) <= not(layer0_outputs(3178));
    layer1_outputs(1689) <= layer0_outputs(4907);
    layer1_outputs(1690) <= (layer0_outputs(1304)) and not (layer0_outputs(4642));
    layer1_outputs(1691) <= not(layer0_outputs(2241));
    layer1_outputs(1692) <= (layer0_outputs(1418)) and (layer0_outputs(1227));
    layer1_outputs(1693) <= (layer0_outputs(1916)) xor (layer0_outputs(3905));
    layer1_outputs(1694) <= layer0_outputs(2706);
    layer1_outputs(1695) <= (layer0_outputs(2864)) and not (layer0_outputs(933));
    layer1_outputs(1696) <= not(layer0_outputs(2244));
    layer1_outputs(1697) <= layer0_outputs(4047);
    layer1_outputs(1698) <= not((layer0_outputs(3865)) or (layer0_outputs(4856)));
    layer1_outputs(1699) <= not(layer0_outputs(3629));
    layer1_outputs(1700) <= (layer0_outputs(4199)) and not (layer0_outputs(2141));
    layer1_outputs(1701) <= layer0_outputs(2096);
    layer1_outputs(1702) <= layer0_outputs(3407);
    layer1_outputs(1703) <= not((layer0_outputs(319)) or (layer0_outputs(2187)));
    layer1_outputs(1704) <= (layer0_outputs(3123)) and (layer0_outputs(3348));
    layer1_outputs(1705) <= (layer0_outputs(2730)) and (layer0_outputs(3547));
    layer1_outputs(1706) <= not(layer0_outputs(2000)) or (layer0_outputs(2768));
    layer1_outputs(1707) <= layer0_outputs(5024);
    layer1_outputs(1708) <= (layer0_outputs(1618)) and not (layer0_outputs(1776));
    layer1_outputs(1709) <= not(layer0_outputs(2378));
    layer1_outputs(1710) <= (layer0_outputs(1280)) and not (layer0_outputs(2982));
    layer1_outputs(1711) <= (layer0_outputs(2720)) and (layer0_outputs(2353));
    layer1_outputs(1712) <= (layer0_outputs(2582)) and not (layer0_outputs(5067));
    layer1_outputs(1713) <= (layer0_outputs(869)) and (layer0_outputs(4154));
    layer1_outputs(1714) <= '0';
    layer1_outputs(1715) <= not(layer0_outputs(146)) or (layer0_outputs(893));
    layer1_outputs(1716) <= not((layer0_outputs(1644)) or (layer0_outputs(2960)));
    layer1_outputs(1717) <= layer0_outputs(3744);
    layer1_outputs(1718) <= (layer0_outputs(1413)) and (layer0_outputs(3524));
    layer1_outputs(1719) <= not((layer0_outputs(2096)) or (layer0_outputs(2907)));
    layer1_outputs(1720) <= (layer0_outputs(2508)) and (layer0_outputs(3790));
    layer1_outputs(1721) <= not((layer0_outputs(3297)) or (layer0_outputs(1815)));
    layer1_outputs(1722) <= not((layer0_outputs(707)) xor (layer0_outputs(3539)));
    layer1_outputs(1723) <= (layer0_outputs(3360)) and not (layer0_outputs(2532));
    layer1_outputs(1724) <= (layer0_outputs(912)) or (layer0_outputs(271));
    layer1_outputs(1725) <= (layer0_outputs(2947)) or (layer0_outputs(1506));
    layer1_outputs(1726) <= not(layer0_outputs(2272));
    layer1_outputs(1727) <= (layer0_outputs(2519)) and (layer0_outputs(610));
    layer1_outputs(1728) <= (layer0_outputs(1006)) and not (layer0_outputs(4522));
    layer1_outputs(1729) <= layer0_outputs(2106);
    layer1_outputs(1730) <= not((layer0_outputs(2010)) xor (layer0_outputs(2704)));
    layer1_outputs(1731) <= '0';
    layer1_outputs(1732) <= not((layer0_outputs(2630)) xor (layer0_outputs(2768)));
    layer1_outputs(1733) <= (layer0_outputs(3666)) or (layer0_outputs(1439));
    layer1_outputs(1734) <= not((layer0_outputs(5022)) or (layer0_outputs(2422)));
    layer1_outputs(1735) <= not((layer0_outputs(4890)) or (layer0_outputs(3035)));
    layer1_outputs(1736) <= (layer0_outputs(3426)) xor (layer0_outputs(673));
    layer1_outputs(1737) <= not(layer0_outputs(368));
    layer1_outputs(1738) <= (layer0_outputs(4648)) xor (layer0_outputs(1665));
    layer1_outputs(1739) <= not((layer0_outputs(1677)) and (layer0_outputs(690)));
    layer1_outputs(1740) <= (layer0_outputs(1978)) and not (layer0_outputs(3092));
    layer1_outputs(1741) <= not((layer0_outputs(40)) xor (layer0_outputs(3998)));
    layer1_outputs(1742) <= not(layer0_outputs(2200));
    layer1_outputs(1743) <= (layer0_outputs(3659)) and not (layer0_outputs(1689));
    layer1_outputs(1744) <= (layer0_outputs(3871)) and (layer0_outputs(699));
    layer1_outputs(1745) <= not(layer0_outputs(2152)) or (layer0_outputs(1441));
    layer1_outputs(1746) <= not((layer0_outputs(1720)) xor (layer0_outputs(4829)));
    layer1_outputs(1747) <= not(layer0_outputs(2368)) or (layer0_outputs(2200));
    layer1_outputs(1748) <= not(layer0_outputs(392));
    layer1_outputs(1749) <= not(layer0_outputs(3993)) or (layer0_outputs(911));
    layer1_outputs(1750) <= not(layer0_outputs(4126));
    layer1_outputs(1751) <= not(layer0_outputs(2599)) or (layer0_outputs(1924));
    layer1_outputs(1752) <= layer0_outputs(1029);
    layer1_outputs(1753) <= (layer0_outputs(3974)) xor (layer0_outputs(1844));
    layer1_outputs(1754) <= not(layer0_outputs(1104));
    layer1_outputs(1755) <= not((layer0_outputs(1758)) and (layer0_outputs(2977)));
    layer1_outputs(1756) <= not(layer0_outputs(1287)) or (layer0_outputs(2482));
    layer1_outputs(1757) <= not((layer0_outputs(3674)) and (layer0_outputs(2876)));
    layer1_outputs(1758) <= not((layer0_outputs(2736)) or (layer0_outputs(4200)));
    layer1_outputs(1759) <= layer0_outputs(3166);
    layer1_outputs(1760) <= not((layer0_outputs(2612)) xor (layer0_outputs(345)));
    layer1_outputs(1761) <= not(layer0_outputs(2479)) or (layer0_outputs(856));
    layer1_outputs(1762) <= (layer0_outputs(4997)) and not (layer0_outputs(3501));
    layer1_outputs(1763) <= (layer0_outputs(906)) or (layer0_outputs(4356));
    layer1_outputs(1764) <= layer0_outputs(1557);
    layer1_outputs(1765) <= (layer0_outputs(987)) and not (layer0_outputs(1042));
    layer1_outputs(1766) <= layer0_outputs(2960);
    layer1_outputs(1767) <= (layer0_outputs(4850)) or (layer0_outputs(2798));
    layer1_outputs(1768) <= not((layer0_outputs(3959)) or (layer0_outputs(2932)));
    layer1_outputs(1769) <= layer0_outputs(420);
    layer1_outputs(1770) <= not((layer0_outputs(4402)) or (layer0_outputs(4193)));
    layer1_outputs(1771) <= layer0_outputs(1139);
    layer1_outputs(1772) <= layer0_outputs(1838);
    layer1_outputs(1773) <= '1';
    layer1_outputs(1774) <= not(layer0_outputs(3355)) or (layer0_outputs(4383));
    layer1_outputs(1775) <= layer0_outputs(1799);
    layer1_outputs(1776) <= (layer0_outputs(1560)) and not (layer0_outputs(3023));
    layer1_outputs(1777) <= layer0_outputs(4206);
    layer1_outputs(1778) <= layer0_outputs(4204);
    layer1_outputs(1779) <= not(layer0_outputs(2248)) or (layer0_outputs(698));
    layer1_outputs(1780) <= (layer0_outputs(3042)) or (layer0_outputs(4501));
    layer1_outputs(1781) <= layer0_outputs(3995);
    layer1_outputs(1782) <= not(layer0_outputs(3838));
    layer1_outputs(1783) <= not(layer0_outputs(2793));
    layer1_outputs(1784) <= not(layer0_outputs(1116));
    layer1_outputs(1785) <= not((layer0_outputs(3747)) and (layer0_outputs(4953)));
    layer1_outputs(1786) <= not((layer0_outputs(4901)) and (layer0_outputs(411)));
    layer1_outputs(1787) <= (layer0_outputs(1016)) and (layer0_outputs(4182));
    layer1_outputs(1788) <= layer0_outputs(4908);
    layer1_outputs(1789) <= layer0_outputs(489);
    layer1_outputs(1790) <= layer0_outputs(3970);
    layer1_outputs(1791) <= (layer0_outputs(3457)) and (layer0_outputs(4148));
    layer1_outputs(1792) <= not(layer0_outputs(4168));
    layer1_outputs(1793) <= (layer0_outputs(4042)) or (layer0_outputs(3834));
    layer1_outputs(1794) <= layer0_outputs(1543);
    layer1_outputs(1795) <= not(layer0_outputs(2920)) or (layer0_outputs(2898));
    layer1_outputs(1796) <= not(layer0_outputs(621));
    layer1_outputs(1797) <= not(layer0_outputs(2507));
    layer1_outputs(1798) <= (layer0_outputs(5020)) and not (layer0_outputs(2602));
    layer1_outputs(1799) <= layer0_outputs(2376);
    layer1_outputs(1800) <= (layer0_outputs(3881)) and not (layer0_outputs(4061));
    layer1_outputs(1801) <= layer0_outputs(3809);
    layer1_outputs(1802) <= not(layer0_outputs(3517)) or (layer0_outputs(1122));
    layer1_outputs(1803) <= not(layer0_outputs(2980));
    layer1_outputs(1804) <= '0';
    layer1_outputs(1805) <= not(layer0_outputs(3199)) or (layer0_outputs(3240));
    layer1_outputs(1806) <= not((layer0_outputs(2327)) xor (layer0_outputs(4120)));
    layer1_outputs(1807) <= (layer0_outputs(434)) xor (layer0_outputs(4234));
    layer1_outputs(1808) <= not(layer0_outputs(950)) or (layer0_outputs(116));
    layer1_outputs(1809) <= not(layer0_outputs(3536)) or (layer0_outputs(3898));
    layer1_outputs(1810) <= layer0_outputs(3371);
    layer1_outputs(1811) <= layer0_outputs(2535);
    layer1_outputs(1812) <= not(layer0_outputs(5118)) or (layer0_outputs(2386));
    layer1_outputs(1813) <= not((layer0_outputs(334)) or (layer0_outputs(1994)));
    layer1_outputs(1814) <= not(layer0_outputs(1112)) or (layer0_outputs(1605));
    layer1_outputs(1815) <= layer0_outputs(1482);
    layer1_outputs(1816) <= (layer0_outputs(1771)) and not (layer0_outputs(397));
    layer1_outputs(1817) <= (layer0_outputs(2069)) and not (layer0_outputs(55));
    layer1_outputs(1818) <= layer0_outputs(223);
    layer1_outputs(1819) <= layer0_outputs(4114);
    layer1_outputs(1820) <= not(layer0_outputs(3278));
    layer1_outputs(1821) <= layer0_outputs(1741);
    layer1_outputs(1822) <= (layer0_outputs(2035)) and not (layer0_outputs(2669));
    layer1_outputs(1823) <= not((layer0_outputs(1242)) and (layer0_outputs(2077)));
    layer1_outputs(1824) <= (layer0_outputs(4152)) or (layer0_outputs(3740));
    layer1_outputs(1825) <= not(layer0_outputs(2624));
    layer1_outputs(1826) <= layer0_outputs(2500);
    layer1_outputs(1827) <= layer0_outputs(393);
    layer1_outputs(1828) <= layer0_outputs(2028);
    layer1_outputs(1829) <= not(layer0_outputs(2420));
    layer1_outputs(1830) <= (layer0_outputs(3147)) or (layer0_outputs(3257));
    layer1_outputs(1831) <= not((layer0_outputs(3734)) or (layer0_outputs(3698)));
    layer1_outputs(1832) <= not((layer0_outputs(1314)) or (layer0_outputs(710)));
    layer1_outputs(1833) <= layer0_outputs(1754);
    layer1_outputs(1834) <= (layer0_outputs(640)) and (layer0_outputs(3308));
    layer1_outputs(1835) <= (layer0_outputs(230)) and not (layer0_outputs(4725));
    layer1_outputs(1836) <= (layer0_outputs(1828)) and (layer0_outputs(1798));
    layer1_outputs(1837) <= (layer0_outputs(836)) and not (layer0_outputs(3782));
    layer1_outputs(1838) <= not(layer0_outputs(1733));
    layer1_outputs(1839) <= not((layer0_outputs(2026)) or (layer0_outputs(1400)));
    layer1_outputs(1840) <= layer0_outputs(655);
    layer1_outputs(1841) <= not(layer0_outputs(2775));
    layer1_outputs(1842) <= not(layer0_outputs(4076));
    layer1_outputs(1843) <= layer0_outputs(153);
    layer1_outputs(1844) <= not(layer0_outputs(12));
    layer1_outputs(1845) <= not(layer0_outputs(4067)) or (layer0_outputs(2862));
    layer1_outputs(1846) <= not((layer0_outputs(4719)) xor (layer0_outputs(3804)));
    layer1_outputs(1847) <= layer0_outputs(941);
    layer1_outputs(1848) <= not((layer0_outputs(2833)) and (layer0_outputs(4664)));
    layer1_outputs(1849) <= layer0_outputs(4098);
    layer1_outputs(1850) <= '0';
    layer1_outputs(1851) <= layer0_outputs(1460);
    layer1_outputs(1852) <= not((layer0_outputs(4501)) and (layer0_outputs(4821)));
    layer1_outputs(1853) <= (layer0_outputs(1016)) and not (layer0_outputs(4849));
    layer1_outputs(1854) <= layer0_outputs(4860);
    layer1_outputs(1855) <= (layer0_outputs(824)) and not (layer0_outputs(1516));
    layer1_outputs(1856) <= (layer0_outputs(3497)) and (layer0_outputs(549));
    layer1_outputs(1857) <= not(layer0_outputs(593)) or (layer0_outputs(4776));
    layer1_outputs(1858) <= not(layer0_outputs(2301));
    layer1_outputs(1859) <= layer0_outputs(4928);
    layer1_outputs(1860) <= layer0_outputs(1235);
    layer1_outputs(1861) <= (layer0_outputs(4199)) xor (layer0_outputs(465));
    layer1_outputs(1862) <= (layer0_outputs(1261)) or (layer0_outputs(3291));
    layer1_outputs(1863) <= not(layer0_outputs(41));
    layer1_outputs(1864) <= not(layer0_outputs(4864)) or (layer0_outputs(3267));
    layer1_outputs(1865) <= not(layer0_outputs(361)) or (layer0_outputs(752));
    layer1_outputs(1866) <= (layer0_outputs(1617)) and not (layer0_outputs(1124));
    layer1_outputs(1867) <= layer0_outputs(2950);
    layer1_outputs(1868) <= not((layer0_outputs(4975)) and (layer0_outputs(2485)));
    layer1_outputs(1869) <= '1';
    layer1_outputs(1870) <= (layer0_outputs(1714)) and not (layer0_outputs(3186));
    layer1_outputs(1871) <= (layer0_outputs(1378)) or (layer0_outputs(3091));
    layer1_outputs(1872) <= layer0_outputs(1713);
    layer1_outputs(1873) <= layer0_outputs(1352);
    layer1_outputs(1874) <= not(layer0_outputs(3108)) or (layer0_outputs(1792));
    layer1_outputs(1875) <= not(layer0_outputs(1976));
    layer1_outputs(1876) <= layer0_outputs(3065);
    layer1_outputs(1877) <= not(layer0_outputs(542)) or (layer0_outputs(743));
    layer1_outputs(1878) <= not(layer0_outputs(1239));
    layer1_outputs(1879) <= '1';
    layer1_outputs(1880) <= (layer0_outputs(4893)) and not (layer0_outputs(3247));
    layer1_outputs(1881) <= (layer0_outputs(2006)) xor (layer0_outputs(2981));
    layer1_outputs(1882) <= layer0_outputs(4452);
    layer1_outputs(1883) <= not(layer0_outputs(1396));
    layer1_outputs(1884) <= not((layer0_outputs(1177)) and (layer0_outputs(2042)));
    layer1_outputs(1885) <= (layer0_outputs(4538)) or (layer0_outputs(1271));
    layer1_outputs(1886) <= layer0_outputs(3867);
    layer1_outputs(1887) <= not(layer0_outputs(2184)) or (layer0_outputs(28));
    layer1_outputs(1888) <= not((layer0_outputs(2019)) and (layer0_outputs(3692)));
    layer1_outputs(1889) <= layer0_outputs(4244);
    layer1_outputs(1890) <= not(layer0_outputs(2098));
    layer1_outputs(1891) <= not(layer0_outputs(2948)) or (layer0_outputs(5037));
    layer1_outputs(1892) <= layer0_outputs(1944);
    layer1_outputs(1893) <= (layer0_outputs(2890)) and not (layer0_outputs(3521));
    layer1_outputs(1894) <= not(layer0_outputs(2560)) or (layer0_outputs(4130));
    layer1_outputs(1895) <= layer0_outputs(1174);
    layer1_outputs(1896) <= (layer0_outputs(3584)) xor (layer0_outputs(3764));
    layer1_outputs(1897) <= not((layer0_outputs(4279)) and (layer0_outputs(3342)));
    layer1_outputs(1898) <= (layer0_outputs(1265)) and (layer0_outputs(5085));
    layer1_outputs(1899) <= layer0_outputs(3283);
    layer1_outputs(1900) <= not(layer0_outputs(2658));
    layer1_outputs(1901) <= not(layer0_outputs(1308));
    layer1_outputs(1902) <= not(layer0_outputs(3464));
    layer1_outputs(1903) <= layer0_outputs(3237);
    layer1_outputs(1904) <= layer0_outputs(1331);
    layer1_outputs(1905) <= not(layer0_outputs(1190));
    layer1_outputs(1906) <= (layer0_outputs(4106)) or (layer0_outputs(2373));
    layer1_outputs(1907) <= not(layer0_outputs(3155)) or (layer0_outputs(1129));
    layer1_outputs(1908) <= not(layer0_outputs(2966)) or (layer0_outputs(973));
    layer1_outputs(1909) <= not((layer0_outputs(1300)) and (layer0_outputs(976)));
    layer1_outputs(1910) <= layer0_outputs(1480);
    layer1_outputs(1911) <= not((layer0_outputs(2383)) and (layer0_outputs(1885)));
    layer1_outputs(1912) <= not((layer0_outputs(2737)) and (layer0_outputs(2119)));
    layer1_outputs(1913) <= layer0_outputs(3478);
    layer1_outputs(1914) <= not((layer0_outputs(3144)) or (layer0_outputs(3136)));
    layer1_outputs(1915) <= not((layer0_outputs(3763)) and (layer0_outputs(1346)));
    layer1_outputs(1916) <= (layer0_outputs(3234)) xor (layer0_outputs(4998));
    layer1_outputs(1917) <= '0';
    layer1_outputs(1918) <= not((layer0_outputs(1027)) xor (layer0_outputs(1788)));
    layer1_outputs(1919) <= (layer0_outputs(979)) and not (layer0_outputs(3204));
    layer1_outputs(1920) <= not(layer0_outputs(1864));
    layer1_outputs(1921) <= not(layer0_outputs(3296)) or (layer0_outputs(3909));
    layer1_outputs(1922) <= not(layer0_outputs(1599));
    layer1_outputs(1923) <= layer0_outputs(991);
    layer1_outputs(1924) <= not((layer0_outputs(2844)) and (layer0_outputs(2976)));
    layer1_outputs(1925) <= (layer0_outputs(3827)) or (layer0_outputs(528));
    layer1_outputs(1926) <= layer0_outputs(3124);
    layer1_outputs(1927) <= not((layer0_outputs(3159)) and (layer0_outputs(5110)));
    layer1_outputs(1928) <= (layer0_outputs(2535)) or (layer0_outputs(2915));
    layer1_outputs(1929) <= not(layer0_outputs(4355));
    layer1_outputs(1930) <= (layer0_outputs(3126)) or (layer0_outputs(4903));
    layer1_outputs(1931) <= (layer0_outputs(3227)) or (layer0_outputs(4852));
    layer1_outputs(1932) <= (layer0_outputs(788)) and (layer0_outputs(2118));
    layer1_outputs(1933) <= not(layer0_outputs(3587));
    layer1_outputs(1934) <= not(layer0_outputs(5075));
    layer1_outputs(1935) <= not(layer0_outputs(4085)) or (layer0_outputs(2414));
    layer1_outputs(1936) <= (layer0_outputs(1075)) and (layer0_outputs(941));
    layer1_outputs(1937) <= not(layer0_outputs(3704));
    layer1_outputs(1938) <= (layer0_outputs(933)) and not (layer0_outputs(3020));
    layer1_outputs(1939) <= layer0_outputs(3310);
    layer1_outputs(1940) <= (layer0_outputs(3276)) and (layer0_outputs(3601));
    layer1_outputs(1941) <= (layer0_outputs(867)) or (layer0_outputs(2447));
    layer1_outputs(1942) <= not((layer0_outputs(4936)) and (layer0_outputs(4155)));
    layer1_outputs(1943) <= not((layer0_outputs(4687)) and (layer0_outputs(3)));
    layer1_outputs(1944) <= not((layer0_outputs(1619)) or (layer0_outputs(4025)));
    layer1_outputs(1945) <= not(layer0_outputs(3253));
    layer1_outputs(1946) <= not((layer0_outputs(1554)) and (layer0_outputs(2222)));
    layer1_outputs(1947) <= (layer0_outputs(1331)) and (layer0_outputs(1201));
    layer1_outputs(1948) <= '0';
    layer1_outputs(1949) <= not(layer0_outputs(509)) or (layer0_outputs(52));
    layer1_outputs(1950) <= (layer0_outputs(2955)) xor (layer0_outputs(2875));
    layer1_outputs(1951) <= not(layer0_outputs(2683)) or (layer0_outputs(4505));
    layer1_outputs(1952) <= (layer0_outputs(2028)) and not (layer0_outputs(966));
    layer1_outputs(1953) <= not((layer0_outputs(1605)) xor (layer0_outputs(928)));
    layer1_outputs(1954) <= not((layer0_outputs(2034)) and (layer0_outputs(3359)));
    layer1_outputs(1955) <= (layer0_outputs(1311)) or (layer0_outputs(5060));
    layer1_outputs(1956) <= (layer0_outputs(1855)) xor (layer0_outputs(4445));
    layer1_outputs(1957) <= (layer0_outputs(798)) and not (layer0_outputs(619));
    layer1_outputs(1958) <= not(layer0_outputs(1806));
    layer1_outputs(1959) <= layer0_outputs(2370);
    layer1_outputs(1960) <= layer0_outputs(305);
    layer1_outputs(1961) <= not((layer0_outputs(2680)) xor (layer0_outputs(2382)));
    layer1_outputs(1962) <= (layer0_outputs(3245)) or (layer0_outputs(3715));
    layer1_outputs(1963) <= not(layer0_outputs(3089)) or (layer0_outputs(4828));
    layer1_outputs(1964) <= layer0_outputs(2681);
    layer1_outputs(1965) <= not(layer0_outputs(268));
    layer1_outputs(1966) <= (layer0_outputs(1173)) and (layer0_outputs(227));
    layer1_outputs(1967) <= (layer0_outputs(3106)) and not (layer0_outputs(3553));
    layer1_outputs(1968) <= (layer0_outputs(1425)) and not (layer0_outputs(415));
    layer1_outputs(1969) <= not(layer0_outputs(4337)) or (layer0_outputs(2443));
    layer1_outputs(1970) <= (layer0_outputs(87)) xor (layer0_outputs(19));
    layer1_outputs(1971) <= not((layer0_outputs(3271)) or (layer0_outputs(3602)));
    layer1_outputs(1972) <= not((layer0_outputs(4181)) or (layer0_outputs(429)));
    layer1_outputs(1973) <= not(layer0_outputs(931));
    layer1_outputs(1974) <= (layer0_outputs(1144)) and (layer0_outputs(2764));
    layer1_outputs(1975) <= (layer0_outputs(2534)) or (layer0_outputs(1212));
    layer1_outputs(1976) <= not((layer0_outputs(4938)) and (layer0_outputs(266)));
    layer1_outputs(1977) <= layer0_outputs(3189);
    layer1_outputs(1978) <= layer0_outputs(4891);
    layer1_outputs(1979) <= (layer0_outputs(1279)) xor (layer0_outputs(2962));
    layer1_outputs(1980) <= not((layer0_outputs(2986)) xor (layer0_outputs(3925)));
    layer1_outputs(1981) <= (layer0_outputs(1516)) xor (layer0_outputs(4329));
    layer1_outputs(1982) <= layer0_outputs(2411);
    layer1_outputs(1983) <= layer0_outputs(984);
    layer1_outputs(1984) <= (layer0_outputs(3553)) xor (layer0_outputs(4409));
    layer1_outputs(1985) <= layer0_outputs(3127);
    layer1_outputs(1986) <= '1';
    layer1_outputs(1987) <= not(layer0_outputs(4246)) or (layer0_outputs(2779));
    layer1_outputs(1988) <= (layer0_outputs(1332)) and not (layer0_outputs(495));
    layer1_outputs(1989) <= layer0_outputs(2755);
    layer1_outputs(1990) <= not(layer0_outputs(1957)) or (layer0_outputs(3481));
    layer1_outputs(1991) <= (layer0_outputs(4794)) and not (layer0_outputs(2487));
    layer1_outputs(1992) <= (layer0_outputs(3013)) xor (layer0_outputs(1167));
    layer1_outputs(1993) <= '0';
    layer1_outputs(1994) <= not((layer0_outputs(4137)) xor (layer0_outputs(3887)));
    layer1_outputs(1995) <= (layer0_outputs(739)) and not (layer0_outputs(897));
    layer1_outputs(1996) <= layer0_outputs(1249);
    layer1_outputs(1997) <= (layer0_outputs(2625)) and not (layer0_outputs(2025));
    layer1_outputs(1998) <= not((layer0_outputs(4060)) and (layer0_outputs(1768)));
    layer1_outputs(1999) <= '1';
    layer1_outputs(2000) <= (layer0_outputs(2058)) and not (layer0_outputs(2861));
    layer1_outputs(2001) <= not(layer0_outputs(1008));
    layer1_outputs(2002) <= (layer0_outputs(365)) or (layer0_outputs(756));
    layer1_outputs(2003) <= (layer0_outputs(1859)) and not (layer0_outputs(2471));
    layer1_outputs(2004) <= (layer0_outputs(192)) or (layer0_outputs(4414));
    layer1_outputs(2005) <= not(layer0_outputs(4784)) or (layer0_outputs(3240));
    layer1_outputs(2006) <= not((layer0_outputs(1384)) and (layer0_outputs(229)));
    layer1_outputs(2007) <= not((layer0_outputs(4970)) xor (layer0_outputs(2544)));
    layer1_outputs(2008) <= layer0_outputs(4117);
    layer1_outputs(2009) <= (layer0_outputs(3301)) and not (layer0_outputs(2258));
    layer1_outputs(2010) <= not((layer0_outputs(131)) or (layer0_outputs(691)));
    layer1_outputs(2011) <= not((layer0_outputs(2878)) xor (layer0_outputs(4341)));
    layer1_outputs(2012) <= (layer0_outputs(1530)) and not (layer0_outputs(4177));
    layer1_outputs(2013) <= '0';
    layer1_outputs(2014) <= not(layer0_outputs(1511));
    layer1_outputs(2015) <= (layer0_outputs(1203)) xor (layer0_outputs(2355));
    layer1_outputs(2016) <= (layer0_outputs(2540)) and not (layer0_outputs(2068));
    layer1_outputs(2017) <= (layer0_outputs(557)) and (layer0_outputs(607));
    layer1_outputs(2018) <= layer0_outputs(1981);
    layer1_outputs(2019) <= not(layer0_outputs(1965));
    layer1_outputs(2020) <= (layer0_outputs(461)) and (layer0_outputs(615));
    layer1_outputs(2021) <= not(layer0_outputs(2914));
    layer1_outputs(2022) <= '0';
    layer1_outputs(2023) <= (layer0_outputs(603)) and (layer0_outputs(2550));
    layer1_outputs(2024) <= (layer0_outputs(3786)) and (layer0_outputs(450));
    layer1_outputs(2025) <= (layer0_outputs(738)) and not (layer0_outputs(2347));
    layer1_outputs(2026) <= layer0_outputs(1125);
    layer1_outputs(2027) <= not((layer0_outputs(2348)) xor (layer0_outputs(1291)));
    layer1_outputs(2028) <= (layer0_outputs(4524)) and not (layer0_outputs(4202));
    layer1_outputs(2029) <= not((layer0_outputs(2437)) or (layer0_outputs(3585)));
    layer1_outputs(2030) <= (layer0_outputs(1638)) or (layer0_outputs(1216));
    layer1_outputs(2031) <= (layer0_outputs(2426)) xor (layer0_outputs(2810));
    layer1_outputs(2032) <= layer0_outputs(963);
    layer1_outputs(2033) <= (layer0_outputs(4062)) and not (layer0_outputs(4759));
    layer1_outputs(2034) <= not(layer0_outputs(1536));
    layer1_outputs(2035) <= (layer0_outputs(1613)) or (layer0_outputs(5027));
    layer1_outputs(2036) <= not(layer0_outputs(2201));
    layer1_outputs(2037) <= (layer0_outputs(3905)) and (layer0_outputs(2938));
    layer1_outputs(2038) <= (layer0_outputs(3152)) or (layer0_outputs(198));
    layer1_outputs(2039) <= not((layer0_outputs(3387)) and (layer0_outputs(84)));
    layer1_outputs(2040) <= '0';
    layer1_outputs(2041) <= (layer0_outputs(2850)) or (layer0_outputs(5035));
    layer1_outputs(2042) <= layer0_outputs(799);
    layer1_outputs(2043) <= not((layer0_outputs(2133)) and (layer0_outputs(1422)));
    layer1_outputs(2044) <= not(layer0_outputs(565)) or (layer0_outputs(1443));
    layer1_outputs(2045) <= not((layer0_outputs(1970)) xor (layer0_outputs(51)));
    layer1_outputs(2046) <= not(layer0_outputs(206));
    layer1_outputs(2047) <= (layer0_outputs(4885)) and not (layer0_outputs(3879));
    layer1_outputs(2048) <= not(layer0_outputs(4270)) or (layer0_outputs(1879));
    layer1_outputs(2049) <= not(layer0_outputs(3810));
    layer1_outputs(2050) <= not(layer0_outputs(27));
    layer1_outputs(2051) <= not(layer0_outputs(4247));
    layer1_outputs(2052) <= layer0_outputs(4798);
    layer1_outputs(2053) <= not(layer0_outputs(3030));
    layer1_outputs(2054) <= not(layer0_outputs(1755));
    layer1_outputs(2055) <= '1';
    layer1_outputs(2056) <= layer0_outputs(1105);
    layer1_outputs(2057) <= (layer0_outputs(1191)) and not (layer0_outputs(4927));
    layer1_outputs(2058) <= (layer0_outputs(3885)) or (layer0_outputs(186));
    layer1_outputs(2059) <= not(layer0_outputs(4717));
    layer1_outputs(2060) <= layer0_outputs(4400);
    layer1_outputs(2061) <= not((layer0_outputs(1429)) and (layer0_outputs(1214)));
    layer1_outputs(2062) <= (layer0_outputs(760)) and (layer0_outputs(1037));
    layer1_outputs(2063) <= not(layer0_outputs(2094));
    layer1_outputs(2064) <= layer0_outputs(4112);
    layer1_outputs(2065) <= (layer0_outputs(3884)) or (layer0_outputs(3402));
    layer1_outputs(2066) <= not((layer0_outputs(4679)) xor (layer0_outputs(4147)));
    layer1_outputs(2067) <= not(layer0_outputs(1416));
    layer1_outputs(2068) <= not((layer0_outputs(2821)) and (layer0_outputs(2230)));
    layer1_outputs(2069) <= not(layer0_outputs(3393)) or (layer0_outputs(780));
    layer1_outputs(2070) <= (layer0_outputs(2805)) and not (layer0_outputs(2312));
    layer1_outputs(2071) <= not((layer0_outputs(2411)) or (layer0_outputs(4549)));
    layer1_outputs(2072) <= '1';
    layer1_outputs(2073) <= not((layer0_outputs(4242)) or (layer0_outputs(3690)));
    layer1_outputs(2074) <= not(layer0_outputs(4463));
    layer1_outputs(2075) <= not(layer0_outputs(578));
    layer1_outputs(2076) <= not(layer0_outputs(126));
    layer1_outputs(2077) <= (layer0_outputs(3370)) or (layer0_outputs(3641));
    layer1_outputs(2078) <= (layer0_outputs(1088)) xor (layer0_outputs(2267));
    layer1_outputs(2079) <= (layer0_outputs(4872)) and (layer0_outputs(1588));
    layer1_outputs(2080) <= (layer0_outputs(1131)) and not (layer0_outputs(4857));
    layer1_outputs(2081) <= not(layer0_outputs(3591));
    layer1_outputs(2082) <= (layer0_outputs(803)) and not (layer0_outputs(4567));
    layer1_outputs(2083) <= not(layer0_outputs(3132));
    layer1_outputs(2084) <= (layer0_outputs(1680)) or (layer0_outputs(1344));
    layer1_outputs(2085) <= (layer0_outputs(3253)) or (layer0_outputs(4917));
    layer1_outputs(2086) <= (layer0_outputs(2908)) or (layer0_outputs(4892));
    layer1_outputs(2087) <= not(layer0_outputs(1905)) or (layer0_outputs(721));
    layer1_outputs(2088) <= '0';
    layer1_outputs(2089) <= not((layer0_outputs(3145)) or (layer0_outputs(4192)));
    layer1_outputs(2090) <= (layer0_outputs(2293)) and not (layer0_outputs(3317));
    layer1_outputs(2091) <= (layer0_outputs(1338)) and not (layer0_outputs(5101));
    layer1_outputs(2092) <= (layer0_outputs(352)) and (layer0_outputs(348));
    layer1_outputs(2093) <= not(layer0_outputs(1050));
    layer1_outputs(2094) <= not(layer0_outputs(3255));
    layer1_outputs(2095) <= layer0_outputs(4935);
    layer1_outputs(2096) <= not(layer0_outputs(1499)) or (layer0_outputs(2132));
    layer1_outputs(2097) <= (layer0_outputs(2890)) and (layer0_outputs(683));
    layer1_outputs(2098) <= not((layer0_outputs(865)) or (layer0_outputs(1229)));
    layer1_outputs(2099) <= (layer0_outputs(3108)) and (layer0_outputs(3081));
    layer1_outputs(2100) <= not(layer0_outputs(1329));
    layer1_outputs(2101) <= layer0_outputs(120);
    layer1_outputs(2102) <= not((layer0_outputs(3559)) and (layer0_outputs(1428)));
    layer1_outputs(2103) <= (layer0_outputs(2254)) or (layer0_outputs(1469));
    layer1_outputs(2104) <= not(layer0_outputs(3465));
    layer1_outputs(2105) <= not((layer0_outputs(3401)) and (layer0_outputs(4486)));
    layer1_outputs(2106) <= (layer0_outputs(2739)) and not (layer0_outputs(2867));
    layer1_outputs(2107) <= (layer0_outputs(1277)) xor (layer0_outputs(3876));
    layer1_outputs(2108) <= (layer0_outputs(4174)) and not (layer0_outputs(424));
    layer1_outputs(2109) <= (layer0_outputs(1670)) xor (layer0_outputs(4559));
    layer1_outputs(2110) <= '0';
    layer1_outputs(2111) <= (layer0_outputs(2016)) and not (layer0_outputs(1688));
    layer1_outputs(2112) <= layer0_outputs(2608);
    layer1_outputs(2113) <= (layer0_outputs(4558)) and (layer0_outputs(1684));
    layer1_outputs(2114) <= not((layer0_outputs(1599)) and (layer0_outputs(4314)));
    layer1_outputs(2115) <= not(layer0_outputs(3857));
    layer1_outputs(2116) <= layer0_outputs(1749);
    layer1_outputs(2117) <= not(layer0_outputs(4138)) or (layer0_outputs(324));
    layer1_outputs(2118) <= not(layer0_outputs(4336)) or (layer0_outputs(2196));
    layer1_outputs(2119) <= (layer0_outputs(113)) or (layer0_outputs(2995));
    layer1_outputs(2120) <= (layer0_outputs(3030)) and (layer0_outputs(4659));
    layer1_outputs(2121) <= (layer0_outputs(3536)) and not (layer0_outputs(207));
    layer1_outputs(2122) <= not((layer0_outputs(4297)) and (layer0_outputs(3027)));
    layer1_outputs(2123) <= not(layer0_outputs(1963));
    layer1_outputs(2124) <= layer0_outputs(2231);
    layer1_outputs(2125) <= not((layer0_outputs(3424)) and (layer0_outputs(3317)));
    layer1_outputs(2126) <= not((layer0_outputs(339)) xor (layer0_outputs(77)));
    layer1_outputs(2127) <= not((layer0_outputs(2924)) or (layer0_outputs(2530)));
    layer1_outputs(2128) <= not((layer0_outputs(4986)) xor (layer0_outputs(572)));
    layer1_outputs(2129) <= (layer0_outputs(1050)) or (layer0_outputs(1176));
    layer1_outputs(2130) <= (layer0_outputs(1931)) and not (layer0_outputs(3531));
    layer1_outputs(2131) <= not((layer0_outputs(2340)) xor (layer0_outputs(3275)));
    layer1_outputs(2132) <= not(layer0_outputs(2489));
    layer1_outputs(2133) <= not(layer0_outputs(3300)) or (layer0_outputs(2667));
    layer1_outputs(2134) <= not(layer0_outputs(2533));
    layer1_outputs(2135) <= (layer0_outputs(1241)) xor (layer0_outputs(2889));
    layer1_outputs(2136) <= (layer0_outputs(599)) and (layer0_outputs(4593));
    layer1_outputs(2137) <= not(layer0_outputs(280)) or (layer0_outputs(1252));
    layer1_outputs(2138) <= not(layer0_outputs(375)) or (layer0_outputs(3266));
    layer1_outputs(2139) <= layer0_outputs(3049);
    layer1_outputs(2140) <= (layer0_outputs(2521)) xor (layer0_outputs(4863));
    layer1_outputs(2141) <= (layer0_outputs(2546)) and not (layer0_outputs(2563));
    layer1_outputs(2142) <= layer0_outputs(4703);
    layer1_outputs(2143) <= not((layer0_outputs(2834)) and (layer0_outputs(5084)));
    layer1_outputs(2144) <= not(layer0_outputs(716));
    layer1_outputs(2145) <= (layer0_outputs(1587)) and (layer0_outputs(531));
    layer1_outputs(2146) <= not(layer0_outputs(2945));
    layer1_outputs(2147) <= not(layer0_outputs(1827));
    layer1_outputs(2148) <= (layer0_outputs(544)) and not (layer0_outputs(1393));
    layer1_outputs(2149) <= not((layer0_outputs(4297)) xor (layer0_outputs(3566)));
    layer1_outputs(2150) <= (layer0_outputs(307)) or (layer0_outputs(3542));
    layer1_outputs(2151) <= not((layer0_outputs(4981)) and (layer0_outputs(3333)));
    layer1_outputs(2152) <= (layer0_outputs(4499)) and not (layer0_outputs(2839));
    layer1_outputs(2153) <= (layer0_outputs(3321)) or (layer0_outputs(1623));
    layer1_outputs(2154) <= (layer0_outputs(3201)) and not (layer0_outputs(122));
    layer1_outputs(2155) <= (layer0_outputs(1551)) or (layer0_outputs(1789));
    layer1_outputs(2156) <= layer0_outputs(1986);
    layer1_outputs(2157) <= not((layer0_outputs(3756)) and (layer0_outputs(2433)));
    layer1_outputs(2158) <= '1';
    layer1_outputs(2159) <= not(layer0_outputs(507));
    layer1_outputs(2160) <= layer0_outputs(129);
    layer1_outputs(2161) <= (layer0_outputs(3911)) or (layer0_outputs(3589));
    layer1_outputs(2162) <= not(layer0_outputs(2868)) or (layer0_outputs(4915));
    layer1_outputs(2163) <= not(layer0_outputs(3005));
    layer1_outputs(2164) <= (layer0_outputs(1403)) and not (layer0_outputs(1382));
    layer1_outputs(2165) <= (layer0_outputs(3277)) or (layer0_outputs(4427));
    layer1_outputs(2166) <= (layer0_outputs(2824)) or (layer0_outputs(2772));
    layer1_outputs(2167) <= not((layer0_outputs(2105)) or (layer0_outputs(328)));
    layer1_outputs(2168) <= (layer0_outputs(1787)) xor (layer0_outputs(1797));
    layer1_outputs(2169) <= (layer0_outputs(1001)) and not (layer0_outputs(3520));
    layer1_outputs(2170) <= (layer0_outputs(2857)) and (layer0_outputs(5114));
    layer1_outputs(2171) <= (layer0_outputs(3533)) and not (layer0_outputs(4612));
    layer1_outputs(2172) <= not((layer0_outputs(42)) or (layer0_outputs(4610)));
    layer1_outputs(2173) <= (layer0_outputs(2170)) or (layer0_outputs(874));
    layer1_outputs(2174) <= not((layer0_outputs(4358)) and (layer0_outputs(4698)));
    layer1_outputs(2175) <= (layer0_outputs(733)) or (layer0_outputs(3903));
    layer1_outputs(2176) <= not(layer0_outputs(2539));
    layer1_outputs(2177) <= not(layer0_outputs(2799));
    layer1_outputs(2178) <= not(layer0_outputs(4256)) or (layer0_outputs(540));
    layer1_outputs(2179) <= not((layer0_outputs(4059)) and (layer0_outputs(4672)));
    layer1_outputs(2180) <= not(layer0_outputs(2471));
    layer1_outputs(2181) <= (layer0_outputs(377)) and not (layer0_outputs(1192));
    layer1_outputs(2182) <= '0';
    layer1_outputs(2183) <= not(layer0_outputs(4455));
    layer1_outputs(2184) <= not(layer0_outputs(4668)) or (layer0_outputs(3938));
    layer1_outputs(2185) <= (layer0_outputs(2422)) xor (layer0_outputs(1355));
    layer1_outputs(2186) <= layer0_outputs(869);
    layer1_outputs(2187) <= layer0_outputs(468);
    layer1_outputs(2188) <= not(layer0_outputs(1321));
    layer1_outputs(2189) <= (layer0_outputs(1268)) and not (layer0_outputs(1996));
    layer1_outputs(2190) <= not((layer0_outputs(1903)) and (layer0_outputs(1245)));
    layer1_outputs(2191) <= (layer0_outputs(1660)) and not (layer0_outputs(5042));
    layer1_outputs(2192) <= not((layer0_outputs(163)) and (layer0_outputs(2721)));
    layer1_outputs(2193) <= not(layer0_outputs(3034)) or (layer0_outputs(3043));
    layer1_outputs(2194) <= not(layer0_outputs(69)) or (layer0_outputs(919));
    layer1_outputs(2195) <= not((layer0_outputs(583)) xor (layer0_outputs(4564)));
    layer1_outputs(2196) <= not((layer0_outputs(3384)) and (layer0_outputs(2716)));
    layer1_outputs(2197) <= layer0_outputs(507);
    layer1_outputs(2198) <= (layer0_outputs(1501)) and not (layer0_outputs(2389));
    layer1_outputs(2199) <= not(layer0_outputs(932));
    layer1_outputs(2200) <= not((layer0_outputs(1406)) and (layer0_outputs(2973)));
    layer1_outputs(2201) <= not(layer0_outputs(21)) or (layer0_outputs(211));
    layer1_outputs(2202) <= (layer0_outputs(2080)) xor (layer0_outputs(1540));
    layer1_outputs(2203) <= not(layer0_outputs(3303)) or (layer0_outputs(1588));
    layer1_outputs(2204) <= (layer0_outputs(3586)) or (layer0_outputs(3842));
    layer1_outputs(2205) <= not((layer0_outputs(142)) or (layer0_outputs(1203)));
    layer1_outputs(2206) <= not(layer0_outputs(3796)) or (layer0_outputs(4288));
    layer1_outputs(2207) <= not(layer0_outputs(3784));
    layer1_outputs(2208) <= layer0_outputs(2343);
    layer1_outputs(2209) <= not(layer0_outputs(1669)) or (layer0_outputs(3612));
    layer1_outputs(2210) <= layer0_outputs(3438);
    layer1_outputs(2211) <= not((layer0_outputs(2988)) or (layer0_outputs(823)));
    layer1_outputs(2212) <= layer0_outputs(2043);
    layer1_outputs(2213) <= layer0_outputs(2500);
    layer1_outputs(2214) <= not(layer0_outputs(396));
    layer1_outputs(2215) <= not(layer0_outputs(4803));
    layer1_outputs(2216) <= not(layer0_outputs(3736));
    layer1_outputs(2217) <= layer0_outputs(3852);
    layer1_outputs(2218) <= not((layer0_outputs(3943)) xor (layer0_outputs(3572)));
    layer1_outputs(2219) <= not(layer0_outputs(3662));
    layer1_outputs(2220) <= (layer0_outputs(141)) and not (layer0_outputs(2176));
    layer1_outputs(2221) <= not(layer0_outputs(2001)) or (layer0_outputs(2143));
    layer1_outputs(2222) <= (layer0_outputs(3980)) and (layer0_outputs(3813));
    layer1_outputs(2223) <= layer0_outputs(764);
    layer1_outputs(2224) <= not(layer0_outputs(3195)) or (layer0_outputs(731));
    layer1_outputs(2225) <= layer0_outputs(299);
    layer1_outputs(2226) <= (layer0_outputs(1525)) and not (layer0_outputs(591));
    layer1_outputs(2227) <= (layer0_outputs(2262)) and not (layer0_outputs(5033));
    layer1_outputs(2228) <= (layer0_outputs(3822)) xor (layer0_outputs(1075));
    layer1_outputs(2229) <= not(layer0_outputs(2166));
    layer1_outputs(2230) <= not(layer0_outputs(2371));
    layer1_outputs(2231) <= not(layer0_outputs(3785));
    layer1_outputs(2232) <= layer0_outputs(32);
    layer1_outputs(2233) <= layer0_outputs(1371);
    layer1_outputs(2234) <= not(layer0_outputs(2352)) or (layer0_outputs(2284));
    layer1_outputs(2235) <= not(layer0_outputs(4453));
    layer1_outputs(2236) <= layer0_outputs(5037);
    layer1_outputs(2237) <= (layer0_outputs(2122)) or (layer0_outputs(5108));
    layer1_outputs(2238) <= layer0_outputs(1509);
    layer1_outputs(2239) <= '1';
    layer1_outputs(2240) <= (layer0_outputs(786)) or (layer0_outputs(56));
    layer1_outputs(2241) <= not((layer0_outputs(2911)) and (layer0_outputs(4277)));
    layer1_outputs(2242) <= layer0_outputs(465);
    layer1_outputs(2243) <= (layer0_outputs(3722)) and (layer0_outputs(74));
    layer1_outputs(2244) <= (layer0_outputs(4727)) or (layer0_outputs(427));
    layer1_outputs(2245) <= layer0_outputs(2472);
    layer1_outputs(2246) <= (layer0_outputs(1606)) and not (layer0_outputs(3685));
    layer1_outputs(2247) <= layer0_outputs(2675);
    layer1_outputs(2248) <= (layer0_outputs(4614)) and not (layer0_outputs(5093));
    layer1_outputs(2249) <= not(layer0_outputs(3894));
    layer1_outputs(2250) <= not((layer0_outputs(3567)) or (layer0_outputs(2462)));
    layer1_outputs(2251) <= not(layer0_outputs(2226));
    layer1_outputs(2252) <= not(layer0_outputs(1549));
    layer1_outputs(2253) <= not((layer0_outputs(3557)) or (layer0_outputs(4280)));
    layer1_outputs(2254) <= not(layer0_outputs(723));
    layer1_outputs(2255) <= layer0_outputs(1726);
    layer1_outputs(2256) <= (layer0_outputs(1438)) and not (layer0_outputs(3350));
    layer1_outputs(2257) <= (layer0_outputs(2381)) or (layer0_outputs(4683));
    layer1_outputs(2258) <= (layer0_outputs(179)) or (layer0_outputs(1337));
    layer1_outputs(2259) <= '0';
    layer1_outputs(2260) <= not(layer0_outputs(1453)) or (layer0_outputs(3863));
    layer1_outputs(2261) <= layer0_outputs(157);
    layer1_outputs(2262) <= (layer0_outputs(2273)) or (layer0_outputs(2752));
    layer1_outputs(2263) <= '1';
    layer1_outputs(2264) <= layer0_outputs(2660);
    layer1_outputs(2265) <= (layer0_outputs(1971)) and not (layer0_outputs(1594));
    layer1_outputs(2266) <= layer0_outputs(2637);
    layer1_outputs(2267) <= not((layer0_outputs(709)) xor (layer0_outputs(4888)));
    layer1_outputs(2268) <= (layer0_outputs(4417)) and not (layer0_outputs(4311));
    layer1_outputs(2269) <= layer0_outputs(3607);
    layer1_outputs(2270) <= (layer0_outputs(2469)) and not (layer0_outputs(1841));
    layer1_outputs(2271) <= (layer0_outputs(1091)) xor (layer0_outputs(2855));
    layer1_outputs(2272) <= '0';
    layer1_outputs(2273) <= layer0_outputs(167);
    layer1_outputs(2274) <= (layer0_outputs(1760)) and not (layer0_outputs(1409));
    layer1_outputs(2275) <= not((layer0_outputs(3711)) or (layer0_outputs(193)));
    layer1_outputs(2276) <= not((layer0_outputs(2505)) xor (layer0_outputs(4922)));
    layer1_outputs(2277) <= not((layer0_outputs(4229)) and (layer0_outputs(4400)));
    layer1_outputs(2278) <= layer0_outputs(1076);
    layer1_outputs(2279) <= not((layer0_outputs(4478)) or (layer0_outputs(4761)));
    layer1_outputs(2280) <= not(layer0_outputs(690)) or (layer0_outputs(3174));
    layer1_outputs(2281) <= not((layer0_outputs(2587)) xor (layer0_outputs(2671)));
    layer1_outputs(2282) <= '0';
    layer1_outputs(2283) <= layer0_outputs(970);
    layer1_outputs(2284) <= not((layer0_outputs(1441)) or (layer0_outputs(4172)));
    layer1_outputs(2285) <= not(layer0_outputs(3749));
    layer1_outputs(2286) <= (layer0_outputs(1770)) and not (layer0_outputs(535));
    layer1_outputs(2287) <= '0';
    layer1_outputs(2288) <= not(layer0_outputs(1668));
    layer1_outputs(2289) <= layer0_outputs(2165);
    layer1_outputs(2290) <= (layer0_outputs(3851)) and not (layer0_outputs(2346));
    layer1_outputs(2291) <= not(layer0_outputs(4127)) or (layer0_outputs(1078));
    layer1_outputs(2292) <= (layer0_outputs(3401)) xor (layer0_outputs(2268));
    layer1_outputs(2293) <= not(layer0_outputs(213)) or (layer0_outputs(4178));
    layer1_outputs(2294) <= not(layer0_outputs(3274));
    layer1_outputs(2295) <= not(layer0_outputs(3261)) or (layer0_outputs(4057));
    layer1_outputs(2296) <= not(layer0_outputs(3729));
    layer1_outputs(2297) <= (layer0_outputs(1005)) and not (layer0_outputs(3439));
    layer1_outputs(2298) <= not(layer0_outputs(239));
    layer1_outputs(2299) <= (layer0_outputs(2989)) and not (layer0_outputs(2368));
    layer1_outputs(2300) <= layer0_outputs(1172);
    layer1_outputs(2301) <= not(layer0_outputs(2664));
    layer1_outputs(2302) <= (layer0_outputs(3633)) and not (layer0_outputs(1474));
    layer1_outputs(2303) <= not(layer0_outputs(4980)) or (layer0_outputs(4961));
    layer1_outputs(2304) <= (layer0_outputs(1387)) and (layer0_outputs(4655));
    layer1_outputs(2305) <= (layer0_outputs(4399)) and (layer0_outputs(3044));
    layer1_outputs(2306) <= (layer0_outputs(2563)) and not (layer0_outputs(4651));
    layer1_outputs(2307) <= not(layer0_outputs(1255));
    layer1_outputs(2308) <= not(layer0_outputs(4085));
    layer1_outputs(2309) <= not(layer0_outputs(2148)) or (layer0_outputs(3116));
    layer1_outputs(2310) <= not(layer0_outputs(758)) or (layer0_outputs(4879));
    layer1_outputs(2311) <= (layer0_outputs(1436)) xor (layer0_outputs(2452));
    layer1_outputs(2312) <= layer0_outputs(4135);
    layer1_outputs(2313) <= (layer0_outputs(4104)) xor (layer0_outputs(2416));
    layer1_outputs(2314) <= not((layer0_outputs(3381)) or (layer0_outputs(2597)));
    layer1_outputs(2315) <= not(layer0_outputs(2827)) or (layer0_outputs(1407));
    layer1_outputs(2316) <= layer0_outputs(3927);
    layer1_outputs(2317) <= layer0_outputs(2900);
    layer1_outputs(2318) <= not(layer0_outputs(4270));
    layer1_outputs(2319) <= (layer0_outputs(3222)) xor (layer0_outputs(1036));
    layer1_outputs(2320) <= layer0_outputs(4379);
    layer1_outputs(2321) <= (layer0_outputs(237)) and not (layer0_outputs(5111));
    layer1_outputs(2322) <= not(layer0_outputs(2385));
    layer1_outputs(2323) <= not(layer0_outputs(3523)) or (layer0_outputs(4458));
    layer1_outputs(2324) <= not(layer0_outputs(3249)) or (layer0_outputs(807));
    layer1_outputs(2325) <= layer0_outputs(2311);
    layer1_outputs(2326) <= not(layer0_outputs(4897));
    layer1_outputs(2327) <= '1';
    layer1_outputs(2328) <= (layer0_outputs(3443)) and (layer0_outputs(1790));
    layer1_outputs(2329) <= (layer0_outputs(833)) or (layer0_outputs(4267));
    layer1_outputs(2330) <= not((layer0_outputs(2650)) xor (layer0_outputs(315)));
    layer1_outputs(2331) <= (layer0_outputs(2999)) xor (layer0_outputs(4455));
    layer1_outputs(2332) <= not(layer0_outputs(4291)) or (layer0_outputs(523));
    layer1_outputs(2333) <= not((layer0_outputs(1374)) and (layer0_outputs(872)));
    layer1_outputs(2334) <= not(layer0_outputs(1003));
    layer1_outputs(2335) <= not((layer0_outputs(729)) or (layer0_outputs(4006)));
    layer1_outputs(2336) <= not(layer0_outputs(3268)) or (layer0_outputs(4518));
    layer1_outputs(2337) <= not((layer0_outputs(291)) and (layer0_outputs(178)));
    layer1_outputs(2338) <= not((layer0_outputs(3392)) or (layer0_outputs(3511)));
    layer1_outputs(2339) <= not(layer0_outputs(895));
    layer1_outputs(2340) <= not(layer0_outputs(1065)) or (layer0_outputs(1781));
    layer1_outputs(2341) <= (layer0_outputs(1676)) and (layer0_outputs(5083));
    layer1_outputs(2342) <= not(layer0_outputs(4578));
    layer1_outputs(2343) <= not(layer0_outputs(414));
    layer1_outputs(2344) <= not(layer0_outputs(4778));
    layer1_outputs(2345) <= not((layer0_outputs(4752)) and (layer0_outputs(784)));
    layer1_outputs(2346) <= (layer0_outputs(3229)) or (layer0_outputs(3456));
    layer1_outputs(2347) <= not(layer0_outputs(1598));
    layer1_outputs(2348) <= not(layer0_outputs(4316)) or (layer0_outputs(3083));
    layer1_outputs(2349) <= not(layer0_outputs(3740));
    layer1_outputs(2350) <= layer0_outputs(4694);
    layer1_outputs(2351) <= not((layer0_outputs(140)) or (layer0_outputs(4015)));
    layer1_outputs(2352) <= not((layer0_outputs(813)) or (layer0_outputs(144)));
    layer1_outputs(2353) <= layer0_outputs(3631);
    layer1_outputs(2354) <= not(layer0_outputs(5019));
    layer1_outputs(2355) <= not(layer0_outputs(739));
    layer1_outputs(2356) <= not(layer0_outputs(3852)) or (layer0_outputs(2609));
    layer1_outputs(2357) <= (layer0_outputs(3498)) and not (layer0_outputs(3434));
    layer1_outputs(2358) <= (layer0_outputs(661)) and (layer0_outputs(4255));
    layer1_outputs(2359) <= (layer0_outputs(161)) and not (layer0_outputs(4525));
    layer1_outputs(2360) <= not(layer0_outputs(4369)) or (layer0_outputs(4212));
    layer1_outputs(2361) <= (layer0_outputs(3718)) and (layer0_outputs(2350));
    layer1_outputs(2362) <= '0';
    layer1_outputs(2363) <= (layer0_outputs(115)) or (layer0_outputs(2370));
    layer1_outputs(2364) <= (layer0_outputs(5096)) and not (layer0_outputs(164));
    layer1_outputs(2365) <= not(layer0_outputs(8));
    layer1_outputs(2366) <= not(layer0_outputs(880));
    layer1_outputs(2367) <= layer0_outputs(860);
    layer1_outputs(2368) <= not((layer0_outputs(2979)) and (layer0_outputs(3064)));
    layer1_outputs(2369) <= not(layer0_outputs(339));
    layer1_outputs(2370) <= (layer0_outputs(244)) or (layer0_outputs(3485));
    layer1_outputs(2371) <= not((layer0_outputs(4424)) and (layer0_outputs(1717)));
    layer1_outputs(2372) <= layer0_outputs(613);
    layer1_outputs(2373) <= (layer0_outputs(4301)) and (layer0_outputs(4678));
    layer1_outputs(2374) <= not(layer0_outputs(1781));
    layer1_outputs(2375) <= (layer0_outputs(1877)) and (layer0_outputs(2299));
    layer1_outputs(2376) <= not(layer0_outputs(2212));
    layer1_outputs(2377) <= (layer0_outputs(3404)) and not (layer0_outputs(4040));
    layer1_outputs(2378) <= not((layer0_outputs(63)) xor (layer0_outputs(3323)));
    layer1_outputs(2379) <= not((layer0_outputs(4053)) xor (layer0_outputs(1740)));
    layer1_outputs(2380) <= (layer0_outputs(4328)) and not (layer0_outputs(1659));
    layer1_outputs(2381) <= not(layer0_outputs(5016));
    layer1_outputs(2382) <= layer0_outputs(97);
    layer1_outputs(2383) <= not(layer0_outputs(3630));
    layer1_outputs(2384) <= not((layer0_outputs(4757)) and (layer0_outputs(3987)));
    layer1_outputs(2385) <= not(layer0_outputs(5091));
    layer1_outputs(2386) <= (layer0_outputs(4280)) and not (layer0_outputs(1306));
    layer1_outputs(2387) <= (layer0_outputs(4526)) or (layer0_outputs(1054));
    layer1_outputs(2388) <= not(layer0_outputs(2197));
    layer1_outputs(2389) <= layer0_outputs(3656);
    layer1_outputs(2390) <= (layer0_outputs(3405)) and not (layer0_outputs(2065));
    layer1_outputs(2391) <= not(layer0_outputs(2193));
    layer1_outputs(2392) <= (layer0_outputs(2045)) or (layer0_outputs(1620));
    layer1_outputs(2393) <= (layer0_outputs(1719)) and not (layer0_outputs(4321));
    layer1_outputs(2394) <= not(layer0_outputs(2249));
    layer1_outputs(2395) <= layer0_outputs(4135);
    layer1_outputs(2396) <= layer0_outputs(3671);
    layer1_outputs(2397) <= not(layer0_outputs(2130));
    layer1_outputs(2398) <= not((layer0_outputs(4544)) xor (layer0_outputs(3599)));
    layer1_outputs(2399) <= not(layer0_outputs(4660)) or (layer0_outputs(843));
    layer1_outputs(2400) <= not(layer0_outputs(5017)) or (layer0_outputs(4218));
    layer1_outputs(2401) <= '0';
    layer1_outputs(2402) <= not((layer0_outputs(3711)) and (layer0_outputs(1355)));
    layer1_outputs(2403) <= not(layer0_outputs(4363));
    layer1_outputs(2404) <= (layer0_outputs(125)) or (layer0_outputs(2398));
    layer1_outputs(2405) <= layer0_outputs(404);
    layer1_outputs(2406) <= (layer0_outputs(2333)) and (layer0_outputs(3974));
    layer1_outputs(2407) <= layer0_outputs(1264);
    layer1_outputs(2408) <= not(layer0_outputs(2909));
    layer1_outputs(2409) <= not((layer0_outputs(4511)) and (layer0_outputs(382)));
    layer1_outputs(2410) <= layer0_outputs(2719);
    layer1_outputs(2411) <= not((layer0_outputs(9)) or (layer0_outputs(3527)));
    layer1_outputs(2412) <= not((layer0_outputs(4100)) and (layer0_outputs(4996)));
    layer1_outputs(2413) <= (layer0_outputs(2239)) or (layer0_outputs(3819));
    layer1_outputs(2414) <= (layer0_outputs(1680)) or (layer0_outputs(2421));
    layer1_outputs(2415) <= not(layer0_outputs(2253));
    layer1_outputs(2416) <= not(layer0_outputs(147));
    layer1_outputs(2417) <= (layer0_outputs(5003)) and (layer0_outputs(3096));
    layer1_outputs(2418) <= (layer0_outputs(4832)) and not (layer0_outputs(4723));
    layer1_outputs(2419) <= not(layer0_outputs(3177));
    layer1_outputs(2420) <= (layer0_outputs(4157)) xor (layer0_outputs(3095));
    layer1_outputs(2421) <= '0';
    layer1_outputs(2422) <= not(layer0_outputs(4143));
    layer1_outputs(2423) <= (layer0_outputs(2488)) and not (layer0_outputs(107));
    layer1_outputs(2424) <= not((layer0_outputs(2089)) xor (layer0_outputs(3900)));
    layer1_outputs(2425) <= not(layer0_outputs(4870)) or (layer0_outputs(4716));
    layer1_outputs(2426) <= not(layer0_outputs(817));
    layer1_outputs(2427) <= (layer0_outputs(4674)) and not (layer0_outputs(2044));
    layer1_outputs(2428) <= (layer0_outputs(3372)) and not (layer0_outputs(2326));
    layer1_outputs(2429) <= layer0_outputs(4425);
    layer1_outputs(2430) <= (layer0_outputs(410)) or (layer0_outputs(3972));
    layer1_outputs(2431) <= not(layer0_outputs(2161));
    layer1_outputs(2432) <= not(layer0_outputs(884)) or (layer0_outputs(3162));
    layer1_outputs(2433) <= not((layer0_outputs(587)) or (layer0_outputs(2843)));
    layer1_outputs(2434) <= layer0_outputs(2323);
    layer1_outputs(2435) <= not(layer0_outputs(2923));
    layer1_outputs(2436) <= not(layer0_outputs(4416));
    layer1_outputs(2437) <= '0';
    layer1_outputs(2438) <= not(layer0_outputs(2519)) or (layer0_outputs(1822));
    layer1_outputs(2439) <= not((layer0_outputs(3972)) or (layer0_outputs(3134)));
    layer1_outputs(2440) <= (layer0_outputs(4742)) and not (layer0_outputs(701));
    layer1_outputs(2441) <= (layer0_outputs(995)) or (layer0_outputs(381));
    layer1_outputs(2442) <= layer0_outputs(4310);
    layer1_outputs(2443) <= (layer0_outputs(3071)) and not (layer0_outputs(1789));
    layer1_outputs(2444) <= layer0_outputs(327);
    layer1_outputs(2445) <= not((layer0_outputs(4193)) or (layer0_outputs(524)));
    layer1_outputs(2446) <= not((layer0_outputs(3064)) and (layer0_outputs(3137)));
    layer1_outputs(2447) <= not(layer0_outputs(1910));
    layer1_outputs(2448) <= not(layer0_outputs(150));
    layer1_outputs(2449) <= (layer0_outputs(3356)) and not (layer0_outputs(1395));
    layer1_outputs(2450) <= layer0_outputs(2991);
    layer1_outputs(2451) <= not(layer0_outputs(413)) or (layer0_outputs(1309));
    layer1_outputs(2452) <= not(layer0_outputs(3274));
    layer1_outputs(2453) <= not(layer0_outputs(1872)) or (layer0_outputs(3564));
    layer1_outputs(2454) <= not(layer0_outputs(441));
    layer1_outputs(2455) <= (layer0_outputs(3936)) and (layer0_outputs(3603));
    layer1_outputs(2456) <= '0';
    layer1_outputs(2457) <= not((layer0_outputs(4445)) xor (layer0_outputs(2666)));
    layer1_outputs(2458) <= not((layer0_outputs(1619)) or (layer0_outputs(3236)));
    layer1_outputs(2459) <= not((layer0_outputs(1314)) or (layer0_outputs(2240)));
    layer1_outputs(2460) <= layer0_outputs(1739);
    layer1_outputs(2461) <= (layer0_outputs(2197)) and not (layer0_outputs(2117));
    layer1_outputs(2462) <= (layer0_outputs(871)) and not (layer0_outputs(3701));
    layer1_outputs(2463) <= layer0_outputs(1660);
    layer1_outputs(2464) <= (layer0_outputs(5008)) or (layer0_outputs(1025));
    layer1_outputs(2465) <= '0';
    layer1_outputs(2466) <= (layer0_outputs(1978)) and not (layer0_outputs(1177));
    layer1_outputs(2467) <= layer0_outputs(1744);
    layer1_outputs(2468) <= (layer0_outputs(3473)) and not (layer0_outputs(137));
    layer1_outputs(2469) <= not(layer0_outputs(1887)) or (layer0_outputs(1101));
    layer1_outputs(2470) <= '1';
    layer1_outputs(2471) <= not(layer0_outputs(1012)) or (layer0_outputs(2356));
    layer1_outputs(2472) <= (layer0_outputs(4268)) or (layer0_outputs(3855));
    layer1_outputs(2473) <= (layer0_outputs(3409)) xor (layer0_outputs(235));
    layer1_outputs(2474) <= (layer0_outputs(3851)) and (layer0_outputs(4855));
    layer1_outputs(2475) <= layer0_outputs(1205);
    layer1_outputs(2476) <= not(layer0_outputs(1620));
    layer1_outputs(2477) <= not(layer0_outputs(3197));
    layer1_outputs(2478) <= (layer0_outputs(3012)) xor (layer0_outputs(1043));
    layer1_outputs(2479) <= '1';
    layer1_outputs(2480) <= not(layer0_outputs(2655)) or (layer0_outputs(2361));
    layer1_outputs(2481) <= not(layer0_outputs(396));
    layer1_outputs(2482) <= (layer0_outputs(2979)) and not (layer0_outputs(2151));
    layer1_outputs(2483) <= (layer0_outputs(3618)) xor (layer0_outputs(874));
    layer1_outputs(2484) <= not(layer0_outputs(4842)) or (layer0_outputs(3179));
    layer1_outputs(2485) <= not((layer0_outputs(1751)) or (layer0_outputs(5094)));
    layer1_outputs(2486) <= not((layer0_outputs(2912)) and (layer0_outputs(3634)));
    layer1_outputs(2487) <= (layer0_outputs(3503)) or (layer0_outputs(3667));
    layer1_outputs(2488) <= not((layer0_outputs(2754)) xor (layer0_outputs(3799)));
    layer1_outputs(2489) <= not(layer0_outputs(3831)) or (layer0_outputs(1670));
    layer1_outputs(2490) <= (layer0_outputs(2098)) or (layer0_outputs(4158));
    layer1_outputs(2491) <= (layer0_outputs(4692)) xor (layer0_outputs(1456));
    layer1_outputs(2492) <= not((layer0_outputs(1343)) xor (layer0_outputs(2157)));
    layer1_outputs(2493) <= (layer0_outputs(1410)) and not (layer0_outputs(3839));
    layer1_outputs(2494) <= not((layer0_outputs(3103)) or (layer0_outputs(793)));
    layer1_outputs(2495) <= not(layer0_outputs(4688));
    layer1_outputs(2496) <= not(layer0_outputs(649));
    layer1_outputs(2497) <= (layer0_outputs(3512)) and (layer0_outputs(1480));
    layer1_outputs(2498) <= not((layer0_outputs(219)) or (layer0_outputs(951)));
    layer1_outputs(2499) <= (layer0_outputs(2827)) and not (layer0_outputs(1475));
    layer1_outputs(2500) <= '1';
    layer1_outputs(2501) <= not((layer0_outputs(4697)) and (layer0_outputs(1799)));
    layer1_outputs(2502) <= layer0_outputs(4334);
    layer1_outputs(2503) <= layer0_outputs(4724);
    layer1_outputs(2504) <= not(layer0_outputs(3211)) or (layer0_outputs(2213));
    layer1_outputs(2505) <= (layer0_outputs(778)) and not (layer0_outputs(2833));
    layer1_outputs(2506) <= not(layer0_outputs(1987)) or (layer0_outputs(1348));
    layer1_outputs(2507) <= not(layer0_outputs(681));
    layer1_outputs(2508) <= (layer0_outputs(2336)) or (layer0_outputs(419));
    layer1_outputs(2509) <= not((layer0_outputs(1145)) xor (layer0_outputs(628)));
    layer1_outputs(2510) <= not((layer0_outputs(4943)) and (layer0_outputs(3690)));
    layer1_outputs(2511) <= layer0_outputs(3541);
    layer1_outputs(2512) <= (layer0_outputs(3336)) or (layer0_outputs(4282));
    layer1_outputs(2513) <= not(layer0_outputs(3060));
    layer1_outputs(2514) <= '0';
    layer1_outputs(2515) <= layer0_outputs(3872);
    layer1_outputs(2516) <= not((layer0_outputs(759)) xor (layer0_outputs(2744)));
    layer1_outputs(2517) <= layer0_outputs(1305);
    layer1_outputs(2518) <= layer0_outputs(1137);
    layer1_outputs(2519) <= '0';
    layer1_outputs(2520) <= not(layer0_outputs(3821));
    layer1_outputs(2521) <= not((layer0_outputs(3490)) and (layer0_outputs(4384)));
    layer1_outputs(2522) <= (layer0_outputs(3860)) and (layer0_outputs(2315));
    layer1_outputs(2523) <= (layer0_outputs(4583)) xor (layer0_outputs(1876));
    layer1_outputs(2524) <= (layer0_outputs(4602)) and not (layer0_outputs(835));
    layer1_outputs(2525) <= (layer0_outputs(212)) and not (layer0_outputs(2401));
    layer1_outputs(2526) <= (layer0_outputs(4676)) xor (layer0_outputs(3817));
    layer1_outputs(2527) <= not((layer0_outputs(2263)) or (layer0_outputs(2451)));
    layer1_outputs(2528) <= not(layer0_outputs(850));
    layer1_outputs(2529) <= layer0_outputs(1341);
    layer1_outputs(2530) <= (layer0_outputs(3982)) and not (layer0_outputs(1164));
    layer1_outputs(2531) <= not(layer0_outputs(692));
    layer1_outputs(2532) <= (layer0_outputs(2580)) and (layer0_outputs(2614));
    layer1_outputs(2533) <= (layer0_outputs(3369)) or (layer0_outputs(1906));
    layer1_outputs(2534) <= layer0_outputs(1429);
    layer1_outputs(2535) <= not(layer0_outputs(4288));
    layer1_outputs(2536) <= (layer0_outputs(4860)) or (layer0_outputs(1087));
    layer1_outputs(2537) <= not(layer0_outputs(3281));
    layer1_outputs(2538) <= (layer0_outputs(1840)) and not (layer0_outputs(1543));
    layer1_outputs(2539) <= not(layer0_outputs(1169));
    layer1_outputs(2540) <= not((layer0_outputs(826)) and (layer0_outputs(383)));
    layer1_outputs(2541) <= not((layer0_outputs(2085)) or (layer0_outputs(1901)));
    layer1_outputs(2542) <= not(layer0_outputs(3513));
    layer1_outputs(2543) <= not(layer0_outputs(3297)) or (layer0_outputs(203));
    layer1_outputs(2544) <= not((layer0_outputs(3066)) xor (layer0_outputs(3389)));
    layer1_outputs(2545) <= layer0_outputs(4539);
    layer1_outputs(2546) <= not((layer0_outputs(4749)) and (layer0_outputs(3386)));
    layer1_outputs(2547) <= layer0_outputs(4136);
    layer1_outputs(2548) <= not(layer0_outputs(1989)) or (layer0_outputs(5022));
    layer1_outputs(2549) <= not(layer0_outputs(1118));
    layer1_outputs(2550) <= (layer0_outputs(4570)) or (layer0_outputs(2218));
    layer1_outputs(2551) <= not((layer0_outputs(230)) or (layer0_outputs(891)));
    layer1_outputs(2552) <= '1';
    layer1_outputs(2553) <= (layer0_outputs(753)) or (layer0_outputs(5117));
    layer1_outputs(2554) <= not(layer0_outputs(175)) or (layer0_outputs(1955));
    layer1_outputs(2555) <= not(layer0_outputs(910));
    layer1_outputs(2556) <= not(layer0_outputs(4922));
    layer1_outputs(2557) <= not(layer0_outputs(1778)) or (layer0_outputs(4874));
    layer1_outputs(2558) <= not(layer0_outputs(2606)) or (layer0_outputs(1870));
    layer1_outputs(2559) <= '1';
    layer1_outputs(2560) <= not((layer0_outputs(554)) or (layer0_outputs(1056)));
    layer1_outputs(2561) <= not(layer0_outputs(3691)) or (layer0_outputs(3785));
    layer1_outputs(2562) <= layer0_outputs(4524);
    layer1_outputs(2563) <= (layer0_outputs(4608)) and (layer0_outputs(1914));
    layer1_outputs(2564) <= not(layer0_outputs(907));
    layer1_outputs(2565) <= (layer0_outputs(279)) and not (layer0_outputs(1761));
    layer1_outputs(2566) <= '0';
    layer1_outputs(2567) <= (layer0_outputs(4658)) or (layer0_outputs(4756));
    layer1_outputs(2568) <= not((layer0_outputs(952)) xor (layer0_outputs(1537)));
    layer1_outputs(2569) <= not(layer0_outputs(1035));
    layer1_outputs(2570) <= not((layer0_outputs(4799)) xor (layer0_outputs(2405)));
    layer1_outputs(2571) <= not(layer0_outputs(264));
    layer1_outputs(2572) <= not((layer0_outputs(3812)) xor (layer0_outputs(886)));
    layer1_outputs(2573) <= not(layer0_outputs(2969)) or (layer0_outputs(1956));
    layer1_outputs(2574) <= layer0_outputs(3726);
    layer1_outputs(2575) <= not((layer0_outputs(387)) xor (layer0_outputs(3895)));
    layer1_outputs(2576) <= layer0_outputs(4851);
    layer1_outputs(2577) <= (layer0_outputs(1196)) xor (layer0_outputs(1677));
    layer1_outputs(2578) <= not((layer0_outputs(1415)) and (layer0_outputs(2801)));
    layer1_outputs(2579) <= layer0_outputs(1710);
    layer1_outputs(2580) <= not(layer0_outputs(4098));
    layer1_outputs(2581) <= (layer0_outputs(3024)) xor (layer0_outputs(1183));
    layer1_outputs(2582) <= layer0_outputs(2843);
    layer1_outputs(2583) <= layer0_outputs(1008);
    layer1_outputs(2584) <= (layer0_outputs(2688)) or (layer0_outputs(273));
    layer1_outputs(2585) <= layer0_outputs(2137);
    layer1_outputs(2586) <= (layer0_outputs(3643)) and not (layer0_outputs(5052));
    layer1_outputs(2587) <= (layer0_outputs(4698)) or (layer0_outputs(206));
    layer1_outputs(2588) <= (layer0_outputs(4806)) and not (layer0_outputs(1600));
    layer1_outputs(2589) <= layer0_outputs(4395);
    layer1_outputs(2590) <= (layer0_outputs(336)) and not (layer0_outputs(818));
    layer1_outputs(2591) <= (layer0_outputs(967)) and not (layer0_outputs(4626));
    layer1_outputs(2592) <= not(layer0_outputs(117)) or (layer0_outputs(2225));
    layer1_outputs(2593) <= (layer0_outputs(4141)) and not (layer0_outputs(2212));
    layer1_outputs(2594) <= (layer0_outputs(2355)) and not (layer0_outputs(3107));
    layer1_outputs(2595) <= (layer0_outputs(3558)) and (layer0_outputs(755));
    layer1_outputs(2596) <= not(layer0_outputs(1022));
    layer1_outputs(2597) <= not((layer0_outputs(1211)) or (layer0_outputs(220)));
    layer1_outputs(2598) <= '1';
    layer1_outputs(2599) <= not((layer0_outputs(2105)) and (layer0_outputs(4785)));
    layer1_outputs(2600) <= not(layer0_outputs(1555));
    layer1_outputs(2601) <= (layer0_outputs(2562)) and (layer0_outputs(1720));
    layer1_outputs(2602) <= not(layer0_outputs(43));
    layer1_outputs(2603) <= layer0_outputs(3224);
    layer1_outputs(2604) <= layer0_outputs(2672);
    layer1_outputs(2605) <= not(layer0_outputs(2670));
    layer1_outputs(2606) <= layer0_outputs(4925);
    layer1_outputs(2607) <= not((layer0_outputs(1967)) xor (layer0_outputs(2698)));
    layer1_outputs(2608) <= not(layer0_outputs(579)) or (layer0_outputs(4151));
    layer1_outputs(2609) <= (layer0_outputs(1200)) or (layer0_outputs(1306));
    layer1_outputs(2610) <= (layer0_outputs(3823)) and not (layer0_outputs(3249));
    layer1_outputs(2611) <= (layer0_outputs(3626)) and (layer0_outputs(171));
    layer1_outputs(2612) <= not(layer0_outputs(3819));
    layer1_outputs(2613) <= '0';
    layer1_outputs(2614) <= not(layer0_outputs(4826));
    layer1_outputs(2615) <= layer0_outputs(1095);
    layer1_outputs(2616) <= (layer0_outputs(1223)) and not (layer0_outputs(2555));
    layer1_outputs(2617) <= (layer0_outputs(4911)) or (layer0_outputs(1109));
    layer1_outputs(2618) <= not(layer0_outputs(2270));
    layer1_outputs(2619) <= layer0_outputs(2638);
    layer1_outputs(2620) <= layer0_outputs(2701);
    layer1_outputs(2621) <= not((layer0_outputs(4520)) and (layer0_outputs(3430)));
    layer1_outputs(2622) <= (layer0_outputs(1747)) and not (layer0_outputs(2109));
    layer1_outputs(2623) <= (layer0_outputs(4429)) and (layer0_outputs(2815));
    layer1_outputs(2624) <= not(layer0_outputs(4417));
    layer1_outputs(2625) <= layer0_outputs(768);
    layer1_outputs(2626) <= (layer0_outputs(1013)) and not (layer0_outputs(681));
    layer1_outputs(2627) <= not((layer0_outputs(1014)) or (layer0_outputs(3306)));
    layer1_outputs(2628) <= (layer0_outputs(2959)) and not (layer0_outputs(4843));
    layer1_outputs(2629) <= (layer0_outputs(4802)) xor (layer0_outputs(2642));
    layer1_outputs(2630) <= not(layer0_outputs(4413)) or (layer0_outputs(2576));
    layer1_outputs(2631) <= not(layer0_outputs(2350)) or (layer0_outputs(675));
    layer1_outputs(2632) <= (layer0_outputs(4635)) xor (layer0_outputs(477));
    layer1_outputs(2633) <= not(layer0_outputs(1646));
    layer1_outputs(2634) <= not(layer0_outputs(1401));
    layer1_outputs(2635) <= not(layer0_outputs(1297)) or (layer0_outputs(134));
    layer1_outputs(2636) <= not((layer0_outputs(3934)) and (layer0_outputs(4107)));
    layer1_outputs(2637) <= '1';
    layer1_outputs(2638) <= not(layer0_outputs(477));
    layer1_outputs(2639) <= (layer0_outputs(1263)) and (layer0_outputs(3897));
    layer1_outputs(2640) <= not(layer0_outputs(4167));
    layer1_outputs(2641) <= not(layer0_outputs(1526)) or (layer0_outputs(4820));
    layer1_outputs(2642) <= layer0_outputs(1174);
    layer1_outputs(2643) <= not(layer0_outputs(4619));
    layer1_outputs(2644) <= layer0_outputs(3743);
    layer1_outputs(2645) <= not(layer0_outputs(257));
    layer1_outputs(2646) <= (layer0_outputs(4878)) and (layer0_outputs(1889));
    layer1_outputs(2647) <= '1';
    layer1_outputs(2648) <= layer0_outputs(777);
    layer1_outputs(2649) <= (layer0_outputs(714)) and (layer0_outputs(1690));
    layer1_outputs(2650) <= (layer0_outputs(306)) or (layer0_outputs(4333));
    layer1_outputs(2651) <= (layer0_outputs(327)) and not (layer0_outputs(4927));
    layer1_outputs(2652) <= not(layer0_outputs(483)) or (layer0_outputs(580));
    layer1_outputs(2653) <= not((layer0_outputs(936)) or (layer0_outputs(1399)));
    layer1_outputs(2654) <= (layer0_outputs(4841)) and (layer0_outputs(128));
    layer1_outputs(2655) <= (layer0_outputs(3844)) and not (layer0_outputs(5026));
    layer1_outputs(2656) <= not(layer0_outputs(1570));
    layer1_outputs(2657) <= not(layer0_outputs(151));
    layer1_outputs(2658) <= not(layer0_outputs(726));
    layer1_outputs(2659) <= (layer0_outputs(4188)) and (layer0_outputs(4944));
    layer1_outputs(2660) <= not(layer0_outputs(3554));
    layer1_outputs(2661) <= (layer0_outputs(1728)) and not (layer0_outputs(3289));
    layer1_outputs(2662) <= (layer0_outputs(4031)) or (layer0_outputs(2242));
    layer1_outputs(2663) <= layer0_outputs(2978);
    layer1_outputs(2664) <= not((layer0_outputs(1344)) or (layer0_outputs(3077)));
    layer1_outputs(2665) <= layer0_outputs(1142);
    layer1_outputs(2666) <= layer0_outputs(28);
    layer1_outputs(2667) <= not(layer0_outputs(2752));
    layer1_outputs(2668) <= (layer0_outputs(3083)) and not (layer0_outputs(1681));
    layer1_outputs(2669) <= (layer0_outputs(2160)) and not (layer0_outputs(3969));
    layer1_outputs(2670) <= not(layer0_outputs(2472));
    layer1_outputs(2671) <= not((layer0_outputs(4820)) xor (layer0_outputs(378)));
    layer1_outputs(2672) <= not((layer0_outputs(3723)) and (layer0_outputs(1972)));
    layer1_outputs(2673) <= not((layer0_outputs(3655)) and (layer0_outputs(3814)));
    layer1_outputs(2674) <= '0';
    layer1_outputs(2675) <= not((layer0_outputs(4736)) xor (layer0_outputs(1490)));
    layer1_outputs(2676) <= not(layer0_outputs(2682)) or (layer0_outputs(2504));
    layer1_outputs(2677) <= (layer0_outputs(815)) and not (layer0_outputs(1215));
    layer1_outputs(2678) <= (layer0_outputs(3830)) or (layer0_outputs(85));
    layer1_outputs(2679) <= (layer0_outputs(2305)) and not (layer0_outputs(4410));
    layer1_outputs(2680) <= '1';
    layer1_outputs(2681) <= not(layer0_outputs(4119)) or (layer0_outputs(91));
    layer1_outputs(2682) <= not(layer0_outputs(3428)) or (layer0_outputs(3923));
    layer1_outputs(2683) <= not(layer0_outputs(4130));
    layer1_outputs(2684) <= not((layer0_outputs(3508)) or (layer0_outputs(1520)));
    layer1_outputs(2685) <= layer0_outputs(3063);
    layer1_outputs(2686) <= not((layer0_outputs(438)) xor (layer0_outputs(2905)));
    layer1_outputs(2687) <= not(layer0_outputs(4904)) or (layer0_outputs(3707));
    layer1_outputs(2688) <= not(layer0_outputs(4921)) or (layer0_outputs(1513));
    layer1_outputs(2689) <= (layer0_outputs(3638)) xor (layer0_outputs(4122));
    layer1_outputs(2690) <= not(layer0_outputs(2576)) or (layer0_outputs(1531));
    layer1_outputs(2691) <= not((layer0_outputs(1777)) and (layer0_outputs(4367)));
    layer1_outputs(2692) <= (layer0_outputs(4299)) and not (layer0_outputs(3102));
    layer1_outputs(2693) <= not((layer0_outputs(3596)) and (layer0_outputs(2023)));
    layer1_outputs(2694) <= layer0_outputs(4999);
    layer1_outputs(2695) <= (layer0_outputs(637)) and (layer0_outputs(413));
    layer1_outputs(2696) <= layer0_outputs(966);
    layer1_outputs(2697) <= layer0_outputs(3744);
    layer1_outputs(2698) <= not(layer0_outputs(2383)) or (layer0_outputs(2740));
    layer1_outputs(2699) <= (layer0_outputs(2145)) and not (layer0_outputs(1695));
    layer1_outputs(2700) <= layer0_outputs(2791);
    layer1_outputs(2701) <= not(layer0_outputs(4349)) or (layer0_outputs(4192));
    layer1_outputs(2702) <= not(layer0_outputs(1999));
    layer1_outputs(2703) <= not(layer0_outputs(3340));
    layer1_outputs(2704) <= (layer0_outputs(2430)) and (layer0_outputs(1148));
    layer1_outputs(2705) <= (layer0_outputs(3978)) and (layer0_outputs(2159));
    layer1_outputs(2706) <= not(layer0_outputs(2924));
    layer1_outputs(2707) <= not(layer0_outputs(3717)) or (layer0_outputs(4244));
    layer1_outputs(2708) <= not(layer0_outputs(3753));
    layer1_outputs(2709) <= layer0_outputs(4247);
    layer1_outputs(2710) <= not(layer0_outputs(4152));
    layer1_outputs(2711) <= layer0_outputs(4128);
    layer1_outputs(2712) <= layer0_outputs(2056);
    layer1_outputs(2713) <= not(layer0_outputs(128));
    layer1_outputs(2714) <= not((layer0_outputs(749)) xor (layer0_outputs(2784)));
    layer1_outputs(2715) <= '0';
    layer1_outputs(2716) <= not(layer0_outputs(4614));
    layer1_outputs(2717) <= not((layer0_outputs(372)) xor (layer0_outputs(3597)));
    layer1_outputs(2718) <= not(layer0_outputs(1591)) or (layer0_outputs(4717));
    layer1_outputs(2719) <= (layer0_outputs(2648)) and (layer0_outputs(3258));
    layer1_outputs(2720) <= not((layer0_outputs(1034)) and (layer0_outputs(3260)));
    layer1_outputs(2721) <= (layer0_outputs(3900)) xor (layer0_outputs(3323));
    layer1_outputs(2722) <= not(layer0_outputs(511));
    layer1_outputs(2723) <= not(layer0_outputs(596));
    layer1_outputs(2724) <= not(layer0_outputs(4144)) or (layer0_outputs(2606));
    layer1_outputs(2725) <= not((layer0_outputs(4173)) xor (layer0_outputs(2529)));
    layer1_outputs(2726) <= not(layer0_outputs(863)) or (layer0_outputs(2312));
    layer1_outputs(2727) <= not((layer0_outputs(4051)) xor (layer0_outputs(2759)));
    layer1_outputs(2728) <= layer0_outputs(942);
    layer1_outputs(2729) <= layer0_outputs(4598);
    layer1_outputs(2730) <= not(layer0_outputs(1917));
    layer1_outputs(2731) <= not(layer0_outputs(5029));
    layer1_outputs(2732) <= '0';
    layer1_outputs(2733) <= (layer0_outputs(4607)) and (layer0_outputs(3335));
    layer1_outputs(2734) <= not((layer0_outputs(4265)) xor (layer0_outputs(169)));
    layer1_outputs(2735) <= not((layer0_outputs(1883)) and (layer0_outputs(1601)));
    layer1_outputs(2736) <= (layer0_outputs(4278)) and not (layer0_outputs(2429));
    layer1_outputs(2737) <= not(layer0_outputs(2424)) or (layer0_outputs(321));
    layer1_outputs(2738) <= not(layer0_outputs(1109));
    layer1_outputs(2739) <= not(layer0_outputs(4292)) or (layer0_outputs(1810));
    layer1_outputs(2740) <= layer0_outputs(2130);
    layer1_outputs(2741) <= not((layer0_outputs(3403)) and (layer0_outputs(1663)));
    layer1_outputs(2742) <= not(layer0_outputs(1901));
    layer1_outputs(2743) <= not(layer0_outputs(1067)) or (layer0_outputs(2639));
    layer1_outputs(2744) <= not(layer0_outputs(4262)) or (layer0_outputs(2593));
    layer1_outputs(2745) <= not(layer0_outputs(176)) or (layer0_outputs(4777));
    layer1_outputs(2746) <= layer0_outputs(292);
    layer1_outputs(2747) <= not(layer0_outputs(4670)) or (layer0_outputs(582));
    layer1_outputs(2748) <= not(layer0_outputs(2415)) or (layer0_outputs(4408));
    layer1_outputs(2749) <= (layer0_outputs(1813)) and (layer0_outputs(2820));
    layer1_outputs(2750) <= not((layer0_outputs(3793)) xor (layer0_outputs(1913)));
    layer1_outputs(2751) <= (layer0_outputs(4091)) and not (layer0_outputs(999));
    layer1_outputs(2752) <= '0';
    layer1_outputs(2753) <= (layer0_outputs(2079)) and not (layer0_outputs(1944));
    layer1_outputs(2754) <= not(layer0_outputs(2362));
    layer1_outputs(2755) <= layer0_outputs(3934);
    layer1_outputs(2756) <= layer0_outputs(4432);
    layer1_outputs(2757) <= not(layer0_outputs(1832)) or (layer0_outputs(3133));
    layer1_outputs(2758) <= not(layer0_outputs(4438)) or (layer0_outputs(3534));
    layer1_outputs(2759) <= layer0_outputs(692);
    layer1_outputs(2760) <= not(layer0_outputs(3368));
    layer1_outputs(2761) <= (layer0_outputs(2793)) and (layer0_outputs(2239));
    layer1_outputs(2762) <= layer0_outputs(2759);
    layer1_outputs(2763) <= not(layer0_outputs(2729));
    layer1_outputs(2764) <= (layer0_outputs(2926)) and (layer0_outputs(386));
    layer1_outputs(2765) <= '1';
    layer1_outputs(2766) <= not(layer0_outputs(58)) or (layer0_outputs(3758));
    layer1_outputs(2767) <= not(layer0_outputs(3275));
    layer1_outputs(2768) <= '0';
    layer1_outputs(2769) <= layer0_outputs(2167);
    layer1_outputs(2770) <= (layer0_outputs(3053)) and (layer0_outputs(1939));
    layer1_outputs(2771) <= not((layer0_outputs(3578)) and (layer0_outputs(3098)));
    layer1_outputs(2772) <= not(layer0_outputs(3426));
    layer1_outputs(2773) <= (layer0_outputs(1955)) and not (layer0_outputs(3658));
    layer1_outputs(2774) <= not(layer0_outputs(285));
    layer1_outputs(2775) <= (layer0_outputs(798)) or (layer0_outputs(2954));
    layer1_outputs(2776) <= (layer0_outputs(1968)) and not (layer0_outputs(2775));
    layer1_outputs(2777) <= not(layer0_outputs(2345));
    layer1_outputs(2778) <= layer0_outputs(3914);
    layer1_outputs(2779) <= not(layer0_outputs(505));
    layer1_outputs(2780) <= '1';
    layer1_outputs(2781) <= not(layer0_outputs(4859));
    layer1_outputs(2782) <= layer0_outputs(2178);
    layer1_outputs(2783) <= (layer0_outputs(2771)) or (layer0_outputs(1239));
    layer1_outputs(2784) <= (layer0_outputs(2261)) and not (layer0_outputs(4638));
    layer1_outputs(2785) <= (layer0_outputs(653)) and not (layer0_outputs(1114));
    layer1_outputs(2786) <= (layer0_outputs(2932)) or (layer0_outputs(2746));
    layer1_outputs(2787) <= not(layer0_outputs(4003));
    layer1_outputs(2788) <= layer0_outputs(2935);
    layer1_outputs(2789) <= layer0_outputs(889);
    layer1_outputs(2790) <= not((layer0_outputs(3250)) or (layer0_outputs(2064)));
    layer1_outputs(2791) <= (layer0_outputs(425)) xor (layer0_outputs(290));
    layer1_outputs(2792) <= (layer0_outputs(23)) and not (layer0_outputs(722));
    layer1_outputs(2793) <= (layer0_outputs(1259)) or (layer0_outputs(1057));
    layer1_outputs(2794) <= not(layer0_outputs(2123));
    layer1_outputs(2795) <= not(layer0_outputs(4625));
    layer1_outputs(2796) <= not(layer0_outputs(3847));
    layer1_outputs(2797) <= (layer0_outputs(4092)) and not (layer0_outputs(971));
    layer1_outputs(2798) <= (layer0_outputs(854)) xor (layer0_outputs(2801));
    layer1_outputs(2799) <= not(layer0_outputs(4121)) or (layer0_outputs(4358));
    layer1_outputs(2800) <= layer0_outputs(3694);
    layer1_outputs(2801) <= (layer0_outputs(2569)) xor (layer0_outputs(4165));
    layer1_outputs(2802) <= layer0_outputs(3948);
    layer1_outputs(2803) <= not((layer0_outputs(182)) and (layer0_outputs(49)));
    layer1_outputs(2804) <= not(layer0_outputs(3363)) or (layer0_outputs(3428));
    layer1_outputs(2805) <= not(layer0_outputs(4473)) or (layer0_outputs(3192));
    layer1_outputs(2806) <= layer0_outputs(2644);
    layer1_outputs(2807) <= not(layer0_outputs(2951)) or (layer0_outputs(501));
    layer1_outputs(2808) <= layer0_outputs(5075);
    layer1_outputs(2809) <= (layer0_outputs(1523)) and not (layer0_outputs(1625));
    layer1_outputs(2810) <= not((layer0_outputs(40)) or (layer0_outputs(4365)));
    layer1_outputs(2811) <= not(layer0_outputs(380)) or (layer0_outputs(3054));
    layer1_outputs(2812) <= not(layer0_outputs(1983)) or (layer0_outputs(1784));
    layer1_outputs(2813) <= not(layer0_outputs(1582)) or (layer0_outputs(18));
    layer1_outputs(2814) <= (layer0_outputs(4185)) xor (layer0_outputs(1997));
    layer1_outputs(2815) <= not((layer0_outputs(4559)) xor (layer0_outputs(2836)));
    layer1_outputs(2816) <= not(layer0_outputs(1831));
    layer1_outputs(2817) <= not(layer0_outputs(3098));
    layer1_outputs(2818) <= (layer0_outputs(3420)) or (layer0_outputs(1836));
    layer1_outputs(2819) <= layer0_outputs(1378);
    layer1_outputs(2820) <= (layer0_outputs(2611)) xor (layer0_outputs(3318));
    layer1_outputs(2821) <= (layer0_outputs(2858)) xor (layer0_outputs(959));
    layer1_outputs(2822) <= layer0_outputs(3212);
    layer1_outputs(2823) <= not((layer0_outputs(4567)) or (layer0_outputs(657)));
    layer1_outputs(2824) <= layer0_outputs(2230);
    layer1_outputs(2825) <= not(layer0_outputs(1391));
    layer1_outputs(2826) <= not(layer0_outputs(3779));
    layer1_outputs(2827) <= (layer0_outputs(1180)) and (layer0_outputs(1634));
    layer1_outputs(2828) <= '1';
    layer1_outputs(2829) <= not(layer0_outputs(1104));
    layer1_outputs(2830) <= '1';
    layer1_outputs(2831) <= not((layer0_outputs(3173)) and (layer0_outputs(521)));
    layer1_outputs(2832) <= not((layer0_outputs(4395)) or (layer0_outputs(2719)));
    layer1_outputs(2833) <= (layer0_outputs(2288)) xor (layer0_outputs(4149));
    layer1_outputs(2834) <= not((layer0_outputs(2992)) xor (layer0_outputs(1067)));
    layer1_outputs(2835) <= layer0_outputs(4497);
    layer1_outputs(2836) <= (layer0_outputs(1184)) and not (layer0_outputs(2996));
    layer1_outputs(2837) <= (layer0_outputs(4110)) and not (layer0_outputs(3573));
    layer1_outputs(2838) <= (layer0_outputs(4382)) and not (layer0_outputs(3406));
    layer1_outputs(2839) <= not(layer0_outputs(3580));
    layer1_outputs(2840) <= not((layer0_outputs(195)) or (layer0_outputs(1346)));
    layer1_outputs(2841) <= not((layer0_outputs(3891)) or (layer0_outputs(1638)));
    layer1_outputs(2842) <= (layer0_outputs(2597)) xor (layer0_outputs(4350));
    layer1_outputs(2843) <= layer0_outputs(3466);
    layer1_outputs(2844) <= (layer0_outputs(4561)) or (layer0_outputs(3174));
    layer1_outputs(2845) <= not(layer0_outputs(4071)) or (layer0_outputs(728));
    layer1_outputs(2846) <= (layer0_outputs(265)) and not (layer0_outputs(401));
    layer1_outputs(2847) <= layer0_outputs(1778);
    layer1_outputs(2848) <= layer0_outputs(1626);
    layer1_outputs(2849) <= layer0_outputs(935);
    layer1_outputs(2850) <= not(layer0_outputs(3699)) or (layer0_outputs(734));
    layer1_outputs(2851) <= (layer0_outputs(4919)) and (layer0_outputs(3502));
    layer1_outputs(2852) <= not(layer0_outputs(3219));
    layer1_outputs(2853) <= not((layer0_outputs(239)) and (layer0_outputs(4462)));
    layer1_outputs(2854) <= layer0_outputs(1734);
    layer1_outputs(2855) <= not(layer0_outputs(1586)) or (layer0_outputs(1449));
    layer1_outputs(2856) <= not((layer0_outputs(5021)) or (layer0_outputs(1880)));
    layer1_outputs(2857) <= '1';
    layer1_outputs(2858) <= not(layer0_outputs(4243));
    layer1_outputs(2859) <= '0';
    layer1_outputs(2860) <= not(layer0_outputs(1489)) or (layer0_outputs(1323));
    layer1_outputs(2861) <= not(layer0_outputs(4629));
    layer1_outputs(2862) <= '1';
    layer1_outputs(2863) <= layer0_outputs(4542);
    layer1_outputs(2864) <= (layer0_outputs(2204)) xor (layer0_outputs(4839));
    layer1_outputs(2865) <= (layer0_outputs(3387)) or (layer0_outputs(2492));
    layer1_outputs(2866) <= (layer0_outputs(1667)) and (layer0_outputs(4035));
    layer1_outputs(2867) <= layer0_outputs(190);
    layer1_outputs(2868) <= not(layer0_outputs(1099)) or (layer0_outputs(4032));
    layer1_outputs(2869) <= (layer0_outputs(4752)) and not (layer0_outputs(4338));
    layer1_outputs(2870) <= '0';
    layer1_outputs(2871) <= (layer0_outputs(499)) xor (layer0_outputs(301));
    layer1_outputs(2872) <= not(layer0_outputs(4033));
    layer1_outputs(2873) <= (layer0_outputs(3488)) and not (layer0_outputs(1373));
    layer1_outputs(2874) <= layer0_outputs(3319);
    layer1_outputs(2875) <= layer0_outputs(2378);
    layer1_outputs(2876) <= (layer0_outputs(4396)) and not (layer0_outputs(3324));
    layer1_outputs(2877) <= layer0_outputs(3234);
    layer1_outputs(2878) <= (layer0_outputs(3888)) and not (layer0_outputs(1696));
    layer1_outputs(2879) <= layer0_outputs(3873);
    layer1_outputs(2880) <= (layer0_outputs(838)) xor (layer0_outputs(4966));
    layer1_outputs(2881) <= not(layer0_outputs(1245));
    layer1_outputs(2882) <= not((layer0_outputs(2588)) xor (layer0_outputs(3482)));
    layer1_outputs(2883) <= not(layer0_outputs(955));
    layer1_outputs(2884) <= layer0_outputs(5056);
    layer1_outputs(2885) <= (layer0_outputs(1376)) xor (layer0_outputs(1014));
    layer1_outputs(2886) <= (layer0_outputs(482)) and not (layer0_outputs(1356));
    layer1_outputs(2887) <= '0';
    layer1_outputs(2888) <= not(layer0_outputs(639));
    layer1_outputs(2889) <= (layer0_outputs(1468)) and not (layer0_outputs(2435));
    layer1_outputs(2890) <= (layer0_outputs(4714)) xor (layer0_outputs(1610));
    layer1_outputs(2891) <= (layer0_outputs(3188)) and not (layer0_outputs(4276));
    layer1_outputs(2892) <= not((layer0_outputs(1759)) or (layer0_outputs(3523)));
    layer1_outputs(2893) <= not((layer0_outputs(5047)) or (layer0_outputs(4470)));
    layer1_outputs(2894) <= (layer0_outputs(1544)) and not (layer0_outputs(4979));
    layer1_outputs(2895) <= not(layer0_outputs(4166));
    layer1_outputs(2896) <= not(layer0_outputs(4273));
    layer1_outputs(2897) <= (layer0_outputs(3358)) or (layer0_outputs(1572));
    layer1_outputs(2898) <= not((layer0_outputs(3508)) and (layer0_outputs(2780)));
    layer1_outputs(2899) <= not((layer0_outputs(2341)) or (layer0_outputs(3250)));
    layer1_outputs(2900) <= '0';
    layer1_outputs(2901) <= not((layer0_outputs(3571)) or (layer0_outputs(494)));
    layer1_outputs(2902) <= not(layer0_outputs(3019));
    layer1_outputs(2903) <= '1';
    layer1_outputs(2904) <= not(layer0_outputs(1390)) or (layer0_outputs(3441));
    layer1_outputs(2905) <= (layer0_outputs(4843)) xor (layer0_outputs(1767));
    layer1_outputs(2906) <= not((layer0_outputs(383)) xor (layer0_outputs(4932)));
    layer1_outputs(2907) <= not((layer0_outputs(3272)) or (layer0_outputs(1946)));
    layer1_outputs(2908) <= not(layer0_outputs(999));
    layer1_outputs(2909) <= layer0_outputs(4318);
    layer1_outputs(2910) <= layer0_outputs(4322);
    layer1_outputs(2911) <= (layer0_outputs(5025)) and (layer0_outputs(1365));
    layer1_outputs(2912) <= (layer0_outputs(1621)) and (layer0_outputs(2919));
    layer1_outputs(2913) <= (layer0_outputs(972)) and not (layer0_outputs(3820));
    layer1_outputs(2914) <= not(layer0_outputs(961)) or (layer0_outputs(2051));
    layer1_outputs(2915) <= not(layer0_outputs(2574));
    layer1_outputs(2916) <= (layer0_outputs(1023)) and (layer0_outputs(4354));
    layer1_outputs(2917) <= (layer0_outputs(2486)) or (layer0_outputs(695));
    layer1_outputs(2918) <= (layer0_outputs(1293)) or (layer0_outputs(4467));
    layer1_outputs(2919) <= not(layer0_outputs(2711)) or (layer0_outputs(3131));
    layer1_outputs(2920) <= layer0_outputs(4459);
    layer1_outputs(2921) <= not(layer0_outputs(3848)) or (layer0_outputs(5108));
    layer1_outputs(2922) <= (layer0_outputs(3321)) and (layer0_outputs(2975));
    layer1_outputs(2923) <= not((layer0_outputs(2748)) and (layer0_outputs(2785)));
    layer1_outputs(2924) <= (layer0_outputs(1134)) xor (layer0_outputs(4660));
    layer1_outputs(2925) <= layer0_outputs(4126);
    layer1_outputs(2926) <= (layer0_outputs(3927)) or (layer0_outputs(5034));
    layer1_outputs(2927) <= layer0_outputs(3588);
    layer1_outputs(2928) <= not(layer0_outputs(2417)) or (layer0_outputs(1196));
    layer1_outputs(2929) <= not(layer0_outputs(2969));
    layer1_outputs(2930) <= '1';
    layer1_outputs(2931) <= not((layer0_outputs(2825)) or (layer0_outputs(903)));
    layer1_outputs(2932) <= (layer0_outputs(350)) or (layer0_outputs(1735));
    layer1_outputs(2933) <= (layer0_outputs(3399)) and (layer0_outputs(1201));
    layer1_outputs(2934) <= layer0_outputs(353);
    layer1_outputs(2935) <= layer0_outputs(1265);
    layer1_outputs(2936) <= not(layer0_outputs(444));
    layer1_outputs(2937) <= (layer0_outputs(4929)) and not (layer0_outputs(1849));
    layer1_outputs(2938) <= (layer0_outputs(2269)) and not (layer0_outputs(1350));
    layer1_outputs(2939) <= not(layer0_outputs(3856));
    layer1_outputs(2940) <= not(layer0_outputs(4513));
    layer1_outputs(2941) <= '1';
    layer1_outputs(2942) <= (layer0_outputs(1648)) and not (layer0_outputs(4012));
    layer1_outputs(2943) <= (layer0_outputs(4808)) or (layer0_outputs(2165));
    layer1_outputs(2944) <= layer0_outputs(592);
    layer1_outputs(2945) <= not((layer0_outputs(4804)) xor (layer0_outputs(2442)));
    layer1_outputs(2946) <= (layer0_outputs(4661)) and (layer0_outputs(2185));
    layer1_outputs(2947) <= (layer0_outputs(1462)) and not (layer0_outputs(2427));
    layer1_outputs(2948) <= not((layer0_outputs(1567)) and (layer0_outputs(4087)));
    layer1_outputs(2949) <= not(layer0_outputs(3634));
    layer1_outputs(2950) <= not(layer0_outputs(4604)) or (layer0_outputs(3947));
    layer1_outputs(2951) <= layer0_outputs(2281);
    layer1_outputs(2952) <= (layer0_outputs(94)) xor (layer0_outputs(2748));
    layer1_outputs(2953) <= not((layer0_outputs(1562)) xor (layer0_outputs(2110)));
    layer1_outputs(2954) <= layer0_outputs(2063);
    layer1_outputs(2955) <= not((layer0_outputs(1152)) xor (layer0_outputs(4362)));
    layer1_outputs(2956) <= not(layer0_outputs(5042)) or (layer0_outputs(3766));
    layer1_outputs(2957) <= (layer0_outputs(1315)) and (layer0_outputs(1637));
    layer1_outputs(2958) <= not((layer0_outputs(2297)) xor (layer0_outputs(3942)));
    layer1_outputs(2959) <= not((layer0_outputs(1844)) xor (layer0_outputs(801)));
    layer1_outputs(2960) <= (layer0_outputs(3068)) and not (layer0_outputs(810));
    layer1_outputs(2961) <= (layer0_outputs(3762)) xor (layer0_outputs(4653));
    layer1_outputs(2962) <= not(layer0_outputs(2360));
    layer1_outputs(2963) <= not((layer0_outputs(2353)) or (layer0_outputs(3029)));
    layer1_outputs(2964) <= not(layer0_outputs(46));
    layer1_outputs(2965) <= not((layer0_outputs(366)) xor (layer0_outputs(625)));
    layer1_outputs(2966) <= '1';
    layer1_outputs(2967) <= not((layer0_outputs(4004)) xor (layer0_outputs(3352)));
    layer1_outputs(2968) <= layer0_outputs(3119);
    layer1_outputs(2969) <= not((layer0_outputs(2899)) and (layer0_outputs(3222)));
    layer1_outputs(2970) <= not(layer0_outputs(4463));
    layer1_outputs(2971) <= not((layer0_outputs(1141)) or (layer0_outputs(1667)));
    layer1_outputs(2972) <= not((layer0_outputs(4709)) and (layer0_outputs(642)));
    layer1_outputs(2973) <= (layer0_outputs(436)) and (layer0_outputs(1188));
    layer1_outputs(2974) <= not((layer0_outputs(2724)) and (layer0_outputs(3062)));
    layer1_outputs(2975) <= (layer0_outputs(594)) and (layer0_outputs(1163));
    layer1_outputs(2976) <= not((layer0_outputs(740)) xor (layer0_outputs(89)));
    layer1_outputs(2977) <= (layer0_outputs(4750)) and not (layer0_outputs(1205));
    layer1_outputs(2978) <= not(layer0_outputs(2102));
    layer1_outputs(2979) <= (layer0_outputs(49)) and not (layer0_outputs(257));
    layer1_outputs(2980) <= not(layer0_outputs(3243)) or (layer0_outputs(4486));
    layer1_outputs(2981) <= not(layer0_outputs(830));
    layer1_outputs(2982) <= not(layer0_outputs(4401));
    layer1_outputs(2983) <= (layer0_outputs(4594)) or (layer0_outputs(1614));
    layer1_outputs(2984) <= not(layer0_outputs(3874));
    layer1_outputs(2985) <= layer0_outputs(1342);
    layer1_outputs(2986) <= not(layer0_outputs(168)) or (layer0_outputs(2285));
    layer1_outputs(2987) <= not(layer0_outputs(3957)) or (layer0_outputs(3625));
    layer1_outputs(2988) <= not((layer0_outputs(5046)) and (layer0_outputs(815)));
    layer1_outputs(2989) <= not((layer0_outputs(3985)) xor (layer0_outputs(286)));
    layer1_outputs(2990) <= not((layer0_outputs(1966)) xor (layer0_outputs(2448)));
    layer1_outputs(2991) <= layer0_outputs(4954);
    layer1_outputs(2992) <= layer0_outputs(2331);
    layer1_outputs(2993) <= not(layer0_outputs(4941));
    layer1_outputs(2994) <= (layer0_outputs(3243)) or (layer0_outputs(3463));
    layer1_outputs(2995) <= (layer0_outputs(3046)) and not (layer0_outputs(2235));
    layer1_outputs(2996) <= not(layer0_outputs(2907)) or (layer0_outputs(2330));
    layer1_outputs(2997) <= (layer0_outputs(4259)) and (layer0_outputs(4314));
    layer1_outputs(2998) <= not((layer0_outputs(2605)) or (layer0_outputs(2678)));
    layer1_outputs(2999) <= not((layer0_outputs(3646)) or (layer0_outputs(2578)));
    layer1_outputs(3000) <= not(layer0_outputs(1074));
    layer1_outputs(3001) <= not(layer0_outputs(4340));
    layer1_outputs(3002) <= (layer0_outputs(624)) and not (layer0_outputs(1927));
    layer1_outputs(3003) <= '1';
    layer1_outputs(3004) <= (layer0_outputs(30)) and not (layer0_outputs(4848));
    layer1_outputs(3005) <= '1';
    layer1_outputs(3006) <= not(layer0_outputs(3484)) or (layer0_outputs(3233));
    layer1_outputs(3007) <= not(layer0_outputs(2078)) or (layer0_outputs(3205));
    layer1_outputs(3008) <= not((layer0_outputs(280)) xor (layer0_outputs(3104)));
    layer1_outputs(3009) <= not((layer0_outputs(3839)) or (layer0_outputs(1641)));
    layer1_outputs(3010) <= layer0_outputs(3741);
    layer1_outputs(3011) <= not(layer0_outputs(2756));
    layer1_outputs(3012) <= (layer0_outputs(3792)) and not (layer0_outputs(2530));
    layer1_outputs(3013) <= (layer0_outputs(2959)) and not (layer0_outputs(3805));
    layer1_outputs(3014) <= layer0_outputs(1274);
    layer1_outputs(3015) <= not((layer0_outputs(2103)) xor (layer0_outputs(601)));
    layer1_outputs(3016) <= layer0_outputs(2598);
    layer1_outputs(3017) <= not(layer0_outputs(85));
    layer1_outputs(3018) <= not((layer0_outputs(4185)) xor (layer0_outputs(3758)));
    layer1_outputs(3019) <= not(layer0_outputs(3810));
    layer1_outputs(3020) <= layer0_outputs(219);
    layer1_outputs(3021) <= (layer0_outputs(3776)) and not (layer0_outputs(4150));
    layer1_outputs(3022) <= not(layer0_outputs(4825));
    layer1_outputs(3023) <= '1';
    layer1_outputs(3024) <= (layer0_outputs(5015)) xor (layer0_outputs(539));
    layer1_outputs(3025) <= not(layer0_outputs(5066)) or (layer0_outputs(400));
    layer1_outputs(3026) <= not((layer0_outputs(480)) or (layer0_outputs(4579)));
    layer1_outputs(3027) <= not(layer0_outputs(4859));
    layer1_outputs(3028) <= (layer0_outputs(367)) and (layer0_outputs(4552));
    layer1_outputs(3029) <= not(layer0_outputs(1580));
    layer1_outputs(3030) <= not(layer0_outputs(1710));
    layer1_outputs(3031) <= (layer0_outputs(1133)) or (layer0_outputs(1770));
    layer1_outputs(3032) <= (layer0_outputs(782)) and not (layer0_outputs(2631));
    layer1_outputs(3033) <= '0';
    layer1_outputs(3034) <= (layer0_outputs(114)) and not (layer0_outputs(3720));
    layer1_outputs(3035) <= not(layer0_outputs(1443));
    layer1_outputs(3036) <= (layer0_outputs(4205)) xor (layer0_outputs(2605));
    layer1_outputs(3037) <= layer0_outputs(2572);
    layer1_outputs(3038) <= not((layer0_outputs(225)) and (layer0_outputs(3286)));
    layer1_outputs(3039) <= layer0_outputs(3341);
    layer1_outputs(3040) <= (layer0_outputs(59)) and not (layer0_outputs(3986));
    layer1_outputs(3041) <= not(layer0_outputs(554));
    layer1_outputs(3042) <= not((layer0_outputs(2573)) and (layer0_outputs(2092)));
    layer1_outputs(3043) <= not(layer0_outputs(1904));
    layer1_outputs(3044) <= not(layer0_outputs(611)) or (layer0_outputs(4739));
    layer1_outputs(3045) <= (layer0_outputs(1694)) or (layer0_outputs(3958));
    layer1_outputs(3046) <= not(layer0_outputs(3171)) or (layer0_outputs(1981));
    layer1_outputs(3047) <= not(layer0_outputs(1017)) or (layer0_outputs(4984));
    layer1_outputs(3048) <= (layer0_outputs(3047)) or (layer0_outputs(4780));
    layer1_outputs(3049) <= (layer0_outputs(3468)) and (layer0_outputs(2531));
    layer1_outputs(3050) <= not(layer0_outputs(1240));
    layer1_outputs(3051) <= not(layer0_outputs(2289));
    layer1_outputs(3052) <= layer0_outputs(3340);
    layer1_outputs(3053) <= not((layer0_outputs(1580)) xor (layer0_outputs(4897)));
    layer1_outputs(3054) <= (layer0_outputs(4235)) and not (layer0_outputs(2446));
    layer1_outputs(3055) <= layer0_outputs(2177);
    layer1_outputs(3056) <= not((layer0_outputs(537)) xor (layer0_outputs(4970)));
    layer1_outputs(3057) <= not(layer0_outputs(4336));
    layer1_outputs(3058) <= layer0_outputs(3436);
    layer1_outputs(3059) <= not(layer0_outputs(2030)) or (layer0_outputs(2222));
    layer1_outputs(3060) <= not(layer0_outputs(4816));
    layer1_outputs(3061) <= layer0_outputs(2357);
    layer1_outputs(3062) <= not(layer0_outputs(1236)) or (layer0_outputs(4574));
    layer1_outputs(3063) <= not((layer0_outputs(2949)) or (layer0_outputs(3877)));
    layer1_outputs(3064) <= not(layer0_outputs(2873));
    layer1_outputs(3065) <= not((layer0_outputs(2392)) or (layer0_outputs(940)));
    layer1_outputs(3066) <= not(layer0_outputs(4964)) or (layer0_outputs(988));
    layer1_outputs(3067) <= '1';
    layer1_outputs(3068) <= not(layer0_outputs(1358));
    layer1_outputs(3069) <= '1';
    layer1_outputs(3070) <= (layer0_outputs(3262)) and not (layer0_outputs(4993));
    layer1_outputs(3071) <= not((layer0_outputs(876)) xor (layer0_outputs(4436)));
    layer1_outputs(3072) <= layer0_outputs(3806);
    layer1_outputs(3073) <= not((layer0_outputs(3454)) and (layer0_outputs(3148)));
    layer1_outputs(3074) <= (layer0_outputs(5024)) or (layer0_outputs(1704));
    layer1_outputs(3075) <= '1';
    layer1_outputs(3076) <= not(layer0_outputs(67)) or (layer0_outputs(148));
    layer1_outputs(3077) <= not((layer0_outputs(3449)) or (layer0_outputs(2387)));
    layer1_outputs(3078) <= (layer0_outputs(4818)) xor (layer0_outputs(3619));
    layer1_outputs(3079) <= '1';
    layer1_outputs(3080) <= not(layer0_outputs(2488));
    layer1_outputs(3081) <= layer0_outputs(1202);
    layer1_outputs(3082) <= not(layer0_outputs(2402));
    layer1_outputs(3083) <= not((layer0_outputs(713)) or (layer0_outputs(4707)));
    layer1_outputs(3084) <= not(layer0_outputs(2224)) or (layer0_outputs(3947));
    layer1_outputs(3085) <= layer0_outputs(3444);
    layer1_outputs(3086) <= not(layer0_outputs(3220));
    layer1_outputs(3087) <= layer0_outputs(4497);
    layer1_outputs(3088) <= (layer0_outputs(3160)) or (layer0_outputs(1748));
    layer1_outputs(3089) <= not(layer0_outputs(1028));
    layer1_outputs(3090) <= layer0_outputs(2782);
    layer1_outputs(3091) <= '1';
    layer1_outputs(3092) <= layer0_outputs(2380);
    layer1_outputs(3093) <= layer0_outputs(3298);
    layer1_outputs(3094) <= (layer0_outputs(3288)) and not (layer0_outputs(2502));
    layer1_outputs(3095) <= (layer0_outputs(2857)) and not (layer0_outputs(1517));
    layer1_outputs(3096) <= not((layer0_outputs(210)) or (layer0_outputs(1784)));
    layer1_outputs(3097) <= not((layer0_outputs(3327)) xor (layer0_outputs(3527)));
    layer1_outputs(3098) <= not(layer0_outputs(3526));
    layer1_outputs(3099) <= (layer0_outputs(244)) and not (layer0_outputs(2819));
    layer1_outputs(3100) <= layer0_outputs(2150);
    layer1_outputs(3101) <= not(layer0_outputs(4097)) or (layer0_outputs(4195));
    layer1_outputs(3102) <= layer0_outputs(4132);
    layer1_outputs(3103) <= (layer0_outputs(4562)) xor (layer0_outputs(2525));
    layer1_outputs(3104) <= (layer0_outputs(2155)) and not (layer0_outputs(4918));
    layer1_outputs(3105) <= layer0_outputs(2188);
    layer1_outputs(3106) <= layer0_outputs(1098);
    layer1_outputs(3107) <= not(layer0_outputs(3631));
    layer1_outputs(3108) <= layer0_outputs(3271);
    layer1_outputs(3109) <= not(layer0_outputs(2194));
    layer1_outputs(3110) <= (layer0_outputs(4635)) or (layer0_outputs(664));
    layer1_outputs(3111) <= '0';
    layer1_outputs(3112) <= not((layer0_outputs(1772)) and (layer0_outputs(4409)));
    layer1_outputs(3113) <= (layer0_outputs(3376)) and (layer0_outputs(4384));
    layer1_outputs(3114) <= not((layer0_outputs(3644)) xor (layer0_outputs(2316)));
    layer1_outputs(3115) <= not(layer0_outputs(100));
    layer1_outputs(3116) <= not((layer0_outputs(1679)) and (layer0_outputs(3706)));
    layer1_outputs(3117) <= not((layer0_outputs(2633)) and (layer0_outputs(135)));
    layer1_outputs(3118) <= (layer0_outputs(4770)) and not (layer0_outputs(2493));
    layer1_outputs(3119) <= not((layer0_outputs(950)) and (layer0_outputs(1802)));
    layer1_outputs(3120) <= not(layer0_outputs(521));
    layer1_outputs(3121) <= not(layer0_outputs(3235));
    layer1_outputs(3122) <= layer0_outputs(3449);
    layer1_outputs(3123) <= not(layer0_outputs(4303)) or (layer0_outputs(4730));
    layer1_outputs(3124) <= not(layer0_outputs(4019));
    layer1_outputs(3125) <= not((layer0_outputs(2868)) or (layer0_outputs(934)));
    layer1_outputs(3126) <= (layer0_outputs(1007)) and not (layer0_outputs(4267));
    layer1_outputs(3127) <= not(layer0_outputs(5102));
    layer1_outputs(3128) <= not((layer0_outputs(2077)) and (layer0_outputs(4361)));
    layer1_outputs(3129) <= not(layer0_outputs(2557));
    layer1_outputs(3130) <= (layer0_outputs(797)) and not (layer0_outputs(1793));
    layer1_outputs(3131) <= not(layer0_outputs(2794));
    layer1_outputs(3132) <= (layer0_outputs(4782)) or (layer0_outputs(2218));
    layer1_outputs(3133) <= not((layer0_outputs(1051)) xor (layer0_outputs(2526)));
    layer1_outputs(3134) <= (layer0_outputs(5112)) or (layer0_outputs(772));
    layer1_outputs(3135) <= not(layer0_outputs(3929)) or (layer0_outputs(2713));
    layer1_outputs(3136) <= not((layer0_outputs(4677)) and (layer0_outputs(3537)));
    layer1_outputs(3137) <= not((layer0_outputs(4595)) or (layer0_outputs(3832)));
    layer1_outputs(3138) <= layer0_outputs(2095);
    layer1_outputs(3139) <= (layer0_outputs(4032)) xor (layer0_outputs(2376));
    layer1_outputs(3140) <= not((layer0_outputs(980)) and (layer0_outputs(513)));
    layer1_outputs(3141) <= not(layer0_outputs(4763)) or (layer0_outputs(1354));
    layer1_outputs(3142) <= (layer0_outputs(667)) and not (layer0_outputs(216));
    layer1_outputs(3143) <= not(layer0_outputs(1132));
    layer1_outputs(3144) <= not(layer0_outputs(3197)) or (layer0_outputs(1228));
    layer1_outputs(3145) <= not(layer0_outputs(1119));
    layer1_outputs(3146) <= not((layer0_outputs(2408)) or (layer0_outputs(2377)));
    layer1_outputs(3147) <= not(layer0_outputs(2390)) or (layer0_outputs(4848));
    layer1_outputs(3148) <= '1';
    layer1_outputs(3149) <= (layer0_outputs(395)) and not (layer0_outputs(2934));
    layer1_outputs(3150) <= not(layer0_outputs(1861));
    layer1_outputs(3151) <= (layer0_outputs(3521)) xor (layer0_outputs(3279));
    layer1_outputs(3152) <= layer0_outputs(5030);
    layer1_outputs(3153) <= (layer0_outputs(4589)) and not (layer0_outputs(1635));
    layer1_outputs(3154) <= not(layer0_outputs(3259));
    layer1_outputs(3155) <= not(layer0_outputs(2994)) or (layer0_outputs(4228));
    layer1_outputs(3156) <= (layer0_outputs(2498)) and (layer0_outputs(1156));
    layer1_outputs(3157) <= (layer0_outputs(5006)) and (layer0_outputs(5119));
    layer1_outputs(3158) <= layer0_outputs(5067);
    layer1_outputs(3159) <= not((layer0_outputs(3623)) and (layer0_outputs(3344)));
    layer1_outputs(3160) <= layer0_outputs(2778);
    layer1_outputs(3161) <= not(layer0_outputs(5061));
    layer1_outputs(3162) <= not(layer0_outputs(1225));
    layer1_outputs(3163) <= (layer0_outputs(2044)) and not (layer0_outputs(2849));
    layer1_outputs(3164) <= (layer0_outputs(962)) or (layer0_outputs(4427));
    layer1_outputs(3165) <= (layer0_outputs(3512)) xor (layer0_outputs(3472));
    layer1_outputs(3166) <= (layer0_outputs(3480)) xor (layer0_outputs(4376));
    layer1_outputs(3167) <= (layer0_outputs(737)) or (layer0_outputs(3153));
    layer1_outputs(3168) <= (layer0_outputs(4863)) and not (layer0_outputs(298));
    layer1_outputs(3169) <= not(layer0_outputs(3314));
    layer1_outputs(3170) <= layer0_outputs(1492);
    layer1_outputs(3171) <= not(layer0_outputs(3772));
    layer1_outputs(3172) <= not(layer0_outputs(3359));
    layer1_outputs(3173) <= layer0_outputs(218);
    layer1_outputs(3174) <= not((layer0_outputs(4541)) xor (layer0_outputs(4052)));
    layer1_outputs(3175) <= (layer0_outputs(2067)) and not (layer0_outputs(4639));
    layer1_outputs(3176) <= (layer0_outputs(1252)) and (layer0_outputs(4309));
    layer1_outputs(3177) <= (layer0_outputs(1873)) and (layer0_outputs(1669));
    layer1_outputs(3178) <= (layer0_outputs(595)) xor (layer0_outputs(774));
    layer1_outputs(3179) <= layer0_outputs(2547);
    layer1_outputs(3180) <= not(layer0_outputs(2807));
    layer1_outputs(3181) <= (layer0_outputs(4366)) and not (layer0_outputs(277));
    layer1_outputs(3182) <= not(layer0_outputs(3184));
    layer1_outputs(3183) <= not((layer0_outputs(1829)) and (layer0_outputs(1673)));
    layer1_outputs(3184) <= (layer0_outputs(4357)) or (layer0_outputs(3856));
    layer1_outputs(3185) <= not((layer0_outputs(630)) or (layer0_outputs(2431)));
    layer1_outputs(3186) <= not(layer0_outputs(961));
    layer1_outputs(3187) <= (layer0_outputs(2558)) and (layer0_outputs(4161));
    layer1_outputs(3188) <= (layer0_outputs(2195)) and not (layer0_outputs(4643));
    layer1_outputs(3189) <= not((layer0_outputs(570)) and (layer0_outputs(2394)));
    layer1_outputs(3190) <= not((layer0_outputs(4477)) xor (layer0_outputs(1172)));
    layer1_outputs(3191) <= (layer0_outputs(3493)) or (layer0_outputs(39));
    layer1_outputs(3192) <= not(layer0_outputs(1481)) or (layer0_outputs(2817));
    layer1_outputs(3193) <= not((layer0_outputs(4765)) or (layer0_outputs(258)));
    layer1_outputs(3194) <= not((layer0_outputs(3342)) and (layer0_outputs(928)));
    layer1_outputs(3195) <= not(layer0_outputs(3644)) or (layer0_outputs(2306));
    layer1_outputs(3196) <= (layer0_outputs(2662)) and (layer0_outputs(1301));
    layer1_outputs(3197) <= not(layer0_outputs(2700)) or (layer0_outputs(1065));
    layer1_outputs(3198) <= not(layer0_outputs(272));
    layer1_outputs(3199) <= layer0_outputs(978);
    layer1_outputs(3200) <= (layer0_outputs(4804)) xor (layer0_outputs(5084));
    layer1_outputs(3201) <= layer0_outputs(741);
    layer1_outputs(3202) <= not(layer0_outputs(1511));
    layer1_outputs(3203) <= not(layer0_outputs(2110)) or (layer0_outputs(4363));
    layer1_outputs(3204) <= (layer0_outputs(1234)) and not (layer0_outputs(3299));
    layer1_outputs(3205) <= not((layer0_outputs(1813)) or (layer0_outputs(2997)));
    layer1_outputs(3206) <= layer0_outputs(2299);
    layer1_outputs(3207) <= (layer0_outputs(1049)) and not (layer0_outputs(4885));
    layer1_outputs(3208) <= layer0_outputs(1891);
    layer1_outputs(3209) <= '1';
    layer1_outputs(3210) <= (layer0_outputs(217)) and (layer0_outputs(1634));
    layer1_outputs(3211) <= not(layer0_outputs(1134));
    layer1_outputs(3212) <= (layer0_outputs(5103)) and (layer0_outputs(3573));
    layer1_outputs(3213) <= not(layer0_outputs(4319));
    layer1_outputs(3214) <= (layer0_outputs(1471)) and not (layer0_outputs(3822));
    layer1_outputs(3215) <= not(layer0_outputs(2373)) or (layer0_outputs(789));
    layer1_outputs(3216) <= not(layer0_outputs(1698));
    layer1_outputs(3217) <= (layer0_outputs(2735)) and not (layer0_outputs(659));
    layer1_outputs(3218) <= not(layer0_outputs(2396)) or (layer0_outputs(2330));
    layer1_outputs(3219) <= (layer0_outputs(2668)) and not (layer0_outputs(119));
    layer1_outputs(3220) <= not((layer0_outputs(3060)) and (layer0_outputs(34)));
    layer1_outputs(3221) <= not(layer0_outputs(2828)) or (layer0_outputs(3507));
    layer1_outputs(3222) <= not(layer0_outputs(2331)) or (layer0_outputs(514));
    layer1_outputs(3223) <= not(layer0_outputs(2192));
    layer1_outputs(3224) <= not((layer0_outputs(2300)) or (layer0_outputs(4502)));
    layer1_outputs(3225) <= not(layer0_outputs(4277));
    layer1_outputs(3226) <= (layer0_outputs(3843)) xor (layer0_outputs(4137));
    layer1_outputs(3227) <= layer0_outputs(1865);
    layer1_outputs(3228) <= (layer0_outputs(2723)) and not (layer0_outputs(1581));
    layer1_outputs(3229) <= not((layer0_outputs(4821)) xor (layer0_outputs(3459)));
    layer1_outputs(3230) <= not(layer0_outputs(2080));
    layer1_outputs(3231) <= (layer0_outputs(1668)) and not (layer0_outputs(443));
    layer1_outputs(3232) <= not(layer0_outputs(395)) or (layer0_outputs(1423));
    layer1_outputs(3233) <= layer0_outputs(556);
    layer1_outputs(3234) <= layer0_outputs(3251);
    layer1_outputs(3235) <= not(layer0_outputs(4322)) or (layer0_outputs(92));
    layer1_outputs(3236) <= (layer0_outputs(4509)) and not (layer0_outputs(2522));
    layer1_outputs(3237) <= layer0_outputs(4368);
    layer1_outputs(3238) <= (layer0_outputs(4091)) and (layer0_outputs(2893));
    layer1_outputs(3239) <= not((layer0_outputs(1121)) or (layer0_outputs(927)));
    layer1_outputs(3240) <= (layer0_outputs(2548)) and (layer0_outputs(726));
    layer1_outputs(3241) <= (layer0_outputs(4597)) or (layer0_outputs(2565));
    layer1_outputs(3242) <= not((layer0_outputs(94)) and (layer0_outputs(218)));
    layer1_outputs(3243) <= (layer0_outputs(2766)) and (layer0_outputs(1382));
    layer1_outputs(3244) <= not((layer0_outputs(454)) and (layer0_outputs(2534)));
    layer1_outputs(3245) <= layer0_outputs(2186);
    layer1_outputs(3246) <= not(layer0_outputs(3009)) or (layer0_outputs(662));
    layer1_outputs(3247) <= not(layer0_outputs(1556));
    layer1_outputs(3248) <= not((layer0_outputs(1139)) xor (layer0_outputs(3199)));
    layer1_outputs(3249) <= (layer0_outputs(2357)) and not (layer0_outputs(754));
    layer1_outputs(3250) <= (layer0_outputs(3475)) and not (layer0_outputs(3742));
    layer1_outputs(3251) <= (layer0_outputs(3432)) and (layer0_outputs(5040));
    layer1_outputs(3252) <= (layer0_outputs(2133)) and not (layer0_outputs(4029));
    layer1_outputs(3253) <= (layer0_outputs(2008)) and not (layer0_outputs(2785));
    layer1_outputs(3254) <= not(layer0_outputs(3994));
    layer1_outputs(3255) <= not((layer0_outputs(2169)) or (layer0_outputs(3684)));
    layer1_outputs(3256) <= not((layer0_outputs(3497)) xor (layer0_outputs(3539)));
    layer1_outputs(3257) <= (layer0_outputs(3170)) xor (layer0_outputs(3140));
    layer1_outputs(3258) <= not((layer0_outputs(234)) or (layer0_outputs(4057)));
    layer1_outputs(3259) <= layer0_outputs(3723);
    layer1_outputs(3260) <= not(layer0_outputs(1024));
    layer1_outputs(3261) <= not(layer0_outputs(877));
    layer1_outputs(3262) <= (layer0_outputs(4713)) xor (layer0_outputs(2903));
    layer1_outputs(3263) <= (layer0_outputs(929)) or (layer0_outputs(3811));
    layer1_outputs(3264) <= layer0_outputs(2457);
    layer1_outputs(3265) <= not((layer0_outputs(4913)) or (layer0_outputs(4775)));
    layer1_outputs(3266) <= (layer0_outputs(3602)) and not (layer0_outputs(641));
    layer1_outputs(3267) <= not(layer0_outputs(1444));
    layer1_outputs(3268) <= not((layer0_outputs(1316)) xor (layer0_outputs(4387)));
    layer1_outputs(3269) <= (layer0_outputs(1202)) and not (layer0_outputs(2594));
    layer1_outputs(3270) <= not((layer0_outputs(2260)) and (layer0_outputs(3757)));
    layer1_outputs(3271) <= '1';
    layer1_outputs(3272) <= not(layer0_outputs(4702));
    layer1_outputs(3273) <= layer0_outputs(2777);
    layer1_outputs(3274) <= (layer0_outputs(3136)) xor (layer0_outputs(2503));
    layer1_outputs(3275) <= not((layer0_outputs(2108)) or (layer0_outputs(2037)));
    layer1_outputs(3276) <= not(layer0_outputs(3964));
    layer1_outputs(3277) <= not(layer0_outputs(2685));
    layer1_outputs(3278) <= not((layer0_outputs(3575)) or (layer0_outputs(2722)));
    layer1_outputs(3279) <= layer0_outputs(2050);
    layer1_outputs(3280) <= layer0_outputs(2475);
    layer1_outputs(3281) <= layer0_outputs(1991);
    layer1_outputs(3282) <= layer0_outputs(1544);
    layer1_outputs(3283) <= not(layer0_outputs(2889)) or (layer0_outputs(2732));
    layer1_outputs(3284) <= layer0_outputs(3298);
    layer1_outputs(3285) <= (layer0_outputs(3833)) and not (layer0_outputs(486));
    layer1_outputs(3286) <= not((layer0_outputs(308)) or (layer0_outputs(65)));
    layer1_outputs(3287) <= (layer0_outputs(1662)) and not (layer0_outputs(4633));
    layer1_outputs(3288) <= layer0_outputs(4969);
    layer1_outputs(3289) <= (layer0_outputs(4049)) or (layer0_outputs(1607));
    layer1_outputs(3290) <= (layer0_outputs(2261)) and (layer0_outputs(704));
    layer1_outputs(3291) <= not((layer0_outputs(847)) and (layer0_outputs(3784)));
    layer1_outputs(3292) <= not(layer0_outputs(1933));
    layer1_outputs(3293) <= (layer0_outputs(580)) and (layer0_outputs(4055));
    layer1_outputs(3294) <= not((layer0_outputs(689)) or (layer0_outputs(3560)));
    layer1_outputs(3295) <= layer0_outputs(2442);
    layer1_outputs(3296) <= not(layer0_outputs(5111));
    layer1_outputs(3297) <= not(layer0_outputs(920));
    layer1_outputs(3298) <= not(layer0_outputs(831)) or (layer0_outputs(2379));
    layer1_outputs(3299) <= layer0_outputs(517);
    layer1_outputs(3300) <= not(layer0_outputs(1814));
    layer1_outputs(3301) <= (layer0_outputs(1875)) and (layer0_outputs(1928));
    layer1_outputs(3302) <= not((layer0_outputs(1724)) or (layer0_outputs(3452)));
    layer1_outputs(3303) <= not((layer0_outputs(4306)) and (layer0_outputs(926)));
    layer1_outputs(3304) <= not((layer0_outputs(3565)) and (layer0_outputs(1661)));
    layer1_outputs(3305) <= not(layer0_outputs(4580)) or (layer0_outputs(670));
    layer1_outputs(3306) <= not(layer0_outputs(848)) or (layer0_outputs(3628));
    layer1_outputs(3307) <= (layer0_outputs(1149)) and not (layer0_outputs(1157));
    layer1_outputs(3308) <= not((layer0_outputs(2970)) or (layer0_outputs(65)));
    layer1_outputs(3309) <= not(layer0_outputs(75)) or (layer0_outputs(3069));
    layer1_outputs(3310) <= not((layer0_outputs(2236)) xor (layer0_outputs(736)));
    layer1_outputs(3311) <= (layer0_outputs(3632)) xor (layer0_outputs(1969));
    layer1_outputs(3312) <= not(layer0_outputs(1936));
    layer1_outputs(3313) <= (layer0_outputs(1791)) and not (layer0_outputs(2335));
    layer1_outputs(3314) <= (layer0_outputs(3496)) and (layer0_outputs(1538));
    layer1_outputs(3315) <= not((layer0_outputs(945)) and (layer0_outputs(1168)));
    layer1_outputs(3316) <= not((layer0_outputs(4420)) or (layer0_outputs(1982)));
    layer1_outputs(3317) <= not(layer0_outputs(2613)) or (layer0_outputs(1068));
    layer1_outputs(3318) <= (layer0_outputs(450)) and not (layer0_outputs(4890));
    layer1_outputs(3319) <= (layer0_outputs(4260)) and (layer0_outputs(488));
    layer1_outputs(3320) <= layer0_outputs(1246);
    layer1_outputs(3321) <= layer0_outputs(4636);
    layer1_outputs(3322) <= (layer0_outputs(270)) and not (layer0_outputs(4972));
    layer1_outputs(3323) <= not(layer0_outputs(1434));
    layer1_outputs(3324) <= not(layer0_outputs(2532));
    layer1_outputs(3325) <= not(layer0_outputs(1971)) or (layer0_outputs(1385));
    layer1_outputs(3326) <= not(layer0_outputs(4290)) or (layer0_outputs(1214));
    layer1_outputs(3327) <= not(layer0_outputs(1567));
    layer1_outputs(3328) <= (layer0_outputs(4082)) or (layer0_outputs(5087));
    layer1_outputs(3329) <= not(layer0_outputs(3470)) or (layer0_outputs(74));
    layer1_outputs(3330) <= not(layer0_outputs(2730)) or (layer0_outputs(1808));
    layer1_outputs(3331) <= (layer0_outputs(1915)) and (layer0_outputs(3305));
    layer1_outputs(3332) <= layer0_outputs(663);
    layer1_outputs(3333) <= (layer0_outputs(1564)) or (layer0_outputs(1614));
    layer1_outputs(3334) <= not((layer0_outputs(4673)) or (layer0_outputs(5012)));
    layer1_outputs(3335) <= (layer0_outputs(3993)) or (layer0_outputs(1952));
    layer1_outputs(3336) <= layer0_outputs(1603);
    layer1_outputs(3337) <= not((layer0_outputs(277)) or (layer0_outputs(5073)));
    layer1_outputs(3338) <= not(layer0_outputs(193)) or (layer0_outputs(4606));
    layer1_outputs(3339) <= layer0_outputs(2989);
    layer1_outputs(3340) <= (layer0_outputs(2026)) and not (layer0_outputs(2021));
    layer1_outputs(3341) <= (layer0_outputs(2504)) and not (layer0_outputs(4769));
    layer1_outputs(3342) <= (layer0_outputs(4229)) and not (layer0_outputs(1963));
    layer1_outputs(3343) <= not(layer0_outputs(2709));
    layer1_outputs(3344) <= not(layer0_outputs(132)) or (layer0_outputs(4459));
    layer1_outputs(3345) <= not((layer0_outputs(4022)) and (layer0_outputs(1493)));
    layer1_outputs(3346) <= not(layer0_outputs(356)) or (layer0_outputs(1675));
    layer1_outputs(3347) <= not(layer0_outputs(1898));
    layer1_outputs(3348) <= not(layer0_outputs(3000));
    layer1_outputs(3349) <= (layer0_outputs(3498)) and not (layer0_outputs(930));
    layer1_outputs(3350) <= '0';
    layer1_outputs(3351) <= (layer0_outputs(82)) and not (layer0_outputs(405));
    layer1_outputs(3352) <= not((layer0_outputs(866)) and (layer0_outputs(1757)));
    layer1_outputs(3353) <= not(layer0_outputs(1709));
    layer1_outputs(3354) <= '1';
    layer1_outputs(3355) <= layer0_outputs(4323);
    layer1_outputs(3356) <= not(layer0_outputs(4181));
    layer1_outputs(3357) <= (layer0_outputs(3242)) xor (layer0_outputs(2917));
    layer1_outputs(3358) <= not(layer0_outputs(224));
    layer1_outputs(3359) <= layer0_outputs(4472);
    layer1_outputs(3360) <= layer0_outputs(2601);
    layer1_outputs(3361) <= not((layer0_outputs(1244)) and (layer0_outputs(2057)));
    layer1_outputs(3362) <= not(layer0_outputs(4827));
    layer1_outputs(3363) <= (layer0_outputs(2424)) and not (layer0_outputs(1299));
    layer1_outputs(3364) <= not((layer0_outputs(344)) xor (layer0_outputs(4554)));
    layer1_outputs(3365) <= layer0_outputs(2452);
    layer1_outputs(3366) <= not((layer0_outputs(3016)) and (layer0_outputs(4162)));
    layer1_outputs(3367) <= layer0_outputs(4183);
    layer1_outputs(3368) <= not(layer0_outputs(1715));
    layer1_outputs(3369) <= layer0_outputs(255);
    layer1_outputs(3370) <= (layer0_outputs(3670)) or (layer0_outputs(3966));
    layer1_outputs(3371) <= not(layer0_outputs(248));
    layer1_outputs(3372) <= not(layer0_outputs(1419)) or (layer0_outputs(1073));
    layer1_outputs(3373) <= layer0_outputs(2611);
    layer1_outputs(3374) <= not((layer0_outputs(1562)) and (layer0_outputs(539)));
    layer1_outputs(3375) <= not(layer0_outputs(2941)) or (layer0_outputs(2556));
    layer1_outputs(3376) <= not(layer0_outputs(5112));
    layer1_outputs(3377) <= not(layer0_outputs(1011)) or (layer0_outputs(3446));
    layer1_outputs(3378) <= (layer0_outputs(3257)) and (layer0_outputs(3530));
    layer1_outputs(3379) <= not(layer0_outputs(661));
    layer1_outputs(3380) <= (layer0_outputs(4366)) and not (layer0_outputs(35));
    layer1_outputs(3381) <= not(layer0_outputs(342)) or (layer0_outputs(373));
    layer1_outputs(3382) <= (layer0_outputs(3166)) or (layer0_outputs(3049));
    layer1_outputs(3383) <= not((layer0_outputs(4482)) xor (layer0_outputs(969)));
    layer1_outputs(3384) <= not((layer0_outputs(3889)) xor (layer0_outputs(699)));
    layer1_outputs(3385) <= '0';
    layer1_outputs(3386) <= not(layer0_outputs(3188));
    layer1_outputs(3387) <= layer0_outputs(420);
    layer1_outputs(3388) <= '0';
    layer1_outputs(3389) <= (layer0_outputs(2502)) and not (layer0_outputs(2797));
    layer1_outputs(3390) <= layer0_outputs(597);
    layer1_outputs(3391) <= not((layer0_outputs(1919)) xor (layer0_outputs(131)));
    layer1_outputs(3392) <= not((layer0_outputs(4176)) or (layer0_outputs(2354)));
    layer1_outputs(3393) <= layer0_outputs(5082);
    layer1_outputs(3394) <= not(layer0_outputs(4783));
    layer1_outputs(3395) <= (layer0_outputs(4487)) and not (layer0_outputs(1583));
    layer1_outputs(3396) <= (layer0_outputs(1835)) xor (layer0_outputs(2334));
    layer1_outputs(3397) <= (layer0_outputs(2789)) or (layer0_outputs(2901));
    layer1_outputs(3398) <= not(layer0_outputs(5106));
    layer1_outputs(3399) <= layer0_outputs(3676);
    layer1_outputs(3400) <= not((layer0_outputs(2514)) or (layer0_outputs(3614)));
    layer1_outputs(3401) <= not((layer0_outputs(2810)) or (layer0_outputs(2210)));
    layer1_outputs(3402) <= layer0_outputs(4312);
    layer1_outputs(3403) <= not(layer0_outputs(4694));
    layer1_outputs(3404) <= layer0_outputs(3490);
    layer1_outputs(3405) <= (layer0_outputs(3041)) and not (layer0_outputs(4168));
    layer1_outputs(3406) <= layer0_outputs(4681);
    layer1_outputs(3407) <= (layer0_outputs(2267)) xor (layer0_outputs(2140));
    layer1_outputs(3408) <= layer0_outputs(746);
    layer1_outputs(3409) <= not(layer0_outputs(3977));
    layer1_outputs(3410) <= not(layer0_outputs(78));
    layer1_outputs(3411) <= (layer0_outputs(1581)) xor (layer0_outputs(1335));
    layer1_outputs(3412) <= '1';
    layer1_outputs(3413) <= (layer0_outputs(2280)) xor (layer0_outputs(1595));
    layer1_outputs(3414) <= (layer0_outputs(1970)) or (layer0_outputs(4656));
    layer1_outputs(3415) <= not(layer0_outputs(2872));
    layer1_outputs(3416) <= not(layer0_outputs(4942)) or (layer0_outputs(2279));
    layer1_outputs(3417) <= not(layer0_outputs(464));
    layer1_outputs(3418) <= not((layer0_outputs(2473)) xor (layer0_outputs(746)));
    layer1_outputs(3419) <= not((layer0_outputs(4291)) and (layer0_outputs(3640)));
    layer1_outputs(3420) <= not(layer0_outputs(3014));
    layer1_outputs(3421) <= (layer0_outputs(1327)) and (layer0_outputs(1283));
    layer1_outputs(3422) <= not(layer0_outputs(4510)) or (layer0_outputs(4256));
    layer1_outputs(3423) <= (layer0_outputs(2891)) xor (layer0_outputs(1380));
    layer1_outputs(3424) <= not((layer0_outputs(4195)) xor (layer0_outputs(820)));
    layer1_outputs(3425) <= (layer0_outputs(3434)) and not (layer0_outputs(2263));
    layer1_outputs(3426) <= not((layer0_outputs(4982)) and (layer0_outputs(4680)));
    layer1_outputs(3427) <= not(layer0_outputs(1753)) or (layer0_outputs(3058));
    layer1_outputs(3428) <= not((layer0_outputs(997)) xor (layer0_outputs(1611)));
    layer1_outputs(3429) <= not(layer0_outputs(787)) or (layer0_outputs(3356));
    layer1_outputs(3430) <= '1';
    layer1_outputs(3431) <= layer0_outputs(3466);
    layer1_outputs(3432) <= layer0_outputs(4994);
    layer1_outputs(3433) <= not(layer0_outputs(3581)) or (layer0_outputs(2554));
    layer1_outputs(3434) <= not((layer0_outputs(4768)) or (layer0_outputs(3068)));
    layer1_outputs(3435) <= (layer0_outputs(2696)) and not (layer0_outputs(1051));
    layer1_outputs(3436) <= not(layer0_outputs(4465));
    layer1_outputs(3437) <= not((layer0_outputs(1932)) and (layer0_outputs(104)));
    layer1_outputs(3438) <= '1';
    layer1_outputs(3439) <= (layer0_outputs(1654)) or (layer0_outputs(1262));
    layer1_outputs(3440) <= not((layer0_outputs(4542)) or (layer0_outputs(355)));
    layer1_outputs(3441) <= not(layer0_outputs(4361));
    layer1_outputs(3442) <= not(layer0_outputs(1959)) or (layer0_outputs(3699));
    layer1_outputs(3443) <= not(layer0_outputs(364));
    layer1_outputs(3444) <= not(layer0_outputs(3301)) or (layer0_outputs(4554));
    layer1_outputs(3445) <= (layer0_outputs(916)) xor (layer0_outputs(4249));
    layer1_outputs(3446) <= layer0_outputs(429);
    layer1_outputs(3447) <= not(layer0_outputs(3952));
    layer1_outputs(3448) <= (layer0_outputs(2823)) and (layer0_outputs(2030));
    layer1_outputs(3449) <= (layer0_outputs(2269)) or (layer0_outputs(2641));
    layer1_outputs(3450) <= (layer0_outputs(2169)) or (layer0_outputs(4227));
    layer1_outputs(3451) <= (layer0_outputs(5078)) and (layer0_outputs(3306));
    layer1_outputs(3452) <= not((layer0_outputs(1594)) xor (layer0_outputs(658)));
    layer1_outputs(3453) <= not(layer0_outputs(4295));
    layer1_outputs(3454) <= not((layer0_outputs(1646)) and (layer0_outputs(557)));
    layer1_outputs(3455) <= (layer0_outputs(4775)) and not (layer0_outputs(1320));
    layer1_outputs(3456) <= (layer0_outputs(3890)) xor (layer0_outputs(2691));
    layer1_outputs(3457) <= not(layer0_outputs(2549)) or (layer0_outputs(2290));
    layer1_outputs(3458) <= (layer0_outputs(4805)) xor (layer0_outputs(4456));
    layer1_outputs(3459) <= (layer0_outputs(4105)) xor (layer0_outputs(3788));
    layer1_outputs(3460) <= '0';
    layer1_outputs(3461) <= (layer0_outputs(3499)) and not (layer0_outputs(5107));
    layer1_outputs(3462) <= layer0_outputs(105);
    layer1_outputs(3463) <= not(layer0_outputs(4962)) or (layer0_outputs(4753));
    layer1_outputs(3464) <= (layer0_outputs(2309)) or (layer0_outputs(4960));
    layer1_outputs(3465) <= not((layer0_outputs(492)) xor (layer0_outputs(4456)));
    layer1_outputs(3466) <= (layer0_outputs(3886)) and not (layer0_outputs(602));
    layer1_outputs(3467) <= not(layer0_outputs(820)) or (layer0_outputs(4723));
    layer1_outputs(3468) <= layer0_outputs(792);
    layer1_outputs(3469) <= not(layer0_outputs(758));
    layer1_outputs(3470) <= layer0_outputs(304);
    layer1_outputs(3471) <= not((layer0_outputs(209)) and (layer0_outputs(3150)));
    layer1_outputs(3472) <= not(layer0_outputs(1077));
    layer1_outputs(3473) <= layer0_outputs(456);
    layer1_outputs(3474) <= (layer0_outputs(1187)) or (layer0_outputs(925));
    layer1_outputs(3475) <= not(layer0_outputs(278));
    layer1_outputs(3476) <= (layer0_outputs(2815)) and not (layer0_outputs(767));
    layer1_outputs(3477) <= not((layer0_outputs(2206)) and (layer0_outputs(2156)));
    layer1_outputs(3478) <= not(layer0_outputs(4543)) or (layer0_outputs(3290));
    layer1_outputs(3479) <= (layer0_outputs(2403)) and not (layer0_outputs(3241));
    layer1_outputs(3480) <= (layer0_outputs(3139)) and not (layer0_outputs(2467));
    layer1_outputs(3481) <= layer0_outputs(155);
    layer1_outputs(3482) <= not(layer0_outputs(4965));
    layer1_outputs(3483) <= not(layer0_outputs(185));
    layer1_outputs(3484) <= layer0_outputs(3790);
    layer1_outputs(3485) <= not(layer0_outputs(2586));
    layer1_outputs(3486) <= layer0_outputs(3866);
    layer1_outputs(3487) <= (layer0_outputs(1512)) and (layer0_outputs(3329));
    layer1_outputs(3488) <= not(layer0_outputs(926));
    layer1_outputs(3489) <= not(layer0_outputs(1773)) or (layer0_outputs(735));
    layer1_outputs(3490) <= not(layer0_outputs(391));
    layer1_outputs(3491) <= not(layer0_outputs(178));
    layer1_outputs(3492) <= '1';
    layer1_outputs(3493) <= (layer0_outputs(3752)) and not (layer0_outputs(3377));
    layer1_outputs(3494) <= (layer0_outputs(5115)) and (layer0_outputs(3210));
    layer1_outputs(3495) <= not(layer0_outputs(3616));
    layer1_outputs(3496) <= (layer0_outputs(911)) and not (layer0_outputs(4033));
    layer1_outputs(3497) <= (layer0_outputs(5057)) xor (layer0_outputs(165));
    layer1_outputs(3498) <= layer0_outputs(1102);
    layer1_outputs(3499) <= layer0_outputs(622);
    layer1_outputs(3500) <= (layer0_outputs(2168)) xor (layer0_outputs(1550));
    layer1_outputs(3501) <= layer0_outputs(333);
    layer1_outputs(3502) <= not((layer0_outputs(4370)) and (layer0_outputs(1920)));
    layer1_outputs(3503) <= not(layer0_outputs(4378)) or (layer0_outputs(2445));
    layer1_outputs(3504) <= (layer0_outputs(1795)) or (layer0_outputs(1484));
    layer1_outputs(3505) <= not((layer0_outputs(4790)) and (layer0_outputs(4441)));
    layer1_outputs(3506) <= (layer0_outputs(470)) and not (layer0_outputs(5064));
    layer1_outputs(3507) <= layer0_outputs(734);
    layer1_outputs(3508) <= not((layer0_outputs(1628)) or (layer0_outputs(3983)));
    layer1_outputs(3509) <= not(layer0_outputs(972));
    layer1_outputs(3510) <= '1';
    layer1_outputs(3511) <= not((layer0_outputs(2930)) and (layer0_outputs(397)));
    layer1_outputs(3512) <= not((layer0_outputs(1559)) and (layer0_outputs(3689)));
    layer1_outputs(3513) <= (layer0_outputs(199)) and not (layer0_outputs(1175));
    layer1_outputs(3514) <= (layer0_outputs(921)) and (layer0_outputs(2039));
    layer1_outputs(3515) <= not(layer0_outputs(316));
    layer1_outputs(3516) <= (layer0_outputs(4630)) and (layer0_outputs(2124));
    layer1_outputs(3517) <= (layer0_outputs(3787)) and not (layer0_outputs(440));
    layer1_outputs(3518) <= not((layer0_outputs(4959)) xor (layer0_outputs(358)));
    layer1_outputs(3519) <= (layer0_outputs(4514)) or (layer0_outputs(4279));
    layer1_outputs(3520) <= (layer0_outputs(1411)) xor (layer0_outputs(5100));
    layer1_outputs(3521) <= layer0_outputs(1410);
    layer1_outputs(3522) <= not((layer0_outputs(783)) or (layer0_outputs(482)));
    layer1_outputs(3523) <= not(layer0_outputs(4254));
    layer1_outputs(3524) <= not(layer0_outputs(3517));
    layer1_outputs(3525) <= (layer0_outputs(649)) and not (layer0_outputs(1967));
    layer1_outputs(3526) <= layer0_outputs(2915);
    layer1_outputs(3527) <= (layer0_outputs(2735)) or (layer0_outputs(3868));
    layer1_outputs(3528) <= not(layer0_outputs(4512));
    layer1_outputs(3529) <= (layer0_outputs(4443)) and not (layer0_outputs(4225));
    layer1_outputs(3530) <= not(layer0_outputs(2033)) or (layer0_outputs(2712));
    layer1_outputs(3531) <= (layer0_outputs(3167)) and not (layer0_outputs(5083));
    layer1_outputs(3532) <= not(layer0_outputs(2687)) or (layer0_outputs(3681));
    layer1_outputs(3533) <= not(layer0_outputs(1361)) or (layer0_outputs(3562));
    layer1_outputs(3534) <= not(layer0_outputs(1025));
    layer1_outputs(3535) <= (layer0_outputs(5113)) and (layer0_outputs(294));
    layer1_outputs(3536) <= (layer0_outputs(870)) or (layer0_outputs(3097));
    layer1_outputs(3537) <= layer0_outputs(4573);
    layer1_outputs(3538) <= (layer0_outputs(2501)) and not (layer0_outputs(542));
    layer1_outputs(3539) <= layer0_outputs(4871);
    layer1_outputs(3540) <= (layer0_outputs(1351)) or (layer0_outputs(1370));
    layer1_outputs(3541) <= not(layer0_outputs(3761)) or (layer0_outputs(712));
    layer1_outputs(3542) <= not(layer0_outputs(1160)) or (layer0_outputs(202));
    layer1_outputs(3543) <= layer0_outputs(4080);
    layer1_outputs(3544) <= not(layer0_outputs(3319));
    layer1_outputs(3545) <= (layer0_outputs(4435)) and not (layer0_outputs(15));
    layer1_outputs(3546) <= not(layer0_outputs(2961));
    layer1_outputs(3547) <= (layer0_outputs(2126)) and not (layer0_outputs(423));
    layer1_outputs(3548) <= not(layer0_outputs(1959));
    layer1_outputs(3549) <= (layer0_outputs(3721)) and not (layer0_outputs(2181));
    layer1_outputs(3550) <= not(layer0_outputs(4961));
    layer1_outputs(3551) <= (layer0_outputs(3325)) and not (layer0_outputs(2484));
    layer1_outputs(3552) <= (layer0_outputs(4206)) xor (layer0_outputs(3173));
    layer1_outputs(3553) <= layer0_outputs(4133);
    layer1_outputs(3554) <= (layer0_outputs(4237)) and (layer0_outputs(440));
    layer1_outputs(3555) <= not((layer0_outputs(3954)) xor (layer0_outputs(325)));
    layer1_outputs(3556) <= (layer0_outputs(3832)) or (layer0_outputs(4240));
    layer1_outputs(3557) <= not(layer0_outputs(3503));
    layer1_outputs(3558) <= not((layer0_outputs(1985)) or (layer0_outputs(4844)));
    layer1_outputs(3559) <= '1';
    layer1_outputs(3560) <= not(layer0_outputs(3448)) or (layer0_outputs(16));
    layer1_outputs(3561) <= layer0_outputs(3693);
    layer1_outputs(3562) <= not(layer0_outputs(2315));
    layer1_outputs(3563) <= (layer0_outputs(1288)) or (layer0_outputs(3061));
    layer1_outputs(3564) <= (layer0_outputs(2061)) xor (layer0_outputs(1642));
    layer1_outputs(3565) <= not(layer0_outputs(422)) or (layer0_outputs(4440));
    layer1_outputs(3566) <= not(layer0_outputs(4957)) or (layer0_outputs(3349));
    layer1_outputs(3567) <= layer0_outputs(1113);
    layer1_outputs(3568) <= layer0_outputs(4387);
    layer1_outputs(3569) <= not(layer0_outputs(1862));
    layer1_outputs(3570) <= not((layer0_outputs(217)) or (layer0_outputs(2426)));
    layer1_outputs(3571) <= '1';
    layer1_outputs(3572) <= not((layer0_outputs(2215)) or (layer0_outputs(1809)));
    layer1_outputs(3573) <= not(layer0_outputs(4334)) or (layer0_outputs(3739));
    layer1_outputs(3574) <= not(layer0_outputs(2005));
    layer1_outputs(3575) <= layer0_outputs(88);
    layer1_outputs(3576) <= not(layer0_outputs(4094));
    layer1_outputs(3577) <= not(layer0_outputs(4637)) or (layer0_outputs(2846));
    layer1_outputs(3578) <= layer0_outputs(4446);
    layer1_outputs(3579) <= not(layer0_outputs(1130));
    layer1_outputs(3580) <= not((layer0_outputs(3879)) and (layer0_outputs(3281)));
    layer1_outputs(3581) <= not(layer0_outputs(2294));
    layer1_outputs(3582) <= layer0_outputs(3360);
    layer1_outputs(3583) <= not(layer0_outputs(2004)) or (layer0_outputs(2011));
    layer1_outputs(3584) <= layer0_outputs(1537);
    layer1_outputs(3585) <= not((layer0_outputs(4487)) xor (layer0_outputs(1185)));
    layer1_outputs(3586) <= '1';
    layer1_outputs(3587) <= (layer0_outputs(1004)) and (layer0_outputs(1361));
    layer1_outputs(3588) <= not((layer0_outputs(3335)) or (layer0_outputs(3688)));
    layer1_outputs(3589) <= (layer0_outputs(3887)) and (layer0_outputs(3647));
    layer1_outputs(3590) <= not((layer0_outputs(3056)) or (layer0_outputs(858)));
    layer1_outputs(3591) <= not((layer0_outputs(785)) and (layer0_outputs(872)));
    layer1_outputs(3592) <= not((layer0_outputs(3999)) and (layer0_outputs(3012)));
    layer1_outputs(3593) <= not(layer0_outputs(5016));
    layer1_outputs(3594) <= not(layer0_outputs(978)) or (layer0_outputs(1475));
    layer1_outputs(3595) <= layer0_outputs(1153);
    layer1_outputs(3596) <= layer0_outputs(3670);
    layer1_outputs(3597) <= '1';
    layer1_outputs(3598) <= not(layer0_outputs(5044)) or (layer0_outputs(322));
    layer1_outputs(3599) <= not(layer0_outputs(3733)) or (layer0_outputs(411));
    layer1_outputs(3600) <= not(layer0_outputs(1193)) or (layer0_outputs(3984));
    layer1_outputs(3601) <= (layer0_outputs(4742)) and (layer0_outputs(3370));
    layer1_outputs(3602) <= (layer0_outputs(4054)) or (layer0_outputs(328));
    layer1_outputs(3603) <= (layer0_outputs(4147)) xor (layer0_outputs(1492));
    layer1_outputs(3604) <= layer0_outputs(1270);
    layer1_outputs(3605) <= (layer0_outputs(4813)) and not (layer0_outputs(3164));
    layer1_outputs(3606) <= layer0_outputs(956);
    layer1_outputs(3607) <= '1';
    layer1_outputs(3608) <= (layer0_outputs(400)) and not (layer0_outputs(680));
    layer1_outputs(3609) <= layer0_outputs(2983);
    layer1_outputs(3610) <= not(layer0_outputs(169));
    layer1_outputs(3611) <= (layer0_outputs(1705)) and (layer0_outputs(3729));
    layer1_outputs(3612) <= layer0_outputs(1648);
    layer1_outputs(3613) <= not(layer0_outputs(890)) or (layer0_outputs(3778));
    layer1_outputs(3614) <= not(layer0_outputs(3265));
    layer1_outputs(3615) <= (layer0_outputs(240)) and (layer0_outputs(2310));
    layer1_outputs(3616) <= (layer0_outputs(2120)) and (layer0_outputs(2257));
    layer1_outputs(3617) <= not((layer0_outputs(1425)) or (layer0_outputs(246)));
    layer1_outputs(3618) <= not(layer0_outputs(3788)) or (layer0_outputs(1159));
    layer1_outputs(3619) <= not(layer0_outputs(2984));
    layer1_outputs(3620) <= (layer0_outputs(851)) and not (layer0_outputs(4541));
    layer1_outputs(3621) <= not((layer0_outputs(3650)) xor (layer0_outputs(3273)));
    layer1_outputs(3622) <= not(layer0_outputs(1123)) or (layer0_outputs(3692));
    layer1_outputs(3623) <= (layer0_outputs(1539)) xor (layer0_outputs(2451));
    layer1_outputs(3624) <= '0';
    layer1_outputs(3625) <= (layer0_outputs(379)) and (layer0_outputs(3835));
    layer1_outputs(3626) <= (layer0_outputs(2831)) and not (layer0_outputs(545));
    layer1_outputs(3627) <= not(layer0_outputs(1742));
    layer1_outputs(3628) <= layer0_outputs(4161);
    layer1_outputs(3629) <= '0';
    layer1_outputs(3630) <= not(layer0_outputs(4543)) or (layer0_outputs(3373));
    layer1_outputs(3631) <= layer0_outputs(3315);
    layer1_outputs(3632) <= (layer0_outputs(505)) and (layer0_outputs(3565));
    layer1_outputs(3633) <= not(layer0_outputs(4830));
    layer1_outputs(3634) <= (layer0_outputs(1126)) and (layer0_outputs(1693));
    layer1_outputs(3635) <= layer0_outputs(4838);
    layer1_outputs(3636) <= not((layer0_outputs(4847)) or (layer0_outputs(2260)));
    layer1_outputs(3637) <= layer0_outputs(3760);
    layer1_outputs(3638) <= (layer0_outputs(4762)) or (layer0_outputs(3579));
    layer1_outputs(3639) <= (layer0_outputs(3206)) or (layer0_outputs(4881));
    layer1_outputs(3640) <= not((layer0_outputs(2113)) or (layer0_outputs(1044)));
    layer1_outputs(3641) <= layer0_outputs(3500);
    layer1_outputs(3642) <= (layer0_outputs(1697)) and (layer0_outputs(4011));
    layer1_outputs(3643) <= not(layer0_outputs(2840));
    layer1_outputs(3644) <= not(layer0_outputs(78));
    layer1_outputs(3645) <= not(layer0_outputs(183));
    layer1_outputs(3646) <= (layer0_outputs(4810)) and not (layer0_outputs(2743));
    layer1_outputs(3647) <= not(layer0_outputs(1403));
    layer1_outputs(3648) <= layer0_outputs(2082);
    layer1_outputs(3649) <= not((layer0_outputs(3493)) or (layer0_outputs(5018)));
    layer1_outputs(3650) <= not(layer0_outputs(4613)) or (layer0_outputs(514));
    layer1_outputs(3651) <= not(layer0_outputs(2253));
    layer1_outputs(3652) <= not((layer0_outputs(4393)) xor (layer0_outputs(4757)));
    layer1_outputs(3653) <= not(layer0_outputs(3901)) or (layer0_outputs(670));
    layer1_outputs(3654) <= not(layer0_outputs(3216));
    layer1_outputs(3655) <= (layer0_outputs(1893)) or (layer0_outputs(2581));
    layer1_outputs(3656) <= layer0_outputs(821);
    layer1_outputs(3657) <= not(layer0_outputs(2873)) or (layer0_outputs(753));
    layer1_outputs(3658) <= not((layer0_outputs(646)) and (layer0_outputs(2217)));
    layer1_outputs(3659) <= (layer0_outputs(228)) and (layer0_outputs(4704));
    layer1_outputs(3660) <= (layer0_outputs(1532)) and not (layer0_outputs(3));
    layer1_outputs(3661) <= (layer0_outputs(4433)) and (layer0_outputs(1232));
    layer1_outputs(3662) <= not(layer0_outputs(811));
    layer1_outputs(3663) <= not(layer0_outputs(4634)) or (layer0_outputs(3748));
    layer1_outputs(3664) <= not((layer0_outputs(3095)) or (layer0_outputs(1976)));
    layer1_outputs(3665) <= '0';
    layer1_outputs(3666) <= (layer0_outputs(1930)) or (layer0_outputs(2258));
    layer1_outputs(3667) <= not(layer0_outputs(569));
    layer1_outputs(3668) <= layer0_outputs(3025);
    layer1_outputs(3669) <= not(layer0_outputs(4980)) or (layer0_outputs(965));
    layer1_outputs(3670) <= not(layer0_outputs(593));
    layer1_outputs(3671) <= layer0_outputs(2865);
    layer1_outputs(3672) <= layer0_outputs(2225);
    layer1_outputs(3673) <= not(layer0_outputs(2149));
    layer1_outputs(3674) <= not(layer0_outputs(1550)) or (layer0_outputs(776));
    layer1_outputs(3675) <= (layer0_outputs(4026)) xor (layer0_outputs(3127));
    layer1_outputs(3676) <= not(layer0_outputs(4586)) or (layer0_outputs(960));
    layer1_outputs(3677) <= (layer0_outputs(644)) xor (layer0_outputs(2302));
    layer1_outputs(3678) <= not((layer0_outputs(4419)) or (layer0_outputs(4645)));
    layer1_outputs(3679) <= not(layer0_outputs(1092));
    layer1_outputs(3680) <= layer0_outputs(618);
    layer1_outputs(3681) <= not(layer0_outputs(4283)) or (layer0_outputs(2830));
    layer1_outputs(3682) <= not((layer0_outputs(474)) xor (layer0_outputs(5012)));
    layer1_outputs(3683) <= (layer0_outputs(5021)) and (layer0_outputs(530));
    layer1_outputs(3684) <= not(layer0_outputs(4730));
    layer1_outputs(3685) <= not(layer0_outputs(2031)) or (layer0_outputs(2281));
    layer1_outputs(3686) <= (layer0_outputs(4434)) and not (layer0_outputs(2728));
    layer1_outputs(3687) <= (layer0_outputs(3797)) or (layer0_outputs(3688));
    layer1_outputs(3688) <= layer0_outputs(4112);
    layer1_outputs(3689) <= not(layer0_outputs(4949));
    layer1_outputs(3690) <= not(layer0_outputs(4679)) or (layer0_outputs(1558));
    layer1_outputs(3691) <= not(layer0_outputs(1491));
    layer1_outputs(3692) <= not(layer0_outputs(1278));
    layer1_outputs(3693) <= (layer0_outputs(2480)) and (layer0_outputs(1055));
    layer1_outputs(3694) <= (layer0_outputs(404)) and not (layer0_outputs(4800));
    layer1_outputs(3695) <= (layer0_outputs(489)) and not (layer0_outputs(3907));
    layer1_outputs(3696) <= not(layer0_outputs(3967)) or (layer0_outputs(1500));
    layer1_outputs(3697) <= (layer0_outputs(1973)) or (layer0_outputs(284));
    layer1_outputs(3698) <= '1';
    layer1_outputs(3699) <= not(layer0_outputs(2010));
    layer1_outputs(3700) <= (layer0_outputs(759)) and not (layer0_outputs(3185));
    layer1_outputs(3701) <= '0';
    layer1_outputs(3702) <= not((layer0_outputs(4236)) or (layer0_outputs(3915)));
    layer1_outputs(3703) <= (layer0_outputs(3010)) or (layer0_outputs(2900));
    layer1_outputs(3704) <= (layer0_outputs(2309)) and (layer0_outputs(3295));
    layer1_outputs(3705) <= not((layer0_outputs(2116)) xor (layer0_outputs(886)));
    layer1_outputs(3706) <= (layer0_outputs(3469)) and not (layer0_outputs(4290));
    layer1_outputs(3707) <= layer0_outputs(108);
    layer1_outputs(3708) <= '0';
    layer1_outputs(3709) <= not(layer0_outputs(1764)) or (layer0_outputs(2496));
    layer1_outputs(3710) <= not(layer0_outputs(1850)) or (layer0_outputs(2918));
    layer1_outputs(3711) <= '0';
    layer1_outputs(3712) <= (layer0_outputs(1707)) and not (layer0_outputs(2322));
    layer1_outputs(3713) <= layer0_outputs(352);
    layer1_outputs(3714) <= layer0_outputs(1421);
    layer1_outputs(3715) <= (layer0_outputs(877)) and not (layer0_outputs(879));
    layer1_outputs(3716) <= not(layer0_outputs(1934));
    layer1_outputs(3717) <= not(layer0_outputs(2157));
    layer1_outputs(3718) <= layer0_outputs(1266);
    layer1_outputs(3719) <= not(layer0_outputs(1388)) or (layer0_outputs(1859));
    layer1_outputs(3720) <= layer0_outputs(2940);
    layer1_outputs(3721) <= not((layer0_outputs(296)) or (layer0_outputs(2773)));
    layer1_outputs(3722) <= not((layer0_outputs(1896)) and (layer0_outputs(4911)));
    layer1_outputs(3723) <= (layer0_outputs(639)) xor (layer0_outputs(4043));
    layer1_outputs(3724) <= not((layer0_outputs(180)) or (layer0_outputs(2635)));
    layer1_outputs(3725) <= not(layer0_outputs(2364)) or (layer0_outputs(1814));
    layer1_outputs(3726) <= (layer0_outputs(4849)) and not (layer0_outputs(448));
    layer1_outputs(3727) <= not(layer0_outputs(1366));
    layer1_outputs(3728) <= layer0_outputs(1250);
    layer1_outputs(3729) <= not(layer0_outputs(4997)) or (layer0_outputs(4685));
    layer1_outputs(3730) <= layer0_outputs(3889);
    layer1_outputs(3731) <= (layer0_outputs(586)) or (layer0_outputs(2632));
    layer1_outputs(3732) <= not(layer0_outputs(740)) or (layer0_outputs(4743));
    layer1_outputs(3733) <= layer0_outputs(1446);
    layer1_outputs(3734) <= (layer0_outputs(1729)) or (layer0_outputs(3382));
    layer1_outputs(3735) <= not((layer0_outputs(3753)) and (layer0_outputs(1906)));
    layer1_outputs(3736) <= not((layer0_outputs(208)) and (layer0_outputs(2722)));
    layer1_outputs(3737) <= (layer0_outputs(4261)) or (layer0_outputs(3385));
    layer1_outputs(3738) <= not((layer0_outputs(1629)) or (layer0_outputs(4038)));
    layer1_outputs(3739) <= not(layer0_outputs(3099)) or (layer0_outputs(574));
    layer1_outputs(3740) <= layer0_outputs(2529);
    layer1_outputs(3741) <= not(layer0_outputs(2939)) or (layer0_outputs(2209));
    layer1_outputs(3742) <= layer0_outputs(640);
    layer1_outputs(3743) <= layer0_outputs(1021);
    layer1_outputs(3744) <= layer0_outputs(1577);
    layer1_outputs(3745) <= not(layer0_outputs(3334));
    layer1_outputs(3746) <= not(layer0_outputs(1208));
    layer1_outputs(3747) <= not(layer0_outputs(2128));
    layer1_outputs(3748) <= not(layer0_outputs(2237)) or (layer0_outputs(1998));
    layer1_outputs(3749) <= not((layer0_outputs(2779)) xor (layer0_outputs(330)));
    layer1_outputs(3750) <= not(layer0_outputs(1047)) or (layer0_outputs(2847));
    layer1_outputs(3751) <= layer0_outputs(2551);
    layer1_outputs(3752) <= layer0_outputs(3990);
    layer1_outputs(3753) <= (layer0_outputs(4391)) and not (layer0_outputs(1636));
    layer1_outputs(3754) <= not(layer0_outputs(2627));
    layer1_outputs(3755) <= (layer0_outputs(1247)) and not (layer0_outputs(274));
    layer1_outputs(3756) <= (layer0_outputs(3078)) and (layer0_outputs(154));
    layer1_outputs(3757) <= (layer0_outputs(3777)) xor (layer0_outputs(4251));
    layer1_outputs(3758) <= not(layer0_outputs(1430));
    layer1_outputs(3759) <= (layer0_outputs(3326)) or (layer0_outputs(1972));
    layer1_outputs(3760) <= (layer0_outputs(3836)) and not (layer0_outputs(2842));
    layer1_outputs(3761) <= not(layer0_outputs(1145));
    layer1_outputs(3762) <= not(layer0_outputs(1408)) or (layer0_outputs(4326));
    layer1_outputs(3763) <= layer0_outputs(4271);
    layer1_outputs(3764) <= (layer0_outputs(1381)) and not (layer0_outputs(5097));
    layer1_outputs(3765) <= '0';
    layer1_outputs(3766) <= layer0_outputs(490);
    layer1_outputs(3767) <= layer0_outputs(143);
    layer1_outputs(3768) <= layer0_outputs(1850);
    layer1_outputs(3769) <= not((layer0_outputs(3956)) and (layer0_outputs(1647)));
    layer1_outputs(3770) <= not(layer0_outputs(154));
    layer1_outputs(3771) <= not((layer0_outputs(3623)) or (layer0_outputs(4878)));
    layer1_outputs(3772) <= (layer0_outputs(897)) and not (layer0_outputs(394));
    layer1_outputs(3773) <= '1';
    layer1_outputs(3774) <= layer0_outputs(944);
    layer1_outputs(3775) <= (layer0_outputs(527)) and (layer0_outputs(1834));
    layer1_outputs(3776) <= layer0_outputs(2612);
    layer1_outputs(3777) <= layer0_outputs(1974);
    layer1_outputs(3778) <= not(layer0_outputs(2468));
    layer1_outputs(3779) <= not(layer0_outputs(3285));
    layer1_outputs(3780) <= layer0_outputs(4534);
    layer1_outputs(3781) <= layer0_outputs(3533);
    layer1_outputs(3782) <= not(layer0_outputs(2049));
    layer1_outputs(3783) <= (layer0_outputs(1776)) xor (layer0_outputs(5106));
    layer1_outputs(3784) <= (layer0_outputs(4307)) and not (layer0_outputs(4441));
    layer1_outputs(3785) <= (layer0_outputs(4423)) and not (layer0_outputs(4876));
    layer1_outputs(3786) <= layer0_outputs(1199);
    layer1_outputs(3787) <= (layer0_outputs(2170)) and (layer0_outputs(3583));
    layer1_outputs(3788) <= (layer0_outputs(496)) and not (layer0_outputs(3308));
    layer1_outputs(3789) <= not(layer0_outputs(1040));
    layer1_outputs(3790) <= not(layer0_outputs(4853)) or (layer0_outputs(1964));
    layer1_outputs(3791) <= not((layer0_outputs(2432)) and (layer0_outputs(1455)));
    layer1_outputs(3792) <= not((layer0_outputs(4811)) or (layer0_outputs(2894)));
    layer1_outputs(3793) <= (layer0_outputs(3307)) or (layer0_outputs(4914));
    layer1_outputs(3794) <= not((layer0_outputs(3448)) and (layer0_outputs(2804)));
    layer1_outputs(3795) <= (layer0_outputs(2478)) and (layer0_outputs(3347));
    layer1_outputs(3796) <= (layer0_outputs(3380)) and not (layer0_outputs(1659));
    layer1_outputs(3797) <= layer0_outputs(4801);
    layer1_outputs(3798) <= (layer0_outputs(3687)) and not (layer0_outputs(2138));
    layer1_outputs(3799) <= (layer0_outputs(183)) or (layer0_outputs(1423));
    layer1_outputs(3800) <= not(layer0_outputs(918)) or (layer0_outputs(5028));
    layer1_outputs(3801) <= (layer0_outputs(2397)) or (layer0_outputs(5054));
    layer1_outputs(3802) <= not(layer0_outputs(957)) or (layer0_outputs(604));
    layer1_outputs(3803) <= (layer0_outputs(4496)) and not (layer0_outputs(4923));
    layer1_outputs(3804) <= '0';
    layer1_outputs(3805) <= (layer0_outputs(1858)) or (layer0_outputs(3793));
    layer1_outputs(3806) <= not((layer0_outputs(2020)) xor (layer0_outputs(61)));
    layer1_outputs(3807) <= not(layer0_outputs(1121)) or (layer0_outputs(2547));
    layer1_outputs(3808) <= not(layer0_outputs(1338)) or (layer0_outputs(615));
    layer1_outputs(3809) <= not(layer0_outputs(3578));
    layer1_outputs(3810) <= not((layer0_outputs(771)) xor (layer0_outputs(1437)));
    layer1_outputs(3811) <= (layer0_outputs(3958)) and not (layer0_outputs(96));
    layer1_outputs(3812) <= not((layer0_outputs(2880)) xor (layer0_outputs(2770)));
    layer1_outputs(3813) <= (layer0_outputs(3611)) and not (layer0_outputs(2277));
    layer1_outputs(3814) <= '1';
    layer1_outputs(3815) <= (layer0_outputs(2509)) and not (layer0_outputs(1210));
    layer1_outputs(3816) <= not((layer0_outputs(3777)) xor (layer0_outputs(2841)));
    layer1_outputs(3817) <= not((layer0_outputs(2643)) xor (layer0_outputs(495)));
    layer1_outputs(3818) <= not((layer0_outputs(2590)) or (layer0_outputs(4343)));
    layer1_outputs(3819) <= layer0_outputs(1642);
    layer1_outputs(3820) <= (layer0_outputs(2887)) xor (layer0_outputs(2797));
    layer1_outputs(3821) <= (layer0_outputs(3509)) and not (layer0_outputs(658));
    layer1_outputs(3822) <= (layer0_outputs(4592)) and (layer0_outputs(4082));
    layer1_outputs(3823) <= not(layer0_outputs(998)) or (layer0_outputs(5050));
    layer1_outputs(3824) <= layer0_outputs(841);
    layer1_outputs(3825) <= not(layer0_outputs(1158)) or (layer0_outputs(2219));
    layer1_outputs(3826) <= layer0_outputs(2166);
    layer1_outputs(3827) <= '1';
    layer1_outputs(3828) <= not(layer0_outputs(1389)) or (layer0_outputs(3580));
    layer1_outputs(3829) <= layer0_outputs(4219);
    layer1_outputs(3830) <= (layer0_outputs(2859)) and not (layer0_outputs(360));
    layer1_outputs(3831) <= (layer0_outputs(2284)) and not (layer0_outputs(3795));
    layer1_outputs(3832) <= layer0_outputs(3587);
    layer1_outputs(3833) <= not(layer0_outputs(4326)) or (layer0_outputs(3175));
    layer1_outputs(3834) <= (layer0_outputs(399)) and not (layer0_outputs(3138));
    layer1_outputs(3835) <= not(layer0_outputs(3705));
    layer1_outputs(3836) <= (layer0_outputs(4856)) xor (layer0_outputs(2474));
    layer1_outputs(3837) <= not(layer0_outputs(4898));
    layer1_outputs(3838) <= not((layer0_outputs(4655)) or (layer0_outputs(3911)));
    layer1_outputs(3839) <= not(layer0_outputs(2497));
    layer1_outputs(3840) <= not(layer0_outputs(2266));
    layer1_outputs(3841) <= (layer0_outputs(3007)) and (layer0_outputs(2879));
    layer1_outputs(3842) <= not((layer0_outputs(1658)) xor (layer0_outputs(992)));
    layer1_outputs(3843) <= not((layer0_outputs(1292)) or (layer0_outputs(3567)));
    layer1_outputs(3844) <= not((layer0_outputs(3018)) or (layer0_outputs(3053)));
    layer1_outputs(3845) <= not((layer0_outputs(4142)) xor (layer0_outputs(2575)));
    layer1_outputs(3846) <= layer0_outputs(829);
    layer1_outputs(3847) <= not(layer0_outputs(2155));
    layer1_outputs(3848) <= (layer0_outputs(3410)) and not (layer0_outputs(2289));
    layer1_outputs(3849) <= layer0_outputs(1238);
    layer1_outputs(3850) <= not((layer0_outputs(401)) and (layer0_outputs(5070)));
    layer1_outputs(3851) <= (layer0_outputs(2937)) and not (layer0_outputs(26));
    layer1_outputs(3852) <= layer0_outputs(762);
    layer1_outputs(3853) <= not(layer0_outputs(4159)) or (layer0_outputs(700));
    layer1_outputs(3854) <= layer0_outputs(3820);
    layer1_outputs(3855) <= not(layer0_outputs(834));
    layer1_outputs(3856) <= (layer0_outputs(3473)) xor (layer0_outputs(4070));
    layer1_outputs(3857) <= not(layer0_outputs(1284)) or (layer0_outputs(4900));
    layer1_outputs(3858) <= not((layer0_outputs(3866)) and (layer0_outputs(4906)));
    layer1_outputs(3859) <= layer0_outputs(591);
    layer1_outputs(3860) <= not(layer0_outputs(4916));
    layer1_outputs(3861) <= not(layer0_outputs(2636));
    layer1_outputs(3862) <= (layer0_outputs(3846)) and not (layer0_outputs(3129));
    layer1_outputs(3863) <= layer0_outputs(1650);
    layer1_outputs(3864) <= not(layer0_outputs(498));
    layer1_outputs(3865) <= layer0_outputs(533);
    layer1_outputs(3866) <= (layer0_outputs(1149)) and not (layer0_outputs(3912));
    layer1_outputs(3867) <= layer0_outputs(2708);
    layer1_outputs(3868) <= (layer0_outputs(3792)) and not (layer0_outputs(4814));
    layer1_outputs(3869) <= (layer0_outputs(281)) and not (layer0_outputs(4624));
    layer1_outputs(3870) <= not(layer0_outputs(2060)) or (layer0_outputs(1756));
    layer1_outputs(3871) <= (layer0_outputs(4345)) and (layer0_outputs(849));
    layer1_outputs(3872) <= (layer0_outputs(2699)) or (layer0_outputs(2439));
    layer1_outputs(3873) <= layer0_outputs(1820);
    layer1_outputs(3874) <= not(layer0_outputs(675));
    layer1_outputs(3875) <= (layer0_outputs(1749)) or (layer0_outputs(439));
    layer1_outputs(3876) <= not(layer0_outputs(1702));
    layer1_outputs(3877) <= (layer0_outputs(2609)) and not (layer0_outputs(2905));
    layer1_outputs(3878) <= (layer0_outputs(4078)) and not (layer0_outputs(3767));
    layer1_outputs(3879) <= (layer0_outputs(1938)) and not (layer0_outputs(1334));
    layer1_outputs(3880) <= not(layer0_outputs(1732)) or (layer0_outputs(2031));
    layer1_outputs(3881) <= not(layer0_outputs(1499));
    layer1_outputs(3882) <= (layer0_outputs(5076)) xor (layer0_outputs(821));
    layer1_outputs(3883) <= (layer0_outputs(287)) and (layer0_outputs(3525));
    layer1_outputs(3884) <= layer0_outputs(3380);
    layer1_outputs(3885) <= not((layer0_outputs(898)) or (layer0_outputs(553)));
    layer1_outputs(3886) <= (layer0_outputs(4657)) or (layer0_outputs(4704));
    layer1_outputs(3887) <= (layer0_outputs(2543)) and not (layer0_outputs(3338));
    layer1_outputs(3888) <= '0';
    layer1_outputs(3889) <= not((layer0_outputs(4580)) xor (layer0_outputs(800)));
    layer1_outputs(3890) <= not((layer0_outputs(749)) xor (layer0_outputs(2541)));
    layer1_outputs(3891) <= not(layer0_outputs(4023));
    layer1_outputs(3892) <= (layer0_outputs(4571)) and not (layer0_outputs(2631));
    layer1_outputs(3893) <= (layer0_outputs(1645)) and (layer0_outputs(4536));
    layer1_outputs(3894) <= (layer0_outputs(389)) and not (layer0_outputs(4888));
    layer1_outputs(3895) <= not(layer0_outputs(473));
    layer1_outputs(3896) <= '1';
    layer1_outputs(3897) <= not(layer0_outputs(840));
    layer1_outputs(3898) <= not(layer0_outputs(4990)) or (layer0_outputs(1161));
    layer1_outputs(3899) <= layer0_outputs(782);
    layer1_outputs(3900) <= not(layer0_outputs(2580)) or (layer0_outputs(2163));
    layer1_outputs(3901) <= layer0_outputs(825);
    layer1_outputs(3902) <= not(layer0_outputs(3416));
    layer1_outputs(3903) <= (layer0_outputs(4103)) and (layer0_outputs(1372));
    layer1_outputs(3904) <= (layer0_outputs(3516)) and not (layer0_outputs(469));
    layer1_outputs(3905) <= not(layer0_outputs(2227));
    layer1_outputs(3906) <= not(layer0_outputs(1358));
    layer1_outputs(3907) <= not(layer0_outputs(1487));
    layer1_outputs(3908) <= not((layer0_outputs(2305)) xor (layer0_outputs(4587)));
    layer1_outputs(3909) <= (layer0_outputs(1223)) and not (layer0_outputs(3093));
    layer1_outputs(3910) <= (layer0_outputs(1300)) and (layer0_outputs(231));
    layer1_outputs(3911) <= not(layer0_outputs(2425));
    layer1_outputs(3912) <= '0';
    layer1_outputs(3913) <= not(layer0_outputs(691)) or (layer0_outputs(1461));
    layer1_outputs(3914) <= (layer0_outputs(2494)) xor (layer0_outputs(83));
    layer1_outputs(3915) <= not(layer0_outputs(2747));
    layer1_outputs(3916) <= not((layer0_outputs(187)) or (layer0_outputs(130)));
    layer1_outputs(3917) <= layer0_outputs(1081);
    layer1_outputs(3918) <= (layer0_outputs(500)) or (layer0_outputs(3782));
    layer1_outputs(3919) <= not(layer0_outputs(1928)) or (layer0_outputs(830));
    layer1_outputs(3920) <= not(layer0_outputs(2804));
    layer1_outputs(3921) <= (layer0_outputs(2461)) or (layer0_outputs(1636));
    layer1_outputs(3922) <= (layer0_outputs(3183)) xor (layer0_outputs(2818));
    layer1_outputs(3923) <= not((layer0_outputs(3937)) or (layer0_outputs(839)));
    layer1_outputs(3924) <= layer0_outputs(4887);
    layer1_outputs(3925) <= (layer0_outputs(1652)) xor (layer0_outputs(3279));
    layer1_outputs(3926) <= not(layer0_outputs(313)) or (layer0_outputs(1741));
    layer1_outputs(3927) <= not(layer0_outputs(4633));
    layer1_outputs(3928) <= layer0_outputs(634);
    layer1_outputs(3929) <= not(layer0_outputs(3581));
    layer1_outputs(3930) <= (layer0_outputs(2249)) and not (layer0_outputs(547));
    layer1_outputs(3931) <= not(layer0_outputs(583));
    layer1_outputs(3932) <= not((layer0_outputs(4496)) and (layer0_outputs(116)));
    layer1_outputs(3933) <= not(layer0_outputs(1811));
    layer1_outputs(3934) <= not(layer0_outputs(3976));
    layer1_outputs(3935) <= '0';
    layer1_outputs(3936) <= not((layer0_outputs(4745)) xor (layer0_outputs(1079)));
    layer1_outputs(3937) <= not((layer0_outputs(4328)) or (layer0_outputs(2595)));
    layer1_outputs(3938) <= not(layer0_outputs(819)) or (layer0_outputs(3703));
    layer1_outputs(3939) <= layer0_outputs(4994);
    layer1_outputs(3940) <= layer0_outputs(685);
    layer1_outputs(3941) <= not(layer0_outputs(1231));
    layer1_outputs(3942) <= (layer0_outputs(3003)) and not (layer0_outputs(3181));
    layer1_outputs(3943) <= (layer0_outputs(3172)) or (layer0_outputs(1166));
    layer1_outputs(3944) <= (layer0_outputs(3476)) or (layer0_outputs(1736));
    layer1_outputs(3945) <= not(layer0_outputs(4394)) or (layer0_outputs(698));
    layer1_outputs(3946) <= not(layer0_outputs(5116));
    layer1_outputs(3947) <= (layer0_outputs(4166)) and not (layer0_outputs(2266));
    layer1_outputs(3948) <= (layer0_outputs(2185)) or (layer0_outputs(522));
    layer1_outputs(3949) <= not((layer0_outputs(3239)) xor (layer0_outputs(3885)));
    layer1_outputs(3950) <= (layer0_outputs(4088)) and (layer0_outputs(3112));
    layer1_outputs(3951) <= not(layer0_outputs(51));
    layer1_outputs(3952) <= (layer0_outputs(3187)) and not (layer0_outputs(3755));
    layer1_outputs(3953) <= layer0_outputs(250);
    layer1_outputs(3954) <= layer0_outputs(3545);
    layer1_outputs(3955) <= not((layer0_outputs(1847)) and (layer0_outputs(3783)));
    layer1_outputs(3956) <= not(layer0_outputs(4023)) or (layer0_outputs(566));
    layer1_outputs(3957) <= not(layer0_outputs(283)) or (layer0_outputs(1522));
    layer1_outputs(3958) <= (layer0_outputs(4761)) and not (layer0_outputs(1391));
    layer1_outputs(3959) <= layer0_outputs(4338);
    layer1_outputs(3960) <= not(layer0_outputs(4102));
    layer1_outputs(3961) <= not(layer0_outputs(2679));
    layer1_outputs(3962) <= not((layer0_outputs(1182)) or (layer0_outputs(103)));
    layer1_outputs(3963) <= not((layer0_outputs(3842)) or (layer0_outputs(3659)));
    layer1_outputs(3964) <= not(layer0_outputs(3976)) or (layer0_outputs(1498));
    layer1_outputs(3965) <= (layer0_outputs(1088)) and (layer0_outputs(1841));
    layer1_outputs(3966) <= layer0_outputs(2897);
    layer1_outputs(3967) <= (layer0_outputs(2264)) and not (layer0_outputs(1683));
    layer1_outputs(3968) <= (layer0_outputs(3006)) and not (layer0_outputs(4886));
    layer1_outputs(3969) <= layer0_outputs(100);
    layer1_outputs(3970) <= (layer0_outputs(97)) and not (layer0_outputs(3325));
    layer1_outputs(3971) <= not(layer0_outputs(4773));
    layer1_outputs(3972) <= layer0_outputs(685);
    layer1_outputs(3973) <= (layer0_outputs(723)) and not (layer0_outputs(1452));
    layer1_outputs(3974) <= not((layer0_outputs(3103)) or (layer0_outputs(458)));
    layer1_outputs(3975) <= layer0_outputs(617);
    layer1_outputs(3976) <= (layer0_outputs(476)) or (layer0_outputs(1641));
    layer1_outputs(3977) <= not((layer0_outputs(1830)) xor (layer0_outputs(2684)));
    layer1_outputs(3978) <= not(layer0_outputs(2160));
    layer1_outputs(3979) <= (layer0_outputs(2674)) and (layer0_outputs(4414));
    layer1_outputs(3980) <= not(layer0_outputs(2645));
    layer1_outputs(3981) <= layer0_outputs(2710);
    layer1_outputs(3982) <= not(layer0_outputs(3759));
    layer1_outputs(3983) <= (layer0_outputs(948)) and not (layer0_outputs(4386));
    layer1_outputs(3984) <= not((layer0_outputs(3981)) xor (layer0_outputs(4099)));
    layer1_outputs(3985) <= not(layer0_outputs(3940));
    layer1_outputs(3986) <= not((layer0_outputs(2150)) or (layer0_outputs(2313)));
    layer1_outputs(3987) <= not(layer0_outputs(2245));
    layer1_outputs(3988) <= (layer0_outputs(4155)) and not (layer0_outputs(2069));
    layer1_outputs(3989) <= (layer0_outputs(2761)) xor (layer0_outputs(4649));
    layer1_outputs(3990) <= (layer0_outputs(2503)) xor (layer0_outputs(2211));
    layer1_outputs(3991) <= not(layer0_outputs(622));
    layer1_outputs(3992) <= (layer0_outputs(3320)) or (layer0_outputs(2171));
    layer1_outputs(3993) <= not((layer0_outputs(827)) xor (layer0_outputs(2017)));
    layer1_outputs(3994) <= not((layer0_outputs(1592)) xor (layer0_outputs(4593)));
    layer1_outputs(3995) <= (layer0_outputs(2275)) xor (layer0_outputs(4930));
    layer1_outputs(3996) <= not(layer0_outputs(1485)) or (layer0_outputs(3549));
    layer1_outputs(3997) <= '0';
    layer1_outputs(3998) <= not((layer0_outputs(2410)) and (layer0_outputs(4433)));
    layer1_outputs(3999) <= (layer0_outputs(1387)) and not (layer0_outputs(1466));
    layer1_outputs(4000) <= (layer0_outputs(2161)) and (layer0_outputs(1097));
    layer1_outputs(4001) <= (layer0_outputs(831)) xor (layer0_outputs(1186));
    layer1_outputs(4002) <= layer0_outputs(1484);
    layer1_outputs(4003) <= not((layer0_outputs(2005)) and (layer0_outputs(1125)));
    layer1_outputs(4004) <= (layer0_outputs(4546)) and not (layer0_outputs(374));
    layer1_outputs(4005) <= not(layer0_outputs(1074)) or (layer0_outputs(1564));
    layer1_outputs(4006) <= not((layer0_outputs(4877)) and (layer0_outputs(4461)));
    layer1_outputs(4007) <= not(layer0_outputs(205));
    layer1_outputs(4008) <= (layer0_outputs(1054)) xor (layer0_outputs(4550));
    layer1_outputs(4009) <= layer0_outputs(2073);
    layer1_outputs(4010) <= '1';
    layer1_outputs(4011) <= not(layer0_outputs(3719));
    layer1_outputs(4012) <= (layer0_outputs(338)) and not (layer0_outputs(4590));
    layer1_outputs(4013) <= not(layer0_outputs(1460));
    layer1_outputs(4014) <= not(layer0_outputs(1323));
    layer1_outputs(4015) <= not((layer0_outputs(609)) or (layer0_outputs(1291)));
    layer1_outputs(4016) <= '0';
    layer1_outputs(4017) <= (layer0_outputs(4799)) and not (layer0_outputs(127));
    layer1_outputs(4018) <= (layer0_outputs(708)) and (layer0_outputs(1643));
    layer1_outputs(4019) <= not((layer0_outputs(1246)) or (layer0_outputs(1743)));
    layer1_outputs(4020) <= (layer0_outputs(1867)) xor (layer0_outputs(333));
    layer1_outputs(4021) <= (layer0_outputs(456)) and not (layer0_outputs(696));
    layer1_outputs(4022) <= not((layer0_outputs(2968)) and (layer0_outputs(3226)));
    layer1_outputs(4023) <= not(layer0_outputs(4080)) or (layer0_outputs(3671));
    layer1_outputs(4024) <= not((layer0_outputs(1345)) or (layer0_outputs(817)));
    layer1_outputs(4025) <= not(layer0_outputs(3213)) or (layer0_outputs(1414));
    layer1_outputs(4026) <= layer0_outputs(2189);
    layer1_outputs(4027) <= not((layer0_outputs(901)) and (layer0_outputs(1795)));
    layer1_outputs(4028) <= layer0_outputs(3378);
    layer1_outputs(4029) <= not(layer0_outputs(2048)) or (layer0_outputs(4476));
    layer1_outputs(4030) <= not((layer0_outputs(1692)) and (layer0_outputs(2333)));
    layer1_outputs(4031) <= not((layer0_outputs(3059)) xor (layer0_outputs(1542)));
    layer1_outputs(4032) <= layer0_outputs(862);
    layer1_outputs(4033) <= not(layer0_outputs(4755));
    layer1_outputs(4034) <= '1';
    layer1_outputs(4035) <= (layer0_outputs(3369)) or (layer0_outputs(2516));
    layer1_outputs(4036) <= not(layer0_outputs(2525));
    layer1_outputs(4037) <= (layer0_outputs(1004)) and (layer0_outputs(4905));
    layer1_outputs(4038) <= not((layer0_outputs(3345)) and (layer0_outputs(4211)));
    layer1_outputs(4039) <= not(layer0_outputs(3313)) or (layer0_outputs(2106));
    layer1_outputs(4040) <= (layer0_outputs(2280)) or (layer0_outputs(2549));
    layer1_outputs(4041) <= not(layer0_outputs(828));
    layer1_outputs(4042) <= not(layer0_outputs(4390));
    layer1_outputs(4043) <= layer0_outputs(2362);
    layer1_outputs(4044) <= '0';
    layer1_outputs(4045) <= layer0_outputs(3439);
    layer1_outputs(4046) <= (layer0_outputs(177)) and (layer0_outputs(2578));
    layer1_outputs(4047) <= layer0_outputs(3919);
    layer1_outputs(4048) <= not((layer0_outputs(1577)) xor (layer0_outputs(2184)));
    layer1_outputs(4049) <= not(layer0_outputs(424)) or (layer0_outputs(2177));
    layer1_outputs(4050) <= layer0_outputs(1676);
    layer1_outputs(4051) <= (layer0_outputs(2956)) and not (layer0_outputs(565));
    layer1_outputs(4052) <= '0';
    layer1_outputs(4053) <= not(layer0_outputs(373)) or (layer0_outputs(838));
    layer1_outputs(4054) <= not(layer0_outputs(1183));
    layer1_outputs(4055) <= not(layer0_outputs(4423)) or (layer0_outputs(1929));
    layer1_outputs(4056) <= layer0_outputs(4037);
    layer1_outputs(4057) <= not(layer0_outputs(4464));
    layer1_outputs(4058) <= layer0_outputs(4519);
    layer1_outputs(4059) <= layer0_outputs(1611);
    layer1_outputs(4060) <= not((layer0_outputs(2371)) and (layer0_outputs(2814)));
    layer1_outputs(4061) <= (layer0_outputs(2243)) xor (layer0_outputs(72));
    layer1_outputs(4062) <= (layer0_outputs(1105)) and (layer0_outputs(2103));
    layer1_outputs(4063) <= not(layer0_outputs(847));
    layer1_outputs(4064) <= (layer0_outputs(3442)) or (layer0_outputs(1724));
    layer1_outputs(4065) <= (layer0_outputs(4722)) and not (layer0_outputs(4743));
    layer1_outputs(4066) <= (layer0_outputs(4030)) and not (layer0_outputs(2869));
    layer1_outputs(4067) <= (layer0_outputs(1243)) and not (layer0_outputs(2083));
    layer1_outputs(4068) <= not(layer0_outputs(5055));
    layer1_outputs(4069) <= (layer0_outputs(4250)) and not (layer0_outputs(3867));
    layer1_outputs(4070) <= not(layer0_outputs(346)) or (layer0_outputs(1170));
    layer1_outputs(4071) <= not((layer0_outputs(1309)) xor (layer0_outputs(700)));
    layer1_outputs(4072) <= (layer0_outputs(668)) and (layer0_outputs(2291));
    layer1_outputs(4073) <= not(layer0_outputs(1818));
    layer1_outputs(4074) <= (layer0_outputs(4839)) and not (layer0_outputs(743));
    layer1_outputs(4075) <= (layer0_outputs(5035)) and not (layer0_outputs(1518));
    layer1_outputs(4076) <= not(layer0_outputs(4609));
    layer1_outputs(4077) <= (layer0_outputs(2571)) and (layer0_outputs(188));
    layer1_outputs(4078) <= (layer0_outputs(3368)) and not (layer0_outputs(4283));
    layer1_outputs(4079) <= (layer0_outputs(1207)) and not (layer0_outputs(627));
    layer1_outputs(4080) <= (layer0_outputs(5)) and (layer0_outputs(4683));
    layer1_outputs(4081) <= (layer0_outputs(2982)) or (layer0_outputs(1609));
    layer1_outputs(4082) <= not(layer0_outputs(1565)) or (layer0_outputs(2965));
    layer1_outputs(4083) <= not((layer0_outputs(3899)) and (layer0_outputs(3343)));
    layer1_outputs(4084) <= not(layer0_outputs(2012)) or (layer0_outputs(1288));
    layer1_outputs(4085) <= not(layer0_outputs(2338)) or (layer0_outputs(3330));
    layer1_outputs(4086) <= not(layer0_outputs(775));
    layer1_outputs(4087) <= layer0_outputs(288);
    layer1_outputs(4088) <= not(layer0_outputs(1910));
    layer1_outputs(4089) <= (layer0_outputs(1736)) or (layer0_outputs(878));
    layer1_outputs(4090) <= not(layer0_outputs(2707));
    layer1_outputs(4091) <= (layer0_outputs(423)) and not (layer0_outputs(1803));
    layer1_outputs(4092) <= not((layer0_outputs(2791)) or (layer0_outputs(457)));
    layer1_outputs(4093) <= (layer0_outputs(4705)) xor (layer0_outputs(2782));
    layer1_outputs(4094) <= (layer0_outputs(402)) and not (layer0_outputs(3133));
    layer1_outputs(4095) <= layer0_outputs(893);
    layer1_outputs(4096) <= not(layer0_outputs(3139));
    layer1_outputs(4097) <= (layer0_outputs(3862)) and (layer0_outputs(644));
    layer1_outputs(4098) <= not(layer0_outputs(1404));
    layer1_outputs(4099) <= not(layer0_outputs(1750));
    layer1_outputs(4100) <= not(layer0_outputs(4078)) or (layer0_outputs(4547));
    layer1_outputs(4101) <= (layer0_outputs(3551)) and not (layer0_outputs(2214));
    layer1_outputs(4102) <= not(layer0_outputs(3349));
    layer1_outputs(4103) <= (layer0_outputs(2744)) and not (layer0_outputs(2742));
    layer1_outputs(4104) <= (layer0_outputs(4553)) and not (layer0_outputs(3635));
    layer1_outputs(4105) <= not((layer0_outputs(156)) and (layer0_outputs(4577)));
    layer1_outputs(4106) <= not(layer0_outputs(4797));
    layer1_outputs(4107) <= (layer0_outputs(5043)) and not (layer0_outputs(291));
    layer1_outputs(4108) <= not(layer0_outputs(1471));
    layer1_outputs(4109) <= not((layer0_outputs(4301)) or (layer0_outputs(4163)));
    layer1_outputs(4110) <= layer0_outputs(1231);
    layer1_outputs(4111) <= not(layer0_outputs(5059));
    layer1_outputs(4112) <= not((layer0_outputs(1915)) or (layer0_outputs(1908)));
    layer1_outputs(4113) <= not(layer0_outputs(4502));
    layer1_outputs(4114) <= (layer0_outputs(4058)) and not (layer0_outputs(1691));
    layer1_outputs(4115) <= not(layer0_outputs(1874));
    layer1_outputs(4116) <= (layer0_outputs(796)) and not (layer0_outputs(5095));
    layer1_outputs(4117) <= (layer0_outputs(2725)) and (layer0_outputs(546));
    layer1_outputs(4118) <= layer0_outputs(4209);
    layer1_outputs(4119) <= (layer0_outputs(2113)) and not (layer0_outputs(645));
    layer1_outputs(4120) <= not(layer0_outputs(2933));
    layer1_outputs(4121) <= not(layer0_outputs(5027));
    layer1_outputs(4122) <= not((layer0_outputs(3462)) and (layer0_outputs(2692)));
    layer1_outputs(4123) <= layer0_outputs(3379);
    layer1_outputs(4124) <= (layer0_outputs(2135)) and not (layer0_outputs(6));
    layer1_outputs(4125) <= (layer0_outputs(2463)) and (layer0_outputs(422));
    layer1_outputs(4126) <= not(layer0_outputs(388));
    layer1_outputs(4127) <= (layer0_outputs(1579)) or (layer0_outputs(883));
    layer1_outputs(4128) <= not((layer0_outputs(4494)) or (layer0_outputs(2561)));
    layer1_outputs(4129) <= layer0_outputs(596);
    layer1_outputs(4130) <= not(layer0_outputs(1106));
    layer1_outputs(4131) <= layer0_outputs(2713);
    layer1_outputs(4132) <= layer0_outputs(3389);
    layer1_outputs(4133) <= not((layer0_outputs(3416)) and (layer0_outputs(1103)));
    layer1_outputs(4134) <= layer0_outputs(1591);
    layer1_outputs(4135) <= (layer0_outputs(3727)) xor (layer0_outputs(1584));
    layer1_outputs(4136) <= (layer0_outputs(4115)) and (layer0_outputs(1368));
    layer1_outputs(4137) <= not(layer0_outputs(579)) or (layer0_outputs(3803));
    layer1_outputs(4138) <= (layer0_outputs(4109)) xor (layer0_outputs(3024));
    layer1_outputs(4139) <= layer0_outputs(481);
    layer1_outputs(4140) <= '0';
    layer1_outputs(4141) <= (layer0_outputs(2936)) and (layer0_outputs(2745));
    layer1_outputs(4142) <= not(layer0_outputs(1674)) or (layer0_outputs(551));
    layer1_outputs(4143) <= not(layer0_outputs(541)) or (layer0_outputs(4565));
    layer1_outputs(4144) <= (layer0_outputs(1633)) and (layer0_outputs(2904));
    layer1_outputs(4145) <= not((layer0_outputs(2591)) xor (layer0_outputs(4995)));
    layer1_outputs(4146) <= layer0_outputs(4470);
    layer1_outputs(4147) <= layer0_outputs(1501);
    layer1_outputs(4148) <= not(layer0_outputs(4869)) or (layer0_outputs(1451));
    layer1_outputs(4149) <= (layer0_outputs(2942)) or (layer0_outputs(3506));
    layer1_outputs(4150) <= layer0_outputs(4296);
    layer1_outputs(4151) <= not((layer0_outputs(2276)) or (layer0_outputs(2256)));
    layer1_outputs(4152) <= layer0_outputs(158);
    layer1_outputs(4153) <= (layer0_outputs(2610)) and (layer0_outputs(3717));
    layer1_outputs(4154) <= not(layer0_outputs(940));
    layer1_outputs(4155) <= not(layer0_outputs(4919));
    layer1_outputs(4156) <= not((layer0_outputs(3287)) xor (layer0_outputs(4484)));
    layer1_outputs(4157) <= not(layer0_outputs(1772));
    layer1_outputs(4158) <= layer0_outputs(3285);
    layer1_outputs(4159) <= (layer0_outputs(1730)) and not (layer0_outputs(3952));
    layer1_outputs(4160) <= not(layer0_outputs(3427)) or (layer0_outputs(238));
    layer1_outputs(4161) <= layer0_outputs(4797);
    layer1_outputs(4162) <= not(layer0_outputs(3161));
    layer1_outputs(4163) <= not((layer0_outputs(4139)) or (layer0_outputs(816)));
    layer1_outputs(4164) <= '0';
    layer1_outputs(4165) <= not((layer0_outputs(4857)) and (layer0_outputs(3383)));
    layer1_outputs(4166) <= not(layer0_outputs(4488));
    layer1_outputs(4167) <= (layer0_outputs(2617)) and (layer0_outputs(4209));
    layer1_outputs(4168) <= (layer0_outputs(530)) and not (layer0_outputs(2246));
    layer1_outputs(4169) <= not((layer0_outputs(2164)) or (layer0_outputs(2760)));
    layer1_outputs(4170) <= (layer0_outputs(1787)) and not (layer0_outputs(1249));
    layer1_outputs(4171) <= layer0_outputs(3828);
    layer1_outputs(4172) <= not(layer0_outputs(375));
    layer1_outputs(4173) <= (layer0_outputs(656)) and (layer0_outputs(4894));
    layer1_outputs(4174) <= (layer0_outputs(4597)) or (layer0_outputs(1120));
    layer1_outputs(4175) <= not(layer0_outputs(1606)) or (layer0_outputs(2041));
    layer1_outputs(4176) <= (layer0_outputs(3333)) and (layer0_outputs(4351));
    layer1_outputs(4177) <= layer0_outputs(1483);
    layer1_outputs(4178) <= not((layer0_outputs(3182)) or (layer0_outputs(3001)));
    layer1_outputs(4179) <= (layer0_outputs(703)) and not (layer0_outputs(2301));
    layer1_outputs(4180) <= layer0_outputs(1251);
    layer1_outputs(4181) <= layer0_outputs(4827);
    layer1_outputs(4182) <= not(layer0_outputs(1146)) or (layer0_outputs(3760));
    layer1_outputs(4183) <= (layer0_outputs(3044)) or (layer0_outputs(3037));
    layer1_outputs(4184) <= (layer0_outputs(1160)) and (layer0_outputs(850));
    layer1_outputs(4185) <= not((layer0_outputs(3817)) and (layer0_outputs(4469)));
    layer1_outputs(4186) <= (layer0_outputs(2388)) xor (layer0_outputs(4499));
    layer1_outputs(4187) <= not(layer0_outputs(3045));
    layer1_outputs(4188) <= layer0_outputs(2293);
    layer1_outputs(4189) <= not(layer0_outputs(2053)) or (layer0_outputs(931));
    layer1_outputs(4190) <= not(layer0_outputs(1830));
    layer1_outputs(4191) <= layer0_outputs(2675);
    layer1_outputs(4192) <= not((layer0_outputs(1711)) xor (layer0_outputs(2136)));
    layer1_outputs(4193) <= '1';
    layer1_outputs(4194) <= not(layer0_outputs(1211));
    layer1_outputs(4195) <= (layer0_outputs(4465)) and not (layer0_outputs(369));
    layer1_outputs(4196) <= not((layer0_outputs(4656)) or (layer0_outputs(2191)));
    layer1_outputs(4197) <= (layer0_outputs(952)) or (layer0_outputs(2922));
    layer1_outputs(4198) <= (layer0_outputs(724)) or (layer0_outputs(765));
    layer1_outputs(4199) <= (layer0_outputs(2363)) and not (layer0_outputs(3316));
    layer1_outputs(4200) <= not((layer0_outputs(1007)) or (layer0_outputs(761)));
    layer1_outputs(4201) <= not(layer0_outputs(744));
    layer1_outputs(4202) <= (layer0_outputs(4644)) xor (layer0_outputs(4789));
    layer1_outputs(4203) <= layer0_outputs(4562);
    layer1_outputs(4204) <= not((layer0_outputs(2875)) xor (layer0_outputs(589)));
    layer1_outputs(4205) <= (layer0_outputs(2892)) and not (layer0_outputs(3813));
    layer1_outputs(4206) <= '0';
    layer1_outputs(4207) <= not((layer0_outputs(2247)) and (layer0_outputs(4325)));
    layer1_outputs(4208) <= (layer0_outputs(2144)) and (layer0_outputs(2375));
    layer1_outputs(4209) <= (layer0_outputs(4766)) xor (layer0_outputs(984));
    layer1_outputs(4210) <= (layer0_outputs(4362)) or (layer0_outputs(2493));
    layer1_outputs(4211) <= layer0_outputs(187);
    layer1_outputs(4212) <= not(layer0_outputs(2621));
    layer1_outputs(4213) <= (layer0_outputs(5097)) and not (layer0_outputs(818));
    layer1_outputs(4214) <= not((layer0_outputs(4141)) and (layer0_outputs(1279)));
    layer1_outputs(4215) <= (layer0_outputs(4013)) or (layer0_outputs(1128));
    layer1_outputs(4216) <= not(layer0_outputs(159));
    layer1_outputs(4217) <= layer0_outputs(4822);
    layer1_outputs(4218) <= not(layer0_outputs(4962)) or (layer0_outputs(70));
    layer1_outputs(4219) <= not((layer0_outputs(3945)) and (layer0_outputs(1701)));
    layer1_outputs(4220) <= not(layer0_outputs(1446)) or (layer0_outputs(191));
    layer1_outputs(4221) <= '0';
    layer1_outputs(4222) <= (layer0_outputs(4569)) or (layer0_outputs(3124));
    layer1_outputs(4223) <= not(layer0_outputs(4124));
    layer1_outputs(4224) <= (layer0_outputs(3609)) and not (layer0_outputs(1435));
    layer1_outputs(4225) <= '1';
    layer1_outputs(4226) <= '1';
    layer1_outputs(4227) <= layer0_outputs(2790);
    layer1_outputs(4228) <= not(layer0_outputs(198)) or (layer0_outputs(4988));
    layer1_outputs(4229) <= not(layer0_outputs(4269));
    layer1_outputs(4230) <= not(layer0_outputs(468)) or (layer0_outputs(4769));
    layer1_outputs(4231) <= not((layer0_outputs(1470)) and (layer0_outputs(3870)));
    layer1_outputs(4232) <= layer0_outputs(1569);
    layer1_outputs(4233) <= not(layer0_outputs(4345)) or (layer0_outputs(1664));
    layer1_outputs(4234) <= not((layer0_outputs(852)) and (layer0_outputs(3532)));
    layer1_outputs(4235) <= '1';
    layer1_outputs(4236) <= not((layer0_outputs(943)) and (layer0_outputs(3835)));
    layer1_outputs(4237) <= (layer0_outputs(3975)) and (layer0_outputs(3575));
    layer1_outputs(4238) <= layer0_outputs(647);
    layer1_outputs(4239) <= not(layer0_outputs(2623)) or (layer0_outputs(4913));
    layer1_outputs(4240) <= not((layer0_outputs(2035)) and (layer0_outputs(2870)));
    layer1_outputs(4241) <= not((layer0_outputs(3048)) and (layer0_outputs(3868)));
    layer1_outputs(4242) <= not(layer0_outputs(767));
    layer1_outputs(4243) <= layer0_outputs(4148);
    layer1_outputs(4244) <= layer0_outputs(4699);
    layer1_outputs(4245) <= not((layer0_outputs(3592)) or (layer0_outputs(1450)));
    layer1_outputs(4246) <= not(layer0_outputs(1010)) or (layer0_outputs(561));
    layer1_outputs(4247) <= layer0_outputs(4788);
    layer1_outputs(4248) <= not(layer0_outputs(4521)) or (layer0_outputs(2769));
    layer1_outputs(4249) <= (layer0_outputs(4056)) and not (layer0_outputs(4296));
    layer1_outputs(4250) <= not(layer0_outputs(4013));
    layer1_outputs(4251) <= not((layer0_outputs(4881)) and (layer0_outputs(4219)));
    layer1_outputs(4252) <= not(layer0_outputs(2492)) or (layer0_outputs(4420));
    layer1_outputs(4253) <= not(layer0_outputs(2922));
    layer1_outputs(4254) <= (layer0_outputs(4626)) and not (layer0_outputs(3290));
    layer1_outputs(4255) <= not((layer0_outputs(2151)) and (layer0_outputs(2971)));
    layer1_outputs(4256) <= layer0_outputs(3891);
    layer1_outputs(4257) <= not(layer0_outputs(3278));
    layer1_outputs(4258) <= (layer0_outputs(4304)) and not (layer0_outputs(2153));
    layer1_outputs(4259) <= not(layer0_outputs(3796)) or (layer0_outputs(4705));
    layer1_outputs(4260) <= (layer0_outputs(552)) and (layer0_outputs(1726));
    layer1_outputs(4261) <= (layer0_outputs(657)) and not (layer0_outputs(892));
    layer1_outputs(4262) <= (layer0_outputs(2571)) and not (layer0_outputs(4884));
    layer1_outputs(4263) <= layer0_outputs(4406);
    layer1_outputs(4264) <= '1';
    layer1_outputs(4265) <= not(layer0_outputs(4454)) or (layer0_outputs(5039));
    layer1_outputs(4266) <= layer0_outputs(2491);
    layer1_outputs(4267) <= not(layer0_outputs(4523));
    layer1_outputs(4268) <= layer0_outputs(3224);
    layer1_outputs(4269) <= not((layer0_outputs(4520)) or (layer0_outputs(2845)));
    layer1_outputs(4270) <= (layer0_outputs(1220)) and not (layer0_outputs(2544));
    layer1_outputs(4271) <= not(layer0_outputs(1582));
    layer1_outputs(4272) <= (layer0_outputs(1521)) and (layer0_outputs(3783));
    layer1_outputs(4273) <= not(layer0_outputs(44)) or (layer0_outputs(2352));
    layer1_outputs(4274) <= (layer0_outputs(3609)) and not (layer0_outputs(2538));
    layer1_outputs(4275) <= not((layer0_outputs(1708)) and (layer0_outputs(145)));
    layer1_outputs(4276) <= layer0_outputs(1552);
    layer1_outputs(4277) <= not(layer0_outputs(2136)) or (layer0_outputs(3679));
    layer1_outputs(4278) <= layer0_outputs(1687);
    layer1_outputs(4279) <= not(layer0_outputs(1027)) or (layer0_outputs(1071));
    layer1_outputs(4280) <= not(layer0_outputs(757));
    layer1_outputs(4281) <= layer0_outputs(4875);
    layer1_outputs(4282) <= layer0_outputs(1118);
    layer1_outputs(4283) <= layer0_outputs(757);
    layer1_outputs(4284) <= not(layer0_outputs(4271)) or (layer0_outputs(3394));
    layer1_outputs(4285) <= not(layer0_outputs(1418));
    layer1_outputs(4286) <= not(layer0_outputs(1703));
    layer1_outputs(4287) <= not(layer0_outputs(1275)) or (layer0_outputs(2795));
    layer1_outputs(4288) <= (layer0_outputs(4654)) and (layer0_outputs(3863));
    layer1_outputs(4289) <= not(layer0_outputs(3697));
    layer1_outputs(4290) <= (layer0_outputs(447)) and not (layer0_outputs(290));
    layer1_outputs(4291) <= layer0_outputs(2464);
    layer1_outputs(4292) <= not(layer0_outputs(864));
    layer1_outputs(4293) <= not(layer0_outputs(853));
    layer1_outputs(4294) <= (layer0_outputs(4925)) or (layer0_outputs(4565));
    layer1_outputs(4295) <= layer0_outputs(2993);
    layer1_outputs(4296) <= layer0_outputs(2906);
    layer1_outputs(4297) <= (layer0_outputs(1408)) and not (layer0_outputs(184));
    layer1_outputs(4298) <= (layer0_outputs(326)) and not (layer0_outputs(398));
    layer1_outputs(4299) <= not((layer0_outputs(2665)) or (layer0_outputs(2199)));
    layer1_outputs(4300) <= (layer0_outputs(855)) and (layer0_outputs(110));
    layer1_outputs(4301) <= (layer0_outputs(1191)) and (layer0_outputs(1934));
    layer1_outputs(4302) <= layer0_outputs(5030);
    layer1_outputs(4303) <= layer0_outputs(1119);
    layer1_outputs(4304) <= not((layer0_outputs(2115)) and (layer0_outputs(1042)));
    layer1_outputs(4305) <= (layer0_outputs(3624)) and not (layer0_outputs(810));
    layer1_outputs(4306) <= not((layer0_outputs(4064)) xor (layer0_outputs(3528)));
    layer1_outputs(4307) <= not(layer0_outputs(2600)) or (layer0_outputs(1465));
    layer1_outputs(4308) <= '1';
    layer1_outputs(4309) <= (layer0_outputs(544)) and not (layer0_outputs(4973));
    layer1_outputs(4310) <= layer0_outputs(4492);
    layer1_outputs(4311) <= not(layer0_outputs(307));
    layer1_outputs(4312) <= (layer0_outputs(472)) and not (layer0_outputs(1737));
    layer1_outputs(4313) <= not((layer0_outputs(2349)) and (layer0_outputs(235)));
    layer1_outputs(4314) <= not(layer0_outputs(4762));
    layer1_outputs(4315) <= layer0_outputs(210);
    layer1_outputs(4316) <= (layer0_outputs(4403)) and (layer0_outputs(3898));
    layer1_outputs(4317) <= (layer0_outputs(1208)) and (layer0_outputs(3264));
    layer1_outputs(4318) <= (layer0_outputs(5009)) and (layer0_outputs(2154));
    layer1_outputs(4319) <= not((layer0_outputs(73)) xor (layer0_outputs(633)));
    layer1_outputs(4320) <= (layer0_outputs(3007)) and (layer0_outputs(1563));
    layer1_outputs(4321) <= not((layer0_outputs(2344)) and (layer0_outputs(1760)));
    layer1_outputs(4322) <= not(layer0_outputs(278)) or (layer0_outputs(3864));
    layer1_outputs(4323) <= not(layer0_outputs(2523));
    layer1_outputs(4324) <= layer0_outputs(1162);
    layer1_outputs(4325) <= layer0_outputs(118);
    layer1_outputs(4326) <= not(layer0_outputs(4375)) or (layer0_outputs(3962));
    layer1_outputs(4327) <= not(layer0_outputs(1162));
    layer1_outputs(4328) <= not((layer0_outputs(2954)) and (layer0_outputs(1843)));
    layer1_outputs(4329) <= not((layer0_outputs(264)) xor (layer0_outputs(953)));
    layer1_outputs(4330) <= '0';
    layer1_outputs(4331) <= layer0_outputs(2799);
    layer1_outputs(4332) <= not((layer0_outputs(3120)) or (layer0_outputs(1924)));
    layer1_outputs(4333) <= layer0_outputs(1495);
    layer1_outputs(4334) <= not((layer0_outputs(3187)) xor (layer0_outputs(1393)));
    layer1_outputs(4335) <= layer0_outputs(4086);
    layer1_outputs(4336) <= not(layer0_outputs(4294)) or (layer0_outputs(917));
    layer1_outputs(4337) <= not(layer0_outputs(693)) or (layer0_outputs(3592));
    layer1_outputs(4338) <= (layer0_outputs(1421)) xor (layer0_outputs(4214));
    layer1_outputs(4339) <= (layer0_outputs(564)) and not (layer0_outputs(379));
    layer1_outputs(4340) <= not((layer0_outputs(513)) xor (layer0_outputs(2866)));
    layer1_outputs(4341) <= (layer0_outputs(532)) and (layer0_outputs(4369));
    layer1_outputs(4342) <= not(layer0_outputs(733));
    layer1_outputs(4343) <= (layer0_outputs(1984)) and not (layer0_outputs(2486));
    layer1_outputs(4344) <= not(layer0_outputs(1438));
    layer1_outputs(4345) <= (layer0_outputs(2871)) and (layer0_outputs(2703));
    layer1_outputs(4346) <= (layer0_outputs(1732)) or (layer0_outputs(1824));
    layer1_outputs(4347) <= not(layer0_outputs(765));
    layer1_outputs(4348) <= layer0_outputs(2842);
    layer1_outputs(4349) <= (layer0_outputs(4781)) and (layer0_outputs(1147));
    layer1_outputs(4350) <= (layer0_outputs(1712)) and (layer0_outputs(2629));
    layer1_outputs(4351) <= not(layer0_outputs(3504));
    layer1_outputs(4352) <= not(layer0_outputs(4065)) or (layer0_outputs(1148));
    layer1_outputs(4353) <= not(layer0_outputs(4534)) or (layer0_outputs(913));
    layer1_outputs(4354) <= layer0_outputs(3924);
    layer1_outputs(4355) <= (layer0_outputs(3446)) xor (layer0_outputs(4627));
    layer1_outputs(4356) <= (layer0_outputs(4302)) xor (layer0_outputs(2645));
    layer1_outputs(4357) <= (layer0_outputs(292)) or (layer0_outputs(881));
    layer1_outputs(4358) <= layer0_outputs(4506);
    layer1_outputs(4359) <= not(layer0_outputs(5088)) or (layer0_outputs(2998));
    layer1_outputs(4360) <= (layer0_outputs(2693)) and not (layer0_outputs(3558));
    layer1_outputs(4361) <= (layer0_outputs(4815)) xor (layer0_outputs(92));
    layer1_outputs(4362) <= (layer0_outputs(3869)) and not (layer0_outputs(3294));
    layer1_outputs(4363) <= (layer0_outputs(3161)) and not (layer0_outputs(3899));
    layer1_outputs(4364) <= (layer0_outputs(3058)) xor (layer0_outputs(2247));
    layer1_outputs(4365) <= not(layer0_outputs(2923));
    layer1_outputs(4366) <= not(layer0_outputs(4575)) or (layer0_outputs(1950));
    layer1_outputs(4367) <= '1';
    layer1_outputs(4368) <= (layer0_outputs(4426)) and (layer0_outputs(4305));
    layer1_outputs(4369) <= layer0_outputs(1739);
    layer1_outputs(4370) <= (layer0_outputs(3158)) and not (layer0_outputs(2689));
    layer1_outputs(4371) <= layer0_outputs(5079);
    layer1_outputs(4372) <= not((layer0_outputs(1995)) xor (layer0_outputs(3620)));
    layer1_outputs(4373) <= '0';
    layer1_outputs(4374) <= not((layer0_outputs(1433)) xor (layer0_outputs(853)));
    layer1_outputs(4375) <= (layer0_outputs(785)) and not (layer0_outputs(538));
    layer1_outputs(4376) <= not(layer0_outputs(3074));
    layer1_outputs(4377) <= not(layer0_outputs(2758)) or (layer0_outputs(1151));
    layer1_outputs(4378) <= layer0_outputs(1962);
    layer1_outputs(4379) <= not((layer0_outputs(2475)) and (layer0_outputs(1328)));
    layer1_outputs(4380) <= (layer0_outputs(4616)) and (layer0_outputs(1447));
    layer1_outputs(4381) <= (layer0_outputs(2501)) and (layer0_outputs(318));
    layer1_outputs(4382) <= not(layer0_outputs(1686)) or (layer0_outputs(1518));
    layer1_outputs(4383) <= not((layer0_outputs(2809)) or (layer0_outputs(4852)));
    layer1_outputs(4384) <= not(layer0_outputs(3062)) or (layer0_outputs(3312));
    layer1_outputs(4385) <= '1';
    layer1_outputs(4386) <= (layer0_outputs(90)) xor (layer0_outputs(4162));
    layer1_outputs(4387) <= not(layer0_outputs(3925));
    layer1_outputs(4388) <= not((layer0_outputs(1788)) and (layer0_outputs(4835)));
    layer1_outputs(4389) <= (layer0_outputs(4129)) xor (layer0_outputs(3075));
    layer1_outputs(4390) <= '1';
    layer1_outputs(4391) <= (layer0_outputs(1383)) and not (layer0_outputs(98));
    layer1_outputs(4392) <= layer0_outputs(3828);
    layer1_outputs(4393) <= (layer0_outputs(1392)) and not (layer0_outputs(2577));
    layer1_outputs(4394) <= not(layer0_outputs(1402)) or (layer0_outputs(3961));
    layer1_outputs(4395) <= (layer0_outputs(1719)) or (layer0_outputs(3045));
    layer1_outputs(4396) <= (layer0_outputs(406)) and not (layer0_outputs(968));
    layer1_outputs(4397) <= (layer0_outputs(2066)) and not (layer0_outputs(4643));
    layer1_outputs(4398) <= not((layer0_outputs(1526)) or (layer0_outputs(1649)));
    layer1_outputs(4399) <= not(layer0_outputs(47)) or (layer0_outputs(1846));
    layer1_outputs(4400) <= not((layer0_outputs(4594)) and (layer0_outputs(3009)));
    layer1_outputs(4401) <= not(layer0_outputs(2423));
    layer1_outputs(4402) <= not((layer0_outputs(1657)) xor (layer0_outputs(2232)));
    layer1_outputs(4403) <= (layer0_outputs(2208)) and (layer0_outputs(3985));
    layer1_outputs(4404) <= (layer0_outputs(221)) xor (layer0_outputs(7));
    layer1_outputs(4405) <= (layer0_outputs(4711)) and not (layer0_outputs(2972));
    layer1_outputs(4406) <= (layer0_outputs(4737)) and (layer0_outputs(1407));
    layer1_outputs(4407) <= (layer0_outputs(4838)) or (layer0_outputs(380));
    layer1_outputs(4408) <= not(layer0_outputs(3928));
    layer1_outputs(4409) <= layer0_outputs(3175);
    layer1_outputs(4410) <= not(layer0_outputs(43));
    layer1_outputs(4411) <= layer0_outputs(1571);
    layer1_outputs(4412) <= (layer0_outputs(1666)) and not (layer0_outputs(958));
    layer1_outputs(4413) <= not(layer0_outputs(4108));
    layer1_outputs(4414) <= layer0_outputs(650);
    layer1_outputs(4415) <= (layer0_outputs(3276)) xor (layer0_outputs(1442));
    layer1_outputs(4416) <= (layer0_outputs(1791)) and not (layer0_outputs(3191));
    layer1_outputs(4417) <= (layer0_outputs(946)) or (layer0_outputs(2278));
    layer1_outputs(4418) <= not(layer0_outputs(4294)) or (layer0_outputs(166));
    layer1_outputs(4419) <= (layer0_outputs(4818)) or (layer0_outputs(1991));
    layer1_outputs(4420) <= (layer0_outputs(2367)) xor (layer0_outputs(4802));
    layer1_outputs(4421) <= (layer0_outputs(2034)) and (layer0_outputs(3980));
    layer1_outputs(4422) <= not((layer0_outputs(4996)) and (layer0_outputs(4817)));
    layer1_outputs(4423) <= layer0_outputs(95);
    layer1_outputs(4424) <= (layer0_outputs(300)) xor (layer0_outputs(2138));
    layer1_outputs(4425) <= layer0_outputs(3804);
    layer1_outputs(4426) <= (layer0_outputs(3378)) and not (layer0_outputs(3991));
    layer1_outputs(4427) <= not(layer0_outputs(32));
    layer1_outputs(4428) <= (layer0_outputs(4522)) and not (layer0_outputs(1325));
    layer1_outputs(4429) <= not(layer0_outputs(1128)) or (layer0_outputs(4865));
    layer1_outputs(4430) <= not(layer0_outputs(4099));
    layer1_outputs(4431) <= not((layer0_outputs(1432)) and (layer0_outputs(4377)));
    layer1_outputs(4432) <= not(layer0_outputs(1370));
    layer1_outputs(4433) <= not(layer0_outputs(4965)) or (layer0_outputs(2279));
    layer1_outputs(4434) <= layer0_outputs(1216);
    layer1_outputs(4435) <= (layer0_outputs(1851)) and not (layer0_outputs(3730));
    layer1_outputs(4436) <= not(layer0_outputs(4380));
    layer1_outputs(4437) <= not(layer0_outputs(242));
    layer1_outputs(4438) <= not(layer0_outputs(4471));
    layer1_outputs(4439) <= (layer0_outputs(4021)) or (layer0_outputs(1060));
    layer1_outputs(4440) <= layer0_outputs(1058);
    layer1_outputs(4441) <= (layer0_outputs(4346)) and (layer0_outputs(3115));
    layer1_outputs(4442) <= (layer0_outputs(623)) and (layer0_outputs(294));
    layer1_outputs(4443) <= '1';
    layer1_outputs(4444) <= not(layer0_outputs(267)) or (layer0_outputs(1975));
    layer1_outputs(4445) <= not(layer0_outputs(1807)) or (layer0_outputs(2228));
    layer1_outputs(4446) <= not(layer0_outputs(656)) or (layer0_outputs(3154));
    layer1_outputs(4447) <= not(layer0_outputs(3529)) or (layer0_outputs(924));
    layer1_outputs(4448) <= not(layer0_outputs(1940));
    layer1_outputs(4449) <= (layer0_outputs(4418)) and not (layer0_outputs(892));
    layer1_outputs(4450) <= not(layer0_outputs(713));
    layer1_outputs(4451) <= not(layer0_outputs(4069));
    layer1_outputs(4452) <= not(layer0_outputs(24)) or (layer0_outputs(3445));
    layer1_outputs(4453) <= layer0_outputs(13);
    layer1_outputs(4454) <= (layer0_outputs(5098)) and (layer0_outputs(2132));
    layer1_outputs(4455) <= not(layer0_outputs(1996));
    layer1_outputs(4456) <= not((layer0_outputs(3775)) and (layer0_outputs(5081)));
    layer1_outputs(4457) <= (layer0_outputs(320)) and not (layer0_outputs(4903));
    layer1_outputs(4458) <= not(layer0_outputs(1909));
    layer1_outputs(4459) <= layer0_outputs(4781);
    layer1_outputs(4460) <= '1';
    layer1_outputs(4461) <= not(layer0_outputs(3156)) or (layer0_outputs(4228));
    layer1_outputs(4462) <= layer0_outputs(1882);
    layer1_outputs(4463) <= not(layer0_outputs(1651));
    layer1_outputs(4464) <= (layer0_outputs(4800)) and not (layer0_outputs(467));
    layer1_outputs(4465) <= (layer0_outputs(3309)) and not (layer0_outputs(384));
    layer1_outputs(4466) <= layer0_outputs(4134);
    layer1_outputs(4467) <= layer0_outputs(4673);
    layer1_outputs(4468) <= layer0_outputs(2654);
    layer1_outputs(4469) <= not((layer0_outputs(4428)) or (layer0_outputs(679)));
    layer1_outputs(4470) <= (layer0_outputs(2901)) or (layer0_outputs(1424));
    layer1_outputs(4471) <= not(layer0_outputs(2449));
    layer1_outputs(4472) <= (layer0_outputs(650)) xor (layer0_outputs(4225));
    layer1_outputs(4473) <= not(layer0_outputs(3113));
    layer1_outputs(4474) <= (layer0_outputs(3093)) and not (layer0_outputs(790));
    layer1_outputs(4475) <= (layer0_outputs(526)) xor (layer0_outputs(3425));
    layer1_outputs(4476) <= layer0_outputs(1929);
    layer1_outputs(4477) <= '1';
    layer1_outputs(4478) <= '1';
    layer1_outputs(4479) <= layer0_outputs(1110);
    layer1_outputs(4480) <= (layer0_outputs(3695)) and not (layer0_outputs(619));
    layer1_outputs(4481) <= not(layer0_outputs(1324));
    layer1_outputs(4482) <= '0';
    layer1_outputs(4483) <= (layer0_outputs(1325)) and not (layer0_outputs(387));
    layer1_outputs(4484) <= layer0_outputs(2116);
    layer1_outputs(4485) <= not(layer0_outputs(4370));
    layer1_outputs(4486) <= not((layer0_outputs(460)) and (layer0_outputs(2366)));
    layer1_outputs(4487) <= not(layer0_outputs(3277)) or (layer0_outputs(1297));
    layer1_outputs(4488) <= not(layer0_outputs(3689));
    layer1_outputs(4489) <= not(layer0_outputs(2798));
    layer1_outputs(4490) <= not(layer0_outputs(5079));
    layer1_outputs(4491) <= (layer0_outputs(2945)) and not (layer0_outputs(3598));
    layer1_outputs(4492) <= '0';
    layer1_outputs(4493) <= not(layer0_outputs(1481)) or (layer0_outputs(4759));
    layer1_outputs(4494) <= (layer0_outputs(680)) and (layer0_outputs(1019));
    layer1_outputs(4495) <= (layer0_outputs(631)) and (layer0_outputs(3229));
    layer1_outputs(4496) <= layer0_outputs(2856);
    layer1_outputs(4497) <= (layer0_outputs(1283)) and not (layer0_outputs(4164));
    layer1_outputs(4498) <= not(layer0_outputs(3207));
    layer1_outputs(4499) <= not(layer0_outputs(3189)) or (layer0_outputs(3733));
    layer1_outputs(4500) <= (layer0_outputs(124)) or (layer0_outputs(1171));
    layer1_outputs(4501) <= not((layer0_outputs(1030)) xor (layer0_outputs(1064)));
    layer1_outputs(4502) <= (layer0_outputs(1728)) or (layer0_outputs(2761));
    layer1_outputs(4503) <= not(layer0_outputs(1839)) or (layer0_outputs(862));
    layer1_outputs(4504) <= layer0_outputs(4335);
    layer1_outputs(4505) <= (layer0_outputs(3701)) and (layer0_outputs(3248));
    layer1_outputs(4506) <= (layer0_outputs(3708)) and not (layer0_outputs(4140));
    layer1_outputs(4507) <= layer0_outputs(1882);
    layer1_outputs(4508) <= not((layer0_outputs(133)) xor (layer0_outputs(4622)));
    layer1_outputs(4509) <= (layer0_outputs(2575)) or (layer0_outputs(1256));
    layer1_outputs(4510) <= not(layer0_outputs(4129));
    layer1_outputs(4511) <= not(layer0_outputs(80)) or (layer0_outputs(3345));
    layer1_outputs(4512) <= not(layer0_outputs(3639));
    layer1_outputs(4513) <= not(layer0_outputs(3190));
    layer1_outputs(4514) <= (layer0_outputs(3994)) and (layer0_outputs(571));
    layer1_outputs(4515) <= not((layer0_outputs(4325)) and (layer0_outputs(3400)));
    layer1_outputs(4516) <= not(layer0_outputs(2653));
    layer1_outputs(4517) <= not((layer0_outputs(2721)) and (layer0_outputs(1566)));
    layer1_outputs(4518) <= '0';
    layer1_outputs(4519) <= not(layer0_outputs(3975));
    layer1_outputs(4520) <= not((layer0_outputs(2957)) or (layer0_outputs(4740)));
    layer1_outputs(4521) <= (layer0_outputs(4898)) and not (layer0_outputs(2171));
    layer1_outputs(4522) <= not(layer0_outputs(3557));
    layer1_outputs(4523) <= not(layer0_outputs(2548)) or (layer0_outputs(2898));
    layer1_outputs(4524) <= (layer0_outputs(1881)) or (layer0_outputs(2056));
    layer1_outputs(4525) <= layer0_outputs(4293);
    layer1_outputs(4526) <= (layer0_outputs(852)) and not (layer0_outputs(889));
    layer1_outputs(4527) <= not((layer0_outputs(1170)) or (layer0_outputs(4735)));
    layer1_outputs(4528) <= not(layer0_outputs(1842));
    layer1_outputs(4529) <= layer0_outputs(4240);
    layer1_outputs(4530) <= '0';
    layer1_outputs(4531) <= layer0_outputs(2088);
    layer1_outputs(4532) <= (layer0_outputs(3261)) and (layer0_outputs(3244));
    layer1_outputs(4533) <= not(layer0_outputs(2062)) or (layer0_outputs(735));
    layer1_outputs(4534) <= not((layer0_outputs(4101)) and (layer0_outputs(253)));
    layer1_outputs(4535) <= '1';
    layer1_outputs(4536) <= (layer0_outputs(2948)) and not (layer0_outputs(417));
    layer1_outputs(4537) <= not(layer0_outputs(4841));
    layer1_outputs(4538) <= '1';
    layer1_outputs(4539) <= layer0_outputs(1622);
    layer1_outputs(4540) <= (layer0_outputs(2203)) and (layer0_outputs(603));
    layer1_outputs(4541) <= not(layer0_outputs(5051)) or (layer0_outputs(4844));
    layer1_outputs(4542) <= not((layer0_outputs(1727)) and (layer0_outputs(4858)));
    layer1_outputs(4543) <= not(layer0_outputs(1377));
    layer1_outputs(4544) <= (layer0_outputs(1340)) or (layer0_outputs(1006));
    layer1_outputs(4545) <= not((layer0_outputs(1257)) or (layer0_outputs(3142)));
    layer1_outputs(4546) <= (layer0_outputs(1017)) and not (layer0_outputs(14));
    layer1_outputs(4547) <= not(layer0_outputs(3223));
    layer1_outputs(4548) <= not(layer0_outputs(261)) or (layer0_outputs(3615));
    layer1_outputs(4549) <= (layer0_outputs(1342)) or (layer0_outputs(1585));
    layer1_outputs(4550) <= not(layer0_outputs(2649));
    layer1_outputs(4551) <= not((layer0_outputs(2910)) or (layer0_outputs(3540)));
    layer1_outputs(4552) <= not(layer0_outputs(1992)) or (layer0_outputs(2637));
    layer1_outputs(4553) <= (layer0_outputs(3988)) and (layer0_outputs(2255));
    layer1_outputs(4554) <= not((layer0_outputs(2413)) and (layer0_outputs(4231)));
    layer1_outputs(4555) <= not(layer0_outputs(2100)) or (layer0_outputs(4392));
    layer1_outputs(4556) <= (layer0_outputs(4521)) and not (layer0_outputs(4133));
    layer1_outputs(4557) <= (layer0_outputs(2749)) and not (layer0_outputs(2015));
    layer1_outputs(4558) <= layer0_outputs(4912);
    layer1_outputs(4559) <= not((layer0_outputs(3463)) or (layer0_outputs(1244)));
    layer1_outputs(4560) <= (layer0_outputs(4385)) and not (layer0_outputs(4121));
    layer1_outputs(4561) <= not(layer0_outputs(3146));
    layer1_outputs(4562) <= not(layer0_outputs(2325)) or (layer0_outputs(2131));
    layer1_outputs(4563) <= (layer0_outputs(199)) and (layer0_outputs(152));
    layer1_outputs(4564) <= not((layer0_outputs(1144)) xor (layer0_outputs(7)));
    layer1_outputs(4565) <= not(layer0_outputs(2055));
    layer1_outputs(4566) <= '1';
    layer1_outputs(4567) <= not(layer0_outputs(3225));
    layer1_outputs(4568) <= not(layer0_outputs(1576)) or (layer0_outputs(1106));
    layer1_outputs(4569) <= not(layer0_outputs(1942));
    layer1_outputs(4570) <= (layer0_outputs(289)) xor (layer0_outputs(2325));
    layer1_outputs(4571) <= not(layer0_outputs(149));
    layer1_outputs(4572) <= (layer0_outputs(616)) and (layer0_outputs(2951));
    layer1_outputs(4573) <= '1';
    layer1_outputs(4574) <= (layer0_outputs(1837)) and not (layer0_outputs(1812));
    layer1_outputs(4575) <= not(layer0_outputs(1663));
    layer1_outputs(4576) <= not((layer0_outputs(3865)) xor (layer0_outputs(2180)));
    layer1_outputs(4577) <= layer0_outputs(4975);
    layer1_outputs(4578) <= not(layer0_outputs(3652)) or (layer0_outputs(2079));
    layer1_outputs(4579) <= not(layer0_outputs(3214)) or (layer0_outputs(2074));
    layer1_outputs(4580) <= not((layer0_outputs(431)) and (layer0_outputs(4035)));
    layer1_outputs(4581) <= (layer0_outputs(4493)) or (layer0_outputs(4450));
    layer1_outputs(4582) <= not(layer0_outputs(1987));
    layer1_outputs(4583) <= (layer0_outputs(1500)) xor (layer0_outputs(2483));
    layer1_outputs(4584) <= (layer0_outputs(3636)) and not (layer0_outputs(3037));
    layer1_outputs(4585) <= not((layer0_outputs(4658)) and (layer0_outputs(9)));
    layer1_outputs(4586) <= not((layer0_outputs(2616)) or (layer0_outputs(159)));
    layer1_outputs(4587) <= (layer0_outputs(2282)) or (layer0_outputs(3081));
    layer1_outputs(4588) <= not(layer0_outputs(4868));
    layer1_outputs(4589) <= not(layer0_outputs(2589)) or (layer0_outputs(1083));
    layer1_outputs(4590) <= not((layer0_outputs(3366)) or (layer0_outputs(3829)));
    layer1_outputs(4591) <= not((layer0_outputs(1608)) or (layer0_outputs(1502)));
    layer1_outputs(4592) <= layer0_outputs(3847);
    layer1_outputs(4593) <= (layer0_outputs(1740)) xor (layer0_outputs(1854));
    layer1_outputs(4594) <= not((layer0_outputs(4545)) or (layer0_outputs(3302)));
    layer1_outputs(4595) <= layer0_outputs(3057);
    layer1_outputs(4596) <= (layer0_outputs(157)) and not (layer0_outputs(25));
    layer1_outputs(4597) <= not(layer0_outputs(474)) or (layer0_outputs(1272));
    layer1_outputs(4598) <= layer0_outputs(2272);
    layer1_outputs(4599) <= not(layer0_outputs(3825));
    layer1_outputs(4600) <= '0';
    layer1_outputs(4601) <= not(layer0_outputs(1362)) or (layer0_outputs(1700));
    layer1_outputs(4602) <= not((layer0_outputs(2596)) xor (layer0_outputs(3629)));
    layer1_outputs(4603) <= not((layer0_outputs(4381)) and (layer0_outputs(348)));
    layer1_outputs(4604) <= not(layer0_outputs(4741)) or (layer0_outputs(3100));
    layer1_outputs(4605) <= not(layer0_outputs(4232)) or (layer0_outputs(2632));
    layer1_outputs(4606) <= not((layer0_outputs(1805)) or (layer0_outputs(2306)));
    layer1_outputs(4607) <= not((layer0_outputs(4438)) or (layer0_outputs(790)));
    layer1_outputs(4608) <= not((layer0_outputs(1527)) or (layer0_outputs(4425)));
    layer1_outputs(4609) <= not(layer0_outputs(4215)) or (layer0_outputs(4634));
    layer1_outputs(4610) <= not(layer0_outputs(873));
    layer1_outputs(4611) <= (layer0_outputs(4236)) and not (layer0_outputs(2490));
    layer1_outputs(4612) <= not(layer0_outputs(2622));
    layer1_outputs(4613) <= not((layer0_outputs(536)) and (layer0_outputs(3675)));
    layer1_outputs(4614) <= not(layer0_outputs(1794)) or (layer0_outputs(5100));
    layer1_outputs(4615) <= not((layer0_outputs(4317)) or (layer0_outputs(1141)));
    layer1_outputs(4616) <= layer0_outputs(4153);
    layer1_outputs(4617) <= not(layer0_outputs(4721)) or (layer0_outputs(358));
    layer1_outputs(4618) <= (layer0_outputs(1632)) xor (layer0_outputs(2286));
    layer1_outputs(4619) <= '0';
    layer1_outputs(4620) <= layer0_outputs(2598);
    layer1_outputs(4621) <= not(layer0_outputs(1357));
    layer1_outputs(4622) <= (layer0_outputs(3939)) and not (layer0_outputs(2134));
    layer1_outputs(4623) <= not((layer0_outputs(3055)) or (layer0_outputs(4)));
    layer1_outputs(4624) <= not((layer0_outputs(727)) or (layer0_outputs(3036)));
    layer1_outputs(4625) <= not((layer0_outputs(1318)) or (layer0_outputs(2219)));
    layer1_outputs(4626) <= (layer0_outputs(5056)) xor (layer0_outputs(844));
    layer1_outputs(4627) <= layer0_outputs(1193);
    layer1_outputs(4628) <= not((layer0_outputs(2043)) or (layer0_outputs(1561)));
    layer1_outputs(4629) <= not((layer0_outputs(4261)) and (layer0_outputs(4136)));
    layer1_outputs(4630) <= not(layer0_outputs(4978));
    layer1_outputs(4631) <= not(layer0_outputs(4710));
    layer1_outputs(4632) <= not(layer0_outputs(160));
    layer1_outputs(4633) <= not(layer0_outputs(4739));
    layer1_outputs(4634) <= not(layer0_outputs(4119)) or (layer0_outputs(4159));
    layer1_outputs(4635) <= not((layer0_outputs(10)) xor (layer0_outputs(922)));
    layer1_outputs(4636) <= not(layer0_outputs(234));
    layer1_outputs(4637) <= not(layer0_outputs(1313));
    layer1_outputs(4638) <= not(layer0_outputs(3331)) or (layer0_outputs(3605));
    layer1_outputs(4639) <= '0';
    layer1_outputs(4640) <= not((layer0_outputs(3135)) or (layer0_outputs(4720)));
    layer1_outputs(4641) <= not(layer0_outputs(5)) or (layer0_outputs(4063));
    layer1_outputs(4642) <= not(layer0_outputs(4805)) or (layer0_outputs(568));
    layer1_outputs(4643) <= layer0_outputs(2109);
    layer1_outputs(4644) <= (layer0_outputs(3514)) and not (layer0_outputs(4895));
    layer1_outputs(4645) <= not(layer0_outputs(2680));
    layer1_outputs(4646) <= not(layer0_outputs(2702));
    layer1_outputs(4647) <= not(layer0_outputs(3221));
    layer1_outputs(4648) <= not(layer0_outputs(816));
    layer1_outputs(4649) <= not(layer0_outputs(2251));
    layer1_outputs(4650) <= not(layer0_outputs(2476));
    layer1_outputs(4651) <= not((layer0_outputs(3311)) xor (layer0_outputs(1848)));
    layer1_outputs(4652) <= not(layer0_outputs(3955)) or (layer0_outputs(1059));
    layer1_outputs(4653) <= not(layer0_outputs(2673)) or (layer0_outputs(4464));
    layer1_outputs(4654) <= not(layer0_outputs(67));
    layer1_outputs(4655) <= (layer0_outputs(254)) and not (layer0_outputs(4558));
    layer1_outputs(4656) <= not(layer0_outputs(2072)) or (layer0_outputs(1748));
    layer1_outputs(4657) <= (layer0_outputs(1631)) and not (layer0_outputs(4184));
    layer1_outputs(4658) <= not((layer0_outputs(947)) or (layer0_outputs(2669)));
    layer1_outputs(4659) <= (layer0_outputs(4525)) and not (layer0_outputs(343));
    layer1_outputs(4660) <= (layer0_outputs(2751)) xor (layer0_outputs(3141));
    layer1_outputs(4661) <= (layer0_outputs(2618)) or (layer0_outputs(4732));
    layer1_outputs(4662) <= layer0_outputs(1287);
    layer1_outputs(4663) <= layer0_outputs(4419);
    layer1_outputs(4664) <= not((layer0_outputs(1180)) or (layer0_outputs(4468)));
    layer1_outputs(4665) <= not(layer0_outputs(324)) or (layer0_outputs(920));
    layer1_outputs(4666) <= layer0_outputs(2229);
    layer1_outputs(4667) <= not(layer0_outputs(845)) or (layer0_outputs(3610));
    layer1_outputs(4668) <= (layer0_outputs(3256)) or (layer0_outputs(3509));
    layer1_outputs(4669) <= layer0_outputs(2729);
    layer1_outputs(4670) <= not(layer0_outputs(693)) or (layer0_outputs(2323));
    layer1_outputs(4671) <= layer0_outputs(5053);
    layer1_outputs(4672) <= not(layer0_outputs(1348));
    layer1_outputs(4673) <= '1';
    layer1_outputs(4674) <= not(layer0_outputs(2676));
    layer1_outputs(4675) <= layer0_outputs(684);
    layer1_outputs(4676) <= not(layer0_outputs(2984));
    layer1_outputs(4677) <= not(layer0_outputs(4507));
    layer1_outputs(4678) <= (layer0_outputs(1666)) and not (layer0_outputs(1654));
    layer1_outputs(4679) <= not(layer0_outputs(1697));
    layer1_outputs(4680) <= not(layer0_outputs(2404));
    layer1_outputs(4681) <= not(layer0_outputs(1376)) or (layer0_outputs(1745));
    layer1_outputs(4682) <= layer0_outputs(3332);
    layer1_outputs(4683) <= not((layer0_outputs(4446)) or (layer0_outputs(989)));
    layer1_outputs(4684) <= (layer0_outputs(3217)) and (layer0_outputs(4302));
    layer1_outputs(4685) <= not((layer0_outputs(4809)) or (layer0_outputs(3930)));
    layer1_outputs(4686) <= not((layer0_outputs(1961)) xor (layer0_outputs(4457)));
    layer1_outputs(4687) <= not(layer0_outputs(2537));
    layer1_outputs(4688) <= (layer0_outputs(1613)) and (layer0_outputs(2399));
    layer1_outputs(4689) <= not(layer0_outputs(1270)) or (layer0_outputs(3541));
    layer1_outputs(4690) <= not(layer0_outputs(2423));
    layer1_outputs(4691) <= not((layer0_outputs(1412)) xor (layer0_outputs(669)));
    layer1_outputs(4692) <= layer0_outputs(2949);
    layer1_outputs(4693) <= layer0_outputs(3396);
    layer1_outputs(4694) <= (layer0_outputs(3080)) and not (layer0_outputs(906));
    layer1_outputs(4695) <= not(layer0_outputs(1576));
    layer1_outputs(4696) <= (layer0_outputs(1026)) and not (layer0_outputs(393));
    layer1_outputs(4697) <= layer0_outputs(4351);
    layer1_outputs(4698) <= (layer0_outputs(2233)) xor (layer0_outputs(1165));
    layer1_outputs(4699) <= layer0_outputs(1874);
    layer1_outputs(4700) <= (layer0_outputs(3643)) and not (layer0_outputs(458));
    layer1_outputs(4701) <= not((layer0_outputs(4583)) and (layer0_outputs(2409)));
    layer1_outputs(4702) <= not((layer0_outputs(1282)) or (layer0_outputs(1284)));
    layer1_outputs(4703) <= layer0_outputs(3551);
    layer1_outputs(4704) <= '0';
    layer1_outputs(4705) <= '0';
    layer1_outputs(4706) <= not((layer0_outputs(0)) xor (layer0_outputs(4939)));
    layer1_outputs(4707) <= layer0_outputs(2916);
    layer1_outputs(4708) <= (layer0_outputs(1310)) or (layer0_outputs(4780));
    layer1_outputs(4709) <= not((layer0_outputs(21)) and (layer0_outputs(105)));
    layer1_outputs(4710) <= (layer0_outputs(4289)) xor (layer0_outputs(1243));
    layer1_outputs(4711) <= (layer0_outputs(1571)) or (layer0_outputs(3264));
    layer1_outputs(4712) <= layer0_outputs(2217);
    layer1_outputs(4713) <= not(layer0_outputs(2201));
    layer1_outputs(4714) <= not((layer0_outputs(70)) xor (layer0_outputs(3364)));
    layer1_outputs(4715) <= layer0_outputs(4868);
    layer1_outputs(4716) <= not(layer0_outputs(4183));
    layer1_outputs(4717) <= not((layer0_outputs(770)) and (layer0_outputs(4233)));
    layer1_outputs(4718) <= not((layer0_outputs(3920)) or (layer0_outputs(4388)));
    layer1_outputs(4719) <= not(layer0_outputs(2232));
    layer1_outputs(4720) <= (layer0_outputs(109)) and not (layer0_outputs(4157));
    layer1_outputs(4721) <= (layer0_outputs(2703)) and (layer0_outputs(265));
    layer1_outputs(4722) <= not(layer0_outputs(3654));
    layer1_outputs(4723) <= not(layer0_outputs(4081));
    layer1_outputs(4724) <= not(layer0_outputs(88));
    layer1_outputs(4725) <= not(layer0_outputs(1220));
    layer1_outputs(4726) <= not(layer0_outputs(3430));
    layer1_outputs(4727) <= layer0_outputs(4745);
    layer1_outputs(4728) <= (layer0_outputs(4833)) and not (layer0_outputs(5009));
    layer1_outputs(4729) <= not(layer0_outputs(3566));
    layer1_outputs(4730) <= not(layer0_outputs(4252));
    layer1_outputs(4731) <= not((layer0_outputs(3036)) and (layer0_outputs(832)));
    layer1_outputs(4732) <= (layer0_outputs(4210)) and not (layer0_outputs(4865));
    layer1_outputs(4733) <= layer0_outputs(3801);
    layer1_outputs(4734) <= not(layer0_outputs(4846));
    layer1_outputs(4735) <= layer0_outputs(2062);
    layer1_outputs(4736) <= (layer0_outputs(3712)) or (layer0_outputs(4269));
    layer1_outputs(4737) <= not(layer0_outputs(2677));
    layer1_outputs(4738) <= not((layer0_outputs(905)) and (layer0_outputs(1397)));
    layer1_outputs(4739) <= not(layer0_outputs(1078));
    layer1_outputs(4740) <= layer0_outputs(1985);
    layer1_outputs(4741) <= not(layer0_outputs(724)) or (layer0_outputs(1258));
    layer1_outputs(4742) <= not(layer0_outputs(4472));
    layer1_outputs(4743) <= not((layer0_outputs(1222)) or (layer0_outputs(1980)));
    layer1_outputs(4744) <= not(layer0_outputs(1868));
    layer1_outputs(4745) <= (layer0_outputs(1150)) and (layer0_outputs(3090));
    layer1_outputs(4746) <= layer0_outputs(1868);
    layer1_outputs(4747) <= (layer0_outputs(1899)) and not (layer0_outputs(3526));
    layer1_outputs(4748) <= (layer0_outputs(1212)) or (layer0_outputs(3807));
    layer1_outputs(4749) <= not((layer0_outputs(1757)) or (layer0_outputs(3033)));
    layer1_outputs(4750) <= not(layer0_outputs(1221));
    layer1_outputs(4751) <= not(layer0_outputs(4227));
    layer1_outputs(4752) <= not(layer0_outputs(4000));
    layer1_outputs(4753) <= not(layer0_outputs(4915));
    layer1_outputs(4754) <= not((layer0_outputs(4232)) xor (layer0_outputs(37)));
    layer1_outputs(4755) <= not(layer0_outputs(769)) or (layer0_outputs(2657));
    layer1_outputs(4756) <= not(layer0_outputs(4675)) or (layer0_outputs(1898));
    layer1_outputs(4757) <= layer0_outputs(3522);
    layer1_outputs(4758) <= layer0_outputs(4252);
    layer1_outputs(4759) <= (layer0_outputs(4659)) and not (layer0_outputs(2070));
    layer1_outputs(4760) <= not(layer0_outputs(672));
    layer1_outputs(4761) <= (layer0_outputs(430)) and (layer0_outputs(1476));
    layer1_outputs(4762) <= not((layer0_outputs(569)) or (layer0_outputs(1510)));
    layer1_outputs(4763) <= not((layer0_outputs(3932)) xor (layer0_outputs(1886)));
    layer1_outputs(4764) <= not(layer0_outputs(4516));
    layer1_outputs(4765) <= not((layer0_outputs(376)) or (layer0_outputs(3915)));
    layer1_outputs(4766) <= not(layer0_outputs(1895));
    layer1_outputs(4767) <= not((layer0_outputs(2582)) and (layer0_outputs(4992)));
    layer1_outputs(4768) <= (layer0_outputs(2897)) and not (layer0_outputs(3710));
    layer1_outputs(4769) <= not((layer0_outputs(4842)) and (layer0_outputs(937)));
    layer1_outputs(4770) <= not((layer0_outputs(247)) xor (layer0_outputs(453)));
    layer1_outputs(4771) <= not((layer0_outputs(3248)) and (layer0_outputs(3661)));
    layer1_outputs(4772) <= not(layer0_outputs(2107)) or (layer0_outputs(2365));
    layer1_outputs(4773) <= not(layer0_outputs(469));
    layer1_outputs(4774) <= not((layer0_outputs(3445)) or (layer0_outputs(923)));
    layer1_outputs(4775) <= not((layer0_outputs(1637)) xor (layer0_outputs(4728)));
    layer1_outputs(4776) <= not((layer0_outputs(5050)) xor (layer0_outputs(1107)));
    layer1_outputs(4777) <= layer0_outputs(1076);
    layer1_outputs(4778) <= not(layer0_outputs(1135));
    layer1_outputs(4779) <= layer0_outputs(186);
    layer1_outputs(4780) <= (layer0_outputs(3616)) and not (layer0_outputs(502));
    layer1_outputs(4781) <= (layer0_outputs(138)) and not (layer0_outputs(57));
    layer1_outputs(4782) <= (layer0_outputs(1108)) and not (layer0_outputs(1093));
    layer1_outputs(4783) <= not(layer0_outputs(534));
    layer1_outputs(4784) <= (layer0_outputs(2288)) and (layer0_outputs(5043));
    layer1_outputs(4785) <= (layer0_outputs(1029)) and not (layer0_outputs(2449));
    layer1_outputs(4786) <= not(layer0_outputs(2767));
    layer1_outputs(4787) <= layer0_outputs(228);
    layer1_outputs(4788) <= (layer0_outputs(3358)) xor (layer0_outputs(3787));
    layer1_outputs(4789) <= not(layer0_outputs(1127));
    layer1_outputs(4790) <= layer0_outputs(1540);
    layer1_outputs(4791) <= not((layer0_outputs(62)) and (layer0_outputs(3650)));
    layer1_outputs(4792) <= not(layer0_outputs(3552));
    layer1_outputs(4793) <= not(layer0_outputs(1001));
    layer1_outputs(4794) <= (layer0_outputs(4858)) or (layer0_outputs(5110));
    layer1_outputs(4795) <= not((layer0_outputs(1384)) and (layer0_outputs(227)));
    layer1_outputs(4796) <= not(layer0_outputs(1458)) or (layer0_outputs(31));
    layer1_outputs(4797) <= not((layer0_outputs(1440)) and (layer0_outputs(254)));
    layer1_outputs(4798) <= not((layer0_outputs(80)) xor (layer0_outputs(3881)));
    layer1_outputs(4799) <= not((layer0_outputs(185)) or (layer0_outputs(3590)));
    layer1_outputs(4800) <= not(layer0_outputs(1597));
    layer1_outputs(4801) <= '0';
    layer1_outputs(4802) <= layer0_outputs(4518);
    layer1_outputs(4803) <= (layer0_outputs(1462)) and not (layer0_outputs(1731));
    layer1_outputs(4804) <= not((layer0_outputs(4605)) and (layer0_outputs(2910)));
    layer1_outputs(4805) <= not(layer0_outputs(1072));
    layer1_outputs(4806) <= layer0_outputs(1846);
    layer1_outputs(4807) <= (layer0_outputs(3067)) and not (layer0_outputs(3145));
    layer1_outputs(4808) <= layer0_outputs(63);
    layer1_outputs(4809) <= (layer0_outputs(1780)) and not (layer0_outputs(1867));
    layer1_outputs(4810) <= not((layer0_outputs(2733)) xor (layer0_outputs(1116)));
    layer1_outputs(4811) <= '0';
    layer1_outputs(4812) <= not((layer0_outputs(2564)) or (layer0_outputs(282)));
    layer1_outputs(4813) <= (layer0_outputs(3115)) and not (layer0_outputs(1610));
    layer1_outputs(4814) <= not(layer0_outputs(4230)) or (layer0_outputs(3588));
    layer1_outputs(4815) <= not(layer0_outputs(4946)) or (layer0_outputs(2506));
    layer1_outputs(4816) <= layer0_outputs(2013);
    layer1_outputs(4817) <= not((layer0_outputs(1961)) xor (layer0_outputs(497)));
    layer1_outputs(4818) <= not(layer0_outputs(428)) or (layer0_outputs(2705));
    layer1_outputs(4819) <= '0';
    layer1_outputs(4820) <= not(layer0_outputs(1217));
    layer1_outputs(4821) <= (layer0_outputs(4591)) and not (layer0_outputs(54));
    layer1_outputs(4822) <= (layer0_outputs(1436)) or (layer0_outputs(4511));
    layer1_outputs(4823) <= not(layer0_outputs(3897)) or (layer0_outputs(1507));
    layer1_outputs(4824) <= layer0_outputs(4976);
    layer1_outputs(4825) <= not((layer0_outputs(1181)) xor (layer0_outputs(3163)));
    layer1_outputs(4826) <= not((layer0_outputs(232)) xor (layer0_outputs(3455)));
    layer1_outputs(4827) <= layer0_outputs(3440);
    layer1_outputs(4828) <= (layer0_outputs(4918)) xor (layer0_outputs(2821));
    layer1_outputs(4829) <= not((layer0_outputs(2925)) and (layer0_outputs(2369)));
    layer1_outputs(4830) <= '0';
    layer1_outputs(4831) <= not(layer0_outputs(392));
    layer1_outputs(4832) <= (layer0_outputs(123)) and not (layer0_outputs(39));
    layer1_outputs(4833) <= (layer0_outputs(302)) xor (layer0_outputs(211));
    layer1_outputs(4834) <= not(layer0_outputs(2021));
    layer1_outputs(4835) <= not((layer0_outputs(2071)) or (layer0_outputs(3233)));
    layer1_outputs(4836) <= layer0_outputs(2121);
    layer1_outputs(4837) <= '0';
    layer1_outputs(4838) <= (layer0_outputs(69)) xor (layer0_outputs(4728));
    layer1_outputs(4839) <= not(layer0_outputs(3447)) or (layer0_outputs(4231));
    layer1_outputs(4840) <= not(layer0_outputs(1681));
    layer1_outputs(4841) <= not((layer0_outputs(332)) or (layer0_outputs(1043)));
    layer1_outputs(4842) <= layer0_outputs(2863);
    layer1_outputs(4843) <= not((layer0_outputs(2574)) or (layer0_outputs(19)));
    layer1_outputs(4844) <= '1';
    layer1_outputs(4845) <= not((layer0_outputs(3374)) or (layer0_outputs(1262)));
    layer1_outputs(4846) <= layer0_outputs(4389);
    layer1_outputs(4847) <= layer0_outputs(2418);
    layer1_outputs(4848) <= not((layer0_outputs(4693)) xor (layer0_outputs(4095)));
    layer1_outputs(4849) <= (layer0_outputs(1316)) xor (layer0_outputs(1206));
    layer1_outputs(4850) <= layer0_outputs(4138);
    layer1_outputs(4851) <= '0';
    layer1_outputs(4852) <= layer0_outputs(531);
    layer1_outputs(4853) <= (layer0_outputs(2252)) xor (layer0_outputs(3176));
    layer1_outputs(4854) <= layer0_outputs(388);
    layer1_outputs(4855) <= (layer0_outputs(4627)) and not (layer0_outputs(2601));
    layer1_outputs(4856) <= not(layer0_outputs(3397));
    layer1_outputs(4857) <= not((layer0_outputs(4895)) and (layer0_outputs(4914)));
    layer1_outputs(4858) <= (layer0_outputs(4974)) and (layer0_outputs(313));
    layer1_outputs(4859) <= (layer0_outputs(3892)) and not (layer0_outputs(4983));
    layer1_outputs(4860) <= (layer0_outputs(1503)) or (layer0_outputs(2018));
    layer1_outputs(4861) <= '0';
    layer1_outputs(4862) <= not(layer0_outputs(3451));
    layer1_outputs(4863) <= not(layer0_outputs(3848));
    layer1_outputs(4864) <= not((layer0_outputs(2507)) xor (layer0_outputs(585)));
    layer1_outputs(4865) <= (layer0_outputs(4095)) and (layer0_outputs(1332));
    layer1_outputs(4866) <= layer0_outputs(2274);
    layer1_outputs(4867) <= layer0_outputs(3907);
    layer1_outputs(4868) <= (layer0_outputs(2296)) and (layer0_outputs(590));
    layer1_outputs(4869) <= not(layer0_outputs(1137));
    layer1_outputs(4870) <= (layer0_outputs(1686)) or (layer0_outputs(3918));
    layer1_outputs(4871) <= '0';
    layer1_outputs(4872) <= not(layer0_outputs(4726)) or (layer0_outputs(2241));
    layer1_outputs(4873) <= not(layer0_outputs(50)) or (layer0_outputs(3768));
    layer1_outputs(4874) <= (layer0_outputs(4442)) or (layer0_outputs(635));
    layer1_outputs(4875) <= not((layer0_outputs(3680)) and (layer0_outputs(747)));
    layer1_outputs(4876) <= not(layer0_outputs(3232)) or (layer0_outputs(543));
    layer1_outputs(4877) <= layer0_outputs(279);
    layer1_outputs(4878) <= not(layer0_outputs(3668));
    layer1_outputs(4879) <= (layer0_outputs(1319)) and not (layer0_outputs(2100));
    layer1_outputs(4880) <= layer0_outputs(2754);
    layer1_outputs(4881) <= not(layer0_outputs(3114));
    layer1_outputs(4882) <= (layer0_outputs(1092)) and (layer0_outputs(3104));
    layer1_outputs(4883) <= layer0_outputs(2291);
    layer1_outputs(4884) <= not((layer0_outputs(1529)) or (layer0_outputs(3043)));
    layer1_outputs(4885) <= layer0_outputs(5068);
    layer1_outputs(4886) <= not((layer0_outputs(3731)) and (layer0_outputs(524)));
    layer1_outputs(4887) <= (layer0_outputs(2329)) or (layer0_outputs(498));
    layer1_outputs(4888) <= not(layer0_outputs(4738));
    layer1_outputs(4889) <= (layer0_outputs(2384)) and not (layer0_outputs(609));
    layer1_outputs(4890) <= not((layer0_outputs(2593)) and (layer0_outputs(1189)));
    layer1_outputs(4891) <= layer0_outputs(3015);
    layer1_outputs(4892) <= not(layer0_outputs(3514)) or (layer0_outputs(4611));
    layer1_outputs(4893) <= not((layer0_outputs(3563)) and (layer0_outputs(2965)));
    layer1_outputs(4894) <= (layer0_outputs(4519)) or (layer0_outputs(17));
    layer1_outputs(4895) <= not(layer0_outputs(2434)) or (layer0_outputs(1367));
    layer1_outputs(4896) <= layer0_outputs(2085);
    layer1_outputs(4897) <= (layer0_outputs(2802)) xor (layer0_outputs(2585));
    layer1_outputs(4898) <= '1';
    layer1_outputs(4899) <= not(layer0_outputs(2202));
    layer1_outputs(4900) <= not(layer0_outputs(2929)) or (layer0_outputs(29));
    layer1_outputs(4901) <= not((layer0_outputs(5072)) or (layer0_outputs(4503)));
    layer1_outputs(4902) <= (layer0_outputs(4364)) xor (layer0_outputs(510));
    layer1_outputs(4903) <= (layer0_outputs(3304)) and (layer0_outputs(3999));
    layer1_outputs(4904) <= '1';
    layer1_outputs(4905) <= not((layer0_outputs(2853)) xor (layer0_outputs(2884)));
    layer1_outputs(4906) <= (layer0_outputs(4934)) or (layer0_outputs(275));
    layer1_outputs(4907) <= layer0_outputs(4876);
    layer1_outputs(4908) <= (layer0_outputs(2178)) and not (layer0_outputs(3838));
    layer1_outputs(4909) <= not(layer0_outputs(1834));
    layer1_outputs(4910) <= '0';
    layer1_outputs(4911) <= not((layer0_outputs(754)) or (layer0_outputs(4439)));
    layer1_outputs(4912) <= not(layer0_outputs(4601)) or (layer0_outputs(900));
    layer1_outputs(4913) <= not((layer0_outputs(534)) xor (layer0_outputs(4951)));
    layer1_outputs(4914) <= (layer0_outputs(2555)) and (layer0_outputs(4251));
    layer1_outputs(4915) <= not(layer0_outputs(2899));
    layer1_outputs(4916) <= '1';
    layer1_outputs(4917) <= layer0_outputs(3821);
    layer1_outputs(4918) <= layer0_outputs(3255);
    layer1_outputs(4919) <= '0';
    layer1_outputs(4920) <= layer0_outputs(4625);
    layer1_outputs(4921) <= not(layer0_outputs(3084)) or (layer0_outputs(3535));
    layer1_outputs(4922) <= not(layer0_outputs(1094));
    layer1_outputs(4923) <= not(layer0_outputs(3901));
    layer1_outputs(4924) <= not((layer0_outputs(3050)) and (layer0_outputs(1415)));
    layer1_outputs(4925) <= not(layer0_outputs(2757)) or (layer0_outputs(3413));
    layer1_outputs(4926) <= not((layer0_outputs(936)) or (layer0_outputs(2953)));
    layer1_outputs(4927) <= (layer0_outputs(4198)) and (layer0_outputs(3906));
    layer1_outputs(4928) <= not(layer0_outputs(417)) or (layer0_outputs(4735));
    layer1_outputs(4929) <= not(layer0_outputs(3824));
    layer1_outputs(4930) <= (layer0_outputs(58)) and not (layer0_outputs(2303));
    layer1_outputs(4931) <= (layer0_outputs(4776)) and (layer0_outputs(3334));
    layer1_outputs(4932) <= layer0_outputs(1124);
    layer1_outputs(4933) <= (layer0_outputs(2941)) or (layer0_outputs(5076));
    layer1_outputs(4934) <= not(layer0_outputs(515)) or (layer0_outputs(4344));
    layer1_outputs(4935) <= not(layer0_outputs(3051));
    layer1_outputs(4936) <= layer0_outputs(2521);
    layer1_outputs(4937) <= not(layer0_outputs(1769));
    layer1_outputs(4938) <= not(layer0_outputs(2820)) or (layer0_outputs(2164));
    layer1_outputs(4939) <= (layer0_outputs(716)) and not (layer0_outputs(225));
    layer1_outputs(4940) <= (layer0_outputs(1558)) or (layer0_outputs(2143));
    layer1_outputs(4941) <= not((layer0_outputs(134)) xor (layer0_outputs(1587)));
    layer1_outputs(4942) <= not(layer0_outputs(1156));
    layer1_outputs(4943) <= (layer0_outputs(3721)) or (layer0_outputs(4574));
    layer1_outputs(4944) <= not(layer0_outputs(4807));
    layer1_outputs(4945) <= (layer0_outputs(3364)) or (layer0_outputs(4025));
    layer1_outputs(4946) <= not(layer0_outputs(1292));
    layer1_outputs(4947) <= (layer0_outputs(555)) or (layer0_outputs(1825));
    layer1_outputs(4948) <= (layer0_outputs(4572)) and not (layer0_outputs(3408));
    layer1_outputs(4949) <= not(layer0_outputs(1420));
    layer1_outputs(4950) <= (layer0_outputs(3764)) and not (layer0_outputs(168));
    layer1_outputs(4951) <= (layer0_outputs(1315)) or (layer0_outputs(14));
    layer1_outputs(4952) <= layer0_outputs(3398);
    layer1_outputs(4953) <= (layer0_outputs(4955)) xor (layer0_outputs(3895));
    layer1_outputs(4954) <= (layer0_outputs(1853)) and not (layer0_outputs(3815));
    layer1_outputs(4955) <= not((layer0_outputs(4260)) xor (layer0_outputs(2254)));
    layer1_outputs(4956) <= (layer0_outputs(2455)) and not (layer0_outputs(1557));
    layer1_outputs(4957) <= '0';
    layer1_outputs(4958) <= layer0_outputs(4912);
    layer1_outputs(4959) <= '0';
    layer1_outputs(4960) <= layer0_outputs(3963);
    layer1_outputs(4961) <= (layer0_outputs(5025)) and not (layer0_outputs(1616));
    layer1_outputs(4962) <= not(layer0_outputs(8)) or (layer0_outputs(1182));
    layer1_outputs(4963) <= layer0_outputs(885);
    layer1_outputs(4964) <= layer0_outputs(643);
    layer1_outputs(4965) <= (layer0_outputs(461)) xor (layer0_outputs(4588));
    layer1_outputs(4966) <= not((layer0_outputs(503)) or (layer0_outputs(2221)));
    layer1_outputs(4967) <= (layer0_outputs(2163)) and not (layer0_outputs(340));
    layer1_outputs(4968) <= not(layer0_outputs(430));
    layer1_outputs(4969) <= not(layer0_outputs(4224)) or (layer0_outputs(4850));
    layer1_outputs(4970) <= (layer0_outputs(1052)) and (layer0_outputs(4798));
    layer1_outputs(4971) <= layer0_outputs(676);
    layer1_outputs(4972) <= (layer0_outputs(2831)) and (layer0_outputs(1158));
    layer1_outputs(4973) <= not(layer0_outputs(2927));
    layer1_outputs(4974) <= layer0_outputs(3546);
    layer1_outputs(4975) <= not(layer0_outputs(2528));
    layer1_outputs(4976) <= (layer0_outputs(4019)) xor (layer0_outputs(337));
    layer1_outputs(4977) <= not(layer0_outputs(3186));
    layer1_outputs(4978) <= not(layer0_outputs(3691)) or (layer0_outputs(3481));
    layer1_outputs(4979) <= not((layer0_outputs(2084)) xor (layer0_outputs(3963)));
    layer1_outputs(4980) <= layer0_outputs(236);
    layer1_outputs(4981) <= (layer0_outputs(2023)) and (layer0_outputs(115));
    layer1_outputs(4982) <= (layer0_outputs(1825)) and (layer0_outputs(4790));
    layer1_outputs(4983) <= (layer0_outputs(1927)) and (layer0_outputs(2180));
    layer1_outputs(4984) <= (layer0_outputs(2127)) xor (layer0_outputs(140));
    layer1_outputs(4985) <= not(layer0_outputs(4604)) or (layer0_outputs(4340));
    layer1_outputs(4986) <= (layer0_outputs(4467)) xor (layer0_outputs(868));
    layer1_outputs(4987) <= not((layer0_outputs(3100)) xor (layer0_outputs(992)));
    layer1_outputs(4988) <= '1';
    layer1_outputs(4989) <= (layer0_outputs(4620)) or (layer0_outputs(3713));
    layer1_outputs(4990) <= '0';
    layer1_outputs(4991) <= (layer0_outputs(1832)) and not (layer0_outputs(1545));
    layer1_outputs(4992) <= not((layer0_outputs(676)) or (layer0_outputs(1816)));
    layer1_outputs(4993) <= not((layer0_outputs(3687)) and (layer0_outputs(463)));
    layer1_outputs(4994) <= not(layer0_outputs(1937));
    layer1_outputs(4995) <= layer0_outputs(4893);
    layer1_outputs(4996) <= (layer0_outputs(694)) and not (layer0_outputs(4592));
    layer1_outputs(4997) <= not(layer0_outputs(1607)) or (layer0_outputs(3906));
    layer1_outputs(4998) <= '0';
    layer1_outputs(4999) <= layer0_outputs(4399);
    layer1_outputs(5000) <= (layer0_outputs(1694)) or (layer0_outputs(1765));
    layer1_outputs(5001) <= (layer0_outputs(1777)) and not (layer0_outputs(1858));
    layer1_outputs(5002) <= layer0_outputs(1538);
    layer1_outputs(5003) <= layer0_outputs(2262);
    layer1_outputs(5004) <= not(layer0_outputs(1639));
    layer1_outputs(5005) <= layer0_outputs(5062);
    layer1_outputs(5006) <= (layer0_outputs(1521)) and not (layer0_outputs(1398));
    layer1_outputs(5007) <= (layer0_outputs(913)) and not (layer0_outputs(204));
    layer1_outputs(5008) <= not((layer0_outputs(4349)) xor (layer0_outputs(538)));
    layer1_outputs(5009) <= not(layer0_outputs(3844));
    layer1_outputs(5010) <= layer0_outputs(2127);
    layer1_outputs(5011) <= (layer0_outputs(1341)) xor (layer0_outputs(1657));
    layer1_outputs(5012) <= (layer0_outputs(1805)) or (layer0_outputs(4474));
    layer1_outputs(5013) <= not(layer0_outputs(772)) or (layer0_outputs(4639));
    layer1_outputs(5014) <= (layer0_outputs(4172)) or (layer0_outputs(1553));
    layer1_outputs(5015) <= layer0_outputs(1161);
    layer1_outputs(5016) <= '0';
    layer1_outputs(5017) <= layer0_outputs(4880);
    layer1_outputs(5018) <= not(layer0_outputs(727));
    layer1_outputs(5019) <= layer0_outputs(4090);
    layer1_outputs(5020) <= not((layer0_outputs(3478)) or (layer0_outputs(4588)));
    layer1_outputs(5021) <= layer0_outputs(4123);
    layer1_outputs(5022) <= layer0_outputs(805);
    layer1_outputs(5023) <= layer0_outputs(312);
    layer1_outputs(5024) <= (layer0_outputs(243)) and not (layer0_outputs(2564));
    layer1_outputs(5025) <= not((layer0_outputs(986)) and (layer0_outputs(3528)));
    layer1_outputs(5026) <= not((layer0_outputs(3354)) or (layer0_outputs(2294)));
    layer1_outputs(5027) <= not((layer0_outputs(1622)) or (layer0_outputs(1396)));
    layer1_outputs(5028) <= not((layer0_outputs(2822)) or (layer0_outputs(4493)));
    layer1_outputs(5029) <= not(layer0_outputs(2726));
    layer1_outputs(5030) <= (layer0_outputs(4744)) and not (layer0_outputs(1028));
    layer1_outputs(5031) <= not(layer0_outputs(3241)) or (layer0_outputs(1510));
    layer1_outputs(5032) <= (layer0_outputs(4221)) and (layer0_outputs(1916));
    layer1_outputs(5033) <= layer0_outputs(3494);
    layer1_outputs(5034) <= layer0_outputs(3630);
    layer1_outputs(5035) <= (layer0_outputs(763)) and not (layer0_outputs(4145));
    layer1_outputs(5036) <= not((layer0_outputs(3675)) xor (layer0_outputs(4005)));
    layer1_outputs(5037) <= not((layer0_outputs(3433)) or (layer0_outputs(4408)));
    layer1_outputs(5038) <= not(layer0_outputs(3893));
    layer1_outputs(5039) <= not((layer0_outputs(3006)) or (layer0_outputs(3712)));
    layer1_outputs(5040) <= not(layer0_outputs(3431));
    layer1_outputs(5041) <= layer0_outputs(1635);
    layer1_outputs(5042) <= '1';
    layer1_outputs(5043) <= not((layer0_outputs(3598)) and (layer0_outputs(677)));
    layer1_outputs(5044) <= (layer0_outputs(3467)) and not (layer0_outputs(262));
    layer1_outputs(5045) <= layer0_outputs(2112);
    layer1_outputs(5046) <= not((layer0_outputs(2968)) and (layer0_outputs(1318)));
    layer1_outputs(5047) <= not((layer0_outputs(2855)) xor (layer0_outputs(3280)));
    layer1_outputs(5048) <= (layer0_outputs(5119)) and (layer0_outputs(3725));
    layer1_outputs(5049) <= (layer0_outputs(2135)) and (layer0_outputs(3872));
    layer1_outputs(5050) <= (layer0_outputs(175)) or (layer0_outputs(2003));
    layer1_outputs(5051) <= not((layer0_outputs(3896)) and (layer0_outputs(584)));
    layer1_outputs(5052) <= not(layer0_outputs(1286));
    layer1_outputs(5053) <= (layer0_outputs(1679)) and not (layer0_outputs(1775));
    layer1_outputs(5054) <= not((layer0_outputs(4689)) or (layer0_outputs(3079)));
    layer1_outputs(5055) <= not(layer0_outputs(2974));
    layer1_outputs(5056) <= (layer0_outputs(4164)) or (layer0_outputs(4243));
    layer1_outputs(5057) <= not(layer0_outputs(4928));
    layer1_outputs(5058) <= not(layer0_outputs(1038)) or (layer0_outputs(2176));
    layer1_outputs(5059) <= layer0_outputs(1416);
    layer1_outputs(5060) <= not(layer0_outputs(4607)) or (layer0_outputs(2392));
    layer1_outputs(5061) <= layer0_outputs(3287);
    layer1_outputs(5062) <= not((layer0_outputs(4226)) or (layer0_outputs(3564)));
    layer1_outputs(5063) <= (layer0_outputs(1152)) or (layer0_outputs(501));
    layer1_outputs(5064) <= layer0_outputs(1213);
    layer1_outputs(5065) <= '1';
    layer1_outputs(5066) <= (layer0_outputs(4671)) or (layer0_outputs(2255));
    layer1_outputs(5067) <= (layer0_outputs(1560)) and (layer0_outputs(4715));
    layer1_outputs(5068) <= not((layer0_outputs(3968)) xor (layer0_outputs(2182)));
    layer1_outputs(5069) <= (layer0_outputs(1115)) and not (layer0_outputs(3955));
    layer1_outputs(5070) <= (layer0_outputs(3196)) or (layer0_outputs(4968));
    layer1_outputs(5071) <= not((layer0_outputs(4896)) and (layer0_outputs(2577)));
    layer1_outputs(5072) <= (layer0_outputs(3841)) or (layer0_outputs(4272));
    layer1_outputs(5073) <= not((layer0_outputs(4393)) xor (layer0_outputs(201)));
    layer1_outputs(5074) <= (layer0_outputs(4978)) and not (layer0_outputs(416));
    layer1_outputs(5075) <= not((layer0_outputs(2918)) or (layer0_outputs(3391)));
    layer1_outputs(5076) <= layer0_outputs(1414);
    layer1_outputs(5077) <= (layer0_outputs(2419)) and not (layer0_outputs(3556));
    layer1_outputs(5078) <= (layer0_outputs(1875)) xor (layer0_outputs(4257));
    layer1_outputs(5079) <= (layer0_outputs(1082)) and (layer0_outputs(899));
    layer1_outputs(5080) <= '0';
    layer1_outputs(5081) <= not((layer0_outputs(5118)) or (layer0_outputs(3262)));
    layer1_outputs(5082) <= not((layer0_outputs(2114)) xor (layer0_outputs(4641)));
    layer1_outputs(5083) <= not((layer0_outputs(1298)) or (layer0_outputs(4700)));
    layer1_outputs(5084) <= not(layer0_outputs(4315));
    layer1_outputs(5085) <= (layer0_outputs(4746)) and (layer0_outputs(499));
    layer1_outputs(5086) <= not(layer0_outputs(991));
    layer1_outputs(5087) <= '0';
    layer1_outputs(5088) <= not(layer0_outputs(192)) or (layer0_outputs(4892));
    layer1_outputs(5089) <= not(layer0_outputs(4778));
    layer1_outputs(5090) <= not(layer0_outputs(3196));
    layer1_outputs(5091) <= not(layer0_outputs(4253)) or (layer0_outputs(2516));
    layer1_outputs(5092) <= not((layer0_outputs(5010)) xor (layer0_outputs(439)));
    layer1_outputs(5093) <= not(layer0_outputs(1334)) or (layer0_outputs(2872));
    layer1_outputs(5094) <= not((layer0_outputs(363)) or (layer0_outputs(1782)));
    layer1_outputs(5095) <= not((layer0_outputs(3818)) xor (layer0_outputs(969)));
    layer1_outputs(5096) <= not(layer0_outputs(4737)) or (layer0_outputs(4989));
    layer1_outputs(5097) <= not((layer0_outputs(3779)) and (layer0_outputs(2313)));
    layer1_outputs(5098) <= layer0_outputs(426);
    layer1_outputs(5099) <= (layer0_outputs(2668)) or (layer0_outputs(5102));
    layer1_outputs(5100) <= not((layer0_outputs(3422)) or (layer0_outputs(229)));
    layer1_outputs(5101) <= (layer0_outputs(1059)) xor (layer0_outputs(3702));
    layer1_outputs(5102) <= not(layer0_outputs(2407));
    layer1_outputs(5103) <= layer0_outputs(3953);
    layer1_outputs(5104) <= (layer0_outputs(3959)) and not (layer0_outputs(4495));
    layer1_outputs(5105) <= layer0_outputs(4309);
    layer1_outputs(5106) <= not(layer0_outputs(4313));
    layer1_outputs(5107) <= layer0_outputs(4488);
    layer1_outputs(5108) <= not((layer0_outputs(1835)) or (layer0_outputs(1596)));
    layer1_outputs(5109) <= layer0_outputs(1674);
    layer1_outputs(5110) <= (layer0_outputs(2087)) and not (layer0_outputs(1754));
    layer1_outputs(5111) <= (layer0_outputs(5104)) and not (layer0_outputs(4650));
    layer1_outputs(5112) <= layer0_outputs(3474);
    layer1_outputs(5113) <= layer0_outputs(4066);
    layer1_outputs(5114) <= (layer0_outputs(1509)) and not (layer0_outputs(1563));
    layer1_outputs(5115) <= (layer0_outputs(1864)) or (layer0_outputs(2916));
    layer1_outputs(5116) <= (layer0_outputs(2359)) xor (layer0_outputs(4436));
    layer1_outputs(5117) <= not(layer0_outputs(1900));
    layer1_outputs(5118) <= not(layer0_outputs(1733));
    layer1_outputs(5119) <= not(layer0_outputs(2509)) or (layer0_outputs(995));
    layer2_outputs(0) <= not(layer1_outputs(1783));
    layer2_outputs(1) <= (layer1_outputs(2083)) and not (layer1_outputs(2511));
    layer2_outputs(2) <= layer1_outputs(547);
    layer2_outputs(3) <= (layer1_outputs(2846)) or (layer1_outputs(3378));
    layer2_outputs(4) <= not(layer1_outputs(3743)) or (layer1_outputs(3937));
    layer2_outputs(5) <= not((layer1_outputs(3530)) xor (layer1_outputs(2554)));
    layer2_outputs(6) <= (layer1_outputs(1046)) or (layer1_outputs(141));
    layer2_outputs(7) <= not(layer1_outputs(3896));
    layer2_outputs(8) <= (layer1_outputs(367)) and not (layer1_outputs(2629));
    layer2_outputs(9) <= not(layer1_outputs(2475));
    layer2_outputs(10) <= not(layer1_outputs(4267)) or (layer1_outputs(4810));
    layer2_outputs(11) <= layer1_outputs(2781);
    layer2_outputs(12) <= (layer1_outputs(2249)) and not (layer1_outputs(2385));
    layer2_outputs(13) <= not(layer1_outputs(4843));
    layer2_outputs(14) <= not(layer1_outputs(2947));
    layer2_outputs(15) <= (layer1_outputs(2260)) or (layer1_outputs(1480));
    layer2_outputs(16) <= not(layer1_outputs(491));
    layer2_outputs(17) <= not(layer1_outputs(3868));
    layer2_outputs(18) <= (layer1_outputs(3126)) or (layer1_outputs(4482));
    layer2_outputs(19) <= (layer1_outputs(4487)) xor (layer1_outputs(485));
    layer2_outputs(20) <= (layer1_outputs(699)) xor (layer1_outputs(337));
    layer2_outputs(21) <= (layer1_outputs(3778)) and not (layer1_outputs(2040));
    layer2_outputs(22) <= layer1_outputs(1974);
    layer2_outputs(23) <= not(layer1_outputs(3998)) or (layer1_outputs(4738));
    layer2_outputs(24) <= layer1_outputs(867);
    layer2_outputs(25) <= not(layer1_outputs(250));
    layer2_outputs(26) <= not((layer1_outputs(3882)) and (layer1_outputs(1871)));
    layer2_outputs(27) <= not(layer1_outputs(4061)) or (layer1_outputs(695));
    layer2_outputs(28) <= (layer1_outputs(1684)) or (layer1_outputs(765));
    layer2_outputs(29) <= layer1_outputs(4399);
    layer2_outputs(30) <= (layer1_outputs(1948)) xor (layer1_outputs(707));
    layer2_outputs(31) <= (layer1_outputs(3107)) and (layer1_outputs(2340));
    layer2_outputs(32) <= (layer1_outputs(3647)) and (layer1_outputs(1814));
    layer2_outputs(33) <= layer1_outputs(3019);
    layer2_outputs(34) <= not(layer1_outputs(2750));
    layer2_outputs(35) <= not(layer1_outputs(3283));
    layer2_outputs(36) <= (layer1_outputs(2759)) and not (layer1_outputs(5087));
    layer2_outputs(37) <= not(layer1_outputs(1461));
    layer2_outputs(38) <= (layer1_outputs(3537)) and not (layer1_outputs(3809));
    layer2_outputs(39) <= not(layer1_outputs(3056));
    layer2_outputs(40) <= (layer1_outputs(1120)) xor (layer1_outputs(3856));
    layer2_outputs(41) <= layer1_outputs(1840);
    layer2_outputs(42) <= layer1_outputs(1779);
    layer2_outputs(43) <= not((layer1_outputs(839)) and (layer1_outputs(3206)));
    layer2_outputs(44) <= not(layer1_outputs(725));
    layer2_outputs(45) <= layer1_outputs(1096);
    layer2_outputs(46) <= layer1_outputs(4647);
    layer2_outputs(47) <= (layer1_outputs(4588)) and not (layer1_outputs(4409));
    layer2_outputs(48) <= not(layer1_outputs(4141));
    layer2_outputs(49) <= not(layer1_outputs(1748));
    layer2_outputs(50) <= not(layer1_outputs(712));
    layer2_outputs(51) <= not((layer1_outputs(455)) or (layer1_outputs(5024)));
    layer2_outputs(52) <= not(layer1_outputs(2354));
    layer2_outputs(53) <= not((layer1_outputs(2787)) and (layer1_outputs(418)));
    layer2_outputs(54) <= (layer1_outputs(5091)) xor (layer1_outputs(3395));
    layer2_outputs(55) <= not(layer1_outputs(4732));
    layer2_outputs(56) <= layer1_outputs(2173);
    layer2_outputs(57) <= layer1_outputs(1801);
    layer2_outputs(58) <= layer1_outputs(2535);
    layer2_outputs(59) <= (layer1_outputs(3180)) and (layer1_outputs(3515));
    layer2_outputs(60) <= not((layer1_outputs(2292)) xor (layer1_outputs(573)));
    layer2_outputs(61) <= (layer1_outputs(163)) and (layer1_outputs(4026));
    layer2_outputs(62) <= not(layer1_outputs(918));
    layer2_outputs(63) <= '0';
    layer2_outputs(64) <= layer1_outputs(4930);
    layer2_outputs(65) <= (layer1_outputs(1605)) and not (layer1_outputs(2416));
    layer2_outputs(66) <= (layer1_outputs(250)) xor (layer1_outputs(4193));
    layer2_outputs(67) <= not(layer1_outputs(1428)) or (layer1_outputs(2357));
    layer2_outputs(68) <= not(layer1_outputs(5034));
    layer2_outputs(69) <= not(layer1_outputs(4991));
    layer2_outputs(70) <= not((layer1_outputs(4891)) or (layer1_outputs(898)));
    layer2_outputs(71) <= layer1_outputs(4711);
    layer2_outputs(72) <= layer1_outputs(1004);
    layer2_outputs(73) <= not((layer1_outputs(1578)) and (layer1_outputs(31)));
    layer2_outputs(74) <= layer1_outputs(1753);
    layer2_outputs(75) <= (layer1_outputs(4388)) and not (layer1_outputs(2360));
    layer2_outputs(76) <= (layer1_outputs(2995)) or (layer1_outputs(1851));
    layer2_outputs(77) <= layer1_outputs(3598);
    layer2_outputs(78) <= (layer1_outputs(4135)) and (layer1_outputs(1089));
    layer2_outputs(79) <= not((layer1_outputs(907)) xor (layer1_outputs(2293)));
    layer2_outputs(80) <= not(layer1_outputs(840)) or (layer1_outputs(687));
    layer2_outputs(81) <= not(layer1_outputs(2624));
    layer2_outputs(82) <= (layer1_outputs(3480)) and not (layer1_outputs(4753));
    layer2_outputs(83) <= layer1_outputs(2082);
    layer2_outputs(84) <= (layer1_outputs(2623)) and (layer1_outputs(4717));
    layer2_outputs(85) <= not(layer1_outputs(4701)) or (layer1_outputs(1643));
    layer2_outputs(86) <= layer1_outputs(3954);
    layer2_outputs(87) <= layer1_outputs(3411);
    layer2_outputs(88) <= layer1_outputs(2665);
    layer2_outputs(89) <= layer1_outputs(4401);
    layer2_outputs(90) <= layer1_outputs(3717);
    layer2_outputs(91) <= (layer1_outputs(3123)) and (layer1_outputs(1558));
    layer2_outputs(92) <= (layer1_outputs(4683)) and not (layer1_outputs(841));
    layer2_outputs(93) <= layer1_outputs(4211);
    layer2_outputs(94) <= not(layer1_outputs(3001));
    layer2_outputs(95) <= layer1_outputs(4216);
    layer2_outputs(96) <= layer1_outputs(4728);
    layer2_outputs(97) <= not(layer1_outputs(4799));
    layer2_outputs(98) <= (layer1_outputs(3613)) or (layer1_outputs(3987));
    layer2_outputs(99) <= layer1_outputs(325);
    layer2_outputs(100) <= (layer1_outputs(1173)) or (layer1_outputs(4243));
    layer2_outputs(101) <= not(layer1_outputs(2325));
    layer2_outputs(102) <= not(layer1_outputs(701));
    layer2_outputs(103) <= (layer1_outputs(854)) xor (layer1_outputs(2346));
    layer2_outputs(104) <= layer1_outputs(54);
    layer2_outputs(105) <= not(layer1_outputs(3192));
    layer2_outputs(106) <= layer1_outputs(3997);
    layer2_outputs(107) <= layer1_outputs(2124);
    layer2_outputs(108) <= layer1_outputs(305);
    layer2_outputs(109) <= (layer1_outputs(78)) and not (layer1_outputs(4541));
    layer2_outputs(110) <= layer1_outputs(4784);
    layer2_outputs(111) <= (layer1_outputs(4193)) xor (layer1_outputs(3184));
    layer2_outputs(112) <= not(layer1_outputs(4434));
    layer2_outputs(113) <= not((layer1_outputs(2709)) xor (layer1_outputs(3818)));
    layer2_outputs(114) <= (layer1_outputs(358)) xor (layer1_outputs(3654));
    layer2_outputs(115) <= layer1_outputs(3315);
    layer2_outputs(116) <= not(layer1_outputs(1168));
    layer2_outputs(117) <= not(layer1_outputs(4563)) or (layer1_outputs(640));
    layer2_outputs(118) <= not(layer1_outputs(3721)) or (layer1_outputs(4689));
    layer2_outputs(119) <= layer1_outputs(4331);
    layer2_outputs(120) <= (layer1_outputs(3341)) and not (layer1_outputs(4464));
    layer2_outputs(121) <= '1';
    layer2_outputs(122) <= not((layer1_outputs(2196)) and (layer1_outputs(3977)));
    layer2_outputs(123) <= (layer1_outputs(4113)) and not (layer1_outputs(874));
    layer2_outputs(124) <= not((layer1_outputs(787)) or (layer1_outputs(4884)));
    layer2_outputs(125) <= layer1_outputs(256);
    layer2_outputs(126) <= not(layer1_outputs(4552)) or (layer1_outputs(2691));
    layer2_outputs(127) <= layer1_outputs(563);
    layer2_outputs(128) <= layer1_outputs(1535);
    layer2_outputs(129) <= not((layer1_outputs(3780)) or (layer1_outputs(1431)));
    layer2_outputs(130) <= not(layer1_outputs(4599));
    layer2_outputs(131) <= not(layer1_outputs(1440)) or (layer1_outputs(2170));
    layer2_outputs(132) <= layer1_outputs(1088);
    layer2_outputs(133) <= not(layer1_outputs(561)) or (layer1_outputs(4081));
    layer2_outputs(134) <= not((layer1_outputs(4495)) xor (layer1_outputs(3002)));
    layer2_outputs(135) <= layer1_outputs(3835);
    layer2_outputs(136) <= not((layer1_outputs(3960)) xor (layer1_outputs(3815)));
    layer2_outputs(137) <= not(layer1_outputs(690));
    layer2_outputs(138) <= '0';
    layer2_outputs(139) <= (layer1_outputs(469)) and not (layer1_outputs(1689));
    layer2_outputs(140) <= not(layer1_outputs(464)) or (layer1_outputs(3587));
    layer2_outputs(141) <= not(layer1_outputs(1331)) or (layer1_outputs(4889));
    layer2_outputs(142) <= not(layer1_outputs(1110));
    layer2_outputs(143) <= layer1_outputs(3903);
    layer2_outputs(144) <= not(layer1_outputs(932));
    layer2_outputs(145) <= layer1_outputs(3450);
    layer2_outputs(146) <= (layer1_outputs(619)) and (layer1_outputs(3071));
    layer2_outputs(147) <= (layer1_outputs(2635)) or (layer1_outputs(2653));
    layer2_outputs(148) <= not(layer1_outputs(4982));
    layer2_outputs(149) <= not(layer1_outputs(3574));
    layer2_outputs(150) <= not(layer1_outputs(2882));
    layer2_outputs(151) <= (layer1_outputs(1989)) or (layer1_outputs(2520));
    layer2_outputs(152) <= not(layer1_outputs(5020)) or (layer1_outputs(586));
    layer2_outputs(153) <= not((layer1_outputs(2931)) or (layer1_outputs(3330)));
    layer2_outputs(154) <= not((layer1_outputs(3414)) xor (layer1_outputs(687)));
    layer2_outputs(155) <= layer1_outputs(2798);
    layer2_outputs(156) <= not(layer1_outputs(2904));
    layer2_outputs(157) <= not(layer1_outputs(4144));
    layer2_outputs(158) <= (layer1_outputs(5103)) and not (layer1_outputs(4312));
    layer2_outputs(159) <= (layer1_outputs(4288)) and not (layer1_outputs(1809));
    layer2_outputs(160) <= not((layer1_outputs(25)) and (layer1_outputs(1894)));
    layer2_outputs(161) <= not(layer1_outputs(1055));
    layer2_outputs(162) <= (layer1_outputs(414)) xor (layer1_outputs(4819));
    layer2_outputs(163) <= layer1_outputs(3099);
    layer2_outputs(164) <= not(layer1_outputs(3648));
    layer2_outputs(165) <= layer1_outputs(2836);
    layer2_outputs(166) <= (layer1_outputs(1111)) or (layer1_outputs(4350));
    layer2_outputs(167) <= (layer1_outputs(4302)) xor (layer1_outputs(691));
    layer2_outputs(168) <= not(layer1_outputs(1417));
    layer2_outputs(169) <= layer1_outputs(4007);
    layer2_outputs(170) <= layer1_outputs(1628);
    layer2_outputs(171) <= (layer1_outputs(5034)) and not (layer1_outputs(3645));
    layer2_outputs(172) <= (layer1_outputs(2598)) xor (layer1_outputs(4391));
    layer2_outputs(173) <= layer1_outputs(3548);
    layer2_outputs(174) <= (layer1_outputs(2689)) and not (layer1_outputs(36));
    layer2_outputs(175) <= not(layer1_outputs(3));
    layer2_outputs(176) <= not((layer1_outputs(2840)) or (layer1_outputs(1722)));
    layer2_outputs(177) <= (layer1_outputs(1853)) and (layer1_outputs(1521));
    layer2_outputs(178) <= not(layer1_outputs(1703));
    layer2_outputs(179) <= layer1_outputs(3214);
    layer2_outputs(180) <= layer1_outputs(2773);
    layer2_outputs(181) <= (layer1_outputs(3615)) or (layer1_outputs(1465));
    layer2_outputs(182) <= not((layer1_outputs(4922)) or (layer1_outputs(2983)));
    layer2_outputs(183) <= '0';
    layer2_outputs(184) <= layer1_outputs(913);
    layer2_outputs(185) <= not((layer1_outputs(1257)) and (layer1_outputs(1483)));
    layer2_outputs(186) <= not(layer1_outputs(5016));
    layer2_outputs(187) <= not((layer1_outputs(119)) or (layer1_outputs(1910)));
    layer2_outputs(188) <= not((layer1_outputs(4485)) or (layer1_outputs(3319)));
    layer2_outputs(189) <= layer1_outputs(3990);
    layer2_outputs(190) <= layer1_outputs(1339);
    layer2_outputs(191) <= (layer1_outputs(4048)) xor (layer1_outputs(4758));
    layer2_outputs(192) <= '1';
    layer2_outputs(193) <= (layer1_outputs(953)) and not (layer1_outputs(2303));
    layer2_outputs(194) <= (layer1_outputs(1738)) and (layer1_outputs(679));
    layer2_outputs(195) <= layer1_outputs(3501);
    layer2_outputs(196) <= layer1_outputs(4149);
    layer2_outputs(197) <= layer1_outputs(4473);
    layer2_outputs(198) <= not(layer1_outputs(4901)) or (layer1_outputs(3176));
    layer2_outputs(199) <= layer1_outputs(1417);
    layer2_outputs(200) <= not(layer1_outputs(3362));
    layer2_outputs(201) <= not((layer1_outputs(927)) xor (layer1_outputs(5072)));
    layer2_outputs(202) <= layer1_outputs(2817);
    layer2_outputs(203) <= (layer1_outputs(4526)) xor (layer1_outputs(788));
    layer2_outputs(204) <= layer1_outputs(3360);
    layer2_outputs(205) <= not(layer1_outputs(3538));
    layer2_outputs(206) <= not(layer1_outputs(2728)) or (layer1_outputs(1099));
    layer2_outputs(207) <= (layer1_outputs(4342)) and not (layer1_outputs(2883));
    layer2_outputs(208) <= layer1_outputs(3727);
    layer2_outputs(209) <= layer1_outputs(3151);
    layer2_outputs(210) <= (layer1_outputs(656)) or (layer1_outputs(1900));
    layer2_outputs(211) <= not((layer1_outputs(1355)) xor (layer1_outputs(5)));
    layer2_outputs(212) <= layer1_outputs(641);
    layer2_outputs(213) <= not(layer1_outputs(2735));
    layer2_outputs(214) <= not((layer1_outputs(3307)) or (layer1_outputs(1113)));
    layer2_outputs(215) <= layer1_outputs(1245);
    layer2_outputs(216) <= not((layer1_outputs(376)) xor (layer1_outputs(4758)));
    layer2_outputs(217) <= layer1_outputs(2783);
    layer2_outputs(218) <= (layer1_outputs(138)) and (layer1_outputs(1124));
    layer2_outputs(219) <= not((layer1_outputs(4527)) or (layer1_outputs(1284)));
    layer2_outputs(220) <= (layer1_outputs(2295)) and (layer1_outputs(910));
    layer2_outputs(221) <= not((layer1_outputs(3691)) and (layer1_outputs(3475)));
    layer2_outputs(222) <= not(layer1_outputs(254));
    layer2_outputs(223) <= (layer1_outputs(1291)) xor (layer1_outputs(1736));
    layer2_outputs(224) <= not(layer1_outputs(360));
    layer2_outputs(225) <= not(layer1_outputs(1612));
    layer2_outputs(226) <= not(layer1_outputs(642)) or (layer1_outputs(4813));
    layer2_outputs(227) <= layer1_outputs(385);
    layer2_outputs(228) <= not(layer1_outputs(1626));
    layer2_outputs(229) <= not(layer1_outputs(852));
    layer2_outputs(230) <= not(layer1_outputs(4449));
    layer2_outputs(231) <= (layer1_outputs(1062)) xor (layer1_outputs(3751));
    layer2_outputs(232) <= not((layer1_outputs(739)) xor (layer1_outputs(1600)));
    layer2_outputs(233) <= (layer1_outputs(5017)) and not (layer1_outputs(2365));
    layer2_outputs(234) <= layer1_outputs(3734);
    layer2_outputs(235) <= layer1_outputs(1831);
    layer2_outputs(236) <= layer1_outputs(2658);
    layer2_outputs(237) <= layer1_outputs(2317);
    layer2_outputs(238) <= (layer1_outputs(2147)) and (layer1_outputs(766));
    layer2_outputs(239) <= layer1_outputs(4778);
    layer2_outputs(240) <= '0';
    layer2_outputs(241) <= layer1_outputs(444);
    layer2_outputs(242) <= layer1_outputs(3839);
    layer2_outputs(243) <= '1';
    layer2_outputs(244) <= not(layer1_outputs(1982));
    layer2_outputs(245) <= not(layer1_outputs(2319));
    layer2_outputs(246) <= (layer1_outputs(4630)) and (layer1_outputs(654));
    layer2_outputs(247) <= (layer1_outputs(2671)) and (layer1_outputs(3906));
    layer2_outputs(248) <= layer1_outputs(259);
    layer2_outputs(249) <= (layer1_outputs(1214)) xor (layer1_outputs(2801));
    layer2_outputs(250) <= not(layer1_outputs(4528));
    layer2_outputs(251) <= not((layer1_outputs(3127)) xor (layer1_outputs(2382)));
    layer2_outputs(252) <= not(layer1_outputs(342));
    layer2_outputs(253) <= (layer1_outputs(3880)) and not (layer1_outputs(1518));
    layer2_outputs(254) <= not(layer1_outputs(1271));
    layer2_outputs(255) <= layer1_outputs(1071);
    layer2_outputs(256) <= not(layer1_outputs(1261));
    layer2_outputs(257) <= not(layer1_outputs(3944)) or (layer1_outputs(4272));
    layer2_outputs(258) <= not((layer1_outputs(264)) xor (layer1_outputs(586)));
    layer2_outputs(259) <= layer1_outputs(1250);
    layer2_outputs(260) <= not(layer1_outputs(3889)) or (layer1_outputs(1758));
    layer2_outputs(261) <= (layer1_outputs(4403)) and not (layer1_outputs(2609));
    layer2_outputs(262) <= layer1_outputs(1145);
    layer2_outputs(263) <= layer1_outputs(3461);
    layer2_outputs(264) <= not(layer1_outputs(2342));
    layer2_outputs(265) <= (layer1_outputs(2965)) and not (layer1_outputs(2222));
    layer2_outputs(266) <= layer1_outputs(3995);
    layer2_outputs(267) <= layer1_outputs(1970);
    layer2_outputs(268) <= not(layer1_outputs(1163));
    layer2_outputs(269) <= (layer1_outputs(1038)) and not (layer1_outputs(249));
    layer2_outputs(270) <= (layer1_outputs(1797)) and (layer1_outputs(975));
    layer2_outputs(271) <= not(layer1_outputs(1818));
    layer2_outputs(272) <= layer1_outputs(12);
    layer2_outputs(273) <= layer1_outputs(3105);
    layer2_outputs(274) <= not(layer1_outputs(1582));
    layer2_outputs(275) <= (layer1_outputs(30)) and not (layer1_outputs(674));
    layer2_outputs(276) <= layer1_outputs(1635);
    layer2_outputs(277) <= (layer1_outputs(5016)) xor (layer1_outputs(2122));
    layer2_outputs(278) <= (layer1_outputs(3312)) xor (layer1_outputs(62));
    layer2_outputs(279) <= not(layer1_outputs(2518)) or (layer1_outputs(3972));
    layer2_outputs(280) <= layer1_outputs(3906);
    layer2_outputs(281) <= layer1_outputs(4011);
    layer2_outputs(282) <= not(layer1_outputs(2499)) or (layer1_outputs(4316));
    layer2_outputs(283) <= not((layer1_outputs(4880)) xor (layer1_outputs(316)));
    layer2_outputs(284) <= not(layer1_outputs(1256));
    layer2_outputs(285) <= not(layer1_outputs(1319));
    layer2_outputs(286) <= layer1_outputs(732);
    layer2_outputs(287) <= not((layer1_outputs(2919)) or (layer1_outputs(4504)));
    layer2_outputs(288) <= not(layer1_outputs(531));
    layer2_outputs(289) <= not((layer1_outputs(2436)) xor (layer1_outputs(4276)));
    layer2_outputs(290) <= layer1_outputs(4371);
    layer2_outputs(291) <= not((layer1_outputs(2997)) and (layer1_outputs(3592)));
    layer2_outputs(292) <= (layer1_outputs(3723)) and not (layer1_outputs(3213));
    layer2_outputs(293) <= not(layer1_outputs(4762));
    layer2_outputs(294) <= not(layer1_outputs(2797));
    layer2_outputs(295) <= not((layer1_outputs(4131)) xor (layer1_outputs(2828)));
    layer2_outputs(296) <= not((layer1_outputs(2140)) or (layer1_outputs(3337)));
    layer2_outputs(297) <= not(layer1_outputs(1519)) or (layer1_outputs(3399));
    layer2_outputs(298) <= not(layer1_outputs(95));
    layer2_outputs(299) <= (layer1_outputs(5091)) or (layer1_outputs(1956));
    layer2_outputs(300) <= layer1_outputs(353);
    layer2_outputs(301) <= not(layer1_outputs(3672)) or (layer1_outputs(4634));
    layer2_outputs(302) <= (layer1_outputs(4892)) and not (layer1_outputs(3885));
    layer2_outputs(303) <= (layer1_outputs(2930)) xor (layer1_outputs(550));
    layer2_outputs(304) <= layer1_outputs(395);
    layer2_outputs(305) <= not(layer1_outputs(1176));
    layer2_outputs(306) <= (layer1_outputs(1587)) and (layer1_outputs(2521));
    layer2_outputs(307) <= '0';
    layer2_outputs(308) <= not(layer1_outputs(2721));
    layer2_outputs(309) <= (layer1_outputs(4895)) or (layer1_outputs(3860));
    layer2_outputs(310) <= not((layer1_outputs(2169)) or (layer1_outputs(1069)));
    layer2_outputs(311) <= layer1_outputs(409);
    layer2_outputs(312) <= layer1_outputs(329);
    layer2_outputs(313) <= layer1_outputs(860);
    layer2_outputs(314) <= not(layer1_outputs(383));
    layer2_outputs(315) <= not(layer1_outputs(3441)) or (layer1_outputs(1348));
    layer2_outputs(316) <= not((layer1_outputs(4372)) and (layer1_outputs(3339)));
    layer2_outputs(317) <= layer1_outputs(3512);
    layer2_outputs(318) <= (layer1_outputs(2459)) or (layer1_outputs(1405));
    layer2_outputs(319) <= layer1_outputs(388);
    layer2_outputs(320) <= not(layer1_outputs(4213)) or (layer1_outputs(1832));
    layer2_outputs(321) <= (layer1_outputs(3945)) xor (layer1_outputs(4443));
    layer2_outputs(322) <= not((layer1_outputs(4238)) and (layer1_outputs(3057)));
    layer2_outputs(323) <= (layer1_outputs(2922)) and not (layer1_outputs(734));
    layer2_outputs(324) <= not((layer1_outputs(3660)) and (layer1_outputs(4986)));
    layer2_outputs(325) <= (layer1_outputs(3417)) or (layer1_outputs(1605));
    layer2_outputs(326) <= (layer1_outputs(4017)) or (layer1_outputs(2108));
    layer2_outputs(327) <= (layer1_outputs(3088)) xor (layer1_outputs(781));
    layer2_outputs(328) <= not(layer1_outputs(4025)) or (layer1_outputs(1449));
    layer2_outputs(329) <= layer1_outputs(4623);
    layer2_outputs(330) <= (layer1_outputs(2890)) xor (layer1_outputs(507));
    layer2_outputs(331) <= not(layer1_outputs(516));
    layer2_outputs(332) <= (layer1_outputs(3187)) and not (layer1_outputs(4244));
    layer2_outputs(333) <= (layer1_outputs(2701)) and not (layer1_outputs(336));
    layer2_outputs(334) <= layer1_outputs(1033);
    layer2_outputs(335) <= not(layer1_outputs(2777));
    layer2_outputs(336) <= layer1_outputs(980);
    layer2_outputs(337) <= not(layer1_outputs(598));
    layer2_outputs(338) <= layer1_outputs(351);
    layer2_outputs(339) <= not((layer1_outputs(3726)) and (layer1_outputs(4187)));
    layer2_outputs(340) <= not((layer1_outputs(1566)) or (layer1_outputs(2692)));
    layer2_outputs(341) <= '0';
    layer2_outputs(342) <= not(layer1_outputs(3412)) or (layer1_outputs(4927));
    layer2_outputs(343) <= not(layer1_outputs(1720)) or (layer1_outputs(3139));
    layer2_outputs(344) <= not(layer1_outputs(850)) or (layer1_outputs(4422));
    layer2_outputs(345) <= layer1_outputs(4152);
    layer2_outputs(346) <= not((layer1_outputs(3847)) and (layer1_outputs(2331)));
    layer2_outputs(347) <= (layer1_outputs(5100)) and not (layer1_outputs(574));
    layer2_outputs(348) <= not((layer1_outputs(2675)) or (layer1_outputs(4310)));
    layer2_outputs(349) <= layer1_outputs(195);
    layer2_outputs(350) <= (layer1_outputs(307)) xor (layer1_outputs(14));
    layer2_outputs(351) <= (layer1_outputs(2348)) and not (layer1_outputs(1025));
    layer2_outputs(352) <= (layer1_outputs(3715)) or (layer1_outputs(1670));
    layer2_outputs(353) <= (layer1_outputs(3342)) xor (layer1_outputs(1162));
    layer2_outputs(354) <= layer1_outputs(1877);
    layer2_outputs(355) <= not(layer1_outputs(3645));
    layer2_outputs(356) <= layer1_outputs(2913);
    layer2_outputs(357) <= (layer1_outputs(398)) or (layer1_outputs(2614));
    layer2_outputs(358) <= not((layer1_outputs(5106)) or (layer1_outputs(2025)));
    layer2_outputs(359) <= (layer1_outputs(2994)) and not (layer1_outputs(1327));
    layer2_outputs(360) <= (layer1_outputs(1979)) xor (layer1_outputs(443));
    layer2_outputs(361) <= not(layer1_outputs(4841)) or (layer1_outputs(3805));
    layer2_outputs(362) <= not((layer1_outputs(1742)) or (layer1_outputs(3719)));
    layer2_outputs(363) <= (layer1_outputs(4936)) xor (layer1_outputs(2519));
    layer2_outputs(364) <= (layer1_outputs(1616)) or (layer1_outputs(1283));
    layer2_outputs(365) <= layer1_outputs(1109);
    layer2_outputs(366) <= layer1_outputs(531);
    layer2_outputs(367) <= not(layer1_outputs(2480));
    layer2_outputs(368) <= layer1_outputs(470);
    layer2_outputs(369) <= not(layer1_outputs(4914));
    layer2_outputs(370) <= not((layer1_outputs(394)) or (layer1_outputs(2021)));
    layer2_outputs(371) <= layer1_outputs(1344);
    layer2_outputs(372) <= layer1_outputs(4183);
    layer2_outputs(373) <= not(layer1_outputs(1885));
    layer2_outputs(374) <= (layer1_outputs(271)) or (layer1_outputs(3352));
    layer2_outputs(375) <= (layer1_outputs(3733)) and not (layer1_outputs(3951));
    layer2_outputs(376) <= (layer1_outputs(1934)) or (layer1_outputs(2136));
    layer2_outputs(377) <= layer1_outputs(1054);
    layer2_outputs(378) <= not(layer1_outputs(4681));
    layer2_outputs(379) <= not(layer1_outputs(3683)) or (layer1_outputs(208));
    layer2_outputs(380) <= not((layer1_outputs(2414)) or (layer1_outputs(2758)));
    layer2_outputs(381) <= (layer1_outputs(4505)) and (layer1_outputs(2484));
    layer2_outputs(382) <= layer1_outputs(1808);
    layer2_outputs(383) <= not((layer1_outputs(3185)) xor (layer1_outputs(2833)));
    layer2_outputs(384) <= not(layer1_outputs(300));
    layer2_outputs(385) <= (layer1_outputs(2604)) and (layer1_outputs(939));
    layer2_outputs(386) <= not(layer1_outputs(2948));
    layer2_outputs(387) <= layer1_outputs(378);
    layer2_outputs(388) <= not(layer1_outputs(1019));
    layer2_outputs(389) <= (layer1_outputs(1649)) xor (layer1_outputs(165));
    layer2_outputs(390) <= not(layer1_outputs(1165));
    layer2_outputs(391) <= layer1_outputs(2329);
    layer2_outputs(392) <= '0';
    layer2_outputs(393) <= (layer1_outputs(676)) or (layer1_outputs(662));
    layer2_outputs(394) <= (layer1_outputs(2676)) or (layer1_outputs(3443));
    layer2_outputs(395) <= not(layer1_outputs(179)) or (layer1_outputs(1803));
    layer2_outputs(396) <= not((layer1_outputs(796)) and (layer1_outputs(2788)));
    layer2_outputs(397) <= not(layer1_outputs(3073)) or (layer1_outputs(690));
    layer2_outputs(398) <= not(layer1_outputs(4223)) or (layer1_outputs(1875));
    layer2_outputs(399) <= layer1_outputs(2047);
    layer2_outputs(400) <= (layer1_outputs(4670)) and not (layer1_outputs(60));
    layer2_outputs(401) <= not(layer1_outputs(960));
    layer2_outputs(402) <= not((layer1_outputs(3302)) or (layer1_outputs(4451)));
    layer2_outputs(403) <= not(layer1_outputs(5110));
    layer2_outputs(404) <= not(layer1_outputs(4971)) or (layer1_outputs(3365));
    layer2_outputs(405) <= not(layer1_outputs(3436)) or (layer1_outputs(1425));
    layer2_outputs(406) <= (layer1_outputs(3272)) and not (layer1_outputs(4649));
    layer2_outputs(407) <= (layer1_outputs(1971)) and (layer1_outputs(4594));
    layer2_outputs(408) <= layer1_outputs(3347);
    layer2_outputs(409) <= layer1_outputs(2469);
    layer2_outputs(410) <= not(layer1_outputs(3219));
    layer2_outputs(411) <= (layer1_outputs(1803)) or (layer1_outputs(311));
    layer2_outputs(412) <= not(layer1_outputs(697)) or (layer1_outputs(1987));
    layer2_outputs(413) <= not(layer1_outputs(1912)) or (layer1_outputs(4849));
    layer2_outputs(414) <= not(layer1_outputs(2866));
    layer2_outputs(415) <= not(layer1_outputs(1946)) or (layer1_outputs(1074));
    layer2_outputs(416) <= (layer1_outputs(4130)) and (layer1_outputs(950));
    layer2_outputs(417) <= not((layer1_outputs(2946)) xor (layer1_outputs(1470)));
    layer2_outputs(418) <= not((layer1_outputs(505)) or (layer1_outputs(2310)));
    layer2_outputs(419) <= layer1_outputs(3653);
    layer2_outputs(420) <= (layer1_outputs(2982)) or (layer1_outputs(19));
    layer2_outputs(421) <= (layer1_outputs(3023)) and (layer1_outputs(1887));
    layer2_outputs(422) <= layer1_outputs(3838);
    layer2_outputs(423) <= layer1_outputs(4810);
    layer2_outputs(424) <= layer1_outputs(4274);
    layer2_outputs(425) <= layer1_outputs(3264);
    layer2_outputs(426) <= (layer1_outputs(4142)) and (layer1_outputs(4082));
    layer2_outputs(427) <= not(layer1_outputs(4020)) or (layer1_outputs(18));
    layer2_outputs(428) <= not((layer1_outputs(4073)) xor (layer1_outputs(1325)));
    layer2_outputs(429) <= not((layer1_outputs(1906)) and (layer1_outputs(4274)));
    layer2_outputs(430) <= (layer1_outputs(1845)) xor (layer1_outputs(3873));
    layer2_outputs(431) <= not(layer1_outputs(2832)) or (layer1_outputs(4763));
    layer2_outputs(432) <= layer1_outputs(3212);
    layer2_outputs(433) <= not((layer1_outputs(2622)) or (layer1_outputs(3765)));
    layer2_outputs(434) <= (layer1_outputs(611)) and not (layer1_outputs(199));
    layer2_outputs(435) <= (layer1_outputs(1535)) and not (layer1_outputs(3666));
    layer2_outputs(436) <= layer1_outputs(252);
    layer2_outputs(437) <= not(layer1_outputs(4537));
    layer2_outputs(438) <= (layer1_outputs(1400)) and (layer1_outputs(3764));
    layer2_outputs(439) <= not(layer1_outputs(1751));
    layer2_outputs(440) <= not(layer1_outputs(1812));
    layer2_outputs(441) <= (layer1_outputs(2727)) or (layer1_outputs(2940));
    layer2_outputs(442) <= (layer1_outputs(2686)) xor (layer1_outputs(1036));
    layer2_outputs(443) <= not((layer1_outputs(2663)) xor (layer1_outputs(3656)));
    layer2_outputs(444) <= not(layer1_outputs(613));
    layer2_outputs(445) <= layer1_outputs(2629);
    layer2_outputs(446) <= (layer1_outputs(64)) xor (layer1_outputs(3970));
    layer2_outputs(447) <= layer1_outputs(3305);
    layer2_outputs(448) <= layer1_outputs(1198);
    layer2_outputs(449) <= (layer1_outputs(4632)) or (layer1_outputs(4474));
    layer2_outputs(450) <= not(layer1_outputs(269));
    layer2_outputs(451) <= (layer1_outputs(4705)) xor (layer1_outputs(338));
    layer2_outputs(452) <= not(layer1_outputs(12)) or (layer1_outputs(1089));
    layer2_outputs(453) <= '1';
    layer2_outputs(454) <= (layer1_outputs(2796)) and not (layer1_outputs(2050));
    layer2_outputs(455) <= not(layer1_outputs(1659));
    layer2_outputs(456) <= not(layer1_outputs(3135));
    layer2_outputs(457) <= not(layer1_outputs(259));
    layer2_outputs(458) <= (layer1_outputs(3240)) and not (layer1_outputs(3966));
    layer2_outputs(459) <= layer1_outputs(4108);
    layer2_outputs(460) <= not(layer1_outputs(2544));
    layer2_outputs(461) <= layer1_outputs(295);
    layer2_outputs(462) <= not((layer1_outputs(3132)) xor (layer1_outputs(825)));
    layer2_outputs(463) <= (layer1_outputs(1048)) and not (layer1_outputs(46));
    layer2_outputs(464) <= (layer1_outputs(824)) and not (layer1_outputs(2616));
    layer2_outputs(465) <= '0';
    layer2_outputs(466) <= not((layer1_outputs(947)) or (layer1_outputs(3227)));
    layer2_outputs(467) <= (layer1_outputs(786)) xor (layer1_outputs(294));
    layer2_outputs(468) <= not((layer1_outputs(4777)) xor (layer1_outputs(1692)));
    layer2_outputs(469) <= not(layer1_outputs(3357));
    layer2_outputs(470) <= not(layer1_outputs(2747));
    layer2_outputs(471) <= layer1_outputs(2932);
    layer2_outputs(472) <= not((layer1_outputs(2411)) xor (layer1_outputs(1473)));
    layer2_outputs(473) <= (layer1_outputs(3802)) and not (layer1_outputs(1451));
    layer2_outputs(474) <= not(layer1_outputs(474));
    layer2_outputs(475) <= not(layer1_outputs(2749));
    layer2_outputs(476) <= layer1_outputs(3100);
    layer2_outputs(477) <= not(layer1_outputs(3594));
    layer2_outputs(478) <= '1';
    layer2_outputs(479) <= (layer1_outputs(4876)) or (layer1_outputs(30));
    layer2_outputs(480) <= not(layer1_outputs(4346));
    layer2_outputs(481) <= (layer1_outputs(3566)) and not (layer1_outputs(4932));
    layer2_outputs(482) <= not((layer1_outputs(3356)) or (layer1_outputs(4882)));
    layer2_outputs(483) <= not((layer1_outputs(4892)) and (layer1_outputs(43)));
    layer2_outputs(484) <= (layer1_outputs(3580)) and not (layer1_outputs(2192));
    layer2_outputs(485) <= not(layer1_outputs(1672));
    layer2_outputs(486) <= not((layer1_outputs(4537)) and (layer1_outputs(3201)));
    layer2_outputs(487) <= not(layer1_outputs(2924));
    layer2_outputs(488) <= layer1_outputs(903);
    layer2_outputs(489) <= not(layer1_outputs(1428));
    layer2_outputs(490) <= (layer1_outputs(3009)) or (layer1_outputs(4621));
    layer2_outputs(491) <= not((layer1_outputs(217)) and (layer1_outputs(2276)));
    layer2_outputs(492) <= not(layer1_outputs(4249));
    layer2_outputs(493) <= not((layer1_outputs(4208)) and (layer1_outputs(2825)));
    layer2_outputs(494) <= not((layer1_outputs(3894)) xor (layer1_outputs(2915)));
    layer2_outputs(495) <= layer1_outputs(2482);
    layer2_outputs(496) <= not(layer1_outputs(3238));
    layer2_outputs(497) <= layer1_outputs(3886);
    layer2_outputs(498) <= not(layer1_outputs(1518)) or (layer1_outputs(742));
    layer2_outputs(499) <= (layer1_outputs(1701)) or (layer1_outputs(954));
    layer2_outputs(500) <= layer1_outputs(2578);
    layer2_outputs(501) <= not(layer1_outputs(3874));
    layer2_outputs(502) <= (layer1_outputs(2299)) and not (layer1_outputs(4673));
    layer2_outputs(503) <= '1';
    layer2_outputs(504) <= not((layer1_outputs(1458)) and (layer1_outputs(2306)));
    layer2_outputs(505) <= (layer1_outputs(2208)) xor (layer1_outputs(3012));
    layer2_outputs(506) <= not(layer1_outputs(2142));
    layer2_outputs(507) <= not((layer1_outputs(733)) xor (layer1_outputs(3390)));
    layer2_outputs(508) <= not(layer1_outputs(5012));
    layer2_outputs(509) <= layer1_outputs(289);
    layer2_outputs(510) <= not(layer1_outputs(762));
    layer2_outputs(511) <= not((layer1_outputs(3120)) xor (layer1_outputs(2498)));
    layer2_outputs(512) <= layer1_outputs(3667);
    layer2_outputs(513) <= not(layer1_outputs(372));
    layer2_outputs(514) <= layer1_outputs(957);
    layer2_outputs(515) <= layer1_outputs(10);
    layer2_outputs(516) <= (layer1_outputs(2469)) xor (layer1_outputs(1179));
    layer2_outputs(517) <= (layer1_outputs(271)) and (layer1_outputs(1073));
    layer2_outputs(518) <= not(layer1_outputs(2275)) or (layer1_outputs(3104));
    layer2_outputs(519) <= (layer1_outputs(4622)) and (layer1_outputs(3241));
    layer2_outputs(520) <= not(layer1_outputs(1113)) or (layer1_outputs(191));
    layer2_outputs(521) <= not(layer1_outputs(3900));
    layer2_outputs(522) <= layer1_outputs(988);
    layer2_outputs(523) <= not(layer1_outputs(4588)) or (layer1_outputs(2552));
    layer2_outputs(524) <= not(layer1_outputs(2789));
    layer2_outputs(525) <= not(layer1_outputs(3313));
    layer2_outputs(526) <= not(layer1_outputs(2516));
    layer2_outputs(527) <= not(layer1_outputs(2289)) or (layer1_outputs(3442));
    layer2_outputs(528) <= layer1_outputs(545);
    layer2_outputs(529) <= not(layer1_outputs(827));
    layer2_outputs(530) <= (layer1_outputs(2362)) and (layer1_outputs(2754));
    layer2_outputs(531) <= not(layer1_outputs(793));
    layer2_outputs(532) <= not(layer1_outputs(2172));
    layer2_outputs(533) <= layer1_outputs(5111);
    layer2_outputs(534) <= not(layer1_outputs(4107));
    layer2_outputs(535) <= layer1_outputs(4912);
    layer2_outputs(536) <= (layer1_outputs(2369)) and not (layer1_outputs(4731));
    layer2_outputs(537) <= layer1_outputs(3563);
    layer2_outputs(538) <= not(layer1_outputs(365));
    layer2_outputs(539) <= not(layer1_outputs(5038));
    layer2_outputs(540) <= not((layer1_outputs(1330)) or (layer1_outputs(2703)));
    layer2_outputs(541) <= '0';
    layer2_outputs(542) <= not(layer1_outputs(2619));
    layer2_outputs(543) <= not(layer1_outputs(1256));
    layer2_outputs(544) <= layer1_outputs(2536);
    layer2_outputs(545) <= (layer1_outputs(213)) and not (layer1_outputs(1735));
    layer2_outputs(546) <= not((layer1_outputs(3270)) and (layer1_outputs(2250)));
    layer2_outputs(547) <= not(layer1_outputs(3705));
    layer2_outputs(548) <= not(layer1_outputs(3246));
    layer2_outputs(549) <= not(layer1_outputs(2200)) or (layer1_outputs(4111));
    layer2_outputs(550) <= layer1_outputs(2002);
    layer2_outputs(551) <= not(layer1_outputs(1519));
    layer2_outputs(552) <= not(layer1_outputs(3563));
    layer2_outputs(553) <= layer1_outputs(1171);
    layer2_outputs(554) <= layer1_outputs(603);
    layer2_outputs(555) <= layer1_outputs(2065);
    layer2_outputs(556) <= not(layer1_outputs(2756)) or (layer1_outputs(3864));
    layer2_outputs(557) <= not((layer1_outputs(4066)) xor (layer1_outputs(2161)));
    layer2_outputs(558) <= not(layer1_outputs(3435)) or (layer1_outputs(1171));
    layer2_outputs(559) <= layer1_outputs(4545);
    layer2_outputs(560) <= (layer1_outputs(4673)) and (layer1_outputs(621));
    layer2_outputs(561) <= layer1_outputs(1871);
    layer2_outputs(562) <= not(layer1_outputs(4041)) or (layer1_outputs(950));
    layer2_outputs(563) <= (layer1_outputs(629)) or (layer1_outputs(3536));
    layer2_outputs(564) <= not((layer1_outputs(958)) xor (layer1_outputs(4812)));
    layer2_outputs(565) <= not(layer1_outputs(4394));
    layer2_outputs(566) <= not(layer1_outputs(719)) or (layer1_outputs(3967));
    layer2_outputs(567) <= not(layer1_outputs(3643));
    layer2_outputs(568) <= not((layer1_outputs(1667)) xor (layer1_outputs(4822)));
    layer2_outputs(569) <= (layer1_outputs(4652)) and not (layer1_outputs(3995));
    layer2_outputs(570) <= (layer1_outputs(2419)) and not (layer1_outputs(2858));
    layer2_outputs(571) <= (layer1_outputs(3072)) or (layer1_outputs(2352));
    layer2_outputs(572) <= layer1_outputs(4137);
    layer2_outputs(573) <= (layer1_outputs(2677)) and not (layer1_outputs(2051));
    layer2_outputs(574) <= layer1_outputs(4172);
    layer2_outputs(575) <= (layer1_outputs(3261)) and not (layer1_outputs(513));
    layer2_outputs(576) <= not((layer1_outputs(1213)) and (layer1_outputs(1920)));
    layer2_outputs(577) <= not(layer1_outputs(719));
    layer2_outputs(578) <= not(layer1_outputs(3099));
    layer2_outputs(579) <= not((layer1_outputs(2004)) or (layer1_outputs(1326)));
    layer2_outputs(580) <= not((layer1_outputs(1238)) xor (layer1_outputs(994)));
    layer2_outputs(581) <= not(layer1_outputs(1258));
    layer2_outputs(582) <= not(layer1_outputs(648));
    layer2_outputs(583) <= layer1_outputs(3617);
    layer2_outputs(584) <= not((layer1_outputs(765)) or (layer1_outputs(2965)));
    layer2_outputs(585) <= layer1_outputs(2451);
    layer2_outputs(586) <= not(layer1_outputs(4133));
    layer2_outputs(587) <= not((layer1_outputs(4733)) or (layer1_outputs(251)));
    layer2_outputs(588) <= not(layer1_outputs(3634));
    layer2_outputs(589) <= not(layer1_outputs(4379)) or (layer1_outputs(4398));
    layer2_outputs(590) <= (layer1_outputs(668)) and (layer1_outputs(991));
    layer2_outputs(591) <= layer1_outputs(4864);
    layer2_outputs(592) <= not(layer1_outputs(2454));
    layer2_outputs(593) <= layer1_outputs(1659);
    layer2_outputs(594) <= (layer1_outputs(3141)) and (layer1_outputs(3264));
    layer2_outputs(595) <= (layer1_outputs(2464)) and (layer1_outputs(60));
    layer2_outputs(596) <= (layer1_outputs(302)) or (layer1_outputs(1135));
    layer2_outputs(597) <= not((layer1_outputs(1723)) and (layer1_outputs(4078)));
    layer2_outputs(598) <= (layer1_outputs(1520)) xor (layer1_outputs(1049));
    layer2_outputs(599) <= (layer1_outputs(3020)) and (layer1_outputs(3722));
    layer2_outputs(600) <= (layer1_outputs(3784)) or (layer1_outputs(203));
    layer2_outputs(601) <= layer1_outputs(4519);
    layer2_outputs(602) <= (layer1_outputs(2992)) and not (layer1_outputs(2772));
    layer2_outputs(603) <= not((layer1_outputs(5011)) xor (layer1_outputs(1213)));
    layer2_outputs(604) <= not(layer1_outputs(52)) or (layer1_outputs(597));
    layer2_outputs(605) <= (layer1_outputs(2654)) and (layer1_outputs(3455));
    layer2_outputs(606) <= (layer1_outputs(3692)) and not (layer1_outputs(4582));
    layer2_outputs(607) <= layer1_outputs(3153);
    layer2_outputs(608) <= not(layer1_outputs(830));
    layer2_outputs(609) <= not(layer1_outputs(2792));
    layer2_outputs(610) <= layer1_outputs(1824);
    layer2_outputs(611) <= (layer1_outputs(519)) and not (layer1_outputs(1193));
    layer2_outputs(612) <= (layer1_outputs(2290)) and (layer1_outputs(3893));
    layer2_outputs(613) <= layer1_outputs(2839);
    layer2_outputs(614) <= (layer1_outputs(1921)) and not (layer1_outputs(3247));
    layer2_outputs(615) <= (layer1_outputs(4236)) and (layer1_outputs(4126));
    layer2_outputs(616) <= not(layer1_outputs(1278));
    layer2_outputs(617) <= not(layer1_outputs(473));
    layer2_outputs(618) <= not(layer1_outputs(2332));
    layer2_outputs(619) <= (layer1_outputs(1024)) or (layer1_outputs(4790));
    layer2_outputs(620) <= layer1_outputs(1864);
    layer2_outputs(621) <= (layer1_outputs(2024)) xor (layer1_outputs(1467));
    layer2_outputs(622) <= not(layer1_outputs(2776));
    layer2_outputs(623) <= (layer1_outputs(4661)) or (layer1_outputs(365));
    layer2_outputs(624) <= not(layer1_outputs(2761));
    layer2_outputs(625) <= layer1_outputs(335);
    layer2_outputs(626) <= '1';
    layer2_outputs(627) <= layer1_outputs(1581);
    layer2_outputs(628) <= layer1_outputs(4938);
    layer2_outputs(629) <= not((layer1_outputs(1307)) xor (layer1_outputs(47)));
    layer2_outputs(630) <= (layer1_outputs(2903)) and (layer1_outputs(4700));
    layer2_outputs(631) <= layer1_outputs(4786);
    layer2_outputs(632) <= (layer1_outputs(4033)) and not (layer1_outputs(4476));
    layer2_outputs(633) <= (layer1_outputs(4042)) and not (layer1_outputs(901));
    layer2_outputs(634) <= layer1_outputs(2494);
    layer2_outputs(635) <= layer1_outputs(438);
    layer2_outputs(636) <= not((layer1_outputs(2616)) or (layer1_outputs(3681)));
    layer2_outputs(637) <= not(layer1_outputs(3543));
    layer2_outputs(638) <= (layer1_outputs(3918)) and (layer1_outputs(4160));
    layer2_outputs(639) <= not(layer1_outputs(257));
    layer2_outputs(640) <= layer1_outputs(1063);
    layer2_outputs(641) <= not(layer1_outputs(3696)) or (layer1_outputs(1723));
    layer2_outputs(642) <= not((layer1_outputs(400)) and (layer1_outputs(3070)));
    layer2_outputs(643) <= (layer1_outputs(1604)) or (layer1_outputs(1691));
    layer2_outputs(644) <= not(layer1_outputs(3199));
    layer2_outputs(645) <= not(layer1_outputs(4768));
    layer2_outputs(646) <= not((layer1_outputs(3124)) or (layer1_outputs(1404)));
    layer2_outputs(647) <= not(layer1_outputs(797)) or (layer1_outputs(4521));
    layer2_outputs(648) <= not(layer1_outputs(2909));
    layer2_outputs(649) <= not(layer1_outputs(3453));
    layer2_outputs(650) <= (layer1_outputs(823)) and not (layer1_outputs(2175));
    layer2_outputs(651) <= not(layer1_outputs(1729));
    layer2_outputs(652) <= (layer1_outputs(502)) or (layer1_outputs(4117));
    layer2_outputs(653) <= layer1_outputs(2117);
    layer2_outputs(654) <= layer1_outputs(1237);
    layer2_outputs(655) <= (layer1_outputs(997)) and not (layer1_outputs(1070));
    layer2_outputs(656) <= not(layer1_outputs(501));
    layer2_outputs(657) <= layer1_outputs(4919);
    layer2_outputs(658) <= layer1_outputs(4796);
    layer2_outputs(659) <= layer1_outputs(4966);
    layer2_outputs(660) <= not((layer1_outputs(1994)) and (layer1_outputs(4448)));
    layer2_outputs(661) <= layer1_outputs(3109);
    layer2_outputs(662) <= not(layer1_outputs(2651));
    layer2_outputs(663) <= (layer1_outputs(838)) and not (layer1_outputs(4150));
    layer2_outputs(664) <= (layer1_outputs(2381)) or (layer1_outputs(4016));
    layer2_outputs(665) <= not(layer1_outputs(1523));
    layer2_outputs(666) <= (layer1_outputs(3012)) and not (layer1_outputs(429));
    layer2_outputs(667) <= (layer1_outputs(4605)) and not (layer1_outputs(4715));
    layer2_outputs(668) <= layer1_outputs(280);
    layer2_outputs(669) <= not((layer1_outputs(993)) or (layer1_outputs(893)));
    layer2_outputs(670) <= layer1_outputs(2350);
    layer2_outputs(671) <= layer1_outputs(1053);
    layer2_outputs(672) <= not(layer1_outputs(351));
    layer2_outputs(673) <= layer1_outputs(2128);
    layer2_outputs(674) <= not((layer1_outputs(3019)) or (layer1_outputs(1941)));
    layer2_outputs(675) <= layer1_outputs(995);
    layer2_outputs(676) <= not(layer1_outputs(2821));
    layer2_outputs(677) <= not(layer1_outputs(4467));
    layer2_outputs(678) <= not(layer1_outputs(4018));
    layer2_outputs(679) <= layer1_outputs(3502);
    layer2_outputs(680) <= layer1_outputs(4309);
    layer2_outputs(681) <= not((layer1_outputs(702)) or (layer1_outputs(3060)));
    layer2_outputs(682) <= not(layer1_outputs(4028));
    layer2_outputs(683) <= layer1_outputs(4564);
    layer2_outputs(684) <= not((layer1_outputs(581)) xor (layer1_outputs(921)));
    layer2_outputs(685) <= not((layer1_outputs(3117)) and (layer1_outputs(3223)));
    layer2_outputs(686) <= (layer1_outputs(84)) and not (layer1_outputs(1821));
    layer2_outputs(687) <= not(layer1_outputs(2345));
    layer2_outputs(688) <= layer1_outputs(3724);
    layer2_outputs(689) <= not(layer1_outputs(1480)) or (layer1_outputs(4494));
    layer2_outputs(690) <= layer1_outputs(37);
    layer2_outputs(691) <= not(layer1_outputs(4045));
    layer2_outputs(692) <= not(layer1_outputs(2045)) or (layer1_outputs(3396));
    layer2_outputs(693) <= not((layer1_outputs(1129)) xor (layer1_outputs(4767)));
    layer2_outputs(694) <= (layer1_outputs(1856)) and not (layer1_outputs(2465));
    layer2_outputs(695) <= (layer1_outputs(4676)) xor (layer1_outputs(3968));
    layer2_outputs(696) <= layer1_outputs(2518);
    layer2_outputs(697) <= not(layer1_outputs(1239));
    layer2_outputs(698) <= not(layer1_outputs(3103)) or (layer1_outputs(2819));
    layer2_outputs(699) <= not((layer1_outputs(4933)) xor (layer1_outputs(2206)));
    layer2_outputs(700) <= (layer1_outputs(2213)) and not (layer1_outputs(3165));
    layer2_outputs(701) <= (layer1_outputs(198)) or (layer1_outputs(94));
    layer2_outputs(702) <= not(layer1_outputs(2473));
    layer2_outputs(703) <= layer1_outputs(2755);
    layer2_outputs(704) <= not((layer1_outputs(4994)) or (layer1_outputs(4071)));
    layer2_outputs(705) <= not(layer1_outputs(1787)) or (layer1_outputs(957));
    layer2_outputs(706) <= not((layer1_outputs(2077)) xor (layer1_outputs(112)));
    layer2_outputs(707) <= layer1_outputs(4250);
    layer2_outputs(708) <= not(layer1_outputs(3248)) or (layer1_outputs(2581));
    layer2_outputs(709) <= (layer1_outputs(1808)) and not (layer1_outputs(2979));
    layer2_outputs(710) <= layer1_outputs(1727);
    layer2_outputs(711) <= not(layer1_outputs(1333));
    layer2_outputs(712) <= not(layer1_outputs(4650));
    layer2_outputs(713) <= not((layer1_outputs(1732)) xor (layer1_outputs(1925)));
    layer2_outputs(714) <= layer1_outputs(2449);
    layer2_outputs(715) <= not(layer1_outputs(4426));
    layer2_outputs(716) <= layer1_outputs(1990);
    layer2_outputs(717) <= not(layer1_outputs(3892));
    layer2_outputs(718) <= not((layer1_outputs(5062)) and (layer1_outputs(2219)));
    layer2_outputs(719) <= (layer1_outputs(4655)) or (layer1_outputs(5037));
    layer2_outputs(720) <= not(layer1_outputs(4973));
    layer2_outputs(721) <= layer1_outputs(4628);
    layer2_outputs(722) <= layer1_outputs(4152);
    layer2_outputs(723) <= (layer1_outputs(4864)) and (layer1_outputs(1416));
    layer2_outputs(724) <= not(layer1_outputs(2603));
    layer2_outputs(725) <= (layer1_outputs(4524)) and not (layer1_outputs(776));
    layer2_outputs(726) <= (layer1_outputs(1133)) xor (layer1_outputs(4115));
    layer2_outputs(727) <= (layer1_outputs(4348)) or (layer1_outputs(4520));
    layer2_outputs(728) <= not(layer1_outputs(3300));
    layer2_outputs(729) <= (layer1_outputs(1204)) and not (layer1_outputs(2504));
    layer2_outputs(730) <= layer1_outputs(890);
    layer2_outputs(731) <= not(layer1_outputs(548));
    layer2_outputs(732) <= (layer1_outputs(15)) and not (layer1_outputs(3028));
    layer2_outputs(733) <= not(layer1_outputs(2277));
    layer2_outputs(734) <= (layer1_outputs(4686)) and not (layer1_outputs(858));
    layer2_outputs(735) <= (layer1_outputs(2594)) and not (layer1_outputs(3131));
    layer2_outputs(736) <= not((layer1_outputs(4656)) and (layer1_outputs(2980)));
    layer2_outputs(737) <= (layer1_outputs(4580)) and not (layer1_outputs(2976));
    layer2_outputs(738) <= (layer1_outputs(2700)) and not (layer1_outputs(2324));
    layer2_outputs(739) <= not(layer1_outputs(3546));
    layer2_outputs(740) <= '0';
    layer2_outputs(741) <= (layer1_outputs(3398)) or (layer1_outputs(567));
    layer2_outputs(742) <= (layer1_outputs(961)) and not (layer1_outputs(4597));
    layer2_outputs(743) <= (layer1_outputs(3326)) and not (layer1_outputs(4147));
    layer2_outputs(744) <= layer1_outputs(2220);
    layer2_outputs(745) <= not((layer1_outputs(973)) or (layer1_outputs(4051)));
    layer2_outputs(746) <= not(layer1_outputs(565));
    layer2_outputs(747) <= layer1_outputs(1846);
    layer2_outputs(748) <= (layer1_outputs(2744)) xor (layer1_outputs(3849));
    layer2_outputs(749) <= layer1_outputs(700);
    layer2_outputs(750) <= layer1_outputs(526);
    layer2_outputs(751) <= not((layer1_outputs(4883)) xor (layer1_outputs(2944)));
    layer2_outputs(752) <= not((layer1_outputs(2668)) xor (layer1_outputs(255)));
    layer2_outputs(753) <= (layer1_outputs(162)) and not (layer1_outputs(4007));
    layer2_outputs(754) <= (layer1_outputs(3768)) and (layer1_outputs(4611));
    layer2_outputs(755) <= not(layer1_outputs(1032));
    layer2_outputs(756) <= not(layer1_outputs(216));
    layer2_outputs(757) <= '1';
    layer2_outputs(758) <= (layer1_outputs(1404)) xor (layer1_outputs(197));
    layer2_outputs(759) <= (layer1_outputs(2355)) or (layer1_outputs(3573));
    layer2_outputs(760) <= not(layer1_outputs(2116)) or (layer1_outputs(3066));
    layer2_outputs(761) <= not((layer1_outputs(331)) xor (layer1_outputs(922)));
    layer2_outputs(762) <= (layer1_outputs(316)) and (layer1_outputs(130));
    layer2_outputs(763) <= (layer1_outputs(2023)) and (layer1_outputs(970));
    layer2_outputs(764) <= (layer1_outputs(1286)) and not (layer1_outputs(3610));
    layer2_outputs(765) <= not(layer1_outputs(68)) or (layer1_outputs(2595));
    layer2_outputs(766) <= not(layer1_outputs(217)) or (layer1_outputs(5090));
    layer2_outputs(767) <= layer1_outputs(2800);
    layer2_outputs(768) <= (layer1_outputs(981)) xor (layer1_outputs(1700));
    layer2_outputs(769) <= layer1_outputs(4114);
    layer2_outputs(770) <= (layer1_outputs(1439)) xor (layer1_outputs(4088));
    layer2_outputs(771) <= (layer1_outputs(1721)) or (layer1_outputs(1029));
    layer2_outputs(772) <= (layer1_outputs(3964)) xor (layer1_outputs(3806));
    layer2_outputs(773) <= not(layer1_outputs(2934)) or (layer1_outputs(1126));
    layer2_outputs(774) <= layer1_outputs(2562);
    layer2_outputs(775) <= layer1_outputs(5018);
    layer2_outputs(776) <= (layer1_outputs(3503)) and not (layer1_outputs(1415));
    layer2_outputs(777) <= (layer1_outputs(1645)) and (layer1_outputs(907));
    layer2_outputs(778) <= not((layer1_outputs(3400)) xor (layer1_outputs(2902)));
    layer2_outputs(779) <= layer1_outputs(1429);
    layer2_outputs(780) <= not((layer1_outputs(4128)) xor (layer1_outputs(1799)));
    layer2_outputs(781) <= layer1_outputs(4851);
    layer2_outputs(782) <= not(layer1_outputs(3583));
    layer2_outputs(783) <= not(layer1_outputs(3215)) or (layer1_outputs(799));
    layer2_outputs(784) <= not(layer1_outputs(2378));
    layer2_outputs(785) <= '1';
    layer2_outputs(786) <= (layer1_outputs(844)) and (layer1_outputs(3451));
    layer2_outputs(787) <= layer1_outputs(2943);
    layer2_outputs(788) <= (layer1_outputs(4909)) xor (layer1_outputs(3263));
    layer2_outputs(789) <= layer1_outputs(3821);
    layer2_outputs(790) <= not(layer1_outputs(2406));
    layer2_outputs(791) <= not((layer1_outputs(1426)) and (layer1_outputs(2094)));
    layer2_outputs(792) <= layer1_outputs(2347);
    layer2_outputs(793) <= not(layer1_outputs(1762));
    layer2_outputs(794) <= not(layer1_outputs(1062));
    layer2_outputs(795) <= (layer1_outputs(804)) and not (layer1_outputs(2814));
    layer2_outputs(796) <= (layer1_outputs(189)) or (layer1_outputs(4312));
    layer2_outputs(797) <= layer1_outputs(3410);
    layer2_outputs(798) <= not(layer1_outputs(2579));
    layer2_outputs(799) <= layer1_outputs(2090);
    layer2_outputs(800) <= layer1_outputs(1445);
    layer2_outputs(801) <= layer1_outputs(3308);
    layer2_outputs(802) <= not(layer1_outputs(91));
    layer2_outputs(803) <= (layer1_outputs(82)) and (layer1_outputs(3664));
    layer2_outputs(804) <= not((layer1_outputs(1129)) xor (layer1_outputs(2814)));
    layer2_outputs(805) <= layer1_outputs(1204);
    layer2_outputs(806) <= not(layer1_outputs(3001)) or (layer1_outputs(4035));
    layer2_outputs(807) <= layer1_outputs(3516);
    layer2_outputs(808) <= layer1_outputs(1843);
    layer2_outputs(809) <= not(layer1_outputs(1838)) or (layer1_outputs(4899));
    layer2_outputs(810) <= (layer1_outputs(2541)) and (layer1_outputs(2562));
    layer2_outputs(811) <= not(layer1_outputs(2338));
    layer2_outputs(812) <= layer1_outputs(1338);
    layer2_outputs(813) <= not(layer1_outputs(4854)) or (layer1_outputs(1395));
    layer2_outputs(814) <= layer1_outputs(3482);
    layer2_outputs(815) <= not((layer1_outputs(3029)) and (layer1_outputs(3807)));
    layer2_outputs(816) <= not(layer1_outputs(4860));
    layer2_outputs(817) <= not(layer1_outputs(2839));
    layer2_outputs(818) <= not((layer1_outputs(4406)) or (layer1_outputs(1508)));
    layer2_outputs(819) <= (layer1_outputs(3721)) xor (layer1_outputs(2611));
    layer2_outputs(820) <= not(layer1_outputs(2908));
    layer2_outputs(821) <= layer1_outputs(720);
    layer2_outputs(822) <= (layer1_outputs(4612)) or (layer1_outputs(2753));
    layer2_outputs(823) <= (layer1_outputs(891)) and (layer1_outputs(4363));
    layer2_outputs(824) <= layer1_outputs(290);
    layer2_outputs(825) <= not(layer1_outputs(646));
    layer2_outputs(826) <= not(layer1_outputs(237));
    layer2_outputs(827) <= layer1_outputs(3055);
    layer2_outputs(828) <= layer1_outputs(4037);
    layer2_outputs(829) <= layer1_outputs(1888);
    layer2_outputs(830) <= not(layer1_outputs(4451));
    layer2_outputs(831) <= (layer1_outputs(4667)) or (layer1_outputs(2322));
    layer2_outputs(832) <= layer1_outputs(458);
    layer2_outputs(833) <= not(layer1_outputs(340));
    layer2_outputs(834) <= layer1_outputs(458);
    layer2_outputs(835) <= not(layer1_outputs(262));
    layer2_outputs(836) <= (layer1_outputs(4178)) xor (layer1_outputs(864));
    layer2_outputs(837) <= not(layer1_outputs(747));
    layer2_outputs(838) <= (layer1_outputs(3811)) and not (layer1_outputs(2670));
    layer2_outputs(839) <= not(layer1_outputs(2445));
    layer2_outputs(840) <= (layer1_outputs(2320)) xor (layer1_outputs(777));
    layer2_outputs(841) <= layer1_outputs(4550);
    layer2_outputs(842) <= (layer1_outputs(4063)) or (layer1_outputs(2303));
    layer2_outputs(843) <= (layer1_outputs(190)) and (layer1_outputs(3662));
    layer2_outputs(844) <= layer1_outputs(2162);
    layer2_outputs(845) <= (layer1_outputs(3211)) xor (layer1_outputs(2951));
    layer2_outputs(846) <= (layer1_outputs(483)) and not (layer1_outputs(2809));
    layer2_outputs(847) <= layer1_outputs(1385);
    layer2_outputs(848) <= not((layer1_outputs(3962)) or (layer1_outputs(1405)));
    layer2_outputs(849) <= layer1_outputs(1582);
    layer2_outputs(850) <= (layer1_outputs(716)) and not (layer1_outputs(1609));
    layer2_outputs(851) <= not(layer1_outputs(1795));
    layer2_outputs(852) <= not(layer1_outputs(2166));
    layer2_outputs(853) <= not(layer1_outputs(2936)) or (layer1_outputs(3719));
    layer2_outputs(854) <= not(layer1_outputs(4880));
    layer2_outputs(855) <= (layer1_outputs(2736)) xor (layer1_outputs(626));
    layer2_outputs(856) <= not(layer1_outputs(1804)) or (layer1_outputs(2774));
    layer2_outputs(857) <= not(layer1_outputs(1078)) or (layer1_outputs(569));
    layer2_outputs(858) <= not(layer1_outputs(4416)) or (layer1_outputs(1884));
    layer2_outputs(859) <= layer1_outputs(3776);
    layer2_outputs(860) <= layer1_outputs(3528);
    layer2_outputs(861) <= not(layer1_outputs(4201));
    layer2_outputs(862) <= (layer1_outputs(3240)) and (layer1_outputs(4637));
    layer2_outputs(863) <= '0';
    layer2_outputs(864) <= not((layer1_outputs(3288)) xor (layer1_outputs(3070)));
    layer2_outputs(865) <= layer1_outputs(3690);
    layer2_outputs(866) <= not(layer1_outputs(4355));
    layer2_outputs(867) <= not((layer1_outputs(3386)) or (layer1_outputs(3587)));
    layer2_outputs(868) <= not((layer1_outputs(4095)) or (layer1_outputs(204)));
    layer2_outputs(869) <= not(layer1_outputs(2028));
    layer2_outputs(870) <= not(layer1_outputs(2710));
    layer2_outputs(871) <= not(layer1_outputs(1103)) or (layer1_outputs(5004));
    layer2_outputs(872) <= layer1_outputs(2664);
    layer2_outputs(873) <= not(layer1_outputs(920));
    layer2_outputs(874) <= layer1_outputs(3407);
    layer2_outputs(875) <= '0';
    layer2_outputs(876) <= layer1_outputs(3671);
    layer2_outputs(877) <= layer1_outputs(181);
    layer2_outputs(878) <= layer1_outputs(3295);
    layer2_outputs(879) <= '0';
    layer2_outputs(880) <= layer1_outputs(3136);
    layer2_outputs(881) <= not(layer1_outputs(4601)) or (layer1_outputs(27));
    layer2_outputs(882) <= (layer1_outputs(2063)) and not (layer1_outputs(4153));
    layer2_outputs(883) <= '0';
    layer2_outputs(884) <= not((layer1_outputs(2180)) xor (layer1_outputs(1317)));
    layer2_outputs(885) <= (layer1_outputs(2491)) or (layer1_outputs(279));
    layer2_outputs(886) <= (layer1_outputs(3054)) and (layer1_outputs(570));
    layer2_outputs(887) <= layer1_outputs(1697);
    layer2_outputs(888) <= (layer1_outputs(4046)) and not (layer1_outputs(3505));
    layer2_outputs(889) <= not(layer1_outputs(400));
    layer2_outputs(890) <= (layer1_outputs(3777)) and not (layer1_outputs(393));
    layer2_outputs(891) <= not(layer1_outputs(4950)) or (layer1_outputs(3134));
    layer2_outputs(892) <= (layer1_outputs(3037)) and not (layer1_outputs(352));
    layer2_outputs(893) <= layer1_outputs(3479);
    layer2_outputs(894) <= not((layer1_outputs(1255)) or (layer1_outputs(5096)));
    layer2_outputs(895) <= layer1_outputs(3429);
    layer2_outputs(896) <= layer1_outputs(1660);
    layer2_outputs(897) <= not(layer1_outputs(3490));
    layer2_outputs(898) <= (layer1_outputs(322)) and (layer1_outputs(2656));
    layer2_outputs(899) <= (layer1_outputs(3905)) and not (layer1_outputs(2128));
    layer2_outputs(900) <= not((layer1_outputs(2877)) and (layer1_outputs(2322)));
    layer2_outputs(901) <= not(layer1_outputs(63));
    layer2_outputs(902) <= not(layer1_outputs(4284));
    layer2_outputs(903) <= layer1_outputs(3623);
    layer2_outputs(904) <= not(layer1_outputs(2341));
    layer2_outputs(905) <= layer1_outputs(2398);
    layer2_outputs(906) <= layer1_outputs(1299);
    layer2_outputs(907) <= not((layer1_outputs(2732)) xor (layer1_outputs(2354)));
    layer2_outputs(908) <= (layer1_outputs(1944)) and not (layer1_outputs(3929));
    layer2_outputs(909) <= (layer1_outputs(4876)) and (layer1_outputs(4581));
    layer2_outputs(910) <= layer1_outputs(3268);
    layer2_outputs(911) <= '0';
    layer2_outputs(912) <= (layer1_outputs(1615)) and not (layer1_outputs(4373));
    layer2_outputs(913) <= layer1_outputs(3999);
    layer2_outputs(914) <= layer1_outputs(4089);
    layer2_outputs(915) <= not(layer1_outputs(3304)) or (layer1_outputs(5104));
    layer2_outputs(916) <= (layer1_outputs(266)) xor (layer1_outputs(2643));
    layer2_outputs(917) <= not(layer1_outputs(2657));
    layer2_outputs(918) <= layer1_outputs(5006);
    layer2_outputs(919) <= (layer1_outputs(1985)) xor (layer1_outputs(3242));
    layer2_outputs(920) <= not(layer1_outputs(1348));
    layer2_outputs(921) <= (layer1_outputs(3435)) and not (layer1_outputs(5119));
    layer2_outputs(922) <= not((layer1_outputs(629)) or (layer1_outputs(2495)));
    layer2_outputs(923) <= not(layer1_outputs(2705)) or (layer1_outputs(4096));
    layer2_outputs(924) <= not(layer1_outputs(4300));
    layer2_outputs(925) <= not(layer1_outputs(4746));
    layer2_outputs(926) <= layer1_outputs(1242);
    layer2_outputs(927) <= not(layer1_outputs(4052));
    layer2_outputs(928) <= (layer1_outputs(2215)) and not (layer1_outputs(3802));
    layer2_outputs(929) <= not(layer1_outputs(4760));
    layer2_outputs(930) <= (layer1_outputs(3613)) or (layer1_outputs(1261));
    layer2_outputs(931) <= not(layer1_outputs(1753)) or (layer1_outputs(1731));
    layer2_outputs(932) <= not(layer1_outputs(1281)) or (layer1_outputs(2142));
    layer2_outputs(933) <= not(layer1_outputs(2171)) or (layer1_outputs(2960));
    layer2_outputs(934) <= layer1_outputs(2425);
    layer2_outputs(935) <= (layer1_outputs(2401)) xor (layer1_outputs(2280));
    layer2_outputs(936) <= not(layer1_outputs(2408));
    layer2_outputs(937) <= not(layer1_outputs(1819));
    layer2_outputs(938) <= not(layer1_outputs(3604)) or (layer1_outputs(4837));
    layer2_outputs(939) <= not(layer1_outputs(1310));
    layer2_outputs(940) <= not(layer1_outputs(4091));
    layer2_outputs(941) <= not(layer1_outputs(1857));
    layer2_outputs(942) <= layer1_outputs(3417);
    layer2_outputs(943) <= (layer1_outputs(2043)) xor (layer1_outputs(1736));
    layer2_outputs(944) <= not(layer1_outputs(97));
    layer2_outputs(945) <= (layer1_outputs(4848)) and not (layer1_outputs(2883));
    layer2_outputs(946) <= layer1_outputs(1555);
    layer2_outputs(947) <= (layer1_outputs(152)) or (layer1_outputs(754));
    layer2_outputs(948) <= (layer1_outputs(878)) xor (layer1_outputs(1714));
    layer2_outputs(949) <= not(layer1_outputs(4526));
    layer2_outputs(950) <= (layer1_outputs(4828)) and not (layer1_outputs(4317));
    layer2_outputs(951) <= not(layer1_outputs(1844)) or (layer1_outputs(4985));
    layer2_outputs(952) <= not((layer1_outputs(4380)) xor (layer1_outputs(618)));
    layer2_outputs(953) <= not(layer1_outputs(3757));
    layer2_outputs(954) <= not((layer1_outputs(3774)) and (layer1_outputs(151)));
    layer2_outputs(955) <= layer1_outputs(2872);
    layer2_outputs(956) <= layer1_outputs(1538);
    layer2_outputs(957) <= not(layer1_outputs(1709));
    layer2_outputs(958) <= not(layer1_outputs(2658));
    layer2_outputs(959) <= (layer1_outputs(2426)) and (layer1_outputs(4129));
    layer2_outputs(960) <= not(layer1_outputs(3496));
    layer2_outputs(961) <= (layer1_outputs(823)) and not (layer1_outputs(5117));
    layer2_outputs(962) <= layer1_outputs(1911);
    layer2_outputs(963) <= layer1_outputs(4382);
    layer2_outputs(964) <= layer1_outputs(3526);
    layer2_outputs(965) <= (layer1_outputs(3716)) and (layer1_outputs(3660));
    layer2_outputs(966) <= not((layer1_outputs(994)) or (layer1_outputs(4510)));
    layer2_outputs(967) <= (layer1_outputs(283)) and not (layer1_outputs(1531));
    layer2_outputs(968) <= (layer1_outputs(1599)) or (layer1_outputs(4304));
    layer2_outputs(969) <= not(layer1_outputs(4101));
    layer2_outputs(970) <= layer1_outputs(1601);
    layer2_outputs(971) <= not(layer1_outputs(3183));
    layer2_outputs(972) <= layer1_outputs(3335);
    layer2_outputs(973) <= '0';
    layer2_outputs(974) <= layer1_outputs(4472);
    layer2_outputs(975) <= (layer1_outputs(853)) and not (layer1_outputs(3175));
    layer2_outputs(976) <= layer1_outputs(4480);
    layer2_outputs(977) <= not(layer1_outputs(1044));
    layer2_outputs(978) <= not(layer1_outputs(79)) or (layer1_outputs(3662));
    layer2_outputs(979) <= not(layer1_outputs(4047));
    layer2_outputs(980) <= not(layer1_outputs(4738)) or (layer1_outputs(2277));
    layer2_outputs(981) <= not(layer1_outputs(4224)) or (layer1_outputs(3049));
    layer2_outputs(982) <= layer1_outputs(684);
    layer2_outputs(983) <= not(layer1_outputs(2989));
    layer2_outputs(984) <= not((layer1_outputs(3293)) or (layer1_outputs(5117)));
    layer2_outputs(985) <= (layer1_outputs(3784)) and not (layer1_outputs(4347));
    layer2_outputs(986) <= not((layer1_outputs(3747)) or (layer1_outputs(3200)));
    layer2_outputs(987) <= (layer1_outputs(4776)) and (layer1_outputs(3309));
    layer2_outputs(988) <= layer1_outputs(177);
    layer2_outputs(989) <= not((layer1_outputs(3133)) xor (layer1_outputs(2200)));
    layer2_outputs(990) <= (layer1_outputs(1665)) and not (layer1_outputs(320));
    layer2_outputs(991) <= layer1_outputs(2720);
    layer2_outputs(992) <= '1';
    layer2_outputs(993) <= not((layer1_outputs(4475)) and (layer1_outputs(3145)));
    layer2_outputs(994) <= (layer1_outputs(1043)) or (layer1_outputs(3193));
    layer2_outputs(995) <= (layer1_outputs(3458)) and (layer1_outputs(1876));
    layer2_outputs(996) <= layer1_outputs(4337);
    layer2_outputs(997) <= layer1_outputs(3074);
    layer2_outputs(998) <= not(layer1_outputs(2544));
    layer2_outputs(999) <= layer1_outputs(3057);
    layer2_outputs(1000) <= (layer1_outputs(1297)) and (layer1_outputs(4770));
    layer2_outputs(1001) <= not(layer1_outputs(59));
    layer2_outputs(1002) <= not(layer1_outputs(2392));
    layer2_outputs(1003) <= not(layer1_outputs(3154));
    layer2_outputs(1004) <= not(layer1_outputs(1140));
    layer2_outputs(1005) <= layer1_outputs(4901);
    layer2_outputs(1006) <= not((layer1_outputs(1057)) and (layer1_outputs(952)));
    layer2_outputs(1007) <= layer1_outputs(4915);
    layer2_outputs(1008) <= layer1_outputs(3418);
    layer2_outputs(1009) <= not(layer1_outputs(842));
    layer2_outputs(1010) <= not(layer1_outputs(4807)) or (layer1_outputs(2350));
    layer2_outputs(1011) <= (layer1_outputs(2711)) and (layer1_outputs(3015));
    layer2_outputs(1012) <= (layer1_outputs(1042)) and (layer1_outputs(4210));
    layer2_outputs(1013) <= (layer1_outputs(4442)) or (layer1_outputs(2010));
    layer2_outputs(1014) <= not(layer1_outputs(3630));
    layer2_outputs(1015) <= not(layer1_outputs(2770)) or (layer1_outputs(3328));
    layer2_outputs(1016) <= (layer1_outputs(3330)) or (layer1_outputs(2019));
    layer2_outputs(1017) <= not(layer1_outputs(1164)) or (layer1_outputs(1961));
    layer2_outputs(1018) <= not(layer1_outputs(162)) or (layer1_outputs(2232));
    layer2_outputs(1019) <= layer1_outputs(3844);
    layer2_outputs(1020) <= (layer1_outputs(4969)) or (layer1_outputs(3095));
    layer2_outputs(1021) <= (layer1_outputs(5008)) and not (layer1_outputs(1219));
    layer2_outputs(1022) <= layer1_outputs(5032);
    layer2_outputs(1023) <= layer1_outputs(4977);
    layer2_outputs(1024) <= (layer1_outputs(2825)) xor (layer1_outputs(2470));
    layer2_outputs(1025) <= not(layer1_outputs(880));
    layer2_outputs(1026) <= not(layer1_outputs(3794));
    layer2_outputs(1027) <= (layer1_outputs(1766)) or (layer1_outputs(1287));
    layer2_outputs(1028) <= not(layer1_outputs(982));
    layer2_outputs(1029) <= not((layer1_outputs(3279)) or (layer1_outputs(882)));
    layer2_outputs(1030) <= not(layer1_outputs(4349)) or (layer1_outputs(364));
    layer2_outputs(1031) <= (layer1_outputs(1250)) and not (layer1_outputs(3677));
    layer2_outputs(1032) <= not(layer1_outputs(4095));
    layer2_outputs(1033) <= not((layer1_outputs(2049)) or (layer1_outputs(5095)));
    layer2_outputs(1034) <= '0';
    layer2_outputs(1035) <= not(layer1_outputs(1242)) or (layer1_outputs(2569));
    layer2_outputs(1036) <= not(layer1_outputs(2808));
    layer2_outputs(1037) <= not(layer1_outputs(462));
    layer2_outputs(1038) <= layer1_outputs(2757);
    layer2_outputs(1039) <= (layer1_outputs(4811)) and (layer1_outputs(3287));
    layer2_outputs(1040) <= layer1_outputs(3611);
    layer2_outputs(1041) <= not(layer1_outputs(715)) or (layer1_outputs(4457));
    layer2_outputs(1042) <= (layer1_outputs(3866)) or (layer1_outputs(377));
    layer2_outputs(1043) <= not(layer1_outputs(4413)) or (layer1_outputs(4481));
    layer2_outputs(1044) <= not((layer1_outputs(145)) xor (layer1_outputs(13)));
    layer2_outputs(1045) <= layer1_outputs(4367);
    layer2_outputs(1046) <= not(layer1_outputs(4785));
    layer2_outputs(1047) <= (layer1_outputs(3703)) or (layer1_outputs(722));
    layer2_outputs(1048) <= not(layer1_outputs(2906));
    layer2_outputs(1049) <= layer1_outputs(2009);
    layer2_outputs(1050) <= layer1_outputs(219);
    layer2_outputs(1051) <= not(layer1_outputs(1578));
    layer2_outputs(1052) <= not(layer1_outputs(4645));
    layer2_outputs(1053) <= not(layer1_outputs(123));
    layer2_outputs(1054) <= not(layer1_outputs(1252)) or (layer1_outputs(1782));
    layer2_outputs(1055) <= (layer1_outputs(4522)) and not (layer1_outputs(1005));
    layer2_outputs(1056) <= (layer1_outputs(733)) or (layer1_outputs(4221));
    layer2_outputs(1057) <= not(layer1_outputs(4125)) or (layer1_outputs(4401));
    layer2_outputs(1058) <= not(layer1_outputs(2122));
    layer2_outputs(1059) <= (layer1_outputs(2765)) and (layer1_outputs(2685));
    layer2_outputs(1060) <= not(layer1_outputs(3963));
    layer2_outputs(1061) <= layer1_outputs(4345);
    layer2_outputs(1062) <= layer1_outputs(3428);
    layer2_outputs(1063) <= layer1_outputs(4787);
    layer2_outputs(1064) <= not(layer1_outputs(1757));
    layer2_outputs(1065) <= not(layer1_outputs(2221)) or (layer1_outputs(699));
    layer2_outputs(1066) <= not(layer1_outputs(2395));
    layer2_outputs(1067) <= (layer1_outputs(4781)) and not (layer1_outputs(1370));
    layer2_outputs(1068) <= (layer1_outputs(3143)) or (layer1_outputs(3812));
    layer2_outputs(1069) <= not((layer1_outputs(1629)) or (layer1_outputs(1954)));
    layer2_outputs(1070) <= layer1_outputs(1560);
    layer2_outputs(1071) <= (layer1_outputs(3569)) and (layer1_outputs(3957));
    layer2_outputs(1072) <= not(layer1_outputs(3274)) or (layer1_outputs(3823));
    layer2_outputs(1073) <= layer1_outputs(4500);
    layer2_outputs(1074) <= not(layer1_outputs(577));
    layer2_outputs(1075) <= not((layer1_outputs(3926)) or (layer1_outputs(3862)));
    layer2_outputs(1076) <= not(layer1_outputs(4836));
    layer2_outputs(1077) <= (layer1_outputs(1189)) xor (layer1_outputs(1733));
    layer2_outputs(1078) <= not(layer1_outputs(3414)) or (layer1_outputs(3326));
    layer2_outputs(1079) <= not(layer1_outputs(4298));
    layer2_outputs(1080) <= not(layer1_outputs(1506)) or (layer1_outputs(1583));
    layer2_outputs(1081) <= not((layer1_outputs(4209)) xor (layer1_outputs(4159)));
    layer2_outputs(1082) <= not(layer1_outputs(3037)) or (layer1_outputs(1449));
    layer2_outputs(1083) <= not((layer1_outputs(83)) or (layer1_outputs(1274)));
    layer2_outputs(1084) <= not(layer1_outputs(3729));
    layer2_outputs(1085) <= (layer1_outputs(3371)) or (layer1_outputs(2761));
    layer2_outputs(1086) <= not(layer1_outputs(1236));
    layer2_outputs(1087) <= not(layer1_outputs(3508));
    layer2_outputs(1088) <= layer1_outputs(1579);
    layer2_outputs(1089) <= layer1_outputs(1743);
    layer2_outputs(1090) <= (layer1_outputs(2312)) xor (layer1_outputs(3796));
    layer2_outputs(1091) <= (layer1_outputs(1524)) xor (layer1_outputs(321));
    layer2_outputs(1092) <= layer1_outputs(3189);
    layer2_outputs(1093) <= not((layer1_outputs(4909)) xor (layer1_outputs(3420)));
    layer2_outputs(1094) <= layer1_outputs(4420);
    layer2_outputs(1095) <= not((layer1_outputs(4954)) and (layer1_outputs(3684)));
    layer2_outputs(1096) <= not((layer1_outputs(1806)) xor (layer1_outputs(334)));
    layer2_outputs(1097) <= (layer1_outputs(2230)) xor (layer1_outputs(3901));
    layer2_outputs(1098) <= not((layer1_outputs(2557)) and (layer1_outputs(1686)));
    layer2_outputs(1099) <= layer1_outputs(2841);
    layer2_outputs(1100) <= layer1_outputs(2261);
    layer2_outputs(1101) <= (layer1_outputs(4678)) or (layer1_outputs(2811));
    layer2_outputs(1102) <= layer1_outputs(2251);
    layer2_outputs(1103) <= layer1_outputs(1155);
    layer2_outputs(1104) <= not((layer1_outputs(3616)) xor (layer1_outputs(568)));
    layer2_outputs(1105) <= not((layer1_outputs(55)) or (layer1_outputs(3148)));
    layer2_outputs(1106) <= not(layer1_outputs(2794));
    layer2_outputs(1107) <= (layer1_outputs(2409)) and not (layer1_outputs(2957));
    layer2_outputs(1108) <= not(layer1_outputs(2927));
    layer2_outputs(1109) <= (layer1_outputs(3730)) and not (layer1_outputs(4158));
    layer2_outputs(1110) <= not((layer1_outputs(4232)) xor (layer1_outputs(1845)));
    layer2_outputs(1111) <= (layer1_outputs(1334)) and not (layer1_outputs(3289));
    layer2_outputs(1112) <= layer1_outputs(821);
    layer2_outputs(1113) <= not((layer1_outputs(2738)) and (layer1_outputs(4878)));
    layer2_outputs(1114) <= (layer1_outputs(2046)) and (layer1_outputs(1169));
    layer2_outputs(1115) <= not(layer1_outputs(1880));
    layer2_outputs(1116) <= (layer1_outputs(3483)) and not (layer1_outputs(1661));
    layer2_outputs(1117) <= (layer1_outputs(1423)) and not (layer1_outputs(1490));
    layer2_outputs(1118) <= not(layer1_outputs(4735));
    layer2_outputs(1119) <= not(layer1_outputs(4710));
    layer2_outputs(1120) <= not((layer1_outputs(1553)) xor (layer1_outputs(2137)));
    layer2_outputs(1121) <= not((layer1_outputs(2666)) xor (layer1_outputs(1103)));
    layer2_outputs(1122) <= not(layer1_outputs(3344)) or (layer1_outputs(1234));
    layer2_outputs(1123) <= layer1_outputs(1264);
    layer2_outputs(1124) <= not(layer1_outputs(1172)) or (layer1_outputs(4807));
    layer2_outputs(1125) <= layer1_outputs(1275);
    layer2_outputs(1126) <= not((layer1_outputs(314)) xor (layer1_outputs(1826)));
    layer2_outputs(1127) <= not(layer1_outputs(2609));
    layer2_outputs(1128) <= not(layer1_outputs(1141));
    layer2_outputs(1129) <= not(layer1_outputs(1112)) or (layer1_outputs(1427));
    layer2_outputs(1130) <= not((layer1_outputs(567)) and (layer1_outputs(3009)));
    layer2_outputs(1131) <= not(layer1_outputs(3453));
    layer2_outputs(1132) <= layer1_outputs(2447);
    layer2_outputs(1133) <= layer1_outputs(1341);
    layer2_outputs(1134) <= (layer1_outputs(2944)) and (layer1_outputs(1007));
    layer2_outputs(1135) <= (layer1_outputs(4875)) or (layer1_outputs(4757));
    layer2_outputs(1136) <= not((layer1_outputs(180)) xor (layer1_outputs(4531)));
    layer2_outputs(1137) <= not(layer1_outputs(4938)) or (layer1_outputs(4991));
    layer2_outputs(1138) <= not((layer1_outputs(411)) and (layer1_outputs(4503)));
    layer2_outputs(1139) <= '0';
    layer2_outputs(1140) <= not(layer1_outputs(3988));
    layer2_outputs(1141) <= layer1_outputs(915);
    layer2_outputs(1142) <= not(layer1_outputs(4161));
    layer2_outputs(1143) <= not(layer1_outputs(862));
    layer2_outputs(1144) <= layer1_outputs(4944);
    layer2_outputs(1145) <= not(layer1_outputs(937)) or (layer1_outputs(1119));
    layer2_outputs(1146) <= not((layer1_outputs(549)) xor (layer1_outputs(2191)));
    layer2_outputs(1147) <= (layer1_outputs(3614)) or (layer1_outputs(3943));
    layer2_outputs(1148) <= (layer1_outputs(2865)) and not (layer1_outputs(686));
    layer2_outputs(1149) <= not(layer1_outputs(1168));
    layer2_outputs(1150) <= (layer1_outputs(4050)) and not (layer1_outputs(3619));
    layer2_outputs(1151) <= (layer1_outputs(1515)) and not (layer1_outputs(446));
    layer2_outputs(1152) <= (layer1_outputs(3884)) and not (layer1_outputs(3367));
    layer2_outputs(1153) <= layer1_outputs(430);
    layer2_outputs(1154) <= layer1_outputs(2551);
    layer2_outputs(1155) <= not((layer1_outputs(3930)) or (layer1_outputs(5014)));
    layer2_outputs(1156) <= not(layer1_outputs(3310));
    layer2_outputs(1157) <= not(layer1_outputs(1633));
    layer2_outputs(1158) <= not((layer1_outputs(4103)) or (layer1_outputs(3847)));
    layer2_outputs(1159) <= not(layer1_outputs(3424));
    layer2_outputs(1160) <= not(layer1_outputs(301));
    layer2_outputs(1161) <= not(layer1_outputs(1679));
    layer2_outputs(1162) <= not((layer1_outputs(872)) and (layer1_outputs(1904)));
    layer2_outputs(1163) <= layer1_outputs(1525);
    layer2_outputs(1164) <= layer1_outputs(4754);
    layer2_outputs(1165) <= layer1_outputs(3908);
    layer2_outputs(1166) <= (layer1_outputs(4025)) and not (layer1_outputs(2886));
    layer2_outputs(1167) <= not(layer1_outputs(2593));
    layer2_outputs(1168) <= (layer1_outputs(1435)) and (layer1_outputs(2702));
    layer2_outputs(1169) <= layer1_outputs(1754);
    layer2_outputs(1170) <= not(layer1_outputs(4889));
    layer2_outputs(1171) <= not(layer1_outputs(4932));
    layer2_outputs(1172) <= layer1_outputs(1185);
    layer2_outputs(1173) <= (layer1_outputs(1643)) or (layer1_outputs(4416));
    layer2_outputs(1174) <= (layer1_outputs(4939)) and not (layer1_outputs(1081));
    layer2_outputs(1175) <= not(layer1_outputs(4994));
    layer2_outputs(1176) <= not((layer1_outputs(1467)) and (layer1_outputs(1691)));
    layer2_outputs(1177) <= not(layer1_outputs(3473));
    layer2_outputs(1178) <= layer1_outputs(4432);
    layer2_outputs(1179) <= not(layer1_outputs(587)) or (layer1_outputs(898));
    layer2_outputs(1180) <= (layer1_outputs(3988)) and not (layer1_outputs(3385));
    layer2_outputs(1181) <= not(layer1_outputs(2970));
    layer2_outputs(1182) <= not((layer1_outputs(3523)) and (layer1_outputs(940)));
    layer2_outputs(1183) <= (layer1_outputs(72)) and not (layer1_outputs(608));
    layer2_outputs(1184) <= (layer1_outputs(2640)) and (layer1_outputs(120));
    layer2_outputs(1185) <= (layer1_outputs(4716)) and (layer1_outputs(5074));
    layer2_outputs(1186) <= (layer1_outputs(2584)) and (layer1_outputs(3349));
    layer2_outputs(1187) <= (layer1_outputs(4984)) and not (layer1_outputs(4340));
    layer2_outputs(1188) <= not(layer1_outputs(1517));
    layer2_outputs(1189) <= not((layer1_outputs(2940)) or (layer1_outputs(3922)));
    layer2_outputs(1190) <= layer1_outputs(1538);
    layer2_outputs(1191) <= not(layer1_outputs(1015));
    layer2_outputs(1192) <= (layer1_outputs(2569)) and (layer1_outputs(1335));
    layer2_outputs(1193) <= (layer1_outputs(2165)) or (layer1_outputs(3635));
    layer2_outputs(1194) <= not(layer1_outputs(3316));
    layer2_outputs(1195) <= not(layer1_outputs(2423)) or (layer1_outputs(677));
    layer2_outputs(1196) <= not(layer1_outputs(277));
    layer2_outputs(1197) <= layer1_outputs(1402);
    layer2_outputs(1198) <= not((layer1_outputs(2637)) xor (layer1_outputs(2339)));
    layer2_outputs(1199) <= (layer1_outputs(4395)) or (layer1_outputs(4472));
    layer2_outputs(1200) <= layer1_outputs(3068);
    layer2_outputs(1201) <= layer1_outputs(2621);
    layer2_outputs(1202) <= not(layer1_outputs(1454)) or (layer1_outputs(3004));
    layer2_outputs(1203) <= not((layer1_outputs(1477)) or (layer1_outputs(3606)));
    layer2_outputs(1204) <= not((layer1_outputs(1303)) or (layer1_outputs(3364)));
    layer2_outputs(1205) <= not(layer1_outputs(3561));
    layer2_outputs(1206) <= not(layer1_outputs(350));
    layer2_outputs(1207) <= not(layer1_outputs(4968));
    layer2_outputs(1208) <= not(layer1_outputs(2914));
    layer2_outputs(1209) <= '0';
    layer2_outputs(1210) <= layer1_outputs(817);
    layer2_outputs(1211) <= layer1_outputs(4450);
    layer2_outputs(1212) <= '0';
    layer2_outputs(1213) <= layer1_outputs(1763);
    layer2_outputs(1214) <= not(layer1_outputs(1111));
    layer2_outputs(1215) <= layer1_outputs(3100);
    layer2_outputs(1216) <= not((layer1_outputs(3567)) and (layer1_outputs(3737)));
    layer2_outputs(1217) <= not(layer1_outputs(4509));
    layer2_outputs(1218) <= (layer1_outputs(4456)) xor (layer1_outputs(2282));
    layer2_outputs(1219) <= layer1_outputs(3927);
    layer2_outputs(1220) <= layer1_outputs(2103);
    layer2_outputs(1221) <= not(layer1_outputs(4240)) or (layer1_outputs(1270));
    layer2_outputs(1222) <= not((layer1_outputs(2905)) or (layer1_outputs(709)));
    layer2_outputs(1223) <= layer1_outputs(1085);
    layer2_outputs(1224) <= layer1_outputs(1391);
    layer2_outputs(1225) <= (layer1_outputs(578)) and not (layer1_outputs(1743));
    layer2_outputs(1226) <= layer1_outputs(1441);
    layer2_outputs(1227) <= not(layer1_outputs(412));
    layer2_outputs(1228) <= not((layer1_outputs(3511)) xor (layer1_outputs(234)));
    layer2_outputs(1229) <= not(layer1_outputs(4279)) or (layer1_outputs(2713));
    layer2_outputs(1230) <= (layer1_outputs(2052)) and not (layer1_outputs(1625));
    layer2_outputs(1231) <= (layer1_outputs(5073)) xor (layer1_outputs(2181));
    layer2_outputs(1232) <= (layer1_outputs(1662)) or (layer1_outputs(1617));
    layer2_outputs(1233) <= not(layer1_outputs(61));
    layer2_outputs(1234) <= layer1_outputs(1396);
    layer2_outputs(1235) <= not(layer1_outputs(805));
    layer2_outputs(1236) <= not((layer1_outputs(1992)) and (layer1_outputs(4610)));
    layer2_outputs(1237) <= layer1_outputs(3220);
    layer2_outputs(1238) <= (layer1_outputs(4135)) and not (layer1_outputs(1816));
    layer2_outputs(1239) <= not(layer1_outputs(4049));
    layer2_outputs(1240) <= not((layer1_outputs(2352)) xor (layer1_outputs(1408)));
    layer2_outputs(1241) <= not(layer1_outputs(2123)) or (layer1_outputs(4482));
    layer2_outputs(1242) <= layer1_outputs(2536);
    layer2_outputs(1243) <= not(layer1_outputs(2247)) or (layer1_outputs(1047));
    layer2_outputs(1244) <= not((layer1_outputs(722)) or (layer1_outputs(1953)));
    layer2_outputs(1245) <= not((layer1_outputs(959)) xor (layer1_outputs(3734)));
    layer2_outputs(1246) <= layer1_outputs(1057);
    layer2_outputs(1247) <= (layer1_outputs(1818)) xor (layer1_outputs(617));
    layer2_outputs(1248) <= not((layer1_outputs(1382)) and (layer1_outputs(3373)));
    layer2_outputs(1249) <= layer1_outputs(2115);
    layer2_outputs(1250) <= layer1_outputs(810);
    layer2_outputs(1251) <= (layer1_outputs(3533)) or (layer1_outputs(4806));
    layer2_outputs(1252) <= not(layer1_outputs(1541));
    layer2_outputs(1253) <= not((layer1_outputs(4988)) xor (layer1_outputs(1164)));
    layer2_outputs(1254) <= not(layer1_outputs(3177)) or (layer1_outputs(1107));
    layer2_outputs(1255) <= layer1_outputs(925);
    layer2_outputs(1256) <= (layer1_outputs(647)) and not (layer1_outputs(301));
    layer2_outputs(1257) <= (layer1_outputs(5111)) and not (layer1_outputs(809));
    layer2_outputs(1258) <= (layer1_outputs(25)) or (layer1_outputs(3795));
    layer2_outputs(1259) <= not((layer1_outputs(1571)) xor (layer1_outputs(2541)));
    layer2_outputs(1260) <= layer1_outputs(3840);
    layer2_outputs(1261) <= '0';
    layer2_outputs(1262) <= layer1_outputs(4945);
    layer2_outputs(1263) <= not(layer1_outputs(2216));
    layer2_outputs(1264) <= not(layer1_outputs(4101));
    layer2_outputs(1265) <= not(layer1_outputs(3880)) or (layer1_outputs(561));
    layer2_outputs(1266) <= (layer1_outputs(845)) and (layer1_outputs(1802));
    layer2_outputs(1267) <= not(layer1_outputs(3852)) or (layer1_outputs(1782));
    layer2_outputs(1268) <= not((layer1_outputs(2995)) and (layer1_outputs(2436)));
    layer2_outputs(1269) <= not(layer1_outputs(2176));
    layer2_outputs(1270) <= layer1_outputs(3853);
    layer2_outputs(1271) <= (layer1_outputs(4123)) and not (layer1_outputs(2659));
    layer2_outputs(1272) <= (layer1_outputs(89)) xor (layer1_outputs(2461));
    layer2_outputs(1273) <= (layer1_outputs(2922)) xor (layer1_outputs(1534));
    layer2_outputs(1274) <= layer1_outputs(4157);
    layer2_outputs(1275) <= layer1_outputs(4993);
    layer2_outputs(1276) <= (layer1_outputs(1637)) and (layer1_outputs(2994));
    layer2_outputs(1277) <= layer1_outputs(4067);
    layer2_outputs(1278) <= not(layer1_outputs(244)) or (layer1_outputs(4834));
    layer2_outputs(1279) <= not(layer1_outputs(889));
    layer2_outputs(1280) <= not(layer1_outputs(3096));
    layer2_outputs(1281) <= layer1_outputs(1170);
    layer2_outputs(1282) <= not(layer1_outputs(3744));
    layer2_outputs(1283) <= not((layer1_outputs(1760)) or (layer1_outputs(3438)));
    layer2_outputs(1284) <= (layer1_outputs(641)) or (layer1_outputs(3376));
    layer2_outputs(1285) <= layer1_outputs(4167);
    layer2_outputs(1286) <= (layer1_outputs(119)) or (layer1_outputs(3976));
    layer2_outputs(1287) <= not(layer1_outputs(2404)) or (layer1_outputs(763));
    layer2_outputs(1288) <= layer1_outputs(3174);
    layer2_outputs(1289) <= not((layer1_outputs(1701)) xor (layer1_outputs(4740)));
    layer2_outputs(1290) <= (layer1_outputs(1002)) xor (layer1_outputs(1340));
    layer2_outputs(1291) <= not(layer1_outputs(4753));
    layer2_outputs(1292) <= layer1_outputs(1702);
    layer2_outputs(1293) <= not(layer1_outputs(663)) or (layer1_outputs(3826));
    layer2_outputs(1294) <= not(layer1_outputs(1463));
    layer2_outputs(1295) <= not(layer1_outputs(3518));
    layer2_outputs(1296) <= layer1_outputs(2924);
    layer2_outputs(1297) <= layer1_outputs(5058);
    layer2_outputs(1298) <= not((layer1_outputs(4755)) or (layer1_outputs(1918)));
    layer2_outputs(1299) <= layer1_outputs(1718);
    layer2_outputs(1300) <= not(layer1_outputs(2758));
    layer2_outputs(1301) <= not((layer1_outputs(4584)) xor (layer1_outputs(2522)));
    layer2_outputs(1302) <= not(layer1_outputs(3246));
    layer2_outputs(1303) <= (layer1_outputs(1380)) xor (layer1_outputs(4364));
    layer2_outputs(1304) <= (layer1_outputs(1778)) or (layer1_outputs(949));
    layer2_outputs(1305) <= layer1_outputs(0);
    layer2_outputs(1306) <= not((layer1_outputs(4940)) or (layer1_outputs(888)));
    layer2_outputs(1307) <= (layer1_outputs(1305)) xor (layer1_outputs(1323));
    layer2_outputs(1308) <= not(layer1_outputs(780));
    layer2_outputs(1309) <= not((layer1_outputs(996)) xor (layer1_outputs(1216)));
    layer2_outputs(1310) <= layer1_outputs(997);
    layer2_outputs(1311) <= not(layer1_outputs(1875)) or (layer1_outputs(655));
    layer2_outputs(1312) <= (layer1_outputs(4714)) and not (layer1_outputs(915));
    layer2_outputs(1313) <= layer1_outputs(4078);
    layer2_outputs(1314) <= layer1_outputs(437);
    layer2_outputs(1315) <= not(layer1_outputs(1708));
    layer2_outputs(1316) <= layer1_outputs(1765);
    layer2_outputs(1317) <= not((layer1_outputs(3062)) and (layer1_outputs(3792)));
    layer2_outputs(1318) <= not((layer1_outputs(2583)) or (layer1_outputs(2163)));
    layer2_outputs(1319) <= (layer1_outputs(3168)) and not (layer1_outputs(3406));
    layer2_outputs(1320) <= (layer1_outputs(1622)) and not (layer1_outputs(2490));
    layer2_outputs(1321) <= not(layer1_outputs(439));
    layer2_outputs(1322) <= layer1_outputs(3318);
    layer2_outputs(1323) <= layer1_outputs(2933);
    layer2_outputs(1324) <= (layer1_outputs(2125)) and not (layer1_outputs(297));
    layer2_outputs(1325) <= not((layer1_outputs(3310)) and (layer1_outputs(4375)));
    layer2_outputs(1326) <= (layer1_outputs(3441)) and (layer1_outputs(2608));
    layer2_outputs(1327) <= not(layer1_outputs(3544));
    layer2_outputs(1328) <= (layer1_outputs(1953)) and (layer1_outputs(3533));
    layer2_outputs(1329) <= not(layer1_outputs(2706));
    layer2_outputs(1330) <= not(layer1_outputs(2003));
    layer2_outputs(1331) <= (layer1_outputs(3325)) xor (layer1_outputs(1235));
    layer2_outputs(1332) <= (layer1_outputs(3003)) and not (layer1_outputs(908));
    layer2_outputs(1333) <= (layer1_outputs(45)) xor (layer1_outputs(4712));
    layer2_outputs(1334) <= layer1_outputs(4905);
    layer2_outputs(1335) <= layer1_outputs(783);
    layer2_outputs(1336) <= not((layer1_outputs(3637)) and (layer1_outputs(4823)));
    layer2_outputs(1337) <= layer1_outputs(2874);
    layer2_outputs(1338) <= not(layer1_outputs(1444)) or (layer1_outputs(3573));
    layer2_outputs(1339) <= not((layer1_outputs(798)) or (layer1_outputs(2935)));
    layer2_outputs(1340) <= (layer1_outputs(170)) xor (layer1_outputs(1781));
    layer2_outputs(1341) <= layer1_outputs(4825);
    layer2_outputs(1342) <= (layer1_outputs(3987)) and not (layer1_outputs(2899));
    layer2_outputs(1343) <= not(layer1_outputs(1618));
    layer2_outputs(1344) <= (layer1_outputs(4435)) and (layer1_outputs(4187));
    layer2_outputs(1345) <= not(layer1_outputs(1060));
    layer2_outputs(1346) <= (layer1_outputs(4181)) and not (layer1_outputs(2736));
    layer2_outputs(1347) <= not(layer1_outputs(3671));
    layer2_outputs(1348) <= not(layer1_outputs(4182));
    layer2_outputs(1349) <= not((layer1_outputs(4619)) xor (layer1_outputs(1136)));
    layer2_outputs(1350) <= layer1_outputs(2988);
    layer2_outputs(1351) <= not(layer1_outputs(640));
    layer2_outputs(1352) <= (layer1_outputs(1265)) and not (layer1_outputs(2074));
    layer2_outputs(1353) <= not(layer1_outputs(3478));
    layer2_outputs(1354) <= not(layer1_outputs(4137));
    layer2_outputs(1355) <= not(layer1_outputs(90));
    layer2_outputs(1356) <= (layer1_outputs(1909)) and (layer1_outputs(3278));
    layer2_outputs(1357) <= not((layer1_outputs(4806)) and (layer1_outputs(2120)));
    layer2_outputs(1358) <= not(layer1_outputs(698));
    layer2_outputs(1359) <= (layer1_outputs(1904)) and (layer1_outputs(1183));
    layer2_outputs(1360) <= (layer1_outputs(4606)) and not (layer1_outputs(1031));
    layer2_outputs(1361) <= (layer1_outputs(2166)) and (layer1_outputs(209));
    layer2_outputs(1362) <= (layer1_outputs(4342)) and (layer1_outputs(4));
    layer2_outputs(1363) <= (layer1_outputs(1581)) xor (layer1_outputs(2606));
    layer2_outputs(1364) <= (layer1_outputs(1631)) and (layer1_outputs(2810));
    layer2_outputs(1365) <= (layer1_outputs(4619)) xor (layer1_outputs(4424));
    layer2_outputs(1366) <= not(layer1_outputs(3046));
    layer2_outputs(1367) <= (layer1_outputs(2439)) or (layer1_outputs(1625));
    layer2_outputs(1368) <= not(layer1_outputs(2984));
    layer2_outputs(1369) <= not((layer1_outputs(2706)) or (layer1_outputs(3516)));
    layer2_outputs(1370) <= layer1_outputs(4659);
    layer2_outputs(1371) <= (layer1_outputs(362)) and not (layer1_outputs(544));
    layer2_outputs(1372) <= (layer1_outputs(211)) and (layer1_outputs(3129));
    layer2_outputs(1373) <= (layer1_outputs(971)) and not (layer1_outputs(736));
    layer2_outputs(1374) <= not((layer1_outputs(3891)) xor (layer1_outputs(3837)));
    layer2_outputs(1375) <= (layer1_outputs(2708)) and (layer1_outputs(2750));
    layer2_outputs(1376) <= layer1_outputs(4706);
    layer2_outputs(1377) <= layer1_outputs(4606);
    layer2_outputs(1378) <= (layer1_outputs(1795)) xor (layer1_outputs(1546));
    layer2_outputs(1379) <= layer1_outputs(1199);
    layer2_outputs(1380) <= not(layer1_outputs(4943)) or (layer1_outputs(2243));
    layer2_outputs(1381) <= '1';
    layer2_outputs(1382) <= layer1_outputs(2318);
    layer2_outputs(1383) <= (layer1_outputs(1478)) xor (layer1_outputs(2000));
    layer2_outputs(1384) <= not(layer1_outputs(4648)) or (layer1_outputs(3196));
    layer2_outputs(1385) <= not((layer1_outputs(67)) and (layer1_outputs(3051)));
    layer2_outputs(1386) <= not((layer1_outputs(1621)) xor (layer1_outputs(4062)));
    layer2_outputs(1387) <= layer1_outputs(4997);
    layer2_outputs(1388) <= not((layer1_outputs(1746)) xor (layer1_outputs(66)));
    layer2_outputs(1389) <= layer1_outputs(4435);
    layer2_outputs(1390) <= (layer1_outputs(2073)) xor (layer1_outputs(1055));
    layer2_outputs(1391) <= (layer1_outputs(4886)) and (layer1_outputs(571));
    layer2_outputs(1392) <= (layer1_outputs(1653)) or (layer1_outputs(620));
    layer2_outputs(1393) <= (layer1_outputs(2549)) xor (layer1_outputs(3698));
    layer2_outputs(1394) <= not(layer1_outputs(855));
    layer2_outputs(1395) <= not(layer1_outputs(4972));
    layer2_outputs(1396) <= layer1_outputs(1163);
    layer2_outputs(1397) <= (layer1_outputs(4127)) and not (layer1_outputs(2021));
    layer2_outputs(1398) <= layer1_outputs(2036);
    layer2_outputs(1399) <= layer1_outputs(1067);
    layer2_outputs(1400) <= not(layer1_outputs(1862));
    layer2_outputs(1401) <= not((layer1_outputs(3002)) and (layer1_outputs(2018)));
    layer2_outputs(1402) <= not(layer1_outputs(3655));
    layer2_outputs(1403) <= (layer1_outputs(2955)) and not (layer1_outputs(320));
    layer2_outputs(1404) <= not((layer1_outputs(2450)) or (layer1_outputs(4730)));
    layer2_outputs(1405) <= (layer1_outputs(3126)) or (layer1_outputs(593));
    layer2_outputs(1406) <= (layer1_outputs(4778)) and not (layer1_outputs(3402));
    layer2_outputs(1407) <= layer1_outputs(2575);
    layer2_outputs(1408) <= layer1_outputs(1181);
    layer2_outputs(1409) <= layer1_outputs(4548);
    layer2_outputs(1410) <= (layer1_outputs(3647)) and (layer1_outputs(2011));
    layer2_outputs(1411) <= layer1_outputs(3840);
    layer2_outputs(1412) <= not((layer1_outputs(1158)) and (layer1_outputs(638)));
    layer2_outputs(1413) <= not((layer1_outputs(2012)) xor (layer1_outputs(724)));
    layer2_outputs(1414) <= layer1_outputs(568);
    layer2_outputs(1415) <= not((layer1_outputs(4368)) and (layer1_outputs(1984)));
    layer2_outputs(1416) <= (layer1_outputs(4928)) and not (layer1_outputs(1378));
    layer2_outputs(1417) <= not(layer1_outputs(4587));
    layer2_outputs(1418) <= not((layer1_outputs(107)) xor (layer1_outputs(3649)));
    layer2_outputs(1419) <= not((layer1_outputs(1371)) xor (layer1_outputs(779)));
    layer2_outputs(1420) <= not(layer1_outputs(2826));
    layer2_outputs(1421) <= layer1_outputs(1205);
    layer2_outputs(1422) <= not(layer1_outputs(4473));
    layer2_outputs(1423) <= layer1_outputs(4334);
    layer2_outputs(1424) <= not(layer1_outputs(686));
    layer2_outputs(1425) <= layer1_outputs(509);
    layer2_outputs(1426) <= layer1_outputs(4182);
    layer2_outputs(1427) <= not((layer1_outputs(3332)) and (layer1_outputs(705)));
    layer2_outputs(1428) <= (layer1_outputs(2947)) and not (layer1_outputs(2167));
    layer2_outputs(1429) <= not(layer1_outputs(4952));
    layer2_outputs(1430) <= not(layer1_outputs(2186));
    layer2_outputs(1431) <= layer1_outputs(147);
    layer2_outputs(1432) <= (layer1_outputs(4228)) and (layer1_outputs(297));
    layer2_outputs(1433) <= (layer1_outputs(2301)) xor (layer1_outputs(396));
    layer2_outputs(1434) <= not(layer1_outputs(3086));
    layer2_outputs(1435) <= layer1_outputs(4175);
    layer2_outputs(1436) <= (layer1_outputs(761)) and (layer1_outputs(4032));
    layer2_outputs(1437) <= not((layer1_outputs(606)) and (layer1_outputs(3810)));
    layer2_outputs(1438) <= (layer1_outputs(863)) or (layer1_outputs(3564));
    layer2_outputs(1439) <= (layer1_outputs(5069)) and (layer1_outputs(4970));
    layer2_outputs(1440) <= layer1_outputs(1151);
    layer2_outputs(1441) <= (layer1_outputs(1551)) and (layer1_outputs(4515));
    layer2_outputs(1442) <= not(layer1_outputs(4467));
    layer2_outputs(1443) <= (layer1_outputs(4040)) and not (layer1_outputs(4220));
    layer2_outputs(1444) <= not(layer1_outputs(2537));
    layer2_outputs(1445) <= layer1_outputs(2183);
    layer2_outputs(1446) <= not((layer1_outputs(2842)) or (layer1_outputs(4188)));
    layer2_outputs(1447) <= (layer1_outputs(420)) and (layer1_outputs(2410));
    layer2_outputs(1448) <= (layer1_outputs(1749)) and not (layer1_outputs(1241));
    layer2_outputs(1449) <= (layer1_outputs(2430)) or (layer1_outputs(829));
    layer2_outputs(1450) <= '0';
    layer2_outputs(1451) <= not((layer1_outputs(3199)) and (layer1_outputs(3344)));
    layer2_outputs(1452) <= not((layer1_outputs(3665)) xor (layer1_outputs(932)));
    layer2_outputs(1453) <= layer1_outputs(3445);
    layer2_outputs(1454) <= not(layer1_outputs(5049));
    layer2_outputs(1455) <= not(layer1_outputs(189));
    layer2_outputs(1456) <= layer1_outputs(422);
    layer2_outputs(1457) <= not((layer1_outputs(1786)) xor (layer1_outputs(1822)));
    layer2_outputs(1458) <= not(layer1_outputs(2160)) or (layer1_outputs(3080));
    layer2_outputs(1459) <= not((layer1_outputs(4229)) and (layer1_outputs(541)));
    layer2_outputs(1460) <= (layer1_outputs(2923)) and not (layer1_outputs(911));
    layer2_outputs(1461) <= not(layer1_outputs(3444));
    layer2_outputs(1462) <= layer1_outputs(1891);
    layer2_outputs(1463) <= (layer1_outputs(2402)) xor (layer1_outputs(4308));
    layer2_outputs(1464) <= not(layer1_outputs(2768)) or (layer1_outputs(3271));
    layer2_outputs(1465) <= (layer1_outputs(2556)) or (layer1_outputs(2169));
    layer2_outputs(1466) <= (layer1_outputs(1755)) or (layer1_outputs(225));
    layer2_outputs(1467) <= '0';
    layer2_outputs(1468) <= (layer1_outputs(3541)) xor (layer1_outputs(105));
    layer2_outputs(1469) <= layer1_outputs(5028);
    layer2_outputs(1470) <= '0';
    layer2_outputs(1471) <= (layer1_outputs(2593)) and not (layer1_outputs(168));
    layer2_outputs(1472) <= layer1_outputs(2688);
    layer2_outputs(1473) <= layer1_outputs(3915);
    layer2_outputs(1474) <= layer1_outputs(381);
    layer2_outputs(1475) <= layer1_outputs(2729);
    layer2_outputs(1476) <= not(layer1_outputs(4930));
    layer2_outputs(1477) <= layer1_outputs(683);
    layer2_outputs(1478) <= (layer1_outputs(1785)) or (layer1_outputs(1120));
    layer2_outputs(1479) <= '0';
    layer2_outputs(1480) <= (layer1_outputs(2910)) and (layer1_outputs(1322));
    layer2_outputs(1481) <= (layer1_outputs(2492)) or (layer1_outputs(4995));
    layer2_outputs(1482) <= layer1_outputs(4283);
    layer2_outputs(1483) <= not((layer1_outputs(2424)) and (layer1_outputs(593)));
    layer2_outputs(1484) <= not((layer1_outputs(286)) and (layer1_outputs(2420)));
    layer2_outputs(1485) <= not(layer1_outputs(931));
    layer2_outputs(1486) <= (layer1_outputs(1941)) and (layer1_outputs(101));
    layer2_outputs(1487) <= not(layer1_outputs(1598));
    layer2_outputs(1488) <= layer1_outputs(4793);
    layer2_outputs(1489) <= not((layer1_outputs(4613)) and (layer1_outputs(895)));
    layer2_outputs(1490) <= layer1_outputs(1840);
    layer2_outputs(1491) <= not(layer1_outputs(3405));
    layer2_outputs(1492) <= not((layer1_outputs(1462)) xor (layer1_outputs(681)));
    layer2_outputs(1493) <= (layer1_outputs(1304)) and not (layer1_outputs(2127));
    layer2_outputs(1494) <= layer1_outputs(3366);
    layer2_outputs(1495) <= not(layer1_outputs(2254));
    layer2_outputs(1496) <= not(layer1_outputs(1709));
    layer2_outputs(1497) <= (layer1_outputs(2249)) and not (layer1_outputs(3570));
    layer2_outputs(1498) <= not(layer1_outputs(2069)) or (layer1_outputs(1836));
    layer2_outputs(1499) <= layer1_outputs(1531);
    layer2_outputs(1500) <= not(layer1_outputs(2280));
    layer2_outputs(1501) <= not(layer1_outputs(4551));
    layer2_outputs(1502) <= not(layer1_outputs(1137));
    layer2_outputs(1503) <= layer1_outputs(1476);
    layer2_outputs(1504) <= layer1_outputs(3223);
    layer2_outputs(1505) <= not(layer1_outputs(527)) or (layer1_outputs(3125));
    layer2_outputs(1506) <= (layer1_outputs(4547)) xor (layer1_outputs(2237));
    layer2_outputs(1507) <= layer1_outputs(4321);
    layer2_outputs(1508) <= not(layer1_outputs(5086));
    layer2_outputs(1509) <= layer1_outputs(4389);
    layer2_outputs(1510) <= layer1_outputs(780);
    layer2_outputs(1511) <= not(layer1_outputs(4643));
    layer2_outputs(1512) <= (layer1_outputs(2766)) and (layer1_outputs(3532));
    layer2_outputs(1513) <= (layer1_outputs(669)) and not (layer1_outputs(1419));
    layer2_outputs(1514) <= not(layer1_outputs(710));
    layer2_outputs(1515) <= layer1_outputs(4349);
    layer2_outputs(1516) <= (layer1_outputs(1732)) or (layer1_outputs(533));
    layer2_outputs(1517) <= (layer1_outputs(3395)) and not (layer1_outputs(4934));
    layer2_outputs(1518) <= not(layer1_outputs(2379));
    layer2_outputs(1519) <= (layer1_outputs(918)) and not (layer1_outputs(3393));
    layer2_outputs(1520) <= (layer1_outputs(2716)) or (layer1_outputs(11));
    layer2_outputs(1521) <= not((layer1_outputs(663)) or (layer1_outputs(546)));
    layer2_outputs(1522) <= not((layer1_outputs(3281)) or (layer1_outputs(1868)));
    layer2_outputs(1523) <= (layer1_outputs(4406)) and not (layer1_outputs(4671));
    layer2_outputs(1524) <= layer1_outputs(1916);
    layer2_outputs(1525) <= not(layer1_outputs(1611));
    layer2_outputs(1526) <= (layer1_outputs(804)) xor (layer1_outputs(421));
    layer2_outputs(1527) <= not((layer1_outputs(934)) and (layer1_outputs(235)));
    layer2_outputs(1528) <= layer1_outputs(3331);
    layer2_outputs(1529) <= not((layer1_outputs(2563)) or (layer1_outputs(2265)));
    layer2_outputs(1530) <= not(layer1_outputs(1927)) or (layer1_outputs(2843));
    layer2_outputs(1531) <= (layer1_outputs(1606)) and (layer1_outputs(771));
    layer2_outputs(1532) <= (layer1_outputs(3711)) xor (layer1_outputs(3766));
    layer2_outputs(1533) <= not(layer1_outputs(266)) or (layer1_outputs(3157));
    layer2_outputs(1534) <= layer1_outputs(4141);
    layer2_outputs(1535) <= not(layer1_outputs(3537));
    layer2_outputs(1536) <= layer1_outputs(3312);
    layer2_outputs(1537) <= not(layer1_outputs(4043));
    layer2_outputs(1538) <= not((layer1_outputs(743)) and (layer1_outputs(941)));
    layer2_outputs(1539) <= '0';
    layer2_outputs(1540) <= not((layer1_outputs(1341)) and (layer1_outputs(4680)));
    layer2_outputs(1541) <= not(layer1_outputs(5048)) or (layer1_outputs(4755));
    layer2_outputs(1542) <= not(layer1_outputs(551)) or (layer1_outputs(146));
    layer2_outputs(1543) <= not(layer1_outputs(4438)) or (layer1_outputs(2032));
    layer2_outputs(1544) <= not(layer1_outputs(4538)) or (layer1_outputs(233));
    layer2_outputs(1545) <= (layer1_outputs(1815)) and not (layer1_outputs(2145));
    layer2_outputs(1546) <= layer1_outputs(665);
    layer2_outputs(1547) <= not((layer1_outputs(4541)) xor (layer1_outputs(4984)));
    layer2_outputs(1548) <= (layer1_outputs(2884)) and not (layer1_outputs(1402));
    layer2_outputs(1549) <= not((layer1_outputs(4258)) and (layer1_outputs(800)));
    layer2_outputs(1550) <= not(layer1_outputs(1321));
    layer2_outputs(1551) <= not(layer1_outputs(1600));
    layer2_outputs(1552) <= (layer1_outputs(2585)) or (layer1_outputs(63));
    layer2_outputs(1553) <= not((layer1_outputs(1801)) xor (layer1_outputs(2201)));
    layer2_outputs(1554) <= not(layer1_outputs(3974));
    layer2_outputs(1555) <= layer1_outputs(2802);
    layer2_outputs(1556) <= (layer1_outputs(2744)) and (layer1_outputs(4720));
    layer2_outputs(1557) <= layer1_outputs(4952);
    layer2_outputs(1558) <= not(layer1_outputs(4949));
    layer2_outputs(1559) <= (layer1_outputs(1809)) and not (layer1_outputs(3842));
    layer2_outputs(1560) <= not(layer1_outputs(2348)) or (layer1_outputs(2723));
    layer2_outputs(1561) <= (layer1_outputs(1800)) and not (layer1_outputs(5098));
    layer2_outputs(1562) <= layer1_outputs(2964);
    layer2_outputs(1563) <= '1';
    layer2_outputs(1564) <= not(layer1_outputs(195));
    layer2_outputs(1565) <= not(layer1_outputs(3810));
    layer2_outputs(1566) <= not(layer1_outputs(404));
    layer2_outputs(1567) <= layer1_outputs(3030);
    layer2_outputs(1568) <= layer1_outputs(5003);
    layer2_outputs(1569) <= not(layer1_outputs(3920));
    layer2_outputs(1570) <= (layer1_outputs(3536)) and not (layer1_outputs(4132));
    layer2_outputs(1571) <= (layer1_outputs(293)) and not (layer1_outputs(4542));
    layer2_outputs(1572) <= not(layer1_outputs(4396)) or (layer1_outputs(2816));
    layer2_outputs(1573) <= (layer1_outputs(2613)) xor (layer1_outputs(2136));
    layer2_outputs(1574) <= not(layer1_outputs(2743));
    layer2_outputs(1575) <= not(layer1_outputs(2389));
    layer2_outputs(1576) <= not(layer1_outputs(1983)) or (layer1_outputs(4164));
    layer2_outputs(1577) <= not(layer1_outputs(4687)) or (layer1_outputs(4262));
    layer2_outputs(1578) <= not(layer1_outputs(2287));
    layer2_outputs(1579) <= not(layer1_outputs(3984));
    layer2_outputs(1580) <= layer1_outputs(468);
    layer2_outputs(1581) <= layer1_outputs(4630);
    layer2_outputs(1582) <= layer1_outputs(4089);
    layer2_outputs(1583) <= (layer1_outputs(1266)) xor (layer1_outputs(71));
    layer2_outputs(1584) <= not((layer1_outputs(1719)) or (layer1_outputs(496)));
    layer2_outputs(1585) <= not((layer1_outputs(3883)) and (layer1_outputs(1039)));
    layer2_outputs(1586) <= not(layer1_outputs(873)) or (layer1_outputs(4249));
    layer2_outputs(1587) <= layer1_outputs(2564);
    layer2_outputs(1588) <= not((layer1_outputs(544)) and (layer1_outputs(967)));
    layer2_outputs(1589) <= (layer1_outputs(2415)) and not (layer1_outputs(3456));
    layer2_outputs(1590) <= (layer1_outputs(2533)) and not (layer1_outputs(1757));
    layer2_outputs(1591) <= not(layer1_outputs(4455));
    layer2_outputs(1592) <= (layer1_outputs(3747)) and not (layer1_outputs(2262));
    layer2_outputs(1593) <= layer1_outputs(2314);
    layer2_outputs(1594) <= layer1_outputs(3485);
    layer2_outputs(1595) <= layer1_outputs(3993);
    layer2_outputs(1596) <= (layer1_outputs(2827)) and not (layer1_outputs(2819));
    layer2_outputs(1597) <= (layer1_outputs(2596)) and not (layer1_outputs(2226));
    layer2_outputs(1598) <= (layer1_outputs(1019)) xor (layer1_outputs(2528));
    layer2_outputs(1599) <= layer1_outputs(630);
    layer2_outputs(1600) <= not(layer1_outputs(4233)) or (layer1_outputs(1264));
    layer2_outputs(1601) <= layer1_outputs(49);
    layer2_outputs(1602) <= layer1_outputs(4490);
    layer2_outputs(1603) <= layer1_outputs(486);
    layer2_outputs(1604) <= layer1_outputs(2966);
    layer2_outputs(1605) <= (layer1_outputs(379)) and (layer1_outputs(3799));
    layer2_outputs(1606) <= not(layer1_outputs(2926)) or (layer1_outputs(3706));
    layer2_outputs(1607) <= not(layer1_outputs(1824));
    layer2_outputs(1608) <= not(layer1_outputs(2176));
    layer2_outputs(1609) <= layer1_outputs(2636);
    layer2_outputs(1610) <= layer1_outputs(1863);
    layer2_outputs(1611) <= (layer1_outputs(4774)) or (layer1_outputs(2760));
    layer2_outputs(1612) <= layer1_outputs(2943);
    layer2_outputs(1613) <= (layer1_outputs(3309)) and not (layer1_outputs(2561));
    layer2_outputs(1614) <= layer1_outputs(3260);
    layer2_outputs(1615) <= not(layer1_outputs(609));
    layer2_outputs(1616) <= layer1_outputs(3292);
    layer2_outputs(1617) <= (layer1_outputs(711)) xor (layer1_outputs(4132));
    layer2_outputs(1618) <= not(layer1_outputs(1482));
    layer2_outputs(1619) <= not(layer1_outputs(4723));
    layer2_outputs(1620) <= (layer1_outputs(3504)) and not (layer1_outputs(103));
    layer2_outputs(1621) <= layer1_outputs(3058);
    layer2_outputs(1622) <= not(layer1_outputs(3311));
    layer2_outputs(1623) <= layer1_outputs(4354);
    layer2_outputs(1624) <= '1';
    layer2_outputs(1625) <= layer1_outputs(2910);
    layer2_outputs(1626) <= not(layer1_outputs(3669));
    layer2_outputs(1627) <= '0';
    layer2_outputs(1628) <= not(layer1_outputs(4709));
    layer2_outputs(1629) <= (layer1_outputs(1262)) xor (layer1_outputs(643));
    layer2_outputs(1630) <= not(layer1_outputs(2480));
    layer2_outputs(1631) <= (layer1_outputs(425)) xor (layer1_outputs(1187));
    layer2_outputs(1632) <= (layer1_outputs(2446)) and (layer1_outputs(1349));
    layer2_outputs(1633) <= not((layer1_outputs(2114)) or (layer1_outputs(667)));
    layer2_outputs(1634) <= (layer1_outputs(3096)) and not (layer1_outputs(3817));
    layer2_outputs(1635) <= layer1_outputs(2363);
    layer2_outputs(1636) <= layer1_outputs(2353);
    layer2_outputs(1637) <= (layer1_outputs(2225)) or (layer1_outputs(4246));
    layer2_outputs(1638) <= layer1_outputs(3464);
    layer2_outputs(1639) <= not(layer1_outputs(2855)) or (layer1_outputs(2777));
    layer2_outputs(1640) <= layer1_outputs(93);
    layer2_outputs(1641) <= not((layer1_outputs(2600)) or (layer1_outputs(1929)));
    layer2_outputs(1642) <= (layer1_outputs(2700)) or (layer1_outputs(2092));
    layer2_outputs(1643) <= not(layer1_outputs(5065)) or (layer1_outputs(2171));
    layer2_outputs(1644) <= not(layer1_outputs(617)) or (layer1_outputs(33));
    layer2_outputs(1645) <= layer1_outputs(4549);
    layer2_outputs(1646) <= not(layer1_outputs(3879));
    layer2_outputs(1647) <= not((layer1_outputs(4650)) or (layer1_outputs(1759)));
    layer2_outputs(1648) <= not((layer1_outputs(1646)) and (layer1_outputs(16)));
    layer2_outputs(1649) <= not(layer1_outputs(2390));
    layer2_outputs(1650) <= layer1_outputs(1345);
    layer2_outputs(1651) <= not(layer1_outputs(3575));
    layer2_outputs(1652) <= not((layer1_outputs(1251)) and (layer1_outputs(3415)));
    layer2_outputs(1653) <= layer1_outputs(3946);
    layer2_outputs(1654) <= not(layer1_outputs(2202)) or (layer1_outputs(1179));
    layer2_outputs(1655) <= not((layer1_outputs(2620)) or (layer1_outputs(1576)));
    layer2_outputs(1656) <= not(layer1_outputs(1570));
    layer2_outputs(1657) <= (layer1_outputs(386)) or (layer1_outputs(1107));
    layer2_outputs(1658) <= layer1_outputs(628);
    layer2_outputs(1659) <= (layer1_outputs(5036)) xor (layer1_outputs(3754));
    layer2_outputs(1660) <= layer1_outputs(4641);
    layer2_outputs(1661) <= layer1_outputs(1573);
    layer2_outputs(1662) <= not(layer1_outputs(3730));
    layer2_outputs(1663) <= layer1_outputs(4421);
    layer2_outputs(1664) <= (layer1_outputs(2521)) and not (layer1_outputs(2683));
    layer2_outputs(1665) <= layer1_outputs(177);
    layer2_outputs(1666) <= not(layer1_outputs(1527));
    layer2_outputs(1667) <= layer1_outputs(3611);
    layer2_outputs(1668) <= not(layer1_outputs(4005));
    layer2_outputs(1669) <= (layer1_outputs(2253)) and not (layer1_outputs(339));
    layer2_outputs(1670) <= layer1_outputs(4681);
    layer2_outputs(1671) <= not(layer1_outputs(1317)) or (layer1_outputs(4319));
    layer2_outputs(1672) <= not(layer1_outputs(1985)) or (layer1_outputs(644));
    layer2_outputs(1673) <= layer1_outputs(3366);
    layer2_outputs(1674) <= not((layer1_outputs(1983)) and (layer1_outputs(3803)));
    layer2_outputs(1675) <= not((layer1_outputs(3016)) or (layer1_outputs(2243)));
    layer2_outputs(1676) <= layer1_outputs(1618);
    layer2_outputs(1677) <= layer1_outputs(3294);
    layer2_outputs(1678) <= (layer1_outputs(3465)) and not (layer1_outputs(1398));
    layer2_outputs(1679) <= layer1_outputs(4570);
    layer2_outputs(1680) <= not(layer1_outputs(1267));
    layer2_outputs(1681) <= not(layer1_outputs(673));
    layer2_outputs(1682) <= not(layer1_outputs(1937));
    layer2_outputs(1683) <= not(layer1_outputs(3949));
    layer2_outputs(1684) <= not(layer1_outputs(92));
    layer2_outputs(1685) <= (layer1_outputs(938)) or (layer1_outputs(745));
    layer2_outputs(1686) <= layer1_outputs(2011);
    layer2_outputs(1687) <= not((layer1_outputs(2920)) and (layer1_outputs(2460)));
    layer2_outputs(1688) <= layer1_outputs(4946);
    layer2_outputs(1689) <= not(layer1_outputs(4199)) or (layer1_outputs(874));
    layer2_outputs(1690) <= layer1_outputs(388);
    layer2_outputs(1691) <= '1';
    layer2_outputs(1692) <= not(layer1_outputs(3800));
    layer2_outputs(1693) <= layer1_outputs(4941);
    layer2_outputs(1694) <= not((layer1_outputs(2159)) or (layer1_outputs(4077)));
    layer2_outputs(1695) <= (layer1_outputs(3048)) or (layer1_outputs(2018));
    layer2_outputs(1696) <= not((layer1_outputs(1642)) or (layer1_outputs(3553)));
    layer2_outputs(1697) <= not(layer1_outputs(1528)) or (layer1_outputs(2674));
    layer2_outputs(1698) <= (layer1_outputs(1526)) or (layer1_outputs(1033));
    layer2_outputs(1699) <= layer1_outputs(3639);
    layer2_outputs(1700) <= not(layer1_outputs(2773));
    layer2_outputs(1701) <= not((layer1_outputs(4613)) or (layer1_outputs(1277)));
    layer2_outputs(1702) <= not((layer1_outputs(2305)) xor (layer1_outputs(2389)));
    layer2_outputs(1703) <= not((layer1_outputs(1140)) or (layer1_outputs(812)));
    layer2_outputs(1704) <= layer1_outputs(2274);
    layer2_outputs(1705) <= (layer1_outputs(4705)) or (layer1_outputs(1135));
    layer2_outputs(1706) <= (layer1_outputs(2145)) and not (layer1_outputs(1984));
    layer2_outputs(1707) <= '0';
    layer2_outputs(1708) <= (layer1_outputs(4609)) and not (layer1_outputs(2452));
    layer2_outputs(1709) <= not((layer1_outputs(961)) and (layer1_outputs(1543)));
    layer2_outputs(1710) <= layer1_outputs(1924);
    layer2_outputs(1711) <= layer1_outputs(5059);
    layer2_outputs(1712) <= not(layer1_outputs(4281));
    layer2_outputs(1713) <= layer1_outputs(2960);
    layer2_outputs(1714) <= (layer1_outputs(647)) or (layer1_outputs(439));
    layer2_outputs(1715) <= layer1_outputs(4093);
    layer2_outputs(1716) <= (layer1_outputs(3044)) or (layer1_outputs(4717));
    layer2_outputs(1717) <= not(layer1_outputs(3483));
    layer2_outputs(1718) <= (layer1_outputs(3902)) and not (layer1_outputs(2291));
    layer2_outputs(1719) <= not((layer1_outputs(4789)) xor (layer1_outputs(4243)));
    layer2_outputs(1720) <= not((layer1_outputs(1016)) or (layer1_outputs(1609)));
    layer2_outputs(1721) <= not(layer1_outputs(3226)) or (layer1_outputs(3447));
    layer2_outputs(1722) <= not(layer1_outputs(639));
    layer2_outputs(1723) <= layer1_outputs(4529);
    layer2_outputs(1724) <= not(layer1_outputs(3094)) or (layer1_outputs(2850));
    layer2_outputs(1725) <= layer1_outputs(4516);
    layer2_outputs(1726) <= not(layer1_outputs(2229)) or (layer1_outputs(3036));
    layer2_outputs(1727) <= layer1_outputs(4737);
    layer2_outputs(1728) <= not(layer1_outputs(2475)) or (layer1_outputs(3525));
    layer2_outputs(1729) <= not(layer1_outputs(2552));
    layer2_outputs(1730) <= not((layer1_outputs(885)) and (layer1_outputs(3369)));
    layer2_outputs(1731) <= not((layer1_outputs(465)) or (layer1_outputs(3976)));
    layer2_outputs(1732) <= not(layer1_outputs(1040)) or (layer1_outputs(2810));
    layer2_outputs(1733) <= (layer1_outputs(3216)) xor (layer1_outputs(182));
    layer2_outputs(1734) <= not((layer1_outputs(4946)) and (layer1_outputs(1399)));
    layer2_outputs(1735) <= not(layer1_outputs(2561));
    layer2_outputs(1736) <= layer1_outputs(3454);
    layer2_outputs(1737) <= (layer1_outputs(833)) and not (layer1_outputs(2725));
    layer2_outputs(1738) <= not(layer1_outputs(1324)) or (layer1_outputs(4176));
    layer2_outputs(1739) <= not(layer1_outputs(3843)) or (layer1_outputs(2197));
    layer2_outputs(1740) <= not(layer1_outputs(2851));
    layer2_outputs(1741) <= (layer1_outputs(706)) xor (layer1_outputs(4506));
    layer2_outputs(1742) <= not((layer1_outputs(2361)) xor (layer1_outputs(3080)));
    layer2_outputs(1743) <= layer1_outputs(234);
    layer2_outputs(1744) <= layer1_outputs(622);
    layer2_outputs(1745) <= (layer1_outputs(3140)) and (layer1_outputs(292));
    layer2_outputs(1746) <= layer1_outputs(4097);
    layer2_outputs(1747) <= (layer1_outputs(4235)) and not (layer1_outputs(4296));
    layer2_outputs(1748) <= not(layer1_outputs(4847)) or (layer1_outputs(1725));
    layer2_outputs(1749) <= (layer1_outputs(4858)) or (layer1_outputs(4557));
    layer2_outputs(1750) <= not(layer1_outputs(3562));
    layer2_outputs(1751) <= not(layer1_outputs(4791)) or (layer1_outputs(3076));
    layer2_outputs(1752) <= not(layer1_outputs(3950)) or (layer1_outputs(3961));
    layer2_outputs(1753) <= not((layer1_outputs(3718)) or (layer1_outputs(1489)));
    layer2_outputs(1754) <= not(layer1_outputs(2404)) or (layer1_outputs(3592));
    layer2_outputs(1755) <= layer1_outputs(703);
    layer2_outputs(1756) <= not((layer1_outputs(669)) xor (layer1_outputs(1937)));
    layer2_outputs(1757) <= not(layer1_outputs(1777)) or (layer1_outputs(3180));
    layer2_outputs(1758) <= (layer1_outputs(3912)) xor (layer1_outputs(1950));
    layer2_outputs(1759) <= not((layer1_outputs(4863)) or (layer1_outputs(3007)));
    layer2_outputs(1760) <= not(layer1_outputs(3752));
    layer2_outputs(1761) <= (layer1_outputs(3772)) or (layer1_outputs(4291));
    layer2_outputs(1762) <= (layer1_outputs(2892)) and (layer1_outputs(2523));
    layer2_outputs(1763) <= (layer1_outputs(2580)) and (layer1_outputs(3862));
    layer2_outputs(1764) <= (layer1_outputs(2856)) and not (layer1_outputs(1495));
    layer2_outputs(1765) <= not((layer1_outputs(4344)) xor (layer1_outputs(2737)));
    layer2_outputs(1766) <= not(layer1_outputs(4100)) or (layer1_outputs(3122));
    layer2_outputs(1767) <= not(layer1_outputs(4556));
    layer2_outputs(1768) <= (layer1_outputs(2531)) and not (layer1_outputs(3405));
    layer2_outputs(1769) <= not((layer1_outputs(1485)) or (layer1_outputs(2724)));
    layer2_outputs(1770) <= (layer1_outputs(1473)) or (layer1_outputs(1819));
    layer2_outputs(1771) <= layer1_outputs(1863);
    layer2_outputs(1772) <= layer1_outputs(1924);
    layer2_outputs(1773) <= (layer1_outputs(4787)) and (layer1_outputs(5041));
    layer2_outputs(1774) <= not(layer1_outputs(2063));
    layer2_outputs(1775) <= not(layer1_outputs(455));
    layer2_outputs(1776) <= not(layer1_outputs(451));
    layer2_outputs(1777) <= not(layer1_outputs(4273));
    layer2_outputs(1778) <= layer1_outputs(282);
    layer2_outputs(1779) <= not(layer1_outputs(5116));
    layer2_outputs(1780) <= '0';
    layer2_outputs(1781) <= (layer1_outputs(4222)) and not (layer1_outputs(3053));
    layer2_outputs(1782) <= (layer1_outputs(5007)) or (layer1_outputs(300));
    layer2_outputs(1783) <= layer1_outputs(2548);
    layer2_outputs(1784) <= not((layer1_outputs(3382)) or (layer1_outputs(4587)));
    layer2_outputs(1785) <= not((layer1_outputs(3172)) or (layer1_outputs(1915)));
    layer2_outputs(1786) <= layer1_outputs(3543);
    layer2_outputs(1787) <= not(layer1_outputs(211)) or (layer1_outputs(3143));
    layer2_outputs(1788) <= not(layer1_outputs(1013));
    layer2_outputs(1789) <= not(layer1_outputs(2043));
    layer2_outputs(1790) <= (layer1_outputs(3231)) and not (layer1_outputs(2330));
    layer2_outputs(1791) <= (layer1_outputs(4496)) xor (layer1_outputs(4332));
    layer2_outputs(1792) <= '1';
    layer2_outputs(1793) <= (layer1_outputs(4034)) and (layer1_outputs(580));
    layer2_outputs(1794) <= layer1_outputs(1833);
    layer2_outputs(1795) <= layer1_outputs(166);
    layer2_outputs(1796) <= not((layer1_outputs(2628)) and (layer1_outputs(875)));
    layer2_outputs(1797) <= (layer1_outputs(2143)) or (layer1_outputs(604));
    layer2_outputs(1798) <= not(layer1_outputs(4950)) or (layer1_outputs(490));
    layer2_outputs(1799) <= not(layer1_outputs(52));
    layer2_outputs(1800) <= (layer1_outputs(3517)) xor (layer1_outputs(4513));
    layer2_outputs(1801) <= not((layer1_outputs(2813)) or (layer1_outputs(81)));
    layer2_outputs(1802) <= not((layer1_outputs(943)) xor (layer1_outputs(769)));
    layer2_outputs(1803) <= not(layer1_outputs(1015));
    layer2_outputs(1804) <= not(layer1_outputs(1958)) or (layer1_outputs(1537));
    layer2_outputs(1805) <= not(layer1_outputs(2397));
    layer2_outputs(1806) <= not(layer1_outputs(1339));
    layer2_outputs(1807) <= (layer1_outputs(2493)) and not (layer1_outputs(3084));
    layer2_outputs(1808) <= layer1_outputs(1929);
    layer2_outputs(1809) <= layer1_outputs(4512);
    layer2_outputs(1810) <= (layer1_outputs(3583)) and (layer1_outputs(1767));
    layer2_outputs(1811) <= (layer1_outputs(1387)) xor (layer1_outputs(4297));
    layer2_outputs(1812) <= (layer1_outputs(909)) and (layer1_outputs(1063));
    layer2_outputs(1813) <= not(layer1_outputs(3134));
    layer2_outputs(1814) <= not(layer1_outputs(938));
    layer2_outputs(1815) <= (layer1_outputs(434)) and (layer1_outputs(3236));
    layer2_outputs(1816) <= not(layer1_outputs(4646));
    layer2_outputs(1817) <= (layer1_outputs(880)) or (layer1_outputs(1026));
    layer2_outputs(1818) <= layer1_outputs(1857);
    layer2_outputs(1819) <= layer1_outputs(535);
    layer2_outputs(1820) <= layer1_outputs(487);
    layer2_outputs(1821) <= layer1_outputs(4924);
    layer2_outputs(1822) <= not((layer1_outputs(4165)) xor (layer1_outputs(1638)));
    layer2_outputs(1823) <= layer1_outputs(3444);
    layer2_outputs(1824) <= layer1_outputs(3127);
    layer2_outputs(1825) <= '1';
    layer2_outputs(1826) <= (layer1_outputs(2659)) or (layer1_outputs(842));
    layer2_outputs(1827) <= layer1_outputs(4465);
    layer2_outputs(1828) <= not((layer1_outputs(2222)) and (layer1_outputs(5049)));
    layer2_outputs(1829) <= layer1_outputs(2650);
    layer2_outputs(1830) <= not((layer1_outputs(3262)) and (layer1_outputs(4404)));
    layer2_outputs(1831) <= layer1_outputs(2439);
    layer2_outputs(1832) <= (layer1_outputs(1711)) and (layer1_outputs(1188));
    layer2_outputs(1833) <= layer1_outputs(3918);
    layer2_outputs(1834) <= not(layer1_outputs(4849));
    layer2_outputs(1835) <= (layer1_outputs(4261)) and (layer1_outputs(1293));
    layer2_outputs(1836) <= layer1_outputs(294);
    layer2_outputs(1837) <= (layer1_outputs(802)) or (layer1_outputs(3484));
    layer2_outputs(1838) <= not(layer1_outputs(3243));
    layer2_outputs(1839) <= (layer1_outputs(2990)) xor (layer1_outputs(1491));
    layer2_outputs(1840) <= not((layer1_outputs(1972)) xor (layer1_outputs(2793)));
    layer2_outputs(1841) <= (layer1_outputs(4226)) and (layer1_outputs(2510));
    layer2_outputs(1842) <= not(layer1_outputs(3949));
    layer2_outputs(1843) <= not(layer1_outputs(621));
    layer2_outputs(1844) <= not(layer1_outputs(3427));
    layer2_outputs(1845) <= layer1_outputs(110);
    layer2_outputs(1846) <= not(layer1_outputs(1115));
    layer2_outputs(1847) <= layer1_outputs(2526);
    layer2_outputs(1848) <= not(layer1_outputs(2574));
    layer2_outputs(1849) <= not(layer1_outputs(3712));
    layer2_outputs(1850) <= not(layer1_outputs(717));
    layer2_outputs(1851) <= (layer1_outputs(808)) xor (layer1_outputs(1376));
    layer2_outputs(1852) <= not(layer1_outputs(2917));
    layer2_outputs(1853) <= not((layer1_outputs(4900)) xor (layer1_outputs(445)));
    layer2_outputs(1854) <= not((layer1_outputs(1812)) or (layer1_outputs(4003)));
    layer2_outputs(1855) <= layer1_outputs(3065);
    layer2_outputs(1856) <= (layer1_outputs(563)) or (layer1_outputs(1377));
    layer2_outputs(1857) <= not((layer1_outputs(3833)) xor (layer1_outputs(2059)));
    layer2_outputs(1858) <= layer1_outputs(2403);
    layer2_outputs(1859) <= not(layer1_outputs(897));
    layer2_outputs(1860) <= (layer1_outputs(2539)) or (layer1_outputs(4381));
    layer2_outputs(1861) <= not(layer1_outputs(3065));
    layer2_outputs(1862) <= (layer1_outputs(2641)) and not (layer1_outputs(1949));
    layer2_outputs(1863) <= layer1_outputs(1842);
    layer2_outputs(1864) <= not((layer1_outputs(190)) or (layer1_outputs(2601)));
    layer2_outputs(1865) <= layer1_outputs(3379);
    layer2_outputs(1866) <= not(layer1_outputs(999)) or (layer1_outputs(4086));
    layer2_outputs(1867) <= layer1_outputs(794);
    layer2_outputs(1868) <= not((layer1_outputs(2912)) xor (layer1_outputs(2272)));
    layer2_outputs(1869) <= not(layer1_outputs(172));
    layer2_outputs(1870) <= layer1_outputs(2784);
    layer2_outputs(1871) <= not((layer1_outputs(2365)) or (layer1_outputs(4011)));
    layer2_outputs(1872) <= (layer1_outputs(3718)) and (layer1_outputs(272));
    layer2_outputs(1873) <= (layer1_outputs(4575)) and not (layer1_outputs(3072));
    layer2_outputs(1874) <= not((layer1_outputs(3251)) and (layer1_outputs(2567)));
    layer2_outputs(1875) <= not((layer1_outputs(402)) xor (layer1_outputs(4811)));
    layer2_outputs(1876) <= (layer1_outputs(1754)) and (layer1_outputs(3252));
    layer2_outputs(1877) <= not((layer1_outputs(4111)) xor (layer1_outputs(108)));
    layer2_outputs(1878) <= layer1_outputs(503);
    layer2_outputs(1879) <= not((layer1_outputs(916)) or (layer1_outputs(1892)));
    layer2_outputs(1880) <= not((layer1_outputs(2803)) or (layer1_outputs(4098)));
    layer2_outputs(1881) <= layer1_outputs(1680);
    layer2_outputs(1882) <= (layer1_outputs(4272)) xor (layer1_outputs(555));
    layer2_outputs(1883) <= (layer1_outputs(3698)) and not (layer1_outputs(543));
    layer2_outputs(1884) <= not((layer1_outputs(3136)) and (layer1_outputs(2153)));
    layer2_outputs(1885) <= (layer1_outputs(2824)) xor (layer1_outputs(4533));
    layer2_outputs(1886) <= layer1_outputs(4328);
    layer2_outputs(1887) <= not(layer1_outputs(4859));
    layer2_outputs(1888) <= layer1_outputs(3217);
    layer2_outputs(1889) <= not((layer1_outputs(2718)) or (layer1_outputs(143)));
    layer2_outputs(1890) <= not(layer1_outputs(4682)) or (layer1_outputs(4063));
    layer2_outputs(1891) <= (layer1_outputs(2301)) and not (layer1_outputs(494));
    layer2_outputs(1892) <= (layer1_outputs(920)) xor (layer1_outputs(1607));
    layer2_outputs(1893) <= not(layer1_outputs(3820)) or (layer1_outputs(5106));
    layer2_outputs(1894) <= not(layer1_outputs(5005));
    layer2_outputs(1895) <= (layer1_outputs(147)) and (layer1_outputs(3786));
    layer2_outputs(1896) <= (layer1_outputs(3252)) and not (layer1_outputs(4530));
    layer2_outputs(1897) <= layer1_outputs(1944);
    layer2_outputs(1898) <= layer1_outputs(392);
    layer2_outputs(1899) <= not((layer1_outputs(4303)) and (layer1_outputs(1903)));
    layer2_outputs(1900) <= not((layer1_outputs(988)) or (layer1_outputs(4639)));
    layer2_outputs(1901) <= (layer1_outputs(112)) xor (layer1_outputs(4348));
    layer2_outputs(1902) <= (layer1_outputs(2996)) or (layer1_outputs(627));
    layer2_outputs(1903) <= (layer1_outputs(3568)) or (layer1_outputs(2194));
    layer2_outputs(1904) <= not(layer1_outputs(4683)) or (layer1_outputs(2081));
    layer2_outputs(1905) <= (layer1_outputs(3045)) xor (layer1_outputs(3682));
    layer2_outputs(1906) <= not(layer1_outputs(179));
    layer2_outputs(1907) <= not((layer1_outputs(1314)) or (layer1_outputs(2288)));
    layer2_outputs(1908) <= layer1_outputs(3869);
    layer2_outputs(1909) <= not((layer1_outputs(4973)) xor (layer1_outputs(126)));
    layer2_outputs(1910) <= not(layer1_outputs(1856));
    layer2_outputs(1911) <= '1';
    layer2_outputs(1912) <= not(layer1_outputs(4795));
    layer2_outputs(1913) <= layer1_outputs(4273);
    layer2_outputs(1914) <= layer1_outputs(4391);
    layer2_outputs(1915) <= layer1_outputs(114);
    layer2_outputs(1916) <= layer1_outputs(524);
    layer2_outputs(1917) <= (layer1_outputs(514)) xor (layer1_outputs(2150));
    layer2_outputs(1918) <= not(layer1_outputs(965));
    layer2_outputs(1919) <= layer1_outputs(98);
    layer2_outputs(1920) <= not((layer1_outputs(581)) or (layer1_outputs(498)));
    layer2_outputs(1921) <= layer1_outputs(2044);
    layer2_outputs(1922) <= not(layer1_outputs(192));
    layer2_outputs(1923) <= not(layer1_outputs(3578));
    layer2_outputs(1924) <= (layer1_outputs(24)) and (layer1_outputs(3742));
    layer2_outputs(1925) <= not((layer1_outputs(4322)) xor (layer1_outputs(1333)));
    layer2_outputs(1926) <= layer1_outputs(3387);
    layer2_outputs(1927) <= not((layer1_outputs(2953)) or (layer1_outputs(3641)));
    layer2_outputs(1928) <= layer1_outputs(1083);
    layer2_outputs(1929) <= not((layer1_outputs(1020)) or (layer1_outputs(3527)));
    layer2_outputs(1930) <= not(layer1_outputs(2606));
    layer2_outputs(1931) <= not(layer1_outputs(3783));
    layer2_outputs(1932) <= layer1_outputs(3978);
    layer2_outputs(1933) <= (layer1_outputs(2867)) or (layer1_outputs(314));
    layer2_outputs(1934) <= not((layer1_outputs(1190)) xor (layer1_outputs(4163)));
    layer2_outputs(1935) <= layer1_outputs(256);
    layer2_outputs(1936) <= not(layer1_outputs(1855)) or (layer1_outputs(451));
    layer2_outputs(1937) <= not((layer1_outputs(4834)) xor (layer1_outputs(4642)));
    layer2_outputs(1938) <= not(layer1_outputs(4764)) or (layer1_outputs(1296));
    layer2_outputs(1939) <= not((layer1_outputs(5088)) xor (layer1_outputs(2895)));
    layer2_outputs(1940) <= (layer1_outputs(2534)) and not (layer1_outputs(4796));
    layer2_outputs(1941) <= (layer1_outputs(2989)) and (layer1_outputs(1319));
    layer2_outputs(1942) <= not(layer1_outputs(1268)) or (layer1_outputs(682));
    layer2_outputs(1943) <= not((layer1_outputs(3641)) xor (layer1_outputs(3907)));
    layer2_outputs(1944) <= (layer1_outputs(3977)) or (layer1_outputs(5060));
    layer2_outputs(1945) <= layer1_outputs(4469);
    layer2_outputs(1946) <= not(layer1_outputs(3651));
    layer2_outputs(1947) <= (layer1_outputs(4174)) or (layer1_outputs(4902));
    layer2_outputs(1948) <= not(layer1_outputs(3625)) or (layer1_outputs(4230));
    layer2_outputs(1949) <= not(layer1_outputs(3550));
    layer2_outputs(1950) <= not(layer1_outputs(2625));
    layer2_outputs(1951) <= (layer1_outputs(2088)) xor (layer1_outputs(1418));
    layer2_outputs(1952) <= not(layer1_outputs(2234));
    layer2_outputs(1953) <= not((layer1_outputs(707)) xor (layer1_outputs(4562)));
    layer2_outputs(1954) <= not(layer1_outputs(2248));
    layer2_outputs(1955) <= '0';
    layer2_outputs(1956) <= not(layer1_outputs(789));
    layer2_outputs(1957) <= layer1_outputs(415);
    layer2_outputs(1958) <= not((layer1_outputs(3960)) and (layer1_outputs(2906)));
    layer2_outputs(1959) <= layer1_outputs(125);
    layer2_outputs(1960) <= not((layer1_outputs(85)) and (layer1_outputs(2699)));
    layer2_outputs(1961) <= layer1_outputs(1201);
    layer2_outputs(1962) <= (layer1_outputs(3140)) xor (layer1_outputs(1357));
    layer2_outputs(1963) <= not(layer1_outputs(1928));
    layer2_outputs(1964) <= (layer1_outputs(2364)) and (layer1_outputs(156));
    layer2_outputs(1965) <= (layer1_outputs(1867)) xor (layer1_outputs(540));
    layer2_outputs(1966) <= not(layer1_outputs(4293));
    layer2_outputs(1967) <= '0';
    layer2_outputs(1968) <= not(layer1_outputs(4958));
    layer2_outputs(1969) <= not((layer1_outputs(145)) xor (layer1_outputs(4593)));
    layer2_outputs(1970) <= not(layer1_outputs(2939));
    layer2_outputs(1971) <= not(layer1_outputs(4171)) or (layer1_outputs(3779));
    layer2_outputs(1972) <= layer1_outputs(4635);
    layer2_outputs(1973) <= layer1_outputs(1035);
    layer2_outputs(1974) <= not(layer1_outputs(3609));
    layer2_outputs(1975) <= not((layer1_outputs(607)) and (layer1_outputs(4440)));
    layer2_outputs(1976) <= (layer1_outputs(1389)) and not (layer1_outputs(1021));
    layer2_outputs(1977) <= layer1_outputs(3715);
    layer2_outputs(1978) <= (layer1_outputs(2898)) and not (layer1_outputs(2006));
    layer2_outputs(1979) <= (layer1_outputs(1805)) or (layer1_outputs(1667));
    layer2_outputs(1980) <= (layer1_outputs(1257)) xor (layer1_outputs(683));
    layer2_outputs(1981) <= not(layer1_outputs(188));
    layer2_outputs(1982) <= not(layer1_outputs(585));
    layer2_outputs(1983) <= not(layer1_outputs(2435)) or (layer1_outputs(5110));
    layer2_outputs(1984) <= not(layer1_outputs(5030));
    layer2_outputs(1985) <= not(layer1_outputs(3214)) or (layer1_outputs(1563));
    layer2_outputs(1986) <= not(layer1_outputs(4996));
    layer2_outputs(1987) <= (layer1_outputs(3786)) and not (layer1_outputs(4743));
    layer2_outputs(1988) <= not(layer1_outputs(4440));
    layer2_outputs(1989) <= not(layer1_outputs(4397));
    layer2_outputs(1990) <= not((layer1_outputs(433)) and (layer1_outputs(826)));
    layer2_outputs(1991) <= not((layer1_outputs(4313)) or (layer1_outputs(1285)));
    layer2_outputs(1992) <= layer1_outputs(284);
    layer2_outputs(1993) <= not(layer1_outputs(2845)) or (layer1_outputs(1917));
    layer2_outputs(1994) <= not(layer1_outputs(2459));
    layer2_outputs(1995) <= not((layer1_outputs(4963)) or (layer1_outputs(3429)));
    layer2_outputs(1996) <= not(layer1_outputs(1504));
    layer2_outputs(1997) <= (layer1_outputs(4326)) and not (layer1_outputs(1699));
    layer2_outputs(1998) <= layer1_outputs(3035);
    layer2_outputs(1999) <= (layer1_outputs(2406)) or (layer1_outputs(934));
    layer2_outputs(2000) <= not((layer1_outputs(3109)) and (layer1_outputs(2974)));
    layer2_outputs(2001) <= layer1_outputs(3162);
    layer2_outputs(2002) <= not(layer1_outputs(1848));
    layer2_outputs(2003) <= (layer1_outputs(1431)) xor (layer1_outputs(4197));
    layer2_outputs(2004) <= not(layer1_outputs(1705)) or (layer1_outputs(2397));
    layer2_outputs(2005) <= layer1_outputs(2655);
    layer2_outputs(2006) <= not(layer1_outputs(3114));
    layer2_outputs(2007) <= not(layer1_outputs(2526));
    layer2_outputs(2008) <= not(layer1_outputs(3290));
    layer2_outputs(2009) <= not(layer1_outputs(4343));
    layer2_outputs(2010) <= (layer1_outputs(2869)) or (layer1_outputs(1099));
    layer2_outputs(2011) <= not(layer1_outputs(2065));
    layer2_outputs(2012) <= (layer1_outputs(525)) or (layer1_outputs(4896));
    layer2_outputs(2013) <= not((layer1_outputs(4223)) xor (layer1_outputs(3111)));
    layer2_outputs(2014) <= not((layer1_outputs(4563)) and (layer1_outputs(4050)));
    layer2_outputs(2015) <= not(layer1_outputs(4402));
    layer2_outputs(2016) <= not(layer1_outputs(3426));
    layer2_outputs(2017) <= layer1_outputs(386);
    layer2_outputs(2018) <= not(layer1_outputs(1633));
    layer2_outputs(2019) <= layer1_outputs(3722);
    layer2_outputs(2020) <= '1';
    layer2_outputs(2021) <= not((layer1_outputs(1994)) xor (layer1_outputs(4339)));
    layer2_outputs(2022) <= (layer1_outputs(4436)) and (layer1_outputs(933));
    layer2_outputs(2023) <= layer1_outputs(3346);
    layer2_outputs(2024) <= (layer1_outputs(5094)) and not (layer1_outputs(3849));
    layer2_outputs(2025) <= not(layer1_outputs(3542));
    layer2_outputs(2026) <= not(layer1_outputs(3000)) or (layer1_outputs(866));
    layer2_outputs(2027) <= layer1_outputs(3206);
    layer2_outputs(2028) <= (layer1_outputs(3636)) xor (layer1_outputs(3308));
    layer2_outputs(2029) <= not((layer1_outputs(670)) or (layer1_outputs(2209)));
    layer2_outputs(2030) <= (layer1_outputs(3940)) and not (layer1_outputs(326));
    layer2_outputs(2031) <= not(layer1_outputs(2297));
    layer2_outputs(2032) <= not(layer1_outputs(2615));
    layer2_outputs(2033) <= not(layer1_outputs(44)) or (layer1_outputs(3599));
    layer2_outputs(2034) <= layer1_outputs(188);
    layer2_outputs(2035) <= (layer1_outputs(2586)) and not (layer1_outputs(3254));
    layer2_outputs(2036) <= (layer1_outputs(2422)) and not (layer1_outputs(865));
    layer2_outputs(2037) <= not(layer1_outputs(4969)) or (layer1_outputs(773));
    layer2_outputs(2038) <= (layer1_outputs(3622)) and (layer1_outputs(868));
    layer2_outputs(2039) <= layer1_outputs(110);
    layer2_outputs(2040) <= not(layer1_outputs(4124)) or (layer1_outputs(3234));
    layer2_outputs(2041) <= layer1_outputs(1654);
    layer2_outputs(2042) <= not((layer1_outputs(1334)) or (layer1_outputs(1385)));
    layer2_outputs(2043) <= (layer1_outputs(1230)) and not (layer1_outputs(2570));
    layer2_outputs(2044) <= (layer1_outputs(136)) or (layer1_outputs(1217));
    layer2_outputs(2045) <= (layer1_outputs(1131)) and (layer1_outputs(4386));
    layer2_outputs(2046) <= not(layer1_outputs(1424));
    layer2_outputs(2047) <= layer1_outputs(3650);
    layer2_outputs(2048) <= (layer1_outputs(5089)) and not (layer1_outputs(4000));
    layer2_outputs(2049) <= not((layer1_outputs(2893)) xor (layer1_outputs(684)));
    layer2_outputs(2050) <= layer1_outputs(3601);
    layer2_outputs(2051) <= (layer1_outputs(1433)) xor (layer1_outputs(777));
    layer2_outputs(2052) <= not(layer1_outputs(3054)) or (layer1_outputs(13));
    layer2_outputs(2053) <= layer1_outputs(3904);
    layer2_outputs(2054) <= layer1_outputs(2418);
    layer2_outputs(2055) <= not((layer1_outputs(1775)) and (layer1_outputs(4014)));
    layer2_outputs(2056) <= not(layer1_outputs(423)) or (layer1_outputs(3942));
    layer2_outputs(2057) <= layer1_outputs(436);
    layer2_outputs(2058) <= not(layer1_outputs(580));
    layer2_outputs(2059) <= (layer1_outputs(2326)) xor (layer1_outputs(3323));
    layer2_outputs(2060) <= not((layer1_outputs(109)) xor (layer1_outputs(2565)));
    layer2_outputs(2061) <= not(layer1_outputs(1699));
    layer2_outputs(2062) <= layer1_outputs(1951);
    layer2_outputs(2063) <= not((layer1_outputs(1532)) xor (layer1_outputs(954)));
    layer2_outputs(2064) <= (layer1_outputs(4694)) and not (layer1_outputs(446));
    layer2_outputs(2065) <= (layer1_outputs(4241)) and not (layer1_outputs(4139));
    layer2_outputs(2066) <= (layer1_outputs(5089)) and not (layer1_outputs(1540));
    layer2_outputs(2067) <= not(layer1_outputs(3513));
    layer2_outputs(2068) <= not(layer1_outputs(2311));
    layer2_outputs(2069) <= not((layer1_outputs(4881)) or (layer1_outputs(2417)));
    layer2_outputs(2070) <= not((layer1_outputs(1143)) or (layer1_outputs(785)));
    layer2_outputs(2071) <= not((layer1_outputs(2782)) or (layer1_outputs(1789)));
    layer2_outputs(2072) <= (layer1_outputs(1320)) or (layer1_outputs(4974));
    layer2_outputs(2073) <= (layer1_outputs(1938)) and not (layer1_outputs(1435));
    layer2_outputs(2074) <= not(layer1_outputs(1999)) or (layer1_outputs(1908));
    layer2_outputs(2075) <= not(layer1_outputs(4350));
    layer2_outputs(2076) <= (layer1_outputs(3374)) or (layer1_outputs(1766));
    layer2_outputs(2077) <= not((layer1_outputs(2039)) or (layer1_outputs(2015)));
    layer2_outputs(2078) <= layer1_outputs(3916);
    layer2_outputs(2079) <= layer1_outputs(5099);
    layer2_outputs(2080) <= (layer1_outputs(1263)) and not (layer1_outputs(3636));
    layer2_outputs(2081) <= not(layer1_outputs(462));
    layer2_outputs(2082) <= (layer1_outputs(4546)) xor (layer1_outputs(1207));
    layer2_outputs(2083) <= not(layer1_outputs(1329)) or (layer1_outputs(1642));
    layer2_outputs(2084) <= (layer1_outputs(3861)) xor (layer1_outputs(5000));
    layer2_outputs(2085) <= not(layer1_outputs(3250));
    layer2_outputs(2086) <= (layer1_outputs(4322)) and (layer1_outputs(660));
    layer2_outputs(2087) <= (layer1_outputs(1472)) and not (layer1_outputs(1243));
    layer2_outputs(2088) <= not(layer1_outputs(1077));
    layer2_outputs(2089) <= not((layer1_outputs(623)) and (layer1_outputs(891)));
    layer2_outputs(2090) <= not(layer1_outputs(648));
    layer2_outputs(2091) <= (layer1_outputs(4060)) and not (layer1_outputs(3727));
    layer2_outputs(2092) <= not(layer1_outputs(2928));
    layer2_outputs(2093) <= layer1_outputs(1865);
    layer2_outputs(2094) <= layer1_outputs(460);
    layer2_outputs(2095) <= not((layer1_outputs(1195)) xor (layer1_outputs(4585)));
    layer2_outputs(2096) <= not(layer1_outputs(4218));
    layer2_outputs(2097) <= not(layer1_outputs(3861));
    layer2_outputs(2098) <= layer1_outputs(3695);
    layer2_outputs(2099) <= '1';
    layer2_outputs(2100) <= layer1_outputs(40);
    layer2_outputs(2101) <= not((layer1_outputs(2796)) xor (layer1_outputs(244)));
    layer2_outputs(2102) <= (layer1_outputs(4639)) xor (layer1_outputs(3222));
    layer2_outputs(2103) <= not(layer1_outputs(1568));
    layer2_outputs(2104) <= layer1_outputs(4724);
    layer2_outputs(2105) <= not(layer1_outputs(1534));
    layer2_outputs(2106) <= (layer1_outputs(4517)) and not (layer1_outputs(5006));
    layer2_outputs(2107) <= layer1_outputs(4162);
    layer2_outputs(2108) <= not(layer1_outputs(3631)) or (layer1_outputs(929));
    layer2_outputs(2109) <= layer1_outputs(4418);
    layer2_outputs(2110) <= (layer1_outputs(2321)) xor (layer1_outputs(364));
    layer2_outputs(2111) <= (layer1_outputs(32)) and not (layer1_outputs(3479));
    layer2_outputs(2112) <= '0';
    layer2_outputs(2113) <= not(layer1_outputs(4008));
    layer2_outputs(2114) <= not(layer1_outputs(1415)) or (layer1_outputs(1945));
    layer2_outputs(2115) <= (layer1_outputs(3481)) or (layer1_outputs(1029));
    layer2_outputs(2116) <= layer1_outputs(962);
    layer2_outputs(2117) <= layer1_outputs(3926);
    layer2_outputs(2118) <= layer1_outputs(1123);
    layer2_outputs(2119) <= (layer1_outputs(2765)) and (layer1_outputs(1947));
    layer2_outputs(2120) <= (layer1_outputs(3884)) and not (layer1_outputs(5010));
    layer2_outputs(2121) <= not(layer1_outputs(4625));
    layer2_outputs(2122) <= layer1_outputs(1098);
    layer2_outputs(2123) <= not((layer1_outputs(3039)) or (layer1_outputs(4311)));
    layer2_outputs(2124) <= not(layer1_outputs(1131));
    layer2_outputs(2125) <= not(layer1_outputs(637));
    layer2_outputs(2126) <= (layer1_outputs(664)) xor (layer1_outputs(3656));
    layer2_outputs(2127) <= layer1_outputs(1314);
    layer2_outputs(2128) <= layer1_outputs(296);
    layer2_outputs(2129) <= not(layer1_outputs(2587));
    layer2_outputs(2130) <= layer1_outputs(4709);
    layer2_outputs(2131) <= not(layer1_outputs(2838));
    layer2_outputs(2132) <= (layer1_outputs(4119)) and (layer1_outputs(4030));
    layer2_outputs(2133) <= not(layer1_outputs(11)) or (layer1_outputs(4821));
    layer2_outputs(2134) <= not(layer1_outputs(433));
    layer2_outputs(2135) <= '0';
    layer2_outputs(2136) <= (layer1_outputs(2601)) and not (layer1_outputs(3341));
    layer2_outputs(2137) <= layer1_outputs(3369);
    layer2_outputs(2138) <= not(layer1_outputs(4820));
    layer2_outputs(2139) <= layer1_outputs(2949);
    layer2_outputs(2140) <= not((layer1_outputs(1027)) or (layer1_outputs(4829)));
    layer2_outputs(2141) <= (layer1_outputs(1262)) and (layer1_outputs(1322));
    layer2_outputs(2142) <= layer1_outputs(1109);
    layer2_outputs(2143) <= (layer1_outputs(1927)) and not (layer1_outputs(90));
    layer2_outputs(2144) <= not(layer1_outputs(2217)) or (layer1_outputs(214));
    layer2_outputs(2145) <= layer1_outputs(1094);
    layer2_outputs(2146) <= layer1_outputs(2138);
    layer2_outputs(2147) <= (layer1_outputs(703)) and not (layer1_outputs(1510));
    layer2_outputs(2148) <= not((layer1_outputs(1225)) xor (layer1_outputs(2016)));
    layer2_outputs(2149) <= not((layer1_outputs(1361)) or (layer1_outputs(4756)));
    layer2_outputs(2150) <= (layer1_outputs(4742)) and (layer1_outputs(4458));
    layer2_outputs(2151) <= layer1_outputs(2678);
    layer2_outputs(2152) <= not(layer1_outputs(1282)) or (layer1_outputs(1465));
    layer2_outputs(2153) <= layer1_outputs(328);
    layer2_outputs(2154) <= layer1_outputs(4280);
    layer2_outputs(2155) <= (layer1_outputs(3760)) and (layer1_outputs(2532));
    layer2_outputs(2156) <= (layer1_outputs(616)) and (layer1_outputs(2513));
    layer2_outputs(2157) <= layer1_outputs(3273);
    layer2_outputs(2158) <= layer1_outputs(942);
    layer2_outputs(2159) <= not(layer1_outputs(3361));
    layer2_outputs(2160) <= (layer1_outputs(308)) or (layer1_outputs(1376));
    layer2_outputs(2161) <= (layer1_outputs(3845)) and not (layer1_outputs(5018));
    layer2_outputs(2162) <= not(layer1_outputs(2548));
    layer2_outputs(2163) <= layer1_outputs(1156);
    layer2_outputs(2164) <= '1';
    layer2_outputs(2165) <= not((layer1_outputs(3346)) and (layer1_outputs(3282)));
    layer2_outputs(2166) <= not(layer1_outputs(2497));
    layer2_outputs(2167) <= layer1_outputs(579);
    layer2_outputs(2168) <= (layer1_outputs(1949)) xor (layer1_outputs(3600));
    layer2_outputs(2169) <= layer1_outputs(860);
    layer2_outputs(2170) <= not(layer1_outputs(1815)) or (layer1_outputs(4236));
    layer2_outputs(2171) <= '1';
    layer2_outputs(2172) <= (layer1_outputs(1389)) or (layer1_outputs(1118));
    layer2_outputs(2173) <= layer1_outputs(2379);
    layer2_outputs(2174) <= not((layer1_outputs(4301)) xor (layer1_outputs(3218)));
    layer2_outputs(2175) <= (layer1_outputs(2599)) or (layer1_outputs(4371));
    layer2_outputs(2176) <= not(layer1_outputs(3735)) or (layer1_outputs(3535));
    layer2_outputs(2177) <= (layer1_outputs(2088)) or (layer1_outputs(3332));
    layer2_outputs(2178) <= not(layer1_outputs(4961)) or (layer1_outputs(1783));
    layer2_outputs(2179) <= (layer1_outputs(4913)) and not (layer1_outputs(1463));
    layer2_outputs(2180) <= '0';
    layer2_outputs(2181) <= layer1_outputs(4488);
    layer2_outputs(2182) <= layer1_outputs(302);
    layer2_outputs(2183) <= (layer1_outputs(1407)) xor (layer1_outputs(756));
    layer2_outputs(2184) <= not(layer1_outputs(4486)) or (layer1_outputs(3102));
    layer2_outputs(2185) <= not(layer1_outputs(1378));
    layer2_outputs(2186) <= (layer1_outputs(5022)) and not (layer1_outputs(3106));
    layer2_outputs(2187) <= not((layer1_outputs(1156)) xor (layer1_outputs(1910)));
    layer2_outputs(2188) <= layer1_outputs(103);
    layer2_outputs(2189) <= (layer1_outputs(3225)) and not (layer1_outputs(3007));
    layer2_outputs(2190) <= not(layer1_outputs(3150));
    layer2_outputs(2191) <= not((layer1_outputs(3081)) xor (layer1_outputs(4805)));
    layer2_outputs(2192) <= (layer1_outputs(4305)) or (layer1_outputs(1424));
    layer2_outputs(2193) <= not(layer1_outputs(3955));
    layer2_outputs(2194) <= not((layer1_outputs(3643)) or (layer1_outputs(3269)));
    layer2_outputs(2195) <= not((layer1_outputs(3403)) and (layer1_outputs(4737)));
    layer2_outputs(2196) <= layer1_outputs(2812);
    layer2_outputs(2197) <= layer1_outputs(1461);
    layer2_outputs(2198) <= not(layer1_outputs(3948));
    layer2_outputs(2199) <= not(layer1_outputs(3842));
    layer2_outputs(2200) <= layer1_outputs(1221);
    layer2_outputs(2201) <= not(layer1_outputs(4972));
    layer2_outputs(2202) <= not((layer1_outputs(3377)) and (layer1_outputs(123)));
    layer2_outputs(2203) <= layer1_outputs(4049);
    layer2_outputs(2204) <= not((layer1_outputs(4332)) or (layer1_outputs(9)));
    layer2_outputs(2205) <= layer1_outputs(2183);
    layer2_outputs(2206) <= layer1_outputs(646);
    layer2_outputs(2207) <= layer1_outputs(1304);
    layer2_outputs(2208) <= not(layer1_outputs(3237));
    layer2_outputs(2209) <= (layer1_outputs(1716)) and not (layer1_outputs(450));
    layer2_outputs(2210) <= not(layer1_outputs(4387));
    layer2_outputs(2211) <= not(layer1_outputs(2620)) or (layer1_outputs(1524));
    layer2_outputs(2212) <= not(layer1_outputs(2654)) or (layer1_outputs(3509));
    layer2_outputs(2213) <= layer1_outputs(2220);
    layer2_outputs(2214) <= layer1_outputs(3736);
    layer2_outputs(2215) <= not(layer1_outputs(3614));
    layer2_outputs(2216) <= layer1_outputs(2438);
    layer2_outputs(2217) <= layer1_outputs(1711);
    layer2_outputs(2218) <= not((layer1_outputs(1572)) xor (layer1_outputs(3567)));
    layer2_outputs(2219) <= not(layer1_outputs(4922));
    layer2_outputs(2220) <= not(layer1_outputs(3766));
    layer2_outputs(2221) <= layer1_outputs(3544);
    layer2_outputs(2222) <= not(layer1_outputs(5031)) or (layer1_outputs(4553));
    layer2_outputs(2223) <= not(layer1_outputs(4627));
    layer2_outputs(2224) <= not(layer1_outputs(3952));
    layer2_outputs(2225) <= (layer1_outputs(4625)) and not (layer1_outputs(660));
    layer2_outputs(2226) <= not(layer1_outputs(2483));
    layer2_outputs(2227) <= not((layer1_outputs(1496)) and (layer1_outputs(2512)));
    layer2_outputs(2228) <= not(layer1_outputs(1508));
    layer2_outputs(2229) <= layer1_outputs(4300);
    layer2_outputs(2230) <= not(layer1_outputs(4167)) or (layer1_outputs(4918));
    layer2_outputs(2231) <= not(layer1_outputs(1184)) or (layer1_outputs(2702));
    layer2_outputs(2232) <= (layer1_outputs(4351)) xor (layer1_outputs(428));
    layer2_outputs(2233) <= layer1_outputs(955);
    layer2_outputs(2234) <= (layer1_outputs(4898)) and (layer1_outputs(4430));
    layer2_outputs(2235) <= not(layer1_outputs(2664));
    layer2_outputs(2236) <= (layer1_outputs(2239)) xor (layer1_outputs(2246));
    layer2_outputs(2237) <= not(layer1_outputs(4655));
    layer2_outputs(2238) <= not(layer1_outputs(3630)) or (layer1_outputs(3808));
    layer2_outputs(2239) <= layer1_outputs(3358);
    layer2_outputs(2240) <= layer1_outputs(511);
    layer2_outputs(2241) <= not(layer1_outputs(1301));
    layer2_outputs(2242) <= layer1_outputs(3040);
    layer2_outputs(2243) <= not(layer1_outputs(1368)) or (layer1_outputs(401));
    layer2_outputs(2244) <= not(layer1_outputs(1657));
    layer2_outputs(2245) <= not(layer1_outputs(4276));
    layer2_outputs(2246) <= (layer1_outputs(2062)) and not (layer1_outputs(2464));
    layer2_outputs(2247) <= layer1_outputs(4369);
    layer2_outputs(2248) <= (layer1_outputs(246)) xor (layer1_outputs(1963));
    layer2_outputs(2249) <= (layer1_outputs(2978)) and (layer1_outputs(4546));
    layer2_outputs(2250) <= (layer1_outputs(1988)) and not (layer1_outputs(2985));
    layer2_outputs(2251) <= (layer1_outputs(522)) or (layer1_outputs(4635));
    layer2_outputs(2252) <= layer1_outputs(470);
    layer2_outputs(2253) <= not((layer1_outputs(3267)) xor (layer1_outputs(1076)));
    layer2_outputs(2254) <= (layer1_outputs(4175)) and (layer1_outputs(4644));
    layer2_outputs(2255) <= not(layer1_outputs(2102));
    layer2_outputs(2256) <= layer1_outputs(1095);
    layer2_outputs(2257) <= not(layer1_outputs(3674));
    layer2_outputs(2258) <= layer1_outputs(1013);
    layer2_outputs(2259) <= (layer1_outputs(278)) or (layer1_outputs(3917));
    layer2_outputs(2260) <= (layer1_outputs(4052)) or (layer1_outputs(48));
    layer2_outputs(2261) <= not(layer1_outputs(3757));
    layer2_outputs(2262) <= not(layer1_outputs(1689)) or (layer1_outputs(2779));
    layer2_outputs(2263) <= layer1_outputs(2754);
    layer2_outputs(2264) <= not((layer1_outputs(1247)) or (layer1_outputs(2356)));
    layer2_outputs(2265) <= not((layer1_outputs(2256)) or (layer1_outputs(4266)));
    layer2_outputs(2266) <= (layer1_outputs(4220)) and not (layer1_outputs(2174));
    layer2_outputs(2267) <= not((layer1_outputs(928)) and (layer1_outputs(78)));
    layer2_outputs(2268) <= (layer1_outputs(3713)) and (layer1_outputs(1855));
    layer2_outputs(2269) <= not(layer1_outputs(1677));
    layer2_outputs(2270) <= layer1_outputs(139);
    layer2_outputs(2271) <= not((layer1_outputs(1752)) or (layer1_outputs(1793)));
    layer2_outputs(2272) <= not(layer1_outputs(970)) or (layer1_outputs(2257));
    layer2_outputs(2273) <= not(layer1_outputs(2430));
    layer2_outputs(2274) <= (layer1_outputs(3895)) and not (layer1_outputs(3275));
    layer2_outputs(2275) <= layer1_outputs(3652);
    layer2_outputs(2276) <= not(layer1_outputs(2232)) or (layer1_outputs(1867));
    layer2_outputs(2277) <= not(layer1_outputs(3558));
    layer2_outputs(2278) <= layer1_outputs(3927);
    layer2_outputs(2279) <= layer1_outputs(4214);
    layer2_outputs(2280) <= not(layer1_outputs(2268)) or (layer1_outputs(3213));
    layer2_outputs(2281) <= layer1_outputs(1071);
    layer2_outputs(2282) <= '1';
    layer2_outputs(2283) <= (layer1_outputs(1954)) or (layer1_outputs(1481));
    layer2_outputs(2284) <= layer1_outputs(4385);
    layer2_outputs(2285) <= layer1_outputs(3890);
    layer2_outputs(2286) <= (layer1_outputs(1822)) or (layer1_outputs(3425));
    layer2_outputs(2287) <= not((layer1_outputs(2067)) or (layer1_outputs(472)));
    layer2_outputs(2288) <= not(layer1_outputs(3433));
    layer2_outputs(2289) <= not(layer1_outputs(645));
    layer2_outputs(2290) <= not(layer1_outputs(1433)) or (layer1_outputs(2071));
    layer2_outputs(2291) <= (layer1_outputs(2983)) and not (layer1_outputs(792));
    layer2_outputs(2292) <= layer1_outputs(3045);
    layer2_outputs(2293) <= layer1_outputs(3934);
    layer2_outputs(2294) <= layer1_outputs(194);
    layer2_outputs(2295) <= not(layer1_outputs(2506)) or (layer1_outputs(1785));
    layer2_outputs(2296) <= layer1_outputs(3261);
    layer2_outputs(2297) <= not(layer1_outputs(2358));
    layer2_outputs(2298) <= layer1_outputs(4291);
    layer2_outputs(2299) <= (layer1_outputs(3085)) and not (layer1_outputs(4855));
    layer2_outputs(2300) <= not((layer1_outputs(2178)) and (layer1_outputs(3291)));
    layer2_outputs(2301) <= (layer1_outputs(3673)) and not (layer1_outputs(1222));
    layer2_outputs(2302) <= not((layer1_outputs(2611)) xor (layer1_outputs(678)));
    layer2_outputs(2303) <= layer1_outputs(4661);
    layer2_outputs(2304) <= layer1_outputs(239);
    layer2_outputs(2305) <= layer1_outputs(4544);
    layer2_outputs(2306) <= not((layer1_outputs(4218)) or (layer1_outputs(3236)));
    layer2_outputs(2307) <= not(layer1_outputs(4412));
    layer2_outputs(2308) <= layer1_outputs(2268);
    layer2_outputs(2309) <= not(layer1_outputs(2388));
    layer2_outputs(2310) <= (layer1_outputs(1413)) and not (layer1_outputs(4355));
    layer2_outputs(2311) <= (layer1_outputs(4495)) or (layer1_outputs(4173));
    layer2_outputs(2312) <= layer1_outputs(4725);
    layer2_outputs(2313) <= (layer1_outputs(5031)) and not (layer1_outputs(2938));
    layer2_outputs(2314) <= not(layer1_outputs(484)) or (layer1_outputs(3868));
    layer2_outputs(2315) <= (layer1_outputs(2632)) or (layer1_outputs(2259));
    layer2_outputs(2316) <= not(layer1_outputs(1092));
    layer2_outputs(2317) <= layer1_outputs(4832);
    layer2_outputs(2318) <= not(layer1_outputs(4627));
    layer2_outputs(2319) <= (layer1_outputs(3026)) and not (layer1_outputs(2373));
    layer2_outputs(2320) <= '1';
    layer2_outputs(2321) <= not(layer1_outputs(2912));
    layer2_outputs(2322) <= (layer1_outputs(1142)) and (layer1_outputs(981));
    layer2_outputs(2323) <= not(layer1_outputs(2029));
    layer2_outputs(2324) <= (layer1_outputs(3582)) or (layer1_outputs(3555));
    layer2_outputs(2325) <= not(layer1_outputs(3848));
    layer2_outputs(2326) <= layer1_outputs(3363);
    layer2_outputs(2327) <= not((layer1_outputs(29)) and (layer1_outputs(4788)));
    layer2_outputs(2328) <= not(layer1_outputs(1820));
    layer2_outputs(2329) <= not(layer1_outputs(5078)) or (layer1_outputs(5027));
    layer2_outputs(2330) <= layer1_outputs(472);
    layer2_outputs(2331) <= not((layer1_outputs(327)) xor (layer1_outputs(2192)));
    layer2_outputs(2332) <= (layer1_outputs(935)) and not (layer1_outputs(407));
    layer2_outputs(2333) <= not((layer1_outputs(3433)) or (layer1_outputs(4155)));
    layer2_outputs(2334) <= (layer1_outputs(4893)) and (layer1_outputs(1073));
    layer2_outputs(2335) <= not(layer1_outputs(16)) or (layer1_outputs(192));
    layer2_outputs(2336) <= (layer1_outputs(5009)) and not (layer1_outputs(296));
    layer2_outputs(2337) <= (layer1_outputs(4975)) or (layer1_outputs(3919));
    layer2_outputs(2338) <= (layer1_outputs(1817)) xor (layer1_outputs(1406));
    layer2_outputs(2339) <= not((layer1_outputs(1592)) and (layer1_outputs(3166)));
    layer2_outputs(2340) <= not(layer1_outputs(4026));
    layer2_outputs(2341) <= not((layer1_outputs(2193)) xor (layer1_outputs(1669)));
    layer2_outputs(2342) <= layer1_outputs(2730);
    layer2_outputs(2343) <= not((layer1_outputs(4106)) and (layer1_outputs(5073)));
    layer2_outputs(2344) <= not(layer1_outputs(2117));
    layer2_outputs(2345) <= not(layer1_outputs(1681));
    layer2_outputs(2346) <= layer1_outputs(4581);
    layer2_outputs(2347) <= not(layer1_outputs(3133));
    layer2_outputs(2348) <= not(layer1_outputs(2996));
    layer2_outputs(2349) <= (layer1_outputs(3599)) and (layer1_outputs(4461));
    layer2_outputs(2350) <= not((layer1_outputs(3903)) or (layer1_outputs(1612)));
    layer2_outputs(2351) <= (layer1_outputs(4417)) and (layer1_outputs(3459));
    layer2_outputs(2352) <= layer1_outputs(1682);
    layer2_outputs(2353) <= not(layer1_outputs(3736)) or (layer1_outputs(2844));
    layer2_outputs(2354) <= layer1_outputs(1569);
    layer2_outputs(2355) <= not(layer1_outputs(3855));
    layer2_outputs(2356) <= not(layer1_outputs(3925));
    layer2_outputs(2357) <= layer1_outputs(3776);
    layer2_outputs(2358) <= (layer1_outputs(1361)) or (layer1_outputs(1849));
    layer2_outputs(2359) <= (layer1_outputs(3345)) xor (layer1_outputs(5063));
    layer2_outputs(2360) <= not((layer1_outputs(4200)) xor (layer1_outputs(2822)));
    layer2_outputs(2361) <= (layer1_outputs(3055)) and (layer1_outputs(4609));
    layer2_outputs(2362) <= not((layer1_outputs(1343)) xor (layer1_outputs(32)));
    layer2_outputs(2363) <= layer1_outputs(1672);
    layer2_outputs(2364) <= not(layer1_outputs(4945)) or (layer1_outputs(2260));
    layer2_outputs(2365) <= (layer1_outputs(3625)) and not (layer1_outputs(2038));
    layer2_outputs(2366) <= not(layer1_outputs(2913));
    layer2_outputs(2367) <= (layer1_outputs(672)) and not (layer1_outputs(358));
    layer2_outputs(2368) <= not(layer1_outputs(735));
    layer2_outputs(2369) <= not(layer1_outputs(2863));
    layer2_outputs(2370) <= (layer1_outputs(2066)) xor (layer1_outputs(5038));
    layer2_outputs(2371) <= layer1_outputs(2271);
    layer2_outputs(2372) <= not((layer1_outputs(1839)) or (layer1_outputs(2462)));
    layer2_outputs(2373) <= not((layer1_outputs(2711)) and (layer1_outputs(3115)));
    layer2_outputs(2374) <= (layer1_outputs(1499)) or (layer1_outputs(317));
    layer2_outputs(2375) <= layer1_outputs(4574);
    layer2_outputs(2376) <= not(layer1_outputs(2367));
    layer2_outputs(2377) <= (layer1_outputs(3299)) or (layer1_outputs(4136));
    layer2_outputs(2378) <= not(layer1_outputs(1933));
    layer2_outputs(2379) <= not(layer1_outputs(4468));
    layer2_outputs(2380) <= not(layer1_outputs(3283));
    layer2_outputs(2381) <= layer1_outputs(1085);
    layer2_outputs(2382) <= not(layer1_outputs(1893));
    layer2_outputs(2383) <= (layer1_outputs(3210)) and (layer1_outputs(4386));
    layer2_outputs(2384) <= (layer1_outputs(2254)) and not (layer1_outputs(4212));
    layer2_outputs(2385) <= not(layer1_outputs(1023)) or (layer1_outputs(4169));
    layer2_outputs(2386) <= not(layer1_outputs(4666));
    layer2_outputs(2387) <= (layer1_outputs(1330)) and (layer1_outputs(4288));
    layer2_outputs(2388) <= layer1_outputs(712);
    layer2_outputs(2389) <= (layer1_outputs(4410)) and not (layer1_outputs(3746));
    layer2_outputs(2390) <= layer1_outputs(3600);
    layer2_outputs(2391) <= not((layer1_outputs(2805)) xor (layer1_outputs(868)));
    layer2_outputs(2392) <= not(layer1_outputs(4191));
    layer2_outputs(2393) <= not((layer1_outputs(1585)) xor (layer1_outputs(883)));
    layer2_outputs(2394) <= layer1_outputs(3110);
    layer2_outputs(2395) <= (layer1_outputs(1930)) and not (layer1_outputs(1260));
    layer2_outputs(2396) <= layer1_outputs(468);
    layer2_outputs(2397) <= not((layer1_outputs(2500)) xor (layer1_outputs(1529)));
    layer2_outputs(2398) <= not((layer1_outputs(1240)) xor (layer1_outputs(1876)));
    layer2_outputs(2399) <= not(layer1_outputs(1525));
    layer2_outputs(2400) <= not(layer1_outputs(4561)) or (layer1_outputs(2288));
    layer2_outputs(2401) <= (layer1_outputs(4290)) and (layer1_outputs(1995));
    layer2_outputs(2402) <= not(layer1_outputs(668));
    layer2_outputs(2403) <= (layer1_outputs(4870)) xor (layer1_outputs(4857));
    layer2_outputs(2404) <= not(layer1_outputs(161));
    layer2_outputs(2405) <= layer1_outputs(3558);
    layer2_outputs(2406) <= not(layer1_outputs(4143));
    layer2_outputs(2407) <= not(layer1_outputs(1346)) or (layer1_outputs(483));
    layer2_outputs(2408) <= not(layer1_outputs(3365));
    layer2_outputs(2409) <= not(layer1_outputs(1016)) or (layer1_outputs(4046));
    layer2_outputs(2410) <= not(layer1_outputs(187)) or (layer1_outputs(4906));
    layer2_outputs(2411) <= (layer1_outputs(2441)) and not (layer1_outputs(4453));
    layer2_outputs(2412) <= layer1_outputs(2090);
    layer2_outputs(2413) <= not(layer1_outputs(40));
    layer2_outputs(2414) <= layer1_outputs(4151);
    layer2_outputs(2415) <= layer1_outputs(3190);
    layer2_outputs(2416) <= not(layer1_outputs(3059));
    layer2_outputs(2417) <= not(layer1_outputs(341));
    layer2_outputs(2418) <= layer1_outputs(3431);
    layer2_outputs(2419) <= '0';
    layer2_outputs(2420) <= layer1_outputs(3752);
    layer2_outputs(2421) <= not(layer1_outputs(1758)) or (layer1_outputs(3755));
    layer2_outputs(2422) <= not(layer1_outputs(277)) or (layer1_outputs(1644));
    layer2_outputs(2423) <= not(layer1_outputs(2829));
    layer2_outputs(2424) <= (layer1_outputs(4484)) and (layer1_outputs(951));
    layer2_outputs(2425) <= layer1_outputs(2768);
    layer2_outputs(2426) <= not(layer1_outputs(3648)) or (layer1_outputs(3391));
    layer2_outputs(2427) <= not(layer1_outputs(5017));
    layer2_outputs(2428) <= (layer1_outputs(2539)) and not (layer1_outputs(4765));
    layer2_outputs(2429) <= not(layer1_outputs(3230));
    layer2_outputs(2430) <= layer1_outputs(2133);
    layer2_outputs(2431) <= not(layer1_outputs(4119));
    layer2_outputs(2432) <= not(layer1_outputs(2035)) or (layer1_outputs(1957));
    layer2_outputs(2433) <= not(layer1_outputs(459));
    layer2_outputs(2434) <= not((layer1_outputs(2970)) and (layer1_outputs(3061)));
    layer2_outputs(2435) <= not(layer1_outputs(318));
    layer2_outputs(2436) <= not((layer1_outputs(445)) or (layer1_outputs(2225)));
    layer2_outputs(2437) <= not(layer1_outputs(709));
    layer2_outputs(2438) <= not(layer1_outputs(3609));
    layer2_outputs(2439) <= layer1_outputs(368);
    layer2_outputs(2440) <= layer1_outputs(3548);
    layer2_outputs(2441) <= (layer1_outputs(1363)) and not (layer1_outputs(4598));
    layer2_outputs(2442) <= not(layer1_outputs(3743)) or (layer1_outputs(4244));
    layer2_outputs(2443) <= not((layer1_outputs(627)) and (layer1_outputs(4713)));
    layer2_outputs(2444) <= not(layer1_outputs(4333)) or (layer1_outputs(205));
    layer2_outputs(2445) <= (layer1_outputs(2871)) xor (layer1_outputs(4176));
    layer2_outputs(2446) <= not(layer1_outputs(3832));
    layer2_outputs(2447) <= layer1_outputs(1902);
    layer2_outputs(2448) <= not(layer1_outputs(2236));
    layer2_outputs(2449) <= not((layer1_outputs(1444)) xor (layer1_outputs(2923)));
    layer2_outputs(2450) <= not((layer1_outputs(2442)) and (layer1_outputs(1882)));
    layer2_outputs(2451) <= not(layer1_outputs(2177));
    layer2_outputs(2452) <= not(layer1_outputs(412));
    layer2_outputs(2453) <= (layer1_outputs(998)) and (layer1_outputs(3340));
    layer2_outputs(2454) <= (layer1_outputs(2850)) and not (layer1_outputs(956));
    layer2_outputs(2455) <= layer1_outputs(1545);
    layer2_outputs(2456) <= not(layer1_outputs(560));
    layer2_outputs(2457) <= layer1_outputs(394);
    layer2_outputs(2458) <= layer1_outputs(4483);
    layer2_outputs(2459) <= not((layer1_outputs(3371)) and (layer1_outputs(1565)));
    layer2_outputs(2460) <= (layer1_outputs(4804)) or (layer1_outputs(3772));
    layer2_outputs(2461) <= layer1_outputs(2549);
    layer2_outputs(2462) <= (layer1_outputs(1252)) and (layer1_outputs(1831));
    layer2_outputs(2463) <= (layer1_outputs(2973)) or (layer1_outputs(1177));
    layer2_outputs(2464) <= not((layer1_outputs(1915)) and (layer1_outputs(387)));
    layer2_outputs(2465) <= layer1_outputs(204);
    layer2_outputs(2466) <= not((layer1_outputs(3506)) and (layer1_outputs(2015)));
    layer2_outputs(2467) <= not(layer1_outputs(2785));
    layer2_outputs(2468) <= not(layer1_outputs(430));
    layer2_outputs(2469) <= layer1_outputs(2726);
    layer2_outputs(2470) <= layer1_outputs(95);
    layer2_outputs(2471) <= '1';
    layer2_outputs(2472) <= not(layer1_outputs(4582));
    layer2_outputs(2473) <= not((layer1_outputs(825)) xor (layer1_outputs(466)));
    layer2_outputs(2474) <= layer1_outputs(3475);
    layer2_outputs(2475) <= not((layer1_outputs(926)) and (layer1_outputs(2511)));
    layer2_outputs(2476) <= (layer1_outputs(4045)) and not (layer1_outputs(235));
    layer2_outputs(2477) <= layer1_outputs(1121);
    layer2_outputs(2478) <= not((layer1_outputs(902)) xor (layer1_outputs(4092)));
    layer2_outputs(2479) <= layer1_outputs(2719);
    layer2_outputs(2480) <= (layer1_outputs(91)) and (layer1_outputs(4664));
    layer2_outputs(2481) <= (layer1_outputs(2671)) xor (layer1_outputs(3372));
    layer2_outputs(2482) <= not(layer1_outputs(476));
    layer2_outputs(2483) <= not(layer1_outputs(2557)) or (layer1_outputs(931));
    layer2_outputs(2484) <= (layer1_outputs(878)) or (layer1_outputs(1122));
    layer2_outputs(2485) <= not(layer1_outputs(2690));
    layer2_outputs(2486) <= (layer1_outputs(3322)) or (layer1_outputs(3447));
    layer2_outputs(2487) <= not((layer1_outputs(5086)) and (layer1_outputs(396)));
    layer2_outputs(2488) <= not((layer1_outputs(2732)) xor (layer1_outputs(2517)));
    layer2_outputs(2489) <= not((layer1_outputs(1551)) and (layer1_outputs(2501)));
    layer2_outputs(2490) <= (layer1_outputs(1266)) and (layer1_outputs(327));
    layer2_outputs(2491) <= (layer1_outputs(4489)) and not (layer1_outputs(2143));
    layer2_outputs(2492) <= not(layer1_outputs(1494));
    layer2_outputs(2493) <= not((layer1_outputs(1126)) or (layer1_outputs(922)));
    layer2_outputs(2494) <= layer1_outputs(79);
    layer2_outputs(2495) <= not((layer1_outputs(3576)) and (layer1_outputs(3750)));
    layer2_outputs(2496) <= not(layer1_outputs(2602));
    layer2_outputs(2497) <= layer1_outputs(3709);
    layer2_outputs(2498) <= not(layer1_outputs(990));
    layer2_outputs(2499) <= not(layer1_outputs(425));
    layer2_outputs(2500) <= not((layer1_outputs(2264)) or (layer1_outputs(2284)));
    layer2_outputs(2501) <= not((layer1_outputs(3894)) and (layer1_outputs(4868)));
    layer2_outputs(2502) <= not(layer1_outputs(4356));
    layer2_outputs(2503) <= (layer1_outputs(5053)) and (layer1_outputs(4183));
    layer2_outputs(2504) <= (layer1_outputs(4070)) xor (layer1_outputs(1566));
    layer2_outputs(2505) <= layer1_outputs(4826);
    layer2_outputs(2506) <= (layer1_outputs(3491)) and not (layer1_outputs(3284));
    layer2_outputs(2507) <= not(layer1_outputs(1613));
    layer2_outputs(2508) <= not(layer1_outputs(5068));
    layer2_outputs(2509) <= not(layer1_outputs(2298)) or (layer1_outputs(4059));
    layer2_outputs(2510) <= not(layer1_outputs(3189)) or (layer1_outputs(2921));
    layer2_outputs(2511) <= (layer1_outputs(4942)) and not (layer1_outputs(1682));
    layer2_outputs(2512) <= layer1_outputs(1360);
    layer2_outputs(2513) <= (layer1_outputs(4362)) or (layer1_outputs(2399));
    layer2_outputs(2514) <= layer1_outputs(1170);
    layer2_outputs(2515) <= not(layer1_outputs(4489));
    layer2_outputs(2516) <= layer1_outputs(2098);
    layer2_outputs(2517) <= layer1_outputs(1440);
    layer2_outputs(2518) <= (layer1_outputs(2742)) and not (layer1_outputs(601));
    layer2_outputs(2519) <= (layer1_outputs(3503)) and not (layer1_outputs(203));
    layer2_outputs(2520) <= not((layer1_outputs(4330)) and (layer1_outputs(3234)));
    layer2_outputs(2521) <= not(layer1_outputs(4850)) or (layer1_outputs(4085));
    layer2_outputs(2522) <= (layer1_outputs(4504)) or (layer1_outputs(4832));
    layer2_outputs(2523) <= not(layer1_outputs(2928));
    layer2_outputs(2524) <= not(layer1_outputs(4855));
    layer2_outputs(2525) <= not(layer1_outputs(3921));
    layer2_outputs(2526) <= (layer1_outputs(3992)) or (layer1_outputs(4303));
    layer2_outputs(2527) <= not((layer1_outputs(2151)) and (layer1_outputs(4023)));
    layer2_outputs(2528) <= not(layer1_outputs(1962));
    layer2_outputs(2529) <= (layer1_outputs(1893)) and not (layer1_outputs(1226));
    layer2_outputs(2530) <= not((layer1_outputs(4821)) xor (layer1_outputs(1931)));
    layer2_outputs(2531) <= (layer1_outputs(4571)) xor (layer1_outputs(959));
    layer2_outputs(2532) <= not(layer1_outputs(2927));
    layer2_outputs(2533) <= not(layer1_outputs(4580));
    layer2_outputs(2534) <= layer1_outputs(1134);
    layer2_outputs(2535) <= layer1_outputs(1123);
    layer2_outputs(2536) <= not(layer1_outputs(613));
    layer2_outputs(2537) <= not(layer1_outputs(2551));
    layer2_outputs(2538) <= layer1_outputs(3956);
    layer2_outputs(2539) <= not((layer1_outputs(2030)) xor (layer1_outputs(4815)));
    layer2_outputs(2540) <= layer1_outputs(4022);
    layer2_outputs(2541) <= not(layer1_outputs(4038));
    layer2_outputs(2542) <= (layer1_outputs(4890)) or (layer1_outputs(4241));
    layer2_outputs(2543) <= layer1_outputs(969);
    layer2_outputs(2544) <= layer1_outputs(794);
    layer2_outputs(2545) <= not((layer1_outputs(2359)) or (layer1_outputs(632)));
    layer2_outputs(2546) <= not((layer1_outputs(1874)) xor (layer1_outputs(4873)));
    layer2_outputs(2547) <= (layer1_outputs(665)) and (layer1_outputs(2224));
    layer2_outputs(2548) <= not((layer1_outputs(2039)) xor (layer1_outputs(5025)));
    layer2_outputs(2549) <= layer1_outputs(1555);
    layer2_outputs(2550) <= not(layer1_outputs(947));
    layer2_outputs(2551) <= not(layer1_outputs(3596)) or (layer1_outputs(1209));
    layer2_outputs(2552) <= (layer1_outputs(4400)) or (layer1_outputs(4294));
    layer2_outputs(2553) <= layer1_outputs(4346);
    layer2_outputs(2554) <= not((layer1_outputs(5055)) xor (layer1_outputs(3462)));
    layer2_outputs(2555) <= not((layer1_outputs(2468)) or (layer1_outputs(2640)));
    layer2_outputs(2556) <= (layer1_outputs(4792)) and not (layer1_outputs(673));
    layer2_outputs(2557) <= not(layer1_outputs(4963));
    layer2_outputs(2558) <= layer1_outputs(1730);
    layer2_outputs(2559) <= not(layer1_outputs(1730)) or (layer1_outputs(5023));
    layer2_outputs(2560) <= layer1_outputs(4151);
    layer2_outputs(2561) <= (layer1_outputs(2127)) or (layer1_outputs(1127));
    layer2_outputs(2562) <= layer1_outputs(4698);
    layer2_outputs(2563) <= (layer1_outputs(1443)) xor (layer1_outputs(2073));
    layer2_outputs(2564) <= not(layer1_outputs(1522));
    layer2_outputs(2565) <= '1';
    layer2_outputs(2566) <= not(layer1_outputs(4550));
    layer2_outputs(2567) <= not(layer1_outputs(4448));
    layer2_outputs(2568) <= not((layer1_outputs(1484)) and (layer1_outputs(3819)));
    layer2_outputs(2569) <= not(layer1_outputs(1390));
    layer2_outputs(2570) <= not((layer1_outputs(5065)) and (layer1_outputs(4940)));
    layer2_outputs(2571) <= layer1_outputs(3822);
    layer2_outputs(2572) <= (layer1_outputs(2457)) and not (layer1_outputs(1773));
    layer2_outputs(2573) <= (layer1_outputs(3970)) and not (layer1_outputs(2233));
    layer2_outputs(2574) <= not((layer1_outputs(4378)) or (layer1_outputs(2666)));
    layer2_outputs(2575) <= (layer1_outputs(3448)) and not (layer1_outputs(890));
    layer2_outputs(2576) <= (layer1_outputs(3267)) and not (layer1_outputs(566));
    layer2_outputs(2577) <= not(layer1_outputs(538)) or (layer1_outputs(3218));
    layer2_outputs(2578) <= not(layer1_outputs(5083));
    layer2_outputs(2579) <= (layer1_outputs(2626)) or (layer1_outputs(3090));
    layer2_outputs(2580) <= (layer1_outputs(2146)) and (layer1_outputs(2144));
    layer2_outputs(2581) <= not(layer1_outputs(4181)) or (layer1_outputs(1713));
    layer2_outputs(2582) <= not(layer1_outputs(3644));
    layer2_outputs(2583) <= (layer1_outputs(2669)) and not (layer1_outputs(2505));
    layer2_outputs(2584) <= not(layer1_outputs(3230));
    layer2_outputs(2585) <= not(layer1_outputs(1645));
    layer2_outputs(2586) <= not(layer1_outputs(4179));
    layer2_outputs(2587) <= not(layer1_outputs(3572));
    layer2_outputs(2588) <= layer1_outputs(1536);
    layer2_outputs(2589) <= layer1_outputs(3879);
    layer2_outputs(2590) <= (layer1_outputs(3147)) or (layer1_outputs(3857));
    layer2_outputs(2591) <= layer1_outputs(4022);
    layer2_outputs(2592) <= not(layer1_outputs(1886));
    layer2_outputs(2593) <= (layer1_outputs(1452)) and not (layer1_outputs(697));
    layer2_outputs(2594) <= layer1_outputs(1035);
    layer2_outputs(2595) <= not((layer1_outputs(5044)) xor (layer1_outputs(4566)));
    layer2_outputs(2596) <= not(layer1_outputs(3455));
    layer2_outputs(2597) <= not(layer1_outputs(4798));
    layer2_outputs(2598) <= layer1_outputs(708);
    layer2_outputs(2599) <= not(layer1_outputs(2366));
    layer2_outputs(2600) <= not(layer1_outputs(901));
    layer2_outputs(2601) <= not((layer1_outputs(2349)) xor (layer1_outputs(3902)));
    layer2_outputs(2602) <= not((layer1_outputs(3052)) xor (layer1_outputs(4352)));
    layer2_outputs(2603) <= not(layer1_outputs(3812));
    layer2_outputs(2604) <= (layer1_outputs(5064)) and not (layer1_outputs(2836));
    layer2_outputs(2605) <= (layer1_outputs(1939)) xor (layer1_outputs(4122));
    layer2_outputs(2606) <= not(layer1_outputs(1695));
    layer2_outputs(2607) <= (layer1_outputs(3978)) and (layer1_outputs(2972));
    layer2_outputs(2608) <= (layer1_outputs(5042)) and not (layer1_outputs(1653));
    layer2_outputs(2609) <= layer1_outputs(2333);
    layer2_outputs(2610) <= not(layer1_outputs(1427));
    layer2_outputs(2611) <= (layer1_outputs(1540)) or (layer1_outputs(1122));
    layer2_outputs(2612) <= layer1_outputs(2488);
    layer2_outputs(2613) <= not((layer1_outputs(1027)) or (layer1_outputs(2106)));
    layer2_outputs(2614) <= not((layer1_outputs(4558)) or (layer1_outputs(4449)));
    layer2_outputs(2615) <= not(layer1_outputs(1680));
    layer2_outputs(2616) <= not(layer1_outputs(3319)) or (layer1_outputs(1279));
    layer2_outputs(2617) <= (layer1_outputs(3489)) and not (layer1_outputs(1053));
    layer2_outputs(2618) <= (layer1_outputs(3729)) and (layer1_outputs(4000));
    layer2_outputs(2619) <= not(layer1_outputs(1727)) or (layer1_outputs(4978));
    layer2_outputs(2620) <= (layer1_outputs(2323)) xor (layer1_outputs(3770));
    layer2_outputs(2621) <= not((layer1_outputs(2809)) xor (layer1_outputs(3551)));
    layer2_outputs(2622) <= layer1_outputs(3116);
    layer2_outputs(2623) <= layer1_outputs(4306);
    layer2_outputs(2624) <= layer1_outputs(292);
    layer2_outputs(2625) <= not(layer1_outputs(418));
    layer2_outputs(2626) <= (layer1_outputs(2915)) xor (layer1_outputs(3941));
    layer2_outputs(2627) <= layer1_outputs(1895);
    layer2_outputs(2628) <= layer1_outputs(4615);
    layer2_outputs(2629) <= not(layer1_outputs(3422));
    layer2_outputs(2630) <= not(layer1_outputs(2261));
    layer2_outputs(2631) <= not(layer1_outputs(1472));
    layer2_outputs(2632) <= layer1_outputs(4654);
    layer2_outputs(2633) <= layer1_outputs(5051);
    layer2_outputs(2634) <= not(layer1_outputs(2172));
    layer2_outputs(2635) <= not((layer1_outputs(1973)) and (layer1_outputs(4436)));
    layer2_outputs(2636) <= layer1_outputs(357);
    layer2_outputs(2637) <= not((layer1_outputs(1501)) or (layer1_outputs(3268)));
    layer2_outputs(2638) <= layer1_outputs(2214);
    layer2_outputs(2639) <= (layer1_outputs(4960)) and (layer1_outputs(1087));
    layer2_outputs(2640) <= layer1_outputs(1648);
    layer2_outputs(2641) <= not(layer1_outputs(2823)) or (layer1_outputs(3118));
    layer2_outputs(2642) <= (layer1_outputs(1445)) xor (layer1_outputs(4518));
    layer2_outputs(2643) <= not(layer1_outputs(1251));
    layer2_outputs(2644) <= not(layer1_outputs(2498));
    layer2_outputs(2645) <= (layer1_outputs(3324)) and not (layer1_outputs(2292));
    layer2_outputs(2646) <= not((layer1_outputs(1357)) or (layer1_outputs(1338)));
    layer2_outputs(2647) <= not(layer1_outputs(2934));
    layer2_outputs(2648) <= layer1_outputs(4462);
    layer2_outputs(2649) <= (layer1_outputs(453)) and not (layer1_outputs(1254));
    layer2_outputs(2650) <= layer1_outputs(4056);
    layer2_outputs(2651) <= not(layer1_outputs(603));
    layer2_outputs(2652) <= (layer1_outputs(1636)) xor (layer1_outputs(3277));
    layer2_outputs(2653) <= layer1_outputs(2781);
    layer2_outputs(2654) <= not(layer1_outputs(2137)) or (layer1_outputs(226));
    layer2_outputs(2655) <= (layer1_outputs(3526)) or (layer1_outputs(2661));
    layer2_outputs(2656) <= layer1_outputs(3555);
    layer2_outputs(2657) <= (layer1_outputs(276)) and (layer1_outputs(4861));
    layer2_outputs(2658) <= not(layer1_outputs(2432)) or (layer1_outputs(3470));
    layer2_outputs(2659) <= (layer1_outputs(2919)) and (layer1_outputs(1248));
    layer2_outputs(2660) <= (layer1_outputs(2641)) xor (layer1_outputs(1125));
    layer2_outputs(2661) <= layer1_outputs(1616);
    layer2_outputs(2662) <= not(layer1_outputs(3850));
    layer2_outputs(2663) <= not(layer1_outputs(2721));
    layer2_outputs(2664) <= not((layer1_outputs(2485)) and (layer1_outputs(738)));
    layer2_outputs(2665) <= not(layer1_outputs(3725));
    layer2_outputs(2666) <= not(layer1_outputs(3472));
    layer2_outputs(2667) <= layer1_outputs(819);
    layer2_outputs(2668) <= not(layer1_outputs(4015));
    layer2_outputs(2669) <= not((layer1_outputs(3646)) or (layer1_outputs(3996)));
    layer2_outputs(2670) <= not((layer1_outputs(1403)) and (layer1_outputs(1001)));
    layer2_outputs(2671) <= (layer1_outputs(241)) and not (layer1_outputs(4722));
    layer2_outputs(2672) <= layer1_outputs(1351);
    layer2_outputs(2673) <= not(layer1_outputs(2745));
    layer2_outputs(2674) <= layer1_outputs(2987);
    layer2_outputs(2675) <= not(layer1_outputs(3305));
    layer2_outputs(2676) <= not(layer1_outputs(2909));
    layer2_outputs(2677) <= not(layer1_outputs(3082)) or (layer1_outputs(1561));
    layer2_outputs(2678) <= layer1_outputs(4341);
    layer2_outputs(2679) <= not((layer1_outputs(2440)) and (layer1_outputs(2974)));
    layer2_outputs(2680) <= not(layer1_outputs(2331)) or (layer1_outputs(1143));
    layer2_outputs(2681) <= layer1_outputs(2734);
    layer2_outputs(2682) <= (layer1_outputs(1587)) or (layer1_outputs(3642));
    layer2_outputs(2683) <= not(layer1_outputs(452));
    layer2_outputs(2684) <= not(layer1_outputs(594));
    layer2_outputs(2685) <= not(layer1_outputs(2391)) or (layer1_outputs(3581));
    layer2_outputs(2686) <= (layer1_outputs(3835)) and not (layer1_outputs(2718));
    layer2_outputs(2687) <= not((layer1_outputs(4771)) xor (layer1_outputs(252)));
    layer2_outputs(2688) <= layer1_outputs(4234);
    layer2_outputs(2689) <= (layer1_outputs(1697)) xor (layer1_outputs(3665));
    layer2_outputs(2690) <= (layer1_outputs(4339)) and not (layer1_outputs(4278));
    layer2_outputs(2691) <= not((layer1_outputs(530)) xor (layer1_outputs(4854)));
    layer2_outputs(2692) <= layer1_outputs(1943);
    layer2_outputs(2693) <= not(layer1_outputs(176));
    layer2_outputs(2694) <= not(layer1_outputs(2377)) or (layer1_outputs(2961));
    layer2_outputs(2695) <= not(layer1_outputs(3830)) or (layer1_outputs(1485));
    layer2_outputs(2696) <= not((layer1_outputs(2253)) and (layer1_outputs(3738)));
    layer2_outputs(2697) <= (layer1_outputs(210)) and not (layer1_outputs(4130));
    layer2_outputs(2698) <= layer1_outputs(4102);
    layer2_outputs(2699) <= not((layer1_outputs(1384)) and (layer1_outputs(2977)));
    layer2_outputs(2700) <= '0';
    layer2_outputs(2701) <= not((layer1_outputs(4240)) and (layer1_outputs(384)));
    layer2_outputs(2702) <= not(layer1_outputs(614));
    layer2_outputs(2703) <= not(layer1_outputs(172));
    layer2_outputs(2704) <= not(layer1_outputs(1666));
    layer2_outputs(2705) <= not((layer1_outputs(1995)) or (layer1_outputs(1000)));
    layer2_outputs(2706) <= not((layer1_outputs(4314)) xor (layer1_outputs(1138)));
    layer2_outputs(2707) <= layer1_outputs(2962);
    layer2_outputs(2708) <= not(layer1_outputs(4917));
    layer2_outputs(2709) <= (layer1_outputs(2121)) and not (layer1_outputs(3496));
    layer2_outputs(2710) <= layer1_outputs(4604);
    layer2_outputs(2711) <= not(layer1_outputs(2113));
    layer2_outputs(2712) <= not(layer1_outputs(2001));
    layer2_outputs(2713) <= not((layer1_outputs(1601)) and (layer1_outputs(2914)));
    layer2_outputs(2714) <= (layer1_outputs(2187)) and not (layer1_outputs(405));
    layer2_outputs(2715) <= layer1_outputs(930);
    layer2_outputs(2716) <= not(layer1_outputs(3408));
    layer2_outputs(2717) <= (layer1_outputs(806)) or (layer1_outputs(2842));
    layer2_outputs(2718) <= not(layer1_outputs(3407));
    layer2_outputs(2719) <= not(layer1_outputs(3320));
    layer2_outputs(2720) <= not((layer1_outputs(1805)) or (layer1_outputs(3805)));
    layer2_outputs(2721) <= not((layer1_outputs(62)) and (layer1_outputs(3605)));
    layer2_outputs(2722) <= not((layer1_outputs(1326)) xor (layer1_outputs(3289)));
    layer2_outputs(2723) <= not(layer1_outputs(5096));
    layer2_outputs(2724) <= not(layer1_outputs(2997)) or (layer1_outputs(447));
    layer2_outputs(2725) <= not(layer1_outputs(2279));
    layer2_outputs(2726) <= not(layer1_outputs(4397));
    layer2_outputs(2727) <= not(layer1_outputs(1507));
    layer2_outputs(2728) <= layer1_outputs(4548);
    layer2_outputs(2729) <= (layer1_outputs(1663)) and not (layer1_outputs(3732));
    layer2_outputs(2730) <= not(layer1_outputs(3043));
    layer2_outputs(2731) <= layer1_outputs(1299);
    layer2_outputs(2732) <= not(layer1_outputs(3823));
    layer2_outputs(2733) <= not(layer1_outputs(293));
    layer2_outputs(2734) <= not(layer1_outputs(4695));
    layer2_outputs(2735) <= not(layer1_outputs(442));
    layer2_outputs(2736) <= not(layer1_outputs(3042));
    layer2_outputs(2737) <= (layer1_outputs(1742)) and not (layer1_outputs(3077));
    layer2_outputs(2738) <= layer1_outputs(3426);
    layer2_outputs(2739) <= (layer1_outputs(2860)) and not (layer1_outputs(3699));
    layer2_outputs(2740) <= layer1_outputs(3164);
    layer2_outputs(2741) <= (layer1_outputs(606)) xor (layer1_outputs(904));
    layer2_outputs(2742) <= (layer1_outputs(2007)) and not (layer1_outputs(117));
    layer2_outputs(2743) <= not(layer1_outputs(857));
    layer2_outputs(2744) <= not(layer1_outputs(2701));
    layer2_outputs(2745) <= not(layer1_outputs(3504));
    layer2_outputs(2746) <= not(layer1_outputs(3135));
    layer2_outputs(2747) <= not(layer1_outputs(966));
    layer2_outputs(2748) <= not(layer1_outputs(4906));
    layer2_outputs(2749) <= (layer1_outputs(4115)) and not (layer1_outputs(4956));
    layer2_outputs(2750) <= layer1_outputs(4700);
    layer2_outputs(2751) <= layer1_outputs(485);
    layer2_outputs(2752) <= layer1_outputs(479);
    layer2_outputs(2753) <= '1';
    layer2_outputs(2754) <= not((layer1_outputs(889)) xor (layer1_outputs(2297)));
    layer2_outputs(2755) <= not(layer1_outputs(4715));
    layer2_outputs(2756) <= not(layer1_outputs(3659)) or (layer1_outputs(4292));
    layer2_outputs(2757) <= layer1_outputs(4178);
    layer2_outputs(2758) <= not(layer1_outputs(1933)) or (layer1_outputs(3704));
    layer2_outputs(2759) <= layer1_outputs(1576);
    layer2_outputs(2760) <= (layer1_outputs(4887)) and (layer1_outputs(3769));
    layer2_outputs(2761) <= not((layer1_outputs(4693)) and (layer1_outputs(1157)));
    layer2_outputs(2762) <= not(layer1_outputs(4927));
    layer2_outputs(2763) <= not((layer1_outputs(4161)) or (layer1_outputs(3955)));
    layer2_outputs(2764) <= (layer1_outputs(3403)) xor (layer1_outputs(2558));
    layer2_outputs(2765) <= not(layer1_outputs(1491));
    layer2_outputs(2766) <= layer1_outputs(1324);
    layer2_outputs(2767) <= layer1_outputs(4376);
    layer2_outputs(2768) <= layer1_outputs(1509);
    layer2_outputs(2769) <= (layer1_outputs(1386)) xor (layer1_outputs(1200));
    layer2_outputs(2770) <= not((layer1_outputs(682)) xor (layer1_outputs(2121)));
    layer2_outputs(2771) <= not((layer1_outputs(4253)) xor (layer1_outputs(337)));
    layer2_outputs(2772) <= not((layer1_outputs(2281)) or (layer1_outputs(1228)));
    layer2_outputs(2773) <= layer1_outputs(4657);
    layer2_outputs(2774) <= (layer1_outputs(3832)) and not (layer1_outputs(1939));
    layer2_outputs(2775) <= not(layer1_outputs(229)) or (layer1_outputs(2105));
    layer2_outputs(2776) <= not((layer1_outputs(298)) or (layer1_outputs(3530)));
    layer2_outputs(2777) <= (layer1_outputs(2447)) and (layer1_outputs(4816));
    layer2_outputs(2778) <= '0';
    layer2_outputs(2779) <= not((layer1_outputs(1554)) or (layer1_outputs(3560)));
    layer2_outputs(2780) <= (layer1_outputs(1558)) and (layer1_outputs(4776));
    layer2_outputs(2781) <= not((layer1_outputs(5039)) and (layer1_outputs(1654)));
    layer2_outputs(2782) <= not(layer1_outputs(1437));
    layer2_outputs(2783) <= (layer1_outputs(3041)) and (layer1_outputs(4147));
    layer2_outputs(2784) <= not(layer1_outputs(2645)) or (layer1_outputs(3649));
    layer2_outputs(2785) <= layer1_outputs(3954);
    layer2_outputs(2786) <= (layer1_outputs(3350)) xor (layer1_outputs(4818));
    layer2_outputs(2787) <= not((layer1_outputs(117)) and (layer1_outputs(4558)));
    layer2_outputs(2788) <= not(layer1_outputs(1276));
    layer2_outputs(2789) <= (layer1_outputs(3627)) and not (layer1_outputs(3657));
    layer2_outputs(2790) <= not(layer1_outputs(1527)) or (layer1_outputs(3525));
    layer2_outputs(2791) <= layer1_outputs(2306);
    layer2_outputs(2792) <= layer1_outputs(161);
    layer2_outputs(2793) <= layer1_outputs(4696);
    layer2_outputs(2794) <= not((layer1_outputs(4902)) or (layer1_outputs(284)));
    layer2_outputs(2795) <= not(layer1_outputs(2653)) or (layer1_outputs(3728));
    layer2_outputs(2796) <= layer1_outputs(5103);
    layer2_outputs(2797) <= not(layer1_outputs(3152));
    layer2_outputs(2798) <= not(layer1_outputs(3789)) or (layer1_outputs(3509));
    layer2_outputs(2799) <= not(layer1_outputs(149));
    layer2_outputs(2800) <= (layer1_outputs(2476)) or (layer1_outputs(3276));
    layer2_outputs(2801) <= (layer1_outputs(3255)) xor (layer1_outputs(3673));
    layer2_outputs(2802) <= (layer1_outputs(5056)) and not (layer1_outputs(3316));
    layer2_outputs(2803) <= not(layer1_outputs(2679));
    layer2_outputs(2804) <= not(layer1_outputs(2941));
    layer2_outputs(2805) <= (layer1_outputs(4602)) and (layer1_outputs(2476));
    layer2_outputs(2806) <= layer1_outputs(3934);
    layer2_outputs(2807) <= not((layer1_outputs(3569)) and (layer1_outputs(4494)));
    layer2_outputs(2808) <= not(layer1_outputs(353)) or (layer1_outputs(820));
    layer2_outputs(2809) <= layer1_outputs(1762);
    layer2_outputs(2810) <= not(layer1_outputs(2398));
    layer2_outputs(2811) <= not((layer1_outputs(1716)) and (layer1_outputs(1843)));
    layer2_outputs(2812) <= not((layer1_outputs(4747)) or (layer1_outputs(2101)));
    layer2_outputs(2813) <= layer1_outputs(175);
    layer2_outputs(2814) <= not(layer1_outputs(651)) or (layer1_outputs(1728));
    layer2_outputs(2815) <= not(layer1_outputs(1367)) or (layer1_outputs(2334));
    layer2_outputs(2816) <= not(layer1_outputs(1798));
    layer2_outputs(2817) <= not(layer1_outputs(3036));
    layer2_outputs(2818) <= not(layer1_outputs(4053)) or (layer1_outputs(2787));
    layer2_outputs(2819) <= (layer1_outputs(3716)) and (layer1_outputs(4987));
    layer2_outputs(2820) <= not((layer1_outputs(3825)) and (layer1_outputs(345)));
    layer2_outputs(2821) <= not(layer1_outputs(306));
    layer2_outputs(2822) <= (layer1_outputs(4384)) and (layer1_outputs(3245));
    layer2_outputs(2823) <= not(layer1_outputs(122));
    layer2_outputs(2824) <= (layer1_outputs(473)) and (layer1_outputs(2165));
    layer2_outputs(2825) <= layer1_outputs(4502);
    layer2_outputs(2826) <= layer1_outputs(387);
    layer2_outputs(2827) <= (layer1_outputs(4703)) and not (layer1_outputs(4231));
    layer2_outputs(2828) <= (layer1_outputs(167)) and (layer1_outputs(3876));
    layer2_outputs(2829) <= layer1_outputs(784);
    layer2_outputs(2830) <= not(layer1_outputs(3454));
    layer2_outputs(2831) <= not(layer1_outputs(3315));
    layer2_outputs(2832) <= not(layer1_outputs(2682)) or (layer1_outputs(2513));
    layer2_outputs(2833) <= not((layer1_outputs(943)) xor (layer1_outputs(3969)));
    layer2_outputs(2834) <= (layer1_outputs(4385)) xor (layer1_outputs(508));
    layer2_outputs(2835) <= not((layer1_outputs(2289)) and (layer1_outputs(291)));
    layer2_outputs(2836) <= not((layer1_outputs(1289)) or (layer1_outputs(923)));
    layer2_outputs(2837) <= not(layer1_outputs(3797)) or (layer1_outputs(3392));
    layer2_outputs(2838) <= not(layer1_outputs(3481));
    layer2_outputs(2839) <= layer1_outputs(1746);
    layer2_outputs(2840) <= not((layer1_outputs(1830)) or (layer1_outputs(3215)));
    layer2_outputs(2841) <= (layer1_outputs(2516)) and not (layer1_outputs(4967));
    layer2_outputs(2842) <= layer1_outputs(4708);
    layer2_outputs(2843) <= (layer1_outputs(2223)) and (layer1_outputs(4189));
    layer2_outputs(2844) <= not(layer1_outputs(3105));
    layer2_outputs(2845) <= (layer1_outputs(645)) and (layer1_outputs(1309));
    layer2_outputs(2846) <= (layer1_outputs(3738)) and not (layer1_outputs(1548));
    layer2_outputs(2847) <= layer1_outputs(73);
    layer2_outputs(2848) <= not(layer1_outputs(1978));
    layer2_outputs(2849) <= not((layer1_outputs(791)) xor (layer1_outputs(3720)));
    layer2_outputs(2850) <= not(layer1_outputs(1942));
    layer2_outputs(2851) <= layer1_outputs(1134);
    layer2_outputs(2852) <= (layer1_outputs(4577)) and (layer1_outputs(881));
    layer2_outputs(2853) <= layer1_outputs(760);
    layer2_outputs(2854) <= not(layer1_outputs(1022));
    layer2_outputs(2855) <= layer1_outputs(3170);
    layer2_outputs(2856) <= not(layer1_outputs(1161));
    layer2_outputs(2857) <= (layer1_outputs(795)) or (layer1_outputs(1767));
    layer2_outputs(2858) <= not(layer1_outputs(1666));
    layer2_outputs(2859) <= not(layer1_outputs(4544));
    layer2_outputs(2860) <= not((layer1_outputs(2806)) and (layer1_outputs(4369)));
    layer2_outputs(2861) <= not(layer1_outputs(4209));
    layer2_outputs(2862) <= (layer1_outputs(380)) and not (layer1_outputs(1260));
    layer2_outputs(2863) <= not(layer1_outputs(1190));
    layer2_outputs(2864) <= not(layer1_outputs(493)) or (layer1_outputs(5020));
    layer2_outputs(2865) <= layer1_outputs(1836);
    layer2_outputs(2866) <= not((layer1_outputs(2283)) xor (layer1_outputs(1530)));
    layer2_outputs(2867) <= not(layer1_outputs(154));
    layer2_outputs(2868) <= layer1_outputs(118);
    layer2_outputs(2869) <= (layer1_outputs(1505)) xor (layer1_outputs(4967));
    layer2_outputs(2870) <= layer1_outputs(4691);
    layer2_outputs(2871) <= layer1_outputs(4059);
    layer2_outputs(2872) <= layer1_outputs(2622);
    layer2_outputs(2873) <= (layer1_outputs(312)) or (layer1_outputs(4688));
    layer2_outputs(2874) <= layer1_outputs(1640);
    layer2_outputs(2875) <= layer1_outputs(1982);
    layer2_outputs(2876) <= not(layer1_outputs(615));
    layer2_outputs(2877) <= (layer1_outputs(1712)) and not (layer1_outputs(1575));
    layer2_outputs(2878) <= (layer1_outputs(4477)) or (layer1_outputs(1012));
    layer2_outputs(2879) <= not((layer1_outputs(2443)) and (layer1_outputs(3185)));
    layer2_outputs(2880) <= not(layer1_outputs(4336));
    layer2_outputs(2881) <= not(layer1_outputs(173)) or (layer1_outputs(99));
    layer2_outputs(2882) <= (layer1_outputs(1368)) and (layer1_outputs(2131));
    layer2_outputs(2883) <= not((layer1_outputs(4335)) or (layer1_outputs(1308)));
    layer2_outputs(2884) <= (layer1_outputs(4569)) and not (layer1_outputs(164));
    layer2_outputs(2885) <= layer1_outputs(4911);
    layer2_outputs(2886) <= not((layer1_outputs(1034)) or (layer1_outputs(4824)));
    layer2_outputs(2887) <= not((layer1_outputs(2708)) and (layer1_outputs(480)));
    layer2_outputs(2888) <= layer1_outputs(330);
    layer2_outputs(2889) <= (layer1_outputs(615)) or (layer1_outputs(4019));
    layer2_outputs(2890) <= layer1_outputs(2820);
    layer2_outputs(2891) <= not(layer1_outputs(3803));
    layer2_outputs(2892) <= (layer1_outputs(2875)) and not (layer1_outputs(3150));
    layer2_outputs(2893) <= not(layer1_outputs(3633)) or (layer1_outputs(3553));
    layer2_outputs(2894) <= (layer1_outputs(3550)) and not (layer1_outputs(1675));
    layer2_outputs(2895) <= not(layer1_outputs(9));
    layer2_outputs(2896) <= not((layer1_outputs(3251)) and (layer1_outputs(1356)));
    layer2_outputs(2897) <= (layer1_outputs(4076)) and (layer1_outputs(4298));
    layer2_outputs(2898) <= (layer1_outputs(565)) and not (layer1_outputs(4420));
    layer2_outputs(2899) <= not(layer1_outputs(1006));
    layer2_outputs(2900) <= (layer1_outputs(3936)) and (layer1_outputs(2210));
    layer2_outputs(2901) <= not((layer1_outputs(1237)) or (layer1_outputs(1821)));
    layer2_outputs(2902) <= not(layer1_outputs(42));
    layer2_outputs(2903) <= not((layer1_outputs(3122)) or (layer1_outputs(2816)));
    layer2_outputs(2904) <= (layer1_outputs(221)) and not (layer1_outputs(2879));
    layer2_outputs(2905) <= '0';
    layer2_outputs(2906) <= (layer1_outputs(3940)) xor (layer1_outputs(3521));
    layer2_outputs(2907) <= not(layer1_outputs(1881));
    layer2_outputs(2908) <= not(layer1_outputs(1542)) or (layer1_outputs(4999));
    layer2_outputs(2909) <= (layer1_outputs(153)) and not (layer1_outputs(3683));
    layer2_outputs(2910) <= not(layer1_outputs(4460));
    layer2_outputs(2911) <= layer1_outputs(2936);
    layer2_outputs(2912) <= (layer1_outputs(4746)) and not (layer1_outputs(369));
    layer2_outputs(2913) <= not((layer1_outputs(3658)) and (layer1_outputs(2195)));
    layer2_outputs(2914) <= not(layer1_outputs(428));
    layer2_outputs(2915) <= layer1_outputs(5027);
    layer2_outputs(2916) <= not((layer1_outputs(4937)) xor (layer1_outputs(4211)));
    layer2_outputs(2917) <= layer1_outputs(375);
    layer2_outputs(2918) <= not(layer1_outputs(3260));
    layer2_outputs(2919) <= not(layer1_outputs(1946)) or (layer1_outputs(3258));
    layer2_outputs(2920) <= (layer1_outputs(657)) and not (layer1_outputs(1853));
    layer2_outputs(2921) <= (layer1_outputs(3529)) xor (layer1_outputs(942));
    layer2_outputs(2922) <= layer1_outputs(3254);
    layer2_outputs(2923) <= layer1_outputs(4419);
    layer2_outputs(2924) <= (layer1_outputs(2434)) and (layer1_outputs(4444));
    layer2_outputs(2925) <= layer1_outputs(136);
    layer2_outputs(2926) <= layer1_outputs(2045);
    layer2_outputs(2927) <= (layer1_outputs(5108)) and not (layer1_outputs(4499));
    layer2_outputs(2928) <= (layer1_outputs(4237)) or (layer1_outputs(460));
    layer2_outputs(2929) <= (layer1_outputs(3023)) xor (layer1_outputs(4665));
    layer2_outputs(2930) <= layer1_outputs(92);
    layer2_outputs(2931) <= not((layer1_outputs(3952)) or (layer1_outputs(2458)));
    layer2_outputs(2932) <= layer1_outputs(4586);
    layer2_outputs(2933) <= not((layer1_outputs(1466)) or (layer1_outputs(306)));
    layer2_outputs(2934) <= layer1_outputs(2323);
    layer2_outputs(2935) <= layer1_outputs(1595);
    layer2_outputs(2936) <= not(layer1_outputs(3360));
    layer2_outputs(2937) <= not(layer1_outputs(708));
    layer2_outputs(2938) <= not(layer1_outputs(3250));
    layer2_outputs(2939) <= layer1_outputs(3560);
    layer2_outputs(2940) <= (layer1_outputs(4128)) xor (layer1_outputs(3253));
    layer2_outputs(2941) <= not(layer1_outputs(700));
    layer2_outputs(2942) <= not((layer1_outputs(4437)) or (layer1_outputs(1807)));
    layer2_outputs(2943) <= not(layer1_outputs(2778));
    layer2_outputs(2944) <= (layer1_outputs(940)) and not (layer1_outputs(1641));
    layer2_outputs(2945) <= not(layer1_outputs(4463));
    layer2_outputs(2946) <= layer1_outputs(4624);
    layer2_outputs(2947) <= (layer1_outputs(948)) or (layer1_outputs(4981));
    layer2_outputs(2948) <= layer1_outputs(4093);
    layer2_outputs(2949) <= not(layer1_outputs(104));
    layer2_outputs(2950) <= layer1_outputs(1976);
    layer2_outputs(2951) <= layer1_outputs(397);
    layer2_outputs(2952) <= not(layer1_outputs(1632));
    layer2_outputs(2953) <= not(layer1_outputs(2856));
    layer2_outputs(2954) <= (layer1_outputs(2235)) and (layer1_outputs(941));
    layer2_outputs(2955) <= not(layer1_outputs(3661)) or (layer1_outputs(2546));
    layer2_outputs(2956) <= layer1_outputs(1366);
    layer2_outputs(2957) <= layer1_outputs(2187);
    layer2_outputs(2958) <= (layer1_outputs(290)) xor (layer1_outputs(1112));
    layer2_outputs(2959) <= not(layer1_outputs(2502));
    layer2_outputs(2960) <= not(layer1_outputs(2686));
    layer2_outputs(2961) <= (layer1_outputs(543)) or (layer1_outputs(3361));
    layer2_outputs(2962) <= layer1_outputs(3027);
    layer2_outputs(2963) <= (layer1_outputs(2333)) and (layer1_outputs(1740));
    layer2_outputs(2964) <= not((layer1_outputs(2153)) and (layer1_outputs(2582)));
    layer2_outputs(2965) <= not(layer1_outputs(3169));
    layer2_outputs(2966) <= not((layer1_outputs(5023)) and (layer1_outputs(2324)));
    layer2_outputs(2967) <= not(layer1_outputs(4502)) or (layer1_outputs(1541));
    layer2_outputs(2968) <= not(layer1_outputs(4418));
    layer2_outputs(2969) <= not(layer1_outputs(3420));
    layer2_outputs(2970) <= not(layer1_outputs(463));
    layer2_outputs(2971) <= not(layer1_outputs(5077));
    layer2_outputs(2972) <= (layer1_outputs(3827)) and not (layer1_outputs(1640));
    layer2_outputs(2973) <= (layer1_outputs(3958)) and (layer1_outputs(1705));
    layer2_outputs(2974) <= '1';
    layer2_outputs(2975) <= not(layer1_outputs(1513));
    layer2_outputs(2976) <= (layer1_outputs(3991)) and not (layer1_outputs(3897));
    layer2_outputs(2977) <= (layer1_outputs(4431)) xor (layer1_outputs(143));
    layer2_outputs(2978) <= (layer1_outputs(5055)) and (layer1_outputs(2078));
    layer2_outputs(2979) <= not(layer1_outputs(3570)) or (layer1_outputs(4841));
    layer2_outputs(2980) <= layer1_outputs(3207);
    layer2_outputs(2981) <= not(layer1_outputs(559));
    layer2_outputs(2982) <= layer1_outputs(3923);
    layer2_outputs(2983) <= not(layer1_outputs(3532));
    layer2_outputs(2984) <= not(layer1_outputs(3653));
    layer2_outputs(2985) <= layer1_outputs(4289);
    layer2_outputs(2986) <= layer1_outputs(3311);
    layer2_outputs(2987) <= layer1_outputs(3376);
    layer2_outputs(2988) <= (layer1_outputs(1532)) xor (layer1_outputs(2851));
    layer2_outputs(2989) <= not((layer1_outputs(2092)) xor (layer1_outputs(440)));
    layer2_outputs(2990) <= not(layer1_outputs(1293));
    layer2_outputs(2991) <= not((layer1_outputs(953)) and (layer1_outputs(1776)));
    layer2_outputs(2992) <= layer1_outputs(4097);
    layer2_outputs(2993) <= not(layer1_outputs(625));
    layer2_outputs(2994) <= (layer1_outputs(1986)) or (layer1_outputs(3067));
    layer2_outputs(2995) <= layer1_outputs(4966);
    layer2_outputs(2996) <= not((layer1_outputs(1703)) xor (layer1_outputs(2582)));
    layer2_outputs(2997) <= not((layer1_outputs(1681)) xor (layer1_outputs(2291)));
    layer2_outputs(2998) <= not(layer1_outputs(5054));
    layer2_outputs(2999) <= not((layer1_outputs(344)) xor (layer1_outputs(186)));
    layer2_outputs(3000) <= (layer1_outputs(956)) and (layer1_outputs(5077));
    layer2_outputs(3001) <= not((layer1_outputs(2757)) and (layer1_outputs(1661)));
    layer2_outputs(3002) <= not(layer1_outputs(515)) or (layer1_outputs(4372));
    layer2_outputs(3003) <= '1';
    layer2_outputs(3004) <= not(layer1_outputs(2252));
    layer2_outputs(3005) <= layer1_outputs(3610);
    layer2_outputs(3006) <= (layer1_outputs(4431)) and not (layer1_outputs(2818));
    layer2_outputs(3007) <= (layer1_outputs(4150)) and not (layer1_outputs(4729));
    layer2_outputs(3008) <= layer1_outputs(239);
    layer2_outputs(3009) <= not(layer1_outputs(1380)) or (layer1_outputs(537));
    layer2_outputs(3010) <= (layer1_outputs(1464)) and (layer1_outputs(4735));
    layer2_outputs(3011) <= (layer1_outputs(1069)) and (layer1_outputs(1947));
    layer2_outputs(3012) <= not((layer1_outputs(3484)) xor (layer1_outputs(2462)));
    layer2_outputs(3013) <= '0';
    layer2_outputs(3014) <= not(layer1_outputs(811)) or (layer1_outputs(4539));
    layer2_outputs(3015) <= (layer1_outputs(3147)) xor (layer1_outputs(175));
    layer2_outputs(3016) <= (layer1_outputs(2211)) and not (layer1_outputs(945));
    layer2_outputs(3017) <= not((layer1_outputs(495)) xor (layer1_outputs(3854)));
    layer2_outputs(3018) <= (layer1_outputs(3667)) xor (layer1_outputs(497));
    layer2_outputs(3019) <= layer1_outputs(3542);
    layer2_outputs(3020) <= layer1_outputs(2566);
    layer2_outputs(3021) <= not(layer1_outputs(2953)) or (layer1_outputs(2986));
    layer2_outputs(3022) <= not(layer1_outputs(383));
    layer2_outputs(3023) <= (layer1_outputs(1921)) and not (layer1_outputs(1850));
    layer2_outputs(3024) <= layer1_outputs(715);
    layer2_outputs(3025) <= not((layer1_outputs(4858)) and (layer1_outputs(2267)));
    layer2_outputs(3026) <= layer1_outputs(1679);
    layer2_outputs(3027) <= not((layer1_outputs(2111)) or (layer1_outputs(3409)));
    layer2_outputs(3028) <= not(layer1_outputs(2642)) or (layer1_outputs(264));
    layer2_outputs(3029) <= layer1_outputs(5041);
    layer2_outputs(3030) <= not((layer1_outputs(542)) xor (layer1_outputs(3423)));
    layer2_outputs(3031) <= (layer1_outputs(4357)) or (layer1_outputs(3149));
    layer2_outputs(3032) <= layer1_outputs(4222);
    layer2_outputs(3033) <= (layer1_outputs(1694)) or (layer1_outputs(2146));
    layer2_outputs(3034) <= layer1_outputs(876);
    layer2_outputs(3035) <= not((layer1_outputs(3875)) and (layer1_outputs(2204)));
    layer2_outputs(3036) <= (layer1_outputs(1050)) and not (layer1_outputs(604));
    layer2_outputs(3037) <= layer1_outputs(2244);
    layer2_outputs(3038) <= not(layer1_outputs(3026)) or (layer1_outputs(210));
    layer2_outputs(3039) <= layer1_outputs(3534);
    layer2_outputs(3040) <= not(layer1_outputs(2044));
    layer2_outputs(3041) <= not((layer1_outputs(4105)) or (layer1_outputs(1369)));
    layer2_outputs(3042) <= not((layer1_outputs(4766)) xor (layer1_outputs(3676)));
    layer2_outputs(3043) <= not(layer1_outputs(2218));
    layer2_outputs(3044) <= not(layer1_outputs(4667));
    layer2_outputs(3045) <= layer1_outputs(2889);
    layer2_outputs(3046) <= not(layer1_outputs(4671));
    layer2_outputs(3047) <= layer1_outputs(4302);
    layer2_outputs(3048) <= layer1_outputs(2312);
    layer2_outputs(3049) <= not((layer1_outputs(2951)) and (layer1_outputs(5101)));
    layer2_outputs(3050) <= not((layer1_outputs(3724)) and (layer1_outputs(1734)));
    layer2_outputs(3051) <= not((layer1_outputs(4564)) or (layer1_outputs(137)));
    layer2_outputs(3052) <= not(layer1_outputs(3198));
    layer2_outputs(3053) <= (layer1_outputs(3383)) and not (layer1_outputs(4492));
    layer2_outputs(3054) <= not(layer1_outputs(354));
    layer2_outputs(3055) <= (layer1_outputs(2196)) and not (layer1_outputs(4196));
    layer2_outputs(3056) <= not(layer1_outputs(2265)) or (layer1_outputs(4559));
    layer2_outputs(3057) <= layer1_outputs(125);
    layer2_outputs(3058) <= (layer1_outputs(2876)) and not (layer1_outputs(4918));
    layer2_outputs(3059) <= layer1_outputs(1345);
    layer2_outputs(3060) <= not(layer1_outputs(782));
    layer2_outputs(3061) <= not(layer1_outputs(2407));
    layer2_outputs(3062) <= not(layer1_outputs(2963));
    layer2_outputs(3063) <= not(layer1_outputs(2240));
    layer2_outputs(3064) <= (layer1_outputs(4809)) xor (layer1_outputs(3501));
    layer2_outputs(3065) <= '0';
    layer2_outputs(3066) <= not(layer1_outputs(4551));
    layer2_outputs(3067) <= not((layer1_outputs(3507)) xor (layer1_outputs(1097)));
    layer2_outputs(3068) <= layer1_outputs(3908);
    layer2_outputs(3069) <= layer1_outputs(610);
    layer2_outputs(3070) <= layer1_outputs(4695);
    layer2_outputs(3071) <= not((layer1_outputs(4819)) xor (layer1_outputs(2108)));
    layer2_outputs(3072) <= not(layer1_outputs(2334));
    layer2_outputs(3073) <= not((layer1_outputs(5090)) or (layer1_outputs(2663)));
    layer2_outputs(3074) <= (layer1_outputs(2811)) and (layer1_outputs(1245));
    layer2_outputs(3075) <= not(layer1_outputs(42));
    layer2_outputs(3076) <= (layer1_outputs(1453)) xor (layer1_outputs(4044));
    layer2_outputs(3077) <= not(layer1_outputs(1583)) or (layer1_outputs(198));
    layer2_outputs(3078) <= not(layer1_outputs(511)) or (layer1_outputs(3809));
    layer2_outputs(3079) <= layer1_outputs(3293);
    layer2_outputs(3080) <= not(layer1_outputs(3947));
    layer2_outputs(3081) <= not((layer1_outputs(5076)) or (layer1_outputs(1270)));
    layer2_outputs(3082) <= not(layer1_outputs(2873));
    layer2_outputs(3083) <= (layer1_outputs(975)) xor (layer1_outputs(4262));
    layer2_outputs(3084) <= layer1_outputs(560);
    layer2_outputs(3085) <= layer1_outputs(562);
    layer2_outputs(3086) <= not(layer1_outputs(2084));
    layer2_outputs(3087) <= not((layer1_outputs(7)) and (layer1_outputs(3818)));
    layer2_outputs(3088) <= layer1_outputs(3975);
    layer2_outputs(3089) <= not(layer1_outputs(2481));
    layer2_outputs(3090) <= layer1_outputs(4791);
    layer2_outputs(3091) <= not(layer1_outputs(973));
    layer2_outputs(3092) <= not((layer1_outputs(3758)) or (layer1_outputs(1964)));
    layer2_outputs(3093) <= not(layer1_outputs(4574));
    layer2_outputs(3094) <= layer1_outputs(3628);
    layer2_outputs(3095) <= not(layer1_outputs(3281)) or (layer1_outputs(4202));
    layer2_outputs(3096) <= layer1_outputs(6);
    layer2_outputs(3097) <= not(layer1_outputs(193));
    layer2_outputs(3098) <= not(layer1_outputs(3873));
    layer2_outputs(3099) <= not(layer1_outputs(4726));
    layer2_outputs(3100) <= (layer1_outputs(1367)) or (layer1_outputs(1342));
    layer2_outputs(3101) <= (layer1_outputs(4633)) and (layer1_outputs(4874));
    layer2_outputs(3102) <= (layer1_outputs(2444)) or (layer1_outputs(5002));
    layer2_outputs(3103) <= layer1_outputs(4604);
    layer2_outputs(3104) <= layer1_outputs(1826);
    layer2_outputs(3105) <= layer1_outputs(1647);
    layer2_outputs(3106) <= not(layer1_outputs(4057));
    layer2_outputs(3107) <= not(layer1_outputs(408));
    layer2_outputs(3108) <= layer1_outputs(3468);
    layer2_outputs(3109) <= not((layer1_outputs(1608)) or (layer1_outputs(3229)));
    layer2_outputs(3110) <= not((layer1_outputs(1390)) xor (layer1_outputs(4731)));
    layer2_outputs(3111) <= not(layer1_outputs(2775)) or (layer1_outputs(3577));
    layer2_outputs(3112) <= not(layer1_outputs(978));
    layer2_outputs(3113) <= not(layer1_outputs(2458));
    layer2_outputs(3114) <= (layer1_outputs(1236)) and not (layer1_outputs(2661));
    layer2_outputs(3115) <= (layer1_outputs(4413)) xor (layer1_outputs(2052));
    layer2_outputs(3116) <= not(layer1_outputs(966));
    layer2_outputs(3117) <= (layer1_outputs(3854)) or (layer1_outputs(3640));
    layer2_outputs(3118) <= (layer1_outputs(1740)) and (layer1_outputs(2691));
    layer2_outputs(3119) <= (layer1_outputs(2639)) xor (layer1_outputs(1203));
    layer2_outputs(3120) <= not(layer1_outputs(1548));
    layer2_outputs(3121) <= not(layer1_outputs(884));
    layer2_outputs(3122) <= not(layer1_outputs(4259)) or (layer1_outputs(4185));
    layer2_outputs(3123) <= not(layer1_outputs(4516));
    layer2_outputs(3124) <= not(layer1_outputs(3067)) or (layer1_outputs(2095));
    layer2_outputs(3125) <= not(layer1_outputs(1841)) or (layer1_outputs(578));
    layer2_outputs(3126) <= not((layer1_outputs(2413)) or (layer1_outputs(858)));
    layer2_outputs(3127) <= (layer1_outputs(2545)) and (layer1_outputs(2215));
    layer2_outputs(3128) <= not((layer1_outputs(1872)) and (layer1_outputs(1003)));
    layer2_outputs(3129) <= not(layer1_outputs(744));
    layer2_outputs(3130) <= layer1_outputs(1153);
    layer2_outputs(3131) <= not((layer1_outputs(797)) and (layer1_outputs(633)));
    layer2_outputs(3132) <= (layer1_outputs(2429)) xor (layer1_outputs(4484));
    layer2_outputs(3133) <= layer1_outputs(4116);
    layer2_outputs(3134) <= (layer1_outputs(288)) and not (layer1_outputs(716));
    layer2_outputs(3135) <= not((layer1_outputs(4166)) or (layer1_outputs(2746)));
    layer2_outputs(3136) <= not(layer1_outputs(4072)) or (layer1_outputs(3761));
    layer2_outputs(3137) <= (layer1_outputs(1307)) or (layer1_outputs(2336));
    layer2_outputs(3138) <= not(layer1_outputs(1496));
    layer2_outputs(3139) <= not((layer1_outputs(750)) xor (layer1_outputs(4094)));
    layer2_outputs(3140) <= not(layer1_outputs(4948));
    layer2_outputs(3141) <= (layer1_outputs(2505)) and not (layer1_outputs(461));
    layer2_outputs(3142) <= layer1_outputs(1501);
    layer2_outputs(3143) <= not(layer1_outputs(1639));
    layer2_outputs(3144) <= not(layer1_outputs(3212));
    layer2_outputs(3145) <= not(layer1_outputs(982));
    layer2_outputs(3146) <= layer1_outputs(4565);
    layer2_outputs(3147) <= (layer1_outputs(658)) or (layer1_outputs(3210));
    layer2_outputs(3148) <= not((layer1_outputs(4850)) xor (layer1_outputs(2401)));
    layer2_outputs(3149) <= '0';
    layer2_outputs(3150) <= layer1_outputs(987);
    layer2_outputs(3151) <= (layer1_outputs(4280)) xor (layer1_outputs(3793));
    layer2_outputs(3152) <= layer1_outputs(1631);
    layer2_outputs(3153) <= layer1_outputs(4283);
    layer2_outputs(3154) <= not(layer1_outputs(2163));
    layer2_outputs(3155) <= not((layer1_outputs(3314)) xor (layer1_outputs(3959)));
    layer2_outputs(3156) <= '0';
    layer2_outputs(3157) <= not(layer1_outputs(1219)) or (layer1_outputs(5057));
    layer2_outputs(3158) <= not(layer1_outputs(4714));
    layer2_outputs(3159) <= not(layer1_outputs(456));
    layer2_outputs(3160) <= not((layer1_outputs(4105)) xor (layer1_outputs(2203)));
    layer2_outputs(3161) <= not(layer1_outputs(745));
    layer2_outputs(3162) <= not(layer1_outputs(2771));
    layer2_outputs(3163) <= not((layer1_outputs(4094)) xor (layer1_outputs(1965)));
    layer2_outputs(3164) <= (layer1_outputs(4961)) or (layer1_outputs(3061));
    layer2_outputs(3165) <= (layer1_outputs(2660)) and not (layer1_outputs(4205));
    layer2_outputs(3166) <= (layer1_outputs(4777)) and not (layer1_outputs(2662));
    layer2_outputs(3167) <= layer1_outputs(4454);
    layer2_outputs(3168) <= layer1_outputs(2272);
    layer2_outputs(3169) <= not((layer1_outputs(3893)) and (layer1_outputs(820)));
    layer2_outputs(3170) <= layer1_outputs(352);
    layer2_outputs(3171) <= '1';
    layer2_outputs(3172) <= not(layer1_outputs(1098));
    layer2_outputs(3173) <= layer1_outputs(4549);
    layer2_outputs(3174) <= not((layer1_outputs(4098)) or (layer1_outputs(984)));
    layer2_outputs(3175) <= (layer1_outputs(2494)) xor (layer1_outputs(2068));
    layer2_outputs(3176) <= layer1_outputs(2564);
    layer2_outputs(3177) <= not(layer1_outputs(583)) or (layer1_outputs(1023));
    layer2_outputs(3178) <= not(layer1_outputs(2546));
    layer2_outputs(3179) <= not(layer1_outputs(2973));
    layer2_outputs(3180) <= not(layer1_outputs(736)) or (layer1_outputs(896));
    layer2_outputs(3181) <= layer1_outputs(194);
    layer2_outputs(3182) <= (layer1_outputs(4008)) and not (layer1_outputs(1276));
    layer2_outputs(3183) <= layer1_outputs(1585);
    layer2_outputs(3184) <= layer1_outputs(100);
    layer2_outputs(3185) <= (layer1_outputs(4743)) and (layer1_outputs(2308));
    layer2_outputs(3186) <= not((layer1_outputs(2007)) xor (layer1_outputs(2592)));
    layer2_outputs(3187) <= layer1_outputs(1567);
    layer2_outputs(3188) <= (layer1_outputs(2916)) and not (layer1_outputs(1635));
    layer2_outputs(3189) <= layer1_outputs(1854);
    layer2_outputs(3190) <= (layer1_outputs(1078)) and not (layer1_outputs(3006));
    layer2_outputs(3191) <= not(layer1_outputs(393));
    layer2_outputs(3192) <= (layer1_outputs(1009)) or (layer1_outputs(3457));
    layer2_outputs(3193) <= layer1_outputs(2583);
    layer2_outputs(3194) <= layer1_outputs(223);
    layer2_outputs(3195) <= layer1_outputs(2739);
    layer2_outputs(3196) <= not(layer1_outputs(534));
    layer2_outputs(3197) <= not(layer1_outputs(1865));
    layer2_outputs(3198) <= (layer1_outputs(4041)) and not (layer1_outputs(3808));
    layer2_outputs(3199) <= (layer1_outputs(142)) xor (layer1_outputs(2949));
    layer2_outputs(3200) <= layer1_outputs(4144);
    layer2_outputs(3201) <= not(layer1_outputs(2031)) or (layer1_outputs(1830));
    layer2_outputs(3202) <= not((layer1_outputs(1100)) or (layer1_outputs(1907)));
    layer2_outputs(3203) <= not(layer1_outputs(3108));
    layer2_outputs(3204) <= not(layer1_outputs(19));
    layer2_outputs(3205) <= not(layer1_outputs(1997));
    layer2_outputs(3206) <= not((layer1_outputs(1607)) xor (layer1_outputs(4840)));
    layer2_outputs(3207) <= '1';
    layer2_outputs(3208) <= layer1_outputs(2854);
    layer2_outputs(3209) <= '0';
    layer2_outputs(3210) <= not(layer1_outputs(2532));
    layer2_outputs(3211) <= not((layer1_outputs(3624)) xor (layer1_outputs(738)));
    layer2_outputs(3212) <= layer1_outputs(3851);
    layer2_outputs(3213) <= not(layer1_outputs(1374));
    layer2_outputs(3214) <= layer1_outputs(247);
    layer2_outputs(3215) <= not(layer1_outputs(3539)) or (layer1_outputs(4088));
    layer2_outputs(3216) <= (layer1_outputs(370)) and not (layer1_outputs(4069));
    layer2_outputs(3217) <= layer1_outputs(4491);
    layer2_outputs(3218) <= not(layer1_outputs(4254));
    layer2_outputs(3219) <= layer1_outputs(3760);
    layer2_outputs(3220) <= layer1_outputs(2340);
    layer2_outputs(3221) <= not(layer1_outputs(441));
    layer2_outputs(3222) <= not((layer1_outputs(1914)) and (layer1_outputs(3595)));
    layer2_outputs(3223) <= layer1_outputs(1446);
    layer2_outputs(3224) <= not((layer1_outputs(1447)) and (layer1_outputs(374)));
    layer2_outputs(3225) <= not((layer1_outputs(3276)) or (layer1_outputs(0)));
    layer2_outputs(3226) <= layer1_outputs(3121);
    layer2_outputs(3227) <= (layer1_outputs(2431)) xor (layer1_outputs(3755));
    layer2_outputs(3228) <= layer1_outputs(960);
    layer2_outputs(3229) <= layer1_outputs(1239);
    layer2_outputs(3230) <= (layer1_outputs(3063)) and not (layer1_outputs(1043));
    layer2_outputs(3231) <= not(layer1_outputs(3628)) or (layer1_outputs(4233));
    layer2_outputs(3232) <= not(layer1_outputs(570));
    layer2_outputs(3233) <= not(layer1_outputs(1847)) or (layer1_outputs(4328));
    layer2_outputs(3234) <= (layer1_outputs(1058)) and (layer1_outputs(2925));
    layer2_outputs(3235) <= not((layer1_outputs(2495)) or (layer1_outputs(391)));
    layer2_outputs(3236) <= (layer1_outputs(1478)) and (layer1_outputs(4870));
    layer2_outputs(3237) <= not(layer1_outputs(48)) or (layer1_outputs(2489));
    layer2_outputs(3238) <= (layer1_outputs(3436)) and (layer1_outputs(2769));
    layer2_outputs(3239) <= not((layer1_outputs(1790)) xor (layer1_outputs(3227)));
    layer2_outputs(3240) <= (layer1_outputs(841)) and not (layer1_outputs(3644));
    layer2_outputs(3241) <= not((layer1_outputs(328)) or (layer1_outputs(3677)));
    layer2_outputs(3242) <= layer1_outputs(3257);
    layer2_outputs(3243) <= layer1_outputs(4812);
    layer2_outputs(3244) <= layer1_outputs(4800);
    layer2_outputs(3245) <= layer1_outputs(692);
    layer2_outputs(3246) <= layer1_outputs(2780);
    layer2_outputs(3247) <= (layer1_outputs(288)) and not (layer1_outputs(3746));
    layer2_outputs(3248) <= layer1_outputs(4275);
    layer2_outputs(3249) <= not(layer1_outputs(1719));
    layer2_outputs(3250) <= not(layer1_outputs(746));
    layer2_outputs(3251) <= not(layer1_outputs(4013)) or (layer1_outputs(3891));
    layer2_outputs(3252) <= (layer1_outputs(4184)) xor (layer1_outputs(3793));
    layer2_outputs(3253) <= not(layer1_outputs(2482));
    layer2_outputs(3254) <= layer1_outputs(2832);
    layer2_outputs(3255) <= layer1_outputs(1369);
    layer2_outputs(3256) <= layer1_outputs(4359);
    layer2_outputs(3257) <= not(layer1_outputs(2714));
    layer2_outputs(3258) <= layer1_outputs(2270);
    layer2_outputs(3259) <= layer1_outputs(3923);
    layer2_outputs(3260) <= not(layer1_outputs(1030));
    layer2_outputs(3261) <= (layer1_outputs(464)) or (layer1_outputs(3606));
    layer2_outputs(3262) <= layer1_outputs(4884);
    layer2_outputs(3263) <= (layer1_outputs(3279)) and not (layer1_outputs(3104));
    layer2_outputs(3264) <= (layer1_outputs(1710)) or (layer1_outputs(2896));
    layer2_outputs(3265) <= not(layer1_outputs(2211)) or (layer1_outputs(885));
    layer2_outputs(3266) <= (layer1_outputs(5051)) and not (layer1_outputs(1210));
    layer2_outputs(3267) <= (layer1_outputs(584)) and not (layer1_outputs(656));
    layer2_outputs(3268) <= not(layer1_outputs(2602));
    layer2_outputs(3269) <= not((layer1_outputs(132)) and (layer1_outputs(2259)));
    layer2_outputs(3270) <= not((layer1_outputs(4290)) and (layer1_outputs(557)));
    layer2_outputs(3271) <= (layer1_outputs(1142)) xor (layer1_outputs(1247));
    layer2_outputs(3272) <= not((layer1_outputs(2790)) xor (layer1_outputs(748)));
    layer2_outputs(3273) <= layer1_outputs(4443);
    layer2_outputs(3274) <= (layer1_outputs(4030)) or (layer1_outputs(4959));
    layer2_outputs(3275) <= not(layer1_outputs(3256));
    layer2_outputs(3276) <= not(layer1_outputs(4447)) or (layer1_outputs(1678));
    layer2_outputs(3277) <= not(layer1_outputs(3998));
    layer2_outputs(3278) <= layer1_outputs(3871);
    layer2_outputs(3279) <= layer1_outputs(2360);
    layer2_outputs(3280) <= (layer1_outputs(4080)) and not (layer1_outputs(4289));
    layer2_outputs(3281) <= (layer1_outputs(1200)) and not (layer1_outputs(1255));
    layer2_outputs(3282) <= '0';
    layer2_outputs(3283) <= (layer1_outputs(4866)) or (layer1_outputs(714));
    layer2_outputs(3284) <= not(layer1_outputs(887));
    layer2_outputs(3285) <= not(layer1_outputs(1294));
    layer2_outputs(3286) <= not((layer1_outputs(1288)) or (layer1_outputs(4996)));
    layer2_outputs(3287) <= layer1_outputs(1196);
    layer2_outputs(3288) <= not(layer1_outputs(67));
    layer2_outputs(3289) <= not(layer1_outputs(1835)) or (layer1_outputs(2234));
    layer2_outputs(3290) <= layer1_outputs(753);
    layer2_outputs(3291) <= layer1_outputs(4511);
    layer2_outputs(3292) <= (layer1_outputs(694)) and not (layer1_outputs(1117));
    layer2_outputs(3293) <= not((layer1_outputs(1059)) xor (layer1_outputs(4278)));
    layer2_outputs(3294) <= (layer1_outputs(4056)) xor (layer1_outputs(2559));
    layer2_outputs(3295) <= not(layer1_outputs(4935));
    layer2_outputs(3296) <= not((layer1_outputs(3097)) or (layer1_outputs(3306)));
    layer2_outputs(3297) <= not(layer1_outputs(1873)) or (layer1_outputs(767));
    layer2_outputs(3298) <= (layer1_outputs(1741)) and (layer1_outputs(4586));
    layer2_outputs(3299) <= not(layer1_outputs(3679));
    layer2_outputs(3300) <= layer1_outputs(1268);
    layer2_outputs(3301) <= not(layer1_outputs(835)) or (layer1_outputs(572));
    layer2_outputs(3302) <= not(layer1_outputs(1144));
    layer2_outputs(3303) <= not((layer1_outputs(564)) or (layer1_outputs(764)));
    layer2_outputs(3304) <= layer1_outputs(1552);
    layer2_outputs(3305) <= not(layer1_outputs(1630)) or (layer1_outputs(4164));
    layer2_outputs(3306) <= layer1_outputs(2387);
    layer2_outputs(3307) <= not(layer1_outputs(3092));
    layer2_outputs(3308) <= layer1_outputs(346);
    layer2_outputs(3309) <= not(layer1_outputs(3446)) or (layer1_outputs(3602));
    layer2_outputs(3310) <= layer1_outputs(2650);
    layer2_outputs(3311) <= (layer1_outputs(3589)) and not (layer1_outputs(2547));
    layer2_outputs(3312) <= not((layer1_outputs(38)) or (layer1_outputs(1221)));
    layer2_outputs(3313) <= not(layer1_outputs(1028));
    layer2_outputs(3314) <= not(layer1_outputs(3031));
    layer2_outputs(3315) <= layer1_outputs(1594);
    layer2_outputs(3316) <= layer1_outputs(2898);
    layer2_outputs(3317) <= layer1_outputs(1715);
    layer2_outputs(3318) <= layer1_outputs(993);
    layer2_outputs(3319) <= not(layer1_outputs(4533));
    layer2_outputs(3320) <= layer1_outputs(1796);
    layer2_outputs(3321) <= not(layer1_outputs(332));
    layer2_outputs(3322) <= (layer1_outputs(4310)) xor (layer1_outputs(1573));
    layer2_outputs(3323) <= (layer1_outputs(1745)) and not (layer1_outputs(1481));
    layer2_outputs(3324) <= not(layer1_outputs(3379));
    layer2_outputs(3325) <= not((layer1_outputs(4121)) or (layer1_outputs(1093)));
    layer2_outputs(3326) <= layer1_outputs(4648);
    layer2_outputs(3327) <= not((layer1_outputs(3984)) xor (layer1_outputs(3131)));
    layer2_outputs(3328) <= layer1_outputs(2824);
    layer2_outputs(3329) <= (layer1_outputs(2682)) or (layer1_outputs(3353));
    layer2_outputs(3330) <= layer1_outputs(218);
    layer2_outputs(3331) <= (layer1_outputs(3087)) and not (layer1_outputs(84));
    layer2_outputs(3332) <= (layer1_outputs(1290)) and not (layer1_outputs(1416));
    layer2_outputs(3333) <= not((layer1_outputs(1315)) xor (layer1_outputs(4301)));
    layer2_outputs(3334) <= not(layer1_outputs(1136));
    layer2_outputs(3335) <= (layer1_outputs(4754)) or (layer1_outputs(625));
    layer2_outputs(3336) <= (layer1_outputs(2133)) xor (layer1_outputs(4476));
    layer2_outputs(3337) <= (layer1_outputs(5092)) or (layer1_outputs(2694));
    layer2_outputs(3338) <= layer1_outputs(1411);
    layer2_outputs(3339) <= (layer1_outputs(5070)) and not (layer1_outputs(2399));
    layer2_outputs(3340) <= (layer1_outputs(155)) or (layer1_outputs(3066));
    layer2_outputs(3341) <= layer1_outputs(935);
    layer2_outputs(3342) <= not((layer1_outputs(4525)) xor (layer1_outputs(1722)));
    layer2_outputs(3343) <= (layer1_outputs(1957)) and (layer1_outputs(4847));
    layer2_outputs(3344) <= (layer1_outputs(4596)) and not (layer1_outputs(4189));
    layer2_outputs(3345) <= (layer1_outputs(917)) and not (layer1_outputs(689));
    layer2_outputs(3346) <= (layer1_outputs(3889)) and (layer1_outputs(1363));
    layer2_outputs(3347) <= layer1_outputs(1494);
    layer2_outputs(3348) <= (layer1_outputs(4043)) and not (layer1_outputs(35));
    layer2_outputs(3349) <= not(layer1_outputs(2878)) or (layer1_outputs(286));
    layer2_outputs(3350) <= not(layer1_outputs(2078)) or (layer1_outputs(811));
    layer2_outputs(3351) <= '0';
    layer2_outputs(3352) <= (layer1_outputs(1884)) xor (layer1_outputs(1258));
    layer2_outputs(3353) <= (layer1_outputs(449)) and not (layer1_outputs(1998));
    layer2_outputs(3354) <= layer1_outputs(3881);
    layer2_outputs(3355) <= (layer1_outputs(1769)) xor (layer1_outputs(853));
    layer2_outputs(3356) <= not(layer1_outputs(1550));
    layer2_outputs(3357) <= (layer1_outputs(124)) and not (layer1_outputs(4344));
    layer2_outputs(3358) <= not((layer1_outputs(4388)) xor (layer1_outputs(4976)));
    layer2_outputs(3359) <= not(layer1_outputs(2634));
    layer2_outputs(3360) <= not((layer1_outputs(4913)) or (layer1_outputs(1148)));
    layer2_outputs(3361) <= layer1_outputs(3699);
    layer2_outputs(3362) <= (layer1_outputs(3520)) or (layer1_outputs(4762));
    layer2_outputs(3363) <= (layer1_outputs(4345)) and not (layer1_outputs(4453));
    layer2_outputs(3364) <= (layer1_outputs(3753)) xor (layer1_outputs(3457));
    layer2_outputs(3365) <= not(layer1_outputs(73));
    layer2_outputs(3366) <= layer1_outputs(1454);
    layer2_outputs(3367) <= (layer1_outputs(2349)) and (layer1_outputs(4904));
    layer2_outputs(3368) <= not((layer1_outputs(3899)) or (layer1_outputs(755)));
    layer2_outputs(3369) <= (layer1_outputs(3391)) and not (layer1_outputs(4531));
    layer2_outputs(3370) <= (layer1_outputs(1316)) and not (layer1_outputs(2330));
    layer2_outputs(3371) <= (layer1_outputs(3418)) and (layer1_outputs(4123));
    layer2_outputs(3372) <= (layer1_outputs(4311)) xor (layer1_outputs(521));
    layer2_outputs(3373) <= (layer1_outputs(4246)) xor (layer1_outputs(4955));
    layer2_outputs(3374) <= layer1_outputs(432);
    layer2_outputs(3375) <= (layer1_outputs(4253)) and (layer1_outputs(26));
    layer2_outputs(3376) <= not(layer1_outputs(4908)) or (layer1_outputs(1331));
    layer2_outputs(3377) <= (layer1_outputs(3905)) and (layer1_outputs(837));
    layer2_outputs(3378) <= layer1_outputs(3529);
    layer2_outputs(3379) <= layer1_outputs(624);
    layer2_outputs(3380) <= layer1_outputs(2515);
    layer2_outputs(3381) <= not(layer1_outputs(2376)) or (layer1_outputs(3686));
    layer2_outputs(3382) <= not((layer1_outputs(693)) xor (layer1_outputs(169)));
    layer2_outputs(3383) <= not((layer1_outputs(368)) xor (layer1_outputs(4287)));
    layer2_outputs(3384) <= not((layer1_outputs(2767)) xor (layer1_outputs(1938)));
    layer2_outputs(3385) <= not(layer1_outputs(3829));
    layer2_outputs(3386) <= layer1_outputs(2670);
    layer2_outputs(3387) <= layer1_outputs(3302);
    layer2_outputs(3388) <= not(layer1_outputs(2328));
    layer2_outputs(3389) <= not((layer1_outputs(4264)) xor (layer1_outputs(3689)));
    layer2_outputs(3390) <= not(layer1_outputs(481));
    layer2_outputs(3391) <= layer1_outputs(4002);
    layer2_outputs(3392) <= (layer1_outputs(1312)) and (layer1_outputs(1475));
    layer2_outputs(3393) <= (layer1_outputs(1229)) xor (layer1_outputs(2834));
    layer2_outputs(3394) <= not(layer1_outputs(2094)) or (layer1_outputs(4079));
    layer2_outputs(3395) <= '0';
    layer2_outputs(3396) <= not((layer1_outputs(23)) or (layer1_outputs(96)));
    layer2_outputs(3397) <= not(layer1_outputs(1128));
    layer2_outputs(3398) <= (layer1_outputs(4989)) xor (layer1_outputs(3590));
    layer2_outputs(3399) <= not((layer1_outputs(1272)) xor (layer1_outputs(612)));
    layer2_outputs(3400) <= not(layer1_outputs(1207));
    layer2_outputs(3401) <= (layer1_outputs(1228)) xor (layer1_outputs(1759));
    layer2_outputs(3402) <= not(layer1_outputs(2971));
    layer2_outputs(3403) <= not((layer1_outputs(4794)) xor (layer1_outputs(2576)));
    layer2_outputs(3404) <= (layer1_outputs(183)) and (layer1_outputs(3741));
    layer2_outputs(3405) <= not(layer1_outputs(4177));
    layer2_outputs(3406) <= (layer1_outputs(3626)) and (layer1_outputs(2089));
    layer2_outputs(3407) <= (layer1_outputs(2209)) xor (layer1_outputs(3790));
    layer2_outputs(3408) <= not(layer1_outputs(1249)) or (layer1_outputs(4195));
    layer2_outputs(3409) <= not((layer1_outputs(4277)) xor (layer1_outputs(2579)));
    layer2_outputs(3410) <= not(layer1_outputs(2871));
    layer2_outputs(3411) <= layer1_outputs(240);
    layer2_outputs(3412) <= not(layer1_outputs(1620));
    layer2_outputs(3413) <= not((layer1_outputs(2077)) or (layer1_outputs(2723)));
    layer2_outputs(3414) <= (layer1_outputs(4670)) and (layer1_outputs(4292));
    layer2_outputs(3415) <= layer1_outputs(1712);
    layer2_outputs(3416) <= layer1_outputs(2751);
    layer2_outputs(3417) <= layer1_outputs(3869);
    layer2_outputs(3418) <= not(layer1_outputs(2710));
    layer2_outputs(3419) <= not(layer1_outputs(454));
    layer2_outputs(3420) <= (layer1_outputs(2109)) xor (layer1_outputs(2235));
    layer2_outputs(3421) <= not((layer1_outputs(2154)) or (layer1_outputs(985)));
    layer2_outputs(3422) <= not(layer1_outputs(5035));
    layer2_outputs(3423) <= not(layer1_outputs(3740)) or (layer1_outputs(1724));
    layer2_outputs(3424) <= layer1_outputs(2075);
    layer2_outputs(3425) <= not(layer1_outputs(1503));
    layer2_outputs(3426) <= not(layer1_outputs(967));
    layer2_outputs(3427) <= (layer1_outputs(2026)) or (layer1_outputs(4654));
    layer2_outputs(3428) <= not(layer1_outputs(3327)) or (layer1_outputs(554));
    layer2_outputs(3429) <= (layer1_outputs(1155)) and not (layer1_outputs(1387));
    layer2_outputs(3430) <= layer1_outputs(631);
    layer2_outputs(3431) <= not(layer1_outputs(3358));
    layer2_outputs(3432) <= (layer1_outputs(4173)) and (layer1_outputs(4383));
    layer2_outputs(3433) <= not((layer1_outputs(4660)) xor (layer1_outputs(3073)));
    layer2_outputs(3434) <= not(layer1_outputs(4055));
    layer2_outputs(3435) <= not(layer1_outputs(2560)) or (layer1_outputs(2283));
    layer2_outputs(3436) <= '1';
    layer2_outputs(3437) <= layer1_outputs(4622);
    layer2_outputs(3438) <= (layer1_outputs(1832)) and not (layer1_outputs(4887));
    layer2_outputs(3439) <= not(layer1_outputs(2791)) or (layer1_outputs(1899));
    layer2_outputs(3440) <= not(layer1_outputs(1011));
    layer2_outputs(3441) <= (layer1_outputs(4547)) and not (layer1_outputs(1627));
    layer2_outputs(3442) <= layer1_outputs(1412);
    layer2_outputs(3443) <= not(layer1_outputs(3014));
    layer2_outputs(3444) <= not(layer1_outputs(4877));
    layer2_outputs(3445) <= (layer1_outputs(3913)) xor (layer1_outputs(3912));
    layer2_outputs(3446) <= not(layer1_outputs(3690));
    layer2_outputs(3447) <= not(layer1_outputs(3421)) or (layer1_outputs(373));
    layer2_outputs(3448) <= not(layer1_outputs(833));
    layer2_outputs(3449) <= not(layer1_outputs(3034));
    layer2_outputs(3450) <= '1';
    layer2_outputs(3451) <= layer1_outputs(4065);
    layer2_outputs(3452) <= not(layer1_outputs(1883)) or (layer1_outputs(469));
    layer2_outputs(3453) <= not(layer1_outputs(3466));
    layer2_outputs(3454) <= not((layer1_outputs(2130)) and (layer1_outputs(2385)));
    layer2_outputs(3455) <= not(layer1_outputs(5050));
    layer2_outputs(3456) <= (layer1_outputs(3266)) xor (layer1_outputs(4585));
    layer2_outputs(3457) <= layer1_outputs(2123);
    layer2_outputs(3458) <= not(layer1_outputs(1384));
    layer2_outputs(3459) <= not(layer1_outputs(4522)) or (layer1_outputs(2783));
    layer2_outputs(3460) <= not((layer1_outputs(3380)) xor (layer1_outputs(813)));
    layer2_outputs(3461) <= not(layer1_outputs(3971)) or (layer1_outputs(1189));
    layer2_outputs(3462) <= (layer1_outputs(1086)) and not (layer1_outputs(2184));
    layer2_outputs(3463) <= not(layer1_outputs(2749));
    layer2_outputs(3464) <= layer1_outputs(539);
    layer2_outputs(3465) <= not((layer1_outputs(3437)) and (layer1_outputs(3495)));
    layer2_outputs(3466) <= not(layer1_outputs(4306));
    layer2_outputs(3467) <= (layer1_outputs(1533)) and (layer1_outputs(3033));
    layer2_outputs(3468) <= (layer1_outputs(1271)) and not (layer1_outputs(3350));
    layer2_outputs(3469) <= layer1_outputs(1725);
    layer2_outputs(3470) <= layer1_outputs(1499);
    layer2_outputs(3471) <= not(layer1_outputs(637));
    layer2_outputs(3472) <= layer1_outputs(36);
    layer2_outputs(3473) <= layer1_outputs(1586);
    layer2_outputs(3474) <= not((layer1_outputs(521)) xor (layer1_outputs(1899)));
    layer2_outputs(3475) <= (layer1_outputs(4402)) or (layer1_outputs(4559));
    layer2_outputs(3476) <= not((layer1_outputs(2149)) or (layer1_outputs(4740)));
    layer2_outputs(3477) <= (layer1_outputs(3749)) and (layer1_outputs(1487));
    layer2_outputs(3478) <= not(layer1_outputs(4881));
    layer2_outputs(3479) <= not(layer1_outputs(489));
    layer2_outputs(3480) <= (layer1_outputs(3913)) and not (layer1_outputs(29));
    layer2_outputs(3481) <= not(layer1_outputs(4739));
    layer2_outputs(3482) <= (layer1_outputs(659)) and not (layer1_outputs(3075));
    layer2_outputs(3483) <= not((layer1_outputs(1469)) or (layer1_outputs(989)));
    layer2_outputs(3484) <= layer1_outputs(2195);
    layer2_outputs(3485) <= not(layer1_outputs(4267));
    layer2_outputs(3486) <= layer1_outputs(441);
    layer2_outputs(3487) <= not(layer1_outputs(600));
    layer2_outputs(3488) <= (layer1_outputs(4712)) or (layer1_outputs(3368));
    layer2_outputs(3489) <= (layer1_outputs(215)) or (layer1_outputs(4962));
    layer2_outputs(3490) <= not(layer1_outputs(5010)) or (layer1_outputs(2990));
    layer2_outputs(3491) <= layer1_outputs(2064);
    layer2_outputs(3492) <= not((layer1_outputs(2577)) xor (layer1_outputs(1370)));
    layer2_outputs(3493) <= (layer1_outputs(2520)) or (layer1_outputs(3378));
    layer2_outputs(3494) <= (layer1_outputs(4745)) xor (layer1_outputs(1197));
    layer2_outputs(3495) <= (layer1_outputs(1096)) xor (layer1_outputs(4465));
    layer2_outputs(3496) <= (layer1_outputs(4282)) or (layer1_outputs(2206));
    layer2_outputs(3497) <= (layer1_outputs(5072)) and (layer1_outputs(4180));
    layer2_outputs(3498) <= not(layer1_outputs(3154)) or (layer1_outputs(3013));
    layer2_outputs(3499) <= not(layer1_outputs(2560)) or (layer1_outputs(3650));
    layer2_outputs(3500) <= not(layer1_outputs(3290));
    layer2_outputs(3501) <= not(layer1_outputs(1688));
    layer2_outputs(3502) <= (layer1_outputs(1593)) xor (layer1_outputs(2589));
    layer2_outputs(3503) <= layer1_outputs(1502);
    layer2_outputs(3504) <= not(layer1_outputs(1724));
    layer2_outputs(3505) <= layer1_outputs(3489);
    layer2_outputs(3506) <= layer1_outputs(3449);
    layer2_outputs(3507) <= (layer1_outputs(4375)) or (layer1_outputs(945));
    layer2_outputs(3508) <= not((layer1_outputs(2705)) or (layer1_outputs(2003)));
    layer2_outputs(3509) <= '0';
    layer2_outputs(3510) <= layer1_outputs(3582);
    layer2_outputs(3511) <= (layer1_outputs(4392)) and not (layer1_outputs(238));
    layer2_outputs(3512) <= layer1_outputs(2603);
    layer2_outputs(3513) <= layer1_outputs(591);
    layer2_outputs(3514) <= not((layer1_outputs(3870)) xor (layer1_outputs(3731)));
    layer2_outputs(3515) <= not(layer1_outputs(4248));
    layer2_outputs(3516) <= layer1_outputs(2678);
    layer2_outputs(3517) <= (layer1_outputs(4907)) or (layer1_outputs(4797));
    layer2_outputs(3518) <= (layer1_outputs(4134)) and (layer1_outputs(4200));
    layer2_outputs(3519) <= not(layer1_outputs(575));
    layer2_outputs(3520) <= not((layer1_outputs(2848)) xor (layer1_outputs(1220)));
    layer2_outputs(3521) <= not((layer1_outputs(3519)) and (layer1_outputs(1223)));
    layer2_outputs(3522) <= layer1_outputs(482);
    layer2_outputs(3523) <= not((layer1_outputs(215)) xor (layer1_outputs(2525)));
    layer2_outputs(3524) <= not((layer1_outputs(685)) or (layer1_outputs(5068)));
    layer2_outputs(3525) <= (layer1_outputs(3545)) or (layer1_outputs(3969));
    layer2_outputs(3526) <= layer1_outputs(1673);
    layer2_outputs(3527) <= (layer1_outputs(4538)) and not (layer1_outputs(3817));
    layer2_outputs(3528) <= layer1_outputs(2489);
    layer2_outputs(3529) <= not(layer1_outputs(2168));
    layer2_outputs(3530) <= (layer1_outputs(2623)) and not (layer1_outputs(4662));
    layer2_outputs(3531) <= not(layer1_outputs(4696));
    layer2_outputs(3532) <= (layer1_outputs(900)) or (layer1_outputs(3714));
    layer2_outputs(3533) <= (layer1_outputs(1161)) xor (layer1_outputs(652));
    layer2_outputs(3534) <= (layer1_outputs(4500)) xor (layer1_outputs(2487));
    layer2_outputs(3535) <= not(layer1_outputs(1381));
    layer2_outputs(3536) <= '1';
    layer2_outputs(3537) <= (layer1_outputs(2479)) xor (layer1_outputs(1588));
    layer2_outputs(3538) <= not(layer1_outputs(5113));
    layer2_outputs(3539) <= (layer1_outputs(2575)) and not (layer1_outputs(1));
    layer2_outputs(3540) <= layer1_outputs(1175);
    layer2_outputs(3541) <= not(layer1_outputs(2648));
    layer2_outputs(3542) <= not(layer1_outputs(2966)) or (layer1_outputs(1589));
    layer2_outputs(3543) <= not(layer1_outputs(4803));
    layer2_outputs(3544) <= not(layer1_outputs(4478)) or (layer1_outputs(4510));
    layer2_outputs(3545) <= not(layer1_outputs(579));
    layer2_outputs(3546) <= layer1_outputs(4721);
    layer2_outputs(3547) <= (layer1_outputs(4438)) or (layer1_outputs(4804));
    layer2_outputs(3548) <= layer1_outputs(4012);
    layer2_outputs(3549) <= layer1_outputs(2588);
    layer2_outputs(3550) <= (layer1_outputs(2782)) and not (layer1_outputs(2600));
    layer2_outputs(3551) <= (layer1_outputs(2302)) or (layer1_outputs(3745));
    layer2_outputs(3552) <= not((layer1_outputs(1975)) and (layer1_outputs(4446)));
    layer2_outputs(3553) <= not(layer1_outputs(342));
    layer2_outputs(3554) <= not(layer1_outputs(4221));
    layer2_outputs(3555) <= layer1_outputs(2838);
    layer2_outputs(3556) <= layer1_outputs(2715);
    layer2_outputs(3557) <= layer1_outputs(532);
    layer2_outputs(3558) <= (layer1_outputs(2359)) and not (layer1_outputs(1913));
    layer2_outputs(3559) <= (layer1_outputs(790)) or (layer1_outputs(1536));
    layer2_outputs(3560) <= not(layer1_outputs(4981));
    layer2_outputs(3561) <= (layer1_outputs(3089)) and (layer1_outputs(2725));
    layer2_outputs(3562) <= (layer1_outputs(4266)) and not (layer1_outputs(504));
    layer2_outputs(3563) <= (layer1_outputs(3182)) and (layer1_outputs(257));
    layer2_outputs(3564) <= not(layer1_outputs(3524)) or (layer1_outputs(3580));
    layer2_outputs(3565) <= layer1_outputs(3710);
    layer2_outputs(3566) <= not(layer1_outputs(140)) or (layer1_outputs(3514));
    layer2_outputs(3567) <= not(layer1_outputs(4739));
    layer2_outputs(3568) <= layer1_outputs(4726);
    layer2_outputs(3569) <= layer1_outputs(1744);
    layer2_outputs(3570) <= layer1_outputs(924);
    layer2_outputs(3571) <= (layer1_outputs(3171)) xor (layer1_outputs(3593));
    layer2_outputs(3572) <= not(layer1_outputs(150));
    layer2_outputs(3573) <= not(layer1_outputs(17)) or (layer1_outputs(2012));
    layer2_outputs(3574) <= not(layer1_outputs(4042));
    layer2_outputs(3575) <= not(layer1_outputs(693));
    layer2_outputs(3576) <= (layer1_outputs(2049)) or (layer1_outputs(4692));
    layer2_outputs(3577) <= not((layer1_outputs(461)) xor (layer1_outputs(4442)));
    layer2_outputs(3578) <= (layer1_outputs(4779)) and not (layer1_outputs(1492));
    layer2_outputs(3579) <= not(layer1_outputs(3239)) or (layer1_outputs(749));
    layer2_outputs(3580) <= (layer1_outputs(1108)) and not (layer1_outputs(1623));
    layer2_outputs(3581) <= (layer1_outputs(2527)) or (layer1_outputs(2829));
    layer2_outputs(3582) <= not((layer1_outputs(4414)) xor (layer1_outputs(1199)));
    layer2_outputs(3583) <= layer1_outputs(1936);
    layer2_outputs(3584) <= not(layer1_outputs(4536)) or (layer1_outputs(1974));
    layer2_outputs(3585) <= layer1_outputs(1375);
    layer2_outputs(3586) <= (layer1_outputs(4112)) and (layer1_outputs(3771));
    layer2_outputs(3587) <= (layer1_outputs(4377)) and not (layer1_outputs(1104));
    layer2_outputs(3588) <= layer1_outputs(363);
    layer2_outputs(3589) <= (layer1_outputs(536)) and not (layer1_outputs(1706));
    layer2_outputs(3590) <= '0';
    layer2_outputs(3591) <= not((layer1_outputs(1040)) and (layer1_outputs(2429)));
    layer2_outputs(3592) <= layer1_outputs(1079);
    layer2_outputs(3593) <= (layer1_outputs(1745)) xor (layer1_outputs(1351));
    layer2_outputs(3594) <= layer1_outputs(3348);
    layer2_outputs(3595) <= not((layer1_outputs(2367)) or (layer1_outputs(488)));
    layer2_outputs(3596) <= layer1_outputs(529);
    layer2_outputs(3597) <= layer1_outputs(262);
    layer2_outputs(3598) <= (layer1_outputs(2138)) and (layer1_outputs(1564));
    layer2_outputs(3599) <= layer1_outputs(5105);
    layer2_outputs(3600) <= not((layer1_outputs(3404)) xor (layer1_outputs(2963)));
    layer2_outputs(3601) <= (layer1_outputs(2058)) and not (layer1_outputs(701));
    layer2_outputs(3602) <= not((layer1_outputs(1346)) and (layer1_outputs(3825)));
    layer2_outputs(3603) <= '0';
    layer2_outputs(3604) <= not((layer1_outputs(2470)) xor (layer1_outputs(1687)));
    layer2_outputs(3605) <= not(layer1_outputs(2607));
    layer2_outputs(3606) <= not(layer1_outputs(4749));
    layer2_outputs(3607) <= (layer1_outputs(3336)) and not (layer1_outputs(150));
    layer2_outputs(3608) <= layer1_outputs(1720);
    layer2_outputs(3609) <= layer1_outputs(4802);
    layer2_outputs(3610) <= '0';
    layer2_outputs(3611) <= not(layer1_outputs(3691));
    layer2_outputs(3612) <= layer1_outputs(3156);
    layer2_outputs(3613) <= (layer1_outputs(5058)) and (layer1_outputs(1907));
    layer2_outputs(3614) <= not((layer1_outputs(4034)) xor (layer1_outputs(4772)));
    layer2_outputs(3615) <= layer1_outputs(1684);
    layer2_outputs(3616) <= not(layer1_outputs(4228));
    layer2_outputs(3617) <= not(layer1_outputs(2508)) or (layer1_outputs(2148));
    layer2_outputs(3618) <= not(layer1_outputs(1382)) or (layer1_outputs(260));
    layer2_outputs(3619) <= layer1_outputs(3973);
    layer2_outputs(3620) <= not(layer1_outputs(340));
    layer2_outputs(3621) <= not(layer1_outputs(3490));
    layer2_outputs(3622) <= layer1_outputs(1495);
    layer2_outputs(3623) <= (layer1_outputs(4888)) and (layer1_outputs(86));
    layer2_outputs(3624) <= not((layer1_outputs(1842)) or (layer1_outputs(747)));
    layer2_outputs(3625) <= (layer1_outputs(2481)) and not (layer1_outputs(506));
    layer2_outputs(3626) <= layer1_outputs(4408);
    layer2_outputs(3627) <= not(layer1_outputs(2497));
    layer2_outputs(3628) <= (layer1_outputs(3566)) and (layer1_outputs(2457));
    layer2_outputs(3629) <= layer1_outputs(4354);
    layer2_outputs(3630) <= layer1_outputs(946);
    layer2_outputs(3631) <= not((layer1_outputs(2660)) xor (layer1_outputs(2441)));
    layer2_outputs(3632) <= not(layer1_outputs(4156));
    layer2_outputs(3633) <= layer1_outputs(1174);
    layer2_outputs(3634) <= (layer1_outputs(3588)) and not (layer1_outputs(1462));
    layer2_outputs(3635) <= not((layer1_outputs(2812)) and (layer1_outputs(2634)));
    layer2_outputs(3636) <= not(layer1_outputs(2964));
    layer2_outputs(3637) <= not(layer1_outputs(3384)) or (layer1_outputs(4146));
    layer2_outputs(3638) <= layer1_outputs(1180);
    layer2_outputs(3639) <= not((layer1_outputs(157)) or (layer1_outputs(3638)));
    layer2_outputs(3640) <= not((layer1_outputs(4982)) and (layer1_outputs(1147)));
    layer2_outputs(3641) <= (layer1_outputs(4486)) and not (layer1_outputs(4577));
    layer2_outputs(3642) <= not(layer1_outputs(3992));
    layer2_outputs(3643) <= not(layer1_outputs(200));
    layer2_outputs(3644) <= not(layer1_outputs(2433));
    layer2_outputs(3645) <= not(layer1_outputs(4814));
    layer2_outputs(3646) <= not(layer1_outputs(514)) or (layer1_outputs(4433));
    layer2_outputs(3647) <= layer1_outputs(3174);
    layer2_outputs(3648) <= layer1_outputs(4359);
    layer2_outputs(3649) <= not(layer1_outputs(1959));
    layer2_outputs(3650) <= not((layer1_outputs(1657)) xor (layer1_outputs(3878)));
    layer2_outputs(3651) <= (layer1_outputs(824)) and (layer1_outputs(2010));
    layer2_outputs(3652) <= layer1_outputs(5070);
    layer2_outputs(3653) <= not(layer1_outputs(4954));
    layer2_outputs(3654) <= layer1_outputs(1707);
    layer2_outputs(3655) <= layer1_outputs(3226);
    layer2_outputs(3656) <= not(layer1_outputs(1011)) or (layer1_outputs(1688));
    layer2_outputs(3657) <= not((layer1_outputs(3668)) xor (layer1_outputs(2672)));
    layer2_outputs(3658) <= layer1_outputs(4835);
    layer2_outputs(3659) <= not((layer1_outputs(1772)) or (layer1_outputs(1668)));
    layer2_outputs(3660) <= (layer1_outputs(3702)) and not (layer1_outputs(5008));
    layer2_outputs(3661) <= (layer1_outputs(3228)) and not (layer1_outputs(1216));
    layer2_outputs(3662) <= (layer1_outputs(3816)) or (layer1_outputs(1273));
    layer2_outputs(3663) <= not(layer1_outputs(1908)) or (layer1_outputs(129));
    layer2_outputs(3664) <= layer1_outputs(2103);
    layer2_outputs(3665) <= layer1_outputs(5061);
    layer2_outputs(3666) <= not(layer1_outputs(3153));
    layer2_outputs(3667) <= layer1_outputs(4009);
    layer2_outputs(3668) <= not(layer1_outputs(5043)) or (layer1_outputs(1923));
    layer2_outputs(3669) <= not((layer1_outputs(2273)) or (layer1_outputs(491)));
    layer2_outputs(3670) <= layer1_outputs(1045);
    layer2_outputs(3671) <= layer1_outputs(926);
    layer2_outputs(3672) <= not(layer1_outputs(666)) or (layer1_outputs(774));
    layer2_outputs(3673) <= not(layer1_outputs(986)) or (layer1_outputs(1358));
    layer2_outputs(3674) <= (layer1_outputs(70)) xor (layer1_outputs(2207));
    layer2_outputs(3675) <= not(layer1_outputs(3491));
    layer2_outputs(3676) <= (layer1_outputs(222)) and not (layer1_outputs(376));
    layer2_outputs(3677) <= (layer1_outputs(454)) and not (layer1_outputs(2763));
    layer2_outputs(3678) <= layer1_outputs(3950);
    layer2_outputs(3679) <= '1';
    layer2_outputs(3680) <= (layer1_outputs(3824)) xor (layer1_outputs(2647));
    layer2_outputs(3681) <= not(layer1_outputs(2208));
    layer2_outputs(3682) <= layer1_outputs(2083);
    layer2_outputs(3683) <= '0';
    layer2_outputs(3684) <= not((layer1_outputs(1647)) xor (layer1_outputs(1890)));
    layer2_outputs(3685) <= not((layer1_outputs(4571)) or (layer1_outputs(643)));
    layer2_outputs(3686) <= not(layer1_outputs(3985));
    layer2_outputs(3687) <= not((layer1_outputs(1212)) or (layer1_outputs(2240)));
    layer2_outputs(3688) <= not(layer1_outputs(1379));
    layer2_outputs(3689) <= not(layer1_outputs(1090)) or (layer1_outputs(1104));
    layer2_outputs(3690) <= not(layer1_outputs(3159)) or (layer1_outputs(2394));
    layer2_outputs(3691) <= not(layer1_outputs(5075)) or (layer1_outputs(3672));
    layer2_outputs(3692) <= layer1_outputs(2975);
    layer2_outputs(3693) <= not(layer1_outputs(419));
    layer2_outputs(3694) <= not((layer1_outputs(1940)) xor (layer1_outputs(827)));
    layer2_outputs(3695) <= layer1_outputs(2590);
    layer2_outputs(3696) <= layer1_outputs(1718);
    layer2_outputs(3697) <= layer1_outputs(1677);
    layer2_outputs(3698) <= not((layer1_outputs(4493)) and (layer1_outputs(5066)));
    layer2_outputs(3699) <= not((layer1_outputs(3855)) or (layer1_outputs(4087)));
    layer2_outputs(3700) <= (layer1_outputs(1660)) and not (layer1_outputs(4100));
    layer2_outputs(3701) <= '1';
    layer2_outputs(3702) <= (layer1_outputs(457)) and not (layer1_outputs(4361));
    layer2_outputs(3703) <= layer1_outputs(4327);
    layer2_outputs(3704) <= not(layer1_outputs(1776));
    layer2_outputs(3705) <= not(layer1_outputs(3413));
    layer2_outputs(3706) <= not((layer1_outputs(5026)) or (layer1_outputs(3982)));
    layer2_outputs(3707) <= layer1_outputs(4155);
    layer2_outputs(3708) <= not(layer1_outputs(28));
    layer2_outputs(3709) <= not(layer1_outputs(5015));
    layer2_outputs(3710) <= layer1_outputs(4744);
    layer2_outputs(3711) <= (layer1_outputs(3313)) and not (layer1_outputs(3652));
    layer2_outputs(3712) <= '0';
    layer2_outputs(3713) <= layer1_outputs(2184);
    layer2_outputs(3714) <= not((layer1_outputs(1175)) or (layer1_outputs(2097)));
    layer2_outputs(3715) <= not((layer1_outputs(772)) and (layer1_outputs(2890)));
    layer2_outputs(3716) <= not(layer1_outputs(2102)) or (layer1_outputs(830));
    layer2_outputs(3717) <= (layer1_outputs(768)) or (layer1_outputs(3588));
    layer2_outputs(3718) <= not((layer1_outputs(263)) xor (layer1_outputs(1514)));
    layer2_outputs(3719) <= not(layer1_outputs(75));
    layer2_outputs(3720) <= (layer1_outputs(1564)) and not (layer1_outputs(1829));
    layer2_outputs(3721) <= not(layer1_outputs(4092));
    layer2_outputs(3722) <= (layer1_outputs(3331)) or (layer1_outputs(1861));
    layer2_outputs(3723) <= (layer1_outputs(2378)) and (layer1_outputs(1018));
    layer2_outputs(3724) <= not(layer1_outputs(4027));
    layer2_outputs(3725) <= layer1_outputs(323);
    layer2_outputs(3726) <= not(layer1_outputs(1198)) or (layer1_outputs(4305));
    layer2_outputs(3727) <= not(layer1_outputs(3549));
    layer2_outputs(3728) <= not(layer1_outputs(1364)) or (layer1_outputs(1671));
    layer2_outputs(3729) <= (layer1_outputs(2862)) and not (layer1_outputs(4424));
    layer2_outputs(3730) <= layer1_outputs(1301);
    layer2_outputs(3731) <= layer1_outputs(718);
    layer2_outputs(3732) <= not(layer1_outputs(3274));
    layer2_outputs(3733) <= '0';
    layer2_outputs(3734) <= not(layer1_outputs(2080));
    layer2_outputs(3735) <= (layer1_outputs(507)) or (layer1_outputs(3225));
    layer2_outputs(3736) <= not(layer1_outputs(831));
    layer2_outputs(3737) <= layer1_outputs(3806);
    layer2_outputs(3738) <= (layer1_outputs(522)) or (layer1_outputs(3999));
    layer2_outputs(3739) <= not(layer1_outputs(601));
    layer2_outputs(3740) <= not(layer1_outputs(3768));
    layer2_outputs(3741) <= (layer1_outputs(3244)) xor (layer1_outputs(2095));
    layer2_outputs(3742) <= layer1_outputs(3498);
    layer2_outputs(3743) <= not(layer1_outputs(3615));
    layer2_outputs(3744) <= layer1_outputs(3572);
    layer2_outputs(3745) <= not(layer1_outputs(4168));
    layer2_outputs(3746) <= not(layer1_outputs(1562));
    layer2_outputs(3747) <= not(layer1_outputs(2921)) or (layer1_outputs(1506));
    layer2_outputs(3748) <= layer1_outputs(556);
    layer2_outputs(3749) <= layer1_outputs(4785);
    layer2_outputs(3750) <= '1';
    layer2_outputs(3751) <= layer1_outputs(2542);
    layer2_outputs(3752) <= not(layer1_outputs(2956));
    layer2_outputs(3753) <= not(layer1_outputs(3478));
    layer2_outputs(3754) <= not((layer1_outputs(1174)) xor (layer1_outputs(5021)));
    layer2_outputs(3755) <= not((layer1_outputs(2097)) or (layer1_outputs(1116)));
    layer2_outputs(3756) <= (layer1_outputs(2408)) and not (layer1_outputs(596));
    layer2_outputs(3757) <= not(layer1_outputs(3409));
    layer2_outputs(3758) <= not(layer1_outputs(2057));
    layer2_outputs(3759) <= layer1_outputs(1154);
    layer2_outputs(3760) <= (layer1_outputs(4329)) xor (layer1_outputs(2053));
    layer2_outputs(3761) <= not(layer1_outputs(2086));
    layer2_outputs(3762) <= not(layer1_outputs(4479));
    layer2_outputs(3763) <= layer1_outputs(1733);
    layer2_outputs(3764) <= (layer1_outputs(564)) xor (layer1_outputs(4610));
    layer2_outputs(3765) <= not((layer1_outputs(4414)) or (layer1_outputs(2173)));
    layer2_outputs(3766) <= not(layer1_outputs(2891));
    layer2_outputs(3767) <= not((layer1_outputs(1209)) or (layer1_outputs(3591)));
    layer2_outputs(3768) <= (layer1_outputs(3711)) and not (layer1_outputs(4911));
    layer2_outputs(3769) <= (layer1_outputs(4286)) and not (layer1_outputs(4539));
    layer2_outputs(3770) <= not((layer1_outputs(4040)) xor (layer1_outputs(1091)));
    layer2_outputs(3771) <= (layer1_outputs(3584)) and (layer1_outputs(546));
    layer2_outputs(3772) <= not(layer1_outputs(995));
    layer2_outputs(3773) <= not(layer1_outputs(3577));
    layer2_outputs(3774) <= not((layer1_outputs(720)) or (layer1_outputs(1685)));
    layer2_outputs(3775) <= not(layer1_outputs(178)) or (layer1_outputs(4783));
    layer2_outputs(3776) <= not(layer1_outputs(4067));
    layer2_outputs(3777) <= not(layer1_outputs(2320)) or (layer1_outputs(3586));
    layer2_outputs(3778) <= not(layer1_outputs(381));
    layer2_outputs(3779) <= (layer1_outputs(4929)) xor (layer1_outputs(2124));
    layer2_outputs(3780) <= (layer1_outputs(762)) or (layer1_outputs(3339));
    layer2_outputs(3781) <= (layer1_outputs(1747)) or (layer1_outputs(1038));
    layer2_outputs(3782) <= not(layer1_outputs(3182));
    layer2_outputs(3783) <= layer1_outputs(782);
    layer2_outputs(3784) <= not((layer1_outputs(2752)) or (layer1_outputs(114)));
    layer2_outputs(3785) <= (layer1_outputs(1817)) and not (layer1_outputs(3370));
    layer2_outputs(3786) <= not(layer1_outputs(3325));
    layer2_outputs(3787) <= not(layer1_outputs(3953)) or (layer1_outputs(4));
    layer2_outputs(3788) <= layer1_outputs(2064);
    layer2_outputs(3789) <= layer1_outputs(1327);
    layer2_outputs(3790) <= not(layer1_outputs(4517)) or (layer1_outputs(2040));
    layer2_outputs(3791) <= (layer1_outputs(4112)) xor (layer1_outputs(4341));
    layer2_outputs(3792) <= not(layer1_outputs(3120));
    layer2_outputs(3793) <= not((layer1_outputs(1991)) xor (layer1_outputs(3562)));
    layer2_outputs(3794) <= not((layer1_outputs(3423)) or (layer1_outputs(4356)));
    layer2_outputs(3795) <= not(layer1_outputs(3595));
    layer2_outputs(3796) <= (layer1_outputs(2387)) xor (layer1_outputs(778));
    layer2_outputs(3797) <= not(layer1_outputs(4106)) or (layer1_outputs(1630));
    layer2_outputs(3798) <= (layer1_outputs(1178)) and not (layer1_outputs(590));
    layer2_outputs(3799) <= '1';
    layer2_outputs(3800) <= layer1_outputs(4817);
    layer2_outputs(3801) <= not((layer1_outputs(912)) or (layer1_outputs(5012)));
    layer2_outputs(3802) <= not(layer1_outputs(4514));
    layer2_outputs(3803) <= (layer1_outputs(1211)) and (layer1_outputs(1146));
    layer2_outputs(3804) <= '0';
    layer2_outputs(3805) <= (layer1_outputs(3284)) or (layer1_outputs(70));
    layer2_outputs(3806) <= not(layer1_outputs(3257));
    layer2_outputs(3807) <= (layer1_outputs(3585)) and (layer1_outputs(278));
    layer2_outputs(3808) <= not(layer1_outputs(5050));
    layer2_outputs(3809) <= not(layer1_outputs(2999));
    layer2_outputs(3810) <= not(layer1_outputs(227));
    layer2_outputs(3811) <= layer1_outputs(755);
    layer2_outputs(3812) <= layer1_outputs(3200);
    layer2_outputs(3813) <= not(layer1_outputs(2688)) or (layer1_outputs(3682));
    layer2_outputs(3814) <= not(layer1_outputs(3399)) or (layer1_outputs(847));
    layer2_outputs(3815) <= not(layer1_outputs(2822));
    layer2_outputs(3816) <= (layer1_outputs(1106)) and (layer1_outputs(2118));
    layer2_outputs(3817) <= (layer1_outputs(4912)) and not (layer1_outputs(718));
    layer2_outputs(3818) <= (layer1_outputs(4631)) xor (layer1_outputs(892));
    layer2_outputs(3819) <= not((layer1_outputs(231)) xor (layer1_outputs(3351)));
    layer2_outputs(3820) <= (layer1_outputs(4808)) xor (layer1_outputs(347));
    layer2_outputs(3821) <= not(layer1_outputs(4384)) or (layer1_outputs(3531));
    layer2_outputs(3822) <= not(layer1_outputs(972));
    layer2_outputs(3823) <= (layer1_outputs(937)) and not (layer1_outputs(2182));
    layer2_outputs(3824) <= '1';
    layer2_outputs(3825) <= layer1_outputs(2407);
    layer2_outputs(3826) <= (layer1_outputs(2558)) xor (layer1_outputs(4520));
    layer2_outputs(3827) <= (layer1_outputs(1008)) and (layer1_outputs(206));
    layer2_outputs(3828) <= not(layer1_outputs(618));
    layer2_outputs(3829) <= layer1_outputs(2967);
    layer2_outputs(3830) <= not((layer1_outputs(1544)) xor (layer1_outputs(3857)));
    layer2_outputs(3831) <= not((layer1_outputs(3664)) xor (layer1_outputs(1217)));
    layer2_outputs(3832) <= not((layer1_outputs(3901)) or (layer1_outputs(1883)));
    layer2_outputs(3833) <= not((layer1_outputs(3021)) xor (layer1_outputs(4699)));
    layer2_outputs(3834) <= not(layer1_outputs(3994));
    layer2_outputs(3835) <= not(layer1_outputs(4215)) or (layer1_outputs(2307));
    layer2_outputs(3836) <= layer1_outputs(3811);
    layer2_outputs(3837) <= not(layer1_outputs(2442));
    layer2_outputs(3838) <= layer1_outputs(2971);
    layer2_outputs(3839) <= not((layer1_outputs(2599)) and (layer1_outputs(4603)));
    layer2_outputs(3840) <= (layer1_outputs(5)) or (layer1_outputs(4701));
    layer2_outputs(3841) <= not((layer1_outputs(4470)) or (layer1_outputs(431)));
    layer2_outputs(3842) <= layer1_outputs(2014);
    layer2_outputs(3843) <= not(layer1_outputs(2190));
    layer2_outputs(3844) <= not((layer1_outputs(3034)) and (layer1_outputs(3675)));
    layer2_outputs(3845) <= not(layer1_outputs(2535));
    layer2_outputs(3846) <= (layer1_outputs(3291)) or (layer1_outputs(4459));
    layer2_outputs(3847) <= not(layer1_outputs(5071));
    layer2_outputs(3848) <= (layer1_outputs(3152)) and (layer1_outputs(2540));
    layer2_outputs(3849) <= (layer1_outputs(3828)) or (layer1_outputs(2987));
    layer2_outputs(3850) <= not((layer1_outputs(1735)) xor (layer1_outputs(2870)));
    layer2_outputs(3851) <= not((layer1_outputs(775)) and (layer1_outputs(2624)));
    layer2_outputs(3852) <= layer1_outputs(139);
    layer2_outputs(3853) <= not(layer1_outputs(3373));
    layer2_outputs(3854) <= not(layer1_outputs(5102));
    layer2_outputs(3855) <= not(layer1_outputs(541)) or (layer1_outputs(2694));
    layer2_outputs(3856) <= layer1_outputs(3317);
    layer2_outputs(3857) <= not((layer1_outputs(528)) xor (layer1_outputs(4493)));
    layer2_outputs(3858) <= not(layer1_outputs(5113));
    layer2_outputs(3859) <= (layer1_outputs(2763)) xor (layer1_outputs(4159));
    layer2_outputs(3860) <= layer1_outputs(127);
    layer2_outputs(3861) <= not(layer1_outputs(287));
    layer2_outputs(3862) <= not(layer1_outputs(4660));
    layer2_outputs(3863) <= not((layer1_outputs(4125)) xor (layer1_outputs(5062)));
    layer2_outputs(3864) <= not((layer1_outputs(3440)) xor (layer1_outputs(4327)));
    layer2_outputs(3865) <= not((layer1_outputs(1248)) and (layer1_outputs(2185)));
    layer2_outputs(3866) <= layer1_outputs(1598);
    layer2_outputs(3867) <= not(layer1_outputs(1459)) or (layer1_outputs(4856));
    layer2_outputs(3868) <= not(layer1_outputs(4216));
    layer2_outputs(3869) <= (layer1_outputs(1028)) and not (layer1_outputs(246));
    layer2_outputs(3870) <= not(layer1_outputs(1010));
    layer2_outputs(3871) <= not(layer1_outputs(1194)) or (layer1_outputs(2368));
    layer2_outputs(3872) <= not((layer1_outputs(1166)) and (layer1_outputs(3077)));
    layer2_outputs(3873) <= not(layer1_outputs(2717));
    layer2_outputs(3874) <= (layer1_outputs(1176)) or (layer1_outputs(100));
    layer2_outputs(3875) <= '1';
    layer2_outputs(3876) <= layer1_outputs(732);
    layer2_outputs(3877) <= (layer1_outputs(440)) or (layer1_outputs(135));
    layer2_outputs(3878) <= not((layer1_outputs(3401)) xor (layer1_outputs(3552)));
    layer2_outputs(3879) <= not(layer1_outputs(1007));
    layer2_outputs(3880) <= not((layer1_outputs(2695)) and (layer1_outputs(1779)));
    layer2_outputs(3881) <= layer1_outputs(4362);
    layer2_outputs(3882) <= (layer1_outputs(4053)) xor (layer1_outputs(1787));
    layer2_outputs(3883) <= layer1_outputs(4257);
    layer2_outputs(3884) <= (layer1_outputs(4886)) xor (layer1_outputs(4703));
    layer2_outputs(3885) <= not((layer1_outputs(3836)) xor (layer1_outputs(4756)));
    layer2_outputs(3886) <= not(layer1_outputs(3255));
    layer2_outputs(3887) <= layer1_outputs(2417);
    layer2_outputs(3888) <= not(layer1_outputs(3936)) or (layer1_outputs(4269));
    layer2_outputs(3889) <= not(layer1_outputs(389)) or (layer1_outputs(3078));
    layer2_outputs(3890) <= layer1_outputs(3434);
    layer2_outputs(3891) <= layer1_outputs(5078);
    layer2_outputs(3892) <= layer1_outputs(1814);
    layer2_outputs(3893) <= layer1_outputs(4818);
    layer2_outputs(3894) <= layer1_outputs(2361);
    layer2_outputs(3895) <= layer1_outputs(3942);
    layer2_outputs(3896) <= not(layer1_outputs(2099));
    layer2_outputs(3897) <= not(layer1_outputs(635)) or (layer1_outputs(2205));
    layer2_outputs(3898) <= (layer1_outputs(4247)) and not (layer1_outputs(2843));
    layer2_outputs(3899) <= layer1_outputs(3139);
    layer2_outputs(3900) <= layer1_outputs(3657);
    layer2_outputs(3901) <= not(layer1_outputs(4845)) or (layer1_outputs(3694));
    layer2_outputs(3902) <= not(layer1_outputs(4970));
    layer2_outputs(3903) <= (layer1_outputs(3186)) xor (layer1_outputs(2313));
    layer2_outputs(3904) <= layer1_outputs(274);
    layer2_outputs(3905) <= not(layer1_outputs(2999));
    layer2_outputs(3906) <= (layer1_outputs(371)) and not (layer1_outputs(1145));
    layer2_outputs(3907) <= not(layer1_outputs(401));
    layer2_outputs(3908) <= not(layer1_outputs(4395));
    layer2_outputs(3909) <= (layer1_outputs(626)) and not (layer1_outputs(1092));
    layer2_outputs(3910) <= not((layer1_outputs(361)) xor (layer1_outputs(2380)));
    layer2_outputs(3911) <= (layer1_outputs(1399)) and not (layer1_outputs(1989));
    layer2_outputs(3912) <= not((layer1_outputs(2309)) and (layer1_outputs(818)));
    layer2_outputs(3913) <= '0';
    layer2_outputs(3914) <= (layer1_outputs(910)) and (layer1_outputs(2503));
    layer2_outputs(3915) <= layer1_outputs(5109);
    layer2_outputs(3916) <= (layer1_outputs(39)) and (layer1_outputs(987));
    layer2_outputs(3917) <= not(layer1_outputs(4358));
    layer2_outputs(3918) <= layer1_outputs(1943);
    layer2_outputs(3919) <= not(layer1_outputs(5005));
    layer2_outputs(3920) <= not((layer1_outputs(3877)) xor (layer1_outputs(289)));
    layer2_outputs(3921) <= not(layer1_outputs(4829));
    layer2_outputs(3922) <= (layer1_outputs(2061)) and not (layer1_outputs(2304));
    layer2_outputs(3923) <= layer1_outputs(2625);
    layer2_outputs(3924) <= not(layer1_outputs(3515)) or (layer1_outputs(3546));
    layer2_outputs(3925) <= not((layer1_outputs(106)) and (layer1_outputs(3087)));
    layer2_outputs(3926) <= (layer1_outputs(2911)) and not (layer1_outputs(1047));
    layer2_outputs(3927) <= not(layer1_outputs(558));
    layer2_outputs(3928) <= not(layer1_outputs(3163)) or (layer1_outputs(2060));
    layer2_outputs(3929) <= not(layer1_outputs(2769)) or (layer1_outputs(2514));
    layer2_outputs(3930) <= (layer1_outputs(2798)) and not (layer1_outputs(3898));
    layer2_outputs(3931) <= (layer1_outputs(2264)) and not (layer1_outputs(619));
    layer2_outputs(3932) <= (layer1_outputs(517)) xor (layer1_outputs(4271));
    layer2_outputs(3933) <= (layer1_outputs(1504)) xor (layer1_outputs(3262));
    layer2_outputs(3934) <= not(layer1_outputs(2125)) or (layer1_outputs(2132));
    layer2_outputs(3935) <= not(layer1_outputs(4168));
    layer2_outputs(3936) <= not((layer1_outputs(575)) xor (layer1_outputs(4487)));
    layer2_outputs(3937) <= not(layer1_outputs(822));
    layer2_outputs(3938) <= '1';
    layer2_outputs(3939) <= not(layer1_outputs(4676));
    layer2_outputs(3940) <= not(layer1_outputs(4480));
    layer2_outputs(3941) <= not(layer1_outputs(1079));
    layer2_outputs(3942) <= (layer1_outputs(341)) xor (layer1_outputs(4865));
    layer2_outputs(3943) <= (layer1_outputs(4177)) xor (layer1_outputs(3078));
    layer2_outputs(3944) <= '0';
    layer2_outputs(3945) <= layer1_outputs(3864);
    layer2_outputs(3946) <= not(layer1_outputs(3178)) or (layer1_outputs(4616));
    layer2_outputs(3947) <= not(layer1_outputs(4248));
    layer2_outputs(3948) <= not((layer1_outputs(2514)) and (layer1_outputs(2880)));
    layer2_outputs(3949) <= not(layer1_outputs(3828));
    layer2_outputs(3950) <= not(layer1_outputs(3301));
    layer2_outputs(3951) <= not(layer1_outputs(919));
    layer2_outputs(3952) <= not(layer1_outputs(2483));
    layer2_outputs(3953) <= layer1_outputs(2413);
    layer2_outputs(3954) <= not(layer1_outputs(1003)) or (layer1_outputs(1969));
    layer2_outputs(3955) <= not(layer1_outputs(4225)) or (layer1_outputs(432));
    layer2_outputs(3956) <= layer1_outputs(3285);
    layer2_outputs(3957) <= not(layer1_outputs(1451));
    layer2_outputs(3958) <= not(layer1_outputs(4153));
    layer2_outputs(3959) <= not(layer1_outputs(2778));
    layer2_outputs(3960) <= (layer1_outputs(3014)) and (layer1_outputs(374));
    layer2_outputs(3961) <= (layer1_outputs(3694)) or (layer1_outputs(4374));
    layer2_outputs(3962) <= layer1_outputs(4333);
    layer2_outputs(3963) <= (layer1_outputs(4329)) and not (layer1_outputs(345));
    layer2_outputs(3964) <= not(layer1_outputs(2968));
    layer2_outputs(3965) <= not(layer1_outputs(4925)) or (layer1_outputs(4387));
    layer2_outputs(3966) <= layer1_outputs(2338);
    layer2_outputs(3967) <= not(layer1_outputs(3981)) or (layer1_outputs(232));
    layer2_outputs(3968) <= not((layer1_outputs(523)) or (layer1_outputs(1533)));
    layer2_outputs(3969) <= not((layer1_outputs(1734)) and (layer1_outputs(3749)));
    layer2_outputs(3970) <= not(layer1_outputs(602));
    layer2_outputs(3971) <= not(layer1_outputs(2803));
    layer2_outputs(3972) <= layer1_outputs(3161);
    layer2_outputs(3973) <= (layer1_outputs(2339)) and not (layer1_outputs(3787));
    layer2_outputs(3974) <= layer1_outputs(555);
    layer2_outputs(3975) <= layer1_outputs(2847);
    layer2_outputs(3976) <= (layer1_outputs(1686)) and (layer1_outputs(1610));
    layer2_outputs(3977) <= not(layer1_outputs(3485));
    layer2_outputs(3978) <= not((layer1_outputs(916)) or (layer1_outputs(3020)));
    layer2_outputs(3979) <= layer1_outputs(846);
    layer2_outputs(3980) <= not(layer1_outputs(3353));
    layer2_outputs(3981) <= (layer1_outputs(944)) or (layer1_outputs(1897));
    layer2_outputs(3982) <= (layer1_outputs(3557)) and (layer1_outputs(2852));
    layer2_outputs(3983) <= layer1_outputs(2384);
    layer2_outputs(3984) <= not(layer1_outputs(1468));
    layer2_outputs(3985) <= not((layer1_outputs(2866)) xor (layer1_outputs(1328)));
    layer2_outputs(3986) <= not(layer1_outputs(3739));
    layer2_outputs(3987) <= layer1_outputs(4672);
    layer2_outputs(3988) <= layer1_outputs(1590);
    layer2_outputs(3989) <= (layer1_outputs(510)) xor (layer1_outputs(3050));
    layer2_outputs(3990) <= not(layer1_outputs(398));
    layer2_outputs(3991) <= not((layer1_outputs(3137)) or (layer1_outputs(729)));
    layer2_outputs(3992) <= not(layer1_outputs(1556));
    layer2_outputs(3993) <= (layer1_outputs(4823)) or (layer1_outputs(4979));
    layer2_outputs(3994) <= (layer1_outputs(958)) and (layer1_outputs(614));
    layer2_outputs(3995) <= (layer1_outputs(2845)) and not (layer1_outputs(2032));
    layer2_outputs(3996) <= not(layer1_outputs(964));
    layer2_outputs(3997) <= not(layer1_outputs(548)) or (layer1_outputs(8));
    layer2_outputs(3998) <= (layer1_outputs(638)) and (layer1_outputs(3324));
    layer2_outputs(3999) <= not(layer1_outputs(914));
    layer2_outputs(4000) <= not((layer1_outputs(3980)) or (layer1_outputs(2571)));
    layer2_outputs(4001) <= not(layer1_outputs(706));
    layer2_outputs(4002) <= not(layer1_outputs(1106));
    layer2_outputs(4003) <= not(layer1_outputs(2327));
    layer2_outputs(4004) <= (layer1_outputs(1858)) and not (layer1_outputs(4017));
    layer2_outputs(4005) <= layer1_outputs(770);
    layer2_outputs(4006) <= (layer1_outputs(4013)) and (layer1_outputs(955));
    layer2_outputs(4007) <= not(layer1_outputs(449));
    layer2_outputs(4008) <= not(layer1_outputs(3114));
    layer2_outputs(4009) <= not((layer1_outputs(1364)) xor (layer1_outputs(3434)));
    layer2_outputs(4010) <= not(layer1_outputs(2589));
    layer2_outputs(4011) <= not(layer1_outputs(3695));
    layer2_outputs(4012) <= not(layer1_outputs(3848));
    layer2_outputs(4013) <= layer1_outputs(457);
    layer2_outputs(4014) <= not(layer1_outputs(517)) or (layer1_outputs(2764));
    layer2_outputs(4015) <= not((layer1_outputs(2881)) or (layer1_outputs(1235)));
    layer2_outputs(4016) <= layer1_outputs(3968);
    layer2_outputs(4017) <= (layer1_outputs(1132)) xor (layer1_outputs(1665));
    layer2_outputs(4018) <= not(layer1_outputs(3228));
    layer2_outputs(4019) <= (layer1_outputs(1761)) and not (layer1_outputs(2504));
    layer2_outputs(4020) <= (layer1_outputs(258)) xor (layer1_outputs(2179));
    layer2_outputs(4021) <= layer1_outputs(1448);
    layer2_outputs(4022) <= not(layer1_outputs(3839));
    layer2_outputs(4023) <= not(layer1_outputs(1347));
    layer2_outputs(4024) <= not(layer1_outputs(1760));
    layer2_outputs(4025) <= not(layer1_outputs(426));
    layer2_outputs(4026) <= layer1_outputs(4527);
    layer2_outputs(4027) <= layer1_outputs(3904);
    layer2_outputs(4028) <= not(layer1_outputs(3910));
    layer2_outputs(4029) <= layer1_outputs(3938);
    layer2_outputs(4030) <= not(layer1_outputs(680)) or (layer1_outputs(304));
    layer2_outputs(4031) <= not(layer1_outputs(5030));
    layer2_outputs(4032) <= not(layer1_outputs(4207));
    layer2_outputs(4033) <= '1';
    layer2_outputs(4034) <= not(layer1_outputs(2870));
    layer2_outputs(4035) <= (layer1_outputs(3495)) and (layer1_outputs(2676));
    layer2_outputs(4036) <= layer1_outputs(1594);
    layer2_outputs(4037) <= layer1_outputs(3201);
    layer2_outputs(4038) <= (layer1_outputs(4381)) xor (layer1_outputs(3961));
    layer2_outputs(4039) <= not((layer1_outputs(5097)) or (layer1_outputs(4060)));
    layer2_outputs(4040) <= not((layer1_outputs(4871)) xor (layer1_outputs(1243)));
    layer2_outputs(4041) <= layer1_outputs(2719);
    layer2_outputs(4042) <= layer1_outputs(2394);
    layer2_outputs(4043) <= not((layer1_outputs(2)) xor (layer1_outputs(140)));
    layer2_outputs(4044) <= not(layer1_outputs(2448));
    layer2_outputs(4045) <= not(layer1_outputs(4998));
    layer2_outputs(4046) <= (layer1_outputs(3028)) or (layer1_outputs(1651));
    layer2_outputs(4047) <= (layer1_outputs(2139)) or (layer1_outputs(4437));
    layer2_outputs(4048) <= not((layer1_outputs(3430)) and (layer1_outputs(2864)));
    layer2_outputs(4049) <= not(layer1_outputs(4724));
    layer2_outputs(4050) <= not(layer1_outputs(1870)) or (layer1_outputs(2656));
    layer2_outputs(4051) <= not(layer1_outputs(2472));
    layer2_outputs(4052) <= not(layer1_outputs(1059));
    layer2_outputs(4053) <= (layer1_outputs(4958)) and not (layer1_outputs(4935));
    layer2_outputs(4054) <= layer1_outputs(559);
    layer2_outputs(4055) <= (layer1_outputs(4866)) and not (layer1_outputs(2287));
    layer2_outputs(4056) <= not(layer1_outputs(4090)) or (layer1_outputs(325));
    layer2_outputs(4057) <= not(layer1_outputs(3445)) or (layer1_outputs(751));
    layer2_outputs(4058) <= layer1_outputs(984);
    layer2_outputs(4059) <= layer1_outputs(2451);
    layer2_outputs(4060) <= not(layer1_outputs(1611)) or (layer1_outputs(3337));
    layer2_outputs(4061) <= not((layer1_outputs(4227)) xor (layer1_outputs(3838)));
    layer2_outputs(4062) <= not((layer1_outputs(459)) xor (layer1_outputs(3836)));
    layer2_outputs(4063) <= (layer1_outputs(4450)) and not (layer1_outputs(3593));
    layer2_outputs(4064) <= (layer1_outputs(380)) and not (layer1_outputs(3616));
    layer2_outputs(4065) <= not((layer1_outputs(1913)) xor (layer1_outputs(4872)));
    layer2_outputs(4066) <= layer1_outputs(2709);
    layer2_outputs(4067) <= not(layer1_outputs(4374));
    layer2_outputs(4068) <= (layer1_outputs(2853)) and not (layer1_outputs(3980));
    layer2_outputs(4069) <= not(layer1_outputs(413));
    layer2_outputs(4070) <= layer1_outputs(1656);
    layer2_outputs(4071) <= (layer1_outputs(3335)) and (layer1_outputs(4129));
    layer2_outputs(4072) <= not((layer1_outputs(4860)) xor (layer1_outputs(4824)));
    layer2_outputs(4073) <= (layer1_outputs(3118)) and (layer1_outputs(609));
    layer2_outputs(4074) <= not(layer1_outputs(2296));
    layer2_outputs(4075) <= layer1_outputs(2892);
    layer2_outputs(4076) <= layer1_outputs(904);
    layer2_outputs(4077) <= (layer1_outputs(877)) and not (layer1_outputs(2612));
    layer2_outputs(4078) <= not((layer1_outputs(866)) or (layer1_outputs(2296)));
    layer2_outputs(4079) <= not(layer1_outputs(1493)) or (layer1_outputs(1934));
    layer2_outputs(4080) <= not(layer1_outputs(632));
    layer2_outputs(4081) <= (layer1_outputs(2388)) or (layer1_outputs(2318));
    layer2_outputs(4082) <= not((layer1_outputs(2161)) xor (layer1_outputs(2069)));
    layer2_outputs(4083) <= not((layer1_outputs(2608)) and (layer1_outputs(2855)));
    layer2_outputs(4084) <= '1';
    layer2_outputs(4085) <= not(layer1_outputs(4481));
    layer2_outputs(4086) <= not(layer1_outputs(2181)) or (layer1_outputs(1411));
    layer2_outputs(4087) <= layer1_outputs(3016);
    layer2_outputs(4088) <= (layer1_outputs(1403)) and not (layer1_outputs(2425));
    layer2_outputs(4089) <= not(layer1_outputs(2164));
    layer2_outputs(4090) <= layer1_outputs(1446);
    layer2_outputs(4091) <= not(layer1_outputs(1180));
    layer2_outputs(4092) <= layer1_outputs(3156);
    layer2_outputs(4093) <= not(layer1_outputs(2932));
    layer2_outputs(4094) <= (layer1_outputs(685)) or (layer1_outputs(3928));
    layer2_outputs(4095) <= not(layer1_outputs(3717)) or (layer1_outputs(1056));
    layer2_outputs(4096) <= (layer1_outputs(3375)) and (layer1_outputs(4843));
    layer2_outputs(4097) <= (layer1_outputs(4054)) xor (layer1_outputs(2453));
    layer2_outputs(4098) <= layer1_outputs(35);
    layer2_outputs(4099) <= (layer1_outputs(1852)) and (layer1_outputs(490));
    layer2_outputs(4100) <= not(layer1_outputs(4985)) or (layer1_outputs(4464));
    layer2_outputs(4101) <= not(layer1_outputs(1592));
    layer2_outputs(4102) <= not((layer1_outputs(107)) xor (layer1_outputs(1218)));
    layer2_outputs(4103) <= not(layer1_outputs(1790));
    layer2_outputs(4104) <= layer1_outputs(305);
    layer2_outputs(4105) <= layer1_outputs(2929);
    layer2_outputs(4106) <= layer1_outputs(4620);
    layer2_outputs(4107) <= (layer1_outputs(2488)) xor (layer1_outputs(1547));
    layer2_outputs(4108) <= layer1_outputs(4427);
    layer2_outputs(4109) <= not((layer1_outputs(503)) and (layer1_outputs(1799)));
    layer2_outputs(4110) <= layer1_outputs(3117);
    layer2_outputs(4111) <= not(layer1_outputs(979));
    layer2_outputs(4112) <= (layer1_outputs(4102)) or (layer1_outputs(2067));
    layer2_outputs(4113) <= layer1_outputs(1184);
    layer2_outputs(4114) <= not(layer1_outputs(760));
    layer2_outputs(4115) <= not(layer1_outputs(3846));
    layer2_outputs(4116) <= not(layer1_outputs(3348));
    layer2_outputs(4117) <= layer1_outputs(159);
    layer2_outputs(4118) <= '0';
    layer2_outputs(4119) <= layer1_outputs(4380);
    layer2_outputs(4120) <= (layer1_outputs(1806)) xor (layer1_outputs(1381));
    layer2_outputs(4121) <= not(layer1_outputs(3830));
    layer2_outputs(4122) <= layer1_outputs(2466);
    layer2_outputs(4123) <= (layer1_outputs(448)) and not (layer1_outputs(1479));
    layer2_outputs(4124) <= not(layer1_outputs(4421));
    layer2_outputs(4125) <= not(layer1_outputs(1263));
    layer2_outputs(4126) <= not(layer1_outputs(1116));
    layer2_outputs(4127) <= layer1_outputs(1886);
    layer2_outputs(4128) <= not(layer1_outputs(869));
    layer2_outputs(4129) <= not(layer1_outputs(1909));
    layer2_outputs(4130) <= not(layer1_outputs(2157)) or (layer1_outputs(2779));
    layer2_outputs(4131) <= not((layer1_outputs(154)) xor (layer1_outputs(2834)));
    layer2_outputs(4132) <= not((layer1_outputs(2790)) or (layer1_outputs(88)));
    layer2_outputs(4133) <= (layer1_outputs(2104)) or (layer1_outputs(1765));
    layer2_outputs(4134) <= (layer1_outputs(2342)) and not (layer1_outputs(3396));
    layer2_outputs(4135) <= layer1_outputs(4951);
    layer2_outputs(4136) <= not((layer1_outputs(4589)) xor (layer1_outputs(4697)));
    layer2_outputs(4137) <= not((layer1_outputs(2159)) or (layer1_outputs(639)));
    layer2_outputs(4138) <= (layer1_outputs(1965)) and not (layer1_outputs(1412));
    layer2_outputs(4139) <= not(layer1_outputs(5047)) or (layer1_outputs(2313));
    layer2_outputs(4140) <= (layer1_outputs(1669)) or (layer1_outputs(163));
    layer2_outputs(4141) <= (layer1_outputs(4415)) xor (layer1_outputs(3497));
    layer2_outputs(4142) <= (layer1_outputs(1312)) or (layer1_outputs(3972));
    layer2_outputs(4143) <= (layer1_outputs(213)) and not (layer1_outputs(3163));
    layer2_outputs(4144) <= not(layer1_outputs(2412));
    layer2_outputs(4145) <= not(layer1_outputs(4833)) or (layer1_outputs(279));
    layer2_outputs(4146) <= layer1_outputs(4751);
    layer2_outputs(4147) <= (layer1_outputs(4364)) or (layer1_outputs(4579));
    layer2_outputs(4148) <= not(layer1_outputs(347));
    layer2_outputs(4149) <= not((layer1_outputs(1080)) and (layer1_outputs(43)));
    layer2_outputs(4150) <= (layer1_outputs(2087)) and not (layer1_outputs(974));
    layer2_outputs(4151) <= not(layer1_outputs(4867));
    layer2_outputs(4152) <= not((layer1_outputs(41)) and (layer1_outputs(1981)));
    layer2_outputs(4153) <= not(layer1_outputs(1191));
    layer2_outputs(4154) <= not((layer1_outputs(4992)) or (layer1_outputs(3661)));
    layer2_outputs(4155) <= (layer1_outputs(903)) or (layer1_outputs(3237));
    layer2_outputs(4156) <= (layer1_outputs(4445)) and not (layer1_outputs(3183));
    layer2_outputs(4157) <= not((layer1_outputs(130)) xor (layer1_outputs(2941)));
    layer2_outputs(4158) <= not((layer1_outputs(4790)) xor (layer1_outputs(2605)));
    layer2_outputs(4159) <= not(layer1_outputs(749));
    layer2_outputs(4160) <= layer1_outputs(4949);
    layer2_outputs(4161) <= not((layer1_outputs(3777)) xor (layer1_outputs(2685)));
    layer2_outputs(4162) <= (layer1_outputs(3388)) and not (layer1_outputs(815));
    layer2_outputs(4163) <= (layer1_outputs(572)) xor (layer1_outputs(229));
    layer2_outputs(4164) <= not(layer1_outputs(2219));
    layer2_outputs(4165) <= layer1_outputs(131);
    layer2_outputs(4166) <= not(layer1_outputs(4104)) or (layer1_outputs(134));
    layer2_outputs(4167) <= layer1_outputs(1457);
    layer2_outputs(4168) <= (layer1_outputs(4568)) or (layer1_outputs(429));
    layer2_outputs(4169) <= not(layer1_outputs(4252));
    layer2_outputs(4170) <= not(layer1_outputs(4977)) or (layer1_outputs(2808));
    layer2_outputs(4171) <= layer1_outputs(2112);
    layer2_outputs(4172) <= not(layer1_outputs(588));
    layer2_outputs(4173) <= (layer1_outputs(1206)) and not (layer1_outputs(4651));
    layer2_outputs(4174) <= layer1_outputs(1159);
    layer2_outputs(4175) <= layer1_outputs(4663);
    layer2_outputs(4176) <= layer1_outputs(2626);
    layer2_outputs(4177) <= not(layer1_outputs(1032));
    layer2_outputs(4178) <= (layer1_outputs(803)) xor (layer1_outputs(1784));
    layer2_outputs(4179) <= not(layer1_outputs(1296));
    layer2_outputs(4180) <= not(layer1_outputs(3428));
    layer2_outputs(4181) <= not((layer1_outputs(3759)) or (layer1_outputs(2717)));
    layer2_outputs(4182) <= not((layer1_outputs(2357)) or (layer1_outputs(3042)));
    layer2_outputs(4183) <= (layer1_outputs(2411)) or (layer1_outputs(248));
    layer2_outputs(4184) <= layer1_outputs(3452);
    layer2_outputs(4185) <= '0';
    layer2_outputs(4186) <= not(layer1_outputs(185));
    layer2_outputs(4187) <= '0';
    layer2_outputs(4188) <= not(layer1_outputs(403));
    layer2_outputs(4189) <= not(layer1_outputs(963));
    layer2_outputs(4190) <= layer1_outputs(2061);
    layer2_outputs(4191) <= not(layer1_outputs(4154));
    layer2_outputs(4192) <= not(layer1_outputs(2911)) or (layer1_outputs(4718));
    layer2_outputs(4193) <= not(layer1_outputs(3579));
    layer2_outputs(4194) <= (layer1_outputs(1118)) or (layer1_outputs(4307));
    layer2_outputs(4195) <= not((layer1_outputs(4636)) and (layer1_outputs(3965)));
    layer2_outputs(4196) <= not(layer1_outputs(1641)) or (layer1_outputs(2748));
    layer2_outputs(4197) <= not((layer1_outputs(5080)) xor (layer1_outputs(4234)));
    layer2_outputs(4198) <= not((layer1_outputs(3476)) or (layer1_outputs(3235)));
    layer2_outputs(4199) <= not((layer1_outputs(5043)) and (layer1_outputs(399)));
    layer2_outputs(4200) <= not(layer1_outputs(4891));
    layer2_outputs(4201) <= layer1_outputs(4512);
    layer2_outputs(4202) <= not(layer1_outputs(2001));
    layer2_outputs(4203) <= not(layer1_outputs(2630));
    layer2_outputs(4204) <= not((layer1_outputs(2383)) or (layer1_outputs(3083)));
    layer2_outputs(4205) <= not(layer1_outputs(1912));
    layer2_outputs(4206) <= (layer1_outputs(89)) xor (layer1_outputs(2358));
    layer2_outputs(4207) <= (layer1_outputs(4741)) xor (layer1_outputs(905));
    layer2_outputs(4208) <= (layer1_outputs(390)) or (layer1_outputs(2178));
    layer2_outputs(4209) <= not(layer1_outputs(894)) or (layer1_outputs(2633));
    layer2_outputs(4210) <= layer1_outputs(921);
    layer2_outputs(4211) <= not(layer1_outputs(4353));
    layer2_outputs(4212) <= not(layer1_outputs(4617)) or (layer1_outputs(424));
    layer2_outputs(4213) <= '0';
    layer2_outputs(4214) <= not(layer1_outputs(4208));
    layer2_outputs(4215) <= not(layer1_outputs(4475)) or (layer1_outputs(5045));
    layer2_outputs(4216) <= (layer1_outputs(4936)) or (layer1_outputs(2189));
    layer2_outputs(4217) <= (layer1_outputs(4687)) and not (layer1_outputs(3064));
    layer2_outputs(4218) <= (layer1_outputs(846)) or (layer1_outputs(2917));
    layer2_outputs(4219) <= not((layer1_outputs(1835)) xor (layer1_outputs(962)));
    layer2_outputs(4220) <= not(layer1_outputs(2591));
    layer2_outputs(4221) <= not((layer1_outputs(3389)) xor (layer1_outputs(3374)));
    layer2_outputs(4222) <= not(layer1_outputs(4643));
    layer2_outputs(4223) <= not(layer1_outputs(133)) or (layer1_outputs(1559));
    layer2_outputs(4224) <= not((layer1_outputs(3875)) and (layer1_outputs(4229)));
    layer2_outputs(4225) <= (layer1_outputs(391)) and (layer1_outputs(3557));
    layer2_outputs(4226) <= not((layer1_outputs(3084)) xor (layer1_outputs(2107)));
    layer2_outputs(4227) <= (layer1_outputs(3735)) and not (layer1_outputs(56));
    layer2_outputs(4228) <= not((layer1_outputs(4825)) and (layer1_outputs(2835)));
    layer2_outputs(4229) <= not(layer1_outputs(4118));
    layer2_outputs(4230) <= not(layer1_outputs(4540));
    layer2_outputs(4231) <= layer1_outputs(3951);
    layer2_outputs(4232) <= not(layer1_outputs(3208));
    layer2_outputs(4233) <= layer1_outputs(4862);
    layer2_outputs(4234) <= not(layer1_outputs(4202));
    layer2_outputs(4235) <= not((layer1_outputs(236)) or (layer1_outputs(2614)));
    layer2_outputs(4236) <= (layer1_outputs(4138)) and not (layer1_outputs(2644));
    layer2_outputs(4237) <= not(layer1_outputs(4800));
    layer2_outputs(4238) <= layer1_outputs(4759);
    layer2_outputs(4239) <= not(layer1_outputs(2036)) or (layer1_outputs(3767));
    layer2_outputs(4240) <= not(layer1_outputs(4659));
    layer2_outputs(4241) <= layer1_outputs(170);
    layer2_outputs(4242) <= not((layer1_outputs(2374)) and (layer1_outputs(4396)));
    layer2_outputs(4243) <= not((layer1_outputs(3397)) xor (layer1_outputs(2900)));
    layer2_outputs(4244) <= (layer1_outputs(2472)) and not (layer1_outputs(1511));
    layer2_outputs(4245) <= not((layer1_outputs(1872)) xor (layer1_outputs(4039)));
    layer2_outputs(4246) <= not(layer1_outputs(1409));
    layer2_outputs(4247) <= layer1_outputs(4075);
    layer2_outputs(4248) <= layer1_outputs(4279);
    layer2_outputs(4249) <= not(layer1_outputs(2286));
    layer2_outputs(4250) <= (layer1_outputs(4242)) xor (layer1_outputs(928));
    layer2_outputs(4251) <= (layer1_outputs(577)) and not (layer1_outputs(4324));
    layer2_outputs(4252) <= layer1_outputs(3239);
    layer2_outputs(4253) <= not(layer1_outputs(899));
    layer2_outputs(4254) <= not((layer1_outputs(2907)) xor (layer1_outputs(851)));
    layer2_outputs(4255) <= not((layer1_outputs(1426)) and (layer1_outputs(864)));
    layer2_outputs(4256) <= not((layer1_outputs(5082)) xor (layer1_outputs(438)));
    layer2_outputs(4257) <= not(layer1_outputs(1044));
    layer2_outputs(4258) <= (layer1_outputs(4400)) and (layer1_outputs(2105));
    layer2_outputs(4259) <= layer1_outputs(3211);
    layer2_outputs(4260) <= layer1_outputs(3670);
    layer2_outputs(4261) <= not(layer1_outputs(291));
    layer2_outputs(4262) <= (layer1_outputs(1291)) xor (layer1_outputs(3221));
    layer2_outputs(4263) <= not(layer1_outputs(4784));
    layer2_outputs(4264) <= (layer1_outputs(1231)) and not (layer1_outputs(3021));
    layer2_outputs(4265) <= layer1_outputs(3038);
    layer2_outputs(4266) <= not((layer1_outputs(1498)) and (layer1_outputs(3488)));
    layer2_outputs(4267) <= (layer1_outputs(82)) and (layer1_outputs(3556));
    layer2_outputs(4268) <= not((layer1_outputs(2804)) and (layer1_outputs(610)));
    layer2_outputs(4269) <= '1';
    layer2_outputs(4270) <= layer1_outputs(99);
    layer2_outputs(4271) <= not((layer1_outputs(1275)) xor (layer1_outputs(792)));
    layer2_outputs(4272) <= not((layer1_outputs(4415)) and (layer1_outputs(3781)));
    layer2_outputs(4273) <= not(layer1_outputs(2016));
    layer2_outputs(4274) <= layer1_outputs(2419);
    layer2_outputs(4275) <= (layer1_outputs(4439)) and not (layer1_outputs(3460));
    layer2_outputs(4276) <= (layer1_outputs(1031)) and not (layer1_outputs(1911));
    layer2_outputs(4277) <= not((layer1_outputs(4307)) or (layer1_outputs(2630)));
    layer2_outputs(4278) <= not(layer1_outputs(911));
    layer2_outputs(4279) <= layer1_outputs(3232);
    layer2_outputs(4280) <= not(layer1_outputs(2285));
    layer2_outputs(4281) <= layer1_outputs(2543);
    layer2_outputs(4282) <= not(layer1_outputs(2802)) or (layer1_outputs(2099));
    layer2_outputs(4283) <= not((layer1_outputs(2477)) or (layer1_outputs(1810)));
    layer2_outputs(4284) <= not(layer1_outputs(4669)) or (layer1_outputs(2618));
    layer2_outputs(4285) <= (layer1_outputs(1004)) and not (layer1_outputs(326));
    layer2_outputs(4286) <= not((layer1_outputs(4230)) and (layer1_outputs(1839)));
    layer2_outputs(4287) <= layer1_outputs(5044);
    layer2_outputs(4288) <= (layer1_outputs(4644)) xor (layer1_outputs(4231));
    layer2_outputs(4289) <= layer1_outputs(2667);
    layer2_outputs(4290) <= not(layer1_outputs(1945)) or (layer1_outputs(1967));
    layer2_outputs(4291) <= layer1_outputs(582);
    layer2_outputs(4292) <= (layer1_outputs(2096)) and not (layer1_outputs(1002));
    layer2_outputs(4293) <= not((layer1_outputs(404)) or (layer1_outputs(3788)));
    layer2_outputs(4294) <= layer1_outputs(4103);
    layer2_outputs(4295) <= (layer1_outputs(50)) and not (layer1_outputs(3765));
    layer2_outputs(4296) <= not(layer1_outputs(1914));
    layer2_outputs(4297) <= not(layer1_outputs(1973));
    layer2_outputs(4298) <= layer1_outputs(919);
    layer2_outputs(4299) <= (layer1_outputs(3419)) and not (layer1_outputs(1202));
    layer2_outputs(4300) <= layer1_outputs(2028);
    layer2_outputs(4301) <= not((layer1_outputs(3965)) or (layer1_outputs(882)));
    layer2_outputs(4302) <= '1';
    layer2_outputs(4303) <= layer1_outputs(4728);
    layer2_outputs(4304) <= layer1_outputs(1372);
    layer2_outputs(4305) <= (layer1_outputs(4318)) or (layer1_outputs(2000));
    layer2_outputs(4306) <= not(layer1_outputs(4560));
    layer2_outputs(4307) <= not((layer1_outputs(193)) xor (layer1_outputs(2217)));
    layer2_outputs(4308) <= not((layer1_outputs(4795)) or (layer1_outputs(4295)));
    layer2_outputs(4309) <= not((layer1_outputs(2828)) and (layer1_outputs(2950)));
    layer2_outputs(4310) <= not((layer1_outputs(2618)) and (layer1_outputs(4842)));
    layer2_outputs(4311) <= not((layer1_outputs(4079)) xor (layer1_outputs(3494)));
    layer2_outputs(4312) <= not((layer1_outputs(2735)) and (layer1_outputs(4749)));
    layer2_outputs(4313) <= not(layer1_outputs(2652));
    layer2_outputs(4314) <= (layer1_outputs(3043)) and (layer1_outputs(1793));
    layer2_outputs(4315) <= '0';
    layer2_outputs(4316) <= not(layer1_outputs(3243));
    layer2_outputs(4317) <= not((layer1_outputs(2375)) or (layer1_outputs(1698)));
    layer2_outputs(4318) <= (layer1_outputs(1227)) xor (layer1_outputs(1859));
    layer2_outputs(4319) <= (layer1_outputs(3273)) and (layer1_outputs(24));
    layer2_outputs(4320) <= (layer1_outputs(3277)) and (layer1_outputs(4146));
    layer2_outputs(4321) <= layer1_outputs(4675);
    layer2_outputs(4322) <= not(layer1_outputs(499)) or (layer1_outputs(4441));
    layer2_outputs(4323) <= (layer1_outputs(2986)) and (layer1_outputs(1160));
    layer2_outputs(4324) <= layer1_outputs(856);
    layer2_outputs(4325) <= not((layer1_outputs(980)) and (layer1_outputs(4035)));
    layer2_outputs(4326) <= not((layer1_outputs(4185)) or (layer1_outputs(253)));
    layer2_outputs(4327) <= (layer1_outputs(4856)) and not (layer1_outputs(3687));
    layer2_outputs(4328) <= not((layer1_outputs(2978)) and (layer1_outputs(2888)));
    layer2_outputs(4329) <= not(layer1_outputs(1878));
    layer2_outputs(4330) <= not(layer1_outputs(2841));
    layer2_outputs(4331) <= not(layer1_outputs(2738));
    layer2_outputs(4332) <= not(layer1_outputs(1662));
    layer2_outputs(4333) <= not((layer1_outputs(3535)) or (layer1_outputs(1866)));
    layer2_outputs(4334) <= layer1_outputs(3688);
    layer2_outputs(4335) <= layer1_outputs(3733);
    layer2_outputs(4336) <= layer1_outputs(1852);
    layer2_outputs(4337) <= layer1_outputs(2474);
    layer2_outputs(4338) <= (layer1_outputs(2699)) and (layer1_outputs(4769));
    layer2_outputs(4339) <= '1';
    layer2_outputs(4340) <= not(layer1_outputs(4470)) or (layer1_outputs(33));
    layer2_outputs(4341) <= '0';
    layer2_outputs(4342) <= not((layer1_outputs(168)) xor (layer1_outputs(2315)));
    layer2_outputs(4343) <= not((layer1_outputs(1178)) and (layer1_outputs(2300)));
    layer2_outputs(4344) <= (layer1_outputs(3186)) xor (layer1_outputs(3047));
    layer2_outputs(4345) <= not((layer1_outputs(1360)) or (layer1_outputs(1951)));
    layer2_outputs(4346) <= not(layer1_outputs(54)) or (layer1_outputs(1354));
    layer2_outputs(4347) <= not((layer1_outputs(4264)) xor (layer1_outputs(4657)));
    layer2_outputs(4348) <= not(layer1_outputs(3132)) or (layer1_outputs(605));
    layer2_outputs(4349) <= (layer1_outputs(4068)) and not (layer1_outputs(1926));
    layer2_outputs(4350) <= not((layer1_outputs(45)) or (layer1_outputs(1286)));
    layer2_outputs(4351) <= layer1_outputs(3876);
    layer2_outputs(4352) <= (layer1_outputs(3307)) xor (layer1_outputs(4370));
    layer2_outputs(4353) <= layer1_outputs(800);
    layer2_outputs(4354) <= not(layer1_outputs(113));
    layer2_outputs(4355) <= not(layer1_outputs(2596));
    layer2_outputs(4356) <= '0';
    layer2_outputs(4357) <= not(layer1_outputs(2645));
    layer2_outputs(4358) <= not(layer1_outputs(1964));
    layer2_outputs(4359) <= not(layer1_outputs(3851));
    layer2_outputs(4360) <= (layer1_outputs(310)) or (layer1_outputs(1476));
    layer2_outputs(4361) <= (layer1_outputs(3035)) and not (layer1_outputs(744));
    layer2_outputs(4362) <= layer1_outputs(1530);
    layer2_outputs(4363) <= (layer1_outputs(1903)) xor (layer1_outputs(2827));
    layer2_outputs(4364) <= layer1_outputs(1148);
    layer2_outputs(4365) <= layer1_outputs(4210);
    layer2_outputs(4366) <= not(layer1_outputs(3946));
    layer2_outputs(4367) <= not(layer1_outputs(2186));
    layer2_outputs(4368) <= (layer1_outputs(4521)) xor (layer1_outputs(2274));
    layer2_outputs(4369) <= layer1_outputs(1967);
    layer2_outputs(4370) <= layer1_outputs(2344);
    layer2_outputs(4371) <= not(layer1_outputs(1274));
    layer2_outputs(4372) <= not(layer1_outputs(1186));
    layer2_outputs(4373) <= not(layer1_outputs(1080));
    layer2_outputs(4374) <= not(layer1_outputs(3044));
    layer2_outputs(4375) <= not((layer1_outputs(1860)) and (layer1_outputs(1797)));
    layer2_outputs(4376) <= not(layer1_outputs(5054));
    layer2_outputs(4377) <= '0';
    layer2_outputs(4378) <= layer1_outputs(1868);
    layer2_outputs(4379) <= (layer1_outputs(879)) or (layer1_outputs(3172));
    layer2_outputs(4380) <= (layer1_outputs(156)) and not (layer1_outputs(2977));
    layer2_outputs(4381) <= (layer1_outputs(2155)) or (layer1_outputs(1065));
    layer2_outputs(4382) <= not(layer1_outputs(1280));
    layer2_outputs(4383) <= not((layer1_outputs(3705)) and (layer1_outputs(658)));
    layer2_outputs(4384) <= layer1_outputs(2703);
    layer2_outputs(4385) <= (layer1_outputs(4074)) xor (layer1_outputs(4201));
    layer2_outputs(4386) <= not((layer1_outputs(661)) xor (layer1_outputs(1751)));
    layer2_outputs(4387) <= layer1_outputs(3222);
    layer2_outputs(4388) <= (layer1_outputs(2958)) or (layer1_outputs(4062));
    layer2_outputs(4389) <= layer1_outputs(989);
    layer2_outputs(4390) <= layer1_outputs(2054);
    layer2_outputs(4391) <= not(layer1_outputs(4171)) or (layer1_outputs(135));
    layer2_outputs(4392) <= layer1_outputs(3517);
    layer2_outputs(4393) <= layer1_outputs(2409);
    layer2_outputs(4394) <= (layer1_outputs(3018)) xor (layer1_outputs(4566));
    layer2_outputs(4395) <= not((layer1_outputs(1614)) and (layer1_outputs(87)));
    layer2_outputs(4396) <= not(layer1_outputs(992)) or (layer1_outputs(2027));
    layer2_outputs(4397) <= layer1_outputs(1337);
    layer2_outputs(4398) <= (layer1_outputs(4066)) and (layer1_outputs(1849));
    layer2_outputs(4399) <= not(layer1_outputs(3282));
    layer2_outputs(4400) <= not(layer1_outputs(3166)) or (layer1_outputs(105));
    layer2_outputs(4401) <= layer1_outputs(2955);
    layer2_outputs(4402) <= layer1_outputs(1503);
    layer2_outputs(4403) <= not((layer1_outputs(4727)) and (layer1_outputs(1956)));
    layer2_outputs(4404) <= layer1_outputs(1254);
    layer2_outputs(4405) <= layer1_outputs(4678);
    layer2_outputs(4406) <= not(layer1_outputs(1401));
    layer2_outputs(4407) <= not(layer1_outputs(4831)) or (layer1_outputs(2821));
    layer2_outputs(4408) <= layer1_outputs(1515);
    layer2_outputs(4409) <= (layer1_outputs(2071)) or (layer1_outputs(4055));
    layer2_outputs(4410) <= layer1_outputs(4757);
    layer2_outputs(4411) <= (layer1_outputs(4702)) or (layer1_outputs(3979));
    layer2_outputs(4412) <= not(layer1_outputs(512));
    layer2_outputs(4413) <= layer1_outputs(798);
    layer2_outputs(4414) <= not(layer1_outputs(3318));
    layer2_outputs(4415) <= not(layer1_outputs(2450));
    layer2_outputs(4416) <= not(layer1_outputs(1698));
    layer2_outputs(4417) <= layer1_outputs(1707);
    layer2_outputs(4418) <= (layer1_outputs(2502)) xor (layer1_outputs(1290));
    layer2_outputs(4419) <= not(layer1_outputs(3756));
    layer2_outputs(4420) <= not(layer1_outputs(3911)) or (layer1_outputs(3863));
    layer2_outputs(4421) <= not(layer1_outputs(4761));
    layer2_outputs(4422) <= layer1_outputs(2743);
    layer2_outputs(4423) <= (layer1_outputs(2276)) and not (layer1_outputs(2801));
    layer2_outputs(4424) <= not(layer1_outputs(1810));
    layer2_outputs(4425) <= not(layer1_outputs(1037)) or (layer1_outputs(4682));
    layer2_outputs(4426) <= not(layer1_outputs(1628));
    layer2_outputs(4427) <= not((layer1_outputs(653)) or (layer1_outputs(2568)));
    layer2_outputs(4428) <= not(layer1_outputs(4838));
    layer2_outputs(4429) <= not(layer1_outputs(877));
    layer2_outputs(4430) <= not((layer1_outputs(1281)) xor (layer1_outputs(1738)));
    layer2_outputs(4431) <= not((layer1_outputs(4456)) and (layer1_outputs(253)));
    layer2_outputs(4432) <= not(layer1_outputs(3944));
    layer2_outputs(4433) <= layer1_outputs(2980);
    layer2_outputs(4434) <= not(layer1_outputs(3463)) or (layer1_outputs(4207));
    layer2_outputs(4435) <= not((layer1_outputs(3680)) and (layer1_outputs(3742)));
    layer2_outputs(4436) <= layer1_outputs(818);
    layer2_outputs(4437) <= layer1_outputs(4263);
    layer2_outputs(4438) <= layer1_outputs(806);
    layer2_outputs(4439) <= (layer1_outputs(58)) xor (layer1_outputs(4532));
    layer2_outputs(4440) <= (layer1_outputs(53)) or (layer1_outputs(160));
    layer2_outputs(4441) <= (layer1_outputs(2466)) or (layer1_outputs(4794));
    layer2_outputs(4442) <= not((layer1_outputs(4361)) xor (layer1_outputs(1072)));
    layer2_outputs(4443) <= (layer1_outputs(2081)) or (layer1_outputs(3063));
    layer2_outputs(4444) <= not((layer1_outputs(1584)) xor (layer1_outputs(1620)));
    layer2_outputs(4445) <= layer1_outputs(1763);
    layer2_outputs(4446) <= (layer1_outputs(4747)) and not (layer1_outputs(124));
    layer2_outputs(4447) <= not((layer1_outputs(1466)) xor (layer1_outputs(1442)));
    layer2_outputs(4448) <= not((layer1_outputs(1935)) xor (layer1_outputs(4921)));
    layer2_outputs(4449) <= layer1_outputs(680);
    layer2_outputs(4450) <= not((layer1_outputs(1650)) xor (layer1_outputs(3684)));
    layer2_outputs(4451) <= layer1_outputs(1336);
    layer2_outputs(4452) <= not(layer1_outputs(3867));
    layer2_outputs(4453) <= layer1_outputs(1141);
    layer2_outputs(4454) <= not(layer1_outputs(3256));
    layer2_outputs(4455) <= not(layer1_outputs(304)) or (layer1_outputs(1042));
    layer2_outputs(4456) <= layer1_outputs(4054);
    layer2_outputs(4457) <= not(layer1_outputs(2395));
    layer2_outputs(4458) <= (layer1_outputs(1512)) xor (layer1_outputs(4116));
    layer2_outputs(4459) <= not(layer1_outputs(2884));
    layer2_outputs(4460) <= (layer1_outputs(4422)) xor (layer1_outputs(2669));
    layer2_outputs(4461) <= not(layer1_outputs(1332)) or (layer1_outputs(2586));
    layer2_outputs(4462) <= layer1_outputs(2093);
    layer2_outputs(4463) <= (layer1_outputs(2329)) and not (layer1_outputs(3188));
    layer2_outputs(4464) <= '0';
    layer2_outputs(4465) <= not(layer1_outputs(2972));
    layer2_outputs(4466) <= layer1_outputs(4826);
    layer2_outputs(4467) <= layer1_outputs(312);
    layer2_outputs(4468) <= not(layer1_outputs(2530)) or (layer1_outputs(3655));
    layer2_outputs(4469) <= (layer1_outputs(3091)) and (layer1_outputs(969));
    layer2_outputs(4470) <= (layer1_outputs(4874)) and not (layer1_outputs(81));
    layer2_outputs(4471) <= not(layer1_outputs(3229));
    layer2_outputs(4472) <= not(layer1_outputs(908));
    layer2_outputs(4473) <= not(layer1_outputs(3498));
    layer2_outputs(4474) <= '0';
    layer2_outputs(4475) <= layer1_outputs(3981);
    layer2_outputs(4476) <= layer1_outputs(4608);
    layer2_outputs(4477) <= not((layer1_outputs(2455)) xor (layer1_outputs(2055)));
    layer2_outputs(4478) <= not(layer1_outputs(174));
    layer2_outputs(4479) <= (layer1_outputs(5069)) and not (layer1_outputs(3191));
    layer2_outputs(4480) <= not(layer1_outputs(3297));
    layer2_outputs(4481) <= not(layer1_outputs(4897)) or (layer1_outputs(2372));
    layer2_outputs(4482) <= (layer1_outputs(2925)) and not (layer1_outputs(3259));
    layer2_outputs(4483) <= layer1_outputs(3510);
    layer2_outputs(4484) <= (layer1_outputs(3477)) xor (layer1_outputs(2992));
    layer2_outputs(4485) <= not(layer1_outputs(1789));
    layer2_outputs(4486) <= not(layer1_outputs(3266));
    layer2_outputs(4487) <= not(layer1_outputs(467)) or (layer1_outputs(4136));
    layer2_outputs(4488) <= not(layer1_outputs(3157)) or (layer1_outputs(237));
    layer2_outputs(4489) <= layer1_outputs(939);
    layer2_outputs(4490) <= not(layer1_outputs(1802)) or (layer1_outputs(2449));
    layer2_outputs(4491) <= (layer1_outputs(871)) or (layer1_outputs(4598));
    layer2_outputs(4492) <= (layer1_outputs(2988)) and (layer1_outputs(1224));
    layer2_outputs(4493) <= not(layer1_outputs(1437));
    layer2_outputs(4494) <= not(layer1_outputs(2958));
    layer2_outputs(4495) <= not(layer1_outputs(4411));
    layer2_outputs(4496) <= layer1_outputs(2714);
    layer2_outputs(4497) <= (layer1_outputs(2129)) xor (layer1_outputs(2255));
    layer2_outputs(4498) <= not((layer1_outputs(228)) or (layer1_outputs(1768)));
    layer2_outputs(4499) <= not((layer1_outputs(1673)) or (layer1_outputs(2962)));
    layer2_outputs(4500) <= (layer1_outputs(976)) and not (layer1_outputs(1308));
    layer2_outputs(4501) <= not(layer1_outputs(322));
    layer2_outputs(4502) <= (layer1_outputs(191)) and (layer1_outputs(1920));
    layer2_outputs(4503) <= not(layer1_outputs(4626)) or (layer1_outputs(4942));
    layer2_outputs(4504) <= layer1_outputs(5028);
    layer2_outputs(4505) <= not(layer1_outputs(4032));
    layer2_outputs(4506) <= not(layer1_outputs(4677)) or (layer1_outputs(2791));
    layer2_outputs(4507) <= (layer1_outputs(3559)) and not (layer1_outputs(2317));
    layer2_outputs(4508) <= not(layer1_outputs(3632));
    layer2_outputs(4509) <= layer1_outputs(2435);
    layer2_outputs(4510) <= (layer1_outputs(1172)) and not (layer1_outputs(2724));
    layer2_outputs(4511) <= not(layer1_outputs(3575));
    layer2_outputs(4512) <= not(layer1_outputs(1400)) or (layer1_outputs(3621));
    layer2_outputs(4513) <= (layer1_outputs(4073)) xor (layer1_outputs(3922));
    layer2_outputs(4514) <= layer1_outputs(2888);
    layer2_outputs(4515) <= layer1_outputs(3686);
    layer2_outputs(4516) <= layer1_outputs(4786);
    layer2_outputs(4517) <= '0';
    layer2_outputs(4518) <= (layer1_outputs(1739)) and not (layer1_outputs(317));
    layer2_outputs(4519) <= layer1_outputs(2501);
    layer2_outputs(4520) <= layer1_outputs(1265);
    layer2_outputs(4521) <= not((layer1_outputs(2174)) xor (layer1_outputs(2266)));
    layer2_outputs(4522) <= layer1_outputs(3973);
    layer2_outputs(4523) <= (layer1_outputs(810)) or (layer1_outputs(1066));
    layer2_outputs(4524) <= layer1_outputs(2072);
    layer2_outputs(4525) <= not((layer1_outputs(1226)) xor (layer1_outputs(3748)));
    layer2_outputs(4526) <= (layer1_outputs(3286)) xor (layer1_outputs(3380));
    layer2_outputs(4527) <= (layer1_outputs(4004)) and (layer1_outputs(1664));
    layer2_outputs(4528) <= not((layer1_outputs(2891)) or (layer1_outputs(1455)));
    layer2_outputs(4529) <= not(layer1_outputs(4917));
    layer2_outputs(4530) <= layer1_outputs(3601);
    layer2_outputs(4531) <= layer1_outputs(977);
    layer2_outputs(4532) <= layer1_outputs(4254);
    layer2_outputs(4533) <= (layer1_outputs(1305)) xor (layer1_outputs(4723));
    layer2_outputs(4534) <= '0';
    layer2_outputs(4535) <= layer1_outputs(2060);
    layer2_outputs(4536) <= layer1_outputs(2867);
    layer2_outputs(4537) <= layer1_outputs(2054);
    layer2_outputs(4538) <= not(layer1_outputs(4774)) or (layer1_outputs(4324));
    layer2_outputs(4539) <= (layer1_outputs(4562)) and not (layer1_outputs(949));
    layer2_outputs(4540) <= layer1_outputs(3340);
    layer2_outputs(4541) <= not(layer1_outputs(1997));
    layer2_outputs(4542) <= not(layer1_outputs(5067));
    layer2_outputs(4543) <= (layer1_outputs(3554)) and not (layer1_outputs(2968));
    layer2_outputs(4544) <= not(layer1_outputs(4270));
    layer2_outputs(4545) <= layer1_outputs(1353);
    layer2_outputs(4546) <= not(layer1_outputs(3623));
    layer2_outputs(4547) <= (layer1_outputs(3071)) or (layer1_outputs(2227));
    layer2_outputs(4548) <= not(layer1_outputs(879));
    layer2_outputs(4549) <= layer1_outputs(3947);
    layer2_outputs(4550) <= not(layer1_outputs(3790));
    layer2_outputs(4551) <= layer1_outputs(2916);
    layer2_outputs(4552) <= not(layer1_outputs(270));
    layer2_outputs(4553) <= layer1_outputs(2493);
    layer2_outputs(4554) <= not(layer1_outputs(743));
    layer2_outputs(4555) <= layer1_outputs(122);
    layer2_outputs(4556) <= not((layer1_outputs(1438)) xor (layer1_outputs(3898)));
    layer2_outputs(4557) <= not(layer1_outputs(1820));
    layer2_outputs(4558) <= (layer1_outputs(4666)) and (layer1_outputs(1414));
    layer2_outputs(4559) <= layer1_outputs(589);
    layer2_outputs(4560) <= layer1_outputs(1550);
    layer2_outputs(4561) <= layer1_outputs(2299);
    layer2_outputs(4562) <= not((layer1_outputs(4268)) or (layer1_outputs(3939)));
    layer2_outputs(4563) <= (layer1_outputs(3512)) or (layer1_outputs(3967));
    layer2_outputs(4564) <= not(layer1_outputs(4085));
    layer2_outputs(4565) <= not(layer1_outputs(1224)) or (layer1_outputs(2110));
    layer2_outputs(4566) <= not(layer1_outputs(4198)) or (layer1_outputs(3144));
    layer2_outputs(4567) <= not((layer1_outputs(4058)) and (layer1_outputs(3858)));
    layer2_outputs(4568) <= not(layer1_outputs(2567));
    layer2_outputs(4569) <= not((layer1_outputs(3463)) and (layer1_outputs(1068)));
    layer2_outputs(4570) <= layer1_outputs(4971);
    layer2_outputs(4571) <= not(layer1_outputs(258));
    layer2_outputs(4572) <= not(layer1_outputs(1549));
    layer2_outputs(4573) <= not(layer1_outputs(4720));
    layer2_outputs(4574) <= layer1_outputs(1756);
    layer2_outputs(4575) <= layer1_outputs(1497);
    layer2_outputs(4576) <= not(layer1_outputs(3845));
    layer2_outputs(4577) <= (layer1_outputs(1310)) and not (layer1_outputs(1371));
    layer2_outputs(4578) <= (layer1_outputs(4640)) and not (layer1_outputs(4072));
    layer2_outputs(4579) <= layer1_outputs(4131);
    layer2_outputs(4580) <= layer1_outputs(3386);
    layer2_outputs(4581) <= not(layer1_outputs(5097));
    layer2_outputs(4582) <= layer1_outputs(2300);
    layer2_outputs(4583) <= not(layer1_outputs(3775));
    layer2_outputs(4584) <= not((layer1_outputs(2741)) and (layer1_outputs(5011)));
    layer2_outputs(4585) <= layer1_outputs(1127);
    layer2_outputs(4586) <= not((layer1_outputs(379)) and (layer1_outputs(69)));
    layer2_outputs(4587) <= not(layer1_outputs(583));
    layer2_outputs(4588) <= not(layer1_outputs(4498));
    layer2_outputs(4589) <= (layer1_outputs(2731)) and not (layer1_outputs(537));
    layer2_outputs(4590) <= not((layer1_outputs(1075)) xor (layer1_outputs(4896)));
    layer2_outputs(4591) <= (layer1_outputs(4507)) xor (layer1_outputs(2343));
    layer2_outputs(4592) <= layer1_outputs(1764);
    layer2_outputs(4593) <= '1';
    layer2_outputs(4594) <= not((layer1_outputs(1429)) xor (layer1_outputs(34)));
    layer2_outputs(4595) <= not(layer1_outputs(2224));
    layer2_outputs(4596) <= (layer1_outputs(3603)) and not (layer1_outputs(3068));
    layer2_outputs(4597) <= not((layer1_outputs(3607)) or (layer1_outputs(356)));
    layer2_outputs(4598) <= not(layer1_outputs(657));
    layer2_outputs(4599) <= not((layer1_outputs(1119)) xor (layer1_outputs(3425)));
    layer2_outputs(4600) <= (layer1_outputs(475)) xor (layer1_outputs(57));
    layer2_outputs(4601) <= not(layer1_outputs(2227)) or (layer1_outputs(1749));
    layer2_outputs(4602) <= (layer1_outputs(1878)) and not (layer1_outputs(2581));
    layer2_outputs(4603) <= layer1_outputs(3253);
    layer2_outputs(4604) <= (layer1_outputs(452)) and not (layer1_outputs(612));
    layer2_outputs(4605) <= not(layer1_outputs(2155));
    layer2_outputs(4606) <= (layer1_outputs(2487)) and (layer1_outputs(3024));
    layer2_outputs(4607) <= not((layer1_outputs(419)) xor (layer1_outputs(1756)));
    layer2_outputs(4608) <= (layer1_outputs(4281)) xor (layer1_outputs(2239));
    layer2_outputs(4609) <= layer1_outputs(4084);
    layer2_outputs(4610) <= (layer1_outputs(4169)) and not (layer1_outputs(4525));
    layer2_outputs(4611) <= layer1_outputs(1375);
    layer2_outputs(4612) <= not(layer1_outputs(166));
    layer2_outputs(4613) <= not(layer1_outputs(2556)) or (layer1_outputs(1121));
    layer2_outputs(4614) <= layer1_outputs(636);
    layer2_outputs(4615) <= (layer1_outputs(5022)) or (layer1_outputs(840));
    layer2_outputs(4616) <= not(layer1_outputs(2675));
    layer2_outputs(4617) <= not(layer1_outputs(2201));
    layer2_outputs(4618) <= layer1_outputs(4875);
    layer2_outputs(4619) <= layer1_outputs(2188);
    layer2_outputs(4620) <= (layer1_outputs(3689)) and not (layer1_outputs(2311));
    layer2_outputs(4621) <= not((layer1_outputs(2852)) and (layer1_outputs(2831)));
    layer2_outputs(4622) <= not(layer1_outputs(3024));
    layer2_outputs(4623) <= not(layer1_outputs(642)) or (layer1_outputs(3333));
    layer2_outputs(4624) <= not(layer1_outputs(3431));
    layer2_outputs(4625) <= '1';
    layer2_outputs(4626) <= layer1_outputs(1088);
    layer2_outputs(4627) <= (layer1_outputs(1153)) and not (layer1_outputs(363));
    layer2_outputs(4628) <= (layer1_outputs(5107)) and not (layer1_outputs(2135));
    layer2_outputs(4629) <= not(layer1_outputs(249));
    layer2_outputs(4630) <= not((layer1_outputs(3304)) and (layer1_outputs(3897)));
    layer2_outputs(4631) <= not(layer1_outputs(1318)) or (layer1_outputs(1018));
    layer2_outputs(4632) <= layer1_outputs(243);
    layer2_outputs(4633) <= '1';
    layer2_outputs(4634) <= layer1_outputs(1406);
    layer2_outputs(4635) <= not((layer1_outputs(200)) or (layer1_outputs(4798)));
    layer2_outputs(4636) <= (layer1_outputs(869)) xor (layer1_outputs(1410));
    layer2_outputs(4637) <= not((layer1_outputs(2933)) and (layer1_outputs(3008)));
    layer2_outputs(4638) <= (layer1_outputs(2100)) xor (layer1_outputs(2382));
    layer2_outputs(4639) <= (layer1_outputs(3394)) and (layer1_outputs(265));
    layer2_outputs(4640) <= not((layer1_outputs(1923)) xor (layer1_outputs(4192)));
    layer2_outputs(4641) <= layer1_outputs(5061);
    layer2_outputs(4642) <= layer1_outputs(2704);
    layer2_outputs(4643) <= not(layer1_outputs(1152));
    layer2_outputs(4644) <= (layer1_outputs(1748)) and not (layer1_outputs(4488));
    layer2_outputs(4645) <= (layer1_outputs(4572)) and not (layer1_outputs(4989));
    layer2_outputs(4646) <= not(layer1_outputs(4907));
    layer2_outputs(4647) <= not(layer1_outputs(4653));
    layer2_outputs(4648) <= layer1_outputs(1892);
    layer2_outputs(4649) <= not((layer1_outputs(4722)) and (layer1_outputs(3856)));
    layer2_outputs(4650) <= not(layer1_outputs(1075));
    layer2_outputs(4651) <= layer1_outputs(207);
    layer2_outputs(4652) <= not((layer1_outputs(1991)) xor (layer1_outputs(4992)));
    layer2_outputs(4653) <= layer1_outputs(1599);
    layer2_outputs(4654) <= (layer1_outputs(1303)) or (layer1_outputs(3193));
    layer2_outputs(4655) <= not(layer1_outputs(399)) or (layer1_outputs(3286));
    layer2_outputs(4656) <= layer1_outputs(410);
    layer2_outputs(4657) <= not(layer1_outputs(2405)) or (layer1_outputs(481));
    layer2_outputs(4658) <= not(layer1_outputs(2017)) or (layer1_outputs(4309));
    layer2_outputs(4659) <= not(layer1_outputs(31)) or (layer1_outputs(2573));
    layer2_outputs(4660) <= not(layer1_outputs(1917)) or (layer1_outputs(1493));
    layer2_outputs(4661) <= layer1_outputs(925);
    layer2_outputs(4662) <= not(layer1_outputs(1298));
    layer2_outputs(4663) <= (layer1_outputs(3700)) or (layer1_outputs(141));
    layer2_outputs(4664) <= layer1_outputs(205);
    layer2_outputs(4665) <= not(layer1_outputs(232));
    layer2_outputs(4666) <= layer1_outputs(4012);
    layer2_outputs(4667) <= (layer1_outputs(3056)) and (layer1_outputs(4565));
    layer2_outputs(4668) <= not((layer1_outputs(3549)) xor (layer1_outputs(1638)));
    layer2_outputs(4669) <= not(layer1_outputs(4452));
    layer2_outputs(4670) <= not(layer1_outputs(4417)) or (layer1_outputs(3843));
    layer2_outputs(4671) <= layer1_outputs(2687);
    layer2_outputs(4672) <= layer1_outputs(2975);
    layer2_outputs(4673) <= not((layer1_outputs(3111)) or (layer1_outputs(2823)));
    layer2_outputs(4674) <= (layer1_outputs(3663)) or (layer1_outputs(829));
    layer2_outputs(4675) <= not((layer1_outputs(4853)) and (layer1_outputs(248)));
    layer2_outputs(4676) <= not(layer1_outputs(96));
    layer2_outputs(4677) <= not(layer1_outputs(4647));
    layer2_outputs(4678) <= not(layer1_outputs(1502));
    layer2_outputs(4679) <= (layer1_outputs(873)) and not (layer1_outputs(228));
    layer2_outputs(4680) <= (layer1_outputs(3565)) xor (layer1_outputs(409));
    layer2_outputs(4681) <= layer1_outputs(223);
    layer2_outputs(4682) <= (layer1_outputs(513)) and not (layer1_outputs(4170));
    layer2_outputs(4683) <= not(layer1_outputs(3232));
    layer2_outputs(4684) <= layer1_outputs(15);
    layer2_outputs(4685) <= layer1_outputs(5112);
    layer2_outputs(4686) <= layer1_outputs(3931);
    layer2_outputs(4687) <= not(layer1_outputs(1430)) or (layer1_outputs(2191));
    layer2_outputs(4688) <= not((layer1_outputs(1603)) and (layer1_outputs(3130)));
    layer2_outputs(4689) <= not(layer1_outputs(2471));
    layer2_outputs(4690) <= layer1_outputs(3060);
    layer2_outputs(4691) <= (layer1_outputs(2079)) xor (layer1_outputs(2374));
    layer2_outputs(4692) <= not(layer1_outputs(3089));
    layer2_outputs(4693) <= (layer1_outputs(688)) or (layer1_outputs(913));
    layer2_outputs(4694) <= (layer1_outputs(529)) xor (layer1_outputs(3292));
    layer2_outputs(4695) <= not((layer1_outputs(2068)) xor (layer1_outputs(2190)));
    layer2_outputs(4696) <= (layer1_outputs(4750)) and (layer1_outputs(622));
    layer2_outputs(4697) <= not(layer1_outputs(2014)) or (layer1_outputs(2248));
    layer2_outputs(4698) <= not((layer1_outputs(809)) and (layer1_outputs(634)));
    layer2_outputs(4699) <= layer1_outputs(4340);
    layer2_outputs(4700) <= (layer1_outputs(3301)) and not (layer1_outputs(2727));
    layer2_outputs(4701) <= not(layer1_outputs(4047));
    layer2_outputs(4702) <= not((layer1_outputs(2605)) and (layer1_outputs(4744)));
    layer2_outputs(4703) <= not(layer1_outputs(3247));
    layer2_outputs(4704) <= not((layer1_outputs(1000)) xor (layer1_outputs(2496)));
    layer2_outputs(4705) <= (layer1_outputs(4506)) xor (layer1_outputs(4578));
    layer2_outputs(4706) <= (layer1_outputs(93)) and not (layer1_outputs(1486));
    layer2_outputs(4707) <= (layer1_outputs(837)) and not (layer1_outputs(3775));
    layer2_outputs(4708) <= layer1_outputs(2635);
    layer2_outputs(4709) <= not(layer1_outputs(1998)) or (layer1_outputs(2662));
    layer2_outputs(4710) <= not(layer1_outputs(783));
    layer2_outputs(4711) <= not(layer1_outputs(2180)) or (layer1_outputs(1218));
    layer2_outputs(4712) <= not(layer1_outputs(4353));
    layer2_outputs(4713) <= (layer1_outputs(3466)) and not (layer1_outputs(4110));
    layer2_outputs(4714) <= (layer1_outputs(5118)) and not (layer1_outputs(3177));
    layer2_outputs(4715) <= not((layer1_outputs(3059)) and (layer1_outputs(1432)));
    layer2_outputs(4716) <= layer1_outputs(553);
    layer2_outputs(4717) <= not((layer1_outputs(116)) or (layer1_outputs(2101)));
    layer2_outputs(4718) <= (layer1_outputs(4732)) or (layer1_outputs(4515));
    layer2_outputs(4719) <= not(layer1_outputs(1847));
    layer2_outputs(4720) <= not((layer1_outputs(1394)) xor (layer1_outputs(1750)));
    layer2_outputs(4721) <= layer1_outputs(2885);
    layer2_outputs(4722) <= (layer1_outputs(5001)) and not (layer1_outputs(4195));
    layer2_outputs(4723) <= (layer1_outputs(3697)) xor (layer1_outputs(854));
    layer2_outputs(4724) <= not(layer1_outputs(3792)) or (layer1_outputs(3203));
    layer2_outputs(4725) <= layer1_outputs(1273);
    layer2_outputs(4726) <= not(layer1_outputs(2109));
    layer2_outputs(4727) <= layer1_outputs(2942);
    layer2_outputs(4728) <= not(layer1_outputs(2818));
    layer2_outputs(4729) <= (layer1_outputs(3596)) and (layer1_outputs(3646));
    layer2_outputs(4730) <= not(layer1_outputs(1151));
    layer2_outputs(4731) <= layer1_outputs(482);
    layer2_outputs(4732) <= not(layer1_outputs(4859));
    layer2_outputs(4733) <= (layer1_outputs(2737)) xor (layer1_outputs(835));
    layer2_outputs(4734) <= (layer1_outputs(4877)) and not (layer1_outputs(4575));
    layer2_outputs(4735) <= (layer1_outputs(80)) and (layer1_outputs(1574));
    layer2_outputs(4736) <= '1';
    layer2_outputs(4737) <= not(layer1_outputs(2461)) or (layer1_outputs(1615));
    layer2_outputs(4738) <= not((layer1_outputs(1460)) or (layer1_outputs(1352)));
    layer2_outputs(4739) <= (layer1_outputs(1744)) xor (layer1_outputs(4766));
    layer2_outputs(4740) <= '0';
    layer2_outputs(4741) <= layer1_outputs(4410);
    layer2_outputs(4742) <= layer1_outputs(3076);
    layer2_outputs(4743) <= (layer1_outputs(3460)) and not (layer1_outputs(2499));
    layer2_outputs(4744) <= not(layer1_outputs(4780));
    layer2_outputs(4745) <= (layer1_outputs(3748)) and not (layer1_outputs(1267));
    layer2_outputs(4746) <= not(layer1_outputs(2636));
    layer2_outputs(4747) <= (layer1_outputs(1149)) and not (layer1_outputs(1897));
    layer2_outputs(4748) <= not(layer1_outputs(5079)) or (layer1_outputs(3605));
    layer2_outputs(4749) <= (layer1_outputs(516)) or (layer1_outputs(3470));
    layer2_outputs(4750) <= (layer1_outputs(3093)) xor (layer1_outputs(3939));
    layer2_outputs(4751) <= not((layer1_outputs(3242)) xor (layer1_outputs(2134)));
    layer2_outputs(4752) <= not(layer1_outputs(4197));
    layer2_outputs(4753) <= not(layer1_outputs(1942)) or (layer1_outputs(3513));
    layer2_outputs(4754) <= layer1_outputs(61);
    layer2_outputs(4755) <= not(layer1_outputs(2053)) or (layer1_outputs(4219));
    layer2_outputs(4756) <= layer1_outputs(4511);
    layer2_outputs(4757) <= not((layer1_outputs(4048)) xor (layer1_outputs(3899)));
    layer2_outputs(4758) <= (layer1_outputs(5033)) and (layer1_outputs(4154));
    layer2_outputs(4759) <= not((layer1_outputs(1280)) or (layer1_outputs(1420)));
    layer2_outputs(4760) <= '1';
    layer2_outputs(4761) <= (layer1_outputs(2902)) or (layer1_outputs(574));
    layer2_outputs(4762) <= not(layer1_outputs(2305));
    layer2_outputs(4763) <= not((layer1_outputs(3763)) or (layer1_outputs(2657)));
    layer2_outputs(4764) <= layer1_outputs(1441);
    layer2_outputs(4765) <= (layer1_outputs(1391)) and (layer1_outputs(2555));
    layer2_outputs(4766) <= (layer1_outputs(502)) and not (layer1_outputs(549));
    layer2_outputs(4767) <= not(layer1_outputs(3025));
    layer2_outputs(4768) <= (layer1_outputs(4573)) and (layer1_outputs(3085));
    layer2_outputs(4769) <= layer1_outputs(173);
    layer2_outputs(4770) <= (layer1_outputs(3488)) and not (layer1_outputs(1655));
    layer2_outputs(4771) <= layer1_outputs(3813);
    layer2_outputs(4772) <= (layer1_outputs(4872)) and (layer1_outputs(2278));
    layer2_outputs(4773) <= not(layer1_outputs(4534));
    layer2_outputs(4774) <= not(layer1_outputs(3370)) or (layer1_outputs(4763));
    layer2_outputs(4775) <= not(layer1_outputs(4929)) or (layer1_outputs(536));
    layer2_outputs(4776) <= not((layer1_outputs(1571)) and (layer1_outputs(1693)));
    layer2_outputs(4777) <= not(layer1_outputs(111));
    layer2_outputs(4778) <= (layer1_outputs(1197)) and not (layer1_outputs(4252));
    layer2_outputs(4779) <= (layer1_outputs(4745)) or (layer1_outputs(4321));
    layer2_outputs(4780) <= not(layer1_outputs(2246));
    layer2_outputs(4781) <= layer1_outputs(964);
    layer2_outputs(4782) <= (layer1_outputs(508)) and not (layer1_outputs(4931));
    layer2_outputs(4783) <= '0';
    layer2_outputs(4784) <= not(layer1_outputs(415)) or (layer1_outputs(330));
    layer2_outputs(4785) <= layer1_outputs(4205);
    layer2_outputs(4786) <= (layer1_outputs(113)) xor (layer1_outputs(2894));
    layer2_outputs(4787) <= (layer1_outputs(1557)) and (layer1_outputs(4552));
    layer2_outputs(4788) <= not(layer1_outputs(4638));
    layer2_outputs(4789) <= (layer1_outputs(799)) and not (layer1_outputs(4299));
    layer2_outputs(4790) <= not((layer1_outputs(768)) xor (layer1_outputs(3865)));
    layer2_outputs(4791) <= not(layer1_outputs(275));
    layer2_outputs(4792) <= not(layer1_outputs(1139));
    layer2_outputs(4793) <= not(layer1_outputs(737)) or (layer1_outputs(1192));
    layer2_outputs(4794) <= (layer1_outputs(4299)) or (layer1_outputs(5107));
    layer2_outputs(4795) <= not(layer1_outputs(2696)) or (layer1_outputs(4923));
    layer2_outputs(4796) <= not(layer1_outputs(2383));
    layer2_outputs(4797) <= layer1_outputs(5085);
    layer2_outputs(4798) <= layer1_outputs(3368);
    layer2_outputs(4799) <= layer1_outputs(4802);
    layer2_outputs(4800) <= not(layer1_outputs(309)) or (layer1_outputs(3833));
    layer2_outputs(4801) <= not((layer1_outputs(1464)) and (layer1_outputs(698)));
    layer2_outputs(4802) <= layer1_outputs(4036);
    layer2_outputs(4803) <= layer1_outputs(5000);
    layer2_outputs(4804) <= not(layer1_outputs(4628));
    layer2_outputs(4805) <= (layer1_outputs(1488)) and not (layer1_outputs(1788));
    layer2_outputs(4806) <= not((layer1_outputs(1827)) xor (layer1_outputs(5040)));
    layer2_outputs(4807) <= not(layer1_outputs(121));
    layer2_outputs(4808) <= (layer1_outputs(1926)) xor (layer1_outputs(3050));
    layer2_outputs(4809) <= not(layer1_outputs(654));
    layer2_outputs(4810) <= not(layer1_outputs(4020));
    layer2_outputs(4811) <= not(layer1_outputs(4039));
    layer2_outputs(4812) <= (layer1_outputs(1837)) and not (layer1_outputs(1791));
    layer2_outputs(4813) <= layer1_outputs(1311);
    layer2_outputs(4814) <= (layer1_outputs(3442)) and (layer1_outputs(659));
    layer2_outputs(4815) <= (layer1_outputs(1895)) and not (layer1_outputs(3355));
    layer2_outputs(4816) <= not(layer1_outputs(4736));
    layer2_outputs(4817) <= not((layer1_outputs(2008)) xor (layer1_outputs(4323)));
    layer2_outputs(4818) <= not(layer1_outputs(4270));
    layer2_outputs(4819) <= not(layer1_outputs(2119));
    layer2_outputs(4820) <= layer1_outputs(133);
    layer2_outputs(4821) <= (layer1_outputs(59)) and not (layer1_outputs(247));
    layer2_outputs(4822) <= not((layer1_outputs(3381)) or (layer1_outputs(4616)));
    layer2_outputs(4823) <= not(layer1_outputs(2400));
    layer2_outputs(4824) <= not(layer1_outputs(1287));
    layer2_outputs(4825) <= layer1_outputs(1058);
    layer2_outputs(4826) <= not(layer1_outputs(3561)) or (layer1_outputs(4044));
    layer2_outputs(4827) <= not(layer1_outputs(127));
    layer2_outputs(4828) <= not(layer1_outputs(3953));
    layer2_outputs(4829) <= not(layer1_outputs(146));
    layer2_outputs(4830) <= (layer1_outputs(655)) or (layer1_outputs(148));
    layer2_outputs(4831) <= layer1_outputs(275);
    layer2_outputs(4832) <= not(layer1_outputs(2336));
    layer2_outputs(4833) <= layer1_outputs(1936);
    layer2_outputs(4834) <= (layer1_outputs(3217)) and not (layer1_outputs(4001));
    layer2_outputs(4835) <= not(layer1_outputs(5014));
    layer2_outputs(4836) <= layer1_outputs(308);
    layer2_outputs(4837) <= layer1_outputs(435);
    layer2_outputs(4838) <= not((layer1_outputs(4075)) or (layer1_outputs(4699)));
    layer2_outputs(4839) <= (layer1_outputs(169)) xor (layer1_outputs(2667));
    layer2_outputs(4840) <= not(layer1_outputs(611)) or (layer1_outputs(4157));
    layer2_outputs(4841) <= not((layer1_outputs(479)) or (layer1_outputs(3389)));
    layer2_outputs(4842) <= layer1_outputs(2740);
    layer2_outputs(4843) <= (layer1_outputs(3841)) and not (layer1_outputs(1591));
    layer2_outputs(4844) <= not(layer1_outputs(4903)) or (layer1_outputs(1678));
    layer2_outputs(4845) <= layer1_outputs(4968);
    layer2_outputs(4846) <= (layer1_outputs(324)) and (layer1_outputs(378));
    layer2_outputs(4847) <= (layer1_outputs(1623)) or (layer1_outputs(2126));
    layer2_outputs(4848) <= (layer1_outputs(3773)) xor (layer1_outputs(3591));
    layer2_outputs(4849) <= not(layer1_outputs(2707)) or (layer1_outputs(1837));
    layer2_outputs(4850) <= not((layer1_outputs(4629)) xor (layer1_outputs(2226)));
    layer2_outputs(4851) <= layer1_outputs(4198);
    layer2_outputs(4852) <= not((layer1_outputs(4623)) xor (layer1_outputs(4788)));
    layer2_outputs(4853) <= (layer1_outputs(4184)) and not (layer1_outputs(4389));
    layer2_outputs(4854) <= not((layer1_outputs(2115)) or (layer1_outputs(4620)));
    layer2_outputs(4855) <= not(layer1_outputs(3459));
    layer2_outputs(4856) <= (layer1_outputs(2729)) and not (layer1_outputs(2979));
    layer2_outputs(4857) <= (layer1_outputs(4404)) and (layer1_outputs(770));
    layer2_outputs(4858) <= not(layer1_outputs(1366));
    layer2_outputs(4859) <= not(layer1_outputs(1460));
    layer2_outputs(4860) <= (layer1_outputs(951)) xor (layer1_outputs(477));
    layer2_outputs(4861) <= not((layer1_outputs(4534)) and (layer1_outputs(4121)));
    layer2_outputs(4862) <= layer1_outputs(1882);
    layer2_outputs(4863) <= layer1_outputs(1149);
    layer2_outputs(4864) <= (layer1_outputs(2104)) and not (layer1_outputs(2460));
    layer2_outputs(4865) <= not((layer1_outputs(1196)) and (layer1_outputs(4138)));
    layer2_outputs(4866) <= not((layer1_outputs(3584)) and (layer1_outputs(2448)));
    layer2_outputs(4867) <= (layer1_outputs(4352)) and (layer1_outputs(3921));
    layer2_outputs(4868) <= layer1_outputs(1595);
    layer2_outputs(4869) <= not(layer1_outputs(3106));
    layer2_outputs(4870) <= (layer1_outputs(1230)) xor (layer1_outputs(914));
    layer2_outputs(4871) <= not(layer1_outputs(2242));
    layer2_outputs(4872) <= (layer1_outputs(4006)) and (layer1_outputs(2868));
    layer2_outputs(4873) <= layer1_outputs(1966);
    layer2_outputs(4874) <= layer1_outputs(2410);
    layer2_outputs(4875) <= not(layer1_outputs(2087));
    layer2_outputs(4876) <= layer1_outputs(1452);
    layer2_outputs(4877) <= layer1_outputs(1671);
    layer2_outputs(4878) <= not((layer1_outputs(3351)) and (layer1_outputs(1962)));
    layer2_outputs(4879) <= not(layer1_outputs(1492));
    layer2_outputs(4880) <= not(layer1_outputs(3627));
    layer2_outputs(4881) <= (layer1_outputs(4752)) and not (layer1_outputs(1861));
    layer2_outputs(4882) <= not((layer1_outputs(674)) xor (layer1_outputs(4194)));
    layer2_outputs(4883) <= (layer1_outputs(4203)) and (layer1_outputs(4446));
    layer2_outputs(4884) <= not(layer1_outputs(3964)) or (layer1_outputs(1784));
    layer2_outputs(4885) <= not(layer1_outputs(4496));
    layer2_outputs(4886) <= (layer1_outputs(2597)) xor (layer1_outputs(1337));
    layer2_outputs(4887) <= (layer1_outputs(450)) and not (layer1_outputs(4591));
    layer2_outputs(4888) <= not(layer1_outputs(3956));
    layer2_outputs(4889) <= not(layer1_outputs(1683));
    layer2_outputs(4890) <= layer1_outputs(1008);
    layer2_outputs(4891) <= not(layer1_outputs(2509));
    layer2_outputs(4892) <= layer1_outputs(1036);
    layer2_outputs(4893) <= not(layer1_outputs(1891));
    layer2_outputs(4894) <= not(layer1_outputs(3146));
    layer2_outputs(4895) <= layer1_outputs(2325);
    layer2_outputs(4896) <= not(layer1_outputs(790));
    layer2_outputs(4897) <= not(layer1_outputs(5085));
    layer2_outputs(4898) <= (layer1_outputs(4474)) xor (layer1_outputs(4323));
    layer2_outputs(4899) <= (layer1_outputs(2858)) and (layer1_outputs(1225));
    layer2_outputs(4900) <= not(layer1_outputs(4076)) or (layer1_outputs(4259));
    layer2_outputs(4901) <= layer1_outputs(861);
    layer2_outputs(4902) <= not(layer1_outputs(500)) or (layer1_outputs(343));
    layer2_outputs(4903) <= (layer1_outputs(1124)) and (layer1_outputs(1054));
    layer2_outputs(4904) <= not((layer1_outputs(1352)) and (layer1_outputs(4656)));
    layer2_outputs(4905) <= layer1_outputs(2515);
    layer2_outputs(4906) <= not(layer1_outputs(3994));
    layer2_outputs(4907) <= not((layer1_outputs(1796)) and (layer1_outputs(492)));
    layer2_outputs(4908) <= not(layer1_outputs(4408)) or (layer1_outputs(3678));
    layer2_outputs(4909) <= layer1_outputs(1130);
    layer2_outputs(4910) <= not(layer1_outputs(281));
    layer2_outputs(4911) <= layer1_outputs(267);
    layer2_outputs(4912) <= layer1_outputs(2716);
    layer2_outputs(4913) <= layer1_outputs(2642);
    layer2_outputs(4914) <= (layer1_outputs(562)) and (layer1_outputs(3750));
    layer2_outputs(4915) <= layer1_outputs(2844);
    layer2_outputs(4916) <= (layer1_outputs(4662)) and (layer1_outputs(4904));
    layer2_outputs(4917) <= not(layer1_outputs(224)) or (layer1_outputs(1823));
    layer2_outputs(4918) <= (layer1_outputs(1778)) and not (layer1_outputs(851));
    layer2_outputs(4919) <= (layer1_outputs(3051)) and not (layer1_outputs(4595));
    layer2_outputs(4920) <= not(layer1_outputs(2089));
    layer2_outputs(4921) <= layer1_outputs(4031);
    layer2_outputs(4922) <= layer1_outputs(3486);
    layer2_outputs(4923) <= layer1_outputs(377);
    layer2_outputs(4924) <= not((layer1_outputs(4297)) or (layer1_outputs(3545)));
    layer2_outputs(4925) <= layer1_outputs(3986);
    layer2_outputs(4926) <= not(layer1_outputs(3626));
    layer2_outputs(4927) <= not(layer1_outputs(2722)) or (layer1_outputs(4242));
    layer2_outputs(4928) <= (layer1_outputs(651)) and not (layer1_outputs(4611));
    layer2_outputs(4929) <= (layer1_outputs(1208)) and not (layer1_outputs(2302));
    layer2_outputs(4930) <= layer1_outputs(5100);
    layer2_outputs(4931) <= not((layer1_outputs(1300)) or (layer1_outputs(3728)));
    layer2_outputs(4932) <= not(layer1_outputs(2384));
    layer2_outputs(4933) <= (layer1_outputs(2673)) and (layer1_outputs(539));
    layer2_outputs(4934) <= not(layer1_outputs(3712)) or (layer1_outputs(34));
    layer2_outputs(4935) <= not(layer1_outputs(4271));
    layer2_outputs(4936) <= not((layer1_outputs(5056)) or (layer1_outputs(4165)));
    layer2_outputs(4937) <= not((layer1_outputs(826)) xor (layer1_outputs(4809)));
    layer2_outputs(4938) <= not(layer1_outputs(97));
    layer2_outputs(4939) <= (layer1_outputs(3508)) and not (layer1_outputs(731));
    layer2_outputs(4940) <= not(layer1_outputs(3170));
    layer2_outputs(4941) <= layer1_outputs(1468);
    layer2_outputs(4942) <= not(layer1_outputs(2847));
    layer2_outputs(4943) <= (layer1_outputs(741)) xor (layer1_outputs(1374));
    layer2_outputs(4944) <= layer1_outputs(4645);
    layer2_outputs(4945) <= not(layer1_outputs(494)) or (layer1_outputs(1866));
    layer2_outputs(4946) <= not(layer1_outputs(667)) or (layer1_outputs(906));
    layer2_outputs(4947) <= layer1_outputs(795);
    layer2_outputs(4948) <= (layer1_outputs(5109)) and not (layer1_outputs(1160));
    layer2_outputs(4949) <= not(layer1_outputs(1901)) or (layer1_outputs(771));
    layer2_outputs(4950) <= layer1_outputs(3979);
    layer2_outputs(4951) <= not((layer1_outputs(2009)) and (layer1_outputs(828)));
    layer2_outputs(4952) <= not(layer1_outputs(2627));
    layer2_outputs(4953) <= not(layer1_outputs(1117)) or (layer1_outputs(3169));
    layer2_outputs(4954) <= (layer1_outputs(2570)) or (layer1_outputs(3477));
    layer2_outputs(4955) <= not(layer1_outputs(2831));
    layer2_outputs(4956) <= layer1_outputs(1774);
    layer2_outputs(4957) <= (layer1_outputs(4976)) and (layer1_outputs(80));
    layer2_outputs(4958) <= not(layer1_outputs(1041));
    layer2_outputs(4959) <= layer1_outputs(3091);
    layer2_outputs(4960) <= not(layer1_outputs(276));
    layer2_outputs(4961) <= not(layer1_outputs(588)) or (layer1_outputs(4513));
    layer2_outputs(4962) <= (layer1_outputs(3831)) or (layer1_outputs(4820));
    layer2_outputs(4963) <= (layer1_outputs(4190)) and not (layer1_outputs(1474));
    layer2_outputs(4964) <= not(layer1_outputs(844));
    layer2_outputs(4965) <= (layer1_outputs(349)) xor (layer1_outputs(2813));
    layer2_outputs(4966) <= not((layer1_outputs(4460)) and (layer1_outputs(1557)));
    layer2_outputs(4967) <= not(layer1_outputs(4817));
    layer2_outputs(4968) <= not(layer1_outputs(3666));
    layer2_outputs(4969) <= layer1_outputs(3249);
    layer2_outputs(4970) <= layer1_outputs(4779);
    layer2_outputs(4971) <= not((layer1_outputs(4003)) or (layer1_outputs(819)));
    layer2_outputs(4972) <= layer1_outputs(3224);
    layer2_outputs(4973) <= not((layer1_outputs(2730)) or (layer1_outputs(2386)));
    layer2_outputs(4974) <= layer1_outputs(3486);
    layer2_outputs(4975) <= not((layer1_outputs(359)) xor (layer1_outputs(4674)));
    layer2_outputs(4976) <= (layer1_outputs(1294)) or (layer1_outputs(5015));
    layer2_outputs(4977) <= not(layer1_outputs(3359));
    layer2_outputs(4978) <= (layer1_outputs(3464)) and not (layer1_outputs(4990));
    layer2_outputs(4979) <= not((layer1_outputs(2468)) xor (layer1_outputs(1834)));
    layer2_outputs(4980) <= layer1_outputs(1621);
    layer2_outputs(4981) <= not(layer1_outputs(3781)) or (layer1_outputs(2848));
    layer2_outputs(4982) <= not((layer1_outputs(1597)) or (layer1_outputs(2648)));
    layer2_outputs(4983) <= layer1_outputs(2550);
    layer2_outputs(4984) <= (layer1_outputs(4684)) and not (layer1_outputs(4038));
    layer2_outputs(4985) <= not((layer1_outputs(152)) xor (layer1_outputs(355)));
    layer2_outputs(4986) <= layer1_outputs(867);
    layer2_outputs(4987) <= not(layer1_outputs(3149));
    layer2_outputs(4988) <= layer1_outputs(5052);
    layer2_outputs(4989) <= not(layer1_outputs(3400));
    layer2_outputs(4990) <= not(layer1_outputs(4583)) or (layer1_outputs(1523));
    layer2_outputs(4991) <= not(layer1_outputs(3564));
    layer2_outputs(4992) <= layer1_outputs(197);
    layer2_outputs(4993) <= layer1_outputs(3285);
    layer2_outputs(4994) <= (layer1_outputs(2770)) xor (layer1_outputs(4492));
    layer2_outputs(4995) <= not(layer1_outputs(5029)) or (layer1_outputs(1422));
    layer2_outputs(4996) <= (layer1_outputs(4561)) xor (layer1_outputs(3107));
    layer2_outputs(4997) <= layer1_outputs(1488);
    layer2_outputs(4998) <= not(layer1_outputs(4669));
    layer2_outputs(4999) <= not(layer1_outputs(896));
    layer2_outputs(5000) <= not(layer1_outputs(3751));
    layer2_outputs(5001) <= layer1_outputs(1916);
    layer2_outputs(5002) <= not(layer1_outputs(214));
    layer2_outputs(5003) <= layer1_outputs(813);
    layer2_outputs(5004) <= not((layer1_outputs(4149)) xor (layer1_outputs(2453)));
    layer2_outputs(5005) <= not(layer1_outputs(2527));
    layer2_outputs(5006) <= layer1_outputs(789);
    layer2_outputs(5007) <= not((layer1_outputs(1844)) or (layer1_outputs(4638)));
    layer2_outputs(5008) <= not(layer1_outputs(4498));
    layer2_outputs(5009) <= not(layer1_outputs(1030));
    layer2_outputs(5010) <= (layer1_outputs(3675)) and (layer1_outputs(3989));
    layer2_outputs(5011) <= (layer1_outputs(2647)) and (layer1_outputs(4536));
    layer2_outputs(5012) <= (layer1_outputs(2543)) and not (layer1_outputs(1955));
    layer2_outputs(5013) <= layer1_outputs(4903);
    layer2_outputs(5014) <= layer1_outputs(4974);
    layer2_outputs(5015) <= (layer1_outputs(740)) and not (layer1_outputs(4962));
    layer2_outputs(5016) <= layer1_outputs(2197);
    layer2_outputs(5017) <= (layer1_outputs(4601)) and not (layer1_outputs(1165));
    layer2_outputs(5018) <= (layer1_outputs(2267)) and not (layer1_outputs(1694));
    layer2_outputs(5019) <= (layer1_outputs(6)) and not (layer1_outputs(1648));
    layer2_outputs(5020) <= layer1_outputs(1372);
    layer2_outputs(5021) <= (layer1_outputs(3155)) and (layer1_outputs(2681));
    layer2_outputs(5022) <= not(layer1_outputs(4937)) or (layer1_outputs(1959));
    layer2_outputs(5023) <= not(layer1_outputs(4885)) or (layer1_outputs(4931));
    layer2_outputs(5024) <= not(layer1_outputs(2162)) or (layer1_outputs(3287));
    layer2_outputs(5025) <= not(layer1_outputs(1976));
    layer2_outputs(5026) <= layer1_outputs(4560);
    layer2_outputs(5027) <= layer1_outputs(2229);
    layer2_outputs(5028) <= not(layer1_outputs(1750));
    layer2_outputs(5029) <= not(layer1_outputs(1316));
    layer2_outputs(5030) <= (layer1_outputs(4646)) and not (layer1_outputs(3837));
    layer2_outputs(5031) <= layer1_outputs(554);
    layer2_outputs(5032) <= not(layer1_outputs(4668));
    layer2_outputs(5033) <= layer1_outputs(2188);
    layer2_outputs(5034) <= not(layer1_outputs(1186));
    layer2_outputs(5035) <= not(layer1_outputs(4607));
    layer2_outputs(5036) <= not(layer1_outputs(4668)) or (layer1_outputs(77));
    layer2_outputs(5037) <= not(layer1_outputs(2082));
    layer2_outputs(5038) <= not(layer1_outputs(1498));
    layer2_outputs(5039) <= not((layer1_outputs(1469)) xor (layer1_outputs(2079)));
    layer2_outputs(5040) <= not((layer1_outputs(4069)) xor (layer1_outputs(4179)));
    layer2_outputs(5041) <= layer1_outputs(4862);
    layer2_outputs(5042) <= not(layer1_outputs(1182)) or (layer1_outputs(4827));
    layer2_outputs(5043) <= not((layer1_outputs(2530)) xor (layer1_outputs(3432)));
    layer2_outputs(5044) <= not(layer1_outputs(4058));
    layer2_outputs(5045) <= not(layer1_outputs(1138));
    layer2_outputs(5046) <= layer1_outputs(1419);
    layer2_outputs(5047) <= not(layer1_outputs(313));
    layer2_outputs(5048) <= not(layer1_outputs(159));
    layer2_outputs(5049) <= (layer1_outputs(1183)) or (layer1_outputs(3473));
    layer2_outputs(5050) <= (layer1_outputs(3541)) and (layer1_outputs(4980));
    layer2_outputs(5051) <= layer1_outputs(3933);
    layer2_outputs(5052) <= (layer1_outputs(737)) and not (layer1_outputs(4908));
    layer2_outputs(5053) <= not((layer1_outputs(2945)) xor (layer1_outputs(1295)));
    layer2_outputs(5054) <= not((layer1_outputs(4166)) and (layer1_outputs(986)));
    layer2_outputs(5055) <= (layer1_outputs(2800)) and not (layer1_outputs(2786));
    layer2_outputs(5056) <= not(layer1_outputs(4797));
    layer2_outputs(5057) <= layer1_outputs(1056);
    layer2_outputs(5058) <= (layer1_outputs(465)) and (layer1_outputs(3754));
    layer2_outputs(5059) <= layer1_outputs(1306);
    layer2_outputs(5060) <= (layer1_outputs(1888)) xor (layer1_outputs(5019));
    layer2_outputs(5061) <= not(layer1_outputs(2697)) or (layer1_outputs(4827));
    layer2_outputs(5062) <= layer1_outputs(515);
    layer2_outputs(5063) <= not(layer1_outputs(4160)) or (layer1_outputs(407));
    layer2_outputs(5064) <= (layer1_outputs(952)) xor (layer1_outputs(1477));
    layer2_outputs(5065) <= not(layer1_outputs(1408));
    layer2_outputs(5066) <= not((layer1_outputs(1588)) or (layer1_outputs(120)));
    layer2_outputs(5067) <= (layer1_outputs(1788)) and (layer1_outputs(108));
    layer2_outputs(5068) <= not((layer1_outputs(1715)) or (layer1_outputs(75)));
    layer2_outputs(5069) <= (layer1_outputs(87)) and not (layer1_outputs(17));
    layer2_outputs(5070) <= (layer1_outputs(3408)) and (layer1_outputs(4928));
    layer2_outputs(5071) <= (layer1_outputs(4710)) and not (layer1_outputs(3974));
    layer2_outputs(5072) <= (layer1_outputs(3639)) and (layer1_outputs(2649));
    layer2_outputs(5073) <= (layer1_outputs(1205)) xor (layer1_outputs(4686));
    layer2_outputs(5074) <= not(layer1_outputs(83));
    layer2_outputs(5075) <= layer1_outputs(1231);
    layer2_outputs(5076) <= not(layer1_outputs(144)) or (layer1_outputs(3321));
    layer2_outputs(5077) <= layer1_outputs(3581);
    layer2_outputs(5078) <= (layer1_outputs(523)) and not (layer1_outputs(1439));
    layer2_outputs(5079) <= not(layer1_outputs(1827));
    layer2_outputs(5080) <= layer1_outputs(3006);
    layer2_outputs(5081) <= not(layer1_outputs(4599));
    layer2_outputs(5082) <= (layer1_outputs(3343)) and not (layer1_outputs(492));
    layer2_outputs(5083) <= not(layer1_outputs(2328));
    layer2_outputs(5084) <= layer1_outputs(1902);
    layer2_outputs(5085) <= (layer1_outputs(3574)) and (layer1_outputs(1202));
    layer2_outputs(5086) <= not(layer1_outputs(1157));
    layer2_outputs(5087) <= (layer1_outputs(3343)) and not (layer1_outputs(2820));
    layer2_outputs(5088) <= not(layer1_outputs(2733));
    layer2_outputs(5089) <= not((layer1_outputs(2985)) xor (layer1_outputs(4378)));
    layer2_outputs(5090) <= not(layer1_outputs(4261)) or (layer1_outputs(2649));
    layer2_outputs(5091) <= not(layer1_outputs(478));
    layer2_outputs(5092) <= (layer1_outputs(518)) xor (layer1_outputs(2861));
    layer2_outputs(5093) <= not((layer1_outputs(4920)) and (layer1_outputs(3364)));
    layer2_outputs(5094) <= layer1_outputs(3916);
    layer2_outputs(5095) <= not(layer1_outputs(4407));
    layer2_outputs(5096) <= (layer1_outputs(936)) and (layer1_outputs(1070));
    layer2_outputs(5097) <= layer1_outputs(3443);
    layer2_outputs(5098) <= not(layer1_outputs(3759)) or (layer1_outputs(1306));
    layer2_outputs(5099) <= not(layer1_outputs(2271));
    layer2_outputs(5100) <= not(layer1_outputs(753));
    layer2_outputs(5101) <= (layer1_outputs(3095)) and not (layer1_outputs(4366));
    layer2_outputs(5102) <= not(layer1_outputs(128));
    layer2_outputs(5103) <= layer1_outputs(1553);
    layer2_outputs(5104) <= not(layer1_outputs(3482));
    layer2_outputs(5105) <= not(layer1_outputs(1272));
    layer2_outputs(5106) <= not((layer1_outputs(4245)) or (layer1_outputs(199)));
    layer2_outputs(5107) <= not(layer1_outputs(493)) or (layer1_outputs(1253));
    layer2_outputs(5108) <= layer1_outputs(4591);
    layer2_outputs(5109) <= layer1_outputs(1147);
    layer2_outputs(5110) <= (layer1_outputs(3011)) or (layer1_outputs(3161));
    layer2_outputs(5111) <= not(layer1_outputs(4848));
    layer2_outputs(5112) <= layer1_outputs(1851);
    layer2_outputs(5113) <= layer1_outputs(4636);
    layer2_outputs(5114) <= layer1_outputs(694);
    layer2_outputs(5115) <= not(layer1_outputs(1414));
    layer2_outputs(5116) <= not(layer1_outputs(505));
    layer2_outputs(5117) <= layer1_outputs(600);
    layer2_outputs(5118) <= layer1_outputs(3919);
    layer2_outputs(5119) <= layer1_outputs(2369);
    outputs(0) <= layer2_outputs(489);
    outputs(1) <= layer2_outputs(4432);
    outputs(2) <= not(layer2_outputs(2188));
    outputs(3) <= not(layer2_outputs(1084));
    outputs(4) <= (layer2_outputs(2982)) or (layer2_outputs(4409));
    outputs(5) <= layer2_outputs(2009);
    outputs(6) <= not(layer2_outputs(4962));
    outputs(7) <= layer2_outputs(4612);
    outputs(8) <= layer2_outputs(1451);
    outputs(9) <= layer2_outputs(3071);
    outputs(10) <= not(layer2_outputs(1141));
    outputs(11) <= not(layer2_outputs(544));
    outputs(12) <= layer2_outputs(1140);
    outputs(13) <= (layer2_outputs(3545)) xor (layer2_outputs(3639));
    outputs(14) <= not((layer2_outputs(3555)) xor (layer2_outputs(2396)));
    outputs(15) <= not(layer2_outputs(2094));
    outputs(16) <= not(layer2_outputs(1285));
    outputs(17) <= layer2_outputs(1786);
    outputs(18) <= layer2_outputs(398);
    outputs(19) <= not((layer2_outputs(1272)) xor (layer2_outputs(4542)));
    outputs(20) <= not((layer2_outputs(2573)) xor (layer2_outputs(412)));
    outputs(21) <= not(layer2_outputs(2072)) or (layer2_outputs(2470));
    outputs(22) <= layer2_outputs(2852);
    outputs(23) <= (layer2_outputs(3103)) xor (layer2_outputs(4877));
    outputs(24) <= not(layer2_outputs(3449));
    outputs(25) <= layer2_outputs(2100);
    outputs(26) <= not((layer2_outputs(2143)) xor (layer2_outputs(3349)));
    outputs(27) <= (layer2_outputs(2493)) xor (layer2_outputs(1593));
    outputs(28) <= not((layer2_outputs(5095)) or (layer2_outputs(4879)));
    outputs(29) <= not(layer2_outputs(1428));
    outputs(30) <= not(layer2_outputs(4349));
    outputs(31) <= not(layer2_outputs(1060));
    outputs(32) <= not(layer2_outputs(3634));
    outputs(33) <= not(layer2_outputs(361));
    outputs(34) <= not(layer2_outputs(4608));
    outputs(35) <= not(layer2_outputs(1866));
    outputs(36) <= not(layer2_outputs(3844));
    outputs(37) <= not(layer2_outputs(1284));
    outputs(38) <= not(layer2_outputs(4425));
    outputs(39) <= not(layer2_outputs(2908));
    outputs(40) <= (layer2_outputs(2199)) xor (layer2_outputs(4872));
    outputs(41) <= not(layer2_outputs(238));
    outputs(42) <= not(layer2_outputs(2167));
    outputs(43) <= (layer2_outputs(2287)) xor (layer2_outputs(1618));
    outputs(44) <= layer2_outputs(3684);
    outputs(45) <= layer2_outputs(247);
    outputs(46) <= not(layer2_outputs(1040));
    outputs(47) <= layer2_outputs(3251);
    outputs(48) <= layer2_outputs(1696);
    outputs(49) <= not((layer2_outputs(4995)) xor (layer2_outputs(2277)));
    outputs(50) <= not(layer2_outputs(4838));
    outputs(51) <= layer2_outputs(1808);
    outputs(52) <= layer2_outputs(3916);
    outputs(53) <= (layer2_outputs(4922)) xor (layer2_outputs(3845));
    outputs(54) <= layer2_outputs(4207);
    outputs(55) <= (layer2_outputs(810)) xor (layer2_outputs(1209));
    outputs(56) <= not(layer2_outputs(2735));
    outputs(57) <= not(layer2_outputs(5020));
    outputs(58) <= layer2_outputs(4326);
    outputs(59) <= not(layer2_outputs(3838));
    outputs(60) <= (layer2_outputs(4936)) or (layer2_outputs(5097));
    outputs(61) <= not(layer2_outputs(1197));
    outputs(62) <= layer2_outputs(449);
    outputs(63) <= (layer2_outputs(4022)) and (layer2_outputs(4288));
    outputs(64) <= not(layer2_outputs(2582));
    outputs(65) <= not((layer2_outputs(2479)) xor (layer2_outputs(4792)));
    outputs(66) <= not((layer2_outputs(2273)) and (layer2_outputs(4416)));
    outputs(67) <= layer2_outputs(360);
    outputs(68) <= not(layer2_outputs(1650));
    outputs(69) <= not(layer2_outputs(1953)) or (layer2_outputs(1412));
    outputs(70) <= (layer2_outputs(1475)) xor (layer2_outputs(1431));
    outputs(71) <= not(layer2_outputs(3170));
    outputs(72) <= layer2_outputs(2187);
    outputs(73) <= not(layer2_outputs(3017)) or (layer2_outputs(1495));
    outputs(74) <= not(layer2_outputs(1543));
    outputs(75) <= not((layer2_outputs(1922)) xor (layer2_outputs(3203)));
    outputs(76) <= (layer2_outputs(863)) xor (layer2_outputs(3616));
    outputs(77) <= not(layer2_outputs(4599));
    outputs(78) <= (layer2_outputs(2564)) xor (layer2_outputs(4534));
    outputs(79) <= not((layer2_outputs(4751)) xor (layer2_outputs(5003)));
    outputs(80) <= layer2_outputs(3293);
    outputs(81) <= not(layer2_outputs(325));
    outputs(82) <= layer2_outputs(4364);
    outputs(83) <= (layer2_outputs(3471)) and (layer2_outputs(4857));
    outputs(84) <= not((layer2_outputs(1490)) xor (layer2_outputs(3073)));
    outputs(85) <= not(layer2_outputs(2085));
    outputs(86) <= not(layer2_outputs(1229));
    outputs(87) <= not(layer2_outputs(3734)) or (layer2_outputs(1499));
    outputs(88) <= not((layer2_outputs(1120)) or (layer2_outputs(1117)));
    outputs(89) <= not(layer2_outputs(4200));
    outputs(90) <= not(layer2_outputs(4594));
    outputs(91) <= not(layer2_outputs(3747));
    outputs(92) <= layer2_outputs(4866);
    outputs(93) <= layer2_outputs(859);
    outputs(94) <= '0';
    outputs(95) <= not(layer2_outputs(3146));
    outputs(96) <= (layer2_outputs(185)) and (layer2_outputs(3079));
    outputs(97) <= not((layer2_outputs(5042)) xor (layer2_outputs(1679)));
    outputs(98) <= not(layer2_outputs(1584));
    outputs(99) <= not(layer2_outputs(3228));
    outputs(100) <= layer2_outputs(4280);
    outputs(101) <= layer2_outputs(1116);
    outputs(102) <= not((layer2_outputs(4551)) and (layer2_outputs(4201)));
    outputs(103) <= not(layer2_outputs(3666));
    outputs(104) <= layer2_outputs(1522);
    outputs(105) <= not((layer2_outputs(3276)) or (layer2_outputs(655)));
    outputs(106) <= not(layer2_outputs(1712)) or (layer2_outputs(3575));
    outputs(107) <= not(layer2_outputs(2378));
    outputs(108) <= (layer2_outputs(3906)) or (layer2_outputs(1073));
    outputs(109) <= not(layer2_outputs(710));
    outputs(110) <= (layer2_outputs(2868)) xor (layer2_outputs(4405));
    outputs(111) <= not(layer2_outputs(2926));
    outputs(112) <= not(layer2_outputs(2956));
    outputs(113) <= layer2_outputs(24);
    outputs(114) <= (layer2_outputs(2854)) and (layer2_outputs(2934));
    outputs(115) <= not(layer2_outputs(759)) or (layer2_outputs(1864));
    outputs(116) <= not(layer2_outputs(3747));
    outputs(117) <= (layer2_outputs(496)) and (layer2_outputs(3485));
    outputs(118) <= not(layer2_outputs(3921));
    outputs(119) <= layer2_outputs(4324);
    outputs(120) <= not(layer2_outputs(4588));
    outputs(121) <= (layer2_outputs(4178)) xor (layer2_outputs(1701));
    outputs(122) <= (layer2_outputs(4755)) and not (layer2_outputs(2416));
    outputs(123) <= not((layer2_outputs(2197)) xor (layer2_outputs(385)));
    outputs(124) <= layer2_outputs(368);
    outputs(125) <= not(layer2_outputs(3641));
    outputs(126) <= not(layer2_outputs(2962));
    outputs(127) <= layer2_outputs(2897);
    outputs(128) <= layer2_outputs(3166);
    outputs(129) <= layer2_outputs(1004);
    outputs(130) <= not(layer2_outputs(375));
    outputs(131) <= not(layer2_outputs(3372));
    outputs(132) <= not(layer2_outputs(1179));
    outputs(133) <= not(layer2_outputs(1027));
    outputs(134) <= not((layer2_outputs(3123)) xor (layer2_outputs(2279)));
    outputs(135) <= (layer2_outputs(2683)) and (layer2_outputs(797));
    outputs(136) <= layer2_outputs(5069);
    outputs(137) <= not(layer2_outputs(1330));
    outputs(138) <= layer2_outputs(371);
    outputs(139) <= layer2_outputs(4821);
    outputs(140) <= layer2_outputs(2446);
    outputs(141) <= layer2_outputs(4741);
    outputs(142) <= not(layer2_outputs(4112));
    outputs(143) <= layer2_outputs(3304);
    outputs(144) <= not(layer2_outputs(4564));
    outputs(145) <= layer2_outputs(68);
    outputs(146) <= not(layer2_outputs(3048));
    outputs(147) <= layer2_outputs(1847);
    outputs(148) <= layer2_outputs(1639);
    outputs(149) <= not(layer2_outputs(3699));
    outputs(150) <= layer2_outputs(336);
    outputs(151) <= not((layer2_outputs(311)) xor (layer2_outputs(1593)));
    outputs(152) <= not(layer2_outputs(4619));
    outputs(153) <= (layer2_outputs(274)) xor (layer2_outputs(4206));
    outputs(154) <= layer2_outputs(3789);
    outputs(155) <= not(layer2_outputs(4536)) or (layer2_outputs(4011));
    outputs(156) <= layer2_outputs(1051);
    outputs(157) <= layer2_outputs(3202);
    outputs(158) <= not(layer2_outputs(119));
    outputs(159) <= layer2_outputs(1365);
    outputs(160) <= not((layer2_outputs(1512)) or (layer2_outputs(3419)));
    outputs(161) <= not(layer2_outputs(1031));
    outputs(162) <= not(layer2_outputs(2163));
    outputs(163) <= layer2_outputs(3661);
    outputs(164) <= layer2_outputs(944);
    outputs(165) <= not((layer2_outputs(3105)) or (layer2_outputs(3682)));
    outputs(166) <= layer2_outputs(3034);
    outputs(167) <= layer2_outputs(3019);
    outputs(168) <= not(layer2_outputs(1992));
    outputs(169) <= (layer2_outputs(2510)) or (layer2_outputs(4643));
    outputs(170) <= layer2_outputs(4989);
    outputs(171) <= (layer2_outputs(1946)) and (layer2_outputs(2731));
    outputs(172) <= layer2_outputs(3006);
    outputs(173) <= not(layer2_outputs(1744)) or (layer2_outputs(1373));
    outputs(174) <= layer2_outputs(4218);
    outputs(175) <= not(layer2_outputs(3160));
    outputs(176) <= layer2_outputs(3056);
    outputs(177) <= not(layer2_outputs(954));
    outputs(178) <= not(layer2_outputs(276));
    outputs(179) <= (layer2_outputs(3055)) and not (layer2_outputs(4913));
    outputs(180) <= not(layer2_outputs(1314));
    outputs(181) <= layer2_outputs(4955);
    outputs(182) <= (layer2_outputs(3674)) and not (layer2_outputs(1002));
    outputs(183) <= not(layer2_outputs(1665)) or (layer2_outputs(1251));
    outputs(184) <= not(layer2_outputs(2901));
    outputs(185) <= not((layer2_outputs(629)) xor (layer2_outputs(4893)));
    outputs(186) <= layer2_outputs(2666);
    outputs(187) <= layer2_outputs(3440);
    outputs(188) <= not(layer2_outputs(1101));
    outputs(189) <= layer2_outputs(4287);
    outputs(190) <= not((layer2_outputs(907)) and (layer2_outputs(3100)));
    outputs(191) <= layer2_outputs(3533);
    outputs(192) <= not(layer2_outputs(3444));
    outputs(193) <= layer2_outputs(2930);
    outputs(194) <= not((layer2_outputs(3393)) xor (layer2_outputs(4092)));
    outputs(195) <= layer2_outputs(3696);
    outputs(196) <= not(layer2_outputs(3328)) or (layer2_outputs(2786));
    outputs(197) <= not((layer2_outputs(3633)) and (layer2_outputs(2396)));
    outputs(198) <= not(layer2_outputs(1521));
    outputs(199) <= not(layer2_outputs(1664));
    outputs(200) <= not(layer2_outputs(3882)) or (layer2_outputs(83));
    outputs(201) <= layer2_outputs(4387);
    outputs(202) <= not(layer2_outputs(1681));
    outputs(203) <= layer2_outputs(208);
    outputs(204) <= (layer2_outputs(1091)) xor (layer2_outputs(3318));
    outputs(205) <= layer2_outputs(1361);
    outputs(206) <= layer2_outputs(2088);
    outputs(207) <= (layer2_outputs(922)) xor (layer2_outputs(2976));
    outputs(208) <= not(layer2_outputs(3597));
    outputs(209) <= not(layer2_outputs(3578));
    outputs(210) <= (layer2_outputs(2847)) xor (layer2_outputs(3185));
    outputs(211) <= not(layer2_outputs(1275));
    outputs(212) <= not(layer2_outputs(1230));
    outputs(213) <= not(layer2_outputs(2428));
    outputs(214) <= not(layer2_outputs(47));
    outputs(215) <= layer2_outputs(1888);
    outputs(216) <= not((layer2_outputs(840)) xor (layer2_outputs(1419)));
    outputs(217) <= not(layer2_outputs(1460));
    outputs(218) <= not(layer2_outputs(1642));
    outputs(219) <= (layer2_outputs(3816)) and not (layer2_outputs(3204));
    outputs(220) <= layer2_outputs(4618);
    outputs(221) <= layer2_outputs(1340);
    outputs(222) <= not(layer2_outputs(1965)) or (layer2_outputs(4857));
    outputs(223) <= not(layer2_outputs(1493)) or (layer2_outputs(1546));
    outputs(224) <= layer2_outputs(3664);
    outputs(225) <= not(layer2_outputs(3346));
    outputs(226) <= not((layer2_outputs(4758)) xor (layer2_outputs(3334)));
    outputs(227) <= layer2_outputs(3806);
    outputs(228) <= layer2_outputs(2887);
    outputs(229) <= not((layer2_outputs(1139)) xor (layer2_outputs(390)));
    outputs(230) <= layer2_outputs(4802);
    outputs(231) <= layer2_outputs(906);
    outputs(232) <= not(layer2_outputs(4024));
    outputs(233) <= not(layer2_outputs(3260));
    outputs(234) <= not(layer2_outputs(2368));
    outputs(235) <= not(layer2_outputs(4723));
    outputs(236) <= not((layer2_outputs(5061)) and (layer2_outputs(3187)));
    outputs(237) <= not(layer2_outputs(3047));
    outputs(238) <= layer2_outputs(4519);
    outputs(239) <= (layer2_outputs(1542)) and not (layer2_outputs(1816));
    outputs(240) <= not(layer2_outputs(550));
    outputs(241) <= not(layer2_outputs(5018));
    outputs(242) <= not(layer2_outputs(4832));
    outputs(243) <= not(layer2_outputs(5117));
    outputs(244) <= not(layer2_outputs(3316));
    outputs(245) <= not(layer2_outputs(4325)) or (layer2_outputs(1615));
    outputs(246) <= not(layer2_outputs(4180));
    outputs(247) <= not(layer2_outputs(1562));
    outputs(248) <= (layer2_outputs(4310)) and not (layer2_outputs(2163));
    outputs(249) <= not(layer2_outputs(2855));
    outputs(250) <= not(layer2_outputs(2116));
    outputs(251) <= layer2_outputs(2002);
    outputs(252) <= not(layer2_outputs(955));
    outputs(253) <= layer2_outputs(606);
    outputs(254) <= layer2_outputs(1554);
    outputs(255) <= not(layer2_outputs(1206));
    outputs(256) <= layer2_outputs(2125);
    outputs(257) <= layer2_outputs(2863);
    outputs(258) <= (layer2_outputs(3690)) and (layer2_outputs(141));
    outputs(259) <= not(layer2_outputs(3980));
    outputs(260) <= layer2_outputs(2847);
    outputs(261) <= not((layer2_outputs(465)) xor (layer2_outputs(4842)));
    outputs(262) <= layer2_outputs(4799);
    outputs(263) <= layer2_outputs(3229);
    outputs(264) <= layer2_outputs(3877);
    outputs(265) <= not(layer2_outputs(163));
    outputs(266) <= layer2_outputs(1200);
    outputs(267) <= (layer2_outputs(2203)) xor (layer2_outputs(2950));
    outputs(268) <= layer2_outputs(1988);
    outputs(269) <= layer2_outputs(156);
    outputs(270) <= not(layer2_outputs(3728));
    outputs(271) <= (layer2_outputs(2985)) and not (layer2_outputs(4213));
    outputs(272) <= not(layer2_outputs(3441));
    outputs(273) <= not(layer2_outputs(1683));
    outputs(274) <= (layer2_outputs(3421)) and not (layer2_outputs(2142));
    outputs(275) <= not(layer2_outputs(1178));
    outputs(276) <= not(layer2_outputs(155));
    outputs(277) <= not(layer2_outputs(4148));
    outputs(278) <= layer2_outputs(3637);
    outputs(279) <= (layer2_outputs(4726)) xor (layer2_outputs(2187));
    outputs(280) <= layer2_outputs(4739);
    outputs(281) <= not(layer2_outputs(461));
    outputs(282) <= not((layer2_outputs(121)) xor (layer2_outputs(462)));
    outputs(283) <= layer2_outputs(953);
    outputs(284) <= layer2_outputs(2321);
    outputs(285) <= not(layer2_outputs(1685));
    outputs(286) <= not(layer2_outputs(3763));
    outputs(287) <= layer2_outputs(1994);
    outputs(288) <= layer2_outputs(2176);
    outputs(289) <= (layer2_outputs(256)) xor (layer2_outputs(2770));
    outputs(290) <= not(layer2_outputs(4202));
    outputs(291) <= '1';
    outputs(292) <= layer2_outputs(3900);
    outputs(293) <= not(layer2_outputs(2212));
    outputs(294) <= (layer2_outputs(280)) and (layer2_outputs(2771));
    outputs(295) <= (layer2_outputs(3502)) xor (layer2_outputs(700));
    outputs(296) <= not(layer2_outputs(2562));
    outputs(297) <= not(layer2_outputs(2744));
    outputs(298) <= layer2_outputs(2683);
    outputs(299) <= not((layer2_outputs(4016)) and (layer2_outputs(2642)));
    outputs(300) <= layer2_outputs(1287);
    outputs(301) <= layer2_outputs(2485);
    outputs(302) <= (layer2_outputs(2164)) xor (layer2_outputs(3743));
    outputs(303) <= layer2_outputs(543);
    outputs(304) <= layer2_outputs(4034);
    outputs(305) <= layer2_outputs(3677);
    outputs(306) <= layer2_outputs(13);
    outputs(307) <= layer2_outputs(2290);
    outputs(308) <= (layer2_outputs(2195)) and (layer2_outputs(228));
    outputs(309) <= layer2_outputs(2353);
    outputs(310) <= layer2_outputs(2706);
    outputs(311) <= not((layer2_outputs(227)) and (layer2_outputs(4601)));
    outputs(312) <= not(layer2_outputs(3319));
    outputs(313) <= not(layer2_outputs(5052));
    outputs(314) <= layer2_outputs(239);
    outputs(315) <= layer2_outputs(3274);
    outputs(316) <= (layer2_outputs(1751)) and not (layer2_outputs(2022));
    outputs(317) <= not(layer2_outputs(4101));
    outputs(318) <= not(layer2_outputs(3833));
    outputs(319) <= not(layer2_outputs(959));
    outputs(320) <= (layer2_outputs(1067)) or (layer2_outputs(1888));
    outputs(321) <= not((layer2_outputs(3719)) and (layer2_outputs(735)));
    outputs(322) <= not(layer2_outputs(1229));
    outputs(323) <= not((layer2_outputs(3588)) xor (layer2_outputs(4860)));
    outputs(324) <= not(layer2_outputs(1094));
    outputs(325) <= not((layer2_outputs(1160)) xor (layer2_outputs(587)));
    outputs(326) <= (layer2_outputs(314)) and not (layer2_outputs(1332));
    outputs(327) <= not(layer2_outputs(1621)) or (layer2_outputs(764));
    outputs(328) <= not(layer2_outputs(3037));
    outputs(329) <= (layer2_outputs(3398)) xor (layer2_outputs(4467));
    outputs(330) <= layer2_outputs(608);
    outputs(331) <= layer2_outputs(892);
    outputs(332) <= layer2_outputs(4722);
    outputs(333) <= layer2_outputs(2637);
    outputs(334) <= not(layer2_outputs(4851));
    outputs(335) <= not((layer2_outputs(2795)) xor (layer2_outputs(1160)));
    outputs(336) <= not(layer2_outputs(2413));
    outputs(337) <= not(layer2_outputs(1915));
    outputs(338) <= layer2_outputs(4938);
    outputs(339) <= layer2_outputs(644);
    outputs(340) <= not(layer2_outputs(4425)) or (layer2_outputs(1219));
    outputs(341) <= layer2_outputs(639);
    outputs(342) <= not(layer2_outputs(1999));
    outputs(343) <= not((layer2_outputs(4371)) and (layer2_outputs(943)));
    outputs(344) <= not(layer2_outputs(913)) or (layer2_outputs(4522));
    outputs(345) <= not(layer2_outputs(3525)) or (layer2_outputs(1950));
    outputs(346) <= layer2_outputs(3154);
    outputs(347) <= layer2_outputs(944);
    outputs(348) <= not(layer2_outputs(2456));
    outputs(349) <= not((layer2_outputs(1414)) xor (layer2_outputs(4909)));
    outputs(350) <= not(layer2_outputs(1584));
    outputs(351) <= layer2_outputs(3605);
    outputs(352) <= layer2_outputs(2818);
    outputs(353) <= not(layer2_outputs(1917));
    outputs(354) <= not((layer2_outputs(178)) and (layer2_outputs(3500)));
    outputs(355) <= not(layer2_outputs(4274));
    outputs(356) <= layer2_outputs(1530);
    outputs(357) <= (layer2_outputs(1434)) or (layer2_outputs(1073));
    outputs(358) <= layer2_outputs(2101);
    outputs(359) <= layer2_outputs(713);
    outputs(360) <= layer2_outputs(376);
    outputs(361) <= layer2_outputs(2754);
    outputs(362) <= layer2_outputs(1574);
    outputs(363) <= layer2_outputs(3819);
    outputs(364) <= not(layer2_outputs(69));
    outputs(365) <= not(layer2_outputs(726));
    outputs(366) <= layer2_outputs(1219);
    outputs(367) <= not(layer2_outputs(4716));
    outputs(368) <= not(layer2_outputs(1734)) or (layer2_outputs(2587));
    outputs(369) <= not(layer2_outputs(1953));
    outputs(370) <= not((layer2_outputs(3366)) xor (layer2_outputs(920)));
    outputs(371) <= not(layer2_outputs(70));
    outputs(372) <= layer2_outputs(730);
    outputs(373) <= not(layer2_outputs(2829)) or (layer2_outputs(291));
    outputs(374) <= not(layer2_outputs(3642));
    outputs(375) <= layer2_outputs(4176);
    outputs(376) <= not(layer2_outputs(3449));
    outputs(377) <= not((layer2_outputs(183)) xor (layer2_outputs(2015)));
    outputs(378) <= not((layer2_outputs(1015)) and (layer2_outputs(4966)));
    outputs(379) <= not(layer2_outputs(2442));
    outputs(380) <= layer2_outputs(1204);
    outputs(381) <= layer2_outputs(5112);
    outputs(382) <= not(layer2_outputs(4753));
    outputs(383) <= layer2_outputs(4761);
    outputs(384) <= not(layer2_outputs(3969)) or (layer2_outputs(4820));
    outputs(385) <= not((layer2_outputs(2613)) or (layer2_outputs(4659)));
    outputs(386) <= (layer2_outputs(1395)) and not (layer2_outputs(331));
    outputs(387) <= not(layer2_outputs(2206));
    outputs(388) <= (layer2_outputs(683)) xor (layer2_outputs(3464));
    outputs(389) <= (layer2_outputs(188)) and not (layer2_outputs(3572));
    outputs(390) <= layer2_outputs(1609);
    outputs(391) <= layer2_outputs(2050);
    outputs(392) <= (layer2_outputs(3988)) or (layer2_outputs(2190));
    outputs(393) <= layer2_outputs(2614);
    outputs(394) <= layer2_outputs(3821);
    outputs(395) <= not(layer2_outputs(4450));
    outputs(396) <= not((layer2_outputs(4272)) or (layer2_outputs(3456)));
    outputs(397) <= layer2_outputs(744);
    outputs(398) <= not(layer2_outputs(104));
    outputs(399) <= not(layer2_outputs(2319)) or (layer2_outputs(1657));
    outputs(400) <= layer2_outputs(567);
    outputs(401) <= layer2_outputs(4014);
    outputs(402) <= layer2_outputs(1066);
    outputs(403) <= not(layer2_outputs(4830));
    outputs(404) <= not(layer2_outputs(872));
    outputs(405) <= not(layer2_outputs(1798));
    outputs(406) <= not((layer2_outputs(3481)) and (layer2_outputs(4945)));
    outputs(407) <= not(layer2_outputs(1431));
    outputs(408) <= not(layer2_outputs(4252));
    outputs(409) <= not(layer2_outputs(697));
    outputs(410) <= layer2_outputs(4782);
    outputs(411) <= not(layer2_outputs(2065));
    outputs(412) <= (layer2_outputs(2620)) or (layer2_outputs(2535));
    outputs(413) <= not(layer2_outputs(3675));
    outputs(414) <= layer2_outputs(2601);
    outputs(415) <= layer2_outputs(1500);
    outputs(416) <= not(layer2_outputs(3037));
    outputs(417) <= layer2_outputs(2161);
    outputs(418) <= (layer2_outputs(1499)) or (layer2_outputs(2071));
    outputs(419) <= not(layer2_outputs(2079));
    outputs(420) <= layer2_outputs(4798);
    outputs(421) <= layer2_outputs(4434);
    outputs(422) <= not(layer2_outputs(4895));
    outputs(423) <= not(layer2_outputs(1347));
    outputs(424) <= not(layer2_outputs(3939));
    outputs(425) <= layer2_outputs(236);
    outputs(426) <= layer2_outputs(3538);
    outputs(427) <= layer2_outputs(3995);
    outputs(428) <= not(layer2_outputs(3583));
    outputs(429) <= not((layer2_outputs(232)) xor (layer2_outputs(3412)));
    outputs(430) <= not(layer2_outputs(4165));
    outputs(431) <= not(layer2_outputs(2305));
    outputs(432) <= not(layer2_outputs(1226)) or (layer2_outputs(1835));
    outputs(433) <= (layer2_outputs(3427)) or (layer2_outputs(209));
    outputs(434) <= layer2_outputs(957);
    outputs(435) <= layer2_outputs(101);
    outputs(436) <= layer2_outputs(582);
    outputs(437) <= (layer2_outputs(4142)) xor (layer2_outputs(1578));
    outputs(438) <= not(layer2_outputs(1650));
    outputs(439) <= layer2_outputs(986);
    outputs(440) <= not((layer2_outputs(1925)) xor (layer2_outputs(4007)));
    outputs(441) <= layer2_outputs(1495);
    outputs(442) <= layer2_outputs(1406);
    outputs(443) <= not(layer2_outputs(4528));
    outputs(444) <= layer2_outputs(660);
    outputs(445) <= not(layer2_outputs(1269));
    outputs(446) <= layer2_outputs(981);
    outputs(447) <= layer2_outputs(5072);
    outputs(448) <= (layer2_outputs(1034)) xor (layer2_outputs(4369));
    outputs(449) <= layer2_outputs(2209);
    outputs(450) <= not((layer2_outputs(3527)) xor (layer2_outputs(1539)));
    outputs(451) <= layer2_outputs(398);
    outputs(452) <= layer2_outputs(2276);
    outputs(453) <= not((layer2_outputs(989)) or (layer2_outputs(1134)));
    outputs(454) <= not(layer2_outputs(3735)) or (layer2_outputs(2704));
    outputs(455) <= (layer2_outputs(5039)) and not (layer2_outputs(2793));
    outputs(456) <= not(layer2_outputs(3085)) or (layer2_outputs(2054));
    outputs(457) <= (layer2_outputs(3138)) xor (layer2_outputs(3846));
    outputs(458) <= (layer2_outputs(1466)) xor (layer2_outputs(910));
    outputs(459) <= layer2_outputs(4362);
    outputs(460) <= layer2_outputs(529);
    outputs(461) <= not(layer2_outputs(3128));
    outputs(462) <= not(layer2_outputs(4073));
    outputs(463) <= not(layer2_outputs(3827));
    outputs(464) <= layer2_outputs(3497);
    outputs(465) <= not(layer2_outputs(904)) or (layer2_outputs(4030));
    outputs(466) <= layer2_outputs(2870);
    outputs(467) <= not((layer2_outputs(392)) or (layer2_outputs(107)));
    outputs(468) <= not(layer2_outputs(3042));
    outputs(469) <= not(layer2_outputs(4855));
    outputs(470) <= layer2_outputs(3474);
    outputs(471) <= not((layer2_outputs(2757)) xor (layer2_outputs(3848)));
    outputs(472) <= not(layer2_outputs(2695));
    outputs(473) <= not(layer2_outputs(954));
    outputs(474) <= not(layer2_outputs(690));
    outputs(475) <= layer2_outputs(3443);
    outputs(476) <= not(layer2_outputs(1217));
    outputs(477) <= layer2_outputs(2048);
    outputs(478) <= (layer2_outputs(2986)) and not (layer2_outputs(2007));
    outputs(479) <= not(layer2_outputs(464)) or (layer2_outputs(1118));
    outputs(480) <= not(layer2_outputs(264));
    outputs(481) <= layer2_outputs(2769);
    outputs(482) <= (layer2_outputs(1119)) and not (layer2_outputs(424));
    outputs(483) <= layer2_outputs(4019);
    outputs(484) <= layer2_outputs(2736);
    outputs(485) <= not(layer2_outputs(4842));
    outputs(486) <= not(layer2_outputs(2236));
    outputs(487) <= not(layer2_outputs(4395)) or (layer2_outputs(4755));
    outputs(488) <= layer2_outputs(591);
    outputs(489) <= layer2_outputs(4297);
    outputs(490) <= (layer2_outputs(209)) and not (layer2_outputs(565));
    outputs(491) <= not(layer2_outputs(3707));
    outputs(492) <= not(layer2_outputs(175));
    outputs(493) <= layer2_outputs(2588);
    outputs(494) <= not(layer2_outputs(3162));
    outputs(495) <= not(layer2_outputs(3196));
    outputs(496) <= (layer2_outputs(1228)) and not (layer2_outputs(4879));
    outputs(497) <= not((layer2_outputs(1007)) xor (layer2_outputs(4054)));
    outputs(498) <= layer2_outputs(5027);
    outputs(499) <= not(layer2_outputs(5064));
    outputs(500) <= not(layer2_outputs(1680));
    outputs(501) <= not(layer2_outputs(4808));
    outputs(502) <= not((layer2_outputs(1305)) or (layer2_outputs(4121)));
    outputs(503) <= not(layer2_outputs(1206));
    outputs(504) <= not(layer2_outputs(1351)) or (layer2_outputs(5066));
    outputs(505) <= layer2_outputs(235);
    outputs(506) <= (layer2_outputs(2958)) xor (layer2_outputs(3652));
    outputs(507) <= not(layer2_outputs(4171));
    outputs(508) <= (layer2_outputs(2713)) and (layer2_outputs(1066));
    outputs(509) <= not(layer2_outputs(2234));
    outputs(510) <= (layer2_outputs(1877)) and not (layer2_outputs(3430));
    outputs(511) <= (layer2_outputs(1228)) and not (layer2_outputs(2512));
    outputs(512) <= not((layer2_outputs(3494)) or (layer2_outputs(3958)));
    outputs(513) <= layer2_outputs(3303);
    outputs(514) <= (layer2_outputs(182)) and (layer2_outputs(932));
    outputs(515) <= not(layer2_outputs(1594));
    outputs(516) <= not(layer2_outputs(4817));
    outputs(517) <= layer2_outputs(4682);
    outputs(518) <= (layer2_outputs(2946)) and not (layer2_outputs(5102));
    outputs(519) <= (layer2_outputs(4162)) xor (layer2_outputs(2630));
    outputs(520) <= (layer2_outputs(2989)) and not (layer2_outputs(3396));
    outputs(521) <= layer2_outputs(3267);
    outputs(522) <= (layer2_outputs(4331)) and not (layer2_outputs(3932));
    outputs(523) <= not((layer2_outputs(2252)) or (layer2_outputs(4813)));
    outputs(524) <= layer2_outputs(417);
    outputs(525) <= layer2_outputs(5058);
    outputs(526) <= (layer2_outputs(153)) and not (layer2_outputs(2450));
    outputs(527) <= not(layer2_outputs(4247));
    outputs(528) <= (layer2_outputs(1266)) and (layer2_outputs(587));
    outputs(529) <= not(layer2_outputs(2108));
    outputs(530) <= (layer2_outputs(2889)) and not (layer2_outputs(1573));
    outputs(531) <= not((layer2_outputs(328)) or (layer2_outputs(2380)));
    outputs(532) <= '0';
    outputs(533) <= not(layer2_outputs(5108));
    outputs(534) <= layer2_outputs(2324);
    outputs(535) <= not((layer2_outputs(4930)) or (layer2_outputs(534)));
    outputs(536) <= not((layer2_outputs(1536)) xor (layer2_outputs(3792)));
    outputs(537) <= not((layer2_outputs(4234)) xor (layer2_outputs(876)));
    outputs(538) <= not(layer2_outputs(580));
    outputs(539) <= layer2_outputs(823);
    outputs(540) <= layer2_outputs(1729);
    outputs(541) <= not(layer2_outputs(778));
    outputs(542) <= not((layer2_outputs(4343)) and (layer2_outputs(1705)));
    outputs(543) <= not((layer2_outputs(4607)) xor (layer2_outputs(4480)));
    outputs(544) <= (layer2_outputs(1815)) and not (layer2_outputs(793));
    outputs(545) <= layer2_outputs(4993);
    outputs(546) <= (layer2_outputs(4431)) and not (layer2_outputs(3380));
    outputs(547) <= not((layer2_outputs(431)) or (layer2_outputs(1182)));
    outputs(548) <= not(layer2_outputs(835));
    outputs(549) <= not(layer2_outputs(729));
    outputs(550) <= not(layer2_outputs(5080));
    outputs(551) <= not((layer2_outputs(514)) or (layer2_outputs(4402)));
    outputs(552) <= not(layer2_outputs(4730));
    outputs(553) <= layer2_outputs(2774);
    outputs(554) <= not((layer2_outputs(651)) xor (layer2_outputs(3564)));
    outputs(555) <= layer2_outputs(2575);
    outputs(556) <= (layer2_outputs(116)) and not (layer2_outputs(5096));
    outputs(557) <= layer2_outputs(1172);
    outputs(558) <= (layer2_outputs(4859)) and not (layer2_outputs(1848));
    outputs(559) <= not((layer2_outputs(3946)) or (layer2_outputs(3347)));
    outputs(560) <= layer2_outputs(4053);
    outputs(561) <= not((layer2_outputs(493)) or (layer2_outputs(3494)));
    outputs(562) <= (layer2_outputs(3612)) and not (layer2_outputs(2601));
    outputs(563) <= not(layer2_outputs(3163));
    outputs(564) <= not(layer2_outputs(3674));
    outputs(565) <= (layer2_outputs(3151)) xor (layer2_outputs(2371));
    outputs(566) <= not(layer2_outputs(2262));
    outputs(567) <= (layer2_outputs(1844)) and not (layer2_outputs(352));
    outputs(568) <= (layer2_outputs(3605)) and not (layer2_outputs(4273));
    outputs(569) <= layer2_outputs(1345);
    outputs(570) <= layer2_outputs(4096);
    outputs(571) <= not(layer2_outputs(1135));
    outputs(572) <= (layer2_outputs(976)) xor (layer2_outputs(4032));
    outputs(573) <= (layer2_outputs(4949)) xor (layer2_outputs(3435));
    outputs(574) <= (layer2_outputs(2578)) and (layer2_outputs(1471));
    outputs(575) <= not((layer2_outputs(4748)) or (layer2_outputs(1274)));
    outputs(576) <= layer2_outputs(4885);
    outputs(577) <= (layer2_outputs(4632)) xor (layer2_outputs(2142));
    outputs(578) <= layer2_outputs(3782);
    outputs(579) <= not((layer2_outputs(904)) or (layer2_outputs(1818)));
    outputs(580) <= (layer2_outputs(3708)) and not (layer2_outputs(37));
    outputs(581) <= (layer2_outputs(3952)) and not (layer2_outputs(815));
    outputs(582) <= not((layer2_outputs(1864)) or (layer2_outputs(812)));
    outputs(583) <= layer2_outputs(4027);
    outputs(584) <= (layer2_outputs(4016)) and not (layer2_outputs(2310));
    outputs(585) <= not(layer2_outputs(3252));
    outputs(586) <= not((layer2_outputs(4136)) or (layer2_outputs(4687)));
    outputs(587) <= (layer2_outputs(2429)) and not (layer2_outputs(598));
    outputs(588) <= layer2_outputs(3580);
    outputs(589) <= not(layer2_outputs(4460));
    outputs(590) <= (layer2_outputs(1546)) and (layer2_outputs(1430));
    outputs(591) <= not((layer2_outputs(3081)) xor (layer2_outputs(5006)));
    outputs(592) <= not(layer2_outputs(1826));
    outputs(593) <= (layer2_outputs(886)) and not (layer2_outputs(3669));
    outputs(594) <= (layer2_outputs(2403)) and not (layer2_outputs(2695));
    outputs(595) <= (layer2_outputs(2297)) and (layer2_outputs(988));
    outputs(596) <= layer2_outputs(242);
    outputs(597) <= not((layer2_outputs(419)) or (layer2_outputs(933)));
    outputs(598) <= (layer2_outputs(1562)) and (layer2_outputs(1559));
    outputs(599) <= (layer2_outputs(2404)) and (layer2_outputs(4296));
    outputs(600) <= not(layer2_outputs(1747));
    outputs(601) <= layer2_outputs(3712);
    outputs(602) <= not(layer2_outputs(1231));
    outputs(603) <= layer2_outputs(1664);
    outputs(604) <= (layer2_outputs(2932)) and not (layer2_outputs(3387));
    outputs(605) <= not((layer2_outputs(4280)) or (layer2_outputs(3106)));
    outputs(606) <= not(layer2_outputs(219));
    outputs(607) <= layer2_outputs(4077);
    outputs(608) <= (layer2_outputs(4610)) and not (layer2_outputs(2827));
    outputs(609) <= layer2_outputs(2489);
    outputs(610) <= layer2_outputs(1180);
    outputs(611) <= (layer2_outputs(3970)) xor (layer2_outputs(3668));
    outputs(612) <= not(layer2_outputs(4609));
    outputs(613) <= layer2_outputs(3558);
    outputs(614) <= layer2_outputs(1843);
    outputs(615) <= (layer2_outputs(4746)) and (layer2_outputs(2240));
    outputs(616) <= (layer2_outputs(1978)) and not (layer2_outputs(3499));
    outputs(617) <= layer2_outputs(3243);
    outputs(618) <= layer2_outputs(5009);
    outputs(619) <= not(layer2_outputs(596));
    outputs(620) <= (layer2_outputs(3242)) and (layer2_outputs(3952));
    outputs(621) <= not(layer2_outputs(2743));
    outputs(622) <= not((layer2_outputs(2534)) or (layer2_outputs(2080)));
    outputs(623) <= not((layer2_outputs(2205)) or (layer2_outputs(2505)));
    outputs(624) <= (layer2_outputs(1386)) and not (layer2_outputs(410));
    outputs(625) <= not((layer2_outputs(2433)) or (layer2_outputs(1247)));
    outputs(626) <= not((layer2_outputs(2924)) or (layer2_outputs(2896)));
    outputs(627) <= not((layer2_outputs(3873)) or (layer2_outputs(3320)));
    outputs(628) <= not(layer2_outputs(3579));
    outputs(629) <= layer2_outputs(5072);
    outputs(630) <= (layer2_outputs(1324)) and not (layer2_outputs(746));
    outputs(631) <= layer2_outputs(4350);
    outputs(632) <= layer2_outputs(3861);
    outputs(633) <= layer2_outputs(4305);
    outputs(634) <= (layer2_outputs(3862)) and not (layer2_outputs(489));
    outputs(635) <= not(layer2_outputs(924));
    outputs(636) <= not((layer2_outputs(2474)) or (layer2_outputs(4905)));
    outputs(637) <= (layer2_outputs(2967)) and (layer2_outputs(1795));
    outputs(638) <= layer2_outputs(1222);
    outputs(639) <= layer2_outputs(2910);
    outputs(640) <= not(layer2_outputs(3961));
    outputs(641) <= (layer2_outputs(2053)) and not (layer2_outputs(1082));
    outputs(642) <= not(layer2_outputs(3169));
    outputs(643) <= layer2_outputs(2069);
    outputs(644) <= not((layer2_outputs(1876)) and (layer2_outputs(4396)));
    outputs(645) <= not((layer2_outputs(3948)) or (layer2_outputs(2492)));
    outputs(646) <= not((layer2_outputs(1817)) xor (layer2_outputs(3450)));
    outputs(647) <= not((layer2_outputs(1192)) or (layer2_outputs(4683)));
    outputs(648) <= layer2_outputs(4271);
    outputs(649) <= not(layer2_outputs(4927));
    outputs(650) <= (layer2_outputs(594)) and (layer2_outputs(3843));
    outputs(651) <= not(layer2_outputs(4724));
    outputs(652) <= layer2_outputs(3064);
    outputs(653) <= not(layer2_outputs(4774));
    outputs(654) <= (layer2_outputs(2478)) and not (layer2_outputs(1188));
    outputs(655) <= not(layer2_outputs(1247));
    outputs(656) <= (layer2_outputs(4729)) and (layer2_outputs(4839));
    outputs(657) <= not(layer2_outputs(1766));
    outputs(658) <= (layer2_outputs(1210)) and not (layer2_outputs(1468));
    outputs(659) <= not(layer2_outputs(1482));
    outputs(660) <= not((layer2_outputs(970)) or (layer2_outputs(1893)));
    outputs(661) <= layer2_outputs(4782);
    outputs(662) <= not(layer2_outputs(2521));
    outputs(663) <= layer2_outputs(4252);
    outputs(664) <= not((layer2_outputs(4441)) or (layer2_outputs(4723)));
    outputs(665) <= not(layer2_outputs(3001));
    outputs(666) <= (layer2_outputs(4158)) and not (layer2_outputs(1340));
    outputs(667) <= layer2_outputs(1590);
    outputs(668) <= (layer2_outputs(2902)) and not (layer2_outputs(2978));
    outputs(669) <= layer2_outputs(2038);
    outputs(670) <= (layer2_outputs(1784)) and not (layer2_outputs(512));
    outputs(671) <= layer2_outputs(2734);
    outputs(672) <= layer2_outputs(956);
    outputs(673) <= (layer2_outputs(516)) and not (layer2_outputs(2495));
    outputs(674) <= layer2_outputs(4277);
    outputs(675) <= (layer2_outputs(1108)) and not (layer2_outputs(401));
    outputs(676) <= not(layer2_outputs(3484));
    outputs(677) <= (layer2_outputs(115)) and not (layer2_outputs(4368));
    outputs(678) <= (layer2_outputs(1064)) and not (layer2_outputs(372));
    outputs(679) <= not((layer2_outputs(1035)) xor (layer2_outputs(4468)));
    outputs(680) <= not((layer2_outputs(2231)) or (layer2_outputs(2454)));
    outputs(681) <= (layer2_outputs(740)) or (layer2_outputs(273));
    outputs(682) <= (layer2_outputs(3193)) and not (layer2_outputs(4229));
    outputs(683) <= (layer2_outputs(1364)) or (layer2_outputs(4399));
    outputs(684) <= (layer2_outputs(4933)) and not (layer2_outputs(1585));
    outputs(685) <= (layer2_outputs(1680)) and (layer2_outputs(4578));
    outputs(686) <= not(layer2_outputs(3299));
    outputs(687) <= not(layer2_outputs(621));
    outputs(688) <= not(layer2_outputs(28)) or (layer2_outputs(169));
    outputs(689) <= layer2_outputs(20);
    outputs(690) <= not((layer2_outputs(3688)) xor (layer2_outputs(4725)));
    outputs(691) <= (layer2_outputs(2508)) and not (layer2_outputs(2012));
    outputs(692) <= not((layer2_outputs(4869)) xor (layer2_outputs(1896)));
    outputs(693) <= not(layer2_outputs(2510));
    outputs(694) <= not(layer2_outputs(410));
    outputs(695) <= layer2_outputs(4119);
    outputs(696) <= not(layer2_outputs(4481));
    outputs(697) <= not((layer2_outputs(4566)) or (layer2_outputs(1984)));
    outputs(698) <= not(layer2_outputs(2752));
    outputs(699) <= not(layer2_outputs(850));
    outputs(700) <= not(layer2_outputs(2616));
    outputs(701) <= not(layer2_outputs(3921));
    outputs(702) <= '0';
    outputs(703) <= layer2_outputs(4747);
    outputs(704) <= not((layer2_outputs(1958)) or (layer2_outputs(4215)));
    outputs(705) <= (layer2_outputs(4237)) and not (layer2_outputs(4407));
    outputs(706) <= not(layer2_outputs(4956));
    outputs(707) <= not(layer2_outputs(1020));
    outputs(708) <= not((layer2_outputs(3403)) and (layer2_outputs(5022)));
    outputs(709) <= (layer2_outputs(2592)) and not (layer2_outputs(2717));
    outputs(710) <= (layer2_outputs(5037)) and (layer2_outputs(4962));
    outputs(711) <= (layer2_outputs(990)) and (layer2_outputs(2919));
    outputs(712) <= (layer2_outputs(3438)) and not (layer2_outputs(910));
    outputs(713) <= layer2_outputs(248);
    outputs(714) <= (layer2_outputs(4015)) and (layer2_outputs(1832));
    outputs(715) <= not(layer2_outputs(4979));
    outputs(716) <= layer2_outputs(4258);
    outputs(717) <= (layer2_outputs(1945)) and (layer2_outputs(874));
    outputs(718) <= not(layer2_outputs(3506));
    outputs(719) <= not(layer2_outputs(2631));
    outputs(720) <= not((layer2_outputs(1934)) or (layer2_outputs(4382)));
    outputs(721) <= not(layer2_outputs(4926));
    outputs(722) <= not(layer2_outputs(3726));
    outputs(723) <= (layer2_outputs(826)) and not (layer2_outputs(1090));
    outputs(724) <= not((layer2_outputs(2444)) or (layer2_outputs(600)));
    outputs(725) <= not(layer2_outputs(3584));
    outputs(726) <= (layer2_outputs(4448)) and not (layer2_outputs(968));
    outputs(727) <= (layer2_outputs(3486)) and not (layer2_outputs(628));
    outputs(728) <= (layer2_outputs(1722)) and not (layer2_outputs(236));
    outputs(729) <= not((layer2_outputs(4451)) or (layer2_outputs(130)));
    outputs(730) <= not(layer2_outputs(3640));
    outputs(731) <= (layer2_outputs(2856)) xor (layer2_outputs(2905));
    outputs(732) <= layer2_outputs(1075);
    outputs(733) <= (layer2_outputs(3613)) and not (layer2_outputs(67));
    outputs(734) <= layer2_outputs(3769);
    outputs(735) <= not(layer2_outputs(3433));
    outputs(736) <= not((layer2_outputs(2450)) or (layer2_outputs(1349)));
    outputs(737) <= layer2_outputs(986);
    outputs(738) <= (layer2_outputs(686)) and not (layer2_outputs(3373));
    outputs(739) <= layer2_outputs(2264);
    outputs(740) <= (layer2_outputs(391)) and (layer2_outputs(4062));
    outputs(741) <= not(layer2_outputs(1979));
    outputs(742) <= layer2_outputs(3118);
    outputs(743) <= layer2_outputs(1360);
    outputs(744) <= layer2_outputs(4941);
    outputs(745) <= (layer2_outputs(926)) and not (layer2_outputs(365));
    outputs(746) <= (layer2_outputs(1444)) and not (layer2_outputs(2211));
    outputs(747) <= not(layer2_outputs(118)) or (layer2_outputs(4880));
    outputs(748) <= not(layer2_outputs(3893));
    outputs(749) <= (layer2_outputs(945)) xor (layer2_outputs(1759));
    outputs(750) <= (layer2_outputs(2727)) xor (layer2_outputs(4227));
    outputs(751) <= '0';
    outputs(752) <= not(layer2_outputs(343));
    outputs(753) <= (layer2_outputs(4919)) and (layer2_outputs(3369));
    outputs(754) <= not((layer2_outputs(2261)) or (layer2_outputs(1847)));
    outputs(755) <= layer2_outputs(4599);
    outputs(756) <= (layer2_outputs(994)) and (layer2_outputs(900));
    outputs(757) <= (layer2_outputs(3923)) and not (layer2_outputs(636));
    outputs(758) <= not(layer2_outputs(4847));
    outputs(759) <= not(layer2_outputs(1062));
    outputs(760) <= (layer2_outputs(184)) xor (layer2_outputs(3255));
    outputs(761) <= layer2_outputs(4173);
    outputs(762) <= layer2_outputs(4602);
    outputs(763) <= (layer2_outputs(4450)) or (layer2_outputs(2729));
    outputs(764) <= layer2_outputs(1881);
    outputs(765) <= not((layer2_outputs(3805)) or (layer2_outputs(4324)));
    outputs(766) <= not(layer2_outputs(2590)) or (layer2_outputs(3583));
    outputs(767) <= layer2_outputs(1011);
    outputs(768) <= not(layer2_outputs(3062)) or (layer2_outputs(4679));
    outputs(769) <= not((layer2_outputs(3812)) or (layer2_outputs(4488)));
    outputs(770) <= not(layer2_outputs(2040));
    outputs(771) <= (layer2_outputs(1709)) and not (layer2_outputs(272));
    outputs(772) <= not((layer2_outputs(4133)) xor (layer2_outputs(4500)));
    outputs(773) <= not((layer2_outputs(4398)) or (layer2_outputs(964)));
    outputs(774) <= (layer2_outputs(1773)) and (layer2_outputs(2747));
    outputs(775) <= (layer2_outputs(4072)) and (layer2_outputs(4886));
    outputs(776) <= (layer2_outputs(3638)) xor (layer2_outputs(3294));
    outputs(777) <= layer2_outputs(2091);
    outputs(778) <= (layer2_outputs(2351)) and (layer2_outputs(1225));
    outputs(779) <= not(layer2_outputs(2655));
    outputs(780) <= layer2_outputs(4823);
    outputs(781) <= layer2_outputs(2015);
    outputs(782) <= not((layer2_outputs(4299)) xor (layer2_outputs(518)));
    outputs(783) <= layer2_outputs(655);
    outputs(784) <= layer2_outputs(880);
    outputs(785) <= not((layer2_outputs(3589)) xor (layer2_outputs(3553)));
    outputs(786) <= (layer2_outputs(1939)) xor (layer2_outputs(1540));
    outputs(787) <= not(layer2_outputs(2144));
    outputs(788) <= not(layer2_outputs(4947));
    outputs(789) <= layer2_outputs(286);
    outputs(790) <= not(layer2_outputs(1740));
    outputs(791) <= layer2_outputs(1420);
    outputs(792) <= (layer2_outputs(3660)) xor (layer2_outputs(2970));
    outputs(793) <= layer2_outputs(2453);
    outputs(794) <= not((layer2_outputs(1169)) or (layer2_outputs(4094)));
    outputs(795) <= (layer2_outputs(1079)) and not (layer2_outputs(2010));
    outputs(796) <= (layer2_outputs(544)) and not (layer2_outputs(4884));
    outputs(797) <= (layer2_outputs(1868)) and (layer2_outputs(1443));
    outputs(798) <= (layer2_outputs(3254)) and (layer2_outputs(2585));
    outputs(799) <= (layer2_outputs(1439)) and (layer2_outputs(1150));
    outputs(800) <= not(layer2_outputs(1928));
    outputs(801) <= (layer2_outputs(3406)) and not (layer2_outputs(792));
    outputs(802) <= not(layer2_outputs(4900));
    outputs(803) <= (layer2_outputs(2273)) and not (layer2_outputs(1841));
    outputs(804) <= (layer2_outputs(4293)) and not (layer2_outputs(2361));
    outputs(805) <= (layer2_outputs(1942)) xor (layer2_outputs(3540));
    outputs(806) <= layer2_outputs(795);
    outputs(807) <= not(layer2_outputs(1598));
    outputs(808) <= layer2_outputs(3473);
    outputs(809) <= not(layer2_outputs(3875));
    outputs(810) <= not((layer2_outputs(1580)) or (layer2_outputs(3887)));
    outputs(811) <= (layer2_outputs(1717)) and (layer2_outputs(3789));
    outputs(812) <= layer2_outputs(2234);
    outputs(813) <= layer2_outputs(3660);
    outputs(814) <= not((layer2_outputs(3104)) or (layer2_outputs(2898)));
    outputs(815) <= (layer2_outputs(2780)) and not (layer2_outputs(4221));
    outputs(816) <= not(layer2_outputs(1911));
    outputs(817) <= '0';
    outputs(818) <= not(layer2_outputs(2526));
    outputs(819) <= (layer2_outputs(577)) xor (layer2_outputs(1589));
    outputs(820) <= (layer2_outputs(2487)) xor (layer2_outputs(820));
    outputs(821) <= not(layer2_outputs(2094));
    outputs(822) <= not(layer2_outputs(4177)) or (layer2_outputs(4700));
    outputs(823) <= (layer2_outputs(890)) and (layer2_outputs(1742));
    outputs(824) <= not((layer2_outputs(3501)) xor (layer2_outputs(2627)));
    outputs(825) <= layer2_outputs(5019);
    outputs(826) <= not(layer2_outputs(723));
    outputs(827) <= not((layer2_outputs(2061)) xor (layer2_outputs(1215)));
    outputs(828) <= not((layer2_outputs(4435)) or (layer2_outputs(2511)));
    outputs(829) <= not(layer2_outputs(4246));
    outputs(830) <= not(layer2_outputs(1171));
    outputs(831) <= not(layer2_outputs(2810));
    outputs(832) <= (layer2_outputs(1797)) xor (layer2_outputs(295));
    outputs(833) <= (layer2_outputs(1000)) and not (layer2_outputs(1074));
    outputs(834) <= (layer2_outputs(1527)) xor (layer2_outputs(3090));
    outputs(835) <= not(layer2_outputs(2803));
    outputs(836) <= not(layer2_outputs(1796));
    outputs(837) <= not(layer2_outputs(3201));
    outputs(838) <= (layer2_outputs(4159)) and not (layer2_outputs(4156));
    outputs(839) <= (layer2_outputs(1907)) and (layer2_outputs(1523));
    outputs(840) <= (layer2_outputs(3656)) xor (layer2_outputs(200));
    outputs(841) <= not(layer2_outputs(2373));
    outputs(842) <= not(layer2_outputs(1028));
    outputs(843) <= not((layer2_outputs(598)) or (layer2_outputs(1682)));
    outputs(844) <= (layer2_outputs(1924)) and (layer2_outputs(3611));
    outputs(845) <= layer2_outputs(1940);
    outputs(846) <= not(layer2_outputs(1363));
    outputs(847) <= (layer2_outputs(490)) xor (layer2_outputs(571));
    outputs(848) <= layer2_outputs(1344);
    outputs(849) <= not(layer2_outputs(1688));
    outputs(850) <= (layer2_outputs(2840)) and not (layer2_outputs(3984));
    outputs(851) <= (layer2_outputs(4179)) and (layer2_outputs(3838));
    outputs(852) <= not(layer2_outputs(1054));
    outputs(853) <= not((layer2_outputs(3745)) xor (layer2_outputs(3127)));
    outputs(854) <= not((layer2_outputs(2701)) xor (layer2_outputs(1997)));
    outputs(855) <= not((layer2_outputs(4656)) or (layer2_outputs(2567)));
    outputs(856) <= (layer2_outputs(3945)) and not (layer2_outputs(3057));
    outputs(857) <= not((layer2_outputs(1750)) or (layer2_outputs(2871)));
    outputs(858) <= (layer2_outputs(3051)) and (layer2_outputs(4576));
    outputs(859) <= (layer2_outputs(2385)) xor (layer2_outputs(4583));
    outputs(860) <= (layer2_outputs(2315)) and not (layer2_outputs(330));
    outputs(861) <= (layer2_outputs(2472)) and not (layer2_outputs(3858));
    outputs(862) <= (layer2_outputs(1905)) or (layer2_outputs(4118));
    outputs(863) <= not((layer2_outputs(3654)) or (layer2_outputs(3145)));
    outputs(864) <= (layer2_outputs(555)) and (layer2_outputs(3503));
    outputs(865) <= not(layer2_outputs(891));
    outputs(866) <= (layer2_outputs(4248)) xor (layer2_outputs(663));
    outputs(867) <= layer2_outputs(1326);
    outputs(868) <= (layer2_outputs(4258)) and not (layer2_outputs(4920));
    outputs(869) <= layer2_outputs(4558);
    outputs(870) <= not((layer2_outputs(843)) or (layer2_outputs(4455)));
    outputs(871) <= (layer2_outputs(1963)) and not (layer2_outputs(3377));
    outputs(872) <= not(layer2_outputs(716));
    outputs(873) <= (layer2_outputs(990)) and not (layer2_outputs(1772));
    outputs(874) <= not(layer2_outputs(2067));
    outputs(875) <= not(layer2_outputs(2625));
    outputs(876) <= (layer2_outputs(874)) and (layer2_outputs(5070));
    outputs(877) <= (layer2_outputs(1553)) and not (layer2_outputs(2835));
    outputs(878) <= not((layer2_outputs(1830)) or (layer2_outputs(3098)));
    outputs(879) <= not(layer2_outputs(191));
    outputs(880) <= not(layer2_outputs(1060));
    outputs(881) <= not(layer2_outputs(1657));
    outputs(882) <= not(layer2_outputs(2740));
    outputs(883) <= (layer2_outputs(8)) xor (layer2_outputs(4586));
    outputs(884) <= (layer2_outputs(4855)) xor (layer2_outputs(585));
    outputs(885) <= layer2_outputs(698);
    outputs(886) <= not((layer2_outputs(4397)) xor (layer2_outputs(3009)));
    outputs(887) <= not((layer2_outputs(2527)) xor (layer2_outputs(2779)));
    outputs(888) <= (layer2_outputs(305)) and (layer2_outputs(890));
    outputs(889) <= not(layer2_outputs(3487));
    outputs(890) <= not(layer2_outputs(3901)) or (layer2_outputs(882));
    outputs(891) <= (layer2_outputs(1443)) and not (layer2_outputs(2933));
    outputs(892) <= layer2_outputs(4717);
    outputs(893) <= (layer2_outputs(2041)) xor (layer2_outputs(2480));
    outputs(894) <= not(layer2_outputs(3737));
    outputs(895) <= not((layer2_outputs(4639)) or (layer2_outputs(2509)));
    outputs(896) <= not(layer2_outputs(3713));
    outputs(897) <= (layer2_outputs(3289)) xor (layer2_outputs(1520));
    outputs(898) <= not(layer2_outputs(1654));
    outputs(899) <= not((layer2_outputs(567)) or (layer2_outputs(4621)));
    outputs(900) <= not((layer2_outputs(682)) or (layer2_outputs(3415)));
    outputs(901) <= layer2_outputs(1158);
    outputs(902) <= (layer2_outputs(2190)) xor (layer2_outputs(1026));
    outputs(903) <= (layer2_outputs(3937)) and not (layer2_outputs(2724));
    outputs(904) <= (layer2_outputs(3878)) and (layer2_outputs(5015));
    outputs(905) <= layer2_outputs(2890);
    outputs(906) <= (layer2_outputs(4577)) and (layer2_outputs(4305));
    outputs(907) <= layer2_outputs(4065);
    outputs(908) <= not(layer2_outputs(641));
    outputs(909) <= layer2_outputs(262);
    outputs(910) <= not(layer2_outputs(4228));
    outputs(911) <= not((layer2_outputs(4055)) or (layer2_outputs(4080)));
    outputs(912) <= not((layer2_outputs(4702)) xor (layer2_outputs(4932)));
    outputs(913) <= not(layer2_outputs(3150));
    outputs(914) <= (layer2_outputs(3869)) and not (layer2_outputs(849));
    outputs(915) <= (layer2_outputs(51)) and not (layer2_outputs(511));
    outputs(916) <= not(layer2_outputs(3713));
    outputs(917) <= (layer2_outputs(193)) and not (layer2_outputs(604));
    outputs(918) <= layer2_outputs(612);
    outputs(919) <= not(layer2_outputs(3636));
    outputs(920) <= (layer2_outputs(1746)) xor (layer2_outputs(4816));
    outputs(921) <= (layer2_outputs(3295)) xor (layer2_outputs(1927));
    outputs(922) <= layer2_outputs(1872);
    outputs(923) <= not((layer2_outputs(2968)) or (layer2_outputs(3784)));
    outputs(924) <= not(layer2_outputs(1724));
    outputs(925) <= (layer2_outputs(1310)) and (layer2_outputs(456));
    outputs(926) <= (layer2_outputs(941)) and not (layer2_outputs(562));
    outputs(927) <= (layer2_outputs(3549)) and (layer2_outputs(242));
    outputs(928) <= layer2_outputs(1614);
    outputs(929) <= layer2_outputs(4292);
    outputs(930) <= (layer2_outputs(4815)) and (layer2_outputs(2735));
    outputs(931) <= not(layer2_outputs(3559));
    outputs(932) <= not((layer2_outputs(2621)) or (layer2_outputs(3828)));
    outputs(933) <= layer2_outputs(1963);
    outputs(934) <= not((layer2_outputs(2466)) or (layer2_outputs(4749)));
    outputs(935) <= not(layer2_outputs(2410));
    outputs(936) <= layer2_outputs(1827);
    outputs(937) <= (layer2_outputs(2239)) and not (layer2_outputs(4512));
    outputs(938) <= (layer2_outputs(3550)) and not (layer2_outputs(719));
    outputs(939) <= not(layer2_outputs(222));
    outputs(940) <= not(layer2_outputs(788));
    outputs(941) <= not(layer2_outputs(951)) or (layer2_outputs(4398));
    outputs(942) <= not(layer2_outputs(1604));
    outputs(943) <= not(layer2_outputs(4348));
    outputs(944) <= (layer2_outputs(2714)) and not (layer2_outputs(4134));
    outputs(945) <= layer2_outputs(1929);
    outputs(946) <= layer2_outputs(4279);
    outputs(947) <= layer2_outputs(1579);
    outputs(948) <= not(layer2_outputs(1130));
    outputs(949) <= (layer2_outputs(1096)) and not (layer2_outputs(1436));
    outputs(950) <= (layer2_outputs(4649)) xor (layer2_outputs(4865));
    outputs(951) <= not(layer2_outputs(484));
    outputs(952) <= (layer2_outputs(3991)) and not (layer2_outputs(485));
    outputs(953) <= not((layer2_outputs(1830)) or (layer2_outputs(2014)));
    outputs(954) <= (layer2_outputs(4818)) and not (layer2_outputs(2786));
    outputs(955) <= layer2_outputs(4644);
    outputs(956) <= layer2_outputs(3859);
    outputs(957) <= not(layer2_outputs(4631));
    outputs(958) <= (layer2_outputs(4891)) and not (layer2_outputs(4724));
    outputs(959) <= not((layer2_outputs(2108)) or (layer2_outputs(1758)));
    outputs(960) <= not(layer2_outputs(2599));
    outputs(961) <= not((layer2_outputs(566)) or (layer2_outputs(3654)));
    outputs(962) <= not((layer2_outputs(1338)) or (layer2_outputs(2458)));
    outputs(963) <= layer2_outputs(2149);
    outputs(964) <= not(layer2_outputs(1998));
    outputs(965) <= (layer2_outputs(2746)) xor (layer2_outputs(3344));
    outputs(966) <= (layer2_outputs(3033)) and not (layer2_outputs(537));
    outputs(967) <= layer2_outputs(4526);
    outputs(968) <= not(layer2_outputs(2374));
    outputs(969) <= not((layer2_outputs(83)) or (layer2_outputs(217)));
    outputs(970) <= layer2_outputs(711);
    outputs(971) <= not(layer2_outputs(2848));
    outputs(972) <= (layer2_outputs(4974)) and not (layer2_outputs(5116));
    outputs(973) <= layer2_outputs(4841);
    outputs(974) <= layer2_outputs(3609);
    outputs(975) <= not((layer2_outputs(3253)) or (layer2_outputs(1556)));
    outputs(976) <= (layer2_outputs(978)) xor (layer2_outputs(5087));
    outputs(977) <= (layer2_outputs(2788)) and (layer2_outputs(5032));
    outputs(978) <= (layer2_outputs(4766)) and not (layer2_outputs(4023));
    outputs(979) <= not(layer2_outputs(866));
    outputs(980) <= layer2_outputs(3280);
    outputs(981) <= (layer2_outputs(5011)) and not (layer2_outputs(2417));
    outputs(982) <= layer2_outputs(3989);
    outputs(983) <= layer2_outputs(2784);
    outputs(984) <= not(layer2_outputs(3014));
    outputs(985) <= layer2_outputs(647);
    outputs(986) <= layer2_outputs(1424);
    outputs(987) <= not(layer2_outputs(3233));
    outputs(988) <= layer2_outputs(91);
    outputs(989) <= (layer2_outputs(652)) and (layer2_outputs(1760));
    outputs(990) <= (layer2_outputs(4271)) and not (layer2_outputs(2948));
    outputs(991) <= not((layer2_outputs(3729)) or (layer2_outputs(4978)));
    outputs(992) <= (layer2_outputs(3842)) and not (layer2_outputs(1048));
    outputs(993) <= not(layer2_outputs(3470));
    outputs(994) <= (layer2_outputs(4548)) and not (layer2_outputs(1851));
    outputs(995) <= layer2_outputs(1729);
    outputs(996) <= (layer2_outputs(1807)) and not (layer2_outputs(553));
    outputs(997) <= not(layer2_outputs(1695));
    outputs(998) <= (layer2_outputs(3011)) xor (layer2_outputs(4475));
    outputs(999) <= (layer2_outputs(4886)) and (layer2_outputs(1259));
    outputs(1000) <= not(layer2_outputs(452));
    outputs(1001) <= layer2_outputs(1006);
    outputs(1002) <= layer2_outputs(5071);
    outputs(1003) <= not(layer2_outputs(4804));
    outputs(1004) <= not(layer2_outputs(1954));
    outputs(1005) <= (layer2_outputs(1467)) xor (layer2_outputs(5045));
    outputs(1006) <= layer2_outputs(177);
    outputs(1007) <= layer2_outputs(5048);
    outputs(1008) <= not(layer2_outputs(2551));
    outputs(1009) <= not(layer2_outputs(4902));
    outputs(1010) <= not(layer2_outputs(933));
    outputs(1011) <= layer2_outputs(2249);
    outputs(1012) <= not((layer2_outputs(1342)) or (layer2_outputs(4653)));
    outputs(1013) <= not((layer2_outputs(1520)) or (layer2_outputs(4939)));
    outputs(1014) <= not(layer2_outputs(3722));
    outputs(1015) <= not((layer2_outputs(344)) or (layer2_outputs(4783)));
    outputs(1016) <= layer2_outputs(2532);
    outputs(1017) <= (layer2_outputs(1894)) xor (layer2_outputs(1989));
    outputs(1018) <= not((layer2_outputs(5099)) or (layer2_outputs(2635)));
    outputs(1019) <= not(layer2_outputs(1946));
    outputs(1020) <= (layer2_outputs(150)) and not (layer2_outputs(3325));
    outputs(1021) <= layer2_outputs(2670);
    outputs(1022) <= (layer2_outputs(4819)) and not (layer2_outputs(4115));
    outputs(1023) <= layer2_outputs(3982);
    outputs(1024) <= (layer2_outputs(3981)) and not (layer2_outputs(381));
    outputs(1025) <= not(layer2_outputs(2213));
    outputs(1026) <= layer2_outputs(456);
    outputs(1027) <= not((layer2_outputs(3005)) xor (layer2_outputs(4730)));
    outputs(1028) <= not(layer2_outputs(2210));
    outputs(1029) <= not(layer2_outputs(4095));
    outputs(1030) <= layer2_outputs(4211);
    outputs(1031) <= layer2_outputs(347);
    outputs(1032) <= not(layer2_outputs(2550));
    outputs(1033) <= not(layer2_outputs(1530));
    outputs(1034) <= not(layer2_outputs(715));
    outputs(1035) <= not(layer2_outputs(4589)) or (layer2_outputs(2801));
    outputs(1036) <= not(layer2_outputs(3080)) or (layer2_outputs(679));
    outputs(1037) <= not(layer2_outputs(144));
    outputs(1038) <= not(layer2_outputs(664)) or (layer2_outputs(29));
    outputs(1039) <= layer2_outputs(2124);
    outputs(1040) <= (layer2_outputs(2430)) and not (layer2_outputs(442));
    outputs(1041) <= not((layer2_outputs(1968)) or (layer2_outputs(4540)));
    outputs(1042) <= not(layer2_outputs(3107));
    outputs(1043) <= not((layer2_outputs(4022)) xor (layer2_outputs(1597)));
    outputs(1044) <= not((layer2_outputs(3268)) xor (layer2_outputs(1992)));
    outputs(1045) <= layer2_outputs(3165);
    outputs(1046) <= not((layer2_outputs(1496)) or (layer2_outputs(887)));
    outputs(1047) <= not(layer2_outputs(1353));
    outputs(1048) <= layer2_outputs(4600);
    outputs(1049) <= (layer2_outputs(4137)) or (layer2_outputs(1462));
    outputs(1050) <= not(layer2_outputs(4319));
    outputs(1051) <= layer2_outputs(4489);
    outputs(1052) <= not(layer2_outputs(1269)) or (layer2_outputs(3063));
    outputs(1053) <= not(layer2_outputs(2025));
    outputs(1054) <= not(layer2_outputs(670));
    outputs(1055) <= not(layer2_outputs(3678));
    outputs(1056) <= (layer2_outputs(4752)) or (layer2_outputs(1450));
    outputs(1057) <= layer2_outputs(4051);
    outputs(1058) <= layer2_outputs(1585);
    outputs(1059) <= layer2_outputs(1700);
    outputs(1060) <= not((layer2_outputs(1981)) and (layer2_outputs(2115)));
    outputs(1061) <= layer2_outputs(431);
    outputs(1062) <= not(layer2_outputs(683));
    outputs(1063) <= not(layer2_outputs(2078));
    outputs(1064) <= layer2_outputs(3357);
    outputs(1065) <= layer2_outputs(2267);
    outputs(1066) <= not(layer2_outputs(535));
    outputs(1067) <= layer2_outputs(2686);
    outputs(1068) <= layer2_outputs(2445);
    outputs(1069) <= layer2_outputs(3832);
    outputs(1070) <= not(layer2_outputs(404)) or (layer2_outputs(1571));
    outputs(1071) <= (layer2_outputs(3823)) xor (layer2_outputs(685));
    outputs(1072) <= layer2_outputs(4999);
    outputs(1073) <= not(layer2_outputs(1861));
    outputs(1074) <= layer2_outputs(5085);
    outputs(1075) <= layer2_outputs(3401);
    outputs(1076) <= not((layer2_outputs(478)) xor (layer2_outputs(963)));
    outputs(1077) <= not(layer2_outputs(1163));
    outputs(1078) <= layer2_outputs(3115);
    outputs(1079) <= (layer2_outputs(4624)) and (layer2_outputs(3972));
    outputs(1080) <= layer2_outputs(3035);
    outputs(1081) <= layer2_outputs(3698);
    outputs(1082) <= not(layer2_outputs(4275));
    outputs(1083) <= not((layer2_outputs(849)) or (layer2_outputs(3917)));
    outputs(1084) <= layer2_outputs(3474);
    outputs(1085) <= (layer2_outputs(109)) xor (layer2_outputs(1415));
    outputs(1086) <= not((layer2_outputs(1306)) xor (layer2_outputs(2097)));
    outputs(1087) <= layer2_outputs(1606);
    outputs(1088) <= not(layer2_outputs(2518));
    outputs(1089) <= layer2_outputs(1346);
    outputs(1090) <= layer2_outputs(3811);
    outputs(1091) <= not(layer2_outputs(1324));
    outputs(1092) <= (layer2_outputs(1092)) or (layer2_outputs(3565));
    outputs(1093) <= (layer2_outputs(1581)) or (layer2_outputs(3288));
    outputs(1094) <= layer2_outputs(4488);
    outputs(1095) <= not((layer2_outputs(4814)) and (layer2_outputs(3214)));
    outputs(1096) <= not(layer2_outputs(1485));
    outputs(1097) <= not(layer2_outputs(4182));
    outputs(1098) <= layer2_outputs(1867);
    outputs(1099) <= not(layer2_outputs(2300));
    outputs(1100) <= not(layer2_outputs(1360)) or (layer2_outputs(4652));
    outputs(1101) <= not(layer2_outputs(3133));
    outputs(1102) <= layer2_outputs(1866);
    outputs(1103) <= layer2_outputs(2946);
    outputs(1104) <= (layer2_outputs(2775)) and (layer2_outputs(1301));
    outputs(1105) <= not(layer2_outputs(493));
    outputs(1106) <= not(layer2_outputs(3897));
    outputs(1107) <= (layer2_outputs(4775)) or (layer2_outputs(2579));
    outputs(1108) <= not(layer2_outputs(1914)) or (layer2_outputs(3965));
    outputs(1109) <= layer2_outputs(4991);
    outputs(1110) <= (layer2_outputs(2436)) or (layer2_outputs(1741));
    outputs(1111) <= (layer2_outputs(2060)) and not (layer2_outputs(4188));
    outputs(1112) <= layer2_outputs(3966);
    outputs(1113) <= not(layer2_outputs(472)) or (layer2_outputs(416));
    outputs(1114) <= not(layer2_outputs(4817));
    outputs(1115) <= not(layer2_outputs(2166));
    outputs(1116) <= not(layer2_outputs(2660));
    outputs(1117) <= (layer2_outputs(1891)) xor (layer2_outputs(4386));
    outputs(1118) <= layer2_outputs(4846);
    outputs(1119) <= not(layer2_outputs(253));
    outputs(1120) <= (layer2_outputs(2961)) xor (layer2_outputs(2524));
    outputs(1121) <= layer2_outputs(878);
    outputs(1122) <= not(layer2_outputs(689)) or (layer2_outputs(1733));
    outputs(1123) <= not(layer2_outputs(1005)) or (layer2_outputs(2995));
    outputs(1124) <= not(layer2_outputs(3323));
    outputs(1125) <= not(layer2_outputs(2176));
    outputs(1126) <= not(layer2_outputs(2328));
    outputs(1127) <= not(layer2_outputs(4268)) or (layer2_outputs(445));
    outputs(1128) <= not(layer2_outputs(5095)) or (layer2_outputs(3188));
    outputs(1129) <= (layer2_outputs(4688)) xor (layer2_outputs(2286));
    outputs(1130) <= not((layer2_outputs(4268)) and (layer2_outputs(1647)));
    outputs(1131) <= layer2_outputs(425);
    outputs(1132) <= layer2_outputs(2167);
    outputs(1133) <= layer2_outputs(95);
    outputs(1134) <= not((layer2_outputs(1754)) xor (layer2_outputs(3376)));
    outputs(1135) <= layer2_outputs(4179);
    outputs(1136) <= (layer2_outputs(539)) and (layer2_outputs(2693));
    outputs(1137) <= not(layer2_outputs(3455));
    outputs(1138) <= not(layer2_outputs(834));
    outputs(1139) <= not(layer2_outputs(2915));
    outputs(1140) <= not((layer2_outputs(1131)) xor (layer2_outputs(2245)));
    outputs(1141) <= (layer2_outputs(3125)) and not (layer2_outputs(2101));
    outputs(1142) <= layer2_outputs(4836);
    outputs(1143) <= not(layer2_outputs(751)) or (layer2_outputs(509));
    outputs(1144) <= not((layer2_outputs(4479)) xor (layer2_outputs(3245)));
    outputs(1145) <= (layer2_outputs(4742)) xor (layer2_outputs(589));
    outputs(1146) <= layer2_outputs(3270);
    outputs(1147) <= not((layer2_outputs(3697)) xor (layer2_outputs(138)));
    outputs(1148) <= not(layer2_outputs(2667));
    outputs(1149) <= (layer2_outputs(52)) and (layer2_outputs(3641));
    outputs(1150) <= (layer2_outputs(1456)) and (layer2_outputs(2711));
    outputs(1151) <= layer2_outputs(300);
    outputs(1152) <= layer2_outputs(181);
    outputs(1153) <= (layer2_outputs(3803)) or (layer2_outputs(4684));
    outputs(1154) <= not(layer2_outputs(2790));
    outputs(1155) <= not((layer2_outputs(8)) xor (layer2_outputs(2773)));
    outputs(1156) <= (layer2_outputs(2610)) and not (layer2_outputs(569));
    outputs(1157) <= not((layer2_outputs(3140)) xor (layer2_outputs(1404)));
    outputs(1158) <= not(layer2_outputs(2481));
    outputs(1159) <= not(layer2_outputs(149));
    outputs(1160) <= not((layer2_outputs(2791)) and (layer2_outputs(1475)));
    outputs(1161) <= not((layer2_outputs(3721)) xor (layer2_outputs(25)));
    outputs(1162) <= layer2_outputs(1016);
    outputs(1163) <= layer2_outputs(1455);
    outputs(1164) <= (layer2_outputs(4335)) xor (layer2_outputs(4487));
    outputs(1165) <= not(layer2_outputs(3248));
    outputs(1166) <= (layer2_outputs(2263)) xor (layer2_outputs(1622));
    outputs(1167) <= not(layer2_outputs(2337));
    outputs(1168) <= layer2_outputs(2018);
    outputs(1169) <= not(layer2_outputs(1611)) or (layer2_outputs(824));
    outputs(1170) <= not((layer2_outputs(1831)) or (layer2_outputs(3762)));
    outputs(1171) <= not(layer2_outputs(4911)) or (layer2_outputs(4862));
    outputs(1172) <= not(layer2_outputs(1382));
    outputs(1173) <= layer2_outputs(1132);
    outputs(1174) <= layer2_outputs(62);
    outputs(1175) <= not(layer2_outputs(2071));
    outputs(1176) <= layer2_outputs(2911);
    outputs(1177) <= not(layer2_outputs(2566));
    outputs(1178) <= not(layer2_outputs(4825));
    outputs(1179) <= not(layer2_outputs(666));
    outputs(1180) <= not(layer2_outputs(169));
    outputs(1181) <= not((layer2_outputs(1343)) xor (layer2_outputs(231)));
    outputs(1182) <= layer2_outputs(4741);
    outputs(1183) <= layer2_outputs(1828);
    outputs(1184) <= not(layer2_outputs(4606));
    outputs(1185) <= not(layer2_outputs(2062)) or (layer2_outputs(1976));
    outputs(1186) <= not(layer2_outputs(3871));
    outputs(1187) <= not(layer2_outputs(4290));
    outputs(1188) <= not(layer2_outputs(2090));
    outputs(1189) <= layer2_outputs(5082);
    outputs(1190) <= (layer2_outputs(739)) and not (layer2_outputs(3116));
    outputs(1191) <= not((layer2_outputs(4250)) and (layer2_outputs(233)));
    outputs(1192) <= not(layer2_outputs(662));
    outputs(1193) <= not((layer2_outputs(3365)) and (layer2_outputs(4509)));
    outputs(1194) <= layer2_outputs(1107);
    outputs(1195) <= not(layer2_outputs(2654));
    outputs(1196) <= not(layer2_outputs(1267));
    outputs(1197) <= not(layer2_outputs(4247));
    outputs(1198) <= not(layer2_outputs(4310));
    outputs(1199) <= (layer2_outputs(2838)) or (layer2_outputs(289));
    outputs(1200) <= (layer2_outputs(2544)) and (layer2_outputs(3907));
    outputs(1201) <= layer2_outputs(3362);
    outputs(1202) <= not((layer2_outputs(4779)) xor (layer2_outputs(4661)));
    outputs(1203) <= not(layer2_outputs(2056));
    outputs(1204) <= not((layer2_outputs(323)) xor (layer2_outputs(4313)));
    outputs(1205) <= not(layer2_outputs(2193));
    outputs(1206) <= layer2_outputs(4345);
    outputs(1207) <= not(layer2_outputs(2438));
    outputs(1208) <= layer2_outputs(1407);
    outputs(1209) <= (layer2_outputs(1780)) xor (layer2_outputs(4117));
    outputs(1210) <= layer2_outputs(790);
    outputs(1211) <= layer2_outputs(4704);
    outputs(1212) <= not(layer2_outputs(3958));
    outputs(1213) <= (layer2_outputs(3766)) and (layer2_outputs(1540));
    outputs(1214) <= not(layer2_outputs(342));
    outputs(1215) <= not(layer2_outputs(2913));
    outputs(1216) <= layer2_outputs(3532);
    outputs(1217) <= (layer2_outputs(838)) or (layer2_outputs(3322));
    outputs(1218) <= layer2_outputs(3682);
    outputs(1219) <= not(layer2_outputs(3626));
    outputs(1220) <= not((layer2_outputs(3835)) xor (layer2_outputs(3522)));
    outputs(1221) <= (layer2_outputs(2541)) and not (layer2_outputs(2332));
    outputs(1222) <= not(layer2_outputs(1869));
    outputs(1223) <= (layer2_outputs(4780)) and (layer2_outputs(3934));
    outputs(1224) <= '1';
    outputs(1225) <= (layer2_outputs(1183)) xor (layer2_outputs(2001));
    outputs(1226) <= (layer2_outputs(1398)) or (layer2_outputs(2080));
    outputs(1227) <= not(layer2_outputs(4942));
    outputs(1228) <= not((layer2_outputs(59)) and (layer2_outputs(2988)));
    outputs(1229) <= (layer2_outputs(1157)) xor (layer2_outputs(261));
    outputs(1230) <= layer2_outputs(1706);
    outputs(1231) <= layer2_outputs(2106);
    outputs(1232) <= not((layer2_outputs(4773)) xor (layer2_outputs(4596)));
    outputs(1233) <= layer2_outputs(4805);
    outputs(1234) <= not((layer2_outputs(3460)) xor (layer2_outputs(767)));
    outputs(1235) <= not((layer2_outputs(1239)) xor (layer2_outputs(4290)));
    outputs(1236) <= not(layer2_outputs(42)) or (layer2_outputs(1574));
    outputs(1237) <= (layer2_outputs(4102)) or (layer2_outputs(4691));
    outputs(1238) <= layer2_outputs(970);
    outputs(1239) <= not((layer2_outputs(3010)) xor (layer2_outputs(3516)));
    outputs(1240) <= layer2_outputs(977);
    outputs(1241) <= (layer2_outputs(2558)) or (layer2_outputs(1900));
    outputs(1242) <= not(layer2_outputs(1821));
    outputs(1243) <= (layer2_outputs(3321)) xor (layer2_outputs(4696));
    outputs(1244) <= (layer2_outputs(3038)) and (layer2_outputs(390));
    outputs(1245) <= not(layer2_outputs(2057));
    outputs(1246) <= not(layer2_outputs(4646));
    outputs(1247) <= not(layer2_outputs(3512));
    outputs(1248) <= not(layer2_outputs(4467));
    outputs(1249) <= not((layer2_outputs(710)) and (layer2_outputs(27)));
    outputs(1250) <= not((layer2_outputs(2738)) xor (layer2_outputs(2092)));
    outputs(1251) <= layer2_outputs(2469);
    outputs(1252) <= not(layer2_outputs(2712)) or (layer2_outputs(4492));
    outputs(1253) <= not(layer2_outputs(2143));
    outputs(1254) <= (layer2_outputs(2201)) and not (layer2_outputs(180));
    outputs(1255) <= not((layer2_outputs(2877)) or (layer2_outputs(294)));
    outputs(1256) <= layer2_outputs(28);
    outputs(1257) <= (layer2_outputs(382)) xor (layer2_outputs(1074));
    outputs(1258) <= not(layer2_outputs(2037)) or (layer2_outputs(4334));
    outputs(1259) <= layer2_outputs(3101);
    outputs(1260) <= layer2_outputs(1442);
    outputs(1261) <= layer2_outputs(4991);
    outputs(1262) <= not(layer2_outputs(2457));
    outputs(1263) <= not(layer2_outputs(4970));
    outputs(1264) <= not(layer2_outputs(3053));
    outputs(1265) <= not((layer2_outputs(4261)) xor (layer2_outputs(1294)));
    outputs(1266) <= layer2_outputs(1052);
    outputs(1267) <= (layer2_outputs(4635)) or (layer2_outputs(3826));
    outputs(1268) <= layer2_outputs(1157);
    outputs(1269) <= not(layer2_outputs(508));
    outputs(1270) <= layer2_outputs(2541);
    outputs(1271) <= layer2_outputs(3552);
    outputs(1272) <= (layer2_outputs(1560)) and not (layer2_outputs(1834));
    outputs(1273) <= layer2_outputs(2179);
    outputs(1274) <= (layer2_outputs(5041)) and not (layer2_outputs(5075));
    outputs(1275) <= not((layer2_outputs(3419)) or (layer2_outputs(2090)));
    outputs(1276) <= layer2_outputs(3690);
    outputs(1277) <= layer2_outputs(2484);
    outputs(1278) <= (layer2_outputs(4009)) and (layer2_outputs(2290));
    outputs(1279) <= layer2_outputs(3081);
    outputs(1280) <= not(layer2_outputs(4313));
    outputs(1281) <= layer2_outputs(4469);
    outputs(1282) <= layer2_outputs(2192);
    outputs(1283) <= (layer2_outputs(5098)) xor (layer2_outputs(2644));
    outputs(1284) <= layer2_outputs(4411);
    outputs(1285) <= not(layer2_outputs(3339));
    outputs(1286) <= not(layer2_outputs(3627));
    outputs(1287) <= layer2_outputs(4261);
    outputs(1288) <= not(layer2_outputs(3661)) or (layer2_outputs(708));
    outputs(1289) <= not(layer2_outputs(1452));
    outputs(1290) <= not(layer2_outputs(2647));
    outputs(1291) <= not(layer2_outputs(3046)) or (layer2_outputs(2513));
    outputs(1292) <= layer2_outputs(366);
    outputs(1293) <= not(layer2_outputs(976));
    outputs(1294) <= not(layer2_outputs(3656));
    outputs(1295) <= layer2_outputs(4099);
    outputs(1296) <= layer2_outputs(2047);
    outputs(1297) <= not(layer2_outputs(4293));
    outputs(1298) <= not(layer2_outputs(3457));
    outputs(1299) <= not(layer2_outputs(3296));
    outputs(1300) <= layer2_outputs(2253);
    outputs(1301) <= layer2_outputs(1910);
    outputs(1302) <= not(layer2_outputs(2756)) or (layer2_outputs(631));
    outputs(1303) <= not(layer2_outputs(210));
    outputs(1304) <= layer2_outputs(1725);
    outputs(1305) <= not(layer2_outputs(2665));
    outputs(1306) <= not(layer2_outputs(4876));
    outputs(1307) <= not(layer2_outputs(3508));
    outputs(1308) <= not(layer2_outputs(869));
    outputs(1309) <= not(layer2_outputs(3159));
    outputs(1310) <= layer2_outputs(3082);
    outputs(1311) <= not(layer2_outputs(3184));
    outputs(1312) <= layer2_outputs(677);
    outputs(1313) <= layer2_outputs(937);
    outputs(1314) <= not(layer2_outputs(4636));
    outputs(1315) <= not(layer2_outputs(4875));
    outputs(1316) <= '1';
    outputs(1317) <= not(layer2_outputs(3872));
    outputs(1318) <= layer2_outputs(534);
    outputs(1319) <= not(layer2_outputs(4721)) or (layer2_outputs(4379));
    outputs(1320) <= layer2_outputs(3728);
    outputs(1321) <= layer2_outputs(641);
    outputs(1322) <= not(layer2_outputs(2181));
    outputs(1323) <= not(layer2_outputs(2113));
    outputs(1324) <= layer2_outputs(75);
    outputs(1325) <= layer2_outputs(2468);
    outputs(1326) <= (layer2_outputs(0)) or (layer2_outputs(3890));
    outputs(1327) <= not(layer2_outputs(1613));
    outputs(1328) <= not(layer2_outputs(2635));
    outputs(1329) <= not(layer2_outputs(4568));
    outputs(1330) <= not(layer2_outputs(4553));
    outputs(1331) <= layer2_outputs(829);
    outputs(1332) <= not(layer2_outputs(3809));
    outputs(1333) <= not((layer2_outputs(3665)) or (layer2_outputs(3712)));
    outputs(1334) <= not(layer2_outputs(2137)) or (layer2_outputs(3947));
    outputs(1335) <= not(layer2_outputs(2113));
    outputs(1336) <= not((layer2_outputs(4520)) xor (layer2_outputs(592)));
    outputs(1337) <= not(layer2_outputs(1386));
    outputs(1338) <= layer2_outputs(4651);
    outputs(1339) <= (layer2_outputs(1435)) and (layer2_outputs(4472));
    outputs(1340) <= layer2_outputs(282);
    outputs(1341) <= not(layer2_outputs(1902));
    outputs(1342) <= layer2_outputs(2854);
    outputs(1343) <= not(layer2_outputs(2286)) or (layer2_outputs(2497));
    outputs(1344) <= layer2_outputs(2794);
    outputs(1345) <= not(layer2_outputs(4990));
    outputs(1346) <= not((layer2_outputs(4244)) xor (layer2_outputs(2352)));
    outputs(1347) <= layer2_outputs(151);
    outputs(1348) <= not(layer2_outputs(4892)) or (layer2_outputs(4278));
    outputs(1349) <= not(layer2_outputs(3122));
    outputs(1350) <= layer2_outputs(259);
    outputs(1351) <= (layer2_outputs(346)) and not (layer2_outputs(7));
    outputs(1352) <= not(layer2_outputs(3286));
    outputs(1353) <= layer2_outputs(2067);
    outputs(1354) <= not((layer2_outputs(830)) xor (layer2_outputs(3076)));
    outputs(1355) <= layer2_outputs(3148);
    outputs(1356) <= not(layer2_outputs(10));
    outputs(1357) <= not(layer2_outputs(2710)) or (layer2_outputs(4610));
    outputs(1358) <= not(layer2_outputs(4059)) or (layer2_outputs(249));
    outputs(1359) <= not(layer2_outputs(727));
    outputs(1360) <= layer2_outputs(2367);
    outputs(1361) <= (layer2_outputs(2339)) or (layer2_outputs(3467));
    outputs(1362) <= not(layer2_outputs(4996)) or (layer2_outputs(761));
    outputs(1363) <= not((layer2_outputs(1837)) xor (layer2_outputs(1926)));
    outputs(1364) <= layer2_outputs(1782);
    outputs(1365) <= not(layer2_outputs(4787));
    outputs(1366) <= not(layer2_outputs(319));
    outputs(1367) <= (layer2_outputs(1668)) xor (layer2_outputs(1515));
    outputs(1368) <= layer2_outputs(772);
    outputs(1369) <= layer2_outputs(2461);
    outputs(1370) <= not(layer2_outputs(796));
    outputs(1371) <= not(layer2_outputs(3416));
    outputs(1372) <= not(layer2_outputs(2011));
    outputs(1373) <= not(layer2_outputs(3523));
    outputs(1374) <= not(layer2_outputs(158));
    outputs(1375) <= (layer2_outputs(546)) and not (layer2_outputs(786));
    outputs(1376) <= not(layer2_outputs(1555));
    outputs(1377) <= not((layer2_outputs(3524)) and (layer2_outputs(238)));
    outputs(1378) <= not(layer2_outputs(1230));
    outputs(1379) <= (layer2_outputs(2709)) or (layer2_outputs(1780));
    outputs(1380) <= not((layer2_outputs(2334)) xor (layer2_outputs(2844)));
    outputs(1381) <= layer2_outputs(3453);
    outputs(1382) <= (layer2_outputs(4408)) xor (layer2_outputs(4122));
    outputs(1383) <= not(layer2_outputs(327));
    outputs(1384) <= not(layer2_outputs(918));
    outputs(1385) <= (layer2_outputs(1769)) xor (layer2_outputs(2117));
    outputs(1386) <= not(layer2_outputs(1393));
    outputs(1387) <= not(layer2_outputs(2780));
    outputs(1388) <= not(layer2_outputs(5119)) or (layer2_outputs(3982));
    outputs(1389) <= not((layer2_outputs(3268)) xor (layer2_outputs(4843)));
    outputs(1390) <= layer2_outputs(358);
    outputs(1391) <= not(layer2_outputs(1473)) or (layer2_outputs(4259));
    outputs(1392) <= (layer2_outputs(927)) xor (layer2_outputs(808));
    outputs(1393) <= not(layer2_outputs(1638)) or (layer2_outputs(5069));
    outputs(1394) <= (layer2_outputs(2805)) or (layer2_outputs(624));
    outputs(1395) <= layer2_outputs(2295);
    outputs(1396) <= not(layer2_outputs(3374));
    outputs(1397) <= not(layer2_outputs(701));
    outputs(1398) <= not((layer2_outputs(2078)) xor (layer2_outputs(4132)));
    outputs(1399) <= not(layer2_outputs(4642));
    outputs(1400) <= layer2_outputs(458);
    outputs(1401) <= not((layer2_outputs(830)) and (layer2_outputs(4822)));
    outputs(1402) <= not(layer2_outputs(2493));
    outputs(1403) <= not(layer2_outputs(3147)) or (layer2_outputs(2136));
    outputs(1404) <= not(layer2_outputs(2134));
    outputs(1405) <= layer2_outputs(3288);
    outputs(1406) <= (layer2_outputs(993)) or (layer2_outputs(2298));
    outputs(1407) <= layer2_outputs(4129);
    outputs(1408) <= not(layer2_outputs(1696));
    outputs(1409) <= not(layer2_outputs(1498));
    outputs(1410) <= layer2_outputs(864);
    outputs(1411) <= layer2_outputs(750);
    outputs(1412) <= layer2_outputs(2862);
    outputs(1413) <= not(layer2_outputs(1134));
    outputs(1414) <= not(layer2_outputs(4504));
    outputs(1415) <= (layer2_outputs(4779)) and (layer2_outputs(1889));
    outputs(1416) <= not(layer2_outputs(2335));
    outputs(1417) <= (layer2_outputs(4355)) xor (layer2_outputs(2891));
    outputs(1418) <= not(layer2_outputs(5006));
    outputs(1419) <= (layer2_outputs(515)) and (layer2_outputs(3181));
    outputs(1420) <= layer2_outputs(3896);
    outputs(1421) <= layer2_outputs(4992);
    outputs(1422) <= layer2_outputs(969);
    outputs(1423) <= (layer2_outputs(1505)) xor (layer2_outputs(2133));
    outputs(1424) <= not(layer2_outputs(3324));
    outputs(1425) <= not((layer2_outputs(646)) xor (layer2_outputs(1740)));
    outputs(1426) <= not((layer2_outputs(620)) and (layer2_outputs(92)));
    outputs(1427) <= (layer2_outputs(3913)) xor (layer2_outputs(3551));
    outputs(1428) <= layer2_outputs(4890);
    outputs(1429) <= not(layer2_outputs(2691));
    outputs(1430) <= not(layer2_outputs(658));
    outputs(1431) <= layer2_outputs(2969);
    outputs(1432) <= not(layer2_outputs(2670)) or (layer2_outputs(1746));
    outputs(1433) <= not((layer2_outputs(2892)) or (layer2_outputs(658)));
    outputs(1434) <= (layer2_outputs(2785)) and (layer2_outputs(1762));
    outputs(1435) <= not((layer2_outputs(3758)) xor (layer2_outputs(4088)));
    outputs(1436) <= (layer2_outputs(1111)) xor (layer2_outputs(3407));
    outputs(1437) <= layer2_outputs(4998);
    outputs(1438) <= layer2_outputs(1863);
    outputs(1439) <= layer2_outputs(3452);
    outputs(1440) <= not((layer2_outputs(2789)) and (layer2_outputs(1314)));
    outputs(1441) <= not(layer2_outputs(1796));
    outputs(1442) <= not((layer2_outputs(961)) and (layer2_outputs(1289)));
    outputs(1443) <= not(layer2_outputs(3954));
    outputs(1444) <= not(layer2_outputs(1136));
    outputs(1445) <= not(layer2_outputs(2169));
    outputs(1446) <= layer2_outputs(4481);
    outputs(1447) <= (layer2_outputs(2088)) xor (layer2_outputs(1302));
    outputs(1448) <= not(layer2_outputs(2344));
    outputs(1449) <= not(layer2_outputs(4642)) or (layer2_outputs(2497));
    outputs(1450) <= not(layer2_outputs(1840));
    outputs(1451) <= not(layer2_outputs(1914));
    outputs(1452) <= not(layer2_outputs(3304));
    outputs(1453) <= not(layer2_outputs(115));
    outputs(1454) <= not(layer2_outputs(2215));
    outputs(1455) <= layer2_outputs(5078);
    outputs(1456) <= (layer2_outputs(903)) and not (layer2_outputs(4168));
    outputs(1457) <= not(layer2_outputs(500)) or (layer2_outputs(2262));
    outputs(1458) <= (layer2_outputs(4241)) and not (layer2_outputs(814));
    outputs(1459) <= layer2_outputs(4300);
    outputs(1460) <= layer2_outputs(4639);
    outputs(1461) <= layer2_outputs(3135);
    outputs(1462) <= not(layer2_outputs(1871));
    outputs(1463) <= layer2_outputs(782);
    outputs(1464) <= layer2_outputs(2969);
    outputs(1465) <= layer2_outputs(2236);
    outputs(1466) <= not((layer2_outputs(1350)) xor (layer2_outputs(2482)));
    outputs(1467) <= layer2_outputs(4896);
    outputs(1468) <= (layer2_outputs(1240)) and not (layer2_outputs(1391));
    outputs(1469) <= not(layer2_outputs(3607));
    outputs(1470) <= layer2_outputs(3161);
    outputs(1471) <= not(layer2_outputs(3759));
    outputs(1472) <= layer2_outputs(1759);
    outputs(1473) <= not(layer2_outputs(3595));
    outputs(1474) <= not(layer2_outputs(2202));
    outputs(1475) <= layer2_outputs(1670);
    outputs(1476) <= layer2_outputs(4492);
    outputs(1477) <= layer2_outputs(4375);
    outputs(1478) <= layer2_outputs(1856);
    outputs(1479) <= not(layer2_outputs(2379)) or (layer2_outputs(3229));
    outputs(1480) <= (layer2_outputs(1989)) xor (layer2_outputs(2153));
    outputs(1481) <= layer2_outputs(1235);
    outputs(1482) <= layer2_outputs(269);
    outputs(1483) <= layer2_outputs(2370);
    outputs(1484) <= (layer2_outputs(1752)) and (layer2_outputs(1018));
    outputs(1485) <= layer2_outputs(147);
    outputs(1486) <= not(layer2_outputs(3189)) or (layer2_outputs(1758));
    outputs(1487) <= not(layer2_outputs(1185));
    outputs(1488) <= not(layer2_outputs(4135));
    outputs(1489) <= not(layer2_outputs(3831));
    outputs(1490) <= not(layer2_outputs(3559));
    outputs(1491) <= (layer2_outputs(4580)) and not (layer2_outputs(1327));
    outputs(1492) <= layer2_outputs(4484);
    outputs(1493) <= layer2_outputs(127);
    outputs(1494) <= layer2_outputs(4073);
    outputs(1495) <= not(layer2_outputs(2319));
    outputs(1496) <= (layer2_outputs(2980)) or (layer2_outputs(1552));
    outputs(1497) <= not(layer2_outputs(2076));
    outputs(1498) <= layer2_outputs(3019);
    outputs(1499) <= layer2_outputs(3412);
    outputs(1500) <= layer2_outputs(4901);
    outputs(1501) <= layer2_outputs(1058);
    outputs(1502) <= layer2_outputs(2022);
    outputs(1503) <= (layer2_outputs(2757)) or (layer2_outputs(4257));
    outputs(1504) <= not(layer2_outputs(4172));
    outputs(1505) <= not(layer2_outputs(1337));
    outputs(1506) <= (layer2_outputs(1921)) and not (layer2_outputs(1964));
    outputs(1507) <= layer2_outputs(2800);
    outputs(1508) <= layer2_outputs(2715);
    outputs(1509) <= (layer2_outputs(66)) and not (layer2_outputs(2315));
    outputs(1510) <= (layer2_outputs(3689)) or (layer2_outputs(3881));
    outputs(1511) <= layer2_outputs(2911);
    outputs(1512) <= layer2_outputs(636);
    outputs(1513) <= not(layer2_outputs(2405));
    outputs(1514) <= not(layer2_outputs(70));
    outputs(1515) <= (layer2_outputs(1019)) and not (layer2_outputs(4275));
    outputs(1516) <= (layer2_outputs(3047)) and not (layer2_outputs(3825));
    outputs(1517) <= not(layer2_outputs(3578));
    outputs(1518) <= layer2_outputs(3830);
    outputs(1519) <= not(layer2_outputs(4037));
    outputs(1520) <= not(layer2_outputs(469)) or (layer2_outputs(457));
    outputs(1521) <= layer2_outputs(572);
    outputs(1522) <= not(layer2_outputs(715));
    outputs(1523) <= not(layer2_outputs(694));
    outputs(1524) <= layer2_outputs(4502);
    outputs(1525) <= not(layer2_outputs(3313)) or (layer2_outputs(1154));
    outputs(1526) <= layer2_outputs(125);
    outputs(1527) <= layer2_outputs(4415);
    outputs(1528) <= (layer2_outputs(4482)) and (layer2_outputs(3219));
    outputs(1529) <= not(layer2_outputs(2692)) or (layer2_outputs(281));
    outputs(1530) <= not((layer2_outputs(4920)) xor (layer2_outputs(4946)));
    outputs(1531) <= layer2_outputs(3049);
    outputs(1532) <= (layer2_outputs(167)) and not (layer2_outputs(3134));
    outputs(1533) <= (layer2_outputs(4428)) or (layer2_outputs(5002));
    outputs(1534) <= not(layer2_outputs(3072));
    outputs(1535) <= (layer2_outputs(184)) and (layer2_outputs(4283));
    outputs(1536) <= not((layer2_outputs(4929)) xor (layer2_outputs(1189)));
    outputs(1537) <= not(layer2_outputs(4321)) or (layer2_outputs(575));
    outputs(1538) <= not(layer2_outputs(3548));
    outputs(1539) <= layer2_outputs(2865);
    outputs(1540) <= not(layer2_outputs(4711));
    outputs(1541) <= not(layer2_outputs(3174));
    outputs(1542) <= layer2_outputs(3052);
    outputs(1543) <= not(layer2_outputs(2350));
    outputs(1544) <= not(layer2_outputs(137));
    outputs(1545) <= layer2_outputs(4607);
    outputs(1546) <= not(layer2_outputs(1235));
    outputs(1547) <= (layer2_outputs(784)) xor (layer2_outputs(4383));
    outputs(1548) <= (layer2_outputs(4839)) and not (layer2_outputs(4235));
    outputs(1549) <= layer2_outputs(4120);
    outputs(1550) <= layer2_outputs(2851);
    outputs(1551) <= not(layer2_outputs(4289));
    outputs(1552) <= not((layer2_outputs(1774)) and (layer2_outputs(853)));
    outputs(1553) <= (layer2_outputs(460)) and not (layer2_outputs(4549));
    outputs(1554) <= (layer2_outputs(3429)) and not (layer2_outputs(673));
    outputs(1555) <= (layer2_outputs(1284)) and not (layer2_outputs(105));
    outputs(1556) <= not(layer2_outputs(1006));
    outputs(1557) <= not(layer2_outputs(1655));
    outputs(1558) <= (layer2_outputs(4248)) and not (layer2_outputs(1524));
    outputs(1559) <= (layer2_outputs(352)) and (layer2_outputs(1743));
    outputs(1560) <= (layer2_outputs(4827)) and not (layer2_outputs(1098));
    outputs(1561) <= layer2_outputs(4810);
    outputs(1562) <= (layer2_outputs(3836)) xor (layer2_outputs(884));
    outputs(1563) <= layer2_outputs(2540);
    outputs(1564) <= layer2_outputs(908);
    outputs(1565) <= layer2_outputs(2242);
    outputs(1566) <= not(layer2_outputs(656)) or (layer2_outputs(4303));
    outputs(1567) <= not((layer2_outputs(126)) xor (layer2_outputs(2477)));
    outputs(1568) <= (layer2_outputs(2701)) and (layer2_outputs(4863));
    outputs(1569) <= not(layer2_outputs(3643));
    outputs(1570) <= layer2_outputs(2348);
    outputs(1571) <= layer2_outputs(537);
    outputs(1572) <= (layer2_outputs(1704)) and (layer2_outputs(100));
    outputs(1573) <= not(layer2_outputs(4539));
    outputs(1574) <= not(layer2_outputs(1954));
    outputs(1575) <= not((layer2_outputs(143)) xor (layer2_outputs(4957)));
    outputs(1576) <= not(layer2_outputs(841));
    outputs(1577) <= (layer2_outputs(4460)) and not (layer2_outputs(4447));
    outputs(1578) <= not(layer2_outputs(1167));
    outputs(1579) <= layer2_outputs(3329);
    outputs(1580) <= (layer2_outputs(873)) and not (layer2_outputs(5117));
    outputs(1581) <= layer2_outputs(287);
    outputs(1582) <= not((layer2_outputs(368)) and (layer2_outputs(1961)));
    outputs(1583) <= not(layer2_outputs(3177));
    outputs(1584) <= not(layer2_outputs(2889));
    outputs(1585) <= layer2_outputs(3649);
    outputs(1586) <= (layer2_outputs(2607)) or (layer2_outputs(4474));
    outputs(1587) <= not(layer2_outputs(2160));
    outputs(1588) <= not(layer2_outputs(471));
    outputs(1589) <= (layer2_outputs(3442)) xor (layer2_outputs(3744));
    outputs(1590) <= not((layer2_outputs(4834)) or (layer2_outputs(2594)));
    outputs(1591) <= not((layer2_outputs(2926)) and (layer2_outputs(1698)));
    outputs(1592) <= (layer2_outputs(1820)) or (layer2_outputs(2032));
    outputs(1593) <= not(layer2_outputs(1557));
    outputs(1594) <= layer2_outputs(758);
    outputs(1595) <= not((layer2_outputs(1025)) xor (layer2_outputs(2621)));
    outputs(1596) <= (layer2_outputs(4153)) xor (layer2_outputs(1401));
    outputs(1597) <= layer2_outputs(4716);
    outputs(1598) <= (layer2_outputs(2434)) and (layer2_outputs(1200));
    outputs(1599) <= layer2_outputs(239);
    outputs(1600) <= not(layer2_outputs(190));
    outputs(1601) <= (layer2_outputs(1081)) and not (layer2_outputs(2806));
    outputs(1602) <= not(layer2_outputs(2514));
    outputs(1603) <= layer2_outputs(1009);
    outputs(1604) <= not(layer2_outputs(395));
    outputs(1605) <= (layer2_outputs(3353)) and not (layer2_outputs(2983));
    outputs(1606) <= not((layer2_outputs(2312)) xor (layer2_outputs(3470)));
    outputs(1607) <= layer2_outputs(1439);
    outputs(1608) <= layer2_outputs(4987);
    outputs(1609) <= layer2_outputs(1016);
    outputs(1610) <= layer2_outputs(2571);
    outputs(1611) <= not(layer2_outputs(1174));
    outputs(1612) <= layer2_outputs(832);
    outputs(1613) <= layer2_outputs(1892);
    outputs(1614) <= (layer2_outputs(356)) and not (layer2_outputs(936));
    outputs(1615) <= not(layer2_outputs(4504));
    outputs(1616) <= layer2_outputs(4449);
    outputs(1617) <= layer2_outputs(1722);
    outputs(1618) <= (layer2_outputs(2441)) xor (layer2_outputs(4705));
    outputs(1619) <= not(layer2_outputs(4997)) or (layer2_outputs(2000));
    outputs(1620) <= not(layer2_outputs(1751));
    outputs(1621) <= (layer2_outputs(1292)) and not (layer2_outputs(4352));
    outputs(1622) <= layer2_outputs(1263);
    outputs(1623) <= not(layer2_outputs(4065));
    outputs(1624) <= layer2_outputs(735);
    outputs(1625) <= not((layer2_outputs(2269)) xor (layer2_outputs(68)));
    outputs(1626) <= layer2_outputs(3518);
    outputs(1627) <= layer2_outputs(3348);
    outputs(1628) <= not((layer2_outputs(4365)) or (layer2_outputs(1845)));
    outputs(1629) <= not(layer2_outputs(3783));
    outputs(1630) <= not(layer2_outputs(275));
    outputs(1631) <= not(layer2_outputs(3194));
    outputs(1632) <= layer2_outputs(3093);
    outputs(1633) <= '1';
    outputs(1634) <= (layer2_outputs(21)) or (layer2_outputs(29));
    outputs(1635) <= layer2_outputs(724);
    outputs(1636) <= not(layer2_outputs(1684));
    outputs(1637) <= layer2_outputs(1290);
    outputs(1638) <= layer2_outputs(3415);
    outputs(1639) <= layer2_outputs(2018);
    outputs(1640) <= (layer2_outputs(645)) xor (layer2_outputs(3208));
    outputs(1641) <= not(layer2_outputs(3593));
    outputs(1642) <= layer2_outputs(684);
    outputs(1643) <= not(layer2_outputs(1825)) or (layer2_outputs(1803));
    outputs(1644) <= (layer2_outputs(4028)) and (layer2_outputs(532));
    outputs(1645) <= (layer2_outputs(3176)) xor (layer2_outputs(4474));
    outputs(1646) <= not(layer2_outputs(4199));
    outputs(1647) <= layer2_outputs(2360);
    outputs(1648) <= layer2_outputs(2965);
    outputs(1649) <= not(layer2_outputs(4155));
    outputs(1650) <= not(layer2_outputs(3356));
    outputs(1651) <= not(layer2_outputs(787));
    outputs(1652) <= not(layer2_outputs(2231)) or (layer2_outputs(311));
    outputs(1653) <= layer2_outputs(5092);
    outputs(1654) <= not(layer2_outputs(1566));
    outputs(1655) <= layer2_outputs(2819);
    outputs(1656) <= layer2_outputs(2288);
    outputs(1657) <= layer2_outputs(1488);
    outputs(1658) <= (layer2_outputs(3283)) and not (layer2_outputs(419));
    outputs(1659) <= layer2_outputs(1588);
    outputs(1660) <= not(layer2_outputs(3242));
    outputs(1661) <= not(layer2_outputs(371));
    outputs(1662) <= (layer2_outputs(3655)) xor (layer2_outputs(2405));
    outputs(1663) <= (layer2_outputs(3337)) xor (layer2_outputs(1331));
    outputs(1664) <= layer2_outputs(11);
    outputs(1665) <= layer2_outputs(3315);
    outputs(1666) <= layer2_outputs(5107);
    outputs(1667) <= (layer2_outputs(2146)) and not (layer2_outputs(4562));
    outputs(1668) <= layer2_outputs(4237);
    outputs(1669) <= layer2_outputs(2679);
    outputs(1670) <= layer2_outputs(3813);
    outputs(1671) <= (layer2_outputs(2083)) or (layer2_outputs(6));
    outputs(1672) <= not(layer2_outputs(2443));
    outputs(1673) <= layer2_outputs(277);
    outputs(1674) <= not(layer2_outputs(1291));
    outputs(1675) <= (layer2_outputs(1292)) and (layer2_outputs(3109));
    outputs(1676) <= not((layer2_outputs(18)) or (layer2_outputs(1901)));
    outputs(1677) <= not(layer2_outputs(491));
    outputs(1678) <= not((layer2_outputs(1919)) or (layer2_outputs(437)));
    outputs(1679) <= not(layer2_outputs(2954)) or (layer2_outputs(4925));
    outputs(1680) <= not(layer2_outputs(4669)) or (layer2_outputs(4898));
    outputs(1681) <= (layer2_outputs(3896)) and (layer2_outputs(280));
    outputs(1682) <= layer2_outputs(422);
    outputs(1683) <= (layer2_outputs(1393)) xor (layer2_outputs(3691));
    outputs(1684) <= not((layer2_outputs(3623)) or (layer2_outputs(3418)));
    outputs(1685) <= layer2_outputs(724);
    outputs(1686) <= not(layer2_outputs(1239));
    outputs(1687) <= not((layer2_outputs(2741)) or (layer2_outputs(2438)));
    outputs(1688) <= not(layer2_outputs(1196));
    outputs(1689) <= layer2_outputs(4452);
    outputs(1690) <= layer2_outputs(3176);
    outputs(1691) <= (layer2_outputs(2922)) and (layer2_outputs(3408));
    outputs(1692) <= not(layer2_outputs(4253));
    outputs(1693) <= not(layer2_outputs(4314));
    outputs(1694) <= (layer2_outputs(1770)) and (layer2_outputs(1312));
    outputs(1695) <= layer2_outputs(3018);
    outputs(1696) <= not((layer2_outputs(2935)) xor (layer2_outputs(4823)));
    outputs(1697) <= not((layer2_outputs(3439)) or (layer2_outputs(4118)));
    outputs(1698) <= not(layer2_outputs(270));
    outputs(1699) <= layer2_outputs(3584);
    outputs(1700) <= not((layer2_outputs(1885)) xor (layer2_outputs(2917)));
    outputs(1701) <= not(layer2_outputs(4332));
    outputs(1702) <= layer2_outputs(1430);
    outputs(1703) <= layer2_outputs(3923);
    outputs(1704) <= layer2_outputs(602);
    outputs(1705) <= layer2_outputs(2330);
    outputs(1706) <= layer2_outputs(32);
    outputs(1707) <= not(layer2_outputs(4391));
    outputs(1708) <= not(layer2_outputs(3657));
    outputs(1709) <= not(layer2_outputs(4035));
    outputs(1710) <= not(layer2_outputs(4737));
    outputs(1711) <= layer2_outputs(847);
    outputs(1712) <= layer2_outputs(602);
    outputs(1713) <= not((layer2_outputs(1965)) and (layer2_outputs(3264)));
    outputs(1714) <= not(layer2_outputs(5039));
    outputs(1715) <= (layer2_outputs(637)) or (layer2_outputs(4664));
    outputs(1716) <= (layer2_outputs(1757)) xor (layer2_outputs(179));
    outputs(1717) <= layer2_outputs(1599);
    outputs(1718) <= (layer2_outputs(526)) and not (layer2_outputs(4605));
    outputs(1719) <= not(layer2_outputs(4008));
    outputs(1720) <= (layer2_outputs(1629)) xor (layer2_outputs(4236));
    outputs(1721) <= not(layer2_outputs(2309)) or (layer2_outputs(1136));
    outputs(1722) <= (layer2_outputs(2711)) xor (layer2_outputs(3095));
    outputs(1723) <= (layer2_outputs(1498)) and not (layer2_outputs(952));
    outputs(1724) <= not(layer2_outputs(2705));
    outputs(1725) <= layer2_outputs(2928);
    outputs(1726) <= not(layer2_outputs(2728));
    outputs(1727) <= layer2_outputs(2098);
    outputs(1728) <= layer2_outputs(790);
    outputs(1729) <= layer2_outputs(3956);
    outputs(1730) <= not((layer2_outputs(664)) and (layer2_outputs(3166)));
    outputs(1731) <= layer2_outputs(2560);
    outputs(1732) <= not(layer2_outputs(282));
    outputs(1733) <= not(layer2_outputs(5026));
    outputs(1734) <= not(layer2_outputs(3528));
    outputs(1735) <= (layer2_outputs(1694)) and not (layer2_outputs(4718));
    outputs(1736) <= not(layer2_outputs(1523));
    outputs(1737) <= layer2_outputs(1149);
    outputs(1738) <= (layer2_outputs(4563)) and (layer2_outputs(2528));
    outputs(1739) <= (layer2_outputs(1351)) and not (layer2_outputs(967));
    outputs(1740) <= layer2_outputs(4551);
    outputs(1741) <= not(layer2_outputs(1122));
    outputs(1742) <= layer2_outputs(734);
    outputs(1743) <= not(layer2_outputs(4035));
    outputs(1744) <= not(layer2_outputs(1265));
    outputs(1745) <= not((layer2_outputs(2416)) xor (layer2_outputs(3913)));
    outputs(1746) <= (layer2_outputs(3259)) xor (layer2_outputs(3993));
    outputs(1747) <= layer2_outputs(2242);
    outputs(1748) <= layer2_outputs(1959);
    outputs(1749) <= not((layer2_outputs(4589)) or (layer2_outputs(1633)));
    outputs(1750) <= not(layer2_outputs(3851)) or (layer2_outputs(3836));
    outputs(1751) <= not(layer2_outputs(2663));
    outputs(1752) <= not(layer2_outputs(126));
    outputs(1753) <= not(layer2_outputs(538));
    outputs(1754) <= not(layer2_outputs(1555));
    outputs(1755) <= not(layer2_outputs(214)) or (layer2_outputs(4570));
    outputs(1756) <= not((layer2_outputs(4854)) xor (layer2_outputs(3131)));
    outputs(1757) <= not(layer2_outputs(1486));
    outputs(1758) <= not(layer2_outputs(1173)) or (layer2_outputs(3723));
    outputs(1759) <= not(layer2_outputs(1128));
    outputs(1760) <= not((layer2_outputs(2975)) xor (layer2_outputs(3136)));
    outputs(1761) <= not(layer2_outputs(3546));
    outputs(1762) <= (layer2_outputs(2504)) and not (layer2_outputs(5008));
    outputs(1763) <= not(layer2_outputs(2916));
    outputs(1764) <= not((layer2_outputs(2202)) xor (layer2_outputs(3731)));
    outputs(1765) <= not(layer2_outputs(1952));
    outputs(1766) <= not(layer2_outputs(4703));
    outputs(1767) <= not(layer2_outputs(638));
    outputs(1768) <= not(layer2_outputs(1805));
    outputs(1769) <= not(layer2_outputs(3936));
    outputs(1770) <= (layer2_outputs(4192)) xor (layer2_outputs(4106));
    outputs(1771) <= not(layer2_outputs(4549));
    outputs(1772) <= (layer2_outputs(3382)) xor (layer2_outputs(4853));
    outputs(1773) <= not(layer2_outputs(3816));
    outputs(1774) <= layer2_outputs(873);
    outputs(1775) <= not(layer2_outputs(3462));
    outputs(1776) <= not((layer2_outputs(272)) xor (layer2_outputs(2084)));
    outputs(1777) <= layer2_outputs(1917);
    outputs(1778) <= not(layer2_outputs(2432)) or (layer2_outputs(995));
    outputs(1779) <= layer2_outputs(219);
    outputs(1780) <= not(layer2_outputs(206));
    outputs(1781) <= not(layer2_outputs(778));
    outputs(1782) <= layer2_outputs(96);
    outputs(1783) <= layer2_outputs(4797);
    outputs(1784) <= layer2_outputs(110);
    outputs(1785) <= (layer2_outputs(845)) xor (layer2_outputs(2976));
    outputs(1786) <= not(layer2_outputs(810));
    outputs(1787) <= (layer2_outputs(1567)) and not (layer2_outputs(4096));
    outputs(1788) <= (layer2_outputs(1485)) xor (layer2_outputs(1732));
    outputs(1789) <= layer2_outputs(5040);
    outputs(1790) <= (layer2_outputs(891)) or (layer2_outputs(2083));
    outputs(1791) <= (layer2_outputs(2685)) and not (layer2_outputs(4017));
    outputs(1792) <= not(layer2_outputs(4359));
    outputs(1793) <= (layer2_outputs(2604)) xor (layer2_outputs(3303));
    outputs(1794) <= not(layer2_outputs(1097));
    outputs(1795) <= layer2_outputs(433);
    outputs(1796) <= layer2_outputs(16);
    outputs(1797) <= layer2_outputs(2560);
    outputs(1798) <= layer2_outputs(3519);
    outputs(1799) <= not((layer2_outputs(328)) xor (layer2_outputs(2320)));
    outputs(1800) <= not((layer2_outputs(4907)) and (layer2_outputs(4861)));
    outputs(1801) <= layer2_outputs(3756);
    outputs(1802) <= not((layer2_outputs(2494)) and (layer2_outputs(4394)));
    outputs(1803) <= layer2_outputs(3771);
    outputs(1804) <= layer2_outputs(4138);
    outputs(1805) <= (layer2_outputs(3244)) xor (layer2_outputs(2460));
    outputs(1806) <= (layer2_outputs(387)) xor (layer2_outputs(1929));
    outputs(1807) <= not(layer2_outputs(4708));
    outputs(1808) <= not(layer2_outputs(4327));
    outputs(1809) <= layer2_outputs(4766);
    outputs(1810) <= (layer2_outputs(4511)) xor (layer2_outputs(1192));
    outputs(1811) <= not((layer2_outputs(736)) xor (layer2_outputs(3168)));
    outputs(1812) <= not(layer2_outputs(4733));
    outputs(1813) <= layer2_outputs(566);
    outputs(1814) <= not(layer2_outputs(1924));
    outputs(1815) <= (layer2_outputs(4636)) and not (layer2_outputs(3687));
    outputs(1816) <= layer2_outputs(4693);
    outputs(1817) <= layer2_outputs(1120);
    outputs(1818) <= not(layer2_outputs(4958));
    outputs(1819) <= not(layer2_outputs(3823));
    outputs(1820) <= not(layer2_outputs(466));
    outputs(1821) <= layer2_outputs(4518);
    outputs(1822) <= not((layer2_outputs(400)) xor (layer2_outputs(3777)));
    outputs(1823) <= (layer2_outputs(3005)) xor (layer2_outputs(3520));
    outputs(1824) <= not(layer2_outputs(1855)) or (layer2_outputs(528));
    outputs(1825) <= layer2_outputs(634);
    outputs(1826) <= not(layer2_outputs(293));
    outputs(1827) <= layer2_outputs(1339);
    outputs(1828) <= layer2_outputs(350);
    outputs(1829) <= not(layer2_outputs(3062)) or (layer2_outputs(3863));
    outputs(1830) <= layer2_outputs(2579);
    outputs(1831) <= not((layer2_outputs(3807)) xor (layer2_outputs(2206)));
    outputs(1832) <= layer2_outputs(3628);
    outputs(1833) <= layer2_outputs(5104);
    outputs(1834) <= not((layer2_outputs(4370)) xor (layer2_outputs(150)));
    outputs(1835) <= layer2_outputs(4658);
    outputs(1836) <= not(layer2_outputs(2065));
    outputs(1837) <= layer2_outputs(1145);
    outputs(1838) <= (layer2_outputs(2650)) and not (layer2_outputs(5115));
    outputs(1839) <= not(layer2_outputs(4897));
    outputs(1840) <= (layer2_outputs(3754)) and not (layer2_outputs(1544));
    outputs(1841) <= not((layer2_outputs(616)) xor (layer2_outputs(3045)));
    outputs(1842) <= not(layer2_outputs(643));
    outputs(1843) <= not(layer2_outputs(1738));
    outputs(1844) <= not(layer2_outputs(2966));
    outputs(1845) <= not(layer2_outputs(437));
    outputs(1846) <= (layer2_outputs(3399)) and not (layer2_outputs(1327));
    outputs(1847) <= not(layer2_outputs(90));
    outputs(1848) <= not((layer2_outputs(1286)) xor (layer2_outputs(2555)));
    outputs(1849) <= (layer2_outputs(4776)) and (layer2_outputs(4086));
    outputs(1850) <= not(layer2_outputs(569)) or (layer2_outputs(3839));
    outputs(1851) <= (layer2_outputs(2762)) xor (layer2_outputs(480));
    outputs(1852) <= not(layer2_outputs(1254)) or (layer2_outputs(1547));
    outputs(1853) <= layer2_outputs(3318);
    outputs(1854) <= layer2_outputs(1784);
    outputs(1855) <= not(layer2_outputs(4708));
    outputs(1856) <= (layer2_outputs(2134)) and not (layer2_outputs(3860));
    outputs(1857) <= not(layer2_outputs(1264));
    outputs(1858) <= layer2_outputs(2732);
    outputs(1859) <= (layer2_outputs(1595)) xor (layer2_outputs(2150));
    outputs(1860) <= (layer2_outputs(3007)) xor (layer2_outputs(4799));
    outputs(1861) <= layer2_outputs(2009);
    outputs(1862) <= (layer2_outputs(3012)) and (layer2_outputs(356));
    outputs(1863) <= layer2_outputs(3939);
    outputs(1864) <= not((layer2_outputs(3041)) or (layer2_outputs(2724)));
    outputs(1865) <= not((layer2_outputs(2225)) xor (layer2_outputs(3435)));
    outputs(1866) <= layer2_outputs(2750);
    outputs(1867) <= not(layer2_outputs(3566));
    outputs(1868) <= not(layer2_outputs(966)) or (layer2_outputs(2626));
    outputs(1869) <= layer2_outputs(1812);
    outputs(1870) <= not((layer2_outputs(972)) and (layer2_outputs(2966)));
    outputs(1871) <= not(layer2_outputs(1635));
    outputs(1872) <= not(layer2_outputs(1166));
    outputs(1873) <= not((layer2_outputs(3253)) or (layer2_outputs(2252)));
    outputs(1874) <= not((layer2_outputs(2866)) and (layer2_outputs(3662)));
    outputs(1875) <= layer2_outputs(867);
    outputs(1876) <= not(layer2_outputs(4253));
    outputs(1877) <= (layer2_outputs(2730)) and not (layer2_outputs(2792));
    outputs(1878) <= (layer2_outputs(2291)) or (layer2_outputs(4975));
    outputs(1879) <= (layer2_outputs(828)) or (layer2_outputs(3364));
    outputs(1880) <= not(layer2_outputs(2589));
    outputs(1881) <= layer2_outputs(4531);
    outputs(1882) <= not(layer2_outputs(2782));
    outputs(1883) <= (layer2_outputs(4224)) and not (layer2_outputs(633));
    outputs(1884) <= (layer2_outputs(2525)) and not (layer2_outputs(4405));
    outputs(1885) <= not(layer2_outputs(2925));
    outputs(1886) <= (layer2_outputs(5)) and not (layer2_outputs(1745));
    outputs(1887) <= (layer2_outputs(2929)) xor (layer2_outputs(3647));
    outputs(1888) <= not((layer2_outputs(2082)) xor (layer2_outputs(839)));
    outputs(1889) <= not(layer2_outputs(1966));
    outputs(1890) <= layer2_outputs(1328);
    outputs(1891) <= not((layer2_outputs(270)) or (layer2_outputs(2453)));
    outputs(1892) <= not(layer2_outputs(2179));
    outputs(1893) <= not(layer2_outputs(1972));
    outputs(1894) <= layer2_outputs(4124);
    outputs(1895) <= not(layer2_outputs(369));
    outputs(1896) <= (layer2_outputs(725)) or (layer2_outputs(819));
    outputs(1897) <= layer2_outputs(2001);
    outputs(1898) <= not(layer2_outputs(178));
    outputs(1899) <= not(layer2_outputs(3860));
    outputs(1900) <= layer2_outputs(3368);
    outputs(1901) <= layer2_outputs(4585);
    outputs(1902) <= not(layer2_outputs(3484));
    outputs(1903) <= not((layer2_outputs(2939)) xor (layer2_outputs(3553)));
    outputs(1904) <= not((layer2_outputs(4112)) and (layer2_outputs(2035)));
    outputs(1905) <= layer2_outputs(2121);
    outputs(1906) <= (layer2_outputs(3857)) and (layer2_outputs(3017));
    outputs(1907) <= not(layer2_outputs(3764));
    outputs(1908) <= (layer2_outputs(366)) or (layer2_outputs(3806));
    outputs(1909) <= layer2_outputs(51);
    outputs(1910) <= not((layer2_outputs(1248)) and (layer2_outputs(103)));
    outputs(1911) <= layer2_outputs(1418);
    outputs(1912) <= (layer2_outputs(3642)) and not (layer2_outputs(1203));
    outputs(1913) <= not(layer2_outputs(1318));
    outputs(1914) <= not(layer2_outputs(3895)) or (layer2_outputs(899));
    outputs(1915) <= (layer2_outputs(4690)) and not (layer2_outputs(3029));
    outputs(1916) <= not(layer2_outputs(331));
    outputs(1917) <= layer2_outputs(1931);
    outputs(1918) <= not(layer2_outputs(4951));
    outputs(1919) <= (layer2_outputs(116)) and not (layer2_outputs(1622));
    outputs(1920) <= not(layer2_outputs(2845));
    outputs(1921) <= not(layer2_outputs(2708));
    outputs(1922) <= not((layer2_outputs(4576)) xor (layer2_outputs(1022)));
    outputs(1923) <= layer2_outputs(4380);
    outputs(1924) <= layer2_outputs(4452);
    outputs(1925) <= (layer2_outputs(4568)) xor (layer2_outputs(1138));
    outputs(1926) <= layer2_outputs(4220);
    outputs(1927) <= not((layer2_outputs(1565)) xor (layer2_outputs(386)));
    outputs(1928) <= (layer2_outputs(3637)) or (layer2_outputs(2690));
    outputs(1929) <= not(layer2_outputs(3998));
    outputs(1930) <= (layer2_outputs(1870)) and (layer2_outputs(767));
    outputs(1931) <= not((layer2_outputs(2672)) xor (layer2_outputs(362)));
    outputs(1932) <= layer2_outputs(929);
    outputs(1933) <= (layer2_outputs(3376)) and (layer2_outputs(779));
    outputs(1934) <= not(layer2_outputs(1545));
    outputs(1935) <= not(layer2_outputs(4899));
    outputs(1936) <= (layer2_outputs(2980)) xor (layer2_outputs(1187));
    outputs(1937) <= not((layer2_outputs(4160)) xor (layer2_outputs(4774)));
    outputs(1938) <= not((layer2_outputs(1375)) and (layer2_outputs(3561)));
    outputs(1939) <= not(layer2_outputs(3493));
    outputs(1940) <= (layer2_outputs(2283)) xor (layer2_outputs(674));
    outputs(1941) <= not(layer2_outputs(3264));
    outputs(1942) <= (layer2_outputs(4123)) or (layer2_outputs(4761));
    outputs(1943) <= (layer2_outputs(4932)) and (layer2_outputs(4709));
    outputs(1944) <= layer2_outputs(820);
    outputs(1945) <= layer2_outputs(1223);
    outputs(1946) <= not(layer2_outputs(1233));
    outputs(1947) <= not(layer2_outputs(4899));
    outputs(1948) <= layer2_outputs(1301);
    outputs(1949) <= layer2_outputs(2500);
    outputs(1950) <= layer2_outputs(409);
    outputs(1951) <= (layer2_outputs(2729)) xor (layer2_outputs(3530));
    outputs(1952) <= not(layer2_outputs(4660)) or (layer2_outputs(989));
    outputs(1953) <= (layer2_outputs(313)) and (layer2_outputs(1920));
    outputs(1954) <= layer2_outputs(4678);
    outputs(1955) <= not(layer2_outputs(5105));
    outputs(1956) <= not(layer2_outputs(4731)) or (layer2_outputs(4175));
    outputs(1957) <= not((layer2_outputs(939)) or (layer2_outputs(4500)));
    outputs(1958) <= layer2_outputs(4794);
    outputs(1959) <= not(layer2_outputs(4289));
    outputs(1960) <= layer2_outputs(4000);
    outputs(1961) <= not(layer2_outputs(324));
    outputs(1962) <= not(layer2_outputs(3597));
    outputs(1963) <= not(layer2_outputs(1278)) or (layer2_outputs(1341));
    outputs(1964) <= not((layer2_outputs(4623)) and (layer2_outputs(4883)));
    outputs(1965) <= not(layer2_outputs(4322));
    outputs(1966) <= layer2_outputs(4330);
    outputs(1967) <= layer2_outputs(1170);
    outputs(1968) <= not(layer2_outputs(1714));
    outputs(1969) <= not((layer2_outputs(2661)) xor (layer2_outputs(4917)));
    outputs(1970) <= not(layer2_outputs(1359));
    outputs(1971) <= layer2_outputs(1148);
    outputs(1972) <= (layer2_outputs(4525)) and not (layer2_outputs(2357));
    outputs(1973) <= not(layer2_outputs(4439));
    outputs(1974) <= layer2_outputs(494);
    outputs(1975) <= not(layer2_outputs(2429));
    outputs(1976) <= not(layer2_outputs(1377));
    outputs(1977) <= (layer2_outputs(243)) xor (layer2_outputs(3077));
    outputs(1978) <= (layer2_outputs(4307)) and not (layer2_outputs(2016));
    outputs(1979) <= layer2_outputs(1620);
    outputs(1980) <= (layer2_outputs(1803)) or (layer2_outputs(4165));
    outputs(1981) <= not(layer2_outputs(3914));
    outputs(1982) <= (layer2_outputs(440)) and not (layer2_outputs(4881));
    outputs(1983) <= layer2_outputs(1094);
    outputs(1984) <= not(layer2_outputs(1884));
    outputs(1985) <= layer2_outputs(198);
    outputs(1986) <= layer2_outputs(4778);
    outputs(1987) <= (layer2_outputs(4795)) or (layer2_outputs(1064));
    outputs(1988) <= not(layer2_outputs(749));
    outputs(1989) <= not(layer2_outputs(3452));
    outputs(1990) <= not(layer2_outputs(1394));
    outputs(1991) <= (layer2_outputs(1534)) xor (layer2_outputs(130));
    outputs(1992) <= layer2_outputs(3550);
    outputs(1993) <= not(layer2_outputs(2790));
    outputs(1994) <= not((layer2_outputs(2522)) or (layer2_outputs(1043)));
    outputs(1995) <= not(layer2_outputs(3635)) or (layer2_outputs(1995));
    outputs(1996) <= layer2_outputs(1791);
    outputs(1997) <= not((layer2_outputs(4968)) xor (layer2_outputs(3970)));
    outputs(1998) <= (layer2_outputs(901)) xor (layer2_outputs(2615));
    outputs(1999) <= not(layer2_outputs(3023));
    outputs(2000) <= not((layer2_outputs(3432)) or (layer2_outputs(4053)));
    outputs(2001) <= not(layer2_outputs(370));
    outputs(2002) <= layer2_outputs(3223);
    outputs(2003) <= not(layer2_outputs(3851));
    outputs(2004) <= (layer2_outputs(429)) and not (layer2_outputs(2454));
    outputs(2005) <= layer2_outputs(4211);
    outputs(2006) <= not(layer2_outputs(2587));
    outputs(2007) <= layer2_outputs(796);
    outputs(2008) <= layer2_outputs(1659);
    outputs(2009) <= not(layer2_outputs(2947));
    outputs(2010) <= not((layer2_outputs(2039)) or (layer2_outputs(269)));
    outputs(2011) <= layer2_outputs(2204);
    outputs(2012) <= not((layer2_outputs(2362)) and (layer2_outputs(3695)));
    outputs(2013) <= not(layer2_outputs(2714));
    outputs(2014) <= not((layer2_outputs(3236)) or (layer2_outputs(579)));
    outputs(2015) <= not(layer2_outputs(2793)) or (layer2_outputs(610));
    outputs(2016) <= not(layer2_outputs(4420));
    outputs(2017) <= not(layer2_outputs(5022));
    outputs(2018) <= layer2_outputs(1748);
    outputs(2019) <= (layer2_outputs(2899)) xor (layer2_outputs(4470));
    outputs(2020) <= not((layer2_outputs(2220)) xor (layer2_outputs(2633)));
    outputs(2021) <= not(layer2_outputs(4346));
    outputs(2022) <= not(layer2_outputs(94));
    outputs(2023) <= layer2_outputs(4947);
    outputs(2024) <= not(layer2_outputs(689));
    outputs(2025) <= (layer2_outputs(2733)) xor (layer2_outputs(1355));
    outputs(2026) <= not(layer2_outputs(9)) or (layer2_outputs(3776));
    outputs(2027) <= not((layer2_outputs(3994)) xor (layer2_outputs(215)));
    outputs(2028) <= layer2_outputs(4422);
    outputs(2029) <= layer2_outputs(2941);
    outputs(2030) <= layer2_outputs(3408);
    outputs(2031) <= not(layer2_outputs(4707));
    outputs(2032) <= layer2_outputs(3365);
    outputs(2033) <= (layer2_outputs(84)) and not (layer2_outputs(4526));
    outputs(2034) <= not(layer2_outputs(1507));
    outputs(2035) <= not((layer2_outputs(3556)) xor (layer2_outputs(3077)));
    outputs(2036) <= not(layer2_outputs(124));
    outputs(2037) <= layer2_outputs(2811);
    outputs(2038) <= not(layer2_outputs(98));
    outputs(2039) <= layer2_outputs(88);
    outputs(2040) <= not((layer2_outputs(3547)) xor (layer2_outputs(232)));
    outputs(2041) <= not((layer2_outputs(1127)) xor (layer2_outputs(1252)));
    outputs(2042) <= not(layer2_outputs(1570));
    outputs(2043) <= layer2_outputs(2428);
    outputs(2044) <= not(layer2_outputs(2055));
    outputs(2045) <= not((layer2_outputs(3740)) xor (layer2_outputs(4003)));
    outputs(2046) <= (layer2_outputs(4878)) and not (layer2_outputs(3805));
    outputs(2047) <= not(layer2_outputs(522));
    outputs(2048) <= not((layer2_outputs(3207)) xor (layer2_outputs(2564)));
    outputs(2049) <= not((layer2_outputs(646)) xor (layer2_outputs(3471)));
    outputs(2050) <= not(layer2_outputs(2766));
    outputs(2051) <= layer2_outputs(4475);
    outputs(2052) <= (layer2_outputs(923)) xor (layer2_outputs(5111));
    outputs(2053) <= layer2_outputs(2573);
    outputs(2054) <= (layer2_outputs(306)) and not (layer2_outputs(1968));
    outputs(2055) <= (layer2_outputs(751)) and (layer2_outputs(648));
    outputs(2056) <= layer2_outputs(1390);
    outputs(2057) <= (layer2_outputs(1608)) and not (layer2_outputs(3615));
    outputs(2058) <= not(layer2_outputs(326));
    outputs(2059) <= layer2_outputs(4715);
    outputs(2060) <= not(layer2_outputs(4754));
    outputs(2061) <= layer2_outputs(2293);
    outputs(2062) <= not(layer2_outputs(2170));
    outputs(2063) <= layer2_outputs(3711);
    outputs(2064) <= not((layer2_outputs(3532)) or (layer2_outputs(1216)));
    outputs(2065) <= layer2_outputs(1570);
    outputs(2066) <= (layer2_outputs(3914)) and not (layer2_outputs(3025));
    outputs(2067) <= layer2_outputs(3343);
    outputs(2068) <= not((layer2_outputs(2781)) and (layer2_outputs(2241)));
    outputs(2069) <= (layer2_outputs(260)) and not (layer2_outputs(4330));
    outputs(2070) <= not(layer2_outputs(886));
    outputs(2071) <= layer2_outputs(1813);
    outputs(2072) <= not(layer2_outputs(4231));
    outputs(2073) <= not(layer2_outputs(2224));
    outputs(2074) <= layer2_outputs(4369);
    outputs(2075) <= layer2_outputs(2600);
    outputs(2076) <= layer2_outputs(1928);
    outputs(2077) <= layer2_outputs(3495);
    outputs(2078) <= (layer2_outputs(404)) and not (layer2_outputs(3108));
    outputs(2079) <= not(layer2_outputs(4574)) or (layer2_outputs(252));
    outputs(2080) <= layer2_outputs(399);
    outputs(2081) <= (layer2_outputs(1125)) xor (layer2_outputs(4260));
    outputs(2082) <= not(layer2_outputs(2053));
    outputs(2083) <= not((layer2_outputs(374)) xor (layer2_outputs(4075)));
    outputs(2084) <= (layer2_outputs(1756)) and (layer2_outputs(1129));
    outputs(2085) <= layer2_outputs(2257);
    outputs(2086) <= (layer2_outputs(4066)) and not (layer2_outputs(4361));
    outputs(2087) <= not(layer2_outputs(3766));
    outputs(2088) <= layer2_outputs(1513);
    outputs(2089) <= (layer2_outputs(196)) and not (layer2_outputs(2292));
    outputs(2090) <= not(layer2_outputs(800)) or (layer2_outputs(2157));
    outputs(2091) <= not(layer2_outputs(1148));
    outputs(2092) <= layer2_outputs(3548);
    outputs(2093) <= not(layer2_outputs(5085));
    outputs(2094) <= (layer2_outputs(4653)) and (layer2_outputs(1634));
    outputs(2095) <= not((layer2_outputs(4316)) or (layer2_outputs(113)));
    outputs(2096) <= (layer2_outputs(4900)) xor (layer2_outputs(3053));
    outputs(2097) <= not((layer2_outputs(4445)) or (layer2_outputs(1710)));
    outputs(2098) <= layer2_outputs(9);
    outputs(2099) <= not(layer2_outputs(446));
    outputs(2100) <= layer2_outputs(1719);
    outputs(2101) <= not(layer2_outputs(3285));
    outputs(2102) <= (layer2_outputs(5090)) and not (layer2_outputs(1132));
    outputs(2103) <= not(layer2_outputs(2815));
    outputs(2104) <= (layer2_outputs(2684)) and (layer2_outputs(4265));
    outputs(2105) <= (layer2_outputs(34)) xor (layer2_outputs(3736));
    outputs(2106) <= layer2_outputs(4746);
    outputs(2107) <= not((layer2_outputs(2513)) or (layer2_outputs(3458)));
    outputs(2108) <= (layer2_outputs(2807)) and (layer2_outputs(1491));
    outputs(2109) <= not((layer2_outputs(2934)) and (layer2_outputs(3576)));
    outputs(2110) <= layer2_outputs(4856);
    outputs(2111) <= not(layer2_outputs(4579));
    outputs(2112) <= (layer2_outputs(415)) xor (layer2_outputs(1935));
    outputs(2113) <= (layer2_outputs(2514)) xor (layer2_outputs(1211));
    outputs(2114) <= not(layer2_outputs(4347));
    outputs(2115) <= not(layer2_outputs(3384));
    outputs(2116) <= layer2_outputs(3151);
    outputs(2117) <= layer2_outputs(1769);
    outputs(2118) <= not(layer2_outputs(1904));
    outputs(2119) <= (layer2_outputs(4056)) xor (layer2_outputs(344));
    outputs(2120) <= (layer2_outputs(5067)) and not (layer2_outputs(3347));
    outputs(2121) <= layer2_outputs(213);
    outputs(2122) <= (layer2_outputs(3621)) and (layer2_outputs(3882));
    outputs(2123) <= (layer2_outputs(1388)) and not (layer2_outputs(5010));
    outputs(2124) <= (layer2_outputs(4337)) xor (layer2_outputs(856));
    outputs(2125) <= layer2_outputs(1723);
    outputs(2126) <= layer2_outputs(3142);
    outputs(2127) <= layer2_outputs(201);
    outputs(2128) <= not(layer2_outputs(1237));
    outputs(2129) <= (layer2_outputs(1700)) and not (layer2_outputs(1));
    outputs(2130) <= layer2_outputs(4074);
    outputs(2131) <= not(layer2_outputs(1149));
    outputs(2132) <= layer2_outputs(1753);
    outputs(2133) <= not(layer2_outputs(4424));
    outputs(2134) <= layer2_outputs(3247);
    outputs(2135) <= not((layer2_outputs(4091)) or (layer2_outputs(2347)));
    outputs(2136) <= not((layer2_outputs(2268)) or (layer2_outputs(509)));
    outputs(2137) <= layer2_outputs(4319);
    outputs(2138) <= not(layer2_outputs(100));
    outputs(2139) <= not((layer2_outputs(3861)) xor (layer2_outputs(5060)));
    outputs(2140) <= (layer2_outputs(1202)) xor (layer2_outputs(3760));
    outputs(2141) <= layer2_outputs(2084);
    outputs(2142) <= not(layer2_outputs(3585));
    outputs(2143) <= not(layer2_outputs(3337));
    outputs(2144) <= not((layer2_outputs(2630)) or (layer2_outputs(3940)));
    outputs(2145) <= layer2_outputs(2383);
    outputs(2146) <= not(layer2_outputs(667));
    outputs(2147) <= (layer2_outputs(2945)) xor (layer2_outputs(2052));
    outputs(2148) <= not(layer2_outputs(2464));
    outputs(2149) <= (layer2_outputs(2440)) and not (layer2_outputs(2708));
    outputs(2150) <= (layer2_outputs(4281)) and (layer2_outputs(4193));
    outputs(2151) <= not((layer2_outputs(4100)) or (layer2_outputs(4754)));
    outputs(2152) <= layer2_outputs(707);
    outputs(2153) <= not((layer2_outputs(3779)) or (layer2_outputs(2662)));
    outputs(2154) <= not(layer2_outputs(2749));
    outputs(2155) <= (layer2_outputs(4154)) xor (layer2_outputs(491));
    outputs(2156) <= not(layer2_outputs(1255));
    outputs(2157) <= layer2_outputs(3203);
    outputs(2158) <= not(layer2_outputs(4797));
    outputs(2159) <= not(layer2_outputs(1772));
    outputs(2160) <= (layer2_outputs(3394)) and (layer2_outputs(339));
    outputs(2161) <= layer2_outputs(125);
    outputs(2162) <= layer2_outputs(197);
    outputs(2163) <= (layer2_outputs(3436)) xor (layer2_outputs(1858));
    outputs(2164) <= not(layer2_outputs(2843));
    outputs(2165) <= not(layer2_outputs(821));
    outputs(2166) <= not(layer2_outputs(2019));
    outputs(2167) <= (layer2_outputs(1652)) xor (layer2_outputs(857));
    outputs(2168) <= not(layer2_outputs(4781));
    outputs(2169) <= (layer2_outputs(4292)) xor (layer2_outputs(568));
    outputs(2170) <= not(layer2_outputs(2141)) or (layer2_outputs(1203));
    outputs(2171) <= not(layer2_outputs(4418));
    outputs(2172) <= (layer2_outputs(1764)) and not (layer2_outputs(3975));
    outputs(2173) <= not(layer2_outputs(145));
    outputs(2174) <= not(layer2_outputs(609));
    outputs(2175) <= layer2_outputs(3611);
    outputs(2176) <= not(layer2_outputs(4546));
    outputs(2177) <= not((layer2_outputs(4264)) xor (layer2_outputs(3964)));
    outputs(2178) <= (layer2_outputs(719)) and not (layer2_outputs(1869));
    outputs(2179) <= not((layer2_outputs(3258)) xor (layer2_outputs(4790)));
    outputs(2180) <= not(layer2_outputs(4712));
    outputs(2181) <= not(layer2_outputs(3022));
    outputs(2182) <= layer2_outputs(723);
    outputs(2183) <= layer2_outputs(3996);
    outputs(2184) <= layer2_outputs(359);
    outputs(2185) <= not(layer2_outputs(247));
    outputs(2186) <= not(layer2_outputs(2304));
    outputs(2187) <= not((layer2_outputs(3648)) or (layer2_outputs(1725)));
    outputs(2188) <= not(layer2_outputs(4345));
    outputs(2189) <= (layer2_outputs(3987)) xor (layer2_outputs(704));
    outputs(2190) <= (layer2_outputs(4393)) and not (layer2_outputs(4471));
    outputs(2191) <= (layer2_outputs(85)) and (layer2_outputs(1138));
    outputs(2192) <= not(layer2_outputs(3959));
    outputs(2193) <= layer2_outputs(2208);
    outputs(2194) <= layer2_outputs(3581);
    outputs(2195) <= not(layer2_outputs(2713));
    outputs(2196) <= layer2_outputs(4811);
    outputs(2197) <= layer2_outputs(2459);
    outputs(2198) <= not(layer2_outputs(1804));
    outputs(2199) <= not(layer2_outputs(1170));
    outputs(2200) <= not(layer2_outputs(4329));
    outputs(2201) <= not(layer2_outputs(750));
    outputs(2202) <= (layer2_outputs(455)) and not (layer2_outputs(4894));
    outputs(2203) <= not(layer2_outputs(1093));
    outputs(2204) <= not(layer2_outputs(4218));
    outputs(2205) <= layer2_outputs(4796);
    outputs(2206) <= not(layer2_outputs(2611));
    outputs(2207) <= layer2_outputs(1632);
    outputs(2208) <= not((layer2_outputs(1030)) xor (layer2_outputs(2214)));
    outputs(2209) <= layer2_outputs(199);
    outputs(2210) <= (layer2_outputs(1183)) or (layer2_outputs(4809));
    outputs(2211) <= not(layer2_outputs(1070));
    outputs(2212) <= not((layer2_outputs(4415)) or (layer2_outputs(286)));
    outputs(2213) <= layer2_outputs(92);
    outputs(2214) <= (layer2_outputs(1098)) xor (layer2_outputs(345));
    outputs(2215) <= not((layer2_outputs(4047)) xor (layer2_outputs(3534)));
    outputs(2216) <= (layer2_outputs(1358)) xor (layer2_outputs(3911));
    outputs(2217) <= not(layer2_outputs(1724)) or (layer2_outputs(4789));
    outputs(2218) <= not(layer2_outputs(1193));
    outputs(2219) <= not(layer2_outputs(3694));
    outputs(2220) <= not((layer2_outputs(1086)) xor (layer2_outputs(1370)));
    outputs(2221) <= layer2_outputs(1702);
    outputs(2222) <= layer2_outputs(1487);
    outputs(2223) <= not(layer2_outputs(2681));
    outputs(2224) <= (layer2_outputs(2628)) xor (layer2_outputs(188));
    outputs(2225) <= layer2_outputs(4847);
    outputs(2226) <= layer2_outputs(903);
    outputs(2227) <= layer2_outputs(4136);
    outputs(2228) <= layer2_outputs(213);
    outputs(2229) <= layer2_outputs(648);
    outputs(2230) <= (layer2_outputs(4717)) xor (layer2_outputs(3541));
    outputs(2231) <= not(layer2_outputs(2665));
    outputs(2232) <= not((layer2_outputs(1656)) xor (layer2_outputs(5060)));
    outputs(2233) <= not((layer2_outputs(3087)) and (layer2_outputs(4149)));
    outputs(2234) <= layer2_outputs(3538);
    outputs(2235) <= not(layer2_outputs(2915));
    outputs(2236) <= layer2_outputs(94);
    outputs(2237) <= layer2_outputs(4931);
    outputs(2238) <= (layer2_outputs(5)) xor (layer2_outputs(316));
    outputs(2239) <= (layer2_outputs(799)) xor (layer2_outputs(3314));
    outputs(2240) <= layer2_outputs(4061);
    outputs(2241) <= layer2_outputs(2881);
    outputs(2242) <= not(layer2_outputs(2569));
    outputs(2243) <= layer2_outputs(630);
    outputs(2244) <= layer2_outputs(380);
    outputs(2245) <= not((layer2_outputs(4116)) or (layer2_outputs(2782)));
    outputs(2246) <= not(layer2_outputs(3969));
    outputs(2247) <= not(layer2_outputs(782)) or (layer2_outputs(2440));
    outputs(2248) <= not(layer2_outputs(1783)) or (layer2_outputs(1019));
    outputs(2249) <= layer2_outputs(2059);
    outputs(2250) <= (layer2_outputs(5086)) and not (layer2_outputs(4712));
    outputs(2251) <= (layer2_outputs(2678)) and not (layer2_outputs(4272));
    outputs(2252) <= (layer2_outputs(1819)) and not (layer2_outputs(3813));
    outputs(2253) <= not((layer2_outputs(1251)) or (layer2_outputs(3352)));
    outputs(2254) <= not((layer2_outputs(2471)) xor (layer2_outputs(3730)));
    outputs(2255) <= layer2_outputs(753);
    outputs(2256) <= not(layer2_outputs(2031));
    outputs(2257) <= not(layer2_outputs(1152));
    outputs(2258) <= (layer2_outputs(45)) or (layer2_outputs(4972));
    outputs(2259) <= (layer2_outputs(955)) xor (layer2_outputs(1250));
    outputs(2260) <= not((layer2_outputs(3940)) xor (layer2_outputs(3572)));
    outputs(2261) <= not(layer2_outputs(1665));
    outputs(2262) <= (layer2_outputs(5109)) and not (layer2_outputs(847));
    outputs(2263) <= (layer2_outputs(2111)) and not (layer2_outputs(2709));
    outputs(2264) <= (layer2_outputs(79)) xor (layer2_outputs(2511));
    outputs(2265) <= not(layer2_outputs(4611));
    outputs(2266) <= not((layer2_outputs(4097)) or (layer2_outputs(334)));
    outputs(2267) <= not((layer2_outputs(2869)) xor (layer2_outputs(207)));
    outputs(2268) <= not(layer2_outputs(1368));
    outputs(2269) <= layer2_outputs(1164);
    outputs(2270) <= (layer2_outputs(120)) and not (layer2_outputs(3582));
    outputs(2271) <= not(layer2_outputs(3609));
    outputs(2272) <= layer2_outputs(691);
    outputs(2273) <= layer2_outputs(1392);
    outputs(2274) <= not(layer2_outputs(3137));
    outputs(2275) <= (layer2_outputs(4788)) and (layer2_outputs(4623));
    outputs(2276) <= not(layer2_outputs(4983)) or (layer2_outputs(4069));
    outputs(2277) <= (layer2_outputs(2949)) xor (layer2_outputs(3050));
    outputs(2278) <= not((layer2_outputs(3283)) or (layer2_outputs(2333)));
    outputs(2279) <= not(layer2_outputs(4208));
    outputs(2280) <= not((layer2_outputs(450)) xor (layer2_outputs(839)));
    outputs(2281) <= not(layer2_outputs(2406));
    outputs(2282) <= (layer2_outputs(3514)) and (layer2_outputs(3704));
    outputs(2283) <= not(layer2_outputs(1829));
    outputs(2284) <= layer2_outputs(2822);
    outputs(2285) <= (layer2_outputs(3381)) and (layer2_outputs(2289));
    outputs(2286) <= not((layer2_outputs(2871)) xor (layer2_outputs(4720)));
    outputs(2287) <= (layer2_outputs(1595)) and not (layer2_outputs(4027));
    outputs(2288) <= (layer2_outputs(175)) xor (layer2_outputs(1242));
    outputs(2289) <= not(layer2_outputs(4206));
    outputs(2290) <= layer2_outputs(1323);
    outputs(2291) <= not(layer2_outputs(1151)) or (layer2_outputs(2095));
    outputs(2292) <= not(layer2_outputs(5075));
    outputs(2293) <= (layer2_outputs(3638)) xor (layer2_outputs(1985));
    outputs(2294) <= layer2_outputs(3551);
    outputs(2295) <= not((layer2_outputs(4831)) and (layer2_outputs(4849)));
    outputs(2296) <= not(layer2_outputs(2767));
    outputs(2297) <= not(layer2_outputs(4428));
    outputs(2298) <= not((layer2_outputs(881)) xor (layer2_outputs(4284)));
    outputs(2299) <= not((layer2_outputs(4950)) or (layer2_outputs(1786)));
    outputs(2300) <= not(layer2_outputs(2348));
    outputs(2301) <= layer2_outputs(3270);
    outputs(2302) <= (layer2_outputs(4912)) and not (layer2_outputs(912));
    outputs(2303) <= layer2_outputs(774);
    outputs(2304) <= not(layer2_outputs(4116));
    outputs(2305) <= not((layer2_outputs(157)) xor (layer2_outputs(3517)));
    outputs(2306) <= not(layer2_outputs(1868));
    outputs(2307) <= (layer2_outputs(1702)) and (layer2_outputs(4725));
    outputs(2308) <= not((layer2_outputs(3478)) xor (layer2_outputs(3032)));
    outputs(2309) <= not(layer2_outputs(2004));
    outputs(2310) <= not(layer2_outputs(4412));
    outputs(2311) <= not(layer2_outputs(1761));
    outputs(2312) <= not(layer2_outputs(2363));
    outputs(2313) <= layer2_outputs(3659);
    outputs(2314) <= (layer2_outputs(2144)) and (layer2_outputs(887));
    outputs(2315) <= (layer2_outputs(114)) and not (layer2_outputs(3390));
    outputs(2316) <= (layer2_outputs(2642)) xor (layer2_outputs(597));
    outputs(2317) <= not(layer2_outputs(3519));
    outputs(2318) <= (layer2_outputs(550)) xor (layer2_outputs(1927));
    outputs(2319) <= not(layer2_outputs(3256));
    outputs(2320) <= (layer2_outputs(1481)) and not (layer2_outputs(373));
    outputs(2321) <= not(layer2_outputs(2334));
    outputs(2322) <= not(layer2_outputs(837));
    outputs(2323) <= not((layer2_outputs(1519)) xor (layer2_outputs(4828)));
    outputs(2324) <= layer2_outputs(1826);
    outputs(2325) <= layer2_outputs(2647);
    outputs(2326) <= (layer2_outputs(351)) xor (layer2_outputs(3729));
    outputs(2327) <= not(layer2_outputs(3030));
    outputs(2328) <= not(layer2_outputs(4737));
    outputs(2329) <= not(layer2_outputs(2668));
    outputs(2330) <= layer2_outputs(4833);
    outputs(2331) <= not(layer2_outputs(2913));
    outputs(2332) <= layer2_outputs(2818);
    outputs(2333) <= not(layer2_outputs(3107)) or (layer2_outputs(1026));
    outputs(2334) <= not(layer2_outputs(2692));
    outputs(2335) <= layer2_outputs(791);
    outputs(2336) <= layer2_outputs(1389);
    outputs(2337) <= layer2_outputs(4350);
    outputs(2338) <= layer2_outputs(521);
    outputs(2339) <= not(layer2_outputs(2040));
    outputs(2340) <= layer2_outputs(1596);
    outputs(2341) <= not(layer2_outputs(3377));
    outputs(2342) <= not(layer2_outputs(625));
    outputs(2343) <= (layer2_outputs(5023)) and (layer2_outputs(2584));
    outputs(2344) <= not((layer2_outputs(1643)) xor (layer2_outputs(3040)));
    outputs(2345) <= not(layer2_outputs(4212)) or (layer2_outputs(1834));
    outputs(2346) <= (layer2_outputs(1426)) and not (layer2_outputs(1423));
    outputs(2347) <= (layer2_outputs(1461)) and (layer2_outputs(4103));
    outputs(2348) <= not(layer2_outputs(2551));
    outputs(2349) <= not(layer2_outputs(335)) or (layer2_outputs(2760));
    outputs(2350) <= not(layer2_outputs(4831));
    outputs(2351) <= layer2_outputs(249);
    outputs(2352) <= (layer2_outputs(1923)) and not (layer2_outputs(1214));
    outputs(2353) <= not(layer2_outputs(2314)) or (layer2_outputs(1482));
    outputs(2354) <= (layer2_outputs(2752)) and (layer2_outputs(133));
    outputs(2355) <= not(layer2_outputs(2435));
    outputs(2356) <= not(layer2_outputs(960)) or (layer2_outputs(605));
    outputs(2357) <= '0';
    outputs(2358) <= layer2_outputs(4225);
    outputs(2359) <= layer2_outputs(5067);
    outputs(2360) <= not((layer2_outputs(2342)) xor (layer2_outputs(1663)));
    outputs(2361) <= not((layer2_outputs(2371)) xor (layer2_outputs(829)));
    outputs(2362) <= (layer2_outputs(1303)) and not (layer2_outputs(4357));
    outputs(2363) <= (layer2_outputs(2459)) and (layer2_outputs(1852));
    outputs(2364) <= not(layer2_outputs(1417));
    outputs(2365) <= not(layer2_outputs(3212));
    outputs(2366) <= not(layer2_outputs(4439));
    outputs(2367) <= (layer2_outputs(2532)) xor (layer2_outputs(237));
    outputs(2368) <= not((layer2_outputs(4390)) or (layer2_outputs(1490)));
    outputs(2369) <= (layer2_outputs(2394)) and not (layer2_outputs(3050));
    outputs(2370) <= not(layer2_outputs(1878));
    outputs(2371) <= (layer2_outputs(2978)) and (layer2_outputs(3571));
    outputs(2372) <= layer2_outputs(4670);
    outputs(2373) <= (layer2_outputs(1454)) xor (layer2_outputs(1261));
    outputs(2374) <= not((layer2_outputs(543)) xor (layer2_outputs(4982)));
    outputs(2375) <= not(layer2_outputs(4100));
    outputs(2376) <= layer2_outputs(727);
    outputs(2377) <= not(layer2_outputs(3847));
    outputs(2378) <= not(layer2_outputs(2937));
    outputs(2379) <= layer2_outputs(365);
    outputs(2380) <= not(layer2_outputs(3115));
    outputs(2381) <= layer2_outputs(1887);
    outputs(2382) <= (layer2_outputs(4463)) xor (layer2_outputs(1578));
    outputs(2383) <= not((layer2_outputs(2675)) and (layer2_outputs(176)));
    outputs(2384) <= not(layer2_outputs(2093));
    outputs(2385) <= layer2_outputs(3888);
    outputs(2386) <= layer2_outputs(2281);
    outputs(2387) <= layer2_outputs(3269);
    outputs(2388) <= not(layer2_outputs(3096));
    outputs(2389) <= not(layer2_outputs(2507));
    outputs(2390) <= not(layer2_outputs(1155));
    outputs(2391) <= not(layer2_outputs(909));
    outputs(2392) <= not(layer2_outputs(2925));
    outputs(2393) <= (layer2_outputs(3179)) xor (layer2_outputs(2825));
    outputs(2394) <= layer2_outputs(1033);
    outputs(2395) <= not((layer2_outputs(3450)) and (layer2_outputs(2081)));
    outputs(2396) <= not(layer2_outputs(1304));
    outputs(2397) <= layer2_outputs(470);
    outputs(2398) <= not(layer2_outputs(3797));
    outputs(2399) <= not(layer2_outputs(1077));
    outputs(2400) <= (layer2_outputs(1242)) and not (layer2_outputs(2044));
    outputs(2401) <= layer2_outputs(222);
    outputs(2402) <= layer2_outputs(4876);
    outputs(2403) <= not(layer2_outputs(1051)) or (layer2_outputs(3068));
    outputs(2404) <= (layer2_outputs(4464)) xor (layer2_outputs(1766));
    outputs(2405) <= (layer2_outputs(3157)) and (layer2_outputs(2079));
    outputs(2406) <= not(layer2_outputs(1733));
    outputs(2407) <= not(layer2_outputs(4940));
    outputs(2408) <= (layer2_outputs(4670)) and not (layer2_outputs(2418));
    outputs(2409) <= layer2_outputs(153);
    outputs(2410) <= not(layer2_outputs(878));
    outputs(2411) <= layer2_outputs(1907);
    outputs(2412) <= layer2_outputs(936);
    outputs(2413) <= not((layer2_outputs(3064)) or (layer2_outputs(764)));
    outputs(2414) <= not(layer2_outputs(3106));
    outputs(2415) <= layer2_outputs(1053);
    outputs(2416) <= layer2_outputs(49);
    outputs(2417) <= layer2_outputs(4561);
    outputs(2418) <= (layer2_outputs(703)) and not (layer2_outputs(4674));
    outputs(2419) <= (layer2_outputs(2182)) and not (layer2_outputs(448));
    outputs(2420) <= not(layer2_outputs(3145));
    outputs(2421) <= not(layer2_outputs(558));
    outputs(2422) <= not((layer2_outputs(35)) xor (layer2_outputs(1899)));
    outputs(2423) <= not((layer2_outputs(3085)) xor (layer2_outputs(3509)));
    outputs(2424) <= layer2_outputs(733);
    outputs(2425) <= not(layer2_outputs(1494));
    outputs(2426) <= not(layer2_outputs(2629));
    outputs(2427) <= not(layer2_outputs(395));
    outputs(2428) <= layer2_outputs(1799);
    outputs(2429) <= not(layer2_outputs(623));
    outputs(2430) <= layer2_outputs(3600);
    outputs(2431) <= layer2_outputs(1099);
    outputs(2432) <= layer2_outputs(2789);
    outputs(2433) <= not(layer2_outputs(2754));
    outputs(2434) <= not(layer2_outputs(4298)) or (layer2_outputs(2140));
    outputs(2435) <= layer2_outputs(1408);
    outputs(2436) <= not(layer2_outputs(3493));
    outputs(2437) <= not(layer2_outputs(583)) or (layer2_outputs(3634));
    outputs(2438) <= layer2_outputs(4986);
    outputs(2439) <= not(layer2_outputs(4469));
    outputs(2440) <= layer2_outputs(4561);
    outputs(2441) <= layer2_outputs(481);
    outputs(2442) <= not(layer2_outputs(3630));
    outputs(2443) <= layer2_outputs(4833);
    outputs(2444) <= not(layer2_outputs(3310));
    outputs(2445) <= not(layer2_outputs(1590));
    outputs(2446) <= layer2_outputs(458);
    outputs(2447) <= (layer2_outputs(1032)) xor (layer2_outputs(3910));
    outputs(2448) <= not(layer2_outputs(1326));
    outputs(2449) <= not((layer2_outputs(2125)) and (layer2_outputs(3889)));
    outputs(2450) <= layer2_outputs(2822);
    outputs(2451) <= (layer2_outputs(1413)) xor (layer2_outputs(2328));
    outputs(2452) <= not(layer2_outputs(4621));
    outputs(2453) <= '1';
    outputs(2454) <= (layer2_outputs(4515)) and not (layer2_outputs(4124));
    outputs(2455) <= not(layer2_outputs(2603));
    outputs(2456) <= (layer2_outputs(1416)) xor (layer2_outputs(1718));
    outputs(2457) <= layer2_outputs(370);
    outputs(2458) <= (layer2_outputs(1433)) xor (layer2_outputs(983));
    outputs(2459) <= (layer2_outputs(1085)) and not (layer2_outputs(3090));
    outputs(2460) <= not(layer2_outputs(3905));
    outputs(2461) <= layer2_outputs(2844);
    outputs(2462) <= layer2_outputs(3434);
    outputs(2463) <= layer2_outputs(3324);
    outputs(2464) <= not(layer2_outputs(2521));
    outputs(2465) <= (layer2_outputs(3570)) and not (layer2_outputs(3852));
    outputs(2466) <= layer2_outputs(40);
    outputs(2467) <= not((layer2_outputs(4523)) and (layer2_outputs(3568)));
    outputs(2468) <= layer2_outputs(3163);
    outputs(2469) <= layer2_outputs(4510);
    outputs(2470) <= not(layer2_outputs(4937));
    outputs(2471) <= layer2_outputs(4432);
    outputs(2472) <= layer2_outputs(1291);
    outputs(2473) <= not(layer2_outputs(1516)) or (layer2_outputs(5008));
    outputs(2474) <= layer2_outputs(5066);
    outputs(2475) <= not((layer2_outputs(4571)) xor (layer2_outputs(2869)));
    outputs(2476) <= (layer2_outputs(4767)) xor (layer2_outputs(60));
    outputs(2477) <= layer2_outputs(1974);
    outputs(2478) <= not(layer2_outputs(1191));
    outputs(2479) <= (layer2_outputs(3054)) and not (layer2_outputs(909));
    outputs(2480) <= (layer2_outputs(2638)) and (layer2_outputs(3335));
    outputs(2481) <= (layer2_outputs(296)) xor (layer2_outputs(1329));
    outputs(2482) <= (layer2_outputs(2781)) and not (layer2_outputs(4611));
    outputs(2483) <= not(layer2_outputs(2661));
    outputs(2484) <= not(layer2_outputs(1673));
    outputs(2485) <= not(layer2_outputs(53));
    outputs(2486) <= (layer2_outputs(1320)) or (layer2_outputs(1288));
    outputs(2487) <= (layer2_outputs(502)) xor (layer2_outputs(3973));
    outputs(2488) <= not((layer2_outputs(1904)) or (layer2_outputs(4208)));
    outputs(2489) <= layer2_outputs(2957);
    outputs(2490) <= not((layer2_outputs(2998)) and (layer2_outputs(741)));
    outputs(2491) <= not(layer2_outputs(3721));
    outputs(2492) <= layer2_outputs(987);
    outputs(2493) <= layer2_outputs(3935);
    outputs(2494) <= not((layer2_outputs(1697)) xor (layer2_outputs(3130)));
    outputs(2495) <= not((layer2_outputs(4457)) or (layer2_outputs(1941)));
    outputs(2496) <= not(layer2_outputs(2287));
    outputs(2497) <= not(layer2_outputs(1843));
    outputs(2498) <= layer2_outputs(3596);
    outputs(2499) <= (layer2_outputs(4308)) or (layer2_outputs(4604));
    outputs(2500) <= not((layer2_outputs(1232)) or (layer2_outputs(48)));
    outputs(2501) <= not(layer2_outputs(4038));
    outputs(2502) <= (layer2_outputs(2191)) and not (layer2_outputs(593));
    outputs(2503) <= layer2_outputs(2116);
    outputs(2504) <= (layer2_outputs(5027)) and not (layer2_outputs(3971));
    outputs(2505) <= layer2_outputs(1667);
    outputs(2506) <= not(layer2_outputs(4844));
    outputs(2507) <= (layer2_outputs(4010)) xor (layer2_outputs(364));
    outputs(2508) <= not(layer2_outputs(2506));
    outputs(2509) <= not((layer2_outputs(5077)) xor (layer2_outputs(663)));
    outputs(2510) <= layer2_outputs(4686);
    outputs(2511) <= (layer2_outputs(3749)) xor (layer2_outputs(2942));
    outputs(2512) <= not(layer2_outputs(1146));
    outputs(2513) <= not(layer2_outputs(136)) or (layer2_outputs(5012));
    outputs(2514) <= (layer2_outputs(112)) xor (layer2_outputs(935));
    outputs(2515) <= (layer2_outputs(2166)) and (layer2_outputs(4978));
    outputs(2516) <= not(layer2_outputs(3986));
    outputs(2517) <= not((layer2_outputs(3518)) or (layer2_outputs(202)));
    outputs(2518) <= not(layer2_outputs(3402));
    outputs(2519) <= not(layer2_outputs(2617));
    outputs(2520) <= layer2_outputs(2185);
    outputs(2521) <= layer2_outputs(4436);
    outputs(2522) <= (layer2_outputs(4433)) xor (layer2_outputs(523));
    outputs(2523) <= layer2_outputs(1920);
    outputs(2524) <= (layer2_outputs(2588)) xor (layer2_outputs(2657));
    outputs(2525) <= layer2_outputs(3941);
    outputs(2526) <= (layer2_outputs(2598)) and (layer2_outputs(4146));
    outputs(2527) <= not(layer2_outputs(980));
    outputs(2528) <= not(layer2_outputs(1979));
    outputs(2529) <= (layer2_outputs(4491)) and (layer2_outputs(424));
    outputs(2530) <= (layer2_outputs(4070)) and not (layer2_outputs(1793));
    outputs(2531) <= layer2_outputs(703);
    outputs(2532) <= not(layer2_outputs(1028));
    outputs(2533) <= layer2_outputs(2414);
    outputs(2534) <= not(layer2_outputs(594));
    outputs(2535) <= (layer2_outputs(3845)) xor (layer2_outputs(1782));
    outputs(2536) <= (layer2_outputs(4158)) and not (layer2_outputs(561));
    outputs(2537) <= not((layer2_outputs(1253)) xor (layer2_outputs(4018)));
    outputs(2538) <= not(layer2_outputs(3809));
    outputs(2539) <= (layer2_outputs(996)) xor (layer2_outputs(220));
    outputs(2540) <= layer2_outputs(4535);
    outputs(2541) <= not(layer2_outputs(499));
    outputs(2542) <= not(layer2_outputs(905));
    outputs(2543) <= not(layer2_outputs(353));
    outputs(2544) <= (layer2_outputs(3737)) and not (layer2_outputs(5033));
    outputs(2545) <= layer2_outputs(4970);
    outputs(2546) <= layer2_outputs(4098);
    outputs(2547) <= not(layer2_outputs(2437));
    outputs(2548) <= layer2_outputs(627);
    outputs(2549) <= not(layer2_outputs(3592));
    outputs(2550) <= not(layer2_outputs(4896));
    outputs(2551) <= layer2_outputs(1378);
    outputs(2552) <= layer2_outputs(165);
    outputs(2553) <= layer2_outputs(1794);
    outputs(2554) <= not((layer2_outputs(3098)) xor (layer2_outputs(3972)));
    outputs(2555) <= not(layer2_outputs(2407));
    outputs(2556) <= not(layer2_outputs(775));
    outputs(2557) <= layer2_outputs(2266);
    outputs(2558) <= layer2_outputs(4604);
    outputs(2559) <= layer2_outputs(4919);
    outputs(2560) <= not((layer2_outputs(1749)) xor (layer2_outputs(1528)));
    outputs(2561) <= not(layer2_outputs(860));
    outputs(2562) <= layer2_outputs(3355);
    outputs(2563) <= not((layer2_outputs(3491)) xor (layer2_outputs(167)));
    outputs(2564) <= not(layer2_outputs(4694)) or (layer2_outputs(101));
    outputs(2565) <= (layer2_outputs(1422)) or (layer2_outputs(1607));
    outputs(2566) <= layer2_outputs(1104);
    outputs(2567) <= not(layer2_outputs(251));
    outputs(2568) <= (layer2_outputs(5094)) and (layer2_outputs(3372));
    outputs(2569) <= (layer2_outputs(1711)) and not (layer2_outputs(3025));
    outputs(2570) <= not(layer2_outputs(895));
    outputs(2571) <= layer2_outputs(1720);
    outputs(2572) <= (layer2_outputs(4554)) or (layer2_outputs(3718));
    outputs(2573) <= layer2_outputs(2965);
    outputs(2574) <= not(layer2_outputs(1463));
    outputs(2575) <= not(layer2_outputs(1226));
    outputs(2576) <= layer2_outputs(4113);
    outputs(2577) <= not(layer2_outputs(2696));
    outputs(2578) <= not(layer2_outputs(824));
    outputs(2579) <= (layer2_outputs(4001)) and not (layer2_outputs(415));
    outputs(2580) <= not((layer2_outputs(982)) xor (layer2_outputs(1760)));
    outputs(2581) <= layer2_outputs(3389);
    outputs(2582) <= layer2_outputs(117);
    outputs(2583) <= not(layer2_outputs(3748));
    outputs(2584) <= layer2_outputs(223);
    outputs(2585) <= layer2_outputs(1104);
    outputs(2586) <= layer2_outputs(4328);
    outputs(2587) <= not(layer2_outputs(3544));
    outputs(2588) <= layer2_outputs(995);
    outputs(2589) <= not(layer2_outputs(1052));
    outputs(2590) <= not((layer2_outputs(1246)) xor (layer2_outputs(3051)));
    outputs(2591) <= (layer2_outputs(4170)) xor (layer2_outputs(3178));
    outputs(2592) <= not(layer2_outputs(1367));
    outputs(2593) <= not(layer2_outputs(5014)) or (layer2_outputs(4219));
    outputs(2594) <= not(layer2_outputs(291));
    outputs(2595) <= layer2_outputs(2017);
    outputs(2596) <= not(layer2_outputs(3880));
    outputs(2597) <= not(layer2_outputs(318));
    outputs(2598) <= not((layer2_outputs(902)) and (layer2_outputs(4338)));
    outputs(2599) <= not(layer2_outputs(3560));
    outputs(2600) <= not(layer2_outputs(33));
    outputs(2601) <= (layer2_outputs(2452)) or (layer2_outputs(4525));
    outputs(2602) <= not(layer2_outputs(1246));
    outputs(2603) <= layer2_outputs(3537);
    outputs(2604) <= not(layer2_outputs(1684));
    outputs(2605) <= not((layer2_outputs(52)) xor (layer2_outputs(4198)));
    outputs(2606) <= (layer2_outputs(1551)) xor (layer2_outputs(640));
    outputs(2607) <= layer2_outputs(37);
    outputs(2608) <= layer2_outputs(684);
    outputs(2609) <= layer2_outputs(1199);
    outputs(2610) <= not(layer2_outputs(413));
    outputs(2611) <= (layer2_outputs(3888)) xor (layer2_outputs(403));
    outputs(2612) <= layer2_outputs(1526);
    outputs(2613) <= (layer2_outputs(5098)) and not (layer2_outputs(3902));
    outputs(2614) <= not(layer2_outputs(862));
    outputs(2615) <= not(layer2_outputs(4827)) or (layer2_outputs(2477));
    outputs(2616) <= (layer2_outputs(1464)) and not (layer2_outputs(695));
    outputs(2617) <= not(layer2_outputs(1535));
    outputs(2618) <= not(layer2_outputs(2833));
    outputs(2619) <= (layer2_outputs(588)) and not (layer2_outputs(1596));
    outputs(2620) <= not((layer2_outputs(1975)) xor (layer2_outputs(2331)));
    outputs(2621) <= not(layer2_outputs(611));
    outputs(2622) <= not((layer2_outputs(420)) xor (layer2_outputs(4333)));
    outputs(2623) <= (layer2_outputs(1587)) xor (layer2_outputs(973));
    outputs(2624) <= not((layer2_outputs(1514)) and (layer2_outputs(524)));
    outputs(2625) <= layer2_outputs(576);
    outputs(2626) <= layer2_outputs(4490);
    outputs(2627) <= layer2_outputs(3078);
    outputs(2628) <= (layer2_outputs(4530)) and not (layer2_outputs(4397));
    outputs(2629) <= not((layer2_outputs(3057)) xor (layer2_outputs(2682)));
    outputs(2630) <= (layer2_outputs(2839)) and (layer2_outputs(4111));
    outputs(2631) <= not(layer2_outputs(1497));
    outputs(2632) <= (layer2_outputs(2841)) and (layer2_outputs(2983));
    outputs(2633) <= layer2_outputs(4750);
    outputs(2634) <= (layer2_outputs(4013)) xor (layer2_outputs(3866));
    outputs(2635) <= not(layer2_outputs(4951));
    outputs(2636) <= not(layer2_outputs(1504));
    outputs(2637) <= layer2_outputs(3129);
    outputs(2638) <= (layer2_outputs(1739)) and not (layer2_outputs(1508));
    outputs(2639) <= (layer2_outputs(3511)) or (layer2_outputs(682));
    outputs(2640) <= layer2_outputs(3220);
    outputs(2641) <= (layer2_outputs(596)) or (layer2_outputs(1844));
    outputs(2642) <= layer2_outputs(1055);
    outputs(2643) <= layer2_outputs(2791);
    outputs(2644) <= not((layer2_outputs(1576)) xor (layer2_outputs(267)));
    outputs(2645) <= not((layer2_outputs(2921)) and (layer2_outputs(274)));
    outputs(2646) <= layer2_outputs(701);
    outputs(2647) <= not(layer2_outputs(3951)) or (layer2_outputs(4320));
    outputs(2648) <= layer2_outputs(3485);
    outputs(2649) <= (layer2_outputs(3918)) and (layer2_outputs(4711));
    outputs(2650) <= not((layer2_outputs(2245)) xor (layer2_outputs(343)));
    outputs(2651) <= not(layer2_outputs(2274));
    outputs(2652) <= (layer2_outputs(3123)) or (layer2_outputs(1704));
    outputs(2653) <= (layer2_outputs(2161)) xor (layer2_outputs(4323));
    outputs(2654) <= (layer2_outputs(2117)) and not (layer2_outputs(363));
    outputs(2655) <= not(layer2_outputs(4529));
    outputs(2656) <= (layer2_outputs(2557)) and (layer2_outputs(1049));
    outputs(2657) <= (layer2_outputs(140)) and not (layer2_outputs(2028));
    outputs(2658) <= not(layer2_outputs(4183));
    outputs(2659) <= not(layer2_outputs(3386));
    outputs(2660) <= not((layer2_outputs(406)) or (layer2_outputs(141)));
    outputs(2661) <= layer2_outputs(3348);
    outputs(2662) <= not(layer2_outputs(1537));
    outputs(2663) <= not((layer2_outputs(1753)) or (layer2_outputs(1940)));
    outputs(2664) <= (layer2_outputs(4190)) or (layer2_outputs(1788));
    outputs(2665) <= not(layer2_outputs(608));
    outputs(2666) <= layer2_outputs(216);
    outputs(2667) <= not(layer2_outputs(2109));
    outputs(2668) <= (layer2_outputs(1093)) xor (layer2_outputs(988));
    outputs(2669) <= (layer2_outputs(4532)) and not (layer2_outputs(2256));
    outputs(2670) <= not(layer2_outputs(271)) or (layer2_outputs(2937));
    outputs(2671) <= layer2_outputs(2132);
    outputs(2672) <= (layer2_outputs(4104)) and (layer2_outputs(4102));
    outputs(2673) <= not(layer2_outputs(3118));
    outputs(2674) <= not(layer2_outputs(1089));
    outputs(2675) <= layer2_outputs(1926);
    outputs(2676) <= not(layer2_outputs(3105));
    outputs(2677) <= layer2_outputs(2409);
    outputs(2678) <= (layer2_outputs(1516)) and not (layer2_outputs(2002));
    outputs(2679) <= not((layer2_outputs(2901)) or (layer2_outputs(3172)));
    outputs(2680) <= not(layer2_outputs(4768));
    outputs(2681) <= not(layer2_outputs(2411)) or (layer2_outputs(2941));
    outputs(2682) <= not(layer2_outputs(1723));
    outputs(2683) <= layer2_outputs(2703);
    outputs(2684) <= not(layer2_outputs(4484));
    outputs(2685) <= layer2_outputs(4904);
    outputs(2686) <= not(layer2_outputs(2406));
    outputs(2687) <= not(layer2_outputs(2919)) or (layer2_outputs(38));
    outputs(2688) <= not(layer2_outputs(5007));
    outputs(2689) <= not((layer2_outputs(38)) xor (layer2_outputs(693)));
    outputs(2690) <= layer2_outputs(4459);
    outputs(2691) <= (layer2_outputs(2538)) and not (layer2_outputs(806));
    outputs(2692) <= layer2_outputs(2894);
    outputs(2693) <= layer2_outputs(3150);
    outputs(2694) <= not(layer2_outputs(3960));
    outputs(2695) <= not((layer2_outputs(3732)) xor (layer2_outputs(4862)));
    outputs(2696) <= layer2_outputs(2614);
    outputs(2697) <= not(layer2_outputs(2313));
    outputs(2698) <= (layer2_outputs(411)) xor (layer2_outputs(2509));
    outputs(2699) <= not((layer2_outputs(4760)) xor (layer2_outputs(3746)));
    outputs(2700) <= not(layer2_outputs(3075));
    outputs(2701) <= (layer2_outputs(1987)) xor (layer2_outputs(4693));
    outputs(2702) <= (layer2_outputs(1334)) xor (layer2_outputs(981));
    outputs(2703) <= layer2_outputs(1995);
    outputs(2704) <= layer2_outputs(2123);
    outputs(2705) <= not(layer2_outputs(1806));
    outputs(2706) <= not((layer2_outputs(2994)) xor (layer2_outputs(4532)));
    outputs(2707) <= (layer2_outputs(1223)) and (layer2_outputs(1638));
    outputs(2708) <= not((layer2_outputs(4713)) xor (layer2_outputs(4240)));
    outputs(2709) <= (layer2_outputs(3511)) or (layer2_outputs(1174));
    outputs(2710) <= not(layer2_outputs(3265));
    outputs(2711) <= (layer2_outputs(1463)) xor (layer2_outputs(4905));
    outputs(2712) <= not(layer2_outputs(1273));
    outputs(2713) <= not(layer2_outputs(30));
    outputs(2714) <= layer2_outputs(2285);
    outputs(2715) <= not((layer2_outputs(414)) or (layer2_outputs(1165)));
    outputs(2716) <= not((layer2_outputs(1472)) xor (layer2_outputs(869)));
    outputs(2717) <= not(layer2_outputs(1605));
    outputs(2718) <= not(layer2_outputs(762));
    outputs(2719) <= not(layer2_outputs(4771));
    outputs(2720) <= (layer2_outputs(2504)) and (layer2_outputs(4152));
    outputs(2721) <= layer2_outputs(4898);
    outputs(2722) <= layer2_outputs(965);
    outputs(2723) <= not((layer2_outputs(2645)) and (layer2_outputs(3999)));
    outputs(2724) <= (layer2_outputs(1313)) xor (layer2_outputs(2663));
    outputs(2725) <= not((layer2_outputs(2140)) or (layer2_outputs(851)));
    outputs(2726) <= not((layer2_outputs(4052)) xor (layer2_outputs(2831)));
    outputs(2727) <= not(layer2_outputs(375));
    outputs(2728) <= not(layer2_outputs(1930));
    outputs(2729) <= not(layer2_outputs(3593));
    outputs(2730) <= layer2_outputs(3180);
    outputs(2731) <= not(layer2_outputs(3198));
    outputs(2732) <= layer2_outputs(2043);
    outputs(2733) <= not((layer2_outputs(3513)) xor (layer2_outputs(977)));
    outputs(2734) <= layer2_outputs(1771);
    outputs(2735) <= layer2_outputs(111);
    outputs(2736) <= not(layer2_outputs(1985)) or (layer2_outputs(5033));
    outputs(2737) <= (layer2_outputs(1858)) and (layer2_outputs(3088));
    outputs(2738) <= layer2_outputs(4620);
    outputs(2739) <= layer2_outputs(32);
    outputs(2740) <= not(layer2_outputs(4538));
    outputs(2741) <= not(layer2_outputs(5034));
    outputs(2742) <= not(layer2_outputs(2963));
    outputs(2743) <= layer2_outputs(4511);
    outputs(2744) <= (layer2_outputs(4878)) and (layer2_outputs(2906));
    outputs(2745) <= (layer2_outputs(2351)) and not (layer2_outputs(2553));
    outputs(2746) <= (layer2_outputs(2042)) and not (layer2_outputs(1411));
    outputs(2747) <= not(layer2_outputs(2006));
    outputs(2748) <= not(layer2_outputs(1850)) or (layer2_outputs(4973));
    outputs(2749) <= not(layer2_outputs(3776));
    outputs(2750) <= (layer2_outputs(5046)) xor (layer2_outputs(4385));
    outputs(2751) <= not((layer2_outputs(1114)) xor (layer2_outputs(4295)));
    outputs(2752) <= layer2_outputs(2783);
    outputs(2753) <= not((layer2_outputs(1059)) xor (layer2_outputs(3319)));
    outputs(2754) <= not(layer2_outputs(1814));
    outputs(2755) <= (layer2_outputs(1517)) xor (layer2_outputs(700));
    outputs(2756) <= not(layer2_outputs(425));
    outputs(2757) <= not(layer2_outputs(600));
    outputs(2758) <= layer2_outputs(73);
    outputs(2759) <= layer2_outputs(2005);
    outputs(2760) <= not((layer2_outputs(2788)) xor (layer2_outputs(1859)));
    outputs(2761) <= not(layer2_outputs(3792));
    outputs(2762) <= layer2_outputs(3727);
    outputs(2763) <= not(layer2_outputs(2536));
    outputs(2764) <= not(layer2_outputs(4764));
    outputs(2765) <= not(layer2_outputs(5091));
    outputs(2766) <= not((layer2_outputs(2244)) xor (layer2_outputs(4926)));
    outputs(2767) <= (layer2_outputs(2720)) or (layer2_outputs(1372));
    outputs(2768) <= not((layer2_outputs(2548)) xor (layer2_outputs(1083)));
    outputs(2769) <= layer2_outputs(529);
    outputs(2770) <= layer2_outputs(2525);
    outputs(2771) <= layer2_outputs(1249);
    outputs(2772) <= layer2_outputs(2155);
    outputs(2773) <= not(layer2_outputs(2012));
    outputs(2774) <= layer2_outputs(731);
    outputs(2775) <= (layer2_outputs(831)) and not (layer2_outputs(3387));
    outputs(2776) <= layer2_outputs(5010);
    outputs(2777) <= layer2_outputs(777);
    outputs(2778) <= not((layer2_outputs(1933)) xor (layer2_outputs(1375)));
    outputs(2779) <= not(layer2_outputs(3371));
    outputs(2780) <= not(layer2_outputs(4354));
    outputs(2781) <= layer2_outputs(4329);
    outputs(2782) <= (layer2_outputs(22)) xor (layer2_outputs(429));
    outputs(2783) <= not(layer2_outputs(706));
    outputs(2784) <= not(layer2_outputs(3291));
    outputs(2785) <= layer2_outputs(1281);
    outputs(2786) <= (layer2_outputs(4667)) xor (layer2_outputs(4649));
    outputs(2787) <= not((layer2_outputs(2638)) xor (layer2_outputs(2068)));
    outputs(2788) <= not(layer2_outputs(2859));
    outputs(2789) <= not(layer2_outputs(4130)) or (layer2_outputs(997));
    outputs(2790) <= (layer2_outputs(2387)) or (layer2_outputs(3726));
    outputs(2791) <= (layer2_outputs(1305)) xor (layer2_outputs(4587));
    outputs(2792) <= layer2_outputs(3662);
    outputs(2793) <= (layer2_outputs(4447)) xor (layer2_outputs(4046));
    outputs(2794) <= layer2_outputs(5030);
    outputs(2795) <= layer2_outputs(2677);
    outputs(2796) <= layer2_outputs(5073);
    outputs(2797) <= not(layer2_outputs(583));
    outputs(2798) <= not((layer2_outputs(804)) xor (layer2_outputs(3834)));
    outputs(2799) <= layer2_outputs(3929);
    outputs(2800) <= (layer2_outputs(3446)) or (layer2_outputs(3589));
    outputs(2801) <= (layer2_outputs(1870)) and not (layer2_outputs(1441));
    outputs(2802) <= not(layer2_outputs(3265));
    outputs(2803) <= layer2_outputs(3224);
    outputs(2804) <= layer2_outputs(4738);
    outputs(2805) <= layer2_outputs(1669);
    outputs(2806) <= (layer2_outputs(4150)) xor (layer2_outputs(1465));
    outputs(2807) <= not(layer2_outputs(2258));
    outputs(2808) <= layer2_outputs(4552);
    outputs(2809) <= layer2_outputs(2195);
    outputs(2810) <= layer2_outputs(4380);
    outputs(2811) <= not((layer2_outputs(2835)) xor (layer2_outputs(397)));
    outputs(2812) <= not(layer2_outputs(3275));
    outputs(2813) <= (layer2_outputs(3780)) and (layer2_outputs(4965));
    outputs(2814) <= not(layer2_outputs(2622));
    outputs(2815) <= not(layer2_outputs(4563));
    outputs(2816) <= layer2_outputs(3475);
    outputs(2817) <= not(layer2_outputs(3354));
    outputs(2818) <= (layer2_outputs(1397)) xor (layer2_outputs(4424));
    outputs(2819) <= not(layer2_outputs(2567));
    outputs(2820) <= not((layer2_outputs(1419)) xor (layer2_outputs(230)));
    outputs(2821) <= layer2_outputs(1607);
    outputs(2822) <= layer2_outputs(2137);
    outputs(2823) <= not(layer2_outputs(44));
    outputs(2824) <= not(layer2_outputs(4087));
    outputs(2825) <= not(layer2_outputs(3560));
    outputs(2826) <= (layer2_outputs(3437)) xor (layer2_outputs(3015));
    outputs(2827) <= (layer2_outputs(4676)) or (layer2_outputs(3495));
    outputs(2828) <= not(layer2_outputs(1209));
    outputs(2829) <= not(layer2_outputs(3561));
    outputs(2830) <= layer2_outputs(2272);
    outputs(2831) <= not(layer2_outputs(1031)) or (layer2_outputs(3580));
    outputs(2832) <= layer2_outputs(3080);
    outputs(2833) <= layer2_outputs(2856);
    outputs(2834) <= layer2_outputs(5059);
    outputs(2835) <= layer2_outputs(3426);
    outputs(2836) <= not(layer2_outputs(4646));
    outputs(2837) <= not(layer2_outputs(3618));
    outputs(2838) <= (layer2_outputs(1407)) xor (layer2_outputs(571));
    outputs(2839) <= layer2_outputs(3297);
    outputs(2840) <= not(layer2_outputs(77));
    outputs(2841) <= not(layer2_outputs(822));
    outputs(2842) <= not(layer2_outputs(448));
    outputs(2843) <= layer2_outputs(931);
    outputs(2844) <= (layer2_outputs(4485)) xor (layer2_outputs(2737));
    outputs(2845) <= (layer2_outputs(3993)) xor (layer2_outputs(5043));
    outputs(2846) <= not(layer2_outputs(1853));
    outputs(2847) <= (layer2_outputs(1166)) xor (layer2_outputs(2320));
    outputs(2848) <= layer2_outputs(3416);
    outputs(2849) <= not((layer2_outputs(2219)) xor (layer2_outputs(949)));
    outputs(2850) <= not(layer2_outputs(848));
    outputs(2851) <= layer2_outputs(1799);
    outputs(2852) <= layer2_outputs(4223);
    outputs(2853) <= layer2_outputs(1245);
    outputs(2854) <= (layer2_outputs(1010)) and not (layer2_outputs(4399));
    outputs(2855) <= not((layer2_outputs(3650)) xor (layer2_outputs(4629)));
    outputs(2856) <= not(layer2_outputs(2932));
    outputs(2857) <= layer2_outputs(1617);
    outputs(2858) <= (layer2_outputs(972)) xor (layer2_outputs(3078));
    outputs(2859) <= not(layer2_outputs(4671));
    outputs(2860) <= not((layer2_outputs(1715)) or (layer2_outputs(2172)));
    outputs(2861) <= not(layer2_outputs(642));
    outputs(2862) <= not(layer2_outputs(2064));
    outputs(2863) <= (layer2_outputs(2298)) xor (layer2_outputs(4591));
    outputs(2864) <= not((layer2_outputs(650)) xor (layer2_outputs(2546)));
    outputs(2865) <= not(layer2_outputs(302));
    outputs(2866) <= layer2_outputs(3211);
    outputs(2867) <= not(layer2_outputs(3883));
    outputs(2868) <= (layer2_outputs(1686)) xor (layer2_outputs(5094));
    outputs(2869) <= not((layer2_outputs(4891)) and (layer2_outputs(2421)));
    outputs(2870) <= layer2_outputs(1518);
    outputs(2871) <= layer2_outputs(1713);
    outputs(2872) <= not(layer2_outputs(1625)) or (layer2_outputs(2644));
    outputs(2873) <= not((layer2_outputs(807)) xor (layer2_outputs(57)));
    outputs(2874) <= (layer2_outputs(3911)) xor (layer2_outputs(2063));
    outputs(2875) <= (layer2_outputs(1406)) xor (layer2_outputs(1815));
    outputs(2876) <= not(layer2_outputs(444));
    outputs(2877) <= layer2_outputs(1345);
    outputs(2878) <= layer2_outputs(3922);
    outputs(2879) <= not((layer2_outputs(2694)) xor (layer2_outputs(949)));
    outputs(2880) <= not(layer2_outputs(2229)) or (layer2_outputs(1677));
    outputs(2881) <= not((layer2_outputs(162)) xor (layer2_outputs(756)));
    outputs(2882) <= layer2_outputs(3933);
    outputs(2883) <= not((layer2_outputs(2200)) xor (layer2_outputs(3278)));
    outputs(2884) <= not(layer2_outputs(2751));
    outputs(2885) <= not((layer2_outputs(557)) xor (layer2_outputs(3491)));
    outputs(2886) <= not((layer2_outputs(3546)) xor (layer2_outputs(3059)));
    outputs(2887) <= layer2_outputs(1438);
    outputs(2888) <= not(layer2_outputs(2928));
    outputs(2889) <= (layer2_outputs(2343)) xor (layer2_outputs(121));
    outputs(2890) <= not((layer2_outputs(4473)) or (layer2_outputs(1319)));
    outputs(2891) <= not(layer2_outputs(2696));
    outputs(2892) <= (layer2_outputs(3967)) and not (layer2_outputs(5055));
    outputs(2893) <= not((layer2_outputs(3298)) xor (layer2_outputs(183)));
    outputs(2894) <= (layer2_outputs(393)) or (layer2_outputs(112));
    outputs(2895) <= (layer2_outputs(3622)) and not (layer2_outputs(1558));
    outputs(2896) <= layer2_outputs(4316);
    outputs(2897) <= not((layer2_outputs(5114)) and (layer2_outputs(4453)));
    outputs(2898) <= (layer2_outputs(1637)) and not (layer2_outputs(1548));
    outputs(2899) <= layer2_outputs(2874);
    outputs(2900) <= not(layer2_outputs(231)) or (layer2_outputs(4565));
    outputs(2901) <= (layer2_outputs(4884)) and (layer2_outputs(3271));
    outputs(2902) <= not((layer2_outputs(4108)) xor (layer2_outputs(3606)));
    outputs(2903) <= not(layer2_outputs(4232));
    outputs(2904) <= layer2_outputs(2940);
    outputs(2905) <= (layer2_outputs(4242)) and not (layer2_outputs(1816));
    outputs(2906) <= not((layer2_outputs(548)) xor (layer2_outputs(4050)));
    outputs(2907) <= not((layer2_outputs(1581)) or (layer2_outputs(508)));
    outputs(2908) <= (layer2_outputs(3949)) and not (layer2_outputs(4143));
    outputs(2909) <= not(layer2_outputs(1818));
    outputs(2910) <= (layer2_outputs(2399)) xor (layer2_outputs(4000));
    outputs(2911) <= layer2_outputs(1647);
    outputs(2912) <= not(layer2_outputs(3218));
    outputs(2913) <= (layer2_outputs(118)) xor (layer2_outputs(1332));
    outputs(2914) <= (layer2_outputs(3392)) xor (layer2_outputs(2743));
    outputs(2915) <= layer2_outputs(4791);
    outputs(2916) <= not((layer2_outputs(1042)) xor (layer2_outputs(4070)));
    outputs(2917) <= not(layer2_outputs(2962));
    outputs(2918) <= layer2_outputs(4025);
    outputs(2919) <= layer2_outputs(1623);
    outputs(2920) <= not(layer2_outputs(4267)) or (layer2_outputs(1249));
    outputs(2921) <= layer2_outputs(894);
    outputs(2922) <= not(layer2_outputs(1629)) or (layer2_outputs(560));
    outputs(2923) <= not(layer2_outputs(257));
    outputs(2924) <= not(layer2_outputs(72));
    outputs(2925) <= (layer2_outputs(1001)) or (layer2_outputs(3917));
    outputs(2926) <= not(layer2_outputs(1348)) or (layer2_outputs(2900));
    outputs(2927) <= not((layer2_outputs(2687)) xor (layer2_outputs(4882)));
    outputs(2928) <= layer2_outputs(1509);
    outputs(2929) <= (layer2_outputs(3755)) xor (layer2_outputs(3210));
    outputs(2930) <= (layer2_outputs(3791)) xor (layer2_outputs(264));
    outputs(2931) <= not(layer2_outputs(3));
    outputs(2932) <= layer2_outputs(2595);
    outputs(2933) <= not(layer2_outputs(2812));
    outputs(2934) <= (layer2_outputs(688)) and (layer2_outputs(892));
    outputs(2935) <= layer2_outputs(1798);
    outputs(2936) <= layer2_outputs(5084);
    outputs(2937) <= layer2_outputs(1944);
    outputs(2938) <= not((layer2_outputs(4645)) xor (layer2_outputs(1956)));
    outputs(2939) <= not((layer2_outputs(913)) or (layer2_outputs(2680)));
    outputs(2940) <= (layer2_outputs(1709)) and not (layer2_outputs(3514));
    outputs(2941) <= (layer2_outputs(2985)) xor (layer2_outputs(3847));
    outputs(2942) <= not((layer2_outputs(1042)) xor (layer2_outputs(3018)));
    outputs(2943) <= not(layer2_outputs(1646));
    outputs(2944) <= not(layer2_outputs(3333)) or (layer2_outputs(2739));
    outputs(2945) <= layer2_outputs(1619);
    outputs(2946) <= (layer2_outputs(3119)) or (layer2_outputs(5041));
    outputs(2947) <= not((layer2_outputs(4856)) xor (layer2_outputs(56)));
    outputs(2948) <= not(layer2_outputs(1768));
    outputs(2949) <= not(layer2_outputs(55)) or (layer2_outputs(4427));
    outputs(2950) <= not((layer2_outputs(4311)) xor (layer2_outputs(950)));
    outputs(2951) <= not(layer2_outputs(507));
    outputs(2952) <= (layer2_outputs(4795)) xor (layer2_outputs(2828));
    outputs(2953) <= not((layer2_outputs(1937)) or (layer2_outputs(2365)));
    outputs(2954) <= not(layer2_outputs(1594));
    outputs(2955) <= layer2_outputs(2882);
    outputs(2956) <= not(layer2_outputs(2806));
    outputs(2957) <= not((layer2_outputs(1385)) or (layer2_outputs(3237)));
    outputs(2958) <= layer2_outputs(928);
    outputs(2959) <= not(layer2_outputs(2314));
    outputs(2960) <= layer2_outputs(661);
    outputs(2961) <= layer2_outputs(2841);
    outputs(2962) <= layer2_outputs(1380);
    outputs(2963) <= not((layer2_outputs(833)) xor (layer2_outputs(2013)));
    outputs(2964) <= (layer2_outputs(2246)) xor (layer2_outputs(1875));
    outputs(2965) <= layer2_outputs(391);
    outputs(2966) <= (layer2_outputs(613)) xor (layer2_outputs(4493));
    outputs(2967) <= not((layer2_outputs(330)) and (layer2_outputs(1113)));
    outputs(2968) <= layer2_outputs(1394);
    outputs(2969) <= layer2_outputs(2447);
    outputs(2970) <= layer2_outputs(607);
    outputs(2971) <= layer2_outputs(4060);
    outputs(2972) <= not(layer2_outputs(81));
    outputs(2973) <= layer2_outputs(283);
    outputs(2974) <= not(layer2_outputs(3420));
    outputs(2975) <= not((layer2_outputs(3226)) or (layer2_outputs(1175)));
    outputs(2976) <= not(layer2_outputs(5103));
    outputs(2977) <= not((layer2_outputs(3330)) xor (layer2_outputs(3316)));
    outputs(2978) <= not((layer2_outputs(4923)) or (layer2_outputs(5103)));
    outputs(2979) <= not(layer2_outputs(3862));
    outputs(2980) <= not((layer2_outputs(4486)) xor (layer2_outputs(3839)));
    outputs(2981) <= (layer2_outputs(893)) xor (layer2_outputs(4141));
    outputs(2982) <= not(layer2_outputs(5049));
    outputs(2983) <= (layer2_outputs(3343)) xor (layer2_outputs(2625));
    outputs(2984) <= (layer2_outputs(137)) and not (layer2_outputs(4994));
    outputs(2985) <= not(layer2_outputs(354)) or (layer2_outputs(734));
    outputs(2986) <= not(layer2_outputs(459));
    outputs(2987) <= layer2_outputs(4410);
    outputs(2988) <= layer2_outputs(2473);
    outputs(2989) <= layer2_outputs(4942);
    outputs(2990) <= layer2_outputs(771);
    outputs(2991) <= layer2_outputs(613);
    outputs(2992) <= (layer2_outputs(2172)) xor (layer2_outputs(2327));
    outputs(2993) <= not((layer2_outputs(4057)) or (layer2_outputs(12)));
    outputs(2994) <= not((layer2_outputs(2189)) and (layer2_outputs(2534)));
    outputs(2995) <= not((layer2_outputs(246)) xor (layer2_outputs(1921)));
    outputs(2996) <= not(layer2_outputs(3329));
    outputs(2997) <= not(layer2_outputs(292));
    outputs(2998) <= (layer2_outputs(3370)) or (layer2_outputs(3255));
    outputs(2999) <= layer2_outputs(814);
    outputs(3000) <= (layer2_outputs(2861)) and not (layer2_outputs(2554));
    outputs(3001) <= (layer2_outputs(4110)) xor (layer2_outputs(3139));
    outputs(3002) <= not((layer2_outputs(421)) or (layer2_outputs(3849)));
    outputs(3003) <= not(layer2_outputs(335)) or (layer2_outputs(1001));
    outputs(3004) <= layer2_outputs(966);
    outputs(3005) <= (layer2_outputs(3425)) xor (layer2_outputs(2075));
    outputs(3006) <= layer2_outputs(255);
    outputs(3007) <= layer2_outputs(1877);
    outputs(3008) <= not(layer2_outputs(2253));
    outputs(3009) <= (layer2_outputs(4444)) or (layer2_outputs(190));
    outputs(3010) <= not(layer2_outputs(4176));
    outputs(3011) <= layer2_outputs(350);
    outputs(3012) <= not(layer2_outputs(1500));
    outputs(3013) <= not((layer2_outputs(2269)) and (layer2_outputs(2609)));
    outputs(3014) <= layer2_outputs(1669);
    outputs(3015) <= (layer2_outputs(4901)) or (layer2_outputs(5100));
    outputs(3016) <= layer2_outputs(53);
    outputs(3017) <= (layer2_outputs(4748)) xor (layer2_outputs(786));
    outputs(3018) <= (layer2_outputs(4418)) xor (layer2_outputs(1560));
    outputs(3019) <= (layer2_outputs(578)) xor (layer2_outputs(4325));
    outputs(3020) <= not((layer2_outputs(71)) or (layer2_outputs(3141)));
    outputs(3021) <= not(layer2_outputs(1925)) or (layer2_outputs(3154));
    outputs(3022) <= layer2_outputs(3327);
    outputs(3023) <= layer2_outputs(2723);
    outputs(3024) <= not(layer2_outputs(4825));
    outputs(3025) <= not((layer2_outputs(155)) xor (layer2_outputs(2016)));
    outputs(3026) <= (layer2_outputs(303)) and (layer2_outputs(1343));
    outputs(3027) <= layer2_outputs(3885);
    outputs(3028) <= not((layer2_outputs(3260)) xor (layer2_outputs(842)));
    outputs(3029) <= (layer2_outputs(2263)) xor (layer2_outputs(1325));
    outputs(3030) <= not(layer2_outputs(2360));
    outputs(3031) <= (layer2_outputs(3650)) xor (layer2_outputs(677));
    outputs(3032) <= not(layer2_outputs(3670)) or (layer2_outputs(4154));
    outputs(3033) <= not((layer2_outputs(1732)) xor (layer2_outputs(475)));
    outputs(3034) <= (layer2_outputs(3501)) and not (layer2_outputs(5052));
    outputs(3035) <= layer2_outputs(4466);
    outputs(3036) <= (layer2_outputs(604)) and not (layer2_outputs(545));
    outputs(3037) <= layer2_outputs(109);
    outputs(3038) <= (layer2_outputs(3132)) or (layer2_outputs(5000));
    outputs(3039) <= (layer2_outputs(1556)) or (layer2_outputs(1838));
    outputs(3040) <= not((layer2_outputs(1577)) or (layer2_outputs(1458)));
    outputs(3041) <= not((layer2_outputs(1106)) xor (layer2_outputs(2402)));
    outputs(3042) <= layer2_outputs(1024);
    outputs(3043) <= (layer2_outputs(1168)) or (layer2_outputs(1205));
    outputs(3044) <= not(layer2_outputs(4400));
    outputs(3045) <= (layer2_outputs(1072)) xor (layer2_outputs(4365));
    outputs(3046) <= not(layer2_outputs(5026));
    outputs(3047) <= not(layer2_outputs(99));
    outputs(3048) <= (layer2_outputs(3487)) and not (layer2_outputs(2897));
    outputs(3049) <= not(layer2_outputs(1980));
    outputs(3050) <= not(layer2_outputs(4301)) or (layer2_outputs(1168));
    outputs(3051) <= not((layer2_outputs(4312)) and (layer2_outputs(473)));
    outputs(3052) <= (layer2_outputs(4205)) xor (layer2_outputs(2171));
    outputs(3053) <= layer2_outputs(3599);
    outputs(3054) <= not(layer2_outputs(4101));
    outputs(3055) <= (layer2_outputs(1156)) and not (layer2_outputs(3828));
    outputs(3056) <= layer2_outputs(3716);
    outputs(3057) <= layer2_outputs(3631);
    outputs(3058) <= not(layer2_outputs(4880));
    outputs(3059) <= not(layer2_outputs(2217));
    outputs(3060) <= (layer2_outputs(273)) and not (layer2_outputs(3707));
    outputs(3061) <= layer2_outputs(3188);
    outputs(3062) <= (layer2_outputs(2112)) xor (layer2_outputs(2886));
    outputs(3063) <= layer2_outputs(3297);
    outputs(3064) <= not((layer2_outputs(897)) xor (layer2_outputs(4384)));
    outputs(3065) <= (layer2_outputs(2636)) xor (layer2_outputs(396));
    outputs(3066) <= (layer2_outputs(958)) xor (layer2_outputs(3692));
    outputs(3067) <= layer2_outputs(586);
    outputs(3068) <= not(layer2_outputs(2593));
    outputs(3069) <= layer2_outputs(2832);
    outputs(3070) <= not(layer2_outputs(258)) or (layer2_outputs(1274));
    outputs(3071) <= not((layer2_outputs(3326)) or (layer2_outputs(64)));
    outputs(3072) <= layer2_outputs(2148);
    outputs(3073) <= (layer2_outputs(1811)) xor (layer2_outputs(4113));
    outputs(3074) <= not(layer2_outputs(2722));
    outputs(3075) <= not((layer2_outputs(632)) xor (layer2_outputs(76)));
    outputs(3076) <= (layer2_outputs(5074)) xor (layer2_outputs(1279));
    outputs(3077) <= (layer2_outputs(4400)) and (layer2_outputs(1176));
    outputs(3078) <= layer2_outputs(5115);
    outputs(3079) <= (layer2_outputs(4953)) and (layer2_outputs(113));
    outputs(3080) <= not((layer2_outputs(546)) xor (layer2_outputs(4317)));
    outputs(3081) <= not(layer2_outputs(3459));
    outputs(3082) <= (layer2_outputs(2637)) and not (layer2_outputs(4803));
    outputs(3083) <= not(layer2_outputs(4988));
    outputs(3084) <= layer2_outputs(1278);
    outputs(3085) <= (layer2_outputs(1509)) xor (layer2_outputs(1619));
    outputs(3086) <= not(layer2_outputs(1508));
    outputs(3087) <= not(layer2_outputs(2049));
    outputs(3088) <= (layer2_outputs(4874)) or (layer2_outputs(4401));
    outputs(3089) <= layer2_outputs(2280);
    outputs(3090) <= not(layer2_outputs(3874));
    outputs(3091) <= (layer2_outputs(81)) xor (layer2_outputs(1885));
    outputs(3092) <= layer2_outputs(3074);
    outputs(3093) <= not((layer2_outputs(3891)) xor (layer2_outputs(4047)));
    outputs(3094) <= not((layer2_outputs(4945)) or (layer2_outputs(4317)));
    outputs(3095) <= not(layer2_outputs(3646)) or (layer2_outputs(4417));
    outputs(3096) <= not((layer2_outputs(3617)) xor (layer2_outputs(1270)));
    outputs(3097) <= not((layer2_outputs(2369)) and (layer2_outputs(4547)));
    outputs(3098) <= (layer2_outputs(2122)) xor (layer2_outputs(1179));
    outputs(3099) <= layer2_outputs(4064);
    outputs(3100) <= not((layer2_outputs(2217)) xor (layer2_outputs(2549)));
    outputs(3101) <= (layer2_outputs(2906)) or (layer2_outputs(159));
    outputs(3102) <= (layer2_outputs(4584)) and (layer2_outputs(4024));
    outputs(3103) <= layer2_outputs(2313);
    outputs(3104) <= (layer2_outputs(45)) xor (layer2_outputs(4063));
    outputs(3105) <= layer2_outputs(4038);
    outputs(3106) <= layer2_outputs(4927);
    outputs(3107) <= (layer2_outputs(940)) and not (layer2_outputs(4059));
    outputs(3108) <= not(layer2_outputs(349));
    outputs(3109) <= not(layer2_outputs(2759));
    outputs(3110) <= not(layer2_outputs(4768));
    outputs(3111) <= layer2_outputs(1603);
    outputs(3112) <= not(layer2_outputs(4028)) or (layer2_outputs(3418));
    outputs(3113) <= not((layer2_outputs(3606)) or (layer2_outputs(3892)));
    outputs(3114) <= not(layer2_outputs(1133));
    outputs(3115) <= not((layer2_outputs(1668)) or (layer2_outputs(3016)));
    outputs(3116) <= not(layer2_outputs(2795));
    outputs(3117) <= layer2_outputs(627);
    outputs(3118) <= layer2_outputs(3327);
    outputs(3119) <= layer2_outputs(1981);
    outputs(3120) <= (layer2_outputs(4445)) xor (layer2_outputs(4466));
    outputs(3121) <= layer2_outputs(654);
    outputs(3122) <= layer2_outputs(1232);
    outputs(3123) <= not(layer2_outputs(2358));
    outputs(3124) <= (layer2_outputs(4577)) and (layer2_outputs(308));
    outputs(3125) <= not(layer2_outputs(78));
    outputs(3126) <= (layer2_outputs(1480)) and not (layer2_outputs(725));
    outputs(3127) <= not(layer2_outputs(513));
    outputs(3128) <= (layer2_outputs(3300)) and (layer2_outputs(2684));
    outputs(3129) <= not(layer2_outputs(41)) or (layer2_outputs(1349));
    outputs(3130) <= (layer2_outputs(651)) and (layer2_outputs(4001));
    outputs(3131) <= not(layer2_outputs(423));
    outputs(3132) <= not(layer2_outputs(2196));
    outputs(3133) <= not((layer2_outputs(1122)) or (layer2_outputs(4005)));
    outputs(3134) <= not((layer2_outputs(4514)) or (layer2_outputs(2953)));
    outputs(3135) <= not(layer2_outputs(4747));
    outputs(3136) <= not(layer2_outputs(971));
    outputs(3137) <= not((layer2_outputs(3765)) or (layer2_outputs(4173)));
    outputs(3138) <= not((layer2_outputs(1178)) xor (layer2_outputs(1243)));
    outputs(3139) <= (layer2_outputs(2361)) and not (layer2_outputs(1396));
    outputs(3140) <= not(layer2_outputs(3423));
    outputs(3141) <= layer2_outputs(1855);
    outputs(3142) <= not(layer2_outputs(772));
    outputs(3143) <= layer2_outputs(4752);
    outputs(3144) <= layer2_outputs(2392);
    outputs(3145) <= layer2_outputs(2679);
    outputs(3146) <= layer2_outputs(672);
    outputs(3147) <= not(layer2_outputs(492));
    outputs(3148) <= not(layer2_outputs(2674));
    outputs(3149) <= layer2_outputs(1220);
    outputs(3150) <= layer2_outputs(1658);
    outputs(3151) <= (layer2_outputs(1004)) and (layer2_outputs(3945));
    outputs(3152) <= layer2_outputs(2444);
    outputs(3153) <= not(layer2_outputs(4570));
    outputs(3154) <= not(layer2_outputs(712));
    outputs(3155) <= not((layer2_outputs(2666)) or (layer2_outputs(495)));
    outputs(3156) <= layer2_outputs(1630);
    outputs(3157) <= not(layer2_outputs(4388));
    outputs(3158) <= not(layer2_outputs(4946)) or (layer2_outputs(2593));
    outputs(3159) <= not(layer2_outputs(2967));
    outputs(3160) <= not(layer2_outputs(3872)) or (layer2_outputs(3859));
    outputs(3161) <= not((layer2_outputs(4673)) or (layer2_outputs(2580)));
    outputs(3162) <= layer2_outputs(1342);
    outputs(3163) <= layer2_outputs(564);
    outputs(3164) <= not(layer2_outputs(1334));
    outputs(3165) <= (layer2_outputs(2823)) and (layer2_outputs(2317));
    outputs(3166) <= not(layer2_outputs(1512));
    outputs(3167) <= not(layer2_outputs(284));
    outputs(3168) <= (layer2_outputs(4912)) and not (layer2_outputs(3211));
    outputs(3169) <= (layer2_outputs(4177)) and (layer2_outputs(75));
    outputs(3170) <= not(layer2_outputs(3279));
    outputs(3171) <= not((layer2_outputs(503)) xor (layer2_outputs(1976)));
    outputs(3172) <= (layer2_outputs(2465)) and not (layer2_outputs(1036));
    outputs(3173) <= not(layer2_outputs(1716));
    outputs(3174) <= (layer2_outputs(321)) and (layer2_outputs(1041));
    outputs(3175) <= not((layer2_outputs(3238)) xor (layer2_outputs(2336)));
    outputs(3176) <= not(layer2_outputs(688));
    outputs(3177) <= not(layer2_outputs(337));
    outputs(3178) <= (layer2_outputs(3529)) or (layer2_outputs(3774));
    outputs(3179) <= (layer2_outputs(630)) xor (layer2_outputs(802));
    outputs(3180) <= not(layer2_outputs(2853));
    outputs(3181) <= layer2_outputs(2420);
    outputs(3182) <= (layer2_outputs(3562)) or (layer2_outputs(434));
    outputs(3183) <= layer2_outputs(3492);
    outputs(3184) <= not(layer2_outputs(4863));
    outputs(3185) <= not(layer2_outputs(4006));
    outputs(3186) <= not((layer2_outputs(1112)) xor (layer2_outputs(2455)));
    outputs(3187) <= layer2_outputs(3968);
    outputs(3188) <= not(layer2_outputs(4541));
    outputs(3189) <= not(layer2_outputs(4191));
    outputs(3190) <= not(layer2_outputs(2233));
    outputs(3191) <= layer2_outputs(3206);
    outputs(3192) <= layer2_outputs(1752);
    outputs(3193) <= not(layer2_outputs(1280));
    outputs(3194) <= layer2_outputs(1260);
    outputs(3195) <= not(layer2_outputs(3263));
    outputs(3196) <= (layer2_outputs(1771)) and not (layer2_outputs(3757));
    outputs(3197) <= not(layer2_outputs(36));
    outputs(3198) <= layer2_outputs(1768);
    outputs(3199) <= (layer2_outputs(938)) and (layer2_outputs(490));
    outputs(3200) <= not(layer2_outputs(3574));
    outputs(3201) <= not(layer2_outputs(1861));
    outputs(3202) <= not((layer2_outputs(4443)) xor (layer2_outputs(1118)));
    outputs(3203) <= not(layer2_outputs(1613));
    outputs(3204) <= not(layer2_outputs(4626)) or (layer2_outputs(591));
    outputs(3205) <= not(layer2_outputs(4013));
    outputs(3206) <= not((layer2_outputs(1245)) or (layer2_outputs(4656)));
    outputs(3207) <= (layer2_outputs(1464)) xor (layer2_outputs(1712));
    outputs(3208) <= (layer2_outputs(2776)) or (layer2_outputs(673));
    outputs(3209) <= not((layer2_outputs(2656)) or (layer2_outputs(3848)));
    outputs(3210) <= not(layer2_outputs(2159));
    outputs(3211) <= layer2_outputs(4494);
    outputs(3212) <= (layer2_outputs(3306)) and not (layer2_outputs(1207));
    outputs(3213) <= not(layer2_outputs(2178));
    outputs(3214) <= layer2_outputs(1564);
    outputs(3215) <= not(layer2_outputs(858));
    outputs(3216) <= layer2_outputs(1013);
    outputs(3217) <= layer2_outputs(3331);
    outputs(3218) <= not(layer2_outputs(4224));
    outputs(3219) <= not((layer2_outputs(4582)) or (layer2_outputs(3573)));
    outputs(3220) <= not(layer2_outputs(1377));
    outputs(3221) <= layer2_outputs(2349);
    outputs(3222) <= not(layer2_outputs(383));
    outputs(3223) <= not((layer2_outputs(1277)) xor (layer2_outputs(4360)));
    outputs(3224) <= layer2_outputs(4161);
    outputs(3225) <= not(layer2_outputs(1137));
    outputs(3226) <= layer2_outputs(3225);
    outputs(3227) <= not(layer2_outputs(4617));
    outputs(3228) <= (layer2_outputs(1408)) and not (layer2_outputs(1762));
    outputs(3229) <= not(layer2_outputs(2346));
    outputs(3230) <= layer2_outputs(1918);
    outputs(3231) <= not(layer2_outputs(2178));
    outputs(3232) <= not(layer2_outputs(2773));
    outputs(3233) <= not(layer2_outputs(47));
    outputs(3234) <= (layer2_outputs(3391)) xor (layer2_outputs(806));
    outputs(3235) <= not((layer2_outputs(1572)) or (layer2_outputs(4963)));
    outputs(3236) <= (layer2_outputs(934)) and (layer2_outputs(4060));
    outputs(3237) <= layer2_outputs(3345);
    outputs(3238) <= not((layer2_outputs(2498)) or (layer2_outputs(2952)));
    outputs(3239) <= layer2_outputs(2935);
    outputs(3240) <= (layer2_outputs(4505)) and not (layer2_outputs(668));
    outputs(3241) <= layer2_outputs(718);
    outputs(3242) <= (layer2_outputs(3523)) xor (layer2_outputs(3153));
    outputs(3243) <= not(layer2_outputs(3205));
    outputs(3244) <= not(layer2_outputs(1791)) or (layer2_outputs(1139));
    outputs(3245) <= not((layer2_outputs(3591)) xor (layer2_outputs(1950)));
    outputs(3246) <= (layer2_outputs(3463)) xor (layer2_outputs(828));
    outputs(3247) <= not(layer2_outputs(1287));
    outputs(3248) <= layer2_outputs(1505);
    outputs(3249) <= not(layer2_outputs(4085));
    outputs(3250) <= layer2_outputs(1100);
    outputs(3251) <= (layer2_outputs(809)) and not (layer2_outputs(3702));
    outputs(3252) <= not(layer2_outputs(3744));
    outputs(3253) <= not((layer2_outputs(3346)) and (layer2_outputs(3201)));
    outputs(3254) <= (layer2_outputs(5020)) xor (layer2_outputs(413));
    outputs(3255) <= not(layer2_outputs(619));
    outputs(3256) <= not(layer2_outputs(1778));
    outputs(3257) <= (layer2_outputs(4071)) and (layer2_outputs(259));
    outputs(3258) <= not(layer2_outputs(2930));
    outputs(3259) <= not(layer2_outputs(2222));
    outputs(3260) <= not(layer2_outputs(19));
    outputs(3261) <= not(layer2_outputs(1919));
    outputs(3262) <= (layer2_outputs(1012)) xor (layer2_outputs(756));
    outputs(3263) <= layer2_outputs(3844);
    outputs(3264) <= layer2_outputs(3864);
    outputs(3265) <= not((layer2_outputs(2554)) or (layer2_outputs(1201)));
    outputs(3266) <= layer2_outputs(1649);
    outputs(3267) <= (layer2_outputs(2165)) xor (layer2_outputs(1765));
    outputs(3268) <= (layer2_outputs(533)) and (layer2_outputs(2039));
    outputs(3269) <= layer2_outputs(3959);
    outputs(3270) <= not((layer2_outputs(3138)) xor (layer2_outputs(996)));
    outputs(3271) <= not((layer2_outputs(1938)) xor (layer2_outputs(4443)));
    outputs(3272) <= not(layer2_outputs(136));
    outputs(3273) <= not(layer2_outputs(4402));
    outputs(3274) <= layer2_outputs(4602);
    outputs(3275) <= not(layer2_outputs(4367));
    outputs(3276) <= not(layer2_outputs(164));
    outputs(3277) <= not(layer2_outputs(4955));
    outputs(3278) <= not(layer2_outputs(2882));
    outputs(3279) <= not(layer2_outputs(4828));
    outputs(3280) <= layer2_outputs(2796);
    outputs(3281) <= (layer2_outputs(3460)) and (layer2_outputs(4359));
    outputs(3282) <= (layer2_outputs(4760)) xor (layer2_outputs(2626));
    outputs(3283) <= (layer2_outputs(2720)) and not (layer2_outputs(1165));
    outputs(3284) <= (layer2_outputs(3104)) and not (layer2_outputs(4910));
    outputs(3285) <= not(layer2_outputs(535));
    outputs(3286) <= not((layer2_outputs(1591)) or (layer2_outputs(2877)));
    outputs(3287) <= not((layer2_outputs(2875)) or (layer2_outputs(4658)));
    outputs(3288) <= not(layer2_outputs(3200)) or (layer2_outputs(5059));
    outputs(3289) <= not((layer2_outputs(3819)) and (layer2_outputs(4705)));
    outputs(3290) <= not(layer2_outputs(3892));
    outputs(3291) <= not(layer2_outputs(4803));
    outputs(3292) <= layer2_outputs(2398);
    outputs(3293) <= not(layer2_outputs(4781)) or (layer2_outputs(2582));
    outputs(3294) <= not(layer2_outputs(5091));
    outputs(3295) <= layer2_outputs(3183);
    outputs(3296) <= not((layer2_outputs(2641)) and (layer2_outputs(2766)));
    outputs(3297) <= not((layer2_outputs(3854)) or (layer2_outputs(1871)));
    outputs(3298) <= not(layer2_outputs(3252));
    outputs(3299) <= not((layer2_outputs(1103)) and (layer2_outputs(3715)));
    outputs(3300) <= layer2_outputs(3798);
    outputs(3301) <= layer2_outputs(1856);
    outputs(3302) <= not(layer2_outputs(2151));
    outputs(3303) <= not((layer2_outputs(224)) xor (layer2_outputs(1005)));
    outputs(3304) <= not(layer2_outputs(487));
    outputs(3305) <= layer2_outputs(5025);
    outputs(3306) <= not((layer2_outputs(1892)) or (layer2_outputs(838)));
    outputs(3307) <= not(layer2_outputs(593));
    outputs(3308) <= not(layer2_outputs(3762));
    outputs(3309) <= (layer2_outputs(3890)) xor (layer2_outputs(3909));
    outputs(3310) <= not((layer2_outputs(402)) or (layer2_outputs(4514)));
    outputs(3311) <= layer2_outputs(2235);
    outputs(3312) <= (layer2_outputs(39)) and not (layer2_outputs(363));
    outputs(3313) <= not(layer2_outputs(4378));
    outputs(3314) <= not((layer2_outputs(1371)) or (layer2_outputs(2226)));
    outputs(3315) <= layer2_outputs(4681);
    outputs(3316) <= not(layer2_outputs(3002));
    outputs(3317) <= layer2_outputs(1763);
    outputs(3318) <= not(layer2_outputs(5032));
    outputs(3319) <= layer2_outputs(1912);
    outputs(3320) <= layer2_outputs(3717);
    outputs(3321) <= not(layer2_outputs(4513));
    outputs(3322) <= not(layer2_outputs(3084));
    outputs(3323) <= layer2_outputs(4775);
    outputs(3324) <= not(layer2_outputs(2892));
    outputs(3325) <= layer2_outputs(2964);
    outputs(3326) <= layer2_outputs(4041);
    outputs(3327) <= layer2_outputs(3698);
    outputs(3328) <= not(layer2_outputs(3763)) or (layer2_outputs(50));
    outputs(3329) <= not(layer2_outputs(3687));
    outputs(3330) <= not(layer2_outputs(607));
    outputs(3331) <= not(layer2_outputs(271));
    outputs(3332) <= not(layer2_outputs(1511)) or (layer2_outputs(3820));
    outputs(3333) <= not(layer2_outputs(2760));
    outputs(3334) <= not(layer2_outputs(4961));
    outputs(3335) <= not(layer2_outputs(402));
    outputs(3336) <= layer2_outputs(4573);
    outputs(3337) <= not(layer2_outputs(1285));
    outputs(3338) <= (layer2_outputs(822)) and not (layer2_outputs(2400));
    outputs(3339) <= layer2_outputs(4438);
    outputs(3340) <= layer2_outputs(1887);
    outputs(3341) <= not(layer2_outputs(3359));
    outputs(3342) <= not(layer2_outputs(3353));
    outputs(3343) <= layer2_outputs(1636);
    outputs(3344) <= not(layer2_outputs(2430)) or (layer2_outputs(1061));
    outputs(3345) <= layer2_outputs(2745);
    outputs(3346) <= layer2_outputs(1295);
    outputs(3347) <= layer2_outputs(3731);
    outputs(3348) <= (layer2_outputs(766)) and not (layer2_outputs(1545));
    outputs(3349) <= not((layer2_outputs(4493)) xor (layer2_outputs(504)));
    outputs(3350) <= not(layer2_outputs(1895));
    outputs(3351) <= not(layer2_outputs(2238));
    outputs(3352) <= layer2_outputs(3321);
    outputs(3353) <= not(layer2_outputs(2484));
    outputs(3354) <= layer2_outputs(2751);
    outputs(3355) <= (layer2_outputs(4669)) or (layer2_outputs(3292));
    outputs(3356) <= layer2_outputs(1048);
    outputs(3357) <= not(layer2_outputs(176));
    outputs(3358) <= layer2_outputs(4647);
    outputs(3359) <= layer2_outputs(4826);
    outputs(3360) <= layer2_outputs(3277);
    outputs(3361) <= not(layer2_outputs(3802));
    outputs(3362) <= not(layer2_outputs(3437));
    outputs(3363) <= not((layer2_outputs(1757)) xor (layer2_outputs(1960)));
    outputs(3364) <= layer2_outputs(1999);
    outputs(3365) <= (layer2_outputs(4095)) xor (layer2_outputs(4509));
    outputs(3366) <= not((layer2_outputs(3887)) or (layer2_outputs(4463)));
    outputs(3367) <= layer2_outputs(3899);
    outputs(3368) <= layer2_outputs(2682);
    outputs(3369) <= not(layer2_outputs(800));
    outputs(3370) <= not(layer2_outputs(698)) or (layer2_outputs(3804));
    outputs(3371) <= not(layer2_outputs(3197));
    outputs(3372) <= layer2_outputs(4344);
    outputs(3373) <= layer2_outputs(679);
    outputs(3374) <= not(layer2_outputs(1068));
    outputs(3375) <= layer2_outputs(809);
    outputs(3376) <= not(layer2_outputs(4952));
    outputs(3377) <= layer2_outputs(1366);
    outputs(3378) <= layer2_outputs(4052);
    outputs(3379) <= not(layer2_outputs(3378));
    outputs(3380) <= (layer2_outputs(2916)) or (layer2_outputs(1708));
    outputs(3381) <= not(layer2_outputs(4067));
    outputs(3382) <= not(layer2_outputs(462)) or (layer2_outputs(4039));
    outputs(3383) <= layer2_outputs(4569);
    outputs(3384) <= layer2_outputs(471);
    outputs(3385) <= (layer2_outputs(4040)) and (layer2_outputs(241));
    outputs(3386) <= not(layer2_outputs(3627));
    outputs(3387) <= (layer2_outputs(3803)) xor (layer2_outputs(2219));
    outputs(3388) <= (layer2_outputs(589)) and not (layer2_outputs(3330));
    outputs(3389) <= (layer2_outputs(4200)) xor (layer2_outputs(2742));
    outputs(3390) <= layer2_outputs(2141);
    outputs(3391) <= (layer2_outputs(2544)) and not (layer2_outputs(3596));
    outputs(3392) <= layer2_outputs(4540);
    outputs(3393) <= (layer2_outputs(496)) and not (layer2_outputs(4537));
    outputs(3394) <= not(layer2_outputs(3088));
    outputs(3395) <= layer2_outputs(959);
    outputs(3396) <= not(layer2_outputs(4408));
    outputs(3397) <= not((layer2_outputs(4569)) xor (layer2_outputs(2184)));
    outputs(3398) <= (layer2_outputs(3239)) and (layer2_outputs(4461));
    outputs(3399) <= layer2_outputs(3066);
    outputs(3400) <= not(layer2_outputs(3630));
    outputs(3401) <= not((layer2_outputs(928)) xor (layer2_outputs(2414)));
    outputs(3402) <= (layer2_outputs(2285)) and not (layer2_outputs(3378));
    outputs(3403) <= layer2_outputs(3614);
    outputs(3404) <= layer2_outputs(2000);
    outputs(3405) <= not(layer2_outputs(2100));
    outputs(3406) <= not((layer2_outputs(557)) xor (layer2_outputs(474)));
    outputs(3407) <= layer2_outputs(1521);
    outputs(3408) <= not(layer2_outputs(1846));
    outputs(3409) <= layer2_outputs(1308);
    outputs(3410) <= layer2_outputs(1023);
    outputs(3411) <= layer2_outputs(4181);
    outputs(3412) <= layer2_outputs(4921);
    outputs(3413) <= not(layer2_outputs(1944));
    outputs(3414) <= not((layer2_outputs(4988)) xor (layer2_outputs(3866)));
    outputs(3415) <= not(layer2_outputs(2652));
    outputs(3416) <= layer2_outputs(614);
    outputs(3417) <= not(layer2_outputs(217));
    outputs(3418) <= (layer2_outputs(1517)) or (layer2_outputs(2931));
    outputs(3419) <= layer2_outputs(1478);
    outputs(3420) <= not(layer2_outputs(2656));
    outputs(3421) <= not(layer2_outputs(420));
    outputs(3422) <= layer2_outputs(3764);
    outputs(3423) <= layer2_outputs(540);
    outputs(3424) <= layer2_outputs(517);
    outputs(3425) <= layer2_outputs(2537);
    outputs(3426) <= layer2_outputs(2463);
    outputs(3427) <= not(layer2_outputs(5086));
    outputs(3428) <= not(layer2_outputs(4309)) or (layer2_outputs(3602));
    outputs(3429) <= layer2_outputs(1023);
    outputs(3430) <= (layer2_outputs(3383)) xor (layer2_outputs(226));
    outputs(3431) <= layer2_outputs(3614);
    outputs(3432) <= (layer2_outputs(2858)) xor (layer2_outputs(1972));
    outputs(3433) <= not(layer2_outputs(142));
    outputs(3434) <= (layer2_outputs(4545)) and (layer2_outputs(1348));
    outputs(3435) <= layer2_outputs(1525);
    outputs(3436) <= (layer2_outputs(1748)) or (layer2_outputs(1295));
    outputs(3437) <= layer2_outputs(3708);
    outputs(3438) <= not(layer2_outputs(2921));
    outputs(3439) <= not(layer2_outputs(3625));
    outputs(3440) <= not(layer2_outputs(4696));
    outputs(3441) <= layer2_outputs(1692);
    outputs(3442) <= not(layer2_outputs(2240)) or (layer2_outputs(3241));
    outputs(3443) <= layer2_outputs(3225);
    outputs(3444) <= layer2_outputs(4950);
    outputs(3445) <= not(layer2_outputs(2276));
    outputs(3446) <= not((layer2_outputs(963)) and (layer2_outputs(3705)));
    outputs(3447) <= layer2_outputs(1763);
    outputs(3448) <= (layer2_outputs(1319)) and not (layer2_outputs(3587));
    outputs(3449) <= layer2_outputs(4984);
    outputs(3450) <= layer2_outputs(1893);
    outputs(3451) <= (layer2_outputs(1243)) and (layer2_outputs(1948));
    outputs(3452) <= (layer2_outputs(2317)) and not (layer2_outputs(1450));
    outputs(3453) <= layer2_outputs(1092);
    outputs(3454) <= layer2_outputs(3089);
    outputs(3455) <= layer2_outputs(2931);
    outputs(3456) <= not(layer2_outputs(3091));
    outputs(3457) <= (layer2_outputs(1672)) and (layer2_outputs(3927));
    outputs(3458) <= not(layer2_outputs(3564)) or (layer2_outputs(1614));
    outputs(3459) <= not(layer2_outputs(166));
    outputs(3460) <= not(layer2_outputs(4335));
    outputs(3461) <= not(layer2_outputs(2369));
    outputs(3462) <= not(layer2_outputs(4045)) or (layer2_outputs(2384));
    outputs(3463) <= (layer2_outputs(4426)) xor (layer2_outputs(1713));
    outputs(3464) <= (layer2_outputs(451)) and (layer2_outputs(1542));
    outputs(3465) <= layer2_outputs(268);
    outputs(3466) <= layer2_outputs(614);
    outputs(3467) <= layer2_outputs(1069);
    outputs(3468) <= layer2_outputs(2035);
    outputs(3469) <= layer2_outputs(4210);
    outputs(3470) <= not(layer2_outputs(1890)) or (layer2_outputs(2769));
    outputs(3471) <= not((layer2_outputs(4673)) or (layer2_outputs(134)));
    outputs(3472) <= (layer2_outputs(1690)) xor (layer2_outputs(4940));
    outputs(3473) <= not(layer2_outputs(4567));
    outputs(3474) <= layer2_outputs(4117);
    outputs(3475) <= layer2_outputs(1402);
    outputs(3476) <= layer2_outputs(709);
    outputs(3477) <= not((layer2_outputs(4209)) and (layer2_outputs(4764)));
    outputs(3478) <= not((layer2_outputs(3756)) xor (layer2_outputs(4283)));
    outputs(3479) <= layer2_outputs(93);
    outputs(3480) <= (layer2_outputs(3004)) and not (layer2_outputs(3686));
    outputs(3481) <= not((layer2_outputs(4023)) xor (layer2_outputs(36)));
    outputs(3482) <= layer2_outputs(2138);
    outputs(3483) <= not(layer2_outputs(61));
    outputs(3484) <= not(layer2_outputs(2938));
    outputs(3485) <= (layer2_outputs(1330)) and not (layer2_outputs(5078));
    outputs(3486) <= not(layer2_outputs(1802));
    outputs(3487) <= (layer2_outputs(89)) and (layer2_outputs(3425));
    outputs(3488) <= not(layer2_outputs(1755));
    outputs(3489) <= not(layer2_outputs(3599));
    outputs(3490) <= not(layer2_outputs(1263));
    outputs(3491) <= not((layer2_outputs(4906)) and (layer2_outputs(1735)));
    outputs(3492) <= not((layer2_outputs(148)) or (layer2_outputs(4513)));
    outputs(3493) <= not(layer2_outputs(3918)) or (layer2_outputs(3963));
    outputs(3494) <= layer2_outputs(3998);
    outputs(3495) <= (layer2_outputs(3143)) xor (layer2_outputs(1198));
    outputs(3496) <= layer2_outputs(426);
    outputs(3497) <= not((layer2_outputs(1787)) xor (layer2_outputs(1288)));
    outputs(3498) <= not((layer2_outputs(3285)) xor (layer2_outputs(3543)));
    outputs(3499) <= (layer2_outputs(4629)) and (layer2_outputs(2824));
    outputs(3500) <= not(layer2_outputs(923));
    outputs(3501) <= (layer2_outputs(230)) and not (layer2_outputs(1378));
    outputs(3502) <= not(layer2_outputs(4980));
    outputs(3503) <= layer2_outputs(2748);
    outputs(3504) <= (layer2_outputs(3748)) and not (layer2_outputs(4903));
    outputs(3505) <= not(layer2_outputs(218));
    outputs(3506) <= not((layer2_outputs(4063)) or (layer2_outputs(2107)));
    outputs(3507) <= not(layer2_outputs(1510));
    outputs(3508) <= layer2_outputs(281);
    outputs(3509) <= not(layer2_outputs(4870));
    outputs(3510) <= (layer2_outputs(1817)) xor (layer2_outputs(3928));
    outputs(3511) <= layer2_outputs(4164);
    outputs(3512) <= layer2_outputs(4256);
    outputs(3513) <= (layer2_outputs(4762)) xor (layer2_outputs(3784));
    outputs(3514) <= not((layer2_outputs(3629)) xor (layer2_outputs(1227)));
    outputs(3515) <= not(layer2_outputs(3516));
    outputs(3516) <= layer2_outputs(1256);
    outputs(3517) <= (layer2_outputs(2291)) or (layer2_outputs(709));
    outputs(3518) <= not(layer2_outputs(1072));
    outputs(3519) <= not((layer2_outputs(495)) xor (layer2_outputs(1316)));
    outputs(3520) <= not((layer2_outputs(969)) xor (layer2_outputs(4772)));
    outputs(3521) <= layer2_outputs(4672);
    outputs(3522) <= not((layer2_outputs(1785)) or (layer2_outputs(1998)));
    outputs(3523) <= not(layer2_outputs(1538));
    outputs(3524) <= not(layer2_outputs(4591));
    outputs(3525) <= (layer2_outputs(3853)) and (layer2_outputs(1437));
    outputs(3526) <= not(layer2_outputs(4227));
    outputs(3527) <= not((layer2_outputs(2540)) xor (layer2_outputs(1379)));
    outputs(3528) <= not(layer2_outputs(665));
    outputs(3529) <= layer2_outputs(618);
    outputs(3530) <= layer2_outputs(3577);
    outputs(3531) <= layer2_outputs(4786);
    outputs(3532) <= layer2_outputs(4544);
    outputs(3533) <= not(layer2_outputs(358));
    outputs(3534) <= layer2_outputs(1176);
    outputs(3535) <= layer2_outputs(3360);
    outputs(3536) <= not(layer2_outputs(3905));
    outputs(3537) <= layer2_outputs(2792);
    outputs(3538) <= not(layer2_outputs(452));
    outputs(3539) <= layer2_outputs(122);
    outputs(3540) <= (layer2_outputs(736)) and not (layer2_outputs(2209));
    outputs(3541) <= not(layer2_outputs(165));
    outputs(3542) <= not(layer2_outputs(4422));
    outputs(3543) <= not(layer2_outputs(4079));
    outputs(3544) <= layer2_outputs(5025);
    outputs(3545) <= layer2_outputs(4417);
    outputs(3546) <= not(layer2_outputs(1445));
    outputs(3547) <= not(layer2_outputs(3359));
    outputs(3548) <= layer2_outputs(4756);
    outputs(3549) <= (layer2_outputs(1425)) or (layer2_outputs(3610));
    outputs(3550) <= not(layer2_outputs(198));
    outputs(3551) <= not(layer2_outputs(1008));
    outputs(3552) <= (layer2_outputs(2098)) xor (layer2_outputs(2476));
    outputs(3553) <= not(layer2_outputs(552));
    outputs(3554) <= (layer2_outputs(3775)) xor (layer2_outputs(4419));
    outputs(3555) <= (layer2_outputs(3350)) xor (layer2_outputs(4537));
    outputs(3556) <= layer2_outputs(86);
    outputs(3557) <= (layer2_outputs(1252)) or (layer2_outputs(2927));
    outputs(3558) <= layer2_outputs(1055);
    outputs(3559) <= not((layer2_outputs(3949)) xor (layer2_outputs(3476)));
    outputs(3560) <= not(layer2_outputs(41));
    outputs(3561) <= not((layer2_outputs(5029)) or (layer2_outputs(1448)));
    outputs(3562) <= not((layer2_outputs(922)) or (layer2_outputs(3732)));
    outputs(3563) <= (layer2_outputs(4444)) and not (layer2_outputs(3714));
    outputs(3564) <= not(layer2_outputs(2207));
    outputs(3565) <= (layer2_outputs(2526)) and not (layer2_outputs(2377));
    outputs(3566) <= not(layer2_outputs(1588));
    outputs(3567) <= layer2_outputs(1491);
    outputs(3568) <= not(layer2_outputs(1011));
    outputs(3569) <= layer2_outputs(2129);
    outputs(3570) <= not((layer2_outputs(2995)) xor (layer2_outputs(4423)));
    outputs(3571) <= not(layer2_outputs(3989)) or (layer2_outputs(4821));
    outputs(3572) <= not(layer2_outputs(384));
    outputs(3573) <= not(layer2_outputs(526));
    outputs(3574) <= not(layer2_outputs(3817));
    outputs(3575) <= not(layer2_outputs(2562)) or (layer2_outputs(2632));
    outputs(3576) <= not(layer2_outputs(4282));
    outputs(3577) <= not(layer2_outputs(3706));
    outputs(3578) <= not(layer2_outputs(132));
    outputs(3579) <= not(layer2_outputs(1761));
    outputs(3580) <= layer2_outputs(2021);
    outputs(3581) <= not(layer2_outputs(17));
    outputs(3582) <= (layer2_outputs(3507)) xor (layer2_outputs(4592));
    outputs(3583) <= layer2_outputs(2618);
    outputs(3584) <= layer2_outputs(446);
    outputs(3585) <= not(layer2_outputs(3158));
    outputs(3586) <= layer2_outputs(4332);
    outputs(3587) <= layer2_outputs(204);
    outputs(3588) <= layer2_outputs(3323);
    outputs(3589) <= not((layer2_outputs(3339)) xor (layer2_outputs(2085)));
    outputs(3590) <= layer2_outputs(143);
    outputs(3591) <= layer2_outputs(2394);
    outputs(3592) <= (layer2_outputs(4192)) and not (layer2_outputs(151));
    outputs(3593) <= (layer2_outputs(521)) and not (layer2_outputs(937));
    outputs(3594) <= not(layer2_outputs(4674));
    outputs(3595) <= not(layer2_outputs(2434));
    outputs(3596) <= layer2_outputs(1238);
    outputs(3597) <= not(layer2_outputs(1960));
    outputs(3598) <= (layer2_outputs(1147)) xor (layer2_outputs(4593));
    outputs(3599) <= layer2_outputs(3624);
    outputs(3600) <= (layer2_outputs(4004)) and (layer2_outputs(1641));
    outputs(3601) <= (layer2_outputs(2175)) and not (layer2_outputs(1454));
    outputs(3602) <= layer2_outputs(4873);
    outputs(3603) <= not(layer2_outputs(2199));
    outputs(3604) <= not(layer2_outputs(4260));
    outputs(3605) <= (layer2_outputs(2828)) and (layer2_outputs(2651));
    outputs(3606) <= layer2_outputs(1551);
    outputs(3607) <= not(layer2_outputs(90));
    outputs(3608) <= layer2_outputs(3667);
    outputs(3609) <= not(layer2_outputs(1587));
    outputs(3610) <= not(layer2_outputs(1077));
    outputs(3611) <= layer2_outputs(3490);
    outputs(3612) <= layer2_outputs(4960);
    outputs(3613) <= not((layer2_outputs(1698)) or (layer2_outputs(278)));
    outputs(3614) <= not((layer2_outputs(3568)) xor (layer2_outputs(3282)));
    outputs(3615) <= not(layer2_outputs(3134));
    outputs(3616) <= layer2_outputs(2809);
    outputs(3617) <= (layer2_outputs(2023)) xor (layer2_outputs(1541));
    outputs(3618) <= not((layer2_outputs(267)) or (layer2_outputs(1194)));
    outputs(3619) <= not(layer2_outputs(1441));
    outputs(3620) <= not(layer2_outputs(4240));
    outputs(3621) <= not(layer2_outputs(527));
    outputs(3622) <= layer2_outputs(3464);
    outputs(3623) <= not((layer2_outputs(2408)) xor (layer2_outputs(2114)));
    outputs(3624) <= not(layer2_outputs(1440));
    outputs(3625) <= not(layer2_outputs(333));
    outputs(3626) <= layer2_outputs(3761);
    outputs(3627) <= (layer2_outputs(4866)) xor (layer2_outputs(1425));
    outputs(3628) <= (layer2_outputs(660)) and not (layer2_outputs(3795));
    outputs(3629) <= layer2_outputs(2153);
    outputs(3630) <= layer2_outputs(3525);
    outputs(3631) <= (layer2_outputs(2322)) and not (layer2_outputs(1728));
    outputs(3632) <= not(layer2_outputs(260));
    outputs(3633) <= not(layer2_outputs(1903));
    outputs(3634) <= layer2_outputs(815);
    outputs(3635) <= layer2_outputs(3441);
    outputs(3636) <= not(layer2_outputs(1434));
    outputs(3637) <= not(layer2_outputs(2716));
    outputs(3638) <= not((layer2_outputs(4675)) xor (layer2_outputs(5047)));
    outputs(3639) <= layer2_outputs(1221);
    outputs(3640) <= not(layer2_outputs(4347));
    outputs(3641) <= (layer2_outputs(2384)) and not (layer2_outputs(4718));
    outputs(3642) <= layer2_outputs(2332);
    outputs(3643) <= (layer2_outputs(1404)) and not (layer2_outputs(4279));
    outputs(3644) <= layer2_outputs(1024);
    outputs(3645) <= (layer2_outputs(322)) and (layer2_outputs(443));
    outputs(3646) <= not(layer2_outputs(3693));
    outputs(3647) <= (layer2_outputs(802)) and (layer2_outputs(2949));
    outputs(3648) <= (layer2_outputs(3671)) and (layer2_outputs(837));
    outputs(3649) <= not(layer2_outputs(1842));
    outputs(3650) <= not((layer2_outputs(1672)) xor (layer2_outputs(4336)));
    outputs(3651) <= layer2_outputs(3290);
    outputs(3652) <= (layer2_outputs(4710)) and (layer2_outputs(2803));
    outputs(3653) <= layer2_outputs(3772);
    outputs(3654) <= not(layer2_outputs(2003));
    outputs(3655) <= layer2_outputs(2529);
    outputs(3656) <= layer2_outputs(329);
    outputs(3657) <= layer2_outputs(3925);
    outputs(3658) <= layer2_outputs(3186);
    outputs(3659) <= (layer2_outputs(2667)) and not (layer2_outputs(780));
    outputs(3660) <= (layer2_outputs(2115)) and (layer2_outputs(2301));
    outputs(3661) <= not(layer2_outputs(2693));
    outputs(3662) <= not(layer2_outputs(476));
    outputs(3663) <= not(layer2_outputs(2745));
    outputs(3664) <= layer2_outputs(488);
    outputs(3665) <= layer2_outputs(2344);
    outputs(3666) <= layer2_outputs(3955);
    outputs(3667) <= not((layer2_outputs(4916)) or (layer2_outputs(3856)));
    outputs(3668) <= (layer2_outputs(3430)) and (layer2_outputs(4732));
    outputs(3669) <= layer2_outputs(3094);
    outputs(3670) <= not((layer2_outputs(3679)) xor (layer2_outputs(945)));
    outputs(3671) <= not(layer2_outputs(1147));
    outputs(3672) <= (layer2_outputs(99)) and not (layer2_outputs(4854));
    outputs(3673) <= (layer2_outputs(3788)) and not (layer2_outputs(3907));
    outputs(3674) <= not((layer2_outputs(187)) xor (layer2_outputs(204)));
    outputs(3675) <= layer2_outputs(877);
    outputs(3676) <= (layer2_outputs(3601)) and (layer2_outputs(1533));
    outputs(3677) <= not(layer2_outputs(4489));
    outputs(3678) <= (layer2_outputs(3700)) and not (layer2_outputs(2798));
    outputs(3679) <= not(layer2_outputs(2321));
    outputs(3680) <= not((layer2_outputs(4239)) or (layer2_outputs(4584)));
    outputs(3681) <= (layer2_outputs(3648)) and not (layer2_outputs(2603));
    outputs(3682) <= not(layer2_outputs(1728));
    outputs(3683) <= not((layer2_outputs(2029)) or (layer2_outputs(3210)));
    outputs(3684) <= layer2_outputs(2374);
    outputs(3685) <= layer2_outputs(1731);
    outputs(3686) <= layer2_outputs(2362);
    outputs(3687) <= layer2_outputs(5054);
    outputs(3688) <= layer2_outputs(1876);
    outputs(3689) <= not(layer2_outputs(3904));
    outputs(3690) <= not((layer2_outputs(2726)) or (layer2_outputs(4699)));
    outputs(3691) <= not(layer2_outputs(998));
    outputs(3692) <= not(layer2_outputs(3950));
    outputs(3693) <= not(layer2_outputs(1461));
    outputs(3694) <= not(layer2_outputs(177));
    outputs(3695) <= not((layer2_outputs(2600)) or (layer2_outputs(2138)));
    outputs(3696) <= not(layer2_outputs(586));
    outputs(3697) <= not(layer2_outputs(2316));
    outputs(3698) <= (layer2_outputs(2960)) and not (layer2_outputs(1152));
    outputs(3699) <= (layer2_outputs(82)) or (layer2_outputs(2220));
    outputs(3700) <= layer2_outputs(3483);
    outputs(3701) <= layer2_outputs(3391);
    outputs(3702) <= not((layer2_outputs(889)) xor (layer2_outputs(1190)));
    outputs(3703) <= not(layer2_outputs(2594));
    outputs(3704) <= not(layer2_outputs(4282));
    outputs(3705) <= (layer2_outputs(2210)) and not (layer2_outputs(3956));
    outputs(3706) <= (layer2_outputs(2989)) and not (layer2_outputs(647));
    outputs(3707) <= not(layer2_outputs(3218));
    outputs(3708) <= (layer2_outputs(752)) and (layer2_outputs(25));
    outputs(3709) <= not(layer2_outputs(2014));
    outputs(3710) <= not(layer2_outputs(554));
    outputs(3711) <= (layer2_outputs(601)) and (layer2_outputs(4160));
    outputs(3712) <= not(layer2_outputs(935));
    outputs(3713) <= layer2_outputs(4169);
    outputs(3714) <= (layer2_outputs(2359)) xor (layer2_outputs(4989));
    outputs(3715) <= (layer2_outputs(3961)) and (layer2_outputs(3209));
    outputs(3716) <= (layer2_outputs(2223)) xor (layer2_outputs(2201));
    outputs(3717) <= (layer2_outputs(2872)) and (layer2_outputs(3865));
    outputs(3718) <= not(layer2_outputs(3981)) or (layer2_outputs(776));
    outputs(3719) <= (layer2_outputs(3486)) and (layer2_outputs(2207));
    outputs(3720) <= not((layer2_outputs(266)) or (layer2_outputs(774)));
    outputs(3721) <= not((layer2_outputs(4270)) or (layer2_outputs(1362)));
    outputs(3722) <= layer2_outputs(2197);
    outputs(3723) <= not((layer2_outputs(3621)) or (layer2_outputs(4410)));
    outputs(3724) <= not(layer2_outputs(1894));
    outputs(3725) <= not((layer2_outputs(108)) and (layer2_outputs(2489)));
    outputs(3726) <= (layer2_outputs(3986)) xor (layer2_outputs(590));
    outputs(3727) <= not((layer2_outputs(950)) xor (layer2_outputs(2859)));
    outputs(3728) <= not(layer2_outputs(2251));
    outputs(3729) <= (layer2_outputs(4155)) and (layer2_outputs(134));
    outputs(3730) <= (layer2_outputs(1156)) and not (layer2_outputs(234));
    outputs(3731) <= not(layer2_outputs(245)) or (layer2_outputs(4081));
    outputs(3732) <= not(layer2_outputs(4245));
    outputs(3733) <= layer2_outputs(2250);
    outputs(3734) <= (layer2_outputs(4068)) or (layer2_outputs(4465));
    outputs(3735) <= (layer2_outputs(4082)) xor (layer2_outputs(3116));
    outputs(3736) <= not((layer2_outputs(877)) xor (layer2_outputs(744)));
    outputs(3737) <= layer2_outputs(1663);
    outputs(3738) <= not(layer2_outputs(2596));
    outputs(3739) <= not(layer2_outputs(525));
    outputs(3740) <= not(layer2_outputs(2478));
    outputs(3741) <= not((layer2_outputs(1164)) or (layer2_outputs(5099)));
    outputs(3742) <= layer2_outputs(2441);
    outputs(3743) <= layer2_outputs(4093);
    outputs(3744) <= not(layer2_outputs(3235));
    outputs(3745) <= layer2_outputs(2809);
    outputs(3746) <= layer2_outputs(2862);
    outputs(3747) <= layer2_outputs(2301);
    outputs(3748) <= not((layer2_outputs(266)) or (layer2_outputs(2333)));
    outputs(3749) <= (layer2_outputs(1262)) xor (layer2_outputs(1867));
    outputs(3750) <= layer2_outputs(615);
    outputs(3751) <= layer2_outputs(435);
    outputs(3752) <= not(layer2_outputs(0)) or (layer2_outputs(3709));
    outputs(3753) <= not(layer2_outputs(2874));
    outputs(3754) <= not(layer2_outputs(5080)) or (layer2_outputs(911));
    outputs(3755) <= layer2_outputs(128);
    outputs(3756) <= (layer2_outputs(1460)) and (layer2_outputs(2923));
    outputs(3757) <= (layer2_outputs(4785)) and (layer2_outputs(671));
    outputs(3758) <= not((layer2_outputs(305)) xor (layer2_outputs(2255)));
    outputs(3759) <= not(layer2_outputs(1372));
    outputs(3760) <= not(layer2_outputs(2131));
    outputs(3761) <= not((layer2_outputs(4805)) or (layer2_outputs(5108)));
    outputs(3762) <= layer2_outputs(4788);
    outputs(3763) <= not(layer2_outputs(833));
    outputs(3764) <= layer2_outputs(80);
    outputs(3765) <= layer2_outputs(4575);
    outputs(3766) <= layer2_outputs(3490);
    outputs(3767) <= not((layer2_outputs(2986)) xor (layer2_outputs(369)));
    outputs(3768) <= layer2_outputs(692);
    outputs(3769) <= layer2_outputs(1632);
    outputs(3770) <= layer2_outputs(4036);
    outputs(3771) <= not(layer2_outputs(4987));
    outputs(3772) <= not(layer2_outputs(3967));
    outputs(3773) <= (layer2_outputs(1289)) and (layer2_outputs(1153));
    outputs(3774) <= (layer2_outputs(4126)) or (layer2_outputs(2639));
    outputs(3775) <= layer2_outputs(1535);
    outputs(3776) <= (layer2_outputs(4342)) and not (layer2_outputs(3400));
    outputs(3777) <= not(layer2_outputs(2885));
    outputs(3778) <= not(layer2_outputs(334));
    outputs(3779) <= layer2_outputs(3059);
    outputs(3780) <= not(layer2_outputs(243)) or (layer2_outputs(359));
    outputs(3781) <= layer2_outputs(119);
    outputs(3782) <= layer2_outputs(3190);
    outputs(3783) <= (layer2_outputs(4871)) xor (layer2_outputs(4414));
    outputs(3784) <= layer2_outputs(4044);
    outputs(3785) <= layer2_outputs(1666);
    outputs(3786) <= not(layer2_outputs(4944));
    outputs(3787) <= (layer2_outputs(1628)) and (layer2_outputs(872));
    outputs(3788) <= (layer2_outputs(4547)) xor (layer2_outputs(2266));
    outputs(3789) <= layer2_outputs(2763);
    outputs(3790) <= not(layer2_outputs(783));
    outputs(3791) <= layer2_outputs(4454);
    outputs(3792) <= layer2_outputs(340);
    outputs(3793) <= (layer2_outputs(3673)) xor (layer2_outputs(1240));
    outputs(3794) <= not((layer2_outputs(1034)) xor (layer2_outputs(527)));
    outputs(3795) <= (layer2_outputs(1566)) and not (layer2_outputs(2152));
    outputs(3796) <= (layer2_outputs(233)) and not (layer2_outputs(3305));
    outputs(3797) <= (layer2_outputs(4679)) and not (layer2_outputs(2354));
    outputs(3798) <= (layer2_outputs(1391)) xor (layer2_outputs(597));
    outputs(3799) <= layer2_outputs(1606);
    outputs(3800) <= (layer2_outputs(3521)) xor (layer2_outputs(3697));
    outputs(3801) <= (layer2_outputs(965)) and not (layer2_outputs(930));
    outputs(3802) <= (layer2_outputs(3099)) and not (layer2_outputs(3767));
    outputs(3803) <= not((layer2_outputs(1376)) xor (layer2_outputs(606)));
    outputs(3804) <= (layer2_outputs(4521)) xor (layer2_outputs(3544));
    outputs(3805) <= layer2_outputs(3832);
    outputs(3806) <= layer2_outputs(1361);
    outputs(3807) <= (layer2_outputs(2845)) and (layer2_outputs(3010));
    outputs(3808) <= (layer2_outputs(2475)) xor (layer2_outputs(1777));
    outputs(3809) <= not(layer2_outputs(5005));
    outputs(3810) <= not((layer2_outputs(4172)) or (layer2_outputs(705)));
    outputs(3811) <= layer2_outputs(687);
    outputs(3812) <= not(layer2_outputs(396)) or (layer2_outputs(742));
    outputs(3813) <= not(layer2_outputs(2984));
    outputs(3814) <= (layer2_outputs(785)) and not (layer2_outputs(4125));
    outputs(3815) <= layer2_outputs(1012);
    outputs(3816) <= (layer2_outputs(3033)) and (layer2_outputs(2036));
    outputs(3817) <= not(layer2_outputs(4495));
    outputs(3818) <= (layer2_outputs(4615)) and not (layer2_outputs(2302));
    outputs(3819) <= not(layer2_outputs(4076));
    outputs(3820) <= layer2_outputs(3788);
    outputs(3821) <= not(layer2_outputs(10));
    outputs(3822) <= layer2_outputs(4759);
    outputs(3823) <= not(layer2_outputs(1009));
    outputs(3824) <= (layer2_outputs(4910)) and (layer2_outputs(1685));
    outputs(3825) <= (layer2_outputs(4807)) and not (layer2_outputs(4468));
    outputs(3826) <= not(layer2_outputs(1616));
    outputs(3827) <= (layer2_outputs(3273)) and (layer2_outputs(3962));
    outputs(3828) <= layer2_outputs(3099);
    outputs(3829) <= not(layer2_outputs(3681));
    outputs(3830) <= (layer2_outputs(2565)) xor (layer2_outputs(1126));
    outputs(3831) <= not(layer2_outputs(3475));
    outputs(3832) <= not((layer2_outputs(4184)) and (layer2_outputs(4010)));
    outputs(3833) <= not((layer2_outputs(3990)) or (layer2_outputs(2894)));
    outputs(3834) <= not((layer2_outputs(4915)) or (layer2_outputs(193)));
    outputs(3835) <= (layer2_outputs(5054)) and not (layer2_outputs(3692));
    outputs(3836) <= (layer2_outputs(2275)) and not (layer2_outputs(3758));
    outputs(3837) <= not(layer2_outputs(978));
    outputs(3838) <= not((layer2_outputs(4163)) xor (layer2_outputs(1608)));
    outputs(3839) <= not(layer2_outputs(1112));
    outputs(3840) <= not(layer2_outputs(4791));
    outputs(3841) <= layer2_outputs(2274);
    outputs(3842) <= layer2_outputs(1369);
    outputs(3843) <= not(layer2_outputs(1180));
    outputs(3844) <= not(layer2_outputs(3424)) or (layer2_outputs(4612));
    outputs(3845) <= layer2_outputs(301);
    outputs(3846) <= layer2_outputs(2904);
    outputs(3847) <= (layer2_outputs(2251)) xor (layer2_outputs(3938));
    outputs(3848) <= layer2_outputs(1906);
    outputs(3849) <= not((layer2_outputs(2694)) xor (layer2_outputs(4085)));
    outputs(3850) <= not((layer2_outputs(355)) xor (layer2_outputs(4893)));
    outputs(3851) <= (layer2_outputs(2492)) and (layer2_outputs(4883));
    outputs(3852) <= not(layer2_outputs(3855));
    outputs(3853) <= layer2_outputs(1037);
    outputs(3854) <= not(layer2_outputs(1567));
    outputs(3855) <= not(layer2_outputs(2903));
    outputs(3856) <= not(layer2_outputs(2490));
    outputs(3857) <= (layer2_outputs(3927)) and not (layer2_outputs(2277));
    outputs(3858) <= layer2_outputs(4009);
    outputs(3859) <= layer2_outputs(2111);
    outputs(3860) <= layer2_outputs(444);
    outputs(3861) <= layer2_outputs(514);
    outputs(3862) <= layer2_outputs(218);
    outputs(3863) <= layer2_outputs(4011);
    outputs(3864) <= not(layer2_outputs(4306));
    outputs(3865) <= layer2_outputs(2299);
    outputs(3866) <= layer2_outputs(5089);
    outputs(3867) <= layer2_outputs(2168);
    outputs(3868) <= (layer2_outputs(2431)) and not (layer2_outputs(2254));
    outputs(3869) <= layer2_outputs(2322);
    outputs(3870) <= (layer2_outputs(3541)) and not (layer2_outputs(2330));
    outputs(3871) <= (layer2_outputs(2908)) and (layer2_outputs(3569));
    outputs(3872) <= layer2_outputs(3428);
    outputs(3873) <= not(layer2_outputs(4263));
    outputs(3874) <= layer2_outputs(1458);
    outputs(3875) <= layer2_outputs(4812);
    outputs(3876) <= not((layer2_outputs(1260)) or (layer2_outputs(2770)));
    outputs(3877) <= not(layer2_outputs(117));
    outputs(3878) <= layer2_outputs(2049);
    outputs(3879) <= (layer2_outputs(592)) and not (layer2_outputs(3414));
    outputs(3880) <= not(layer2_outputs(1190));
    outputs(3881) <= not((layer2_outputs(2462)) or (layer2_outputs(3997)));
    outputs(3882) <= not(layer2_outputs(2888));
    outputs(3883) <= not(layer2_outputs(1973));
    outputs(3884) <= (layer2_outputs(2424)) and not (layer2_outputs(4772));
    outputs(3885) <= not(layer2_outputs(2888));
    outputs(3886) <= layer2_outputs(1809);
    outputs(3887) <= not(layer2_outputs(4054));
    outputs(3888) <= (layer2_outputs(3624)) and not (layer2_outputs(2443));
    outputs(3889) <= not((layer2_outputs(4105)) xor (layer2_outputs(4058)));
    outputs(3890) <= not(layer2_outputs(3093));
    outputs(3891) <= not(layer2_outputs(1346));
    outputs(3892) <= not(layer2_outputs(89));
    outputs(3893) <= (layer2_outputs(3897)) or (layer2_outputs(4765));
    outputs(3894) <= '0';
    outputs(3895) <= not((layer2_outputs(2813)) xor (layer2_outputs(3417)));
    outputs(3896) <= not(layer2_outputs(2378)) or (layer2_outputs(3141));
    outputs(3897) <= layer2_outputs(2653);
    outputs(3898) <= (layer2_outputs(378)) and (layer2_outputs(3613));
    outputs(3899) <= not((layer2_outputs(2104)) xor (layer2_outputs(4654)));
    outputs(3900) <= not(layer2_outputs(4930)) or (layer2_outputs(973));
    outputs(3901) <= (layer2_outputs(2308)) and (layer2_outputs(2389));
    outputs(3902) <= not(layer2_outputs(931));
    outputs(3903) <= layer2_outputs(4358);
    outputs(3904) <= not((layer2_outputs(2561)) or (layer2_outputs(2136)));
    outputs(3905) <= not(layer2_outputs(3181));
    outputs(3906) <= layer2_outputs(105);
    outputs(3907) <= layer2_outputs(1701);
    outputs(3908) <= layer2_outputs(1902);
    outputs(3909) <= (layer2_outputs(1438)) xor (layer2_outputs(4887));
    outputs(3910) <= not(layer2_outputs(4360));
    outputs(3911) <= layer2_outputs(3230);
    outputs(3912) <= layer2_outputs(4333);
    outputs(3913) <= layer2_outputs(3827);
    outputs(3914) <= not(layer2_outputs(4997));
    outputs(3915) <= not(layer2_outputs(4703));
    outputs(3916) <= layer2_outputs(4340);
    outputs(3917) <= (layer2_outputs(4596)) and not (layer2_outputs(3877));
    outputs(3918) <= not(layer2_outputs(880));
    outputs(3919) <= layer2_outputs(477);
    outputs(3920) <= not(layer2_outputs(2649));
    outputs(3921) <= (layer2_outputs(1135)) and (layer2_outputs(4690));
    outputs(3922) <= not((layer2_outputs(44)) xor (layer2_outputs(3071)));
    outputs(3923) <= not(layer2_outputs(5036));
    outputs(3924) <= not(layer2_outputs(1462));
    outputs(3925) <= layer2_outputs(605);
    outputs(3926) <= (layer2_outputs(2375)) and not (layer2_outputs(4162));
    outputs(3927) <= not(layer2_outputs(2372));
    outputs(3928) <= (layer2_outputs(3987)) and not (layer2_outputs(2634));
    outputs(3929) <= (layer2_outputs(3581)) and not (layer2_outputs(3978));
    outputs(3930) <= not((layer2_outputs(4556)) xor (layer2_outputs(805)));
    outputs(3931) <= (layer2_outputs(4092)) and not (layer2_outputs(4613));
    outputs(3932) <= layer2_outputs(472);
    outputs(3933) <= (layer2_outputs(1591)) and not (layer2_outputs(562));
    outputs(3934) <= layer2_outputs(668);
    outputs(3935) <= (layer2_outputs(1895)) and (layer2_outputs(2853));
    outputs(3936) <= not(layer2_outputs(2377));
    outputs(3937) <= not((layer2_outputs(2496)) or (layer2_outputs(2293)));
    outputs(3938) <= not(layer2_outputs(765));
    outputs(3939) <= not(layer2_outputs(2881));
    outputs(3940) <= not(layer2_outputs(1250));
    outputs(3941) <= not((layer2_outputs(2658)) and (layer2_outputs(5076)));
    outputs(3942) <= not(layer2_outputs(2455));
    outputs(3943) <= layer2_outputs(171);
    outputs(3944) <= not(layer2_outputs(3781));
    outputs(3945) <= layer2_outputs(3483);
    outputs(3946) <= (layer2_outputs(71)) and not (layer2_outputs(2192));
    outputs(3947) <= layer2_outputs(4662);
    outputs(3948) <= layer2_outputs(2545);
    outputs(3949) <= layer2_outputs(48);
    outputs(3950) <= layer2_outputs(290);
    outputs(3951) <= (layer2_outputs(3658)) and (layer2_outputs(2715));
    outputs(3952) <= not(layer2_outputs(4924));
    outputs(3953) <= (layer2_outputs(1785)) and not (layer2_outputs(360));
    outputs(3954) <= layer2_outputs(4372);
    outputs(3955) <= (layer2_outputs(4603)) and not (layer2_outputs(505));
    outputs(3956) <= layer2_outputs(1489);
    outputs(3957) <= (layer2_outputs(851)) and (layer2_outputs(4462));
    outputs(3958) <= (layer2_outputs(2606)) and not (layer2_outputs(3919));
    outputs(3959) <= not(layer2_outputs(812));
    outputs(3960) <= layer2_outputs(1978);
    outputs(3961) <= layer2_outputs(2581);
    outputs(3962) <= not((layer2_outputs(3602)) or (layer2_outputs(4676)));
    outputs(3963) <= (layer2_outputs(3091)) and not (layer2_outputs(773));
    outputs(3964) <= (layer2_outputs(486)) and not (layer2_outputs(3121));
    outputs(3965) <= not(layer2_outputs(433));
    outputs(3966) <= (layer2_outputs(1143)) and not (layer2_outputs(3510));
    outputs(3967) <= not(layer2_outputs(3463));
    outputs(3968) <= (layer2_outputs(4083)) xor (layer2_outputs(1032));
    outputs(3969) <= not(layer2_outputs(3592));
    outputs(3970) <= layer2_outputs(4753);
    outputs(3971) <= layer2_outputs(3786);
    outputs(3972) <= layer2_outputs(3870);
    outputs(3973) <= not(layer2_outputs(2233));
    outputs(3974) <= (layer2_outputs(91)) and (layer2_outputs(1793));
    outputs(3975) <= (layer2_outputs(1037)) and (layer2_outputs(1493));
    outputs(3976) <= not(layer2_outputs(4413));
    outputs(3977) <= (layer2_outputs(3894)) or (layer2_outputs(2427));
    outputs(3978) <= not((layer2_outputs(3524)) or (layer2_outputs(5017)));
    outputs(3979) <= (layer2_outputs(3155)) and not (layer2_outputs(780));
    outputs(3980) <= not(layer2_outputs(3192));
    outputs(3981) <= layer2_outputs(2610);
    outputs(3982) <= layer2_outputs(2616);
    outputs(3983) <= not(layer2_outputs(411));
    outputs(3984) <= not((layer2_outputs(3061)) or (layer2_outputs(1586)));
    outputs(3985) <= layer2_outputs(3383);
    outputs(3986) <= not(layer2_outputs(1626));
    outputs(3987) <= not(layer2_outputs(2354)) or (layer2_outputs(2674));
    outputs(3988) <= not(layer2_outputs(2316));
    outputs(3989) <= not((layer2_outputs(26)) xor (layer2_outputs(3220)));
    outputs(3990) <= (layer2_outputs(1937)) and not (layer2_outputs(1670));
    outputs(3991) <= (layer2_outputs(2755)) xor (layer2_outputs(3202));
    outputs(3992) <= layer2_outputs(4832);
    outputs(3993) <= not(layer2_outputs(203));
    outputs(3994) <= (layer2_outputs(5050)) and not (layer2_outputs(1714));
    outputs(3995) <= not((layer2_outputs(5024)) xor (layer2_outputs(2255)));
    outputs(3996) <= (layer2_outputs(3434)) xor (layer2_outputs(4151));
    outputs(3997) <= not(layer2_outputs(3026));
    outputs(3998) <= not(layer2_outputs(5114));
    outputs(3999) <= layer2_outputs(1161);
    outputs(4000) <= (layer2_outputs(4954)) and not (layer2_outputs(5062));
    outputs(4001) <= (layer2_outputs(2074)) and (layer2_outputs(3880));
    outputs(4002) <= not((layer2_outputs(174)) xor (layer2_outputs(212)));
    outputs(4003) <= not(layer2_outputs(728));
    outputs(4004) <= layer2_outputs(3135);
    outputs(4005) <= (layer2_outputs(2494)) and not (layer2_outputs(974));
    outputs(4006) <= (layer2_outputs(4578)) or (layer2_outputs(3227));
    outputs(4007) <= not(layer2_outputs(4251));
    outputs(4008) <= layer2_outputs(4037);
    outputs(4009) <= layer2_outputs(2948);
    outputs(4010) <= layer2_outputs(2270);
    outputs(4011) <= (layer2_outputs(1563)) and (layer2_outputs(4019));
    outputs(4012) <= layer2_outputs(2981);
    outputs(4013) <= (layer2_outputs(4371)) and not (layer2_outputs(2045));
    outputs(4014) <= not(layer2_outputs(676));
    outputs(4015) <= not(layer2_outputs(3399));
    outputs(4016) <= not((layer2_outputs(4331)) xor (layer2_outputs(3132)));
    outputs(4017) <= not(layer2_outputs(2329));
    outputs(4018) <= (layer2_outputs(3685)) xor (layer2_outputs(1676));
    outputs(4019) <= not(layer2_outputs(3869));
    outputs(4020) <= not(layer2_outputs(3345));
    outputs(4021) <= (layer2_outputs(78)) or (layer2_outputs(1781));
    outputs(4022) <= not(layer2_outputs(202));
    outputs(4023) <= layer2_outputs(2491);
    outputs(4024) <= (layer2_outputs(3980)) and (layer2_outputs(4870));
    outputs(4025) <= not((layer2_outputs(2241)) or (layer2_outputs(158)));
    outputs(4026) <= layer2_outputs(408);
    outputs(4027) <= (layer2_outputs(3281)) xor (layer2_outputs(3711));
    outputs(4028) <= (layer2_outputs(4503)) and not (layer2_outputs(173));
    outputs(4029) <= layer2_outputs(1987);
    outputs(4030) <= not(layer2_outputs(2280)) or (layer2_outputs(3209));
    outputs(4031) <= not(layer2_outputs(760));
    outputs(4032) <= not((layer2_outputs(4491)) and (layer2_outputs(23)));
    outputs(4033) <= layer2_outputs(4618);
    outputs(4034) <= layer2_outputs(680);
    outputs(4035) <= not(layer2_outputs(1061));
    outputs(4036) <= layer2_outputs(4671);
    outputs(4037) <= layer2_outputs(3901);
    outputs(4038) <= not(layer2_outputs(992)) or (layer2_outputs(2975));
    outputs(4039) <= (layer2_outputs(3361)) and not (layer2_outputs(4353));
    outputs(4040) <= '0';
    outputs(4041) <= not(layer2_outputs(1845));
    outputs(4042) <= (layer2_outputs(4446)) and not (layer2_outputs(1860));
    outputs(4043) <= not(layer2_outputs(4259));
    outputs(4044) <= (layer2_outputs(499)) and not (layer2_outputs(2194));
    outputs(4045) <= (layer2_outputs(4785)) and not (layer2_outputs(3812));
    outputs(4046) <= (layer2_outputs(4411)) and (layer2_outputs(3700));
    outputs(4047) <= layer2_outputs(4358);
    outputs(4048) <= not(layer2_outputs(2390));
    outputs(4049) <= (layer2_outputs(4867)) and not (layer2_outputs(2723));
    outputs(4050) <= layer2_outputs(1912);
    outputs(4051) <= layer2_outputs(3574);
    outputs(4052) <= (layer2_outputs(3423)) and not (layer2_outputs(1524));
    outputs(4053) <= not(layer2_outputs(2457));
    outputs(4054) <= not(layer2_outputs(379)) or (layer2_outputs(1715));
    outputs(4055) <= layer2_outputs(4436);
    outputs(4056) <= not((layer2_outputs(4202)) xor (layer2_outputs(3968)));
    outputs(4057) <= (layer2_outputs(861)) and not (layer2_outputs(4123));
    outputs(4058) <= layer2_outputs(3117);
    outputs(4059) <= (layer2_outputs(265)) and not (layer2_outputs(4937));
    outputs(4060) <= not((layer2_outputs(541)) xor (layer2_outputs(223)));
    outputs(4061) <= (layer2_outputs(382)) xor (layer2_outputs(1721));
    outputs(4062) <= not(layer2_outputs(653)) or (layer2_outputs(5112));
    outputs(4063) <= (layer2_outputs(4392)) xor (layer2_outputs(3127));
    outputs(4064) <= not(layer2_outputs(4437));
    outputs(4065) <= (layer2_outputs(285)) and not (layer2_outputs(577));
    outputs(4066) <= not(layer2_outputs(3552)) or (layer2_outputs(3052));
    outputs(4067) <= layer2_outputs(611);
    outputs(4068) <= not(layer2_outputs(2038));
    outputs(4069) <= not(layer2_outputs(3693));
    outputs(4070) <= (layer2_outputs(2609)) and not (layer2_outputs(459));
    outputs(4071) <= (layer2_outputs(1808)) xor (layer2_outputs(3865));
    outputs(4072) <= layer2_outputs(1731);
    outputs(4073) <= not((layer2_outputs(132)) xor (layer2_outputs(3871)));
    outputs(4074) <= layer2_outputs(3782);
    outputs(4075) <= (layer2_outputs(1649)) and not (layer2_outputs(540));
    outputs(4076) <= not(layer2_outputs(836)) or (layer2_outputs(441));
    outputs(4077) <= not(layer2_outputs(2082));
    outputs(4078) <= layer2_outputs(2307);
    outputs(4079) <= layer2_outputs(507);
    outputs(4080) <= (layer2_outputs(4583)) and not (layer2_outputs(827));
    outputs(4081) <= (layer2_outputs(4813)) and (layer2_outputs(2221));
    outputs(4082) <= (layer2_outputs(3874)) and not (layer2_outputs(1948));
    outputs(4083) <= not(layer2_outputs(3454));
    outputs(4084) <= layer2_outputs(3110);
    outputs(4085) <= (layer2_outputs(1644)) and not (layer2_outputs(1129));
    outputs(4086) <= not((layer2_outputs(278)) or (layer2_outputs(924)));
    outputs(4087) <= not(layer2_outputs(4284));
    outputs(4088) <= not(layer2_outputs(4681));
    outputs(4089) <= (layer2_outputs(449)) and (layer2_outputs(2449));
    outputs(4090) <= not((layer2_outputs(4726)) or (layer2_outputs(14)));
    outputs(4091) <= not(layer2_outputs(4613));
    outputs(4092) <= layer2_outputs(4881);
    outputs(4093) <= not(layer2_outputs(2353));
    outputs(4094) <= not((layer2_outputs(2556)) xor (layer2_outputs(3179)));
    outputs(4095) <= not(layer2_outputs(4677));
    outputs(4096) <= not(layer2_outputs(4873));
    outputs(4097) <= (layer2_outputs(3453)) xor (layer2_outputs(26));
    outputs(4098) <= layer2_outputs(46);
    outputs(4099) <= not(layer2_outputs(1276));
    outputs(4100) <= layer2_outputs(2168);
    outputs(4101) <= not((layer2_outputs(2502)) xor (layer2_outputs(3722)));
    outputs(4102) <= not(layer2_outputs(4968));
    outputs(4103) <= layer2_outputs(3366);
    outputs(4104) <= not(layer2_outputs(1374));
    outputs(4105) <= not(layer2_outputs(582));
    outputs(4106) <= layer2_outputs(2538);
    outputs(4107) <= layer2_outputs(4262);
    outputs(4108) <= (layer2_outputs(1017)) and (layer2_outputs(13));
    outputs(4109) <= not(layer2_outputs(3308)) or (layer2_outputs(138));
    outputs(4110) <= (layer2_outputs(695)) xor (layer2_outputs(3121));
    outputs(4111) <= not(layer2_outputs(1144));
    outputs(4112) <= not(layer2_outputs(3045));
    outputs(4113) <= not(layer2_outputs(3688));
    outputs(4114) <= (layer2_outputs(4590)) or (layer2_outputs(3196));
    outputs(4115) <= not(layer2_outputs(1198));
    outputs(4116) <= not(layer2_outputs(2812)) or (layer2_outputs(657));
    outputs(4117) <= (layer2_outputs(3174)) xor (layer2_outputs(3312));
    outputs(4118) <= not(layer2_outputs(1903));
    outputs(4119) <= not(layer2_outputs(4204));
    outputs(4120) <= layer2_outputs(702);
    outputs(4121) <= not(layer2_outputs(4684));
    outputs(4122) <= (layer2_outputs(3620)) and not (layer2_outputs(2681));
    outputs(4123) <= not(layer2_outputs(1000));
    outputs(4124) <= layer2_outputs(962);
    outputs(4125) <= not((layer2_outputs(4985)) xor (layer2_outputs(248)));
    outputs(4126) <= not(layer2_outputs(2563));
    outputs(4127) <= layer2_outputs(277);
    outputs(4128) <= not(layer2_outputs(3455));
    outputs(4129) <= (layer2_outputs(794)) and not (layer2_outputs(761));
    outputs(4130) <= not(layer2_outputs(1309));
    outputs(4131) <= not(layer2_outputs(2943)) or (layer2_outputs(4456));
    outputs(4132) <= not(layer2_outputs(1290));
    outputs(4133) <= (layer2_outputs(634)) and not (layer2_outputs(2958));
    outputs(4134) <= layer2_outputs(3513);
    outputs(4135) <= not(layer2_outputs(2248));
    outputs(4136) <= layer2_outputs(4368);
    outputs(4137) <= (layer2_outputs(2385)) xor (layer2_outputs(3868));
    outputs(4138) <= layer2_outputs(4977);
    outputs(4139) <= layer2_outputs(2821);
    outputs(4140) <= not((layer2_outputs(367)) or (layer2_outputs(2214)));
    outputs(4141) <= not((layer2_outputs(2306)) xor (layer2_outputs(4928)));
    outputs(4142) <= (layer2_outputs(3936)) and not (layer2_outputs(3103));
    outputs(4143) <= layer2_outputs(4668);
    outputs(4144) <= layer2_outputs(738);
    outputs(4145) <= not((layer2_outputs(2524)) and (layer2_outputs(2542)));
    outputs(4146) <= not(layer2_outputs(1986));
    outputs(4147) <= not((layer2_outputs(1217)) xor (layer2_outputs(4311)));
    outputs(4148) <= not(layer2_outputs(1653));
    outputs(4149) <= (layer2_outputs(34)) and (layer2_outputs(312));
    outputs(4150) <= not(layer2_outputs(1529));
    outputs(4151) <= (layer2_outputs(2398)) xor (layer2_outputs(4744));
    outputs(4152) <= not((layer2_outputs(686)) xor (layer2_outputs(2458)));
    outputs(4153) <= not(layer2_outputs(1455));
    outputs(4154) <= not(layer2_outputs(1222)) or (layer2_outputs(818));
    outputs(4155) <= not((layer2_outputs(1990)) xor (layer2_outputs(2482)));
    outputs(4156) <= layer2_outputs(4014);
    outputs(4157) <= not(layer2_outputs(4157));
    outputs(4158) <= layer2_outputs(556);
    outputs(4159) <= not((layer2_outputs(720)) and (layer2_outputs(3008)));
    outputs(4160) <= not(layer2_outputs(2536)) or (layer2_outputs(5044));
    outputs(4161) <= not(layer2_outputs(3431));
    outputs(4162) <= not(layer2_outputs(317));
    outputs(4163) <= layer2_outputs(5021);
    outputs(4164) <= layer2_outputs(672);
    outputs(4165) <= not(layer2_outputs(2852));
    outputs(4166) <= layer2_outputs(2863);
    outputs(4167) <= layer2_outputs(2198);
    outputs(4168) <= layer2_outputs(2918);
    outputs(4169) <= layer2_outputs(4389);
    outputs(4170) <= not(layer2_outputs(3666));
    outputs(4171) <= layer2_outputs(2424);
    outputs(4172) <= not(layer2_outputs(1577));
    outputs(4173) <= layer2_outputs(4624);
    outputs(4174) <= not((layer2_outputs(2256)) and (layer2_outputs(376)));
    outputs(4175) <= not((layer2_outputs(3092)) xor (layer2_outputs(3821)));
    outputs(4176) <= not(layer2_outputs(3073)) or (layer2_outputs(4616));
    outputs(4177) <= not(layer2_outputs(3522));
    outputs(4178) <= (layer2_outputs(4976)) xor (layer2_outputs(1645));
    outputs(4179) <= layer2_outputs(5021);
    outputs(4180) <= not((layer2_outputs(2062)) and (layer2_outputs(4145)));
    outputs(4181) <= not(layer2_outputs(1932));
    outputs(4182) <= not(layer2_outputs(1110));
    outputs(4183) <= not(layer2_outputs(2691));
    outputs(4184) <= (layer2_outputs(2591)) or (layer2_outputs(3311));
    outputs(4185) <= not(layer2_outputs(4622));
    outputs(4186) <= layer2_outputs(2177);
    outputs(4187) <= not(layer2_outputs(1266));
    outputs(4188) <= layer2_outputs(1282);
    outputs(4189) <= layer2_outputs(5036);
    outputs(4190) <= not((layer2_outputs(1824)) and (layer2_outputs(2386)));
    outputs(4191) <= layer2_outputs(3375);
    outputs(4192) <= not(layer2_outputs(916));
    outputs(4193) <= (layer2_outputs(1973)) and not (layer2_outputs(3500));
    outputs(4194) <= (layer2_outputs(3791)) or (layer2_outputs(4465));
    outputs(4195) <= layer2_outputs(4628);
    outputs(4196) <= not((layer2_outputs(3573)) xor (layer2_outputs(3575)));
    outputs(4197) <= not(layer2_outputs(4278));
    outputs(4198) <= layer2_outputs(1693);
    outputs(4199) <= layer2_outputs(1648);
    outputs(4200) <= not(layer2_outputs(3608));
    outputs(4201) <= not(layer2_outputs(455)) or (layer2_outputs(2952));
    outputs(4202) <= (layer2_outputs(713)) and (layer2_outputs(388));
    outputs(4203) <= layer2_outputs(2031);
    outputs(4204) <= not(layer2_outputs(2861));
    outputs(4205) <= layer2_outputs(635);
    outputs(4206) <= not(layer2_outputs(197));
    outputs(4207) <= (layer2_outputs(3244)) xor (layer2_outputs(3591));
    outputs(4208) <= not(layer2_outputs(5087));
    outputs(4209) <= (layer2_outputs(3741)) xor (layer2_outputs(3013));
    outputs(4210) <= (layer2_outputs(5031)) xor (layer2_outputs(4109));
    outputs(4211) <= not(layer2_outputs(2133));
    outputs(4212) <= layer2_outputs(2475);
    outputs(4213) <= (layer2_outputs(3930)) xor (layer2_outputs(288));
    outputs(4214) <= not(layer2_outputs(2205));
    outputs(4215) <= not(layer2_outputs(520));
    outputs(4216) <= (layer2_outputs(1453)) and not (layer2_outputs(3526));
    outputs(4217) <= not(layer2_outputs(2486));
    outputs(4218) <= layer2_outputs(2796);
    outputs(4219) <= not(layer2_outputs(1297)) or (layer2_outputs(2673));
    outputs(4220) <= not((layer2_outputs(1955)) or (layer2_outputs(850)));
    outputs(4221) <= (layer2_outputs(863)) xor (layer2_outputs(1409));
    outputs(4222) <= (layer2_outputs(1300)) xor (layer2_outputs(2422));
    outputs(4223) <= not(layer2_outputs(122)) or (layer2_outputs(1335));
    outputs(4224) <= not(layer2_outputs(4505));
    outputs(4225) <= not(layer2_outputs(4385));
    outputs(4226) <= not(layer2_outputs(3388));
    outputs(4227) <= not(layer2_outputs(2944));
    outputs(4228) <= (layer2_outputs(979)) xor (layer2_outputs(2896));
    outputs(4229) <= not(layer2_outputs(3230));
    outputs(4230) <= (layer2_outputs(798)) and not (layer2_outputs(914));
    outputs(4231) <= not(layer2_outputs(1496));
    outputs(4232) <= not(layer2_outputs(2096));
    outputs(4233) <= layer2_outputs(4744);
    outputs(4234) <= not((layer2_outputs(1056)) xor (layer2_outputs(1218)));
    outputs(4235) <= not(layer2_outputs(2517)) or (layer2_outputs(336));
    outputs(4236) <= (layer2_outputs(4249)) xor (layer2_outputs(2379));
    outputs(4237) <= not(layer2_outputs(1908));
    outputs(4238) <= not((layer2_outputs(4351)) or (layer2_outputs(4270)));
    outputs(4239) <= (layer2_outputs(1525)) xor (layer2_outputs(3603));
    outputs(4240) <= not(layer2_outputs(1905));
    outputs(4241) <= layer2_outputs(1880);
    outputs(4242) <= layer2_outputs(1050);
    outputs(4243) <= not(layer2_outputs(1318));
    outputs(4244) <= layer2_outputs(1605);
    outputs(4245) <= not(layer2_outputs(1355));
    outputs(4246) <= not(layer2_outputs(3247)) or (layer2_outputs(4437));
    outputs(4247) <= not(layer2_outputs(2943));
    outputs(4248) <= layer2_outputs(4835);
    outputs(4249) <= layer2_outputs(1272);
    outputs(4250) <= not(layer2_outputs(2851));
    outputs(4251) <= (layer2_outputs(4109)) and not (layer2_outputs(2799));
    outputs(4252) <= not(layer2_outputs(1331));
    outputs(4253) <= (layer2_outputs(3214)) and (layer2_outputs(539));
    outputs(4254) <= not(layer2_outputs(3879));
    outputs(4255) <= not((layer2_outputs(2008)) or (layer2_outputs(1210)));
    outputs(4256) <= not((layer2_outputs(1610)) or (layer2_outputs(2308)));
    outputs(4257) <= layer2_outputs(4390);
    outputs(4258) <= not(layer2_outputs(4078));
    outputs(4259) <= not((layer2_outputs(1029)) xor (layer2_outputs(2817)));
    outputs(4260) <= layer2_outputs(1380);
    outputs(4261) <= not(layer2_outputs(3608));
    outputs(4262) <= not(layer2_outputs(2607));
    outputs(4263) <= layer2_outputs(3983);
    outputs(4264) <= not(layer2_outputs(1779));
    outputs(4265) <= not(layer2_outputs(241)) or (layer2_outputs(4156));
    outputs(4266) <= (layer2_outputs(1411)) or (layer2_outputs(2366));
    outputs(4267) <= not((layer2_outputs(4201)) xor (layer2_outputs(4600)));
    outputs(4268) <= (layer2_outputs(1063)) and (layer2_outputs(1402));
    outputs(4269) <= '1';
    outputs(4270) <= (layer2_outputs(645)) xor (layer2_outputs(154));
    outputs(4271) <= (layer2_outputs(4315)) or (layer2_outputs(799));
    outputs(4272) <= (layer2_outputs(2728)) and not (layer2_outputs(4928));
    outputs(4273) <= not(layer2_outputs(1177)) or (layer2_outputs(3900));
    outputs(4274) <= (layer2_outputs(1602)) and not (layer2_outputs(601));
    outputs(4275) <= (layer2_outputs(4829)) and not (layer2_outputs(2439));
    outputs(4276) <= not(layer2_outputs(2464)) or (layer2_outputs(4667));
    outputs(4277) <= (layer2_outputs(722)) and not (layer2_outputs(2905));
    outputs(4278) <= not(layer2_outputs(3082)) or (layer2_outputs(3672));
    outputs(4279) <= not(layer2_outputs(957));
    outputs(4280) <= not(layer2_outputs(720));
    outputs(4281) <= not(layer2_outputs(2282)) or (layer2_outputs(1436));
    outputs(4282) <= not(layer2_outputs(4454));
    outputs(4283) <= not((layer2_outputs(2558)) xor (layer2_outputs(623)));
    outputs(4284) <= not(layer2_outputs(2951));
    outputs(4285) <= layer2_outputs(513);
    outputs(4286) <= (layer2_outputs(2126)) and (layer2_outputs(644));
    outputs(4287) <= not(layer2_outputs(2069));
    outputs(4288) <= not((layer2_outputs(510)) xor (layer2_outputs(288)));
    outputs(4289) <= layer2_outputs(1421);
    outputs(4290) <= (layer2_outputs(1982)) xor (layer2_outputs(1187));
    outputs(4291) <= not(layer2_outputs(4068)) or (layer2_outputs(4843));
    outputs(4292) <= layer2_outputs(2785);
    outputs(4293) <= not(layer2_outputs(1271));
    outputs(4294) <= not(layer2_outputs(912));
    outputs(4295) <= (layer2_outputs(3710)) and not (layer2_outputs(4187));
    outputs(4296) <= not((layer2_outputs(4657)) and (layer2_outputs(3772)));
    outputs(4297) <= layer2_outputs(1);
    outputs(4298) <= not(layer2_outputs(3173));
    outputs(4299) <= layer2_outputs(1054);
    outputs(4300) <= layer2_outputs(1952);
    outputs(4301) <= layer2_outputs(3320);
    outputs(4302) <= layer2_outputs(4366);
    outputs(4303) <= not(layer2_outputs(916));
    outputs(4304) <= not(layer2_outputs(463)) or (layer2_outputs(2960));
    outputs(4305) <= not(layer2_outputs(39));
    outputs(4306) <= layer2_outputs(4837);
    outputs(4307) <= not(layer2_outputs(2271));
    outputs(4308) <= not(layer2_outputs(1145)) or (layer2_outputs(3367));
    outputs(4309) <= layer2_outputs(5057);
    outputs(4310) <= layer2_outputs(4605);
    outputs(4311) <= layer2_outputs(353);
    outputs(4312) <= (layer2_outputs(4648)) and (layer2_outputs(3340));
    outputs(4313) <= layer2_outputs(2198);
    outputs(4314) <= (layer2_outputs(1939)) and not (layer2_outputs(4276));
    outputs(4315) <= not(layer2_outputs(3431));
    outputs(4316) <= layer2_outputs(3167);
    outputs(4317) <= not(layer2_outputs(2545));
    outputs(4318) <= not(layer2_outputs(3800));
    outputs(4319) <= not(layer2_outputs(4732)) or (layer2_outputs(4790));
    outputs(4320) <= layer2_outputs(4789);
    outputs(4321) <= (layer2_outputs(4557)) and (layer2_outputs(982));
    outputs(4322) <= layer2_outputs(1810);
    outputs(4323) <= not(layer2_outputs(2227));
    outputs(4324) <= not(layer2_outputs(3248));
    outputs(4325) <= (layer2_outputs(4309)) xor (layer2_outputs(4478));
    outputs(4326) <= not(layer2_outputs(3028));
    outputs(4327) <= layer2_outputs(2212);
    outputs(4328) <= not(layer2_outputs(5030));
    outputs(4329) <= not(layer2_outputs(298));
    outputs(4330) <= not(layer2_outputs(4381)) or (layer2_outputs(4388));
    outputs(4331) <= not(layer2_outputs(3271));
    outputs(4332) <= layer2_outputs(1737);
    outputs(4333) <= layer2_outputs(3755);
    outputs(4334) <= layer2_outputs(519);
    outputs(4335) <= not(layer2_outputs(1703));
    outputs(4336) <= not(layer2_outputs(3125)) or (layer2_outputs(2093));
    outputs(4337) <= (layer2_outputs(3672)) or (layer2_outputs(1710));
    outputs(4338) <= not(layer2_outputs(2537));
    outputs(4339) <= layer2_outputs(958);
    outputs(4340) <= not(layer2_outputs(948));
    outputs(4341) <= (layer2_outputs(2884)) and (layer2_outputs(629));
    outputs(4342) <= not((layer2_outputs(4220)) or (layer2_outputs(2592)));
    outputs(4343) <= layer2_outputs(974);
    outputs(4344) <= (layer2_outputs(4894)) and not (layer2_outputs(3771));
    outputs(4345) <= not(layer2_outputs(3622));
    outputs(4346) <= not(layer2_outputs(4098));
    outputs(4347) <= not((layer2_outputs(320)) and (layer2_outputs(4657)));
    outputs(4348) <= not(layer2_outputs(5083));
    outputs(4349) <= not(layer2_outputs(5083));
    outputs(4350) <= layer2_outputs(3678);
    outputs(4351) <= layer2_outputs(2950);
    outputs(4352) <= not(layer2_outputs(2867));
    outputs(4353) <= not(layer2_outputs(1046));
    outputs(4354) <= not(layer2_outputs(2221));
    outputs(4355) <= not((layer2_outputs(1459)) and (layer2_outputs(3226)));
    outputs(4356) <= not(layer2_outputs(2300)) or (layer2_outputs(771));
    outputs(4357) <= not(layer2_outputs(4545)) or (layer2_outputs(2997));
    outputs(4358) <= (layer2_outputs(430)) and not (layer2_outputs(4216));
    outputs(4359) <= (layer2_outputs(2447)) xor (layer2_outputs(3212));
    outputs(4360) <= layer2_outputs(1781);
    outputs(4361) <= (layer2_outputs(5077)) xor (layer2_outputs(4440));
    outputs(4362) <= not((layer2_outputs(2895)) xor (layer2_outputs(4874)));
    outputs(4363) <= not((layer2_outputs(5018)) xor (layer2_outputs(1015)));
    outputs(4364) <= not(layer2_outputs(3331)) or (layer2_outputs(1286));
    outputs(4365) <= layer2_outputs(2355);
    outputs(4366) <= (layer2_outputs(2086)) or (layer2_outputs(2052));
    outputs(4367) <= layer2_outputs(675);
    outputs(4368) <= (layer2_outputs(4091)) xor (layer2_outputs(2412));
    outputs(4369) <= (layer2_outputs(1317)) and not (layer2_outputs(2119));
    outputs(4370) <= not(layer2_outputs(2325));
    outputs(4371) <= not(layer2_outputs(3908));
    outputs(4372) <= not(layer2_outputs(547)) or (layer2_outputs(3841));
    outputs(4373) <= layer2_outputs(1891);
    outputs(4374) <= layer2_outputs(3462);
    outputs(4375) <= not((layer2_outputs(4571)) or (layer2_outputs(2689)));
    outputs(4376) <= layer2_outputs(889);
    outputs(4377) <= layer2_outputs(1162);
    outputs(4378) <= layer2_outputs(1502);
    outputs(4379) <= not((layer2_outputs(3334)) xor (layer2_outputs(3808)));
    outputs(4380) <= layer2_outputs(2392);
    outputs(4381) <= not(layer2_outputs(3182));
    outputs(4382) <= (layer2_outputs(439)) or (layer2_outputs(3160));
    outputs(4383) <= layer2_outputs(4617);
    outputs(4384) <= layer2_outputs(1281);
    outputs(4385) <= layer2_outputs(3240);
    outputs(4386) <= not(layer2_outputs(538));
    outputs(4387) <= not(layer2_outputs(4412)) or (layer2_outputs(3632));
    outputs(4388) <= not(layer2_outputs(4107)) or (layer2_outputs(4770));
    outputs(4389) <= not(layer2_outputs(2597));
    outputs(4390) <= not(layer2_outputs(256));
    outputs(4391) <= layer2_outputs(4985);
    outputs(4392) <= not(layer2_outputs(1633));
    outputs(4393) <= (layer2_outputs(2462)) xor (layer2_outputs(4848));
    outputs(4394) <= not(layer2_outputs(4344)) or (layer2_outputs(1384));
    outputs(4395) <= layer2_outputs(3933);
    outputs(4396) <= layer2_outputs(4148);
    outputs(4397) <= layer2_outputs(4826);
    outputs(4398) <= layer2_outputs(2445);
    outputs(4399) <= not(layer2_outputs(3238));
    outputs(4400) <= layer2_outputs(397);
    outputs(4401) <= not(layer2_outputs(447));
    outputs(4402) <= not(layer2_outputs(3943));
    outputs(4403) <= layer2_outputs(2400);
    outputs(4404) <= not(layer2_outputs(1695));
    outputs(4405) <= not(layer2_outputs(450));
    outputs(4406) <= layer2_outputs(3802);
    outputs(4407) <= not((layer2_outputs(3197)) or (layer2_outputs(1569)));
    outputs(4408) <= not(layer2_outputs(4323));
    outputs(4409) <= (layer2_outputs(947)) and not (layer2_outputs(1879));
    outputs(4410) <= not(layer2_outputs(1945));
    outputs(4411) <= layer2_outputs(1913);
    outputs(4412) <= layer2_outputs(3039);
    outputs(4413) <= not(layer2_outputs(1459));
    outputs(4414) <= layer2_outputs(2716);
    outputs(4415) <= not(layer2_outputs(1089));
    outputs(4416) <= not((layer2_outputs(2109)) and (layer2_outputs(3119)));
    outputs(4417) <= layer2_outputs(1115);
    outputs(4418) <= not(layer2_outputs(2651));
    outputs(4419) <= not(layer2_outputs(4442));
    outputs(4420) <= not(layer2_outputs(3026)) or (layer2_outputs(2499));
    outputs(4421) <= layer2_outputs(2550);
    outputs(4422) <= not(layer2_outputs(4128));
    outputs(4423) <= (layer2_outputs(1942)) and not (layer2_outputs(3770));
    outputs(4424) <= (layer2_outputs(2872)) xor (layer2_outputs(3341));
    outputs(4425) <= not(layer2_outputs(5012));
    outputs(4426) <= layer2_outputs(2498);
    outputs(4427) <= (layer2_outputs(1691)) and not (layer2_outputs(3185));
    outputs(4428) <= (layer2_outputs(1583)) and not (layer2_outputs(4349));
    outputs(4429) <= layer2_outputs(1277);
    outputs(4430) <= not(layer2_outputs(1395));
    outputs(4431) <= (layer2_outputs(574)) and not (layer2_outputs(3502));
    outputs(4432) <= layer2_outputs(2938);
    outputs(4433) <= layer2_outputs(915);
    outputs(4434) <= layer2_outputs(2237);
    outputs(4435) <= (layer2_outputs(773)) and not (layer2_outputs(946));
    outputs(4436) <= layer2_outputs(3974);
    outputs(4437) <= (layer2_outputs(1792)) xor (layer2_outputs(4222));
    outputs(4438) <= (layer2_outputs(721)) xor (layer2_outputs(296));
    outputs(4439) <= not(layer2_outputs(2823));
    outputs(4440) <= layer2_outputs(861);
    outputs(4441) <= not((layer2_outputs(1143)) or (layer2_outputs(3651)));
    outputs(4442) <= not(layer2_outputs(669));
    outputs(4443) <= (layer2_outputs(2947)) and not (layer2_outputs(3388));
    outputs(4444) <= layer2_outputs(3699);
    outputs(4445) <= not((layer2_outputs(4701)) xor (layer2_outputs(1612)));
    outputs(4446) <= (layer2_outputs(1312)) xor (layer2_outputs(3794));
    outputs(4447) <= not((layer2_outputs(485)) and (layer2_outputs(4441)));
    outputs(4448) <= (layer2_outputs(1833)) xor (layer2_outputs(3236));
    outputs(4449) <= not(layer2_outputs(2898));
    outputs(4450) <= not(layer2_outputs(3314));
    outputs(4451) <= (layer2_outputs(5092)) and not (layer2_outputs(2147));
    outputs(4452) <= not(layer2_outputs(297)) or (layer2_outputs(3110));
    outputs(4453) <= layer2_outputs(86);
    outputs(4454) <= not(layer2_outputs(832)) or (layer2_outputs(3390));
    outputs(4455) <= (layer2_outputs(908)) or (layer2_outputs(895));
    outputs(4456) <= layer2_outputs(2239);
    outputs(4457) <= not(layer2_outputs(4266));
    outputs(4458) <= layer2_outputs(251);
    outputs(4459) <= layer2_outputs(836);
    outputs(4460) <= not((layer2_outputs(3670)) and (layer2_outputs(3261)));
    outputs(4461) <= layer2_outputs(2850);
    outputs(4462) <= not(layer2_outputs(3426));
    outputs(4463) <= (layer2_outputs(1405)) xor (layer2_outputs(3294));
    outputs(4464) <= (layer2_outputs(2347)) and not (layer2_outputs(3815));
    outputs(4465) <= (layer2_outputs(4714)) and (layer2_outputs(1079));
    outputs(4466) <= layer2_outputs(4498);
    outputs(4467) <= layer2_outputs(4685);
    outputs(4468) <= not(layer2_outputs(2357)) or (layer2_outputs(3221));
    outputs(4469) <= layer2_outputs(4421);
    outputs(4470) <= layer2_outputs(2627);
    outputs(4471) <= not((layer2_outputs(342)) and (layer2_outputs(1552)));
    outputs(4472) <= (layer2_outputs(704)) or (layer2_outputs(3129));
    outputs(4473) <= (layer2_outputs(2884)) and not (layer2_outputs(2875));
    outputs(4474) <= layer2_outputs(3703);
    outputs(4475) <= not((layer2_outputs(3800)) and (layer2_outputs(3038)));
    outputs(4476) <= not((layer2_outputs(584)) xor (layer2_outputs(1641)));
    outputs(4477) <= layer2_outputs(3237);
    outputs(4478) <= not(layer2_outputs(3778));
    outputs(4479) <= not((layer2_outputs(3540)) or (layer2_outputs(919)));
    outputs(4480) <= not((layer2_outputs(2034)) xor (layer2_outputs(4451)));
    outputs(4481) <= (layer2_outputs(635)) xor (layer2_outputs(5093));
    outputs(4482) <= not(layer2_outputs(1040)) or (layer2_outputs(4948));
    outputs(4483) <= layer2_outputs(1421);
    outputs(4484) <= (layer2_outputs(4300)) and (layer2_outputs(2977));
    outputs(4485) <= layer2_outputs(707);
    outputs(4486) <= not((layer2_outputs(1873)) xor (layer2_outputs(2227)));
    outputs(4487) <= layer2_outputs(3420);
    outputs(4488) <= not(layer2_outputs(649));
    outputs(4489) <= not(layer2_outputs(1044));
    outputs(4490) <= not(layer2_outputs(3029));
    outputs(4491) <= not(layer2_outputs(1445));
    outputs(4492) <= (layer2_outputs(4012)) xor (layer2_outputs(1553));
    outputs(4493) <= (layer2_outputs(4663)) xor (layer2_outputs(1969));
    outputs(4494) <= layer2_outputs(1576);
    outputs(4495) <= not(layer2_outputs(665));
    outputs(4496) <= (layer2_outputs(1896)) xor (layer2_outputs(3232));
    outputs(4497) <= not(layer2_outputs(1204));
    outputs(4498) <= not(layer2_outputs(1390));
    outputs(4499) <= not(layer2_outputs(3001)) or (layer2_outputs(4299));
    outputs(4500) <= layer2_outputs(798);
    outputs(4501) <= layer2_outputs(4829);
    outputs(4502) <= not(layer2_outputs(999));
    outputs(4503) <= layer2_outputs(852);
    outputs(4504) <= (layer2_outputs(1347)) xor (layer2_outputs(3448));
    outputs(4505) <= not(layer2_outputs(351));
    outputs(4506) <= not(layer2_outputs(279));
    outputs(4507) <= not((layer2_outputs(2005)) xor (layer2_outputs(3549)));
    outputs(4508) <= layer2_outputs(4533);
    outputs(4509) <= (layer2_outputs(4964)) or (layer2_outputs(3598));
    outputs(4510) <= layer2_outputs(4733);
    outputs(4511) <= not(layer2_outputs(1477)) or (layer2_outputs(862));
    outputs(4512) <= not((layer2_outputs(315)) xor (layer2_outputs(140)));
    outputs(4513) <= not(layer2_outputs(318));
    outputs(4514) <= not(layer2_outputs(4194));
    outputs(4515) <= layer2_outputs(2956);
    outputs(4516) <= not(layer2_outputs(4680));
    outputs(4517) <= layer2_outputs(4133);
    outputs(4518) <= not(layer2_outputs(907));
    outputs(4519) <= (layer2_outputs(3171)) xor (layer2_outputs(2576));
    outputs(4520) <= not(layer2_outputs(835));
    outputs(4521) <= not(layer2_outputs(1514)) or (layer2_outputs(1609));
    outputs(4522) <= layer2_outputs(816);
    outputs(4523) <= layer2_outputs(4267);
    outputs(4524) <= not(layer2_outputs(2292));
    outputs(4525) <= layer2_outputs(2151);
    outputs(4526) <= not(layer2_outputs(3146));
    outputs(4527) <= not(layer2_outputs(4800));
    outputs(4528) <= (layer2_outputs(2057)) xor (layer2_outputs(3658));
    outputs(4529) <= layer2_outputs(746);
    outputs(4530) <= not(layer2_outputs(3604));
    outputs(4531) <= not(layer2_outputs(180));
    outputs(4532) <= not(layer2_outputs(4090));
    outputs(4533) <= not(layer2_outputs(428));
    outputs(4534) <= not((layer2_outputs(298)) and (layer2_outputs(1984)));
    outputs(4535) <= not(layer2_outputs(3409));
    outputs(4536) <= not(layer2_outputs(1367));
    outputs(4537) <= not(layer2_outputs(154));
    outputs(4538) <= not(layer2_outputs(4041));
    outputs(4539) <= not(layer2_outputs(4031)) or (layer2_outputs(1167));
    outputs(4540) <= not((layer2_outputs(573)) xor (layer2_outputs(2756)));
    outputs(4541) <= layer2_outputs(1181);
    outputs(4542) <= layer2_outputs(3424);
    outputs(4543) <= not(layer2_outputs(2408));
    outputs(4544) <= (layer2_outputs(2619)) xor (layer2_outputs(3557));
    outputs(4545) <= not(layer2_outputs(3198)) or (layer2_outputs(2427));
    outputs(4546) <= not(layer2_outputs(2381));
    outputs(4547) <= not((layer2_outputs(2718)) or (layer2_outputs(2547)));
    outputs(4548) <= layer2_outputs(405);
    outputs(4549) <= not(layer2_outputs(1403));
    outputs(4550) <= (layer2_outputs(2999)) xor (layer2_outputs(1480));
    outputs(4551) <= (layer2_outputs(1518)) and not (layer2_outputs(2817));
    outputs(4552) <= layer2_outputs(362);
    outputs(4553) <= layer2_outputs(2800);
    outputs(4554) <= layer2_outputs(2);
    outputs(4555) <= layer2_outputs(3004);
    outputs(4556) <= not((layer2_outputs(4916)) or (layer2_outputs(1909)));
    outputs(4557) <= layer2_outputs(4546);
    outputs(4558) <= (layer2_outputs(3233)) and not (layer2_outputs(4132));
    outputs(4559) <= not(layer2_outputs(2318));
    outputs(4560) <= (layer2_outputs(4251)) or (layer2_outputs(3300));
    outputs(4561) <= layer2_outputs(3246);
    outputs(4562) <= layer2_outputs(2707);
    outputs(4563) <= (layer2_outputs(1809)) xor (layer2_outputs(240));
    outputs(4564) <= layer2_outputs(4244);
    outputs(4565) <= (layer2_outputs(4543)) or (layer2_outputs(5009));
    outputs(4566) <= not(layer2_outputs(3405));
    outputs(4567) <= layer2_outputs(2329);
    outputs(4568) <= layer2_outputs(3528);
    outputs(4569) <= layer2_outputs(1282);
    outputs(4570) <= not(layer2_outputs(4062));
    outputs(4571) <= (layer2_outputs(345)) and not (layer2_outputs(1675));
    outputs(4572) <= layer2_outputs(4885);
    outputs(4573) <= not(layer2_outputs(3232)) or (layer2_outputs(3102));
    outputs(4574) <= (layer2_outputs(3705)) xor (layer2_outputs(4819));
    outputs(4575) <= layer2_outputs(570);
    outputs(4576) <= (layer2_outputs(792)) or (layer2_outputs(1528));
    outputs(4577) <= (layer2_outputs(3386)) xor (layer2_outputs(221));
    outputs(4578) <= (layer2_outputs(329)) and not (layer2_outputs(2173));
    outputs(4579) <= not(layer2_outputs(1951)) or (layer2_outputs(149));
    outputs(4580) <= (layer2_outputs(2860)) and (layer2_outputs(4654));
    outputs(4581) <= (layer2_outputs(2997)) or (layer2_outputs(1980));
    outputs(4582) <= layer2_outputs(3024);
    outputs(4583) <= not(layer2_outputs(4995));
    outputs(4584) <= (layer2_outputs(2146)) and not (layer2_outputs(2127));
    outputs(4585) <= not((layer2_outputs(5035)) xor (layer2_outputs(2873)));
    outputs(4586) <= layer2_outputs(2307);
    outputs(4587) <= layer2_outputs(476);
    outputs(4588) <= not((layer2_outputs(2077)) xor (layer2_outputs(4745)));
    outputs(4589) <= not(layer2_outputs(4336)) or (layer2_outputs(1643));
    outputs(4590) <= not(layer2_outputs(801));
    outputs(4591) <= (layer2_outputs(1615)) xor (layer2_outputs(427));
    outputs(4592) <= (layer2_outputs(548)) and not (layer2_outputs(2028));
    outputs(4593) <= not(layer2_outputs(610));
    outputs(4594) <= layer2_outputs(314);
    outputs(4595) <= layer2_outputs(2355);
    outputs(4596) <= not((layer2_outputs(3457)) xor (layer2_outputs(4971)));
    outputs(4597) <= not(layer2_outputs(1259));
    outputs(4598) <= not(layer2_outputs(3876));
    outputs(4599) <= layer2_outputs(4966);
    outputs(4600) <= not((layer2_outputs(2302)) and (layer2_outputs(2741)));
    outputs(4601) <= (layer2_outputs(4195)) xor (layer2_outputs(1469));
    outputs(4602) <= (layer2_outputs(3249)) and not (layer2_outputs(898));
    outputs(4603) <= not((layer2_outputs(1107)) xor (layer2_outputs(3643)));
    outputs(4604) <= not(layer2_outputs(310));
    outputs(4605) <= (layer2_outputs(2977)) xor (layer2_outputs(4114));
    outputs(4606) <= layer2_outputs(5017);
    outputs(4607) <= not((layer2_outputs(348)) xor (layer2_outputs(1399)));
    outputs(4608) <= (layer2_outputs(564)) or (layer2_outputs(3213));
    outputs(4609) <= (layer2_outputs(3753)) and not (layer2_outputs(708));
    outputs(4610) <= not((layer2_outputs(4375)) xor (layer2_outputs(3027)));
    outputs(4611) <= (layer2_outputs(4031)) and (layer2_outputs(1352));
    outputs(4612) <= layer2_outputs(2761);
    outputs(4613) <= not(layer2_outputs(1449));
    outputs(4614) <= layer2_outputs(1688);
    outputs(4615) <= layer2_outputs(2660);
    outputs(4616) <= layer2_outputs(5056);
    outputs(4617) <= layer2_outputs(3506);
    outputs(4618) <= layer2_outputs(1068);
    outputs(4619) <= not(layer2_outputs(1216));
    outputs(4620) <= layer2_outputs(1014);
    outputs(4621) <= not(layer2_outputs(1699));
    outputs(4622) <= (layer2_outputs(1776)) and not (layer2_outputs(2899));
    outputs(4623) <= not((layer2_outputs(2527)) xor (layer2_outputs(3246)));
    outputs(4624) <= layer2_outputs(2211);
    outputs(4625) <= not(layer2_outputs(603));
    outputs(4626) <= not((layer2_outputs(1533)) xor (layer2_outputs(706)));
    outputs(4627) <= not((layer2_outputs(4575)) and (layer2_outputs(5065)));
    outputs(4628) <= layer2_outputs(2575);
    outputs(4629) <= layer2_outputs(2698);
    outputs(4630) <= not(layer2_outputs(1983));
    outputs(4631) <= not((layer2_outputs(1747)) and (layer2_outputs(2568)));
    outputs(4632) <= (layer2_outputs(3086)) and not (layer2_outputs(483));
    outputs(4633) <= not((layer2_outputs(4944)) xor (layer2_outputs(1116)));
    outputs(4634) <= not(layer2_outputs(3079));
    outputs(4635) <= layer2_outputs(3942);
    outputs(4636) <= not((layer2_outputs(1857)) and (layer2_outputs(4151)));
    outputs(4637) <= not((layer2_outputs(383)) xor (layer2_outputs(2393)));
    outputs(4638) <= not(layer2_outputs(1336)) or (layer2_outputs(2697));
    outputs(4639) <= not((layer2_outputs(1257)) or (layer2_outputs(483)));
    outputs(4640) <= not(layer2_outputs(4307));
    outputs(4641) <= layer2_outputs(1848);
    outputs(4642) <= not((layer2_outputs(2367)) or (layer2_outputs(4731)));
    outputs(4643) <= not(layer2_outputs(2324));
    outputs(4644) <= (layer2_outputs(2180)) xor (layer2_outputs(524));
    outputs(4645) <= not(layer2_outputs(2323));
    outputs(4646) <= (layer2_outputs(1396)) xor (layer2_outputs(2912));
    outputs(4647) <= layer2_outputs(3342);
    outputs(4648) <= (layer2_outputs(556)) and not (layer2_outputs(2699));
    outputs(4649) <= not(layer2_outputs(1571));
    outputs(4650) <= not(layer2_outputs(2777));
    outputs(4651) <= (layer2_outputs(2023)) and not (layer2_outputs(2634));
    outputs(4652) <= not((layer2_outputs(868)) or (layer2_outputs(254)));
    outputs(4653) <= (layer2_outputs(4721)) and not (layer2_outputs(3165));
    outputs(4654) <= not(layer2_outputs(2019));
    outputs(4655) <= not(layer2_outputs(2259));
    outputs(4656) <= not((layer2_outputs(4448)) or (layer2_outputs(4223)));
    outputs(4657) <= not(layer2_outputs(2483));
    outputs(4658) <= layer2_outputs(2160);
    outputs(4659) <= layer2_outputs(842);
    outputs(4660) <= layer2_outputs(3086);
    outputs(4661) <= layer2_outputs(2046);
    outputs(4662) <= (layer2_outputs(3162)) or (layer2_outputs(3964));
    outputs(4663) <= layer2_outputs(3448);
    outputs(4664) <= (layer2_outputs(902)) and not (layer2_outputs(1478));
    outputs(4665) <= layer2_outputs(2547);
    outputs(4666) <= (layer2_outputs(2972)) and not (layer2_outputs(2798));
    outputs(4667) <= not(layer2_outputs(3043));
    outputs(4668) <= (layer2_outputs(2675)) xor (layer2_outputs(4908));
    outputs(4669) <= not((layer2_outputs(998)) or (layer2_outputs(43)));
    outputs(4670) <= not(layer2_outputs(2017));
    outputs(4671) <= (layer2_outputs(3703)) xor (layer2_outputs(2765));
    outputs(4672) <= not(layer2_outputs(3995));
    outputs(4673) <= not((layer2_outputs(2310)) or (layer2_outputs(2531)));
    outputs(4674) <= not(layer2_outputs(3102)) or (layer2_outputs(5044));
    outputs(4675) <= not(layer2_outputs(2483));
    outputs(4676) <= not(layer2_outputs(1471));
    outputs(4677) <= (layer2_outputs(4587)) and (layer2_outputs(743));
    outputs(4678) <= (layer2_outputs(1671)) and (layer2_outputs(4641));
    outputs(4679) <= not(layer2_outputs(1800));
    outputs(4680) <= layer2_outputs(549);
    outputs(4681) <= layer2_outputs(2216);
    outputs(4682) <= (layer2_outputs(2496)) and (layer2_outputs(795));
    outputs(4683) <= layer2_outputs(754);
    outputs(4684) <= not(layer2_outputs(3619));
    outputs(4685) <= layer2_outputs(769);
    outputs(4686) <= (layer2_outputs(3898)) and not (layer2_outputs(157));
    outputs(4687) <= not((layer2_outputs(4548)) xor (layer2_outputs(412)));
    outputs(4688) <= layer2_outputs(1451);
    outputs(4689) <= not((layer2_outputs(5074)) or (layer2_outputs(1214)));
    outputs(4690) <= (layer2_outputs(3456)) and not (layer2_outputs(1673));
    outputs(4691) <= not(layer2_outputs(4457));
    outputs(4692) <= (layer2_outputs(2998)) and (layer2_outputs(3130));
    outputs(4693) <= (layer2_outputs(3393)) and (layer2_outputs(1121));
    outputs(4694) <= (layer2_outputs(1427)) and not (layer2_outputs(2804));
    outputs(4695) <= layer2_outputs(643);
    outputs(4696) <= (layer2_outputs(2799)) xor (layer2_outputs(4518));
    outputs(4697) <= not(layer2_outputs(979));
    outputs(4698) <= layer2_outputs(380);
    outputs(4699) <= not(layer2_outputs(2051));
    outputs(4700) <= not(layer2_outputs(2797));
    outputs(4701) <= layer2_outputs(4351);
    outputs(4702) <= not((layer2_outputs(1140)) xor (layer2_outputs(1854)));
    outputs(4703) <= not((layer2_outputs(2102)) xor (layer2_outputs(4558)));
    outputs(4704) <= layer2_outputs(3381);
    outputs(4705) <= layer2_outputs(473);
    outputs(4706) <= layer2_outputs(1908);
    outputs(4707) <= not(layer2_outputs(1936));
    outputs(4708) <= (layer2_outputs(4262)) xor (layer2_outputs(4923));
    outputs(4709) <= (layer2_outputs(447)) and not (layer2_outputs(1221));
    outputs(4710) <= not((layer2_outputs(4707)) xor (layer2_outputs(4516)));
    outputs(4711) <= layer2_outputs(1374);
    outputs(4712) <= not(layer2_outputs(1859));
    outputs(4713) <= (layer2_outputs(2574)) xor (layer2_outputs(4020));
    outputs(4714) <= not(layer2_outputs(960));
    outputs(4715) <= layer2_outputs(3566);
    outputs(4716) <= not((layer2_outputs(1812)) or (layer2_outputs(4219)));
    outputs(4717) <= not((layer2_outputs(1865)) or (layer2_outputs(2467)));
    outputs(4718) <= (layer2_outputs(1778)) and not (layer2_outputs(460));
    outputs(4719) <= layer2_outputs(961);
    outputs(4720) <= layer2_outputs(4735);
    outputs(4721) <= layer2_outputs(2846);
    outputs(4722) <= not(layer2_outputs(738));
    outputs(4723) <= not((layer2_outputs(3774)) xor (layer2_outputs(2043)));
    outputs(4724) <= not((layer2_outputs(595)) xor (layer2_outputs(1930)));
    outputs(4725) <= not(layer2_outputs(2375));
    outputs(4726) <= not(layer2_outputs(3565));
    outputs(4727) <= not(layer2_outputs(5100));
    outputs(4728) <= (layer2_outputs(3256)) and not (layer2_outputs(2132));
    outputs(4729) <= layer2_outputs(3477);
    outputs(4730) <= not(layer2_outputs(2833));
    outputs(4731) <= not(layer2_outputs(4367));
    outputs(4732) <= (layer2_outputs(1111)) xor (layer2_outputs(2902));
    outputs(4733) <= not(layer2_outputs(4215));
    outputs(4734) <= (layer2_outputs(1014)) and (layer2_outputs(168));
    outputs(4735) <= (layer2_outputs(2258)) or (layer2_outputs(3781));
    outputs(4736) <= layer2_outputs(2518);
    outputs(4737) <= layer2_outputs(1469);
    outputs(4738) <= (layer2_outputs(2027)) and not (layer2_outputs(1392));
    outputs(4739) <= layer2_outputs(2584);
    outputs(4740) <= not(layer2_outputs(575));
    outputs(4741) <= not(layer2_outputs(1401)) or (layer2_outputs(753));
    outputs(4742) <= not((layer2_outputs(2311)) xor (layer2_outputs(674)));
    outputs(4743) <= not(layer2_outputs(1639));
    outputs(4744) <= not(layer2_outputs(2186));
    outputs(4745) <= not(layer2_outputs(5097));
    outputs(4746) <= not((layer2_outputs(1750)) xor (layer2_outputs(649)));
    outputs(4747) <= layer2_outputs(1388);
    outputs(4748) <= not(layer2_outputs(1437));
    outputs(4749) <= not(layer2_outputs(2463));
    outputs(4750) <= (layer2_outputs(4802)) xor (layer2_outputs(4933));
    outputs(4751) <= (layer2_outputs(3189)) and not (layer2_outputs(1529));
    outputs(4752) <= layer2_outputs(1840);
    outputs(4753) <= layer2_outputs(2204);
    outputs(4754) <= '1';
    outputs(4755) <= (layer2_outputs(4049)) and not (layer2_outputs(1790));
    outputs(4756) <= not(layer2_outputs(2618));
    outputs(4757) <= layer2_outputs(5007);
    outputs(4758) <= layer2_outputs(3685);
    outputs(4759) <= layer2_outputs(865);
    outputs(4760) <= layer2_outputs(4077);
    outputs(4761) <= not((layer2_outputs(5053)) xor (layer2_outputs(2787)));
    outputs(4762) <= layer2_outputs(2157);
    outputs(4763) <= not((layer2_outputs(2654)) or (layer2_outputs(2620)));
    outputs(4764) <= not(layer2_outputs(2893));
    outputs(4765) <= (layer2_outputs(386)) and (layer2_outputs(1726));
    outputs(4766) <= layer2_outputs(2299);
    outputs(4767) <= not((layer2_outputs(1195)) xor (layer2_outputs(2158)));
    outputs(4768) <= (layer2_outputs(3124)) and (layer2_outputs(918));
    outputs(4769) <= not(layer2_outputs(216));
    outputs(4770) <= not((layer2_outputs(4659)) or (layer2_outputs(2395)));
    outputs(4771) <= not(layer2_outputs(1321));
    outputs(4772) <= (layer2_outputs(4)) and not (layer2_outputs(3243));
    outputs(4773) <= not(layer2_outputs(1554));
    outputs(4774) <= (layer2_outputs(4510)) and not (layer2_outputs(2215));
    outputs(4775) <= (layer2_outputs(5011)) and not (layer2_outputs(1690));
    outputs(4776) <= not(layer2_outputs(3742));
    outputs(4777) <= not(layer2_outputs(5004));
    outputs(4778) <= not(layer2_outputs(948));
    outputs(4779) <= not((layer2_outputs(4434)) and (layer2_outputs(4709)));
    outputs(4780) <= (layer2_outputs(991)) and (layer2_outputs(5014));
    outputs(4781) <= layer2_outputs(4685);
    outputs(4782) <= (layer2_outputs(3498)) and (layer2_outputs(1456));
    outputs(4783) <= (layer2_outputs(3689)) xor (layer2_outputs(319));
    outputs(4784) <= (layer2_outputs(2228)) xor (layer2_outputs(1568));
    outputs(4785) <= layer2_outputs(2044);
    outputs(4786) <= layer2_outputs(4722);
    outputs(4787) <= not(layer2_outputs(4087));
    outputs(4788) <= not(layer2_outputs(1800)) or (layer2_outputs(2640));
    outputs(4789) <= layer2_outputs(4453);
    outputs(4790) <= layer2_outputs(2838);
    outputs(4791) <= layer2_outputs(3259);
    outputs(4792) <= (layer2_outputs(1618)) xor (layer2_outputs(434));
    outputs(4793) <= not(layer2_outputs(4180));
    outputs(4794) <= layer2_outputs(3234);
    outputs(4795) <= layer2_outputs(1502);
    outputs(4796) <= layer2_outputs(1923);
    outputs(4797) <= not((layer2_outputs(15)) xor (layer2_outputs(768)));
    outputs(4798) <= not((layer2_outputs(3804)) xor (layer2_outputs(477)));
    outputs(4799) <= not(layer2_outputs(4840));
    outputs(4800) <= not(layer2_outputs(3751));
    outputs(4801) <= not((layer2_outputs(2649)) or (layer2_outputs(4529)));
    outputs(4802) <= not(layer2_outputs(3069));
    outputs(4803) <= not(layer2_outputs(4161));
    outputs(4804) <= not((layer2_outputs(3683)) xor (layer2_outputs(619)));
    outputs(4805) <= (layer2_outputs(168)) xor (layer2_outputs(1561));
    outputs(4806) <= layer2_outputs(3873);
    outputs(4807) <= layer2_outputs(2612);
    outputs(4808) <= not(layer2_outputs(522));
    outputs(4809) <= not((layer2_outputs(2705)) xor (layer2_outputs(4727)));
    outputs(4810) <= (layer2_outputs(3356)) and not (layer2_outputs(4655));
    outputs(4811) <= (layer2_outputs(4508)) and not (layer2_outputs(4379));
    outputs(4812) <= not((layer2_outputs(2864)) xor (layer2_outputs(1736)));
    outputs(4813) <= not((layer2_outputs(3555)) xor (layer2_outputs(503)));
    outputs(4814) <= (layer2_outputs(2106)) xor (layer2_outputs(4838));
    outputs(4815) <= not(layer2_outputs(2294));
    outputs(4816) <= not((layer2_outputs(1789)) xor (layer2_outputs(2338)));
    outputs(4817) <= (layer2_outputs(2671)) or (layer2_outputs(2727));
    outputs(4818) <= layer2_outputs(559);
    outputs(4819) <= not(layer2_outputs(4996));
    outputs(4820) <= not((layer2_outputs(4769)) or (layer2_outputs(1630)));
    outputs(4821) <= layer2_outputs(3032);
    outputs(4822) <= layer2_outputs(3533);
    outputs(4823) <= not(layer2_outputs(4535));
    outputs(4824) <= layer2_outputs(951);
    outputs(4825) <= not(layer2_outputs(486));
    outputs(4826) <= layer2_outputs(4860);
    outputs(4827) <= not(layer2_outputs(2114));
    outputs(4828) <= (layer2_outputs(1420)) xor (layer2_outputs(2539));
    outputs(4829) <= (layer2_outputs(1488)) or (layer2_outputs(984));
    outputs(4830) <= not(layer2_outputs(1197));
    outputs(4831) <= layer2_outputs(2481);
    outputs(4832) <= not((layer2_outputs(3332)) xor (layer2_outputs(1056)));
    outputs(4833) <= (layer2_outputs(1878)) xor (layer2_outputs(925));
    outputs(4834) <= (layer2_outputs(4520)) xor (layer2_outputs(1432));
    outputs(4835) <= not((layer2_outputs(2515)) xor (layer2_outputs(3716)));
    outputs(4836) <= not(layer2_outputs(1839));
    outputs(4837) <= layer2_outputs(4249);
    outputs(4838) <= (layer2_outputs(2955)) and not (layer2_outputs(2680));
    outputs(4839) <= not((layer2_outputs(5024)) xor (layer2_outputs(2029)));
    outputs(4840) <= not(layer2_outputs(1321));
    outputs(4841) <= layer2_outputs(2890);
    outputs(4842) <= not((layer2_outputs(4769)) or (layer2_outputs(4871)));
    outputs(4843) <= layer2_outputs(408);
    outputs(4844) <= layer2_outputs(4770);
    outputs(4845) <= not(layer2_outputs(762));
    outputs(4846) <= not(layer2_outputs(2552));
    outputs(4847) <= not(layer2_outputs(3752));
    outputs(4848) <= not(layer2_outputs(2578));
    outputs(4849) <= layer2_outputs(1363);
    outputs(4850) <= layer2_outputs(4458);
    outputs(4851) <= (layer2_outputs(1883)) and not (layer2_outputs(633));
    outputs(4852) <= layer2_outputs(1300);
    outputs(4853) <= (layer2_outputs(4274)) and not (layer2_outputs(2717));
    outputs(4854) <= (layer2_outputs(3976)) and not (layer2_outputs(4771));
    outputs(4855) <= not(layer2_outputs(4852));
    outputs(4856) <= not(layer2_outputs(3765));
    outputs(4857) <= layer2_outputs(3133);
    outputs(4858) <= layer2_outputs(4485);
    outputs(4859) <= (layer2_outputs(2432)) and not (layer2_outputs(3632));
    outputs(4860) <= (layer2_outputs(3048)) and not (layer2_outputs(2577));
    outputs(4861) <= not(layer2_outputs(985));
    outputs(4862) <= not((layer2_outputs(3022)) or (layer2_outputs(3727)));
    outputs(4863) <= not(layer2_outputs(3333));
    outputs(4864) <= not(layer2_outputs(2267));
    outputs(4865) <= not((layer2_outputs(4134)) xor (layer2_outputs(3628)));
    outputs(4866) <= layer2_outputs(4225);
    outputs(4867) <= not(layer2_outputs(161));
    outputs(4868) <= (layer2_outputs(302)) and not (layer2_outputs(5005));
    outputs(4869) <= not(layer2_outputs(2275)) or (layer2_outputs(2973));
    outputs(4870) <= layer2_outputs(3199);
    outputs(4871) <= not(layer2_outputs(1241)) or (layer2_outputs(1477));
    outputs(4872) <= (layer2_outputs(3569)) xor (layer2_outputs(3413));
    outputs(4873) <= not(layer2_outputs(3886));
    outputs(4874) <= not(layer2_outputs(1828)) or (layer2_outputs(1721));
    outputs(4875) <= layer2_outputs(4627);
    outputs(4876) <= (layer2_outputs(2849)) xor (layer2_outputs(1101));
    outputs(4877) <= not(layer2_outputs(3158));
    outputs(4878) <= not(layer2_outputs(2528));
    outputs(4879) <= not(layer2_outputs(1070));
    outputs(4880) <= (layer2_outputs(228)) or (layer2_outputs(3669));
    outputs(4881) <= not(layer2_outputs(2802));
    outputs(4882) <= layer2_outputs(2250);
    outputs(4883) <= layer2_outputs(4956);
    outputs(4884) <= layer2_outputs(227);
    outputs(4885) <= (layer2_outputs(349)) xor (layer2_outputs(2599));
    outputs(4886) <= (layer2_outputs(3371)) and (layer2_outputs(4915));
    outputs(4887) <= (layer2_outputs(4967)) and not (layer2_outputs(4935));
    outputs(4888) <= not((layer2_outputs(3205)) or (layer2_outputs(3295)));
    outputs(4889) <= layer2_outputs(107);
    outputs(4890) <= not(layer2_outputs(4720));
    outputs(4891) <= (layer2_outputs(1154)) xor (layer2_outputs(5019));
    outputs(4892) <= layer2_outputs(3675);
    outputs(4893) <= not(layer2_outputs(2923));
    outputs(4894) <= not((layer2_outputs(3126)) xor (layer2_outputs(4246)));
    outputs(4895) <= not((layer2_outputs(1201)) xor (layer2_outputs(2920)));
    outputs(4896) <= (layer2_outputs(279)) and not (layer2_outputs(3653));
    outputs(4897) <= layer2_outputs(4122);
    outputs(4898) <= (layer2_outputs(2473)) and not (layer2_outputs(2420));
    outputs(4899) <= layer2_outputs(4665);
    outputs(4900) <= layer2_outputs(3760);
    outputs(4901) <= not((layer2_outputs(4585)) or (layer2_outputs(2730)));
    outputs(4902) <= not((layer2_outputs(638)) xor (layer2_outputs(468)));
    outputs(4903) <= layer2_outputs(283);
    outputs(4904) <= not(layer2_outputs(4864));
    outputs(4905) <= not(layer2_outputs(2777));
    outputs(4906) <= (layer2_outputs(4958)) and (layer2_outputs(82));
    outputs(4907) <= not(layer2_outputs(2278));
    outputs(4908) <= (layer2_outputs(1231)) and not (layer2_outputs(2254));
    outputs(4909) <= layer2_outputs(573);
    outputs(4910) <= (layer2_outputs(3195)) xor (layer2_outputs(5110));
    outputs(4911) <= not((layer2_outputs(418)) xor (layer2_outputs(1568)));
    outputs(4912) <= layer2_outputs(2826);
    outputs(4913) <= (layer2_outputs(2152)) xor (layer2_outputs(315));
    outputs(4914) <= layer2_outputs(817);
    outputs(4915) <= not((layer2_outputs(1831)) xor (layer2_outputs(2490)));
    outputs(4916) <= not(layer2_outputs(4697)) or (layer2_outputs(3034));
    outputs(4917) <= not((layer2_outputs(3938)) xor (layer2_outputs(3204)));
    outputs(4918) <= layer2_outputs(3947);
    outputs(4919) <= layer2_outputs(818);
    outputs(4920) <= layer2_outputs(3374);
    outputs(4921) <= not((layer2_outputs(4539)) xor (layer2_outputs(3465)));
    outputs(4922) <= not(layer2_outputs(4429));
    outputs(4923) <= (layer2_outputs(3117)) and not (layer2_outputs(2303));
    outputs(4924) <= (layer2_outputs(4286)) xor (layer2_outputs(4265));
    outputs(4925) <= layer2_outputs(2883);
    outputs(4926) <= (layer2_outputs(2145)) xor (layer2_outputs(4144));
    outputs(4927) <= not((layer2_outputs(3944)) or (layer2_outputs(4924)));
    outputs(4928) <= layer2_outputs(769);
    outputs(4929) <= layer2_outputs(1185);
    outputs(4930) <= not(layer2_outputs(4383));
    outputs(4931) <= not((layer2_outputs(531)) or (layer2_outputs(1824)));
    outputs(4932) <= (layer2_outputs(377)) and not (layer2_outputs(1616));
    outputs(4933) <= (layer2_outputs(2064)) xor (layer2_outputs(2087));
    outputs(4934) <= (layer2_outputs(4431)) and not (layer2_outputs(4230));
    outputs(4935) <= layer2_outputs(4378);
    outputs(4936) <= (layer2_outputs(3503)) xor (layer2_outputs(2987));
    outputs(4937) <= layer2_outputs(754);
    outputs(4938) <= layer2_outputs(4051);
    outputs(4939) <= (layer2_outputs(1427)) and not (layer2_outputs(1582));
    outputs(4940) <= not(layer2_outputs(306));
    outputs(4941) <= (layer2_outputs(1105)) xor (layer2_outputs(4567));
    outputs(4942) <= not(layer2_outputs(2340));
    outputs(4943) <= layer2_outputs(484);
    outputs(4944) <= layer2_outputs(1745);
    outputs(4945) <= not((layer2_outputs(4214)) xor (layer2_outputs(84)));
    outputs(4946) <= not(layer2_outputs(4528)) or (layer2_outputs(1550));
    outputs(4947) <= not(layer2_outputs(2602));
    outputs(4948) <= (layer2_outputs(3957)) and not (layer2_outputs(3380));
    outputs(4949) <= layer2_outputs(637);
    outputs(4950) <= not(layer2_outputs(1213));
    outputs(4951) <= not((layer2_outputs(4449)) xor (layer2_outputs(4961)));
    outputs(4952) <= (layer2_outputs(1549)) and not (layer2_outputs(4255));
    outputs(4953) <= not(layer2_outputs(4637));
    outputs(4954) <= not(layer2_outputs(4042));
    outputs(4955) <= not(layer2_outputs(3113));
    outputs(4956) <= layer2_outputs(1897);
    outputs(4957) <= layer2_outputs(3563);
    outputs(4958) <= layer2_outputs(1727);
    outputs(4959) <= not((layer2_outputs(3137)) and (layer2_outputs(4233)));
    outputs(4960) <= layer2_outputs(3040);
    outputs(4961) <= not(layer2_outputs(1646));
    outputs(4962) <= not((layer2_outputs(3833)) xor (layer2_outputs(999)));
    outputs(4963) <= not(layer2_outputs(3084));
    outputs(4964) <= (layer2_outputs(3152)) xor (layer2_outputs(2698));
    outputs(4965) <= not(layer2_outputs(4560));
    outputs(4966) <= not(layer2_outputs(3178));
    outputs(4967) <= not(layer2_outputs(4046)) or (layer2_outputs(3481));
    outputs(4968) <= layer2_outputs(3041);
    outputs(4969) <= not((layer2_outputs(4286)) xor (layer2_outputs(4888)));
    outputs(4970) <= (layer2_outputs(1932)) and not (layer2_outputs(2819));
    outputs(4971) <= layer2_outputs(332);
    outputs(4972) <= layer2_outputs(61);
    outputs(4973) <= layer2_outputs(4641);
    outputs(4974) <= layer2_outputs(1764);
    outputs(4975) <= not(layer2_outputs(1303));
    outputs(4976) <= layer2_outputs(4519);
    outputs(4977) <= not(layer2_outputs(3245));
    outputs(4978) <= layer2_outputs(506);
    outputs(4979) <= layer2_outputs(2850);
    outputs(4980) <= not(layer2_outputs(4470));
    outputs(4981) <= layer2_outputs(3363);
    outputs(4982) <= layer2_outputs(4168);
    outputs(4983) <= not(layer2_outputs(3879));
    outputs(4984) <= (layer2_outputs(3530)) xor (layer2_outputs(1829));
    outputs(4985) <= not(layer2_outputs(4626));
    outputs(4986) <= (layer2_outputs(1991)) xor (layer2_outputs(595));
    outputs(4987) <= not(layer2_outputs(4981));
    outputs(4988) <= (layer2_outputs(864)) and not (layer2_outputs(2953));
    outputs(4989) <= layer2_outputs(110);
    outputs(4990) <= layer2_outputs(2612);
    outputs(4991) <= layer2_outputs(3055);
    outputs(4992) <= not(layer2_outputs(3975));
    outputs(4993) <= not((layer2_outputs(1333)) xor (layer2_outputs(2857)));
    outputs(4994) <= (layer2_outputs(2641)) and not (layer2_outputs(1586));
    outputs(4995) <= not(layer2_outputs(1337));
    outputs(4996) <= layer2_outputs(506);
    outputs(4997) <= not(layer2_outputs(846));
    outputs(4998) <= (layer2_outputs(3850)) and not (layer2_outputs(4499));
    outputs(4999) <= not((layer2_outputs(1510)) xor (layer2_outputs(4228)));
    outputs(5000) <= layer2_outputs(338);
    outputs(5001) <= not(layer2_outputs(2970));
    outputs(5002) <= layer2_outputs(4777);
    outputs(5003) <= layer2_outputs(466);
    outputs(5004) <= (layer2_outputs(1256)) and not (layer2_outputs(381));
    outputs(5005) <= not(layer2_outputs(730));
    outputs(5006) <= not((layer2_outputs(1133)) or (layer2_outputs(1955)));
    outputs(5007) <= not(layer2_outputs(808));
    outputs(5008) <= layer2_outputs(743);
    outputs(5009) <= not((layer2_outputs(2409)) and (layer2_outputs(1631)));
    outputs(5010) <= (layer2_outputs(1199)) and not (layer2_outputs(4668));
    outputs(5011) <= not((layer2_outputs(3206)) xor (layer2_outputs(4952)));
    outputs(5012) <= not((layer2_outputs(3730)) xor (layer2_outputs(3783)));
    outputs(5013) <= not((layer2_outputs(510)) or (layer2_outputs(2784)));
    outputs(5014) <= not(layer2_outputs(142));
    outputs(5015) <= layer2_outputs(3278);
    outputs(5016) <= (layer2_outputs(848)) xor (layer2_outputs(2070));
    outputs(5017) <= layer2_outputs(3676);
    outputs(5018) <= not((layer2_outputs(3984)) xor (layer2_outputs(2746)));
    outputs(5019) <= (layer2_outputs(3767)) xor (layer2_outputs(942));
    outputs(5020) <= (layer2_outputs(1035)) xor (layer2_outputs(1627));
    outputs(5021) <= not((layer2_outputs(4914)) xor (layer2_outputs(3796)));
    outputs(5022) <= not(layer2_outputs(1162));
    outputs(5023) <= layer2_outputs(3398);
    outputs(5024) <= not(layer2_outputs(759));
    outputs(5025) <= not(layer2_outputs(4401));
    outputs(5026) <= not(layer2_outputs(1457));
    outputs(5027) <= layer2_outputs(1264);
    outputs(5028) <= (layer2_outputs(2200)) and not (layer2_outputs(4042));
    outputs(5029) <= not((layer2_outputs(1422)) or (layer2_outputs(244)));
    outputs(5030) <= not((layer2_outputs(3035)) or (layer2_outputs(2900)));
    outputs(5031) <= layer2_outputs(262);
    outputs(5032) <= layer2_outputs(4695);
    outputs(5033) <= layer2_outputs(763);
    outputs(5034) <= not(layer2_outputs(1474));
    outputs(5035) <= not(layer2_outputs(3231));
    outputs(5036) <= not(layer2_outputs(2283));
    outputs(5037) <= not((layer2_outputs(2061)) or (layer2_outputs(3488)));
    outputs(5038) <= layer2_outputs(3354);
    outputs(5039) <= layer2_outputs(763);
    outputs(5040) <= not(layer2_outputs(4256));
    outputs(5041) <= layer2_outputs(74);
    outputs(5042) <= (layer2_outputs(3411)) and not (layer2_outputs(4115));
    outputs(5043) <= not(layer2_outputs(1237));
    outputs(5044) <= not(layer2_outputs(2006));
    outputs(5045) <= not(layer2_outputs(4064));
    outputs(5046) <= (layer2_outputs(4903)) and not (layer2_outputs(4362));
    outputs(5047) <= (layer2_outputs(2010)) and (layer2_outputs(1476));
    outputs(5048) <= not(layer2_outputs(642));
    outputs(5049) <= not(layer2_outputs(2734));
    outputs(5050) <= layer2_outputs(2964);
    outputs(5051) <= not((layer2_outputs(3120)) xor (layer2_outputs(940)));
    outputs(5052) <= not(layer2_outputs(2272));
    outputs(5053) <= layer2_outputs(432);
    outputs(5054) <= layer2_outputs(4131);
    outputs(5055) <= not(layer2_outputs(2135));
    outputs(5056) <= layer2_outputs(2628);
    outputs(5057) <= (layer2_outputs(1842)) and not (layer2_outputs(5057));
    outputs(5058) <= (layer2_outputs(3645)) and not (layer2_outputs(4069));
    outputs(5059) <= not((layer2_outputs(4057)) and (layer2_outputs(542)));
    outputs(5060) <= not(layer2_outputs(3350));
    outputs(5061) <= not(layer2_outputs(3364));
    outputs(5062) <= not((layer2_outputs(5053)) xor (layer2_outputs(3539)));
    outputs(5063) <= not(layer2_outputs(1598));
    outputs(5064) <= layer2_outputs(2218);
    outputs(5065) <= not((layer2_outputs(2485)) xor (layer2_outputs(1013)));
    outputs(5066) <= (layer2_outputs(2380)) and not (layer2_outputs(681));
    outputs(5067) <= layer2_outputs(4943);
    outputs(5068) <= layer2_outputs(2368);
    outputs(5069) <= (layer2_outputs(3545)) xor (layer2_outputs(3790));
    outputs(5070) <= layer2_outputs(2042);
    outputs(5071) <= not(layer2_outputs(207)) or (layer2_outputs(1359));
    outputs(5072) <= (layer2_outputs(87)) or (layer2_outputs(3657));
    outputs(5073) <= (layer2_outputs(5034)) and not (layer2_outputs(3539));
    outputs(5074) <= (layer2_outputs(4189)) and not (layer2_outputs(461));
    outputs(5075) <= layer2_outputs(1126);
    outputs(5076) <= (layer2_outputs(4865)) and not (layer2_outputs(235));
    outputs(5077) <= (layer2_outputs(1483)) and not (layer2_outputs(2086));
    outputs(5078) <= not((layer2_outputs(3089)) or (layer2_outputs(4630)));
    outputs(5079) <= not(layer2_outputs(3287));
    outputs(5080) <= layer2_outputs(578);
    outputs(5081) <= not((layer2_outputs(3298)) xor (layer2_outputs(2557)));
    outputs(5082) <= not(layer2_outputs(2479));
    outputs(5083) <= not((layer2_outputs(2337)) xor (layer2_outputs(3438)));
    outputs(5084) <= not((layer2_outputs(3363)) xor (layer2_outputs(4440)));
    outputs(5085) <= (layer2_outputs(3338)) and not (layer2_outputs(2990));
    outputs(5086) <= (layer2_outputs(4965)) xor (layer2_outputs(2147));
    outputs(5087) <= (layer2_outputs(4562)) xor (layer2_outputs(4735));
    outputs(5088) <= (layer2_outputs(1865)) xor (layer2_outputs(2026));
    outputs(5089) <= layer2_outputs(3817);
    outputs(5090) <= layer2_outputs(4888);
    outputs(5091) <= not(layer2_outputs(3489)) or (layer2_outputs(4188));
    outputs(5092) <= not(layer2_outputs(5063));
    outputs(5093) <= not((layer2_outputs(3222)) or (layer2_outputs(1409)));
    outputs(5094) <= (layer2_outputs(1171)) and not (layer2_outputs(868));
    outputs(5095) <= layer2_outputs(4594);
    outputs(5096) <= layer2_outputs(74);
    outputs(5097) <= (layer2_outputs(4979)) and (layer2_outputs(1017));
    outputs(5098) <= not(layer2_outputs(561));
    outputs(5099) <= layer2_outputs(4066);
    outputs(5100) <= not(layer2_outputs(2868));
    outputs(5101) <= (layer2_outputs(1426)) and not (layer2_outputs(400));
    outputs(5102) <= not((layer2_outputs(3482)) xor (layer2_outputs(3478)));
    outputs(5103) <= not(layer2_outputs(4105));
    outputs(5104) <= (layer2_outputs(4127)) and not (layer2_outputs(4630));
    outputs(5105) <= not(layer2_outputs(1241));
    outputs(5106) <= layer2_outputs(3595);
    outputs(5107) <= layer2_outputs(1600);
    outputs(5108) <= not((layer2_outputs(2763)) xor (layer2_outputs(4806)));
    outputs(5109) <= (layer2_outputs(4287)) and not (layer2_outputs(1308));
    outputs(5110) <= layer2_outputs(4476);
    outputs(5111) <= not((layer2_outputs(3680)) xor (layer2_outputs(2559)));
    outputs(5112) <= not(layer2_outputs(4503));
    outputs(5113) <= not(layer2_outputs(3798));
    outputs(5114) <= (layer2_outputs(962)) and (layer2_outputs(3612));
    outputs(5115) <= not(layer2_outputs(3012)) or (layer2_outputs(3422));
    outputs(5116) <= (layer2_outputs(2173)) and (layer2_outputs(4342));
    outputs(5117) <= not(layer2_outputs(3997));
    outputs(5118) <= layer2_outputs(364);
    outputs(5119) <= layer2_outputs(3976);

end Behavioral;
