module logic_network(
    input wire [255:0] inputs,
    output wire [12799:0] outputs
);

    wire [12799:0] layer0_outputs;
    wire [12799:0] layer1_outputs;
    wire [12799:0] layer2_outputs;

    assign layer0_outputs[0] = ~(inputs[220]);
    assign layer0_outputs[1] = ~(inputs[64]);
    assign layer0_outputs[2] = 1'b1;
    assign layer0_outputs[3] = ~(inputs[117]);
    assign layer0_outputs[4] = ~(inputs[25]);
    assign layer0_outputs[5] = inputs[55];
    assign layer0_outputs[6] = ~(inputs[167]);
    assign layer0_outputs[7] = ~((inputs[117]) & (inputs[121]));
    assign layer0_outputs[8] = (inputs[0]) ^ (inputs[107]);
    assign layer0_outputs[9] = ~(inputs[53]);
    assign layer0_outputs[10] = ~(inputs[61]);
    assign layer0_outputs[11] = (inputs[43]) | (inputs[109]);
    assign layer0_outputs[12] = (inputs[210]) ^ (inputs[202]);
    assign layer0_outputs[13] = (inputs[127]) | (inputs[11]);
    assign layer0_outputs[14] = ~(inputs[244]) | (inputs[239]);
    assign layer0_outputs[15] = ~(inputs[65]) | (inputs[145]);
    assign layer0_outputs[16] = (inputs[112]) | (inputs[248]);
    assign layer0_outputs[17] = ~(inputs[245]);
    assign layer0_outputs[18] = ~(inputs[159]);
    assign layer0_outputs[19] = (inputs[145]) | (inputs[7]);
    assign layer0_outputs[20] = ~(inputs[11]) | (inputs[97]);
    assign layer0_outputs[21] = inputs[231];
    assign layer0_outputs[22] = (inputs[47]) | (inputs[77]);
    assign layer0_outputs[23] = inputs[89];
    assign layer0_outputs[24] = (inputs[14]) & (inputs[14]);
    assign layer0_outputs[25] = ~(inputs[173]) | (inputs[48]);
    assign layer0_outputs[26] = (inputs[44]) ^ (inputs[210]);
    assign layer0_outputs[27] = ~((inputs[143]) ^ (inputs[101]));
    assign layer0_outputs[28] = (inputs[245]) | (inputs[205]);
    assign layer0_outputs[29] = (inputs[117]) | (inputs[102]);
    assign layer0_outputs[30] = ~(inputs[115]);
    assign layer0_outputs[31] = (inputs[137]) & ~(inputs[87]);
    assign layer0_outputs[32] = ~((inputs[73]) & (inputs[28]));
    assign layer0_outputs[33] = 1'b0;
    assign layer0_outputs[34] = ~(inputs[76]);
    assign layer0_outputs[35] = ~(inputs[12]) | (inputs[81]);
    assign layer0_outputs[36] = ~((inputs[125]) | (inputs[94]));
    assign layer0_outputs[37] = ~(inputs[219]) | (inputs[21]);
    assign layer0_outputs[38] = ~(inputs[212]) | (inputs[61]);
    assign layer0_outputs[39] = (inputs[49]) ^ (inputs[4]);
    assign layer0_outputs[40] = inputs[196];
    assign layer0_outputs[41] = ~((inputs[145]) ^ (inputs[120]));
    assign layer0_outputs[42] = ~(inputs[120]);
    assign layer0_outputs[43] = ~(inputs[56]) | (inputs[42]);
    assign layer0_outputs[44] = ~((inputs[217]) | (inputs[190]));
    assign layer0_outputs[45] = (inputs[4]) | (inputs[221]);
    assign layer0_outputs[46] = (inputs[200]) & ~(inputs[3]);
    assign layer0_outputs[47] = ~(inputs[120]);
    assign layer0_outputs[48] = (inputs[230]) & ~(inputs[120]);
    assign layer0_outputs[49] = ~(inputs[213]);
    assign layer0_outputs[50] = 1'b0;
    assign layer0_outputs[51] = ~(inputs[213]) | (inputs[54]);
    assign layer0_outputs[52] = ~(inputs[133]) | (inputs[166]);
    assign layer0_outputs[53] = ~(inputs[87]);
    assign layer0_outputs[54] = inputs[151];
    assign layer0_outputs[55] = (inputs[129]) & ~(inputs[80]);
    assign layer0_outputs[56] = (inputs[213]) | (inputs[131]);
    assign layer0_outputs[57] = (inputs[139]) & ~(inputs[70]);
    assign layer0_outputs[58] = 1'b0;
    assign layer0_outputs[59] = ~((inputs[251]) ^ (inputs[107]));
    assign layer0_outputs[60] = (inputs[123]) & ~(inputs[180]);
    assign layer0_outputs[61] = ~((inputs[213]) & (inputs[151]));
    assign layer0_outputs[62] = ~((inputs[103]) | (inputs[22]));
    assign layer0_outputs[63] = ~(inputs[132]) | (inputs[231]);
    assign layer0_outputs[64] = (inputs[252]) ^ (inputs[28]);
    assign layer0_outputs[65] = ~((inputs[94]) ^ (inputs[181]));
    assign layer0_outputs[66] = inputs[34];
    assign layer0_outputs[67] = ~(inputs[94]);
    assign layer0_outputs[68] = 1'b0;
    assign layer0_outputs[69] = inputs[133];
    assign layer0_outputs[70] = ~(inputs[170]) | (inputs[66]);
    assign layer0_outputs[71] = (inputs[10]) & ~(inputs[169]);
    assign layer0_outputs[72] = (inputs[66]) ^ (inputs[49]);
    assign layer0_outputs[73] = ~(inputs[35]);
    assign layer0_outputs[74] = ~(inputs[209]);
    assign layer0_outputs[75] = ~(inputs[100]) | (inputs[9]);
    assign layer0_outputs[76] = (inputs[175]) ^ (inputs[126]);
    assign layer0_outputs[77] = (inputs[213]) | (inputs[195]);
    assign layer0_outputs[78] = inputs[6];
    assign layer0_outputs[79] = ~(inputs[161]);
    assign layer0_outputs[80] = ~(inputs[208]);
    assign layer0_outputs[81] = inputs[71];
    assign layer0_outputs[82] = inputs[109];
    assign layer0_outputs[83] = (inputs[8]) & (inputs[9]);
    assign layer0_outputs[84] = (inputs[159]) ^ (inputs[169]);
    assign layer0_outputs[85] = inputs[176];
    assign layer0_outputs[86] = ~((inputs[173]) ^ (inputs[63]));
    assign layer0_outputs[87] = ~(inputs[227]) | (inputs[154]);
    assign layer0_outputs[88] = ~((inputs[170]) | (inputs[69]));
    assign layer0_outputs[89] = ~(inputs[39]);
    assign layer0_outputs[90] = 1'b1;
    assign layer0_outputs[91] = inputs[161];
    assign layer0_outputs[92] = (inputs[71]) ^ (inputs[23]);
    assign layer0_outputs[93] = ~(inputs[17]) | (inputs[151]);
    assign layer0_outputs[94] = ~(inputs[103]);
    assign layer0_outputs[95] = inputs[2];
    assign layer0_outputs[96] = 1'b1;
    assign layer0_outputs[97] = ~(inputs[76]);
    assign layer0_outputs[98] = ~((inputs[178]) | (inputs[118]));
    assign layer0_outputs[99] = (inputs[87]) & (inputs[95]);
    assign layer0_outputs[100] = inputs[212];
    assign layer0_outputs[101] = 1'b1;
    assign layer0_outputs[102] = ~(inputs[236]) | (inputs[93]);
    assign layer0_outputs[103] = ~(inputs[233]);
    assign layer0_outputs[104] = ~((inputs[21]) ^ (inputs[64]));
    assign layer0_outputs[105] = ~(inputs[90]);
    assign layer0_outputs[106] = (inputs[218]) | (inputs[131]);
    assign layer0_outputs[107] = ~((inputs[48]) | (inputs[180]));
    assign layer0_outputs[108] = (inputs[128]) & ~(inputs[248]);
    assign layer0_outputs[109] = inputs[131];
    assign layer0_outputs[110] = (inputs[133]) | (inputs[213]);
    assign layer0_outputs[111] = 1'b0;
    assign layer0_outputs[112] = ~((inputs[40]) ^ (inputs[255]));
    assign layer0_outputs[113] = ~(inputs[228]);
    assign layer0_outputs[114] = ~(inputs[182]);
    assign layer0_outputs[115] = (inputs[205]) & ~(inputs[249]);
    assign layer0_outputs[116] = (inputs[178]) & ~(inputs[67]);
    assign layer0_outputs[117] = inputs[212];
    assign layer0_outputs[118] = inputs[229];
    assign layer0_outputs[119] = ~(inputs[90]) | (inputs[160]);
    assign layer0_outputs[120] = ~(inputs[35]) | (inputs[25]);
    assign layer0_outputs[121] = 1'b1;
    assign layer0_outputs[122] = (inputs[118]) & ~(inputs[15]);
    assign layer0_outputs[123] = ~((inputs[32]) | (inputs[167]));
    assign layer0_outputs[124] = ~(inputs[50]) | (inputs[202]);
    assign layer0_outputs[125] = 1'b0;
    assign layer0_outputs[126] = ~(inputs[227]) | (inputs[108]);
    assign layer0_outputs[127] = (inputs[52]) & ~(inputs[182]);
    assign layer0_outputs[128] = (inputs[125]) | (inputs[144]);
    assign layer0_outputs[129] = inputs[190];
    assign layer0_outputs[130] = inputs[9];
    assign layer0_outputs[131] = ~((inputs[245]) | (inputs[10]));
    assign layer0_outputs[132] = (inputs[41]) | (inputs[96]);
    assign layer0_outputs[133] = (inputs[56]) & ~(inputs[112]);
    assign layer0_outputs[134] = 1'b0;
    assign layer0_outputs[135] = (inputs[245]) & ~(inputs[218]);
    assign layer0_outputs[136] = inputs[162];
    assign layer0_outputs[137] = (inputs[216]) & ~(inputs[199]);
    assign layer0_outputs[138] = ~(inputs[26]);
    assign layer0_outputs[139] = (inputs[83]) ^ (inputs[134]);
    assign layer0_outputs[140] = 1'b0;
    assign layer0_outputs[141] = (inputs[51]) | (inputs[91]);
    assign layer0_outputs[142] = inputs[76];
    assign layer0_outputs[143] = ~(inputs[57]);
    assign layer0_outputs[144] = ~(inputs[180]);
    assign layer0_outputs[145] = ~((inputs[143]) | (inputs[142]));
    assign layer0_outputs[146] = ~((inputs[91]) | (inputs[171]));
    assign layer0_outputs[147] = ~(inputs[108]);
    assign layer0_outputs[148] = ~(inputs[10]) | (inputs[211]);
    assign layer0_outputs[149] = ~(inputs[85]);
    assign layer0_outputs[150] = ~((inputs[138]) & (inputs[98]));
    assign layer0_outputs[151] = inputs[109];
    assign layer0_outputs[152] = ~(inputs[237]);
    assign layer0_outputs[153] = inputs[205];
    assign layer0_outputs[154] = inputs[55];
    assign layer0_outputs[155] = inputs[106];
    assign layer0_outputs[156] = inputs[25];
    assign layer0_outputs[157] = (inputs[11]) & (inputs[217]);
    assign layer0_outputs[158] = inputs[179];
    assign layer0_outputs[159] = inputs[73];
    assign layer0_outputs[160] = (inputs[44]) & ~(inputs[115]);
    assign layer0_outputs[161] = ~((inputs[131]) & (inputs[60]));
    assign layer0_outputs[162] = (inputs[1]) & (inputs[125]);
    assign layer0_outputs[163] = (inputs[186]) & (inputs[230]);
    assign layer0_outputs[164] = (inputs[239]) & ~(inputs[21]);
    assign layer0_outputs[165] = (inputs[115]) ^ (inputs[7]);
    assign layer0_outputs[166] = (inputs[102]) ^ (inputs[64]);
    assign layer0_outputs[167] = inputs[25];
    assign layer0_outputs[168] = ~(inputs[206]);
    assign layer0_outputs[169] = ~(inputs[84]) | (inputs[175]);
    assign layer0_outputs[170] = (inputs[229]) ^ (inputs[159]);
    assign layer0_outputs[171] = inputs[146];
    assign layer0_outputs[172] = ~((inputs[100]) ^ (inputs[98]));
    assign layer0_outputs[173] = (inputs[83]) & ~(inputs[254]);
    assign layer0_outputs[174] = ~(inputs[166]);
    assign layer0_outputs[175] = ~((inputs[166]) ^ (inputs[95]));
    assign layer0_outputs[176] = ~((inputs[34]) ^ (inputs[203]));
    assign layer0_outputs[177] = (inputs[145]) | (inputs[113]);
    assign layer0_outputs[178] = ~(inputs[152]);
    assign layer0_outputs[179] = ~((inputs[195]) | (inputs[254]));
    assign layer0_outputs[180] = ~(inputs[206]);
    assign layer0_outputs[181] = ~(inputs[148]) | (inputs[253]);
    assign layer0_outputs[182] = (inputs[151]) ^ (inputs[110]);
    assign layer0_outputs[183] = (inputs[113]) | (inputs[3]);
    assign layer0_outputs[184] = inputs[194];
    assign layer0_outputs[185] = ~(inputs[20]) | (inputs[108]);
    assign layer0_outputs[186] = ~(inputs[91]);
    assign layer0_outputs[187] = (inputs[90]) | (inputs[175]);
    assign layer0_outputs[188] = ~((inputs[111]) | (inputs[26]));
    assign layer0_outputs[189] = ~((inputs[145]) & (inputs[43]));
    assign layer0_outputs[190] = inputs[150];
    assign layer0_outputs[191] = (inputs[193]) & ~(inputs[209]);
    assign layer0_outputs[192] = inputs[142];
    assign layer0_outputs[193] = inputs[112];
    assign layer0_outputs[194] = ~(inputs[22]);
    assign layer0_outputs[195] = (inputs[104]) & ~(inputs[145]);
    assign layer0_outputs[196] = ~(inputs[152]);
    assign layer0_outputs[197] = ~((inputs[196]) | (inputs[209]));
    assign layer0_outputs[198] = (inputs[238]) ^ (inputs[189]);
    assign layer0_outputs[199] = ~(inputs[183]) | (inputs[40]);
    assign layer0_outputs[200] = ~((inputs[64]) ^ (inputs[197]));
    assign layer0_outputs[201] = ~((inputs[178]) & (inputs[57]));
    assign layer0_outputs[202] = ~((inputs[20]) ^ (inputs[14]));
    assign layer0_outputs[203] = ~(inputs[166]);
    assign layer0_outputs[204] = (inputs[64]) & ~(inputs[253]);
    assign layer0_outputs[205] = ~((inputs[228]) | (inputs[62]));
    assign layer0_outputs[206] = (inputs[214]) ^ (inputs[174]);
    assign layer0_outputs[207] = (inputs[15]) & ~(inputs[9]);
    assign layer0_outputs[208] = inputs[99];
    assign layer0_outputs[209] = inputs[136];
    assign layer0_outputs[210] = inputs[157];
    assign layer0_outputs[211] = inputs[225];
    assign layer0_outputs[212] = ~(inputs[199]);
    assign layer0_outputs[213] = ~(inputs[157]);
    assign layer0_outputs[214] = (inputs[253]) & ~(inputs[113]);
    assign layer0_outputs[215] = inputs[151];
    assign layer0_outputs[216] = 1'b1;
    assign layer0_outputs[217] = ~((inputs[84]) | (inputs[186]));
    assign layer0_outputs[218] = ~(inputs[235]);
    assign layer0_outputs[219] = ~((inputs[204]) | (inputs[249]));
    assign layer0_outputs[220] = ~(inputs[82]);
    assign layer0_outputs[221] = ~((inputs[86]) ^ (inputs[66]));
    assign layer0_outputs[222] = ~((inputs[247]) | (inputs[192]));
    assign layer0_outputs[223] = inputs[229];
    assign layer0_outputs[224] = ~(inputs[155]);
    assign layer0_outputs[225] = (inputs[10]) ^ (inputs[4]);
    assign layer0_outputs[226] = ~(inputs[9]) | (inputs[16]);
    assign layer0_outputs[227] = ~(inputs[162]) | (inputs[150]);
    assign layer0_outputs[228] = ~((inputs[35]) ^ (inputs[105]));
    assign layer0_outputs[229] = ~((inputs[161]) ^ (inputs[165]));
    assign layer0_outputs[230] = ~((inputs[249]) | (inputs[253]));
    assign layer0_outputs[231] = (inputs[163]) | (inputs[206]);
    assign layer0_outputs[232] = inputs[205];
    assign layer0_outputs[233] = ~(inputs[115]);
    assign layer0_outputs[234] = (inputs[144]) ^ (inputs[40]);
    assign layer0_outputs[235] = (inputs[13]) & ~(inputs[130]);
    assign layer0_outputs[236] = ~((inputs[224]) | (inputs[161]));
    assign layer0_outputs[237] = (inputs[29]) | (inputs[213]);
    assign layer0_outputs[238] = ~((inputs[156]) | (inputs[236]));
    assign layer0_outputs[239] = (inputs[104]) & ~(inputs[213]);
    assign layer0_outputs[240] = ~(inputs[75]);
    assign layer0_outputs[241] = ~(inputs[100]);
    assign layer0_outputs[242] = ~(inputs[41]);
    assign layer0_outputs[243] = (inputs[93]) | (inputs[26]);
    assign layer0_outputs[244] = ~((inputs[248]) & (inputs[129]));
    assign layer0_outputs[245] = inputs[194];
    assign layer0_outputs[246] = ~(inputs[70]);
    assign layer0_outputs[247] = ~((inputs[209]) ^ (inputs[108]));
    assign layer0_outputs[248] = ~((inputs[117]) ^ (inputs[69]));
    assign layer0_outputs[249] = ~(inputs[183]) | (inputs[46]);
    assign layer0_outputs[250] = inputs[136];
    assign layer0_outputs[251] = ~((inputs[158]) ^ (inputs[108]));
    assign layer0_outputs[252] = (inputs[17]) ^ (inputs[32]);
    assign layer0_outputs[253] = ~((inputs[25]) ^ (inputs[176]));
    assign layer0_outputs[254] = ~(inputs[221]);
    assign layer0_outputs[255] = (inputs[202]) & ~(inputs[163]);
    assign layer0_outputs[256] = (inputs[37]) | (inputs[46]);
    assign layer0_outputs[257] = ~((inputs[114]) | (inputs[83]));
    assign layer0_outputs[258] = (inputs[122]) ^ (inputs[174]);
    assign layer0_outputs[259] = 1'b1;
    assign layer0_outputs[260] = (inputs[199]) & ~(inputs[96]);
    assign layer0_outputs[261] = ~((inputs[102]) & (inputs[193]));
    assign layer0_outputs[262] = ~(inputs[161]) | (inputs[192]);
    assign layer0_outputs[263] = (inputs[220]) | (inputs[223]);
    assign layer0_outputs[264] = inputs[21];
    assign layer0_outputs[265] = (inputs[88]) & ~(inputs[255]);
    assign layer0_outputs[266] = (inputs[84]) & ~(inputs[72]);
    assign layer0_outputs[267] = (inputs[229]) ^ (inputs[19]);
    assign layer0_outputs[268] = ~((inputs[207]) | (inputs[119]));
    assign layer0_outputs[269] = inputs[178];
    assign layer0_outputs[270] = (inputs[22]) | (inputs[61]);
    assign layer0_outputs[271] = ~(inputs[77]);
    assign layer0_outputs[272] = ~((inputs[136]) ^ (inputs[103]));
    assign layer0_outputs[273] = inputs[230];
    assign layer0_outputs[274] = (inputs[197]) & ~(inputs[4]);
    assign layer0_outputs[275] = ~(inputs[136]);
    assign layer0_outputs[276] = ~(inputs[76]);
    assign layer0_outputs[277] = ~((inputs[100]) & (inputs[106]));
    assign layer0_outputs[278] = ~(inputs[45]);
    assign layer0_outputs[279] = inputs[145];
    assign layer0_outputs[280] = inputs[164];
    assign layer0_outputs[281] = ~((inputs[98]) ^ (inputs[154]));
    assign layer0_outputs[282] = ~(inputs[79]) | (inputs[172]);
    assign layer0_outputs[283] = ~(inputs[137]);
    assign layer0_outputs[284] = ~((inputs[141]) ^ (inputs[46]));
    assign layer0_outputs[285] = inputs[22];
    assign layer0_outputs[286] = ~(inputs[162]);
    assign layer0_outputs[287] = (inputs[23]) & ~(inputs[29]);
    assign layer0_outputs[288] = ~(inputs[249]) | (inputs[64]);
    assign layer0_outputs[289] = (inputs[8]) | (inputs[239]);
    assign layer0_outputs[290] = inputs[165];
    assign layer0_outputs[291] = ~((inputs[98]) | (inputs[126]));
    assign layer0_outputs[292] = ~(inputs[42]) | (inputs[184]);
    assign layer0_outputs[293] = ~(inputs[81]);
    assign layer0_outputs[294] = ~(inputs[137]);
    assign layer0_outputs[295] = 1'b0;
    assign layer0_outputs[296] = ~(inputs[72]) | (inputs[5]);
    assign layer0_outputs[297] = 1'b0;
    assign layer0_outputs[298] = inputs[170];
    assign layer0_outputs[299] = ~((inputs[63]) ^ (inputs[42]));
    assign layer0_outputs[300] = ~(inputs[99]) | (inputs[235]);
    assign layer0_outputs[301] = (inputs[56]) | (inputs[13]);
    assign layer0_outputs[302] = inputs[29];
    assign layer0_outputs[303] = (inputs[137]) ^ (inputs[131]);
    assign layer0_outputs[304] = inputs[137];
    assign layer0_outputs[305] = (inputs[174]) | (inputs[75]);
    assign layer0_outputs[306] = ~((inputs[197]) | (inputs[128]));
    assign layer0_outputs[307] = (inputs[26]) | (inputs[3]);
    assign layer0_outputs[308] = ~((inputs[4]) & (inputs[67]));
    assign layer0_outputs[309] = ~(inputs[147]);
    assign layer0_outputs[310] = ~((inputs[185]) & (inputs[141]));
    assign layer0_outputs[311] = ~(inputs[97]);
    assign layer0_outputs[312] = ~((inputs[240]) & (inputs[184]));
    assign layer0_outputs[313] = ~(inputs[143]);
    assign layer0_outputs[314] = ~(inputs[184]);
    assign layer0_outputs[315] = ~((inputs[59]) | (inputs[15]));
    assign layer0_outputs[316] = inputs[236];
    assign layer0_outputs[317] = ~(inputs[151]) | (inputs[63]);
    assign layer0_outputs[318] = (inputs[150]) & ~(inputs[12]);
    assign layer0_outputs[319] = ~((inputs[208]) | (inputs[31]));
    assign layer0_outputs[320] = 1'b1;
    assign layer0_outputs[321] = inputs[253];
    assign layer0_outputs[322] = ~((inputs[145]) ^ (inputs[238]));
    assign layer0_outputs[323] = inputs[15];
    assign layer0_outputs[324] = ~((inputs[86]) & (inputs[31]));
    assign layer0_outputs[325] = (inputs[90]) & ~(inputs[176]);
    assign layer0_outputs[326] = inputs[100];
    assign layer0_outputs[327] = (inputs[119]) | (inputs[174]);
    assign layer0_outputs[328] = (inputs[112]) | (inputs[132]);
    assign layer0_outputs[329] = ~(inputs[173]) | (inputs[22]);
    assign layer0_outputs[330] = inputs[63];
    assign layer0_outputs[331] = (inputs[194]) | (inputs[237]);
    assign layer0_outputs[332] = ~(inputs[158]) | (inputs[81]);
    assign layer0_outputs[333] = ~(inputs[38]);
    assign layer0_outputs[334] = (inputs[139]) | (inputs[43]);
    assign layer0_outputs[335] = ~((inputs[45]) | (inputs[238]));
    assign layer0_outputs[336] = ~(inputs[215]);
    assign layer0_outputs[337] = (inputs[172]) & (inputs[233]);
    assign layer0_outputs[338] = (inputs[104]) & ~(inputs[197]);
    assign layer0_outputs[339] = ~((inputs[188]) | (inputs[16]));
    assign layer0_outputs[340] = (inputs[215]) & ~(inputs[131]);
    assign layer0_outputs[341] = ~(inputs[42]) | (inputs[204]);
    assign layer0_outputs[342] = (inputs[161]) & ~(inputs[67]);
    assign layer0_outputs[343] = ~((inputs[60]) & (inputs[81]));
    assign layer0_outputs[344] = 1'b1;
    assign layer0_outputs[345] = inputs[13];
    assign layer0_outputs[346] = ~(inputs[254]) | (inputs[166]);
    assign layer0_outputs[347] = (inputs[65]) ^ (inputs[90]);
    assign layer0_outputs[348] = (inputs[140]) | (inputs[73]);
    assign layer0_outputs[349] = ~(inputs[41]);
    assign layer0_outputs[350] = ~(inputs[196]) | (inputs[34]);
    assign layer0_outputs[351] = ~((inputs[110]) | (inputs[240]));
    assign layer0_outputs[352] = ~(inputs[22]) | (inputs[152]);
    assign layer0_outputs[353] = ~((inputs[54]) ^ (inputs[37]));
    assign layer0_outputs[354] = ~(inputs[248]);
    assign layer0_outputs[355] = ~(inputs[109]);
    assign layer0_outputs[356] = ~(inputs[103]) | (inputs[127]);
    assign layer0_outputs[357] = (inputs[30]) & ~(inputs[79]);
    assign layer0_outputs[358] = inputs[155];
    assign layer0_outputs[359] = ~((inputs[75]) | (inputs[200]));
    assign layer0_outputs[360] = ~(inputs[102]) | (inputs[1]);
    assign layer0_outputs[361] = inputs[137];
    assign layer0_outputs[362] = (inputs[84]) ^ (inputs[81]);
    assign layer0_outputs[363] = inputs[98];
    assign layer0_outputs[364] = (inputs[21]) ^ (inputs[93]);
    assign layer0_outputs[365] = ~((inputs[186]) & (inputs[58]));
    assign layer0_outputs[366] = ~(inputs[88]) | (inputs[191]);
    assign layer0_outputs[367] = inputs[85];
    assign layer0_outputs[368] = (inputs[206]) & ~(inputs[13]);
    assign layer0_outputs[369] = (inputs[146]) & (inputs[219]);
    assign layer0_outputs[370] = ~(inputs[229]);
    assign layer0_outputs[371] = 1'b1;
    assign layer0_outputs[372] = ~(inputs[104]);
    assign layer0_outputs[373] = inputs[90];
    assign layer0_outputs[374] = ~(inputs[115]);
    assign layer0_outputs[375] = (inputs[20]) & (inputs[206]);
    assign layer0_outputs[376] = (inputs[237]) ^ (inputs[206]);
    assign layer0_outputs[377] = inputs[6];
    assign layer0_outputs[378] = (inputs[51]) | (inputs[255]);
    assign layer0_outputs[379] = (inputs[35]) ^ (inputs[72]);
    assign layer0_outputs[380] = ~(inputs[93]);
    assign layer0_outputs[381] = ~(inputs[11]) | (inputs[28]);
    assign layer0_outputs[382] = (inputs[194]) & ~(inputs[0]);
    assign layer0_outputs[383] = ~(inputs[110]) | (inputs[95]);
    assign layer0_outputs[384] = (inputs[236]) | (inputs[103]);
    assign layer0_outputs[385] = (inputs[49]) | (inputs[25]);
    assign layer0_outputs[386] = ~(inputs[6]);
    assign layer0_outputs[387] = ~(inputs[78]);
    assign layer0_outputs[388] = inputs[94];
    assign layer0_outputs[389] = (inputs[197]) & (inputs[255]);
    assign layer0_outputs[390] = (inputs[39]) ^ (inputs[120]);
    assign layer0_outputs[391] = ~((inputs[98]) ^ (inputs[68]));
    assign layer0_outputs[392] = ~(inputs[228]) | (inputs[254]);
    assign layer0_outputs[393] = ~(inputs[94]);
    assign layer0_outputs[394] = (inputs[223]) ^ (inputs[191]);
    assign layer0_outputs[395] = inputs[133];
    assign layer0_outputs[396] = ~((inputs[244]) ^ (inputs[106]));
    assign layer0_outputs[397] = ~(inputs[230]) | (inputs[54]);
    assign layer0_outputs[398] = ~((inputs[114]) | (inputs[30]));
    assign layer0_outputs[399] = inputs[229];
    assign layer0_outputs[400] = (inputs[164]) & (inputs[125]);
    assign layer0_outputs[401] = ~(inputs[146]);
    assign layer0_outputs[402] = inputs[43];
    assign layer0_outputs[403] = ~(inputs[185]);
    assign layer0_outputs[404] = ~((inputs[208]) | (inputs[154]));
    assign layer0_outputs[405] = ~((inputs[22]) | (inputs[236]));
    assign layer0_outputs[406] = (inputs[92]) & ~(inputs[255]);
    assign layer0_outputs[407] = ~(inputs[74]);
    assign layer0_outputs[408] = ~(inputs[232]);
    assign layer0_outputs[409] = ~(inputs[234]);
    assign layer0_outputs[410] = ~(inputs[169]);
    assign layer0_outputs[411] = (inputs[48]) & ~(inputs[179]);
    assign layer0_outputs[412] = (inputs[38]) & (inputs[229]);
    assign layer0_outputs[413] = (inputs[108]) ^ (inputs[4]);
    assign layer0_outputs[414] = ~(inputs[172]) | (inputs[133]);
    assign layer0_outputs[415] = (inputs[242]) | (inputs[212]);
    assign layer0_outputs[416] = (inputs[3]) & ~(inputs[141]);
    assign layer0_outputs[417] = ~((inputs[123]) ^ (inputs[132]));
    assign layer0_outputs[418] = (inputs[88]) & ~(inputs[208]);
    assign layer0_outputs[419] = ~(inputs[160]);
    assign layer0_outputs[420] = 1'b0;
    assign layer0_outputs[421] = ~((inputs[32]) | (inputs[231]));
    assign layer0_outputs[422] = inputs[105];
    assign layer0_outputs[423] = (inputs[63]) | (inputs[45]);
    assign layer0_outputs[424] = ~(inputs[218]);
    assign layer0_outputs[425] = (inputs[52]) & ~(inputs[4]);
    assign layer0_outputs[426] = (inputs[140]) ^ (inputs[175]);
    assign layer0_outputs[427] = ~((inputs[100]) ^ (inputs[3]));
    assign layer0_outputs[428] = (inputs[142]) | (inputs[29]);
    assign layer0_outputs[429] = inputs[214];
    assign layer0_outputs[430] = ~(inputs[83]) | (inputs[252]);
    assign layer0_outputs[431] = (inputs[95]) ^ (inputs[57]);
    assign layer0_outputs[432] = (inputs[34]) ^ (inputs[97]);
    assign layer0_outputs[433] = (inputs[88]) | (inputs[106]);
    assign layer0_outputs[434] = (inputs[111]) ^ (inputs[45]);
    assign layer0_outputs[435] = (inputs[55]) | (inputs[175]);
    assign layer0_outputs[436] = ~(inputs[57]);
    assign layer0_outputs[437] = (inputs[219]) & ~(inputs[94]);
    assign layer0_outputs[438] = (inputs[63]) & ~(inputs[227]);
    assign layer0_outputs[439] = (inputs[29]) & ~(inputs[70]);
    assign layer0_outputs[440] = ~(inputs[165]);
    assign layer0_outputs[441] = ~(inputs[119]);
    assign layer0_outputs[442] = (inputs[156]) & ~(inputs[126]);
    assign layer0_outputs[443] = ~((inputs[79]) | (inputs[104]));
    assign layer0_outputs[444] = (inputs[237]) & (inputs[67]);
    assign layer0_outputs[445] = ~((inputs[253]) ^ (inputs[87]));
    assign layer0_outputs[446] = inputs[111];
    assign layer0_outputs[447] = inputs[182];
    assign layer0_outputs[448] = (inputs[151]) ^ (inputs[33]);
    assign layer0_outputs[449] = ~((inputs[237]) | (inputs[87]));
    assign layer0_outputs[450] = ~((inputs[144]) ^ (inputs[201]));
    assign layer0_outputs[451] = (inputs[121]) & ~(inputs[48]);
    assign layer0_outputs[452] = (inputs[21]) & (inputs[102]);
    assign layer0_outputs[453] = 1'b1;
    assign layer0_outputs[454] = ~((inputs[42]) & (inputs[240]));
    assign layer0_outputs[455] = (inputs[216]) & ~(inputs[56]);
    assign layer0_outputs[456] = ~((inputs[43]) & (inputs[29]));
    assign layer0_outputs[457] = (inputs[123]) | (inputs[227]);
    assign layer0_outputs[458] = (inputs[199]) | (inputs[60]);
    assign layer0_outputs[459] = ~(inputs[102]);
    assign layer0_outputs[460] = ~((inputs[122]) & (inputs[43]));
    assign layer0_outputs[461] = 1'b1;
    assign layer0_outputs[462] = ~(inputs[188]);
    assign layer0_outputs[463] = ~(inputs[61]);
    assign layer0_outputs[464] = ~(inputs[37]);
    assign layer0_outputs[465] = ~(inputs[129]);
    assign layer0_outputs[466] = (inputs[71]) | (inputs[148]);
    assign layer0_outputs[467] = (inputs[74]) & ~(inputs[254]);
    assign layer0_outputs[468] = (inputs[9]) & ~(inputs[208]);
    assign layer0_outputs[469] = ~(inputs[26]) | (inputs[181]);
    assign layer0_outputs[470] = (inputs[64]) & (inputs[77]);
    assign layer0_outputs[471] = (inputs[72]) ^ (inputs[179]);
    assign layer0_outputs[472] = ~((inputs[89]) ^ (inputs[28]));
    assign layer0_outputs[473] = ~(inputs[250]);
    assign layer0_outputs[474] = ~(inputs[171]) | (inputs[35]);
    assign layer0_outputs[475] = 1'b0;
    assign layer0_outputs[476] = ~(inputs[27]);
    assign layer0_outputs[477] = ~(inputs[134]) | (inputs[31]);
    assign layer0_outputs[478] = (inputs[3]) & (inputs[210]);
    assign layer0_outputs[479] = (inputs[167]) | (inputs[110]);
    assign layer0_outputs[480] = ~(inputs[15]);
    assign layer0_outputs[481] = ~((inputs[179]) ^ (inputs[174]));
    assign layer0_outputs[482] = (inputs[7]) & ~(inputs[44]);
    assign layer0_outputs[483] = ~((inputs[225]) | (inputs[201]));
    assign layer0_outputs[484] = 1'b1;
    assign layer0_outputs[485] = ~((inputs[52]) | (inputs[111]));
    assign layer0_outputs[486] = (inputs[36]) ^ (inputs[71]);
    assign layer0_outputs[487] = (inputs[223]) | (inputs[82]);
    assign layer0_outputs[488] = (inputs[38]) & ~(inputs[153]);
    assign layer0_outputs[489] = ~(inputs[94]);
    assign layer0_outputs[490] = (inputs[3]) ^ (inputs[99]);
    assign layer0_outputs[491] = ~((inputs[158]) | (inputs[183]));
    assign layer0_outputs[492] = ~((inputs[36]) | (inputs[76]));
    assign layer0_outputs[493] = ~((inputs[157]) | (inputs[173]));
    assign layer0_outputs[494] = (inputs[160]) & ~(inputs[14]);
    assign layer0_outputs[495] = ~((inputs[174]) | (inputs[132]));
    assign layer0_outputs[496] = ~(inputs[229]);
    assign layer0_outputs[497] = inputs[251];
    assign layer0_outputs[498] = (inputs[237]) | (inputs[186]);
    assign layer0_outputs[499] = (inputs[130]) & ~(inputs[121]);
    assign layer0_outputs[500] = (inputs[135]) & ~(inputs[231]);
    assign layer0_outputs[501] = ~(inputs[134]);
    assign layer0_outputs[502] = inputs[249];
    assign layer0_outputs[503] = ~((inputs[192]) | (inputs[77]));
    assign layer0_outputs[504] = (inputs[7]) | (inputs[219]);
    assign layer0_outputs[505] = (inputs[67]) ^ (inputs[204]);
    assign layer0_outputs[506] = inputs[63];
    assign layer0_outputs[507] = (inputs[119]) & ~(inputs[241]);
    assign layer0_outputs[508] = ~(inputs[83]) | (inputs[24]);
    assign layer0_outputs[509] = 1'b1;
    assign layer0_outputs[510] = ~((inputs[190]) | (inputs[181]));
    assign layer0_outputs[511] = ~(inputs[40]) | (inputs[185]);
    assign layer0_outputs[512] = ~(inputs[202]);
    assign layer0_outputs[513] = ~((inputs[240]) ^ (inputs[156]));
    assign layer0_outputs[514] = ~(inputs[16]);
    assign layer0_outputs[515] = (inputs[67]) | (inputs[82]);
    assign layer0_outputs[516] = ~((inputs[54]) ^ (inputs[105]));
    assign layer0_outputs[517] = ~(inputs[56]) | (inputs[241]);
    assign layer0_outputs[518] = 1'b0;
    assign layer0_outputs[519] = ~((inputs[177]) ^ (inputs[209]));
    assign layer0_outputs[520] = (inputs[202]) & ~(inputs[175]);
    assign layer0_outputs[521] = ~((inputs[214]) & (inputs[222]));
    assign layer0_outputs[522] = ~(inputs[170]);
    assign layer0_outputs[523] = inputs[87];
    assign layer0_outputs[524] = ~((inputs[21]) ^ (inputs[255]));
    assign layer0_outputs[525] = ~((inputs[12]) ^ (inputs[171]));
    assign layer0_outputs[526] = ~((inputs[168]) | (inputs[210]));
    assign layer0_outputs[527] = ~(inputs[158]);
    assign layer0_outputs[528] = inputs[162];
    assign layer0_outputs[529] = (inputs[153]) & ~(inputs[54]);
    assign layer0_outputs[530] = (inputs[133]) | (inputs[84]);
    assign layer0_outputs[531] = ~(inputs[20]) | (inputs[232]);
    assign layer0_outputs[532] = ~(inputs[204]) | (inputs[30]);
    assign layer0_outputs[533] = ~((inputs[169]) & (inputs[163]));
    assign layer0_outputs[534] = 1'b1;
    assign layer0_outputs[535] = ~(inputs[82]);
    assign layer0_outputs[536] = ~(inputs[255]) | (inputs[59]);
    assign layer0_outputs[537] = 1'b0;
    assign layer0_outputs[538] = ~(inputs[71]) | (inputs[16]);
    assign layer0_outputs[539] = ~(inputs[148]) | (inputs[26]);
    assign layer0_outputs[540] = (inputs[247]) & ~(inputs[77]);
    assign layer0_outputs[541] = (inputs[242]) | (inputs[210]);
    assign layer0_outputs[542] = inputs[107];
    assign layer0_outputs[543] = ~((inputs[129]) ^ (inputs[138]));
    assign layer0_outputs[544] = (inputs[50]) & ~(inputs[45]);
    assign layer0_outputs[545] = (inputs[251]) | (inputs[212]);
    assign layer0_outputs[546] = (inputs[241]) | (inputs[135]);
    assign layer0_outputs[547] = ~((inputs[51]) | (inputs[118]));
    assign layer0_outputs[548] = inputs[166];
    assign layer0_outputs[549] = ~(inputs[105]);
    assign layer0_outputs[550] = ~((inputs[171]) & (inputs[200]));
    assign layer0_outputs[551] = ~(inputs[78]);
    assign layer0_outputs[552] = (inputs[189]) ^ (inputs[110]);
    assign layer0_outputs[553] = ~(inputs[253]);
    assign layer0_outputs[554] = (inputs[218]) ^ (inputs[124]);
    assign layer0_outputs[555] = ~(inputs[172]);
    assign layer0_outputs[556] = (inputs[22]) | (inputs[213]);
    assign layer0_outputs[557] = ~((inputs[31]) & (inputs[233]));
    assign layer0_outputs[558] = ~(inputs[113]);
    assign layer0_outputs[559] = inputs[100];
    assign layer0_outputs[560] = ~((inputs[0]) | (inputs[149]));
    assign layer0_outputs[561] = (inputs[226]) | (inputs[65]);
    assign layer0_outputs[562] = ~(inputs[25]);
    assign layer0_outputs[563] = ~(inputs[100]) | (inputs[164]);
    assign layer0_outputs[564] = inputs[215];
    assign layer0_outputs[565] = (inputs[115]) & ~(inputs[58]);
    assign layer0_outputs[566] = (inputs[86]) ^ (inputs[229]);
    assign layer0_outputs[567] = ~(inputs[10]);
    assign layer0_outputs[568] = ~((inputs[88]) & (inputs[54]));
    assign layer0_outputs[569] = ~((inputs[73]) ^ (inputs[95]));
    assign layer0_outputs[570] = ~((inputs[212]) | (inputs[223]));
    assign layer0_outputs[571] = (inputs[102]) & ~(inputs[88]);
    assign layer0_outputs[572] = (inputs[88]) | (inputs[48]);
    assign layer0_outputs[573] = (inputs[223]) | (inputs[218]);
    assign layer0_outputs[574] = ~(inputs[191]);
    assign layer0_outputs[575] = ~(inputs[127]);
    assign layer0_outputs[576] = ~(inputs[145]);
    assign layer0_outputs[577] = ~((inputs[72]) ^ (inputs[179]));
    assign layer0_outputs[578] = (inputs[120]) | (inputs[44]);
    assign layer0_outputs[579] = ~((inputs[67]) ^ (inputs[24]));
    assign layer0_outputs[580] = ~((inputs[203]) ^ (inputs[157]));
    assign layer0_outputs[581] = inputs[114];
    assign layer0_outputs[582] = ~((inputs[176]) | (inputs[206]));
    assign layer0_outputs[583] = (inputs[18]) ^ (inputs[238]);
    assign layer0_outputs[584] = ~((inputs[147]) | (inputs[180]));
    assign layer0_outputs[585] = ~((inputs[57]) | (inputs[161]));
    assign layer0_outputs[586] = ~(inputs[13]);
    assign layer0_outputs[587] = (inputs[136]) & (inputs[233]);
    assign layer0_outputs[588] = ~(inputs[154]);
    assign layer0_outputs[589] = (inputs[37]) & ~(inputs[143]);
    assign layer0_outputs[590] = ~((inputs[45]) ^ (inputs[251]));
    assign layer0_outputs[591] = ~(inputs[154]);
    assign layer0_outputs[592] = ~((inputs[160]) | (inputs[76]));
    assign layer0_outputs[593] = (inputs[223]) ^ (inputs[108]);
    assign layer0_outputs[594] = (inputs[242]) | (inputs[225]);
    assign layer0_outputs[595] = inputs[221];
    assign layer0_outputs[596] = (inputs[253]) & ~(inputs[51]);
    assign layer0_outputs[597] = (inputs[51]) & ~(inputs[165]);
    assign layer0_outputs[598] = ~(inputs[90]) | (inputs[244]);
    assign layer0_outputs[599] = (inputs[246]) & ~(inputs[17]);
    assign layer0_outputs[600] = inputs[60];
    assign layer0_outputs[601] = ~((inputs[212]) | (inputs[76]));
    assign layer0_outputs[602] = ~(inputs[162]);
    assign layer0_outputs[603] = (inputs[36]) | (inputs[12]);
    assign layer0_outputs[604] = ~((inputs[89]) ^ (inputs[91]));
    assign layer0_outputs[605] = (inputs[55]) ^ (inputs[99]);
    assign layer0_outputs[606] = (inputs[105]) & ~(inputs[22]);
    assign layer0_outputs[607] = inputs[102];
    assign layer0_outputs[608] = inputs[109];
    assign layer0_outputs[609] = ~(inputs[72]);
    assign layer0_outputs[610] = ~((inputs[184]) ^ (inputs[178]));
    assign layer0_outputs[611] = 1'b1;
    assign layer0_outputs[612] = ~(inputs[85]);
    assign layer0_outputs[613] = ~(inputs[76]);
    assign layer0_outputs[614] = ~(inputs[247]);
    assign layer0_outputs[615] = ~(inputs[167]) | (inputs[150]);
    assign layer0_outputs[616] = (inputs[68]) ^ (inputs[115]);
    assign layer0_outputs[617] = ~(inputs[114]);
    assign layer0_outputs[618] = ~(inputs[111]) | (inputs[169]);
    assign layer0_outputs[619] = ~((inputs[130]) & (inputs[57]));
    assign layer0_outputs[620] = (inputs[25]) & ~(inputs[126]);
    assign layer0_outputs[621] = (inputs[188]) ^ (inputs[109]);
    assign layer0_outputs[622] = ~(inputs[84]) | (inputs[209]);
    assign layer0_outputs[623] = (inputs[216]) & (inputs[204]);
    assign layer0_outputs[624] = (inputs[99]) | (inputs[45]);
    assign layer0_outputs[625] = ~((inputs[24]) | (inputs[5]));
    assign layer0_outputs[626] = inputs[68];
    assign layer0_outputs[627] = ~(inputs[2]);
    assign layer0_outputs[628] = inputs[13];
    assign layer0_outputs[629] = (inputs[56]) | (inputs[245]);
    assign layer0_outputs[630] = ~((inputs[187]) ^ (inputs[36]));
    assign layer0_outputs[631] = inputs[202];
    assign layer0_outputs[632] = (inputs[103]) & ~(inputs[192]);
    assign layer0_outputs[633] = 1'b1;
    assign layer0_outputs[634] = (inputs[32]) | (inputs[220]);
    assign layer0_outputs[635] = (inputs[58]) ^ (inputs[214]);
    assign layer0_outputs[636] = 1'b1;
    assign layer0_outputs[637] = inputs[5];
    assign layer0_outputs[638] = ~(inputs[18]) | (inputs[221]);
    assign layer0_outputs[639] = ~(inputs[69]) | (inputs[144]);
    assign layer0_outputs[640] = (inputs[225]) & ~(inputs[31]);
    assign layer0_outputs[641] = ~(inputs[38]);
    assign layer0_outputs[642] = (inputs[208]) & ~(inputs[77]);
    assign layer0_outputs[643] = 1'b0;
    assign layer0_outputs[644] = 1'b1;
    assign layer0_outputs[645] = ~(inputs[118]) | (inputs[137]);
    assign layer0_outputs[646] = ~(inputs[81]);
    assign layer0_outputs[647] = ~(inputs[28]);
    assign layer0_outputs[648] = (inputs[1]) ^ (inputs[166]);
    assign layer0_outputs[649] = ~((inputs[173]) | (inputs[232]));
    assign layer0_outputs[650] = ~(inputs[102]);
    assign layer0_outputs[651] = 1'b0;
    assign layer0_outputs[652] = ~(inputs[26]);
    assign layer0_outputs[653] = (inputs[100]) | (inputs[199]);
    assign layer0_outputs[654] = inputs[193];
    assign layer0_outputs[655] = inputs[41];
    assign layer0_outputs[656] = ~(inputs[181]);
    assign layer0_outputs[657] = ~((inputs[184]) & (inputs[164]));
    assign layer0_outputs[658] = ~((inputs[169]) | (inputs[142]));
    assign layer0_outputs[659] = ~(inputs[208]);
    assign layer0_outputs[660] = ~((inputs[41]) | (inputs[75]));
    assign layer0_outputs[661] = 1'b1;
    assign layer0_outputs[662] = (inputs[84]) | (inputs[80]);
    assign layer0_outputs[663] = ~((inputs[112]) | (inputs[37]));
    assign layer0_outputs[664] = (inputs[182]) & (inputs[121]);
    assign layer0_outputs[665] = ~(inputs[196]);
    assign layer0_outputs[666] = ~(inputs[145]) | (inputs[240]);
    assign layer0_outputs[667] = inputs[166];
    assign layer0_outputs[668] = ~((inputs[254]) | (inputs[174]));
    assign layer0_outputs[669] = ~(inputs[154]);
    assign layer0_outputs[670] = ~((inputs[2]) | (inputs[18]));
    assign layer0_outputs[671] = inputs[164];
    assign layer0_outputs[672] = (inputs[205]) & (inputs[44]);
    assign layer0_outputs[673] = ~(inputs[27]) | (inputs[83]);
    assign layer0_outputs[674] = (inputs[207]) | (inputs[110]);
    assign layer0_outputs[675] = (inputs[168]) | (inputs[144]);
    assign layer0_outputs[676] = ~(inputs[53]) | (inputs[17]);
    assign layer0_outputs[677] = inputs[178];
    assign layer0_outputs[678] = (inputs[13]) ^ (inputs[44]);
    assign layer0_outputs[679] = inputs[9];
    assign layer0_outputs[680] = (inputs[12]) & ~(inputs[220]);
    assign layer0_outputs[681] = ~(inputs[113]);
    assign layer0_outputs[682] = (inputs[225]) ^ (inputs[195]);
    assign layer0_outputs[683] = ~((inputs[126]) ^ (inputs[143]));
    assign layer0_outputs[684] = inputs[204];
    assign layer0_outputs[685] = inputs[230];
    assign layer0_outputs[686] = (inputs[9]) & ~(inputs[137]);
    assign layer0_outputs[687] = ~((inputs[58]) & (inputs[157]));
    assign layer0_outputs[688] = 1'b1;
    assign layer0_outputs[689] = (inputs[79]) & ~(inputs[105]);
    assign layer0_outputs[690] = inputs[90];
    assign layer0_outputs[691] = (inputs[62]) & (inputs[95]);
    assign layer0_outputs[692] = (inputs[18]) ^ (inputs[153]);
    assign layer0_outputs[693] = ~(inputs[140]) | (inputs[72]);
    assign layer0_outputs[694] = (inputs[208]) & ~(inputs[124]);
    assign layer0_outputs[695] = 1'b0;
    assign layer0_outputs[696] = (inputs[101]) ^ (inputs[198]);
    assign layer0_outputs[697] = inputs[63];
    assign layer0_outputs[698] = (inputs[212]) | (inputs[104]);
    assign layer0_outputs[699] = (inputs[169]) ^ (inputs[118]);
    assign layer0_outputs[700] = 1'b0;
    assign layer0_outputs[701] = (inputs[10]) & ~(inputs[217]);
    assign layer0_outputs[702] = inputs[127];
    assign layer0_outputs[703] = ~(inputs[99]);
    assign layer0_outputs[704] = (inputs[87]) & ~(inputs[221]);
    assign layer0_outputs[705] = ~(inputs[117]);
    assign layer0_outputs[706] = inputs[154];
    assign layer0_outputs[707] = ~(inputs[174]);
    assign layer0_outputs[708] = (inputs[209]) & (inputs[116]);
    assign layer0_outputs[709] = ~((inputs[189]) | (inputs[23]));
    assign layer0_outputs[710] = ~(inputs[108]) | (inputs[133]);
    assign layer0_outputs[711] = (inputs[230]) & ~(inputs[80]);
    assign layer0_outputs[712] = ~(inputs[100]) | (inputs[94]);
    assign layer0_outputs[713] = ~((inputs[208]) | (inputs[163]));
    assign layer0_outputs[714] = ~(inputs[159]) | (inputs[13]);
    assign layer0_outputs[715] = (inputs[243]) | (inputs[204]);
    assign layer0_outputs[716] = ~((inputs[219]) | (inputs[215]));
    assign layer0_outputs[717] = (inputs[110]) ^ (inputs[14]);
    assign layer0_outputs[718] = ~(inputs[24]);
    assign layer0_outputs[719] = inputs[22];
    assign layer0_outputs[720] = (inputs[74]) & ~(inputs[252]);
    assign layer0_outputs[721] = (inputs[254]) & ~(inputs[40]);
    assign layer0_outputs[722] = ~((inputs[27]) ^ (inputs[153]));
    assign layer0_outputs[723] = ~(inputs[90]);
    assign layer0_outputs[724] = ~(inputs[59]) | (inputs[71]);
    assign layer0_outputs[725] = ~(inputs[85]);
    assign layer0_outputs[726] = (inputs[170]) | (inputs[98]);
    assign layer0_outputs[727] = (inputs[98]) ^ (inputs[115]);
    assign layer0_outputs[728] = ~(inputs[119]) | (inputs[178]);
    assign layer0_outputs[729] = ~((inputs[246]) ^ (inputs[215]));
    assign layer0_outputs[730] = ~(inputs[179]) | (inputs[94]);
    assign layer0_outputs[731] = ~(inputs[48]);
    assign layer0_outputs[732] = ~(inputs[244]);
    assign layer0_outputs[733] = (inputs[251]) ^ (inputs[105]);
    assign layer0_outputs[734] = ~(inputs[38]);
    assign layer0_outputs[735] = (inputs[237]) & ~(inputs[128]);
    assign layer0_outputs[736] = (inputs[214]) ^ (inputs[212]);
    assign layer0_outputs[737] = ~((inputs[47]) & (inputs[32]));
    assign layer0_outputs[738] = ~(inputs[141]);
    assign layer0_outputs[739] = inputs[33];
    assign layer0_outputs[740] = (inputs[156]) & ~(inputs[153]);
    assign layer0_outputs[741] = (inputs[150]) & ~(inputs[220]);
    assign layer0_outputs[742] = (inputs[147]) ^ (inputs[113]);
    assign layer0_outputs[743] = 1'b0;
    assign layer0_outputs[744] = inputs[69];
    assign layer0_outputs[745] = (inputs[150]) & ~(inputs[249]);
    assign layer0_outputs[746] = ~((inputs[143]) | (inputs[138]));
    assign layer0_outputs[747] = (inputs[239]) & ~(inputs[250]);
    assign layer0_outputs[748] = inputs[234];
    assign layer0_outputs[749] = ~((inputs[72]) & (inputs[72]));
    assign layer0_outputs[750] = inputs[168];
    assign layer0_outputs[751] = ~((inputs[25]) ^ (inputs[220]));
    assign layer0_outputs[752] = ~((inputs[251]) | (inputs[198]));
    assign layer0_outputs[753] = (inputs[173]) ^ (inputs[68]);
    assign layer0_outputs[754] = (inputs[158]) | (inputs[225]);
    assign layer0_outputs[755] = ~((inputs[248]) | (inputs[229]));
    assign layer0_outputs[756] = (inputs[196]) ^ (inputs[110]);
    assign layer0_outputs[757] = (inputs[116]) & ~(inputs[245]);
    assign layer0_outputs[758] = (inputs[220]) ^ (inputs[192]);
    assign layer0_outputs[759] = (inputs[62]) ^ (inputs[122]);
    assign layer0_outputs[760] = (inputs[182]) & ~(inputs[58]);
    assign layer0_outputs[761] = (inputs[183]) & ~(inputs[130]);
    assign layer0_outputs[762] = inputs[235];
    assign layer0_outputs[763] = ~(inputs[104]);
    assign layer0_outputs[764] = ~((inputs[64]) ^ (inputs[173]));
    assign layer0_outputs[765] = (inputs[184]) | (inputs[170]);
    assign layer0_outputs[766] = (inputs[137]) & ~(inputs[48]);
    assign layer0_outputs[767] = inputs[23];
    assign layer0_outputs[768] = inputs[154];
    assign layer0_outputs[769] = (inputs[79]) | (inputs[178]);
    assign layer0_outputs[770] = (inputs[213]) & (inputs[71]);
    assign layer0_outputs[771] = (inputs[48]) ^ (inputs[137]);
    assign layer0_outputs[772] = ~(inputs[156]) | (inputs[37]);
    assign layer0_outputs[773] = ~((inputs[194]) | (inputs[4]));
    assign layer0_outputs[774] = ~((inputs[210]) & (inputs[143]));
    assign layer0_outputs[775] = (inputs[191]) & ~(inputs[223]);
    assign layer0_outputs[776] = (inputs[83]) | (inputs[69]);
    assign layer0_outputs[777] = inputs[187];
    assign layer0_outputs[778] = inputs[234];
    assign layer0_outputs[779] = ~(inputs[141]) | (inputs[44]);
    assign layer0_outputs[780] = ~(inputs[79]);
    assign layer0_outputs[781] = ~(inputs[76]) | (inputs[197]);
    assign layer0_outputs[782] = ~(inputs[43]);
    assign layer0_outputs[783] = ~(inputs[181]) | (inputs[166]);
    assign layer0_outputs[784] = ~((inputs[154]) | (inputs[163]));
    assign layer0_outputs[785] = inputs[45];
    assign layer0_outputs[786] = inputs[166];
    assign layer0_outputs[787] = (inputs[26]) | (inputs[208]);
    assign layer0_outputs[788] = (inputs[149]) & (inputs[90]);
    assign layer0_outputs[789] = 1'b1;
    assign layer0_outputs[790] = (inputs[61]) | (inputs[101]);
    assign layer0_outputs[791] = ~((inputs[193]) | (inputs[47]));
    assign layer0_outputs[792] = ~((inputs[175]) | (inputs[166]));
    assign layer0_outputs[793] = (inputs[139]) & (inputs[75]);
    assign layer0_outputs[794] = (inputs[97]) & ~(inputs[106]);
    assign layer0_outputs[795] = ~((inputs[51]) ^ (inputs[102]));
    assign layer0_outputs[796] = ~(inputs[152]) | (inputs[55]);
    assign layer0_outputs[797] = inputs[151];
    assign layer0_outputs[798] = ~(inputs[210]);
    assign layer0_outputs[799] = inputs[75];
    assign layer0_outputs[800] = ~(inputs[28]);
    assign layer0_outputs[801] = ~((inputs[238]) ^ (inputs[106]));
    assign layer0_outputs[802] = ~(inputs[162]);
    assign layer0_outputs[803] = ~(inputs[18]) | (inputs[239]);
    assign layer0_outputs[804] = ~(inputs[167]) | (inputs[116]);
    assign layer0_outputs[805] = ~(inputs[88]) | (inputs[33]);
    assign layer0_outputs[806] = ~(inputs[153]);
    assign layer0_outputs[807] = (inputs[56]) & (inputs[29]);
    assign layer0_outputs[808] = inputs[41];
    assign layer0_outputs[809] = ~(inputs[255]) | (inputs[247]);
    assign layer0_outputs[810] = inputs[167];
    assign layer0_outputs[811] = (inputs[144]) ^ (inputs[104]);
    assign layer0_outputs[812] = inputs[75];
    assign layer0_outputs[813] = ~((inputs[6]) & (inputs[81]));
    assign layer0_outputs[814] = inputs[234];
    assign layer0_outputs[815] = (inputs[198]) & ~(inputs[82]);
    assign layer0_outputs[816] = (inputs[42]) ^ (inputs[61]);
    assign layer0_outputs[817] = ~((inputs[185]) | (inputs[65]));
    assign layer0_outputs[818] = ~((inputs[194]) ^ (inputs[55]));
    assign layer0_outputs[819] = ~(inputs[67]);
    assign layer0_outputs[820] = (inputs[150]) & ~(inputs[175]);
    assign layer0_outputs[821] = (inputs[186]) ^ (inputs[207]);
    assign layer0_outputs[822] = (inputs[232]) | (inputs[249]);
    assign layer0_outputs[823] = ~(inputs[7]) | (inputs[236]);
    assign layer0_outputs[824] = (inputs[40]) & ~(inputs[61]);
    assign layer0_outputs[825] = ~((inputs[111]) ^ (inputs[138]));
    assign layer0_outputs[826] = ~(inputs[87]);
    assign layer0_outputs[827] = ~((inputs[28]) | (inputs[66]));
    assign layer0_outputs[828] = ~(inputs[51]) | (inputs[165]);
    assign layer0_outputs[829] = inputs[4];
    assign layer0_outputs[830] = ~(inputs[122]) | (inputs[131]);
    assign layer0_outputs[831] = (inputs[2]) & (inputs[207]);
    assign layer0_outputs[832] = ~(inputs[79]) | (inputs[48]);
    assign layer0_outputs[833] = ~((inputs[74]) ^ (inputs[0]));
    assign layer0_outputs[834] = (inputs[141]) & ~(inputs[253]);
    assign layer0_outputs[835] = (inputs[144]) & ~(inputs[16]);
    assign layer0_outputs[836] = inputs[152];
    assign layer0_outputs[837] = ~(inputs[228]);
    assign layer0_outputs[838] = 1'b1;
    assign layer0_outputs[839] = ~((inputs[98]) | (inputs[193]));
    assign layer0_outputs[840] = (inputs[20]) & ~(inputs[220]);
    assign layer0_outputs[841] = 1'b1;
    assign layer0_outputs[842] = ~(inputs[80]);
    assign layer0_outputs[843] = ~(inputs[200]);
    assign layer0_outputs[844] = (inputs[171]) ^ (inputs[124]);
    assign layer0_outputs[845] = ~(inputs[231]);
    assign layer0_outputs[846] = (inputs[89]) | (inputs[180]);
    assign layer0_outputs[847] = (inputs[158]) | (inputs[184]);
    assign layer0_outputs[848] = ~((inputs[211]) & (inputs[123]));
    assign layer0_outputs[849] = ~((inputs[163]) ^ (inputs[126]));
    assign layer0_outputs[850] = ~((inputs[241]) ^ (inputs[191]));
    assign layer0_outputs[851] = ~((inputs[212]) | (inputs[189]));
    assign layer0_outputs[852] = inputs[213];
    assign layer0_outputs[853] = (inputs[114]) ^ (inputs[252]);
    assign layer0_outputs[854] = inputs[181];
    assign layer0_outputs[855] = inputs[54];
    assign layer0_outputs[856] = ~(inputs[155]);
    assign layer0_outputs[857] = inputs[51];
    assign layer0_outputs[858] = ~(inputs[204]);
    assign layer0_outputs[859] = inputs[181];
    assign layer0_outputs[860] = ~((inputs[7]) ^ (inputs[26]));
    assign layer0_outputs[861] = inputs[172];
    assign layer0_outputs[862] = (inputs[49]) & ~(inputs[178]);
    assign layer0_outputs[863] = ~((inputs[183]) ^ (inputs[45]));
    assign layer0_outputs[864] = ~(inputs[149]) | (inputs[18]);
    assign layer0_outputs[865] = (inputs[201]) ^ (inputs[209]);
    assign layer0_outputs[866] = (inputs[158]) | (inputs[77]);
    assign layer0_outputs[867] = (inputs[109]) & ~(inputs[98]);
    assign layer0_outputs[868] = (inputs[251]) | (inputs[15]);
    assign layer0_outputs[869] = (inputs[50]) & ~(inputs[35]);
    assign layer0_outputs[870] = ~((inputs[137]) & (inputs[19]));
    assign layer0_outputs[871] = ~(inputs[248]);
    assign layer0_outputs[872] = ~((inputs[83]) ^ (inputs[222]));
    assign layer0_outputs[873] = ~(inputs[38]) | (inputs[44]);
    assign layer0_outputs[874] = ~(inputs[136]);
    assign layer0_outputs[875] = (inputs[154]) | (inputs[51]);
    assign layer0_outputs[876] = ~(inputs[95]);
    assign layer0_outputs[877] = inputs[57];
    assign layer0_outputs[878] = ~((inputs[24]) | (inputs[107]));
    assign layer0_outputs[879] = (inputs[229]) ^ (inputs[190]);
    assign layer0_outputs[880] = (inputs[21]) & ~(inputs[160]);
    assign layer0_outputs[881] = (inputs[115]) & ~(inputs[186]);
    assign layer0_outputs[882] = ~(inputs[23]) | (inputs[181]);
    assign layer0_outputs[883] = (inputs[144]) ^ (inputs[15]);
    assign layer0_outputs[884] = ~((inputs[159]) ^ (inputs[195]));
    assign layer0_outputs[885] = ~(inputs[80]);
    assign layer0_outputs[886] = (inputs[87]) | (inputs[202]);
    assign layer0_outputs[887] = (inputs[192]) ^ (inputs[244]);
    assign layer0_outputs[888] = (inputs[89]) & ~(inputs[32]);
    assign layer0_outputs[889] = inputs[63];
    assign layer0_outputs[890] = ~(inputs[128]);
    assign layer0_outputs[891] = inputs[96];
    assign layer0_outputs[892] = (inputs[211]) | (inputs[178]);
    assign layer0_outputs[893] = 1'b0;
    assign layer0_outputs[894] = inputs[178];
    assign layer0_outputs[895] = ~(inputs[170]);
    assign layer0_outputs[896] = (inputs[251]) | (inputs[98]);
    assign layer0_outputs[897] = inputs[162];
    assign layer0_outputs[898] = ~((inputs[186]) & (inputs[163]));
    assign layer0_outputs[899] = (inputs[17]) ^ (inputs[94]);
    assign layer0_outputs[900] = ~((inputs[98]) | (inputs[172]));
    assign layer0_outputs[901] = (inputs[177]) ^ (inputs[82]);
    assign layer0_outputs[902] = (inputs[184]) & (inputs[141]);
    assign layer0_outputs[903] = ~((inputs[113]) | (inputs[138]));
    assign layer0_outputs[904] = (inputs[219]) | (inputs[20]);
    assign layer0_outputs[905] = 1'b0;
    assign layer0_outputs[906] = (inputs[243]) | (inputs[48]);
    assign layer0_outputs[907] = ~(inputs[36]) | (inputs[206]);
    assign layer0_outputs[908] = ~(inputs[120]);
    assign layer0_outputs[909] = ~(inputs[227]) | (inputs[12]);
    assign layer0_outputs[910] = ~(inputs[169]) | (inputs[68]);
    assign layer0_outputs[911] = ~((inputs[109]) | (inputs[142]));
    assign layer0_outputs[912] = ~(inputs[243]);
    assign layer0_outputs[913] = ~(inputs[218]);
    assign layer0_outputs[914] = (inputs[173]) & ~(inputs[244]);
    assign layer0_outputs[915] = ~(inputs[213]);
    assign layer0_outputs[916] = ~(inputs[224]);
    assign layer0_outputs[917] = ~(inputs[98]);
    assign layer0_outputs[918] = (inputs[62]) & ~(inputs[134]);
    assign layer0_outputs[919] = (inputs[200]) & ~(inputs[47]);
    assign layer0_outputs[920] = ~(inputs[162]) | (inputs[49]);
    assign layer0_outputs[921] = (inputs[247]) & ~(inputs[18]);
    assign layer0_outputs[922] = ~(inputs[206]);
    assign layer0_outputs[923] = inputs[205];
    assign layer0_outputs[924] = ~(inputs[212]);
    assign layer0_outputs[925] = ~(inputs[163]) | (inputs[36]);
    assign layer0_outputs[926] = (inputs[61]) & ~(inputs[210]);
    assign layer0_outputs[927] = ~(inputs[158]);
    assign layer0_outputs[928] = (inputs[61]) ^ (inputs[75]);
    assign layer0_outputs[929] = ~(inputs[228]);
    assign layer0_outputs[930] = ~(inputs[6]);
    assign layer0_outputs[931] = (inputs[186]) & ~(inputs[95]);
    assign layer0_outputs[932] = (inputs[174]) | (inputs[45]);
    assign layer0_outputs[933] = inputs[200];
    assign layer0_outputs[934] = (inputs[61]) ^ (inputs[28]);
    assign layer0_outputs[935] = inputs[64];
    assign layer0_outputs[936] = ~(inputs[233]);
    assign layer0_outputs[937] = ~(inputs[143]) | (inputs[24]);
    assign layer0_outputs[938] = inputs[151];
    assign layer0_outputs[939] = ~(inputs[122]) | (inputs[95]);
    assign layer0_outputs[940] = (inputs[248]) ^ (inputs[208]);
    assign layer0_outputs[941] = ~(inputs[171]);
    assign layer0_outputs[942] = ~((inputs[253]) | (inputs[233]));
    assign layer0_outputs[943] = (inputs[15]) | (inputs[36]);
    assign layer0_outputs[944] = inputs[213];
    assign layer0_outputs[945] = 1'b0;
    assign layer0_outputs[946] = (inputs[104]) ^ (inputs[148]);
    assign layer0_outputs[947] = 1'b0;
    assign layer0_outputs[948] = (inputs[4]) ^ (inputs[115]);
    assign layer0_outputs[949] = ~(inputs[140]) | (inputs[241]);
    assign layer0_outputs[950] = inputs[116];
    assign layer0_outputs[951] = inputs[167];
    assign layer0_outputs[952] = (inputs[159]) & ~(inputs[114]);
    assign layer0_outputs[953] = (inputs[158]) | (inputs[192]);
    assign layer0_outputs[954] = (inputs[35]) & ~(inputs[253]);
    assign layer0_outputs[955] = ~(inputs[218]);
    assign layer0_outputs[956] = ~(inputs[213]);
    assign layer0_outputs[957] = (inputs[165]) ^ (inputs[168]);
    assign layer0_outputs[958] = (inputs[122]) & ~(inputs[65]);
    assign layer0_outputs[959] = inputs[56];
    assign layer0_outputs[960] = ~(inputs[183]) | (inputs[61]);
    assign layer0_outputs[961] = ~(inputs[241]) | (inputs[251]);
    assign layer0_outputs[962] = ~((inputs[255]) & (inputs[138]));
    assign layer0_outputs[963] = (inputs[226]) & ~(inputs[94]);
    assign layer0_outputs[964] = (inputs[76]) & ~(inputs[254]);
    assign layer0_outputs[965] = ~(inputs[8]) | (inputs[240]);
    assign layer0_outputs[966] = (inputs[202]) | (inputs[212]);
    assign layer0_outputs[967] = 1'b0;
    assign layer0_outputs[968] = inputs[123];
    assign layer0_outputs[969] = 1'b1;
    assign layer0_outputs[970] = ~((inputs[36]) ^ (inputs[162]));
    assign layer0_outputs[971] = ~(inputs[167]);
    assign layer0_outputs[972] = (inputs[184]) & (inputs[48]);
    assign layer0_outputs[973] = ~((inputs[11]) ^ (inputs[224]));
    assign layer0_outputs[974] = ~((inputs[26]) ^ (inputs[232]));
    assign layer0_outputs[975] = inputs[93];
    assign layer0_outputs[976] = ~((inputs[20]) | (inputs[5]));
    assign layer0_outputs[977] = ~((inputs[45]) ^ (inputs[59]));
    assign layer0_outputs[978] = ~(inputs[182]);
    assign layer0_outputs[979] = 1'b1;
    assign layer0_outputs[980] = ~(inputs[132]);
    assign layer0_outputs[981] = inputs[168];
    assign layer0_outputs[982] = ~((inputs[118]) | (inputs[192]));
    assign layer0_outputs[983] = ~(inputs[139]) | (inputs[107]);
    assign layer0_outputs[984] = ~((inputs[37]) | (inputs[98]));
    assign layer0_outputs[985] = 1'b0;
    assign layer0_outputs[986] = ~((inputs[101]) | (inputs[233]));
    assign layer0_outputs[987] = ~((inputs[33]) | (inputs[58]));
    assign layer0_outputs[988] = ~(inputs[18]);
    assign layer0_outputs[989] = (inputs[132]) ^ (inputs[112]);
    assign layer0_outputs[990] = (inputs[180]) | (inputs[158]);
    assign layer0_outputs[991] = inputs[8];
    assign layer0_outputs[992] = inputs[144];
    assign layer0_outputs[993] = (inputs[213]) & ~(inputs[39]);
    assign layer0_outputs[994] = ~(inputs[25]);
    assign layer0_outputs[995] = 1'b0;
    assign layer0_outputs[996] = (inputs[118]) ^ (inputs[166]);
    assign layer0_outputs[997] = inputs[232];
    assign layer0_outputs[998] = (inputs[121]) ^ (inputs[2]);
    assign layer0_outputs[999] = 1'b1;
    assign layer0_outputs[1000] = inputs[88];
    assign layer0_outputs[1001] = (inputs[241]) & ~(inputs[140]);
    assign layer0_outputs[1002] = ~(inputs[62]);
    assign layer0_outputs[1003] = (inputs[195]) | (inputs[82]);
    assign layer0_outputs[1004] = (inputs[114]) | (inputs[133]);
    assign layer0_outputs[1005] = ~((inputs[244]) | (inputs[190]));
    assign layer0_outputs[1006] = 1'b1;
    assign layer0_outputs[1007] = inputs[218];
    assign layer0_outputs[1008] = inputs[85];
    assign layer0_outputs[1009] = ~(inputs[77]);
    assign layer0_outputs[1010] = ~(inputs[131]);
    assign layer0_outputs[1011] = (inputs[98]) | (inputs[132]);
    assign layer0_outputs[1012] = inputs[166];
    assign layer0_outputs[1013] = inputs[56];
    assign layer0_outputs[1014] = ~(inputs[104]) | (inputs[114]);
    assign layer0_outputs[1015] = (inputs[117]) & (inputs[39]);
    assign layer0_outputs[1016] = (inputs[151]) | (inputs[2]);
    assign layer0_outputs[1017] = ~(inputs[153]);
    assign layer0_outputs[1018] = (inputs[89]) ^ (inputs[145]);
    assign layer0_outputs[1019] = ~(inputs[229]);
    assign layer0_outputs[1020] = (inputs[229]) ^ (inputs[161]);
    assign layer0_outputs[1021] = (inputs[152]) | (inputs[163]);
    assign layer0_outputs[1022] = inputs[169];
    assign layer0_outputs[1023] = (inputs[255]) | (inputs[141]);
    assign layer0_outputs[1024] = (inputs[171]) & ~(inputs[119]);
    assign layer0_outputs[1025] = ~(inputs[149]) | (inputs[4]);
    assign layer0_outputs[1026] = (inputs[71]) | (inputs[157]);
    assign layer0_outputs[1027] = ~((inputs[227]) | (inputs[233]));
    assign layer0_outputs[1028] = ~(inputs[244]) | (inputs[113]);
    assign layer0_outputs[1029] = ~(inputs[89]);
    assign layer0_outputs[1030] = ~(inputs[165]);
    assign layer0_outputs[1031] = ~(inputs[229]) | (inputs[109]);
    assign layer0_outputs[1032] = inputs[69];
    assign layer0_outputs[1033] = ~(inputs[100]) | (inputs[225]);
    assign layer0_outputs[1034] = ~((inputs[62]) | (inputs[223]));
    assign layer0_outputs[1035] = inputs[173];
    assign layer0_outputs[1036] = ~(inputs[131]);
    assign layer0_outputs[1037] = ~(inputs[39]);
    assign layer0_outputs[1038] = (inputs[166]) ^ (inputs[163]);
    assign layer0_outputs[1039] = ~(inputs[28]);
    assign layer0_outputs[1040] = (inputs[109]) ^ (inputs[60]);
    assign layer0_outputs[1041] = (inputs[237]) & (inputs[143]);
    assign layer0_outputs[1042] = inputs[177];
    assign layer0_outputs[1043] = ~(inputs[56]) | (inputs[173]);
    assign layer0_outputs[1044] = ~(inputs[180]) | (inputs[54]);
    assign layer0_outputs[1045] = ~(inputs[0]) | (inputs[215]);
    assign layer0_outputs[1046] = (inputs[127]) ^ (inputs[65]);
    assign layer0_outputs[1047] = (inputs[49]) ^ (inputs[53]);
    assign layer0_outputs[1048] = ~((inputs[144]) | (inputs[114]));
    assign layer0_outputs[1049] = inputs[122];
    assign layer0_outputs[1050] = inputs[236];
    assign layer0_outputs[1051] = ~((inputs[173]) & (inputs[111]));
    assign layer0_outputs[1052] = inputs[122];
    assign layer0_outputs[1053] = ~(inputs[119]);
    assign layer0_outputs[1054] = (inputs[179]) & (inputs[148]);
    assign layer0_outputs[1055] = (inputs[13]) & (inputs[238]);
    assign layer0_outputs[1056] = ~(inputs[181]) | (inputs[98]);
    assign layer0_outputs[1057] = ~((inputs[166]) & (inputs[119]));
    assign layer0_outputs[1058] = inputs[248];
    assign layer0_outputs[1059] = (inputs[204]) & ~(inputs[29]);
    assign layer0_outputs[1060] = (inputs[67]) & ~(inputs[2]);
    assign layer0_outputs[1061] = (inputs[170]) | (inputs[133]);
    assign layer0_outputs[1062] = ~(inputs[50]) | (inputs[231]);
    assign layer0_outputs[1063] = ~((inputs[125]) ^ (inputs[1]));
    assign layer0_outputs[1064] = (inputs[154]) & ~(inputs[169]);
    assign layer0_outputs[1065] = (inputs[106]) & ~(inputs[227]);
    assign layer0_outputs[1066] = (inputs[58]) & ~(inputs[227]);
    assign layer0_outputs[1067] = ~(inputs[115]);
    assign layer0_outputs[1068] = ~((inputs[155]) & (inputs[39]));
    assign layer0_outputs[1069] = inputs[146];
    assign layer0_outputs[1070] = ~((inputs[31]) ^ (inputs[137]));
    assign layer0_outputs[1071] = ~(inputs[45]);
    assign layer0_outputs[1072] = inputs[130];
    assign layer0_outputs[1073] = ~((inputs[163]) | (inputs[176]));
    assign layer0_outputs[1074] = inputs[116];
    assign layer0_outputs[1075] = ~(inputs[66]);
    assign layer0_outputs[1076] = ~(inputs[91]) | (inputs[123]);
    assign layer0_outputs[1077] = (inputs[35]) | (inputs[234]);
    assign layer0_outputs[1078] = ~(inputs[8]);
    assign layer0_outputs[1079] = ~(inputs[167]);
    assign layer0_outputs[1080] = ~(inputs[126]) | (inputs[174]);
    assign layer0_outputs[1081] = ~((inputs[57]) ^ (inputs[72]));
    assign layer0_outputs[1082] = ~(inputs[42]);
    assign layer0_outputs[1083] = ~((inputs[144]) & (inputs[28]));
    assign layer0_outputs[1084] = ~(inputs[36]);
    assign layer0_outputs[1085] = (inputs[62]) ^ (inputs[79]);
    assign layer0_outputs[1086] = (inputs[70]) & ~(inputs[59]);
    assign layer0_outputs[1087] = inputs[38];
    assign layer0_outputs[1088] = inputs[56];
    assign layer0_outputs[1089] = (inputs[46]) | (inputs[54]);
    assign layer0_outputs[1090] = ~(inputs[67]);
    assign layer0_outputs[1091] = ~(inputs[253]) | (inputs[32]);
    assign layer0_outputs[1092] = inputs[161];
    assign layer0_outputs[1093] = inputs[217];
    assign layer0_outputs[1094] = (inputs[98]) | (inputs[239]);
    assign layer0_outputs[1095] = inputs[250];
    assign layer0_outputs[1096] = 1'b0;
    assign layer0_outputs[1097] = ~(inputs[220]);
    assign layer0_outputs[1098] = 1'b1;
    assign layer0_outputs[1099] = ~(inputs[230]);
    assign layer0_outputs[1100] = ~(inputs[84]);
    assign layer0_outputs[1101] = (inputs[114]) | (inputs[167]);
    assign layer0_outputs[1102] = (inputs[8]) & ~(inputs[3]);
    assign layer0_outputs[1103] = 1'b0;
    assign layer0_outputs[1104] = (inputs[120]) & ~(inputs[33]);
    assign layer0_outputs[1105] = (inputs[200]) & ~(inputs[73]);
    assign layer0_outputs[1106] = 1'b1;
    assign layer0_outputs[1107] = 1'b0;
    assign layer0_outputs[1108] = ~(inputs[7]);
    assign layer0_outputs[1109] = (inputs[177]) ^ (inputs[8]);
    assign layer0_outputs[1110] = ~((inputs[237]) & (inputs[38]));
    assign layer0_outputs[1111] = inputs[87];
    assign layer0_outputs[1112] = ~(inputs[82]);
    assign layer0_outputs[1113] = ~(inputs[168]) | (inputs[90]);
    assign layer0_outputs[1114] = (inputs[118]) | (inputs[68]);
    assign layer0_outputs[1115] = ~(inputs[34]);
    assign layer0_outputs[1116] = ~((inputs[92]) & (inputs[108]));
    assign layer0_outputs[1117] = 1'b0;
    assign layer0_outputs[1118] = ~((inputs[148]) & (inputs[251]));
    assign layer0_outputs[1119] = inputs[246];
    assign layer0_outputs[1120] = 1'b0;
    assign layer0_outputs[1121] = ~((inputs[228]) ^ (inputs[62]));
    assign layer0_outputs[1122] = ~(inputs[57]) | (inputs[83]);
    assign layer0_outputs[1123] = (inputs[139]) ^ (inputs[205]);
    assign layer0_outputs[1124] = ~((inputs[201]) | (inputs[20]));
    assign layer0_outputs[1125] = (inputs[192]) | (inputs[119]);
    assign layer0_outputs[1126] = (inputs[169]) | (inputs[120]);
    assign layer0_outputs[1127] = (inputs[102]) | (inputs[119]);
    assign layer0_outputs[1128] = (inputs[196]) & ~(inputs[78]);
    assign layer0_outputs[1129] = (inputs[251]) ^ (inputs[203]);
    assign layer0_outputs[1130] = ~((inputs[247]) | (inputs[43]));
    assign layer0_outputs[1131] = inputs[76];
    assign layer0_outputs[1132] = inputs[1];
    assign layer0_outputs[1133] = (inputs[83]) | (inputs[239]);
    assign layer0_outputs[1134] = (inputs[20]) ^ (inputs[77]);
    assign layer0_outputs[1135] = (inputs[127]) | (inputs[213]);
    assign layer0_outputs[1136] = inputs[92];
    assign layer0_outputs[1137] = (inputs[60]) ^ (inputs[28]);
    assign layer0_outputs[1138] = (inputs[238]) | (inputs[210]);
    assign layer0_outputs[1139] = ~(inputs[88]) | (inputs[239]);
    assign layer0_outputs[1140] = inputs[50];
    assign layer0_outputs[1141] = 1'b1;
    assign layer0_outputs[1142] = (inputs[1]) | (inputs[187]);
    assign layer0_outputs[1143] = ~((inputs[155]) | (inputs[196]));
    assign layer0_outputs[1144] = ~(inputs[198]) | (inputs[105]);
    assign layer0_outputs[1145] = ~(inputs[60]) | (inputs[71]);
    assign layer0_outputs[1146] = ~((inputs[127]) ^ (inputs[203]));
    assign layer0_outputs[1147] = ~((inputs[62]) | (inputs[37]));
    assign layer0_outputs[1148] = (inputs[239]) ^ (inputs[87]);
    assign layer0_outputs[1149] = 1'b0;
    assign layer0_outputs[1150] = inputs[156];
    assign layer0_outputs[1151] = ~((inputs[73]) | (inputs[226]));
    assign layer0_outputs[1152] = ~(inputs[230]);
    assign layer0_outputs[1153] = (inputs[24]) & ~(inputs[235]);
    assign layer0_outputs[1154] = inputs[201];
    assign layer0_outputs[1155] = inputs[139];
    assign layer0_outputs[1156] = ~((inputs[132]) & (inputs[214]));
    assign layer0_outputs[1157] = ~((inputs[113]) ^ (inputs[68]));
    assign layer0_outputs[1158] = ~((inputs[17]) ^ (inputs[2]));
    assign layer0_outputs[1159] = inputs[93];
    assign layer0_outputs[1160] = ~(inputs[152]) | (inputs[60]);
    assign layer0_outputs[1161] = (inputs[22]) ^ (inputs[157]);
    assign layer0_outputs[1162] = inputs[27];
    assign layer0_outputs[1163] = ~((inputs[10]) & (inputs[216]));
    assign layer0_outputs[1164] = (inputs[127]) | (inputs[183]);
    assign layer0_outputs[1165] = (inputs[86]) ^ (inputs[117]);
    assign layer0_outputs[1166] = ~((inputs[112]) ^ (inputs[210]));
    assign layer0_outputs[1167] = ~(inputs[9]);
    assign layer0_outputs[1168] = ~(inputs[200]);
    assign layer0_outputs[1169] = ~((inputs[107]) & (inputs[139]));
    assign layer0_outputs[1170] = ~(inputs[160]);
    assign layer0_outputs[1171] = inputs[195];
    assign layer0_outputs[1172] = ~(inputs[39]);
    assign layer0_outputs[1173] = ~((inputs[179]) ^ (inputs[26]));
    assign layer0_outputs[1174] = ~((inputs[243]) | (inputs[210]));
    assign layer0_outputs[1175] = ~((inputs[222]) ^ (inputs[21]));
    assign layer0_outputs[1176] = (inputs[244]) ^ (inputs[203]);
    assign layer0_outputs[1177] = (inputs[98]) ^ (inputs[165]);
    assign layer0_outputs[1178] = ~(inputs[62]);
    assign layer0_outputs[1179] = inputs[8];
    assign layer0_outputs[1180] = inputs[52];
    assign layer0_outputs[1181] = (inputs[215]) & (inputs[123]);
    assign layer0_outputs[1182] = ~((inputs[170]) & (inputs[56]));
    assign layer0_outputs[1183] = ~((inputs[199]) & (inputs[202]));
    assign layer0_outputs[1184] = inputs[62];
    assign layer0_outputs[1185] = inputs[145];
    assign layer0_outputs[1186] = (inputs[109]) | (inputs[207]);
    assign layer0_outputs[1187] = inputs[90];
    assign layer0_outputs[1188] = (inputs[189]) & ~(inputs[80]);
    assign layer0_outputs[1189] = ~((inputs[216]) ^ (inputs[11]));
    assign layer0_outputs[1190] = (inputs[0]) & ~(inputs[128]);
    assign layer0_outputs[1191] = (inputs[30]) & ~(inputs[45]);
    assign layer0_outputs[1192] = ~((inputs[57]) ^ (inputs[113]));
    assign layer0_outputs[1193] = ~(inputs[224]) | (inputs[223]);
    assign layer0_outputs[1194] = inputs[214];
    assign layer0_outputs[1195] = (inputs[181]) & ~(inputs[39]);
    assign layer0_outputs[1196] = ~((inputs[38]) ^ (inputs[136]));
    assign layer0_outputs[1197] = ~((inputs[159]) & (inputs[240]));
    assign layer0_outputs[1198] = (inputs[118]) & (inputs[120]);
    assign layer0_outputs[1199] = (inputs[140]) | (inputs[53]);
    assign layer0_outputs[1200] = ~(inputs[38]);
    assign layer0_outputs[1201] = inputs[229];
    assign layer0_outputs[1202] = (inputs[55]) & (inputs[205]);
    assign layer0_outputs[1203] = (inputs[55]) | (inputs[58]);
    assign layer0_outputs[1204] = (inputs[130]) & ~(inputs[243]);
    assign layer0_outputs[1205] = ~(inputs[22]) | (inputs[225]);
    assign layer0_outputs[1206] = inputs[230];
    assign layer0_outputs[1207] = inputs[124];
    assign layer0_outputs[1208] = (inputs[33]) | (inputs[166]);
    assign layer0_outputs[1209] = inputs[141];
    assign layer0_outputs[1210] = inputs[206];
    assign layer0_outputs[1211] = inputs[171];
    assign layer0_outputs[1212] = ~((inputs[168]) | (inputs[98]));
    assign layer0_outputs[1213] = ~(inputs[3]);
    assign layer0_outputs[1214] = ~(inputs[49]);
    assign layer0_outputs[1215] = ~(inputs[132]) | (inputs[251]);
    assign layer0_outputs[1216] = (inputs[161]) ^ (inputs[23]);
    assign layer0_outputs[1217] = inputs[85];
    assign layer0_outputs[1218] = inputs[69];
    assign layer0_outputs[1219] = ~((inputs[79]) | (inputs[162]));
    assign layer0_outputs[1220] = ~((inputs[27]) | (inputs[64]));
    assign layer0_outputs[1221] = ~((inputs[186]) | (inputs[78]));
    assign layer0_outputs[1222] = (inputs[17]) ^ (inputs[168]);
    assign layer0_outputs[1223] = ~(inputs[145]) | (inputs[62]);
    assign layer0_outputs[1224] = (inputs[92]) & ~(inputs[140]);
    assign layer0_outputs[1225] = ~(inputs[54]);
    assign layer0_outputs[1226] = ~((inputs[53]) | (inputs[200]));
    assign layer0_outputs[1227] = ~((inputs[210]) & (inputs[11]));
    assign layer0_outputs[1228] = ~((inputs[131]) ^ (inputs[127]));
    assign layer0_outputs[1229] = (inputs[77]) & ~(inputs[172]);
    assign layer0_outputs[1230] = ~(inputs[135]);
    assign layer0_outputs[1231] = (inputs[242]) ^ (inputs[189]);
    assign layer0_outputs[1232] = (inputs[107]) & ~(inputs[0]);
    assign layer0_outputs[1233] = ~(inputs[133]);
    assign layer0_outputs[1234] = (inputs[191]) | (inputs[84]);
    assign layer0_outputs[1235] = inputs[246];
    assign layer0_outputs[1236] = ~(inputs[53]) | (inputs[93]);
    assign layer0_outputs[1237] = (inputs[146]) | (inputs[51]);
    assign layer0_outputs[1238] = ~((inputs[253]) | (inputs[120]));
    assign layer0_outputs[1239] = ~((inputs[111]) ^ (inputs[5]));
    assign layer0_outputs[1240] = ~((inputs[27]) | (inputs[21]));
    assign layer0_outputs[1241] = inputs[180];
    assign layer0_outputs[1242] = (inputs[51]) ^ (inputs[71]);
    assign layer0_outputs[1243] = ~(inputs[210]);
    assign layer0_outputs[1244] = (inputs[211]) | (inputs[37]);
    assign layer0_outputs[1245] = (inputs[12]) ^ (inputs[2]);
    assign layer0_outputs[1246] = ~((inputs[130]) | (inputs[253]));
    assign layer0_outputs[1247] = ~(inputs[8]) | (inputs[127]);
    assign layer0_outputs[1248] = (inputs[10]) & (inputs[27]);
    assign layer0_outputs[1249] = ~((inputs[172]) | (inputs[100]));
    assign layer0_outputs[1250] = ~(inputs[215]);
    assign layer0_outputs[1251] = ~(inputs[122]) | (inputs[241]);
    assign layer0_outputs[1252] = (inputs[164]) | (inputs[109]);
    assign layer0_outputs[1253] = inputs[198];
    assign layer0_outputs[1254] = ~((inputs[253]) & (inputs[166]));
    assign layer0_outputs[1255] = ~(inputs[86]);
    assign layer0_outputs[1256] = ~((inputs[157]) | (inputs[77]));
    assign layer0_outputs[1257] = ~(inputs[152]) | (inputs[87]);
    assign layer0_outputs[1258] = inputs[72];
    assign layer0_outputs[1259] = (inputs[121]) & ~(inputs[194]);
    assign layer0_outputs[1260] = (inputs[245]) | (inputs[94]);
    assign layer0_outputs[1261] = (inputs[151]) ^ (inputs[34]);
    assign layer0_outputs[1262] = (inputs[189]) & ~(inputs[188]);
    assign layer0_outputs[1263] = (inputs[144]) & ~(inputs[44]);
    assign layer0_outputs[1264] = ~(inputs[137]);
    assign layer0_outputs[1265] = ~(inputs[177]);
    assign layer0_outputs[1266] = ~(inputs[180]);
    assign layer0_outputs[1267] = inputs[209];
    assign layer0_outputs[1268] = (inputs[241]) | (inputs[202]);
    assign layer0_outputs[1269] = (inputs[134]) & (inputs[44]);
    assign layer0_outputs[1270] = ~(inputs[220]);
    assign layer0_outputs[1271] = (inputs[90]) | (inputs[217]);
    assign layer0_outputs[1272] = (inputs[89]) & ~(inputs[23]);
    assign layer0_outputs[1273] = ~((inputs[209]) | (inputs[150]));
    assign layer0_outputs[1274] = inputs[160];
    assign layer0_outputs[1275] = ~(inputs[214]);
    assign layer0_outputs[1276] = ~(inputs[219]);
    assign layer0_outputs[1277] = ~((inputs[19]) | (inputs[92]));
    assign layer0_outputs[1278] = inputs[204];
    assign layer0_outputs[1279] = ~(inputs[237]) | (inputs[227]);
    assign layer0_outputs[1280] = ~((inputs[64]) | (inputs[188]));
    assign layer0_outputs[1281] = ~((inputs[133]) & (inputs[122]));
    assign layer0_outputs[1282] = ~((inputs[176]) | (inputs[156]));
    assign layer0_outputs[1283] = 1'b0;
    assign layer0_outputs[1284] = (inputs[250]) & ~(inputs[0]);
    assign layer0_outputs[1285] = 1'b0;
    assign layer0_outputs[1286] = (inputs[80]) & ~(inputs[223]);
    assign layer0_outputs[1287] = ~(inputs[123]);
    assign layer0_outputs[1288] = inputs[110];
    assign layer0_outputs[1289] = ~(inputs[216]);
    assign layer0_outputs[1290] = ~(inputs[152]) | (inputs[245]);
    assign layer0_outputs[1291] = inputs[116];
    assign layer0_outputs[1292] = (inputs[220]) | (inputs[170]);
    assign layer0_outputs[1293] = (inputs[216]) ^ (inputs[171]);
    assign layer0_outputs[1294] = inputs[94];
    assign layer0_outputs[1295] = ~(inputs[212]);
    assign layer0_outputs[1296] = inputs[91];
    assign layer0_outputs[1297] = inputs[210];
    assign layer0_outputs[1298] = (inputs[183]) ^ (inputs[196]);
    assign layer0_outputs[1299] = ~((inputs[125]) | (inputs[178]));
    assign layer0_outputs[1300] = inputs[236];
    assign layer0_outputs[1301] = ~(inputs[233]) | (inputs[83]);
    assign layer0_outputs[1302] = 1'b0;
    assign layer0_outputs[1303] = (inputs[120]) & ~(inputs[239]);
    assign layer0_outputs[1304] = ~(inputs[218]) | (inputs[143]);
    assign layer0_outputs[1305] = (inputs[99]) | (inputs[29]);
    assign layer0_outputs[1306] = ~(inputs[128]);
    assign layer0_outputs[1307] = ~(inputs[191]);
    assign layer0_outputs[1308] = inputs[158];
    assign layer0_outputs[1309] = ~(inputs[99]);
    assign layer0_outputs[1310] = ~((inputs[237]) | (inputs[199]));
    assign layer0_outputs[1311] = inputs[106];
    assign layer0_outputs[1312] = ~((inputs[193]) & (inputs[222]));
    assign layer0_outputs[1313] = ~(inputs[237]) | (inputs[86]);
    assign layer0_outputs[1314] = ~((inputs[36]) | (inputs[177]));
    assign layer0_outputs[1315] = ~((inputs[211]) & (inputs[38]));
    assign layer0_outputs[1316] = (inputs[62]) ^ (inputs[4]);
    assign layer0_outputs[1317] = (inputs[71]) & ~(inputs[123]);
    assign layer0_outputs[1318] = inputs[119];
    assign layer0_outputs[1319] = ~(inputs[108]) | (inputs[17]);
    assign layer0_outputs[1320] = inputs[73];
    assign layer0_outputs[1321] = ~(inputs[41]);
    assign layer0_outputs[1322] = (inputs[244]) & ~(inputs[219]);
    assign layer0_outputs[1323] = (inputs[183]) & ~(inputs[130]);
    assign layer0_outputs[1324] = ~(inputs[84]) | (inputs[72]);
    assign layer0_outputs[1325] = (inputs[176]) ^ (inputs[138]);
    assign layer0_outputs[1326] = inputs[98];
    assign layer0_outputs[1327] = inputs[37];
    assign layer0_outputs[1328] = (inputs[250]) & ~(inputs[49]);
    assign layer0_outputs[1329] = (inputs[159]) & (inputs[2]);
    assign layer0_outputs[1330] = (inputs[27]) | (inputs[50]);
    assign layer0_outputs[1331] = ~(inputs[122]) | (inputs[42]);
    assign layer0_outputs[1332] = (inputs[206]) | (inputs[202]);
    assign layer0_outputs[1333] = ~(inputs[105]);
    assign layer0_outputs[1334] = (inputs[41]) ^ (inputs[67]);
    assign layer0_outputs[1335] = (inputs[138]) & ~(inputs[166]);
    assign layer0_outputs[1336] = inputs[240];
    assign layer0_outputs[1337] = (inputs[51]) ^ (inputs[164]);
    assign layer0_outputs[1338] = (inputs[62]) & ~(inputs[254]);
    assign layer0_outputs[1339] = ~(inputs[79]);
    assign layer0_outputs[1340] = 1'b1;
    assign layer0_outputs[1341] = (inputs[17]) & ~(inputs[232]);
    assign layer0_outputs[1342] = (inputs[165]) & ~(inputs[111]);
    assign layer0_outputs[1343] = ~(inputs[126]);
    assign layer0_outputs[1344] = ~((inputs[253]) & (inputs[144]));
    assign layer0_outputs[1345] = ~(inputs[122]) | (inputs[27]);
    assign layer0_outputs[1346] = (inputs[107]) | (inputs[48]);
    assign layer0_outputs[1347] = (inputs[172]) ^ (inputs[190]);
    assign layer0_outputs[1348] = ~(inputs[132]) | (inputs[57]);
    assign layer0_outputs[1349] = ~(inputs[84]);
    assign layer0_outputs[1350] = ~(inputs[227]);
    assign layer0_outputs[1351] = ~((inputs[160]) | (inputs[66]));
    assign layer0_outputs[1352] = (inputs[207]) ^ (inputs[250]);
    assign layer0_outputs[1353] = inputs[102];
    assign layer0_outputs[1354] = 1'b1;
    assign layer0_outputs[1355] = (inputs[64]) & (inputs[5]);
    assign layer0_outputs[1356] = inputs[109];
    assign layer0_outputs[1357] = ~(inputs[234]) | (inputs[6]);
    assign layer0_outputs[1358] = (inputs[207]) & (inputs[109]);
    assign layer0_outputs[1359] = ~(inputs[146]) | (inputs[62]);
    assign layer0_outputs[1360] = (inputs[124]) | (inputs[8]);
    assign layer0_outputs[1361] = inputs[126];
    assign layer0_outputs[1362] = (inputs[213]) | (inputs[208]);
    assign layer0_outputs[1363] = ~(inputs[22]);
    assign layer0_outputs[1364] = (inputs[97]) | (inputs[227]);
    assign layer0_outputs[1365] = ~((inputs[174]) & (inputs[204]));
    assign layer0_outputs[1366] = ~(inputs[58]) | (inputs[117]);
    assign layer0_outputs[1367] = ~((inputs[111]) ^ (inputs[239]));
    assign layer0_outputs[1368] = ~(inputs[148]);
    assign layer0_outputs[1369] = (inputs[245]) & (inputs[202]);
    assign layer0_outputs[1370] = ~((inputs[162]) ^ (inputs[233]));
    assign layer0_outputs[1371] = ~(inputs[142]);
    assign layer0_outputs[1372] = inputs[59];
    assign layer0_outputs[1373] = ~((inputs[230]) & (inputs[165]));
    assign layer0_outputs[1374] = ~(inputs[174]) | (inputs[132]);
    assign layer0_outputs[1375] = ~(inputs[106]);
    assign layer0_outputs[1376] = ~((inputs[104]) | (inputs[31]));
    assign layer0_outputs[1377] = inputs[126];
    assign layer0_outputs[1378] = (inputs[29]) | (inputs[120]);
    assign layer0_outputs[1379] = (inputs[85]) & ~(inputs[74]);
    assign layer0_outputs[1380] = ~((inputs[97]) & (inputs[187]));
    assign layer0_outputs[1381] = 1'b1;
    assign layer0_outputs[1382] = ~(inputs[172]);
    assign layer0_outputs[1383] = ~(inputs[6]);
    assign layer0_outputs[1384] = (inputs[74]) & (inputs[100]);
    assign layer0_outputs[1385] = (inputs[231]) & (inputs[226]);
    assign layer0_outputs[1386] = ~(inputs[251]);
    assign layer0_outputs[1387] = 1'b0;
    assign layer0_outputs[1388] = ~(inputs[26]) | (inputs[252]);
    assign layer0_outputs[1389] = ~(inputs[88]);
    assign layer0_outputs[1390] = (inputs[130]) | (inputs[218]);
    assign layer0_outputs[1391] = (inputs[100]) & ~(inputs[126]);
    assign layer0_outputs[1392] = 1'b1;
    assign layer0_outputs[1393] = inputs[43];
    assign layer0_outputs[1394] = ~(inputs[20]) | (inputs[114]);
    assign layer0_outputs[1395] = inputs[126];
    assign layer0_outputs[1396] = 1'b1;
    assign layer0_outputs[1397] = ~(inputs[129]) | (inputs[66]);
    assign layer0_outputs[1398] = ~(inputs[120]) | (inputs[12]);
    assign layer0_outputs[1399] = inputs[209];
    assign layer0_outputs[1400] = ~(inputs[193]);
    assign layer0_outputs[1401] = ~((inputs[15]) ^ (inputs[147]));
    assign layer0_outputs[1402] = (inputs[182]) & ~(inputs[209]);
    assign layer0_outputs[1403] = ~(inputs[70]);
    assign layer0_outputs[1404] = (inputs[240]) ^ (inputs[139]);
    assign layer0_outputs[1405] = ~((inputs[20]) ^ (inputs[81]));
    assign layer0_outputs[1406] = ~((inputs[28]) | (inputs[160]));
    assign layer0_outputs[1407] = (inputs[175]) & ~(inputs[255]);
    assign layer0_outputs[1408] = (inputs[32]) & (inputs[99]);
    assign layer0_outputs[1409] = ~((inputs[116]) | (inputs[61]));
    assign layer0_outputs[1410] = inputs[120];
    assign layer0_outputs[1411] = inputs[239];
    assign layer0_outputs[1412] = inputs[71];
    assign layer0_outputs[1413] = (inputs[184]) & (inputs[9]);
    assign layer0_outputs[1414] = inputs[28];
    assign layer0_outputs[1415] = ~((inputs[30]) ^ (inputs[76]));
    assign layer0_outputs[1416] = 1'b0;
    assign layer0_outputs[1417] = ~((inputs[186]) | (inputs[194]));
    assign layer0_outputs[1418] = (inputs[123]) ^ (inputs[68]);
    assign layer0_outputs[1419] = (inputs[13]) | (inputs[176]);
    assign layer0_outputs[1420] = (inputs[121]) & ~(inputs[168]);
    assign layer0_outputs[1421] = ~(inputs[9]);
    assign layer0_outputs[1422] = (inputs[26]) & ~(inputs[201]);
    assign layer0_outputs[1423] = inputs[113];
    assign layer0_outputs[1424] = ~((inputs[128]) ^ (inputs[231]));
    assign layer0_outputs[1425] = inputs[201];
    assign layer0_outputs[1426] = ~(inputs[94]);
    assign layer0_outputs[1427] = ~(inputs[8]) | (inputs[241]);
    assign layer0_outputs[1428] = (inputs[13]) | (inputs[92]);
    assign layer0_outputs[1429] = (inputs[222]) | (inputs[203]);
    assign layer0_outputs[1430] = ~(inputs[134]) | (inputs[43]);
    assign layer0_outputs[1431] = ~((inputs[148]) ^ (inputs[151]));
    assign layer0_outputs[1432] = ~(inputs[205]) | (inputs[198]);
    assign layer0_outputs[1433] = ~((inputs[167]) & (inputs[110]));
    assign layer0_outputs[1434] = (inputs[69]) | (inputs[130]);
    assign layer0_outputs[1435] = (inputs[203]) & (inputs[95]);
    assign layer0_outputs[1436] = ~(inputs[228]) | (inputs[132]);
    assign layer0_outputs[1437] = ~((inputs[205]) | (inputs[188]));
    assign layer0_outputs[1438] = inputs[152];
    assign layer0_outputs[1439] = ~((inputs[18]) ^ (inputs[26]));
    assign layer0_outputs[1440] = (inputs[7]) | (inputs[109]);
    assign layer0_outputs[1441] = (inputs[231]) & (inputs[181]);
    assign layer0_outputs[1442] = ~(inputs[124]);
    assign layer0_outputs[1443] = ~(inputs[157]);
    assign layer0_outputs[1444] = inputs[134];
    assign layer0_outputs[1445] = (inputs[132]) | (inputs[80]);
    assign layer0_outputs[1446] = inputs[144];
    assign layer0_outputs[1447] = ~((inputs[222]) | (inputs[201]));
    assign layer0_outputs[1448] = ~(inputs[157]) | (inputs[65]);
    assign layer0_outputs[1449] = inputs[202];
    assign layer0_outputs[1450] = (inputs[45]) ^ (inputs[19]);
    assign layer0_outputs[1451] = (inputs[64]) ^ (inputs[126]);
    assign layer0_outputs[1452] = inputs[3];
    assign layer0_outputs[1453] = (inputs[48]) | (inputs[80]);
    assign layer0_outputs[1454] = (inputs[47]) & ~(inputs[255]);
    assign layer0_outputs[1455] = (inputs[101]) | (inputs[143]);
    assign layer0_outputs[1456] = (inputs[150]) | (inputs[164]);
    assign layer0_outputs[1457] = inputs[214];
    assign layer0_outputs[1458] = ~(inputs[199]) | (inputs[97]);
    assign layer0_outputs[1459] = inputs[226];
    assign layer0_outputs[1460] = ~(inputs[40]);
    assign layer0_outputs[1461] = 1'b1;
    assign layer0_outputs[1462] = ~(inputs[137]);
    assign layer0_outputs[1463] = (inputs[183]) | (inputs[86]);
    assign layer0_outputs[1464] = ~(inputs[99]) | (inputs[30]);
    assign layer0_outputs[1465] = inputs[87];
    assign layer0_outputs[1466] = (inputs[226]) & ~(inputs[124]);
    assign layer0_outputs[1467] = ~((inputs[4]) ^ (inputs[60]));
    assign layer0_outputs[1468] = ~(inputs[165]);
    assign layer0_outputs[1469] = (inputs[109]) & ~(inputs[249]);
    assign layer0_outputs[1470] = ~(inputs[41]);
    assign layer0_outputs[1471] = ~(inputs[128]);
    assign layer0_outputs[1472] = ~(inputs[213]) | (inputs[143]);
    assign layer0_outputs[1473] = (inputs[31]) & ~(inputs[129]);
    assign layer0_outputs[1474] = ~(inputs[120]);
    assign layer0_outputs[1475] = ~(inputs[55]);
    assign layer0_outputs[1476] = (inputs[188]) | (inputs[204]);
    assign layer0_outputs[1477] = inputs[96];
    assign layer0_outputs[1478] = (inputs[54]) & ~(inputs[74]);
    assign layer0_outputs[1479] = ~((inputs[186]) & (inputs[179]));
    assign layer0_outputs[1480] = inputs[98];
    assign layer0_outputs[1481] = (inputs[165]) | (inputs[161]);
    assign layer0_outputs[1482] = ~(inputs[120]);
    assign layer0_outputs[1483] = ~((inputs[2]) & (inputs[5]));
    assign layer0_outputs[1484] = (inputs[170]) | (inputs[63]);
    assign layer0_outputs[1485] = (inputs[99]) ^ (inputs[54]);
    assign layer0_outputs[1486] = ~(inputs[206]);
    assign layer0_outputs[1487] = ~((inputs[172]) | (inputs[179]));
    assign layer0_outputs[1488] = ~(inputs[230]);
    assign layer0_outputs[1489] = ~(inputs[59]) | (inputs[250]);
    assign layer0_outputs[1490] = (inputs[106]) | (inputs[12]);
    assign layer0_outputs[1491] = ~(inputs[26]);
    assign layer0_outputs[1492] = 1'b1;
    assign layer0_outputs[1493] = inputs[148];
    assign layer0_outputs[1494] = ~(inputs[188]) | (inputs[223]);
    assign layer0_outputs[1495] = ~(inputs[240]);
    assign layer0_outputs[1496] = ~(inputs[63]);
    assign layer0_outputs[1497] = (inputs[236]) & ~(inputs[228]);
    assign layer0_outputs[1498] = ~((inputs[182]) | (inputs[36]));
    assign layer0_outputs[1499] = (inputs[155]) & ~(inputs[141]);
    assign layer0_outputs[1500] = ~((inputs[82]) | (inputs[72]));
    assign layer0_outputs[1501] = ~(inputs[244]) | (inputs[238]);
    assign layer0_outputs[1502] = (inputs[22]) | (inputs[185]);
    assign layer0_outputs[1503] = (inputs[228]) & ~(inputs[101]);
    assign layer0_outputs[1504] = (inputs[180]) & ~(inputs[79]);
    assign layer0_outputs[1505] = ~((inputs[180]) | (inputs[49]));
    assign layer0_outputs[1506] = ~((inputs[50]) & (inputs[47]));
    assign layer0_outputs[1507] = ~(inputs[143]) | (inputs[171]);
    assign layer0_outputs[1508] = 1'b0;
    assign layer0_outputs[1509] = (inputs[249]) & (inputs[59]);
    assign layer0_outputs[1510] = (inputs[69]) & ~(inputs[178]);
    assign layer0_outputs[1511] = (inputs[58]) | (inputs[118]);
    assign layer0_outputs[1512] = ~((inputs[2]) ^ (inputs[237]));
    assign layer0_outputs[1513] = ~((inputs[64]) & (inputs[234]));
    assign layer0_outputs[1514] = ~(inputs[102]) | (inputs[17]);
    assign layer0_outputs[1515] = ~(inputs[61]);
    assign layer0_outputs[1516] = inputs[37];
    assign layer0_outputs[1517] = inputs[135];
    assign layer0_outputs[1518] = (inputs[160]) ^ (inputs[180]);
    assign layer0_outputs[1519] = inputs[216];
    assign layer0_outputs[1520] = inputs[151];
    assign layer0_outputs[1521] = ~((inputs[1]) ^ (inputs[59]));
    assign layer0_outputs[1522] = (inputs[253]) & (inputs[11]);
    assign layer0_outputs[1523] = (inputs[31]) & (inputs[216]);
    assign layer0_outputs[1524] = (inputs[87]) | (inputs[89]);
    assign layer0_outputs[1525] = ~((inputs[147]) | (inputs[162]));
    assign layer0_outputs[1526] = inputs[59];
    assign layer0_outputs[1527] = (inputs[116]) ^ (inputs[169]);
    assign layer0_outputs[1528] = ~(inputs[246]) | (inputs[138]);
    assign layer0_outputs[1529] = inputs[99];
    assign layer0_outputs[1530] = ~((inputs[21]) & (inputs[155]));
    assign layer0_outputs[1531] = inputs[230];
    assign layer0_outputs[1532] = (inputs[54]) | (inputs[29]);
    assign layer0_outputs[1533] = (inputs[182]) & ~(inputs[252]);
    assign layer0_outputs[1534] = ~((inputs[55]) ^ (inputs[9]));
    assign layer0_outputs[1535] = ~((inputs[184]) ^ (inputs[239]));
    assign layer0_outputs[1536] = inputs[165];
    assign layer0_outputs[1537] = (inputs[210]) | (inputs[80]);
    assign layer0_outputs[1538] = ~(inputs[38]);
    assign layer0_outputs[1539] = (inputs[234]) | (inputs[1]);
    assign layer0_outputs[1540] = (inputs[25]) | (inputs[34]);
    assign layer0_outputs[1541] = ~((inputs[161]) | (inputs[207]));
    assign layer0_outputs[1542] = inputs[9];
    assign layer0_outputs[1543] = ~(inputs[134]) | (inputs[133]);
    assign layer0_outputs[1544] = ~(inputs[107]) | (inputs[25]);
    assign layer0_outputs[1545] = ~(inputs[148]) | (inputs[93]);
    assign layer0_outputs[1546] = ~(inputs[166]);
    assign layer0_outputs[1547] = 1'b1;
    assign layer0_outputs[1548] = inputs[151];
    assign layer0_outputs[1549] = 1'b1;
    assign layer0_outputs[1550] = ~(inputs[203]);
    assign layer0_outputs[1551] = (inputs[12]) | (inputs[128]);
    assign layer0_outputs[1552] = inputs[179];
    assign layer0_outputs[1553] = ~((inputs[198]) & (inputs[186]));
    assign layer0_outputs[1554] = ~(inputs[68]);
    assign layer0_outputs[1555] = inputs[43];
    assign layer0_outputs[1556] = ~(inputs[81]);
    assign layer0_outputs[1557] = inputs[213];
    assign layer0_outputs[1558] = inputs[220];
    assign layer0_outputs[1559] = inputs[239];
    assign layer0_outputs[1560] = ~((inputs[17]) | (inputs[43]));
    assign layer0_outputs[1561] = ~((inputs[83]) | (inputs[52]));
    assign layer0_outputs[1562] = ~(inputs[100]);
    assign layer0_outputs[1563] = ~((inputs[241]) ^ (inputs[119]));
    assign layer0_outputs[1564] = ~(inputs[32]) | (inputs[121]);
    assign layer0_outputs[1565] = ~(inputs[157]);
    assign layer0_outputs[1566] = (inputs[115]) | (inputs[157]);
    assign layer0_outputs[1567] = ~(inputs[102]) | (inputs[223]);
    assign layer0_outputs[1568] = ~(inputs[74]);
    assign layer0_outputs[1569] = ~(inputs[254]);
    assign layer0_outputs[1570] = ~(inputs[233]);
    assign layer0_outputs[1571] = ~((inputs[233]) & (inputs[26]));
    assign layer0_outputs[1572] = inputs[200];
    assign layer0_outputs[1573] = (inputs[238]) & ~(inputs[3]);
    assign layer0_outputs[1574] = inputs[23];
    assign layer0_outputs[1575] = (inputs[14]) & ~(inputs[26]);
    assign layer0_outputs[1576] = ~(inputs[107]) | (inputs[192]);
    assign layer0_outputs[1577] = inputs[26];
    assign layer0_outputs[1578] = (inputs[190]) | (inputs[243]);
    assign layer0_outputs[1579] = ~((inputs[1]) | (inputs[54]));
    assign layer0_outputs[1580] = ~((inputs[197]) & (inputs[90]));
    assign layer0_outputs[1581] = ~((inputs[219]) ^ (inputs[52]));
    assign layer0_outputs[1582] = inputs[25];
    assign layer0_outputs[1583] = inputs[7];
    assign layer0_outputs[1584] = ~((inputs[86]) ^ (inputs[164]));
    assign layer0_outputs[1585] = inputs[92];
    assign layer0_outputs[1586] = (inputs[221]) | (inputs[228]);
    assign layer0_outputs[1587] = ~(inputs[135]);
    assign layer0_outputs[1588] = inputs[120];
    assign layer0_outputs[1589] = (inputs[203]) | (inputs[118]);
    assign layer0_outputs[1590] = 1'b0;
    assign layer0_outputs[1591] = inputs[150];
    assign layer0_outputs[1592] = ~((inputs[228]) | (inputs[233]));
    assign layer0_outputs[1593] = (inputs[7]) & ~(inputs[224]);
    assign layer0_outputs[1594] = ~(inputs[18]);
    assign layer0_outputs[1595] = 1'b1;
    assign layer0_outputs[1596] = inputs[252];
    assign layer0_outputs[1597] = ~((inputs[181]) | (inputs[180]));
    assign layer0_outputs[1598] = ~((inputs[165]) | (inputs[142]));
    assign layer0_outputs[1599] = inputs[103];
    assign layer0_outputs[1600] = 1'b1;
    assign layer0_outputs[1601] = 1'b0;
    assign layer0_outputs[1602] = inputs[200];
    assign layer0_outputs[1603] = (inputs[203]) | (inputs[115]);
    assign layer0_outputs[1604] = ~((inputs[189]) ^ (inputs[143]));
    assign layer0_outputs[1605] = ~(inputs[165]) | (inputs[140]);
    assign layer0_outputs[1606] = inputs[232];
    assign layer0_outputs[1607] = ~((inputs[198]) ^ (inputs[58]));
    assign layer0_outputs[1608] = inputs[126];
    assign layer0_outputs[1609] = (inputs[209]) ^ (inputs[32]);
    assign layer0_outputs[1610] = (inputs[171]) ^ (inputs[253]);
    assign layer0_outputs[1611] = (inputs[205]) ^ (inputs[186]);
    assign layer0_outputs[1612] = inputs[121];
    assign layer0_outputs[1613] = ~(inputs[76]) | (inputs[156]);
    assign layer0_outputs[1614] = (inputs[225]) | (inputs[62]);
    assign layer0_outputs[1615] = 1'b1;
    assign layer0_outputs[1616] = inputs[70];
    assign layer0_outputs[1617] = (inputs[112]) & ~(inputs[218]);
    assign layer0_outputs[1618] = ~(inputs[38]);
    assign layer0_outputs[1619] = (inputs[233]) | (inputs[114]);
    assign layer0_outputs[1620] = (inputs[211]) & ~(inputs[28]);
    assign layer0_outputs[1621] = ~(inputs[198]) | (inputs[94]);
    assign layer0_outputs[1622] = inputs[131];
    assign layer0_outputs[1623] = ~(inputs[219]);
    assign layer0_outputs[1624] = ~((inputs[245]) | (inputs[237]));
    assign layer0_outputs[1625] = ~((inputs[149]) | (inputs[70]));
    assign layer0_outputs[1626] = inputs[190];
    assign layer0_outputs[1627] = inputs[181];
    assign layer0_outputs[1628] = (inputs[227]) | (inputs[48]);
    assign layer0_outputs[1629] = (inputs[116]) ^ (inputs[118]);
    assign layer0_outputs[1630] = ~(inputs[93]) | (inputs[216]);
    assign layer0_outputs[1631] = inputs[133];
    assign layer0_outputs[1632] = (inputs[44]) | (inputs[129]);
    assign layer0_outputs[1633] = ~(inputs[118]) | (inputs[175]);
    assign layer0_outputs[1634] = ~(inputs[102]) | (inputs[218]);
    assign layer0_outputs[1635] = inputs[88];
    assign layer0_outputs[1636] = ~(inputs[102]) | (inputs[74]);
    assign layer0_outputs[1637] = (inputs[6]) | (inputs[129]);
    assign layer0_outputs[1638] = (inputs[214]) | (inputs[230]);
    assign layer0_outputs[1639] = (inputs[216]) & ~(inputs[138]);
    assign layer0_outputs[1640] = (inputs[205]) | (inputs[254]);
    assign layer0_outputs[1641] = (inputs[180]) & (inputs[66]);
    assign layer0_outputs[1642] = ~(inputs[164]);
    assign layer0_outputs[1643] = (inputs[52]) & ~(inputs[202]);
    assign layer0_outputs[1644] = ~(inputs[137]);
    assign layer0_outputs[1645] = (inputs[50]) | (inputs[249]);
    assign layer0_outputs[1646] = (inputs[233]) & ~(inputs[79]);
    assign layer0_outputs[1647] = (inputs[184]) ^ (inputs[146]);
    assign layer0_outputs[1648] = inputs[24];
    assign layer0_outputs[1649] = ~(inputs[132]);
    assign layer0_outputs[1650] = (inputs[78]) & ~(inputs[150]);
    assign layer0_outputs[1651] = ~((inputs[191]) | (inputs[207]));
    assign layer0_outputs[1652] = inputs[201];
    assign layer0_outputs[1653] = (inputs[108]) & ~(inputs[205]);
    assign layer0_outputs[1654] = (inputs[247]) & ~(inputs[113]);
    assign layer0_outputs[1655] = ~(inputs[164]);
    assign layer0_outputs[1656] = ~((inputs[228]) | (inputs[93]));
    assign layer0_outputs[1657] = ~(inputs[69]) | (inputs[93]);
    assign layer0_outputs[1658] = ~((inputs[169]) ^ (inputs[150]));
    assign layer0_outputs[1659] = inputs[18];
    assign layer0_outputs[1660] = (inputs[53]) & ~(inputs[15]);
    assign layer0_outputs[1661] = (inputs[164]) | (inputs[62]);
    assign layer0_outputs[1662] = inputs[91];
    assign layer0_outputs[1663] = ~((inputs[177]) | (inputs[139]));
    assign layer0_outputs[1664] = (inputs[1]) ^ (inputs[21]);
    assign layer0_outputs[1665] = (inputs[77]) ^ (inputs[228]);
    assign layer0_outputs[1666] = (inputs[148]) & (inputs[197]);
    assign layer0_outputs[1667] = ~(inputs[251]);
    assign layer0_outputs[1668] = ~(inputs[70]);
    assign layer0_outputs[1669] = ~((inputs[191]) | (inputs[25]));
    assign layer0_outputs[1670] = 1'b0;
    assign layer0_outputs[1671] = ~((inputs[76]) | (inputs[208]));
    assign layer0_outputs[1672] = ~(inputs[186]) | (inputs[82]);
    assign layer0_outputs[1673] = (inputs[157]) & ~(inputs[66]);
    assign layer0_outputs[1674] = (inputs[200]) & ~(inputs[222]);
    assign layer0_outputs[1675] = ~(inputs[101]) | (inputs[49]);
    assign layer0_outputs[1676] = (inputs[133]) | (inputs[66]);
    assign layer0_outputs[1677] = inputs[78];
    assign layer0_outputs[1678] = ~(inputs[141]);
    assign layer0_outputs[1679] = ~((inputs[58]) ^ (inputs[89]));
    assign layer0_outputs[1680] = (inputs[69]) ^ (inputs[173]);
    assign layer0_outputs[1681] = inputs[246];
    assign layer0_outputs[1682] = ~(inputs[193]) | (inputs[1]);
    assign layer0_outputs[1683] = ~(inputs[70]);
    assign layer0_outputs[1684] = (inputs[108]) | (inputs[23]);
    assign layer0_outputs[1685] = (inputs[96]) ^ (inputs[10]);
    assign layer0_outputs[1686] = ~(inputs[33]);
    assign layer0_outputs[1687] = inputs[56];
    assign layer0_outputs[1688] = (inputs[80]) | (inputs[196]);
    assign layer0_outputs[1689] = (inputs[169]) ^ (inputs[110]);
    assign layer0_outputs[1690] = ~(inputs[248]) | (inputs[2]);
    assign layer0_outputs[1691] = ~(inputs[134]) | (inputs[121]);
    assign layer0_outputs[1692] = (inputs[230]) & ~(inputs[50]);
    assign layer0_outputs[1693] = (inputs[108]) & ~(inputs[226]);
    assign layer0_outputs[1694] = (inputs[77]) & ~(inputs[241]);
    assign layer0_outputs[1695] = ~(inputs[16]);
    assign layer0_outputs[1696] = ~(inputs[172]);
    assign layer0_outputs[1697] = inputs[154];
    assign layer0_outputs[1698] = ~((inputs[208]) & (inputs[234]));
    assign layer0_outputs[1699] = ~((inputs[97]) | (inputs[68]));
    assign layer0_outputs[1700] = inputs[157];
    assign layer0_outputs[1701] = (inputs[192]) | (inputs[155]);
    assign layer0_outputs[1702] = ~((inputs[85]) ^ (inputs[170]));
    assign layer0_outputs[1703] = ~(inputs[151]) | (inputs[132]);
    assign layer0_outputs[1704] = (inputs[191]) & ~(inputs[31]);
    assign layer0_outputs[1705] = (inputs[110]) & ~(inputs[223]);
    assign layer0_outputs[1706] = ~(inputs[150]) | (inputs[112]);
    assign layer0_outputs[1707] = (inputs[196]) ^ (inputs[104]);
    assign layer0_outputs[1708] = ~(inputs[11]) | (inputs[223]);
    assign layer0_outputs[1709] = ~(inputs[26]) | (inputs[182]);
    assign layer0_outputs[1710] = inputs[161];
    assign layer0_outputs[1711] = (inputs[7]) & ~(inputs[163]);
    assign layer0_outputs[1712] = inputs[142];
    assign layer0_outputs[1713] = inputs[115];
    assign layer0_outputs[1714] = ~((inputs[239]) | (inputs[239]));
    assign layer0_outputs[1715] = ~((inputs[39]) | (inputs[29]));
    assign layer0_outputs[1716] = ~((inputs[251]) | (inputs[200]));
    assign layer0_outputs[1717] = inputs[192];
    assign layer0_outputs[1718] = ~(inputs[20]) | (inputs[128]);
    assign layer0_outputs[1719] = inputs[41];
    assign layer0_outputs[1720] = ~(inputs[92]);
    assign layer0_outputs[1721] = inputs[237];
    assign layer0_outputs[1722] = ~(inputs[219]);
    assign layer0_outputs[1723] = 1'b1;
    assign layer0_outputs[1724] = (inputs[33]) ^ (inputs[138]);
    assign layer0_outputs[1725] = 1'b0;
    assign layer0_outputs[1726] = (inputs[27]) & ~(inputs[210]);
    assign layer0_outputs[1727] = ~(inputs[28]) | (inputs[223]);
    assign layer0_outputs[1728] = inputs[152];
    assign layer0_outputs[1729] = ~(inputs[53]) | (inputs[85]);
    assign layer0_outputs[1730] = (inputs[20]) | (inputs[79]);
    assign layer0_outputs[1731] = ~(inputs[78]);
    assign layer0_outputs[1732] = (inputs[14]) ^ (inputs[72]);
    assign layer0_outputs[1733] = (inputs[70]) | (inputs[61]);
    assign layer0_outputs[1734] = (inputs[199]) | (inputs[65]);
    assign layer0_outputs[1735] = ~(inputs[144]);
    assign layer0_outputs[1736] = ~(inputs[4]);
    assign layer0_outputs[1737] = (inputs[108]) & ~(inputs[207]);
    assign layer0_outputs[1738] = ~((inputs[152]) & (inputs[203]));
    assign layer0_outputs[1739] = ~(inputs[142]) | (inputs[229]);
    assign layer0_outputs[1740] = ~(inputs[111]);
    assign layer0_outputs[1741] = (inputs[40]) & ~(inputs[178]);
    assign layer0_outputs[1742] = ~((inputs[96]) ^ (inputs[68]));
    assign layer0_outputs[1743] = ~(inputs[248]) | (inputs[73]);
    assign layer0_outputs[1744] = ~((inputs[50]) | (inputs[9]));
    assign layer0_outputs[1745] = ~(inputs[61]) | (inputs[27]);
    assign layer0_outputs[1746] = 1'b0;
    assign layer0_outputs[1747] = ~((inputs[115]) ^ (inputs[178]));
    assign layer0_outputs[1748] = ~(inputs[191]) | (inputs[251]);
    assign layer0_outputs[1749] = (inputs[191]) | (inputs[31]);
    assign layer0_outputs[1750] = ~(inputs[54]) | (inputs[13]);
    assign layer0_outputs[1751] = (inputs[71]) & ~(inputs[220]);
    assign layer0_outputs[1752] = ~(inputs[231]) | (inputs[53]);
    assign layer0_outputs[1753] = ~((inputs[153]) | (inputs[248]));
    assign layer0_outputs[1754] = (inputs[92]) ^ (inputs[129]);
    assign layer0_outputs[1755] = ~((inputs[152]) ^ (inputs[121]));
    assign layer0_outputs[1756] = inputs[147];
    assign layer0_outputs[1757] = ~(inputs[40]);
    assign layer0_outputs[1758] = (inputs[218]) & (inputs[94]);
    assign layer0_outputs[1759] = inputs[23];
    assign layer0_outputs[1760] = inputs[203];
    assign layer0_outputs[1761] = ~(inputs[229]);
    assign layer0_outputs[1762] = ~((inputs[89]) ^ (inputs[38]));
    assign layer0_outputs[1763] = ~(inputs[231]);
    assign layer0_outputs[1764] = ~(inputs[226]) | (inputs[220]);
    assign layer0_outputs[1765] = (inputs[70]) | (inputs[147]);
    assign layer0_outputs[1766] = ~(inputs[163]) | (inputs[214]);
    assign layer0_outputs[1767] = ~(inputs[87]) | (inputs[24]);
    assign layer0_outputs[1768] = (inputs[94]) | (inputs[8]);
    assign layer0_outputs[1769] = ~(inputs[147]) | (inputs[239]);
    assign layer0_outputs[1770] = ~(inputs[30]);
    assign layer0_outputs[1771] = inputs[180];
    assign layer0_outputs[1772] = (inputs[149]) | (inputs[198]);
    assign layer0_outputs[1773] = inputs[118];
    assign layer0_outputs[1774] = ~((inputs[192]) | (inputs[234]));
    assign layer0_outputs[1775] = (inputs[117]) & ~(inputs[65]);
    assign layer0_outputs[1776] = ~((inputs[3]) ^ (inputs[33]));
    assign layer0_outputs[1777] = ~(inputs[113]) | (inputs[233]);
    assign layer0_outputs[1778] = ~(inputs[16]);
    assign layer0_outputs[1779] = (inputs[183]) & ~(inputs[130]);
    assign layer0_outputs[1780] = ~((inputs[213]) | (inputs[127]));
    assign layer0_outputs[1781] = ~((inputs[151]) & (inputs[231]));
    assign layer0_outputs[1782] = (inputs[8]) & (inputs[73]);
    assign layer0_outputs[1783] = ~((inputs[187]) | (inputs[172]));
    assign layer0_outputs[1784] = ~(inputs[113]) | (inputs[134]);
    assign layer0_outputs[1785] = ~((inputs[0]) | (inputs[8]));
    assign layer0_outputs[1786] = ~(inputs[80]) | (inputs[144]);
    assign layer0_outputs[1787] = ~(inputs[60]) | (inputs[32]);
    assign layer0_outputs[1788] = ~(inputs[56]);
    assign layer0_outputs[1789] = ~(inputs[199]);
    assign layer0_outputs[1790] = (inputs[138]) | (inputs[91]);
    assign layer0_outputs[1791] = 1'b0;
    assign layer0_outputs[1792] = (inputs[94]) | (inputs[60]);
    assign layer0_outputs[1793] = (inputs[97]) ^ (inputs[240]);
    assign layer0_outputs[1794] = (inputs[244]) | (inputs[190]);
    assign layer0_outputs[1795] = ~((inputs[237]) ^ (inputs[173]));
    assign layer0_outputs[1796] = (inputs[75]) & ~(inputs[193]);
    assign layer0_outputs[1797] = (inputs[118]) | (inputs[19]);
    assign layer0_outputs[1798] = (inputs[77]) | (inputs[30]);
    assign layer0_outputs[1799] = (inputs[83]) & (inputs[67]);
    assign layer0_outputs[1800] = ~(inputs[247]);
    assign layer0_outputs[1801] = inputs[240];
    assign layer0_outputs[1802] = ~(inputs[176]) | (inputs[194]);
    assign layer0_outputs[1803] = inputs[236];
    assign layer0_outputs[1804] = ~(inputs[61]);
    assign layer0_outputs[1805] = inputs[42];
    assign layer0_outputs[1806] = (inputs[43]) ^ (inputs[58]);
    assign layer0_outputs[1807] = (inputs[57]) | (inputs[247]);
    assign layer0_outputs[1808] = ~(inputs[85]);
    assign layer0_outputs[1809] = ~(inputs[30]) | (inputs[86]);
    assign layer0_outputs[1810] = (inputs[183]) & ~(inputs[129]);
    assign layer0_outputs[1811] = ~((inputs[213]) & (inputs[173]));
    assign layer0_outputs[1812] = ~((inputs[208]) ^ (inputs[4]));
    assign layer0_outputs[1813] = ~(inputs[19]);
    assign layer0_outputs[1814] = (inputs[212]) & ~(inputs[90]);
    assign layer0_outputs[1815] = ~((inputs[71]) | (inputs[17]));
    assign layer0_outputs[1816] = ~(inputs[168]) | (inputs[63]);
    assign layer0_outputs[1817] = ~(inputs[172]) | (inputs[154]);
    assign layer0_outputs[1818] = ~((inputs[120]) | (inputs[241]));
    assign layer0_outputs[1819] = ~(inputs[69]) | (inputs[121]);
    assign layer0_outputs[1820] = 1'b1;
    assign layer0_outputs[1821] = inputs[206];
    assign layer0_outputs[1822] = (inputs[162]) ^ (inputs[113]);
    assign layer0_outputs[1823] = ~(inputs[210]);
    assign layer0_outputs[1824] = ~(inputs[189]) | (inputs[10]);
    assign layer0_outputs[1825] = ~((inputs[172]) | (inputs[112]));
    assign layer0_outputs[1826] = (inputs[110]) | (inputs[181]);
    assign layer0_outputs[1827] = ~((inputs[179]) | (inputs[111]));
    assign layer0_outputs[1828] = ~((inputs[131]) ^ (inputs[112]));
    assign layer0_outputs[1829] = ~((inputs[73]) | (inputs[187]));
    assign layer0_outputs[1830] = ~(inputs[28]);
    assign layer0_outputs[1831] = inputs[94];
    assign layer0_outputs[1832] = ~(inputs[231]) | (inputs[252]);
    assign layer0_outputs[1833] = (inputs[130]) | (inputs[133]);
    assign layer0_outputs[1834] = ~((inputs[16]) | (inputs[160]));
    assign layer0_outputs[1835] = ~((inputs[94]) ^ (inputs[25]));
    assign layer0_outputs[1836] = (inputs[134]) & ~(inputs[15]);
    assign layer0_outputs[1837] = ~((inputs[161]) ^ (inputs[88]));
    assign layer0_outputs[1838] = inputs[252];
    assign layer0_outputs[1839] = (inputs[88]) & ~(inputs[28]);
    assign layer0_outputs[1840] = ~((inputs[156]) | (inputs[93]));
    assign layer0_outputs[1841] = ~(inputs[116]);
    assign layer0_outputs[1842] = ~((inputs[103]) | (inputs[67]));
    assign layer0_outputs[1843] = (inputs[48]) & ~(inputs[31]);
    assign layer0_outputs[1844] = ~(inputs[233]);
    assign layer0_outputs[1845] = (inputs[19]) | (inputs[218]);
    assign layer0_outputs[1846] = ~(inputs[70]) | (inputs[50]);
    assign layer0_outputs[1847] = (inputs[193]) | (inputs[105]);
    assign layer0_outputs[1848] = ~(inputs[41]) | (inputs[170]);
    assign layer0_outputs[1849] = inputs[177];
    assign layer0_outputs[1850] = (inputs[12]) & ~(inputs[208]);
    assign layer0_outputs[1851] = inputs[155];
    assign layer0_outputs[1852] = ~(inputs[209]);
    assign layer0_outputs[1853] = inputs[126];
    assign layer0_outputs[1854] = ~(inputs[249]);
    assign layer0_outputs[1855] = (inputs[100]) & ~(inputs[142]);
    assign layer0_outputs[1856] = (inputs[161]) | (inputs[227]);
    assign layer0_outputs[1857] = ~(inputs[251]) | (inputs[48]);
    assign layer0_outputs[1858] = ~((inputs[90]) ^ (inputs[119]));
    assign layer0_outputs[1859] = ~(inputs[16]);
    assign layer0_outputs[1860] = (inputs[245]) | (inputs[141]);
    assign layer0_outputs[1861] = ~(inputs[77]);
    assign layer0_outputs[1862] = ~(inputs[37]);
    assign layer0_outputs[1863] = (inputs[239]) ^ (inputs[206]);
    assign layer0_outputs[1864] = inputs[236];
    assign layer0_outputs[1865] = (inputs[237]) & ~(inputs[74]);
    assign layer0_outputs[1866] = ~(inputs[197]) | (inputs[68]);
    assign layer0_outputs[1867] = (inputs[131]) | (inputs[65]);
    assign layer0_outputs[1868] = ~((inputs[187]) | (inputs[37]));
    assign layer0_outputs[1869] = inputs[245];
    assign layer0_outputs[1870] = (inputs[16]) | (inputs[191]);
    assign layer0_outputs[1871] = (inputs[43]) | (inputs[22]);
    assign layer0_outputs[1872] = ~((inputs[149]) | (inputs[229]));
    assign layer0_outputs[1873] = (inputs[228]) & ~(inputs[252]);
    assign layer0_outputs[1874] = (inputs[212]) | (inputs[187]);
    assign layer0_outputs[1875] = (inputs[210]) | (inputs[216]);
    assign layer0_outputs[1876] = ~((inputs[133]) ^ (inputs[152]));
    assign layer0_outputs[1877] = (inputs[193]) & (inputs[193]);
    assign layer0_outputs[1878] = (inputs[139]) ^ (inputs[164]);
    assign layer0_outputs[1879] = inputs[123];
    assign layer0_outputs[1880] = ~((inputs[175]) ^ (inputs[189]));
    assign layer0_outputs[1881] = ~((inputs[183]) & (inputs[252]));
    assign layer0_outputs[1882] = ~(inputs[74]) | (inputs[156]);
    assign layer0_outputs[1883] = (inputs[24]) & ~(inputs[129]);
    assign layer0_outputs[1884] = ~(inputs[67]);
    assign layer0_outputs[1885] = (inputs[78]) & ~(inputs[173]);
    assign layer0_outputs[1886] = ~(inputs[48]);
    assign layer0_outputs[1887] = (inputs[8]) & ~(inputs[164]);
    assign layer0_outputs[1888] = (inputs[86]) ^ (inputs[177]);
    assign layer0_outputs[1889] = (inputs[205]) & ~(inputs[21]);
    assign layer0_outputs[1890] = (inputs[161]) & ~(inputs[150]);
    assign layer0_outputs[1891] = (inputs[107]) & ~(inputs[193]);
    assign layer0_outputs[1892] = ~((inputs[219]) | (inputs[206]));
    assign layer0_outputs[1893] = ~(inputs[117]) | (inputs[92]);
    assign layer0_outputs[1894] = ~(inputs[178]) | (inputs[17]);
    assign layer0_outputs[1895] = ~(inputs[245]);
    assign layer0_outputs[1896] = inputs[97];
    assign layer0_outputs[1897] = ~(inputs[128]);
    assign layer0_outputs[1898] = (inputs[151]) | (inputs[55]);
    assign layer0_outputs[1899] = inputs[147];
    assign layer0_outputs[1900] = (inputs[103]) | (inputs[77]);
    assign layer0_outputs[1901] = (inputs[157]) | (inputs[79]);
    assign layer0_outputs[1902] = (inputs[60]) | (inputs[77]);
    assign layer0_outputs[1903] = ~(inputs[150]);
    assign layer0_outputs[1904] = ~(inputs[252]) | (inputs[252]);
    assign layer0_outputs[1905] = (inputs[21]) | (inputs[121]);
    assign layer0_outputs[1906] = ~(inputs[100]);
    assign layer0_outputs[1907] = (inputs[237]) & ~(inputs[74]);
    assign layer0_outputs[1908] = ~(inputs[8]) | (inputs[15]);
    assign layer0_outputs[1909] = ~(inputs[165]);
    assign layer0_outputs[1910] = (inputs[173]) ^ (inputs[215]);
    assign layer0_outputs[1911] = inputs[37];
    assign layer0_outputs[1912] = (inputs[41]) ^ (inputs[9]);
    assign layer0_outputs[1913] = (inputs[165]) | (inputs[148]);
    assign layer0_outputs[1914] = ~((inputs[37]) ^ (inputs[82]));
    assign layer0_outputs[1915] = ~(inputs[178]);
    assign layer0_outputs[1916] = ~(inputs[193]);
    assign layer0_outputs[1917] = ~(inputs[164]);
    assign layer0_outputs[1918] = ~(inputs[119]) | (inputs[163]);
    assign layer0_outputs[1919] = ~((inputs[49]) | (inputs[192]));
    assign layer0_outputs[1920] = ~(inputs[199]) | (inputs[217]);
    assign layer0_outputs[1921] = (inputs[152]) & ~(inputs[26]);
    assign layer0_outputs[1922] = (inputs[84]) | (inputs[156]);
    assign layer0_outputs[1923] = ~(inputs[47]);
    assign layer0_outputs[1924] = (inputs[208]) | (inputs[192]);
    assign layer0_outputs[1925] = (inputs[205]) & ~(inputs[32]);
    assign layer0_outputs[1926] = ~(inputs[25]);
    assign layer0_outputs[1927] = ~(inputs[51]) | (inputs[168]);
    assign layer0_outputs[1928] = (inputs[161]) | (inputs[178]);
    assign layer0_outputs[1929] = (inputs[208]) | (inputs[5]);
    assign layer0_outputs[1930] = (inputs[128]) ^ (inputs[33]);
    assign layer0_outputs[1931] = ~(inputs[3]);
    assign layer0_outputs[1932] = ~(inputs[115]) | (inputs[17]);
    assign layer0_outputs[1933] = ~((inputs[120]) | (inputs[96]));
    assign layer0_outputs[1934] = (inputs[147]) | (inputs[115]);
    assign layer0_outputs[1935] = ~(inputs[45]) | (inputs[41]);
    assign layer0_outputs[1936] = (inputs[76]) ^ (inputs[235]);
    assign layer0_outputs[1937] = ~(inputs[163]) | (inputs[167]);
    assign layer0_outputs[1938] = (inputs[198]) & ~(inputs[93]);
    assign layer0_outputs[1939] = inputs[141];
    assign layer0_outputs[1940] = ~(inputs[34]) | (inputs[66]);
    assign layer0_outputs[1941] = ~(inputs[135]);
    assign layer0_outputs[1942] = (inputs[106]) ^ (inputs[180]);
    assign layer0_outputs[1943] = ~(inputs[88]) | (inputs[225]);
    assign layer0_outputs[1944] = (inputs[155]) & ~(inputs[110]);
    assign layer0_outputs[1945] = ~(inputs[71]);
    assign layer0_outputs[1946] = (inputs[229]) | (inputs[208]);
    assign layer0_outputs[1947] = ~(inputs[211]) | (inputs[22]);
    assign layer0_outputs[1948] = (inputs[84]) ^ (inputs[21]);
    assign layer0_outputs[1949] = ~((inputs[147]) | (inputs[156]));
    assign layer0_outputs[1950] = (inputs[208]) & ~(inputs[0]);
    assign layer0_outputs[1951] = ~((inputs[169]) | (inputs[150]));
    assign layer0_outputs[1952] = ~(inputs[228]);
    assign layer0_outputs[1953] = ~(inputs[67]);
    assign layer0_outputs[1954] = 1'b1;
    assign layer0_outputs[1955] = ~(inputs[67]);
    assign layer0_outputs[1956] = inputs[123];
    assign layer0_outputs[1957] = ~(inputs[41]) | (inputs[111]);
    assign layer0_outputs[1958] = (inputs[6]) | (inputs[227]);
    assign layer0_outputs[1959] = inputs[4];
    assign layer0_outputs[1960] = inputs[220];
    assign layer0_outputs[1961] = inputs[92];
    assign layer0_outputs[1962] = inputs[171];
    assign layer0_outputs[1963] = (inputs[236]) | (inputs[55]);
    assign layer0_outputs[1964] = inputs[255];
    assign layer0_outputs[1965] = (inputs[118]) | (inputs[251]);
    assign layer0_outputs[1966] = inputs[148];
    assign layer0_outputs[1967] = ~((inputs[112]) | (inputs[247]));
    assign layer0_outputs[1968] = ~(inputs[27]);
    assign layer0_outputs[1969] = ~(inputs[244]) | (inputs[203]);
    assign layer0_outputs[1970] = (inputs[34]) | (inputs[69]);
    assign layer0_outputs[1971] = ~(inputs[87]);
    assign layer0_outputs[1972] = (inputs[130]) & ~(inputs[32]);
    assign layer0_outputs[1973] = (inputs[192]) | (inputs[17]);
    assign layer0_outputs[1974] = (inputs[103]) & ~(inputs[109]);
    assign layer0_outputs[1975] = ~(inputs[106]);
    assign layer0_outputs[1976] = ~((inputs[243]) & (inputs[16]));
    assign layer0_outputs[1977] = (inputs[55]) ^ (inputs[10]);
    assign layer0_outputs[1978] = inputs[141];
    assign layer0_outputs[1979] = (inputs[242]) & ~(inputs[66]);
    assign layer0_outputs[1980] = ~((inputs[146]) | (inputs[179]));
    assign layer0_outputs[1981] = ~((inputs[115]) | (inputs[101]));
    assign layer0_outputs[1982] = ~(inputs[134]) | (inputs[144]);
    assign layer0_outputs[1983] = ~(inputs[82]);
    assign layer0_outputs[1984] = ~(inputs[97]);
    assign layer0_outputs[1985] = ~(inputs[237]);
    assign layer0_outputs[1986] = (inputs[122]) & ~(inputs[81]);
    assign layer0_outputs[1987] = ~(inputs[149]) | (inputs[206]);
    assign layer0_outputs[1988] = 1'b1;
    assign layer0_outputs[1989] = ~(inputs[193]);
    assign layer0_outputs[1990] = ~(inputs[108]) | (inputs[39]);
    assign layer0_outputs[1991] = (inputs[179]) | (inputs[111]);
    assign layer0_outputs[1992] = 1'b0;
    assign layer0_outputs[1993] = ~(inputs[183]) | (inputs[112]);
    assign layer0_outputs[1994] = (inputs[231]) | (inputs[176]);
    assign layer0_outputs[1995] = ~(inputs[104]);
    assign layer0_outputs[1996] = 1'b0;
    assign layer0_outputs[1997] = (inputs[7]) | (inputs[75]);
    assign layer0_outputs[1998] = (inputs[171]) & (inputs[224]);
    assign layer0_outputs[1999] = (inputs[20]) | (inputs[70]);
    assign layer0_outputs[2000] = (inputs[67]) & ~(inputs[65]);
    assign layer0_outputs[2001] = ~((inputs[184]) | (inputs[127]));
    assign layer0_outputs[2002] = ~((inputs[183]) | (inputs[55]));
    assign layer0_outputs[2003] = ~((inputs[180]) ^ (inputs[177]));
    assign layer0_outputs[2004] = ~((inputs[244]) | (inputs[95]));
    assign layer0_outputs[2005] = 1'b0;
    assign layer0_outputs[2006] = 1'b1;
    assign layer0_outputs[2007] = ~((inputs[118]) & (inputs[51]));
    assign layer0_outputs[2008] = ~(inputs[66]) | (inputs[142]);
    assign layer0_outputs[2009] = 1'b0;
    assign layer0_outputs[2010] = (inputs[117]) | (inputs[221]);
    assign layer0_outputs[2011] = ~(inputs[117]) | (inputs[121]);
    assign layer0_outputs[2012] = (inputs[28]) | (inputs[244]);
    assign layer0_outputs[2013] = (inputs[146]) | (inputs[219]);
    assign layer0_outputs[2014] = (inputs[32]) & ~(inputs[79]);
    assign layer0_outputs[2015] = (inputs[242]) | (inputs[194]);
    assign layer0_outputs[2016] = (inputs[9]) ^ (inputs[57]);
    assign layer0_outputs[2017] = ~(inputs[16]);
    assign layer0_outputs[2018] = (inputs[208]) & ~(inputs[200]);
    assign layer0_outputs[2019] = ~(inputs[170]);
    assign layer0_outputs[2020] = (inputs[17]) ^ (inputs[171]);
    assign layer0_outputs[2021] = inputs[14];
    assign layer0_outputs[2022] = ~(inputs[230]);
    assign layer0_outputs[2023] = ~(inputs[167]);
    assign layer0_outputs[2024] = (inputs[56]) | (inputs[228]);
    assign layer0_outputs[2025] = (inputs[31]) | (inputs[43]);
    assign layer0_outputs[2026] = ~((inputs[89]) | (inputs[99]));
    assign layer0_outputs[2027] = (inputs[139]) & ~(inputs[224]);
    assign layer0_outputs[2028] = ~(inputs[239]);
    assign layer0_outputs[2029] = ~((inputs[35]) ^ (inputs[220]));
    assign layer0_outputs[2030] = ~(inputs[35]);
    assign layer0_outputs[2031] = ~((inputs[0]) ^ (inputs[221]));
    assign layer0_outputs[2032] = ~(inputs[25]);
    assign layer0_outputs[2033] = (inputs[171]) & (inputs[245]);
    assign layer0_outputs[2034] = ~(inputs[130]);
    assign layer0_outputs[2035] = ~(inputs[26]);
    assign layer0_outputs[2036] = inputs[168];
    assign layer0_outputs[2037] = (inputs[237]) | (inputs[149]);
    assign layer0_outputs[2038] = ~(inputs[153]);
    assign layer0_outputs[2039] = (inputs[162]) | (inputs[176]);
    assign layer0_outputs[2040] = inputs[254];
    assign layer0_outputs[2041] = ~(inputs[67]);
    assign layer0_outputs[2042] = (inputs[132]) ^ (inputs[149]);
    assign layer0_outputs[2043] = ~(inputs[46]);
    assign layer0_outputs[2044] = ~((inputs[85]) & (inputs[62]));
    assign layer0_outputs[2045] = ~(inputs[228]) | (inputs[53]);
    assign layer0_outputs[2046] = inputs[7];
    assign layer0_outputs[2047] = ~((inputs[146]) | (inputs[175]));
    assign layer0_outputs[2048] = 1'b0;
    assign layer0_outputs[2049] = (inputs[131]) ^ (inputs[21]);
    assign layer0_outputs[2050] = ~(inputs[164]);
    assign layer0_outputs[2051] = ~(inputs[197]);
    assign layer0_outputs[2052] = inputs[178];
    assign layer0_outputs[2053] = (inputs[189]) & ~(inputs[12]);
    assign layer0_outputs[2054] = ~(inputs[255]) | (inputs[122]);
    assign layer0_outputs[2055] = ~((inputs[248]) | (inputs[42]));
    assign layer0_outputs[2056] = ~(inputs[91]);
    assign layer0_outputs[2057] = inputs[93];
    assign layer0_outputs[2058] = ~((inputs[178]) ^ (inputs[232]));
    assign layer0_outputs[2059] = ~(inputs[159]) | (inputs[64]);
    assign layer0_outputs[2060] = inputs[121];
    assign layer0_outputs[2061] = ~(inputs[117]);
    assign layer0_outputs[2062] = inputs[67];
    assign layer0_outputs[2063] = ~(inputs[117]);
    assign layer0_outputs[2064] = ~((inputs[227]) & (inputs[247]));
    assign layer0_outputs[2065] = ~((inputs[214]) ^ (inputs[199]));
    assign layer0_outputs[2066] = (inputs[86]) & ~(inputs[150]);
    assign layer0_outputs[2067] = ~((inputs[65]) | (inputs[164]));
    assign layer0_outputs[2068] = ~(inputs[160]) | (inputs[255]);
    assign layer0_outputs[2069] = ~((inputs[181]) ^ (inputs[208]));
    assign layer0_outputs[2070] = ~(inputs[126]);
    assign layer0_outputs[2071] = ~(inputs[57]);
    assign layer0_outputs[2072] = (inputs[204]) & ~(inputs[41]);
    assign layer0_outputs[2073] = (inputs[128]) & (inputs[210]);
    assign layer0_outputs[2074] = ~((inputs[130]) ^ (inputs[147]));
    assign layer0_outputs[2075] = ~((inputs[203]) ^ (inputs[97]));
    assign layer0_outputs[2076] = (inputs[199]) | (inputs[184]);
    assign layer0_outputs[2077] = 1'b0;
    assign layer0_outputs[2078] = ~((inputs[247]) | (inputs[18]));
    assign layer0_outputs[2079] = ~(inputs[82]) | (inputs[24]);
    assign layer0_outputs[2080] = (inputs[232]) ^ (inputs[113]);
    assign layer0_outputs[2081] = ~((inputs[3]) | (inputs[186]));
    assign layer0_outputs[2082] = ~(inputs[3]) | (inputs[112]);
    assign layer0_outputs[2083] = inputs[81];
    assign layer0_outputs[2084] = (inputs[152]) & ~(inputs[9]);
    assign layer0_outputs[2085] = ~((inputs[254]) | (inputs[253]));
    assign layer0_outputs[2086] = ~(inputs[186]) | (inputs[5]);
    assign layer0_outputs[2087] = ~(inputs[167]) | (inputs[190]);
    assign layer0_outputs[2088] = (inputs[208]) ^ (inputs[212]);
    assign layer0_outputs[2089] = ~(inputs[213]) | (inputs[30]);
    assign layer0_outputs[2090] = inputs[208];
    assign layer0_outputs[2091] = ~(inputs[167]) | (inputs[143]);
    assign layer0_outputs[2092] = inputs[114];
    assign layer0_outputs[2093] = (inputs[23]) | (inputs[124]);
    assign layer0_outputs[2094] = ~(inputs[193]) | (inputs[11]);
    assign layer0_outputs[2095] = 1'b1;
    assign layer0_outputs[2096] = ~((inputs[77]) | (inputs[109]));
    assign layer0_outputs[2097] = ~((inputs[240]) ^ (inputs[154]));
    assign layer0_outputs[2098] = 1'b1;
    assign layer0_outputs[2099] = (inputs[205]) & ~(inputs[112]);
    assign layer0_outputs[2100] = (inputs[28]) ^ (inputs[103]);
    assign layer0_outputs[2101] = ~(inputs[34]) | (inputs[202]);
    assign layer0_outputs[2102] = ~(inputs[41]) | (inputs[224]);
    assign layer0_outputs[2103] = ~((inputs[99]) & (inputs[121]));
    assign layer0_outputs[2104] = inputs[65];
    assign layer0_outputs[2105] = 1'b0;
    assign layer0_outputs[2106] = (inputs[45]) & ~(inputs[241]);
    assign layer0_outputs[2107] = inputs[81];
    assign layer0_outputs[2108] = (inputs[122]) & ~(inputs[97]);
    assign layer0_outputs[2109] = ~(inputs[74]);
    assign layer0_outputs[2110] = (inputs[172]) | (inputs[226]);
    assign layer0_outputs[2111] = (inputs[240]) & ~(inputs[191]);
    assign layer0_outputs[2112] = ~(inputs[222]) | (inputs[114]);
    assign layer0_outputs[2113] = (inputs[243]) | (inputs[208]);
    assign layer0_outputs[2114] = ~((inputs[207]) ^ (inputs[236]));
    assign layer0_outputs[2115] = ~((inputs[91]) | (inputs[236]));
    assign layer0_outputs[2116] = ~((inputs[212]) ^ (inputs[234]));
    assign layer0_outputs[2117] = ~(inputs[7]);
    assign layer0_outputs[2118] = ~(inputs[83]) | (inputs[96]);
    assign layer0_outputs[2119] = ~(inputs[139]);
    assign layer0_outputs[2120] = ~(inputs[108]) | (inputs[223]);
    assign layer0_outputs[2121] = (inputs[127]) & ~(inputs[11]);
    assign layer0_outputs[2122] = ~((inputs[246]) & (inputs[80]));
    assign layer0_outputs[2123] = inputs[182];
    assign layer0_outputs[2124] = ~(inputs[227]) | (inputs[82]);
    assign layer0_outputs[2125] = ~((inputs[225]) | (inputs[152]));
    assign layer0_outputs[2126] = ~((inputs[117]) | (inputs[113]));
    assign layer0_outputs[2127] = ~(inputs[218]) | (inputs[31]);
    assign layer0_outputs[2128] = ~((inputs[3]) | (inputs[96]));
    assign layer0_outputs[2129] = inputs[113];
    assign layer0_outputs[2130] = inputs[72];
    assign layer0_outputs[2131] = 1'b1;
    assign layer0_outputs[2132] = inputs[212];
    assign layer0_outputs[2133] = 1'b1;
    assign layer0_outputs[2134] = ~(inputs[123]);
    assign layer0_outputs[2135] = (inputs[196]) & ~(inputs[76]);
    assign layer0_outputs[2136] = ~((inputs[211]) | (inputs[87]));
    assign layer0_outputs[2137] = inputs[212];
    assign layer0_outputs[2138] = ~(inputs[20]);
    assign layer0_outputs[2139] = ~(inputs[216]) | (inputs[246]);
    assign layer0_outputs[2140] = (inputs[250]) | (inputs[189]);
    assign layer0_outputs[2141] = ~((inputs[139]) ^ (inputs[164]));
    assign layer0_outputs[2142] = (inputs[9]) & ~(inputs[63]);
    assign layer0_outputs[2143] = ~((inputs[196]) | (inputs[112]));
    assign layer0_outputs[2144] = (inputs[46]) & ~(inputs[145]);
    assign layer0_outputs[2145] = ~(inputs[23]);
    assign layer0_outputs[2146] = (inputs[74]) & (inputs[13]);
    assign layer0_outputs[2147] = ~((inputs[30]) & (inputs[123]));
    assign layer0_outputs[2148] = ~((inputs[57]) & (inputs[3]));
    assign layer0_outputs[2149] = (inputs[199]) & ~(inputs[255]);
    assign layer0_outputs[2150] = ~(inputs[198]) | (inputs[16]);
    assign layer0_outputs[2151] = (inputs[160]) & ~(inputs[147]);
    assign layer0_outputs[2152] = ~(inputs[73]);
    assign layer0_outputs[2153] = ~(inputs[182]);
    assign layer0_outputs[2154] = (inputs[205]) ^ (inputs[21]);
    assign layer0_outputs[2155] = (inputs[216]) | (inputs[246]);
    assign layer0_outputs[2156] = ~(inputs[162]);
    assign layer0_outputs[2157] = (inputs[201]) | (inputs[227]);
    assign layer0_outputs[2158] = inputs[234];
    assign layer0_outputs[2159] = ~(inputs[21]) | (inputs[228]);
    assign layer0_outputs[2160] = (inputs[253]) & ~(inputs[187]);
    assign layer0_outputs[2161] = ~((inputs[74]) | (inputs[167]));
    assign layer0_outputs[2162] = ~(inputs[229]) | (inputs[103]);
    assign layer0_outputs[2163] = ~((inputs[15]) | (inputs[4]));
    assign layer0_outputs[2164] = ~((inputs[109]) ^ (inputs[41]));
    assign layer0_outputs[2165] = ~(inputs[48]);
    assign layer0_outputs[2166] = (inputs[80]) | (inputs[9]);
    assign layer0_outputs[2167] = (inputs[194]) | (inputs[249]);
    assign layer0_outputs[2168] = (inputs[104]) & ~(inputs[190]);
    assign layer0_outputs[2169] = (inputs[159]) ^ (inputs[106]);
    assign layer0_outputs[2170] = ~((inputs[107]) & (inputs[37]));
    assign layer0_outputs[2171] = (inputs[236]) | (inputs[173]);
    assign layer0_outputs[2172] = (inputs[166]) & ~(inputs[214]);
    assign layer0_outputs[2173] = (inputs[36]) ^ (inputs[97]);
    assign layer0_outputs[2174] = (inputs[236]) ^ (inputs[10]);
    assign layer0_outputs[2175] = (inputs[89]) ^ (inputs[106]);
    assign layer0_outputs[2176] = inputs[60];
    assign layer0_outputs[2177] = ~(inputs[65]);
    assign layer0_outputs[2178] = ~((inputs[230]) | (inputs[176]));
    assign layer0_outputs[2179] = inputs[232];
    assign layer0_outputs[2180] = inputs[164];
    assign layer0_outputs[2181] = (inputs[229]) & ~(inputs[37]);
    assign layer0_outputs[2182] = (inputs[135]) & ~(inputs[62]);
    assign layer0_outputs[2183] = ~((inputs[69]) ^ (inputs[226]));
    assign layer0_outputs[2184] = inputs[151];
    assign layer0_outputs[2185] = ~((inputs[148]) ^ (inputs[155]));
    assign layer0_outputs[2186] = ~(inputs[86]);
    assign layer0_outputs[2187] = inputs[149];
    assign layer0_outputs[2188] = (inputs[12]) | (inputs[227]);
    assign layer0_outputs[2189] = inputs[27];
    assign layer0_outputs[2190] = ~((inputs[32]) | (inputs[208]));
    assign layer0_outputs[2191] = (inputs[116]) & ~(inputs[0]);
    assign layer0_outputs[2192] = ~(inputs[92]) | (inputs[180]);
    assign layer0_outputs[2193] = (inputs[234]) & ~(inputs[150]);
    assign layer0_outputs[2194] = ~((inputs[117]) ^ (inputs[239]));
    assign layer0_outputs[2195] = (inputs[192]) & ~(inputs[0]);
    assign layer0_outputs[2196] = ~((inputs[175]) | (inputs[158]));
    assign layer0_outputs[2197] = ~((inputs[133]) ^ (inputs[177]));
    assign layer0_outputs[2198] = (inputs[217]) ^ (inputs[163]);
    assign layer0_outputs[2199] = inputs[199];
    assign layer0_outputs[2200] = (inputs[198]) & ~(inputs[208]);
    assign layer0_outputs[2201] = ~((inputs[60]) ^ (inputs[43]));
    assign layer0_outputs[2202] = (inputs[162]) | (inputs[176]);
    assign layer0_outputs[2203] = ~((inputs[155]) | (inputs[52]));
    assign layer0_outputs[2204] = inputs[159];
    assign layer0_outputs[2205] = ~((inputs[190]) | (inputs[150]));
    assign layer0_outputs[2206] = (inputs[220]) & ~(inputs[243]);
    assign layer0_outputs[2207] = (inputs[83]) ^ (inputs[84]);
    assign layer0_outputs[2208] = inputs[234];
    assign layer0_outputs[2209] = ~(inputs[85]);
    assign layer0_outputs[2210] = (inputs[127]) & ~(inputs[251]);
    assign layer0_outputs[2211] = (inputs[130]) & ~(inputs[39]);
    assign layer0_outputs[2212] = inputs[101];
    assign layer0_outputs[2213] = ~((inputs[77]) | (inputs[176]));
    assign layer0_outputs[2214] = ~(inputs[184]);
    assign layer0_outputs[2215] = (inputs[185]) ^ (inputs[80]);
    assign layer0_outputs[2216] = ~(inputs[91]) | (inputs[40]);
    assign layer0_outputs[2217] = inputs[141];
    assign layer0_outputs[2218] = ~(inputs[161]);
    assign layer0_outputs[2219] = inputs[117];
    assign layer0_outputs[2220] = (inputs[64]) ^ (inputs[5]);
    assign layer0_outputs[2221] = ~(inputs[139]);
    assign layer0_outputs[2222] = (inputs[177]) ^ (inputs[136]);
    assign layer0_outputs[2223] = ~((inputs[230]) ^ (inputs[190]));
    assign layer0_outputs[2224] = inputs[127];
    assign layer0_outputs[2225] = ~((inputs[81]) | (inputs[124]));
    assign layer0_outputs[2226] = ~((inputs[0]) | (inputs[30]));
    assign layer0_outputs[2227] = 1'b0;
    assign layer0_outputs[2228] = ~(inputs[19]);
    assign layer0_outputs[2229] = (inputs[88]) & ~(inputs[85]);
    assign layer0_outputs[2230] = inputs[164];
    assign layer0_outputs[2231] = (inputs[56]) & ~(inputs[197]);
    assign layer0_outputs[2232] = (inputs[13]) & (inputs[243]);
    assign layer0_outputs[2233] = ~(inputs[48]);
    assign layer0_outputs[2234] = ~((inputs[198]) | (inputs[47]));
    assign layer0_outputs[2235] = ~(inputs[211]) | (inputs[108]);
    assign layer0_outputs[2236] = (inputs[111]) | (inputs[165]);
    assign layer0_outputs[2237] = inputs[16];
    assign layer0_outputs[2238] = ~((inputs[122]) ^ (inputs[93]));
    assign layer0_outputs[2239] = (inputs[42]) | (inputs[241]);
    assign layer0_outputs[2240] = (inputs[64]) & ~(inputs[173]);
    assign layer0_outputs[2241] = 1'b0;
    assign layer0_outputs[2242] = inputs[220];
    assign layer0_outputs[2243] = ~(inputs[74]);
    assign layer0_outputs[2244] = ~(inputs[10]);
    assign layer0_outputs[2245] = (inputs[213]) ^ (inputs[200]);
    assign layer0_outputs[2246] = ~(inputs[240]) | (inputs[50]);
    assign layer0_outputs[2247] = (inputs[116]) & ~(inputs[4]);
    assign layer0_outputs[2248] = ~(inputs[231]) | (inputs[237]);
    assign layer0_outputs[2249] = (inputs[31]) ^ (inputs[166]);
    assign layer0_outputs[2250] = ~(inputs[140]) | (inputs[61]);
    assign layer0_outputs[2251] = inputs[114];
    assign layer0_outputs[2252] = (inputs[228]) | (inputs[251]);
    assign layer0_outputs[2253] = (inputs[214]) & ~(inputs[15]);
    assign layer0_outputs[2254] = ~(inputs[94]);
    assign layer0_outputs[2255] = (inputs[77]) ^ (inputs[228]);
    assign layer0_outputs[2256] = inputs[66];
    assign layer0_outputs[2257] = (inputs[86]) & ~(inputs[160]);
    assign layer0_outputs[2258] = inputs[175];
    assign layer0_outputs[2259] = (inputs[47]) | (inputs[15]);
    assign layer0_outputs[2260] = (inputs[179]) & ~(inputs[34]);
    assign layer0_outputs[2261] = ~(inputs[109]) | (inputs[154]);
    assign layer0_outputs[2262] = inputs[247];
    assign layer0_outputs[2263] = (inputs[107]) & ~(inputs[205]);
    assign layer0_outputs[2264] = ~((inputs[145]) ^ (inputs[143]));
    assign layer0_outputs[2265] = inputs[157];
    assign layer0_outputs[2266] = ~(inputs[214]);
    assign layer0_outputs[2267] = ~(inputs[163]);
    assign layer0_outputs[2268] = ~(inputs[164]);
    assign layer0_outputs[2269] = ~(inputs[188]);
    assign layer0_outputs[2270] = ~((inputs[194]) | (inputs[31]));
    assign layer0_outputs[2271] = ~(inputs[150]) | (inputs[155]);
    assign layer0_outputs[2272] = ~(inputs[206]) | (inputs[39]);
    assign layer0_outputs[2273] = 1'b1;
    assign layer0_outputs[2274] = inputs[22];
    assign layer0_outputs[2275] = (inputs[145]) ^ (inputs[204]);
    assign layer0_outputs[2276] = ~((inputs[230]) & (inputs[124]));
    assign layer0_outputs[2277] = ~(inputs[56]) | (inputs[247]);
    assign layer0_outputs[2278] = (inputs[1]) ^ (inputs[226]);
    assign layer0_outputs[2279] = (inputs[74]) | (inputs[106]);
    assign layer0_outputs[2280] = (inputs[195]) & ~(inputs[79]);
    assign layer0_outputs[2281] = 1'b0;
    assign layer0_outputs[2282] = inputs[248];
    assign layer0_outputs[2283] = (inputs[27]) ^ (inputs[78]);
    assign layer0_outputs[2284] = ~((inputs[41]) & (inputs[75]));
    assign layer0_outputs[2285] = ~((inputs[130]) ^ (inputs[245]));
    assign layer0_outputs[2286] = ~((inputs[238]) & (inputs[59]));
    assign layer0_outputs[2287] = ~(inputs[129]) | (inputs[181]);
    assign layer0_outputs[2288] = ~(inputs[194]);
    assign layer0_outputs[2289] = ~(inputs[129]);
    assign layer0_outputs[2290] = (inputs[2]) | (inputs[39]);
    assign layer0_outputs[2291] = ~((inputs[202]) & (inputs[242]));
    assign layer0_outputs[2292] = ~((inputs[230]) ^ (inputs[230]));
    assign layer0_outputs[2293] = ~(inputs[84]);
    assign layer0_outputs[2294] = (inputs[129]) ^ (inputs[252]);
    assign layer0_outputs[2295] = (inputs[33]) & ~(inputs[6]);
    assign layer0_outputs[2296] = ~((inputs[150]) | (inputs[82]));
    assign layer0_outputs[2297] = (inputs[116]) & ~(inputs[5]);
    assign layer0_outputs[2298] = (inputs[245]) & ~(inputs[186]);
    assign layer0_outputs[2299] = ~(inputs[180]) | (inputs[160]);
    assign layer0_outputs[2300] = inputs[98];
    assign layer0_outputs[2301] = ~(inputs[55]) | (inputs[38]);
    assign layer0_outputs[2302] = ~((inputs[162]) ^ (inputs[229]));
    assign layer0_outputs[2303] = ~(inputs[74]);
    assign layer0_outputs[2304] = (inputs[157]) & (inputs[144]);
    assign layer0_outputs[2305] = ~(inputs[23]);
    assign layer0_outputs[2306] = ~(inputs[250]) | (inputs[9]);
    assign layer0_outputs[2307] = ~(inputs[91]) | (inputs[208]);
    assign layer0_outputs[2308] = (inputs[57]) & ~(inputs[168]);
    assign layer0_outputs[2309] = ~((inputs[156]) ^ (inputs[35]));
    assign layer0_outputs[2310] = inputs[121];
    assign layer0_outputs[2311] = ~(inputs[99]);
    assign layer0_outputs[2312] = ~((inputs[95]) | (inputs[32]));
    assign layer0_outputs[2313] = 1'b0;
    assign layer0_outputs[2314] = (inputs[96]) & ~(inputs[113]);
    assign layer0_outputs[2315] = (inputs[126]) & (inputs[92]);
    assign layer0_outputs[2316] = inputs[76];
    assign layer0_outputs[2317] = ~(inputs[82]) | (inputs[171]);
    assign layer0_outputs[2318] = ~(inputs[112]) | (inputs[210]);
    assign layer0_outputs[2319] = ~(inputs[154]);
    assign layer0_outputs[2320] = 1'b1;
    assign layer0_outputs[2321] = (inputs[25]) & ~(inputs[155]);
    assign layer0_outputs[2322] = (inputs[137]) | (inputs[170]);
    assign layer0_outputs[2323] = inputs[94];
    assign layer0_outputs[2324] = ~(inputs[30]) | (inputs[10]);
    assign layer0_outputs[2325] = ~(inputs[83]);
    assign layer0_outputs[2326] = ~((inputs[41]) | (inputs[14]));
    assign layer0_outputs[2327] = ~((inputs[107]) ^ (inputs[142]));
    assign layer0_outputs[2328] = ~(inputs[166]) | (inputs[238]);
    assign layer0_outputs[2329] = ~(inputs[1]) | (inputs[207]);
    assign layer0_outputs[2330] = inputs[182];
    assign layer0_outputs[2331] = (inputs[201]) | (inputs[6]);
    assign layer0_outputs[2332] = (inputs[50]) & (inputs[152]);
    assign layer0_outputs[2333] = ~(inputs[238]) | (inputs[87]);
    assign layer0_outputs[2334] = (inputs[227]) & ~(inputs[252]);
    assign layer0_outputs[2335] = ~(inputs[98]) | (inputs[17]);
    assign layer0_outputs[2336] = ~((inputs[146]) ^ (inputs[87]));
    assign layer0_outputs[2337] = ~(inputs[68]);
    assign layer0_outputs[2338] = ~(inputs[213]) | (inputs[146]);
    assign layer0_outputs[2339] = ~(inputs[135]);
    assign layer0_outputs[2340] = (inputs[75]) ^ (inputs[47]);
    assign layer0_outputs[2341] = (inputs[180]) | (inputs[106]);
    assign layer0_outputs[2342] = (inputs[126]) & ~(inputs[19]);
    assign layer0_outputs[2343] = (inputs[71]) | (inputs[71]);
    assign layer0_outputs[2344] = (inputs[64]) & ~(inputs[206]);
    assign layer0_outputs[2345] = (inputs[23]) & ~(inputs[32]);
    assign layer0_outputs[2346] = (inputs[230]) & ~(inputs[152]);
    assign layer0_outputs[2347] = ~(inputs[181]);
    assign layer0_outputs[2348] = (inputs[162]) ^ (inputs[249]);
    assign layer0_outputs[2349] = (inputs[176]) | (inputs[1]);
    assign layer0_outputs[2350] = ~(inputs[91]) | (inputs[158]);
    assign layer0_outputs[2351] = ~(inputs[10]);
    assign layer0_outputs[2352] = ~((inputs[177]) ^ (inputs[20]));
    assign layer0_outputs[2353] = ~((inputs[81]) | (inputs[39]));
    assign layer0_outputs[2354] = ~((inputs[231]) | (inputs[132]));
    assign layer0_outputs[2355] = 1'b0;
    assign layer0_outputs[2356] = (inputs[197]) & ~(inputs[124]);
    assign layer0_outputs[2357] = ~((inputs[137]) | (inputs[63]));
    assign layer0_outputs[2358] = ~(inputs[101]);
    assign layer0_outputs[2359] = ~(inputs[72]);
    assign layer0_outputs[2360] = 1'b1;
    assign layer0_outputs[2361] = (inputs[199]) ^ (inputs[1]);
    assign layer0_outputs[2362] = (inputs[147]) & ~(inputs[93]);
    assign layer0_outputs[2363] = (inputs[83]) ^ (inputs[190]);
    assign layer0_outputs[2364] = ~((inputs[96]) | (inputs[151]));
    assign layer0_outputs[2365] = (inputs[38]) & (inputs[122]);
    assign layer0_outputs[2366] = (inputs[77]) & (inputs[232]);
    assign layer0_outputs[2367] = (inputs[38]) & ~(inputs[70]);
    assign layer0_outputs[2368] = ~(inputs[182]) | (inputs[127]);
    assign layer0_outputs[2369] = ~(inputs[42]);
    assign layer0_outputs[2370] = (inputs[174]) | (inputs[169]);
    assign layer0_outputs[2371] = ~(inputs[99]);
    assign layer0_outputs[2372] = ~(inputs[204]) | (inputs[14]);
    assign layer0_outputs[2373] = (inputs[91]) & (inputs[247]);
    assign layer0_outputs[2374] = (inputs[120]) & ~(inputs[16]);
    assign layer0_outputs[2375] = ~((inputs[97]) ^ (inputs[228]));
    assign layer0_outputs[2376] = (inputs[139]) ^ (inputs[61]);
    assign layer0_outputs[2377] = ~((inputs[254]) | (inputs[46]));
    assign layer0_outputs[2378] = ~((inputs[225]) ^ (inputs[162]));
    assign layer0_outputs[2379] = ~(inputs[77]) | (inputs[235]);
    assign layer0_outputs[2380] = ~((inputs[32]) | (inputs[52]));
    assign layer0_outputs[2381] = ~((inputs[80]) ^ (inputs[84]));
    assign layer0_outputs[2382] = ~(inputs[146]);
    assign layer0_outputs[2383] = ~(inputs[189]);
    assign layer0_outputs[2384] = ~((inputs[81]) | (inputs[211]));
    assign layer0_outputs[2385] = (inputs[8]) & ~(inputs[42]);
    assign layer0_outputs[2386] = inputs[244];
    assign layer0_outputs[2387] = 1'b0;
    assign layer0_outputs[2388] = 1'b1;
    assign layer0_outputs[2389] = (inputs[81]) & (inputs[158]);
    assign layer0_outputs[2390] = ~((inputs[160]) | (inputs[147]));
    assign layer0_outputs[2391] = ~(inputs[41]);
    assign layer0_outputs[2392] = (inputs[76]) | (inputs[101]);
    assign layer0_outputs[2393] = inputs[106];
    assign layer0_outputs[2394] = (inputs[49]) & ~(inputs[15]);
    assign layer0_outputs[2395] = (inputs[52]) ^ (inputs[80]);
    assign layer0_outputs[2396] = 1'b1;
    assign layer0_outputs[2397] = 1'b1;
    assign layer0_outputs[2398] = inputs[32];
    assign layer0_outputs[2399] = ~((inputs[171]) ^ (inputs[218]));
    assign layer0_outputs[2400] = ~(inputs[55]);
    assign layer0_outputs[2401] = inputs[54];
    assign layer0_outputs[2402] = (inputs[135]) | (inputs[122]);
    assign layer0_outputs[2403] = 1'b1;
    assign layer0_outputs[2404] = ~((inputs[248]) ^ (inputs[208]));
    assign layer0_outputs[2405] = ~(inputs[39]);
    assign layer0_outputs[2406] = inputs[168];
    assign layer0_outputs[2407] = ~(inputs[48]);
    assign layer0_outputs[2408] = ~(inputs[84]);
    assign layer0_outputs[2409] = (inputs[119]) & (inputs[159]);
    assign layer0_outputs[2410] = ~((inputs[132]) | (inputs[249]));
    assign layer0_outputs[2411] = ~(inputs[70]) | (inputs[60]);
    assign layer0_outputs[2412] = inputs[63];
    assign layer0_outputs[2413] = ~((inputs[128]) | (inputs[75]));
    assign layer0_outputs[2414] = ~((inputs[8]) & (inputs[222]));
    assign layer0_outputs[2415] = ~((inputs[140]) ^ (inputs[142]));
    assign layer0_outputs[2416] = ~(inputs[106]) | (inputs[185]);
    assign layer0_outputs[2417] = inputs[153];
    assign layer0_outputs[2418] = (inputs[194]) & ~(inputs[11]);
    assign layer0_outputs[2419] = (inputs[110]) ^ (inputs[49]);
    assign layer0_outputs[2420] = ~(inputs[55]);
    assign layer0_outputs[2421] = (inputs[49]) | (inputs[216]);
    assign layer0_outputs[2422] = (inputs[213]) | (inputs[141]);
    assign layer0_outputs[2423] = ~(inputs[100]);
    assign layer0_outputs[2424] = ~(inputs[196]);
    assign layer0_outputs[2425] = ~(inputs[101]) | (inputs[33]);
    assign layer0_outputs[2426] = (inputs[24]) & ~(inputs[135]);
    assign layer0_outputs[2427] = ~(inputs[94]);
    assign layer0_outputs[2428] = 1'b1;
    assign layer0_outputs[2429] = (inputs[40]) ^ (inputs[24]);
    assign layer0_outputs[2430] = ~(inputs[165]);
    assign layer0_outputs[2431] = ~((inputs[59]) ^ (inputs[223]));
    assign layer0_outputs[2432] = ~(inputs[49]);
    assign layer0_outputs[2433] = inputs[140];
    assign layer0_outputs[2434] = (inputs[224]) & ~(inputs[112]);
    assign layer0_outputs[2435] = ~((inputs[41]) ^ (inputs[215]));
    assign layer0_outputs[2436] = (inputs[96]) ^ (inputs[247]);
    assign layer0_outputs[2437] = inputs[235];
    assign layer0_outputs[2438] = inputs[21];
    assign layer0_outputs[2439] = inputs[76];
    assign layer0_outputs[2440] = ~((inputs[186]) ^ (inputs[174]));
    assign layer0_outputs[2441] = ~(inputs[69]);
    assign layer0_outputs[2442] = ~((inputs[78]) | (inputs[40]));
    assign layer0_outputs[2443] = ~((inputs[112]) | (inputs[125]));
    assign layer0_outputs[2444] = ~((inputs[51]) | (inputs[237]));
    assign layer0_outputs[2445] = ~((inputs[233]) & (inputs[77]));
    assign layer0_outputs[2446] = ~(inputs[234]);
    assign layer0_outputs[2447] = ~(inputs[114]) | (inputs[243]);
    assign layer0_outputs[2448] = ~((inputs[170]) | (inputs[8]));
    assign layer0_outputs[2449] = 1'b1;
    assign layer0_outputs[2450] = (inputs[218]) & (inputs[159]);
    assign layer0_outputs[2451] = inputs[160];
    assign layer0_outputs[2452] = (inputs[59]) | (inputs[59]);
    assign layer0_outputs[2453] = ~(inputs[39]);
    assign layer0_outputs[2454] = ~(inputs[114]);
    assign layer0_outputs[2455] = ~((inputs[22]) | (inputs[38]));
    assign layer0_outputs[2456] = (inputs[77]) | (inputs[146]);
    assign layer0_outputs[2457] = (inputs[160]) & ~(inputs[202]);
    assign layer0_outputs[2458] = ~((inputs[171]) ^ (inputs[217]));
    assign layer0_outputs[2459] = (inputs[121]) | (inputs[180]);
    assign layer0_outputs[2460] = ~(inputs[110]);
    assign layer0_outputs[2461] = ~((inputs[87]) | (inputs[237]));
    assign layer0_outputs[2462] = (inputs[125]) ^ (inputs[208]);
    assign layer0_outputs[2463] = inputs[142];
    assign layer0_outputs[2464] = inputs[151];
    assign layer0_outputs[2465] = inputs[17];
    assign layer0_outputs[2466] = ~(inputs[59]);
    assign layer0_outputs[2467] = ~(inputs[123]) | (inputs[72]);
    assign layer0_outputs[2468] = ~(inputs[15]) | (inputs[8]);
    assign layer0_outputs[2469] = (inputs[197]) & ~(inputs[97]);
    assign layer0_outputs[2470] = ~(inputs[74]);
    assign layer0_outputs[2471] = (inputs[30]) & ~(inputs[85]);
    assign layer0_outputs[2472] = (inputs[96]) | (inputs[114]);
    assign layer0_outputs[2473] = (inputs[69]) & ~(inputs[224]);
    assign layer0_outputs[2474] = ~(inputs[116]);
    assign layer0_outputs[2475] = (inputs[157]) & (inputs[58]);
    assign layer0_outputs[2476] = ~(inputs[116]) | (inputs[201]);
    assign layer0_outputs[2477] = 1'b1;
    assign layer0_outputs[2478] = ~((inputs[12]) | (inputs[19]));
    assign layer0_outputs[2479] = (inputs[62]) & ~(inputs[15]);
    assign layer0_outputs[2480] = (inputs[114]) ^ (inputs[137]);
    assign layer0_outputs[2481] = ~((inputs[227]) | (inputs[167]));
    assign layer0_outputs[2482] = ~(inputs[204]) | (inputs[147]);
    assign layer0_outputs[2483] = ~(inputs[53]);
    assign layer0_outputs[2484] = ~(inputs[169]) | (inputs[90]);
    assign layer0_outputs[2485] = ~(inputs[193]);
    assign layer0_outputs[2486] = ~((inputs[224]) | (inputs[145]));
    assign layer0_outputs[2487] = ~((inputs[126]) | (inputs[33]));
    assign layer0_outputs[2488] = ~(inputs[234]);
    assign layer0_outputs[2489] = ~(inputs[33]);
    assign layer0_outputs[2490] = ~(inputs[40]);
    assign layer0_outputs[2491] = (inputs[172]) & (inputs[11]);
    assign layer0_outputs[2492] = ~((inputs[221]) | (inputs[228]));
    assign layer0_outputs[2493] = ~(inputs[187]) | (inputs[253]);
    assign layer0_outputs[2494] = (inputs[165]) | (inputs[182]);
    assign layer0_outputs[2495] = 1'b0;
    assign layer0_outputs[2496] = ~(inputs[196]) | (inputs[241]);
    assign layer0_outputs[2497] = (inputs[17]) ^ (inputs[9]);
    assign layer0_outputs[2498] = ~(inputs[213]) | (inputs[35]);
    assign layer0_outputs[2499] = inputs[203];
    assign layer0_outputs[2500] = inputs[171];
    assign layer0_outputs[2501] = ~(inputs[150]) | (inputs[140]);
    assign layer0_outputs[2502] = ~((inputs[173]) | (inputs[255]));
    assign layer0_outputs[2503] = inputs[248];
    assign layer0_outputs[2504] = (inputs[72]) & ~(inputs[207]);
    assign layer0_outputs[2505] = ~((inputs[209]) | (inputs[97]));
    assign layer0_outputs[2506] = ~(inputs[181]);
    assign layer0_outputs[2507] = ~(inputs[105]) | (inputs[78]);
    assign layer0_outputs[2508] = ~((inputs[184]) | (inputs[200]));
    assign layer0_outputs[2509] = (inputs[105]) | (inputs[237]);
    assign layer0_outputs[2510] = ~(inputs[248]);
    assign layer0_outputs[2511] = ~(inputs[35]) | (inputs[221]);
    assign layer0_outputs[2512] = inputs[116];
    assign layer0_outputs[2513] = ~(inputs[149]) | (inputs[203]);
    assign layer0_outputs[2514] = ~(inputs[230]) | (inputs[239]);
    assign layer0_outputs[2515] = ~(inputs[107]);
    assign layer0_outputs[2516] = inputs[63];
    assign layer0_outputs[2517] = ~(inputs[74]);
    assign layer0_outputs[2518] = (inputs[3]) ^ (inputs[219]);
    assign layer0_outputs[2519] = ~((inputs[202]) | (inputs[246]));
    assign layer0_outputs[2520] = ~((inputs[178]) | (inputs[212]));
    assign layer0_outputs[2521] = (inputs[60]) | (inputs[79]);
    assign layer0_outputs[2522] = ~((inputs[73]) | (inputs[207]));
    assign layer0_outputs[2523] = (inputs[67]) & ~(inputs[165]);
    assign layer0_outputs[2524] = ~(inputs[14]);
    assign layer0_outputs[2525] = ~((inputs[171]) & (inputs[229]));
    assign layer0_outputs[2526] = (inputs[4]) | (inputs[175]);
    assign layer0_outputs[2527] = ~((inputs[187]) | (inputs[248]));
    assign layer0_outputs[2528] = 1'b0;
    assign layer0_outputs[2529] = (inputs[92]) | (inputs[223]);
    assign layer0_outputs[2530] = inputs[100];
    assign layer0_outputs[2531] = inputs[104];
    assign layer0_outputs[2532] = ~(inputs[137]) | (inputs[80]);
    assign layer0_outputs[2533] = (inputs[126]) & ~(inputs[75]);
    assign layer0_outputs[2534] = (inputs[15]) & (inputs[4]);
    assign layer0_outputs[2535] = inputs[180];
    assign layer0_outputs[2536] = ~((inputs[144]) | (inputs[194]));
    assign layer0_outputs[2537] = ~(inputs[24]);
    assign layer0_outputs[2538] = ~(inputs[185]);
    assign layer0_outputs[2539] = ~(inputs[233]);
    assign layer0_outputs[2540] = (inputs[59]) | (inputs[51]);
    assign layer0_outputs[2541] = ~((inputs[93]) | (inputs[4]));
    assign layer0_outputs[2542] = ~(inputs[52]);
    assign layer0_outputs[2543] = inputs[65];
    assign layer0_outputs[2544] = ~((inputs[104]) | (inputs[133]));
    assign layer0_outputs[2545] = (inputs[55]) | (inputs[198]);
    assign layer0_outputs[2546] = inputs[23];
    assign layer0_outputs[2547] = inputs[194];
    assign layer0_outputs[2548] = ~((inputs[52]) | (inputs[108]));
    assign layer0_outputs[2549] = (inputs[88]) | (inputs[216]);
    assign layer0_outputs[2550] = (inputs[196]) & ~(inputs[251]);
    assign layer0_outputs[2551] = (inputs[143]) ^ (inputs[185]);
    assign layer0_outputs[2552] = (inputs[136]) & ~(inputs[175]);
    assign layer0_outputs[2553] = ~(inputs[35]) | (inputs[5]);
    assign layer0_outputs[2554] = 1'b0;
    assign layer0_outputs[2555] = inputs[209];
    assign layer0_outputs[2556] = inputs[61];
    assign layer0_outputs[2557] = 1'b0;
    assign layer0_outputs[2558] = (inputs[184]) & ~(inputs[174]);
    assign layer0_outputs[2559] = ~(inputs[250]);
    assign layer0_outputs[2560] = (inputs[183]) ^ (inputs[126]);
    assign layer0_outputs[2561] = ~((inputs[60]) | (inputs[52]));
    assign layer0_outputs[2562] = ~(inputs[27]) | (inputs[32]);
    assign layer0_outputs[2563] = ~(inputs[53]);
    assign layer0_outputs[2564] = (inputs[9]) ^ (inputs[43]);
    assign layer0_outputs[2565] = inputs[95];
    assign layer0_outputs[2566] = (inputs[70]) ^ (inputs[201]);
    assign layer0_outputs[2567] = (inputs[71]) & ~(inputs[100]);
    assign layer0_outputs[2568] = (inputs[224]) & ~(inputs[228]);
    assign layer0_outputs[2569] = 1'b1;
    assign layer0_outputs[2570] = (inputs[76]) & ~(inputs[186]);
    assign layer0_outputs[2571] = ~(inputs[54]) | (inputs[0]);
    assign layer0_outputs[2572] = ~((inputs[231]) | (inputs[2]));
    assign layer0_outputs[2573] = inputs[113];
    assign layer0_outputs[2574] = 1'b1;
    assign layer0_outputs[2575] = ~(inputs[250]);
    assign layer0_outputs[2576] = ~(inputs[188]);
    assign layer0_outputs[2577] = ~(inputs[214]);
    assign layer0_outputs[2578] = ~((inputs[97]) | (inputs[83]));
    assign layer0_outputs[2579] = 1'b0;
    assign layer0_outputs[2580] = 1'b1;
    assign layer0_outputs[2581] = (inputs[206]) & ~(inputs[39]);
    assign layer0_outputs[2582] = (inputs[109]) | (inputs[114]);
    assign layer0_outputs[2583] = inputs[218];
    assign layer0_outputs[2584] = ~((inputs[92]) ^ (inputs[111]));
    assign layer0_outputs[2585] = (inputs[82]) & ~(inputs[16]);
    assign layer0_outputs[2586] = (inputs[132]) ^ (inputs[24]);
    assign layer0_outputs[2587] = inputs[172];
    assign layer0_outputs[2588] = ~(inputs[156]);
    assign layer0_outputs[2589] = ~(inputs[164]);
    assign layer0_outputs[2590] = ~(inputs[64]);
    assign layer0_outputs[2591] = ~((inputs[150]) ^ (inputs[89]));
    assign layer0_outputs[2592] = (inputs[29]) & ~(inputs[43]);
    assign layer0_outputs[2593] = ~(inputs[5]);
    assign layer0_outputs[2594] = ~(inputs[96]) | (inputs[249]);
    assign layer0_outputs[2595] = inputs[135];
    assign layer0_outputs[2596] = (inputs[85]) & ~(inputs[105]);
    assign layer0_outputs[2597] = (inputs[106]) ^ (inputs[237]);
    assign layer0_outputs[2598] = (inputs[61]) | (inputs[22]);
    assign layer0_outputs[2599] = ~((inputs[170]) ^ (inputs[252]));
    assign layer0_outputs[2600] = inputs[71];
    assign layer0_outputs[2601] = ~(inputs[164]) | (inputs[148]);
    assign layer0_outputs[2602] = 1'b0;
    assign layer0_outputs[2603] = ~(inputs[222]) | (inputs[234]);
    assign layer0_outputs[2604] = ~(inputs[102]);
    assign layer0_outputs[2605] = ~(inputs[148]);
    assign layer0_outputs[2606] = ~(inputs[24]);
    assign layer0_outputs[2607] = ~((inputs[183]) | (inputs[212]));
    assign layer0_outputs[2608] = (inputs[13]) & ~(inputs[115]);
    assign layer0_outputs[2609] = inputs[188];
    assign layer0_outputs[2610] = ~(inputs[115]);
    assign layer0_outputs[2611] = 1'b1;
    assign layer0_outputs[2612] = (inputs[240]) & ~(inputs[145]);
    assign layer0_outputs[2613] = 1'b1;
    assign layer0_outputs[2614] = ~(inputs[66]) | (inputs[55]);
    assign layer0_outputs[2615] = (inputs[136]) & (inputs[123]);
    assign layer0_outputs[2616] = (inputs[226]) | (inputs[193]);
    assign layer0_outputs[2617] = ~(inputs[117]);
    assign layer0_outputs[2618] = ~(inputs[158]);
    assign layer0_outputs[2619] = ~(inputs[121]) | (inputs[53]);
    assign layer0_outputs[2620] = (inputs[122]) ^ (inputs[173]);
    assign layer0_outputs[2621] = 1'b1;
    assign layer0_outputs[2622] = inputs[0];
    assign layer0_outputs[2623] = inputs[176];
    assign layer0_outputs[2624] = ~(inputs[90]);
    assign layer0_outputs[2625] = inputs[152];
    assign layer0_outputs[2626] = ~((inputs[85]) | (inputs[139]));
    assign layer0_outputs[2627] = ~(inputs[253]);
    assign layer0_outputs[2628] = (inputs[80]) | (inputs[4]);
    assign layer0_outputs[2629] = inputs[47];
    assign layer0_outputs[2630] = (inputs[64]) ^ (inputs[147]);
    assign layer0_outputs[2631] = (inputs[57]) ^ (inputs[95]);
    assign layer0_outputs[2632] = (inputs[141]) & ~(inputs[11]);
    assign layer0_outputs[2633] = 1'b0;
    assign layer0_outputs[2634] = inputs[146];
    assign layer0_outputs[2635] = (inputs[12]) ^ (inputs[119]);
    assign layer0_outputs[2636] = inputs[87];
    assign layer0_outputs[2637] = (inputs[55]) & ~(inputs[107]);
    assign layer0_outputs[2638] = ~(inputs[217]);
    assign layer0_outputs[2639] = ~((inputs[146]) ^ (inputs[181]));
    assign layer0_outputs[2640] = inputs[26];
    assign layer0_outputs[2641] = 1'b0;
    assign layer0_outputs[2642] = 1'b0;
    assign layer0_outputs[2643] = ~((inputs[89]) | (inputs[151]));
    assign layer0_outputs[2644] = (inputs[125]) ^ (inputs[123]);
    assign layer0_outputs[2645] = ~((inputs[151]) ^ (inputs[140]));
    assign layer0_outputs[2646] = (inputs[148]) ^ (inputs[102]);
    assign layer0_outputs[2647] = (inputs[208]) | (inputs[222]);
    assign layer0_outputs[2648] = (inputs[81]) | (inputs[248]);
    assign layer0_outputs[2649] = ~((inputs[93]) & (inputs[217]));
    assign layer0_outputs[2650] = (inputs[50]) & ~(inputs[239]);
    assign layer0_outputs[2651] = (inputs[214]) | (inputs[78]);
    assign layer0_outputs[2652] = (inputs[171]) | (inputs[188]);
    assign layer0_outputs[2653] = (inputs[101]) & (inputs[76]);
    assign layer0_outputs[2654] = inputs[214];
    assign layer0_outputs[2655] = (inputs[167]) | (inputs[80]);
    assign layer0_outputs[2656] = ~(inputs[252]) | (inputs[84]);
    assign layer0_outputs[2657] = ~((inputs[78]) | (inputs[208]));
    assign layer0_outputs[2658] = ~((inputs[202]) | (inputs[38]));
    assign layer0_outputs[2659] = ~(inputs[56]);
    assign layer0_outputs[2660] = 1'b0;
    assign layer0_outputs[2661] = inputs[71];
    assign layer0_outputs[2662] = ~(inputs[157]);
    assign layer0_outputs[2663] = ~(inputs[108]) | (inputs[56]);
    assign layer0_outputs[2664] = ~(inputs[219]);
    assign layer0_outputs[2665] = inputs[111];
    assign layer0_outputs[2666] = ~((inputs[218]) | (inputs[217]));
    assign layer0_outputs[2667] = ~(inputs[116]);
    assign layer0_outputs[2668] = (inputs[39]) & ~(inputs[169]);
    assign layer0_outputs[2669] = ~(inputs[147]) | (inputs[248]);
    assign layer0_outputs[2670] = (inputs[53]) & ~(inputs[34]);
    assign layer0_outputs[2671] = ~(inputs[152]);
    assign layer0_outputs[2672] = ~(inputs[163]);
    assign layer0_outputs[2673] = ~(inputs[104]) | (inputs[123]);
    assign layer0_outputs[2674] = (inputs[189]) & ~(inputs[15]);
    assign layer0_outputs[2675] = ~(inputs[123]);
    assign layer0_outputs[2676] = (inputs[76]) & ~(inputs[81]);
    assign layer0_outputs[2677] = ~(inputs[208]);
    assign layer0_outputs[2678] = inputs[64];
    assign layer0_outputs[2679] = inputs[8];
    assign layer0_outputs[2680] = inputs[145];
    assign layer0_outputs[2681] = (inputs[84]) | (inputs[246]);
    assign layer0_outputs[2682] = inputs[22];
    assign layer0_outputs[2683] = (inputs[250]) | (inputs[102]);
    assign layer0_outputs[2684] = 1'b1;
    assign layer0_outputs[2685] = ~(inputs[186]);
    assign layer0_outputs[2686] = inputs[75];
    assign layer0_outputs[2687] = ~((inputs[93]) | (inputs[221]));
    assign layer0_outputs[2688] = ~((inputs[33]) | (inputs[34]));
    assign layer0_outputs[2689] = inputs[77];
    assign layer0_outputs[2690] = (inputs[188]) | (inputs[203]);
    assign layer0_outputs[2691] = (inputs[43]) & ~(inputs[181]);
    assign layer0_outputs[2692] = ~((inputs[120]) & (inputs[115]));
    assign layer0_outputs[2693] = (inputs[195]) | (inputs[15]);
    assign layer0_outputs[2694] = ~(inputs[247]) | (inputs[37]);
    assign layer0_outputs[2695] = ~(inputs[229]) | (inputs[234]);
    assign layer0_outputs[2696] = (inputs[107]) & ~(inputs[197]);
    assign layer0_outputs[2697] = ~((inputs[60]) | (inputs[238]));
    assign layer0_outputs[2698] = inputs[182];
    assign layer0_outputs[2699] = ~(inputs[85]) | (inputs[249]);
    assign layer0_outputs[2700] = inputs[124];
    assign layer0_outputs[2701] = (inputs[116]) | (inputs[60]);
    assign layer0_outputs[2702] = (inputs[220]) & ~(inputs[94]);
    assign layer0_outputs[2703] = 1'b1;
    assign layer0_outputs[2704] = ~((inputs[130]) | (inputs[16]));
    assign layer0_outputs[2705] = (inputs[170]) & ~(inputs[209]);
    assign layer0_outputs[2706] = (inputs[149]) & ~(inputs[13]);
    assign layer0_outputs[2707] = ~(inputs[66]);
    assign layer0_outputs[2708] = (inputs[29]) ^ (inputs[248]);
    assign layer0_outputs[2709] = (inputs[124]) & ~(inputs[222]);
    assign layer0_outputs[2710] = ~(inputs[222]);
    assign layer0_outputs[2711] = 1'b1;
    assign layer0_outputs[2712] = ~(inputs[1]);
    assign layer0_outputs[2713] = (inputs[38]) | (inputs[240]);
    assign layer0_outputs[2714] = ~((inputs[56]) | (inputs[71]));
    assign layer0_outputs[2715] = ~(inputs[22]);
    assign layer0_outputs[2716] = inputs[130];
    assign layer0_outputs[2717] = inputs[66];
    assign layer0_outputs[2718] = ~(inputs[116]) | (inputs[23]);
    assign layer0_outputs[2719] = 1'b0;
    assign layer0_outputs[2720] = ~(inputs[172]) | (inputs[94]);
    assign layer0_outputs[2721] = ~(inputs[18]);
    assign layer0_outputs[2722] = ~((inputs[218]) ^ (inputs[240]));
    assign layer0_outputs[2723] = 1'b1;
    assign layer0_outputs[2724] = (inputs[21]) & ~(inputs[216]);
    assign layer0_outputs[2725] = inputs[193];
    assign layer0_outputs[2726] = (inputs[98]) | (inputs[27]);
    assign layer0_outputs[2727] = inputs[22];
    assign layer0_outputs[2728] = inputs[134];
    assign layer0_outputs[2729] = (inputs[63]) & ~(inputs[242]);
    assign layer0_outputs[2730] = (inputs[79]) & ~(inputs[169]);
    assign layer0_outputs[2731] = (inputs[224]) & ~(inputs[94]);
    assign layer0_outputs[2732] = ~((inputs[36]) | (inputs[2]));
    assign layer0_outputs[2733] = ~((inputs[10]) | (inputs[152]));
    assign layer0_outputs[2734] = inputs[253];
    assign layer0_outputs[2735] = (inputs[110]) | (inputs[204]);
    assign layer0_outputs[2736] = 1'b0;
    assign layer0_outputs[2737] = ~(inputs[57]) | (inputs[225]);
    assign layer0_outputs[2738] = ~((inputs[211]) | (inputs[242]));
    assign layer0_outputs[2739] = ~(inputs[225]);
    assign layer0_outputs[2740] = ~((inputs[28]) | (inputs[34]));
    assign layer0_outputs[2741] = (inputs[113]) ^ (inputs[103]);
    assign layer0_outputs[2742] = ~(inputs[212]);
    assign layer0_outputs[2743] = inputs[255];
    assign layer0_outputs[2744] = (inputs[55]) & ~(inputs[17]);
    assign layer0_outputs[2745] = ~(inputs[232]) | (inputs[93]);
    assign layer0_outputs[2746] = ~(inputs[212]) | (inputs[223]);
    assign layer0_outputs[2747] = ~(inputs[47]) | (inputs[242]);
    assign layer0_outputs[2748] = (inputs[221]) & ~(inputs[67]);
    assign layer0_outputs[2749] = ~((inputs[106]) | (inputs[203]));
    assign layer0_outputs[2750] = (inputs[83]) & ~(inputs[110]);
    assign layer0_outputs[2751] = 1'b0;
    assign layer0_outputs[2752] = ~((inputs[131]) ^ (inputs[69]));
    assign layer0_outputs[2753] = ~(inputs[206]);
    assign layer0_outputs[2754] = ~(inputs[244]);
    assign layer0_outputs[2755] = (inputs[228]) & ~(inputs[14]);
    assign layer0_outputs[2756] = ~((inputs[232]) & (inputs[151]));
    assign layer0_outputs[2757] = (inputs[71]) & ~(inputs[112]);
    assign layer0_outputs[2758] = ~(inputs[205]);
    assign layer0_outputs[2759] = ~(inputs[12]);
    assign layer0_outputs[2760] = ~(inputs[154]);
    assign layer0_outputs[2761] = (inputs[251]) & ~(inputs[73]);
    assign layer0_outputs[2762] = (inputs[24]) & (inputs[52]);
    assign layer0_outputs[2763] = ~((inputs[163]) ^ (inputs[125]));
    assign layer0_outputs[2764] = ~(inputs[9]);
    assign layer0_outputs[2765] = inputs[99];
    assign layer0_outputs[2766] = (inputs[17]) ^ (inputs[2]);
    assign layer0_outputs[2767] = (inputs[207]) & ~(inputs[14]);
    assign layer0_outputs[2768] = ~(inputs[77]);
    assign layer0_outputs[2769] = inputs[15];
    assign layer0_outputs[2770] = ~((inputs[114]) | (inputs[54]));
    assign layer0_outputs[2771] = ~((inputs[26]) | (inputs[27]));
    assign layer0_outputs[2772] = (inputs[83]) & (inputs[83]);
    assign layer0_outputs[2773] = ~((inputs[192]) | (inputs[128]));
    assign layer0_outputs[2774] = ~(inputs[36]);
    assign layer0_outputs[2775] = ~(inputs[114]);
    assign layer0_outputs[2776] = (inputs[240]) & (inputs[167]);
    assign layer0_outputs[2777] = (inputs[230]) | (inputs[47]);
    assign layer0_outputs[2778] = ~((inputs[91]) | (inputs[224]));
    assign layer0_outputs[2779] = (inputs[12]) & ~(inputs[50]);
    assign layer0_outputs[2780] = (inputs[85]) ^ (inputs[111]);
    assign layer0_outputs[2781] = inputs[24];
    assign layer0_outputs[2782] = ~(inputs[159]) | (inputs[215]);
    assign layer0_outputs[2783] = (inputs[135]) | (inputs[105]);
    assign layer0_outputs[2784] = ~(inputs[206]) | (inputs[250]);
    assign layer0_outputs[2785] = ~(inputs[126]) | (inputs[191]);
    assign layer0_outputs[2786] = ~(inputs[45]) | (inputs[225]);
    assign layer0_outputs[2787] = ~(inputs[122]);
    assign layer0_outputs[2788] = ~(inputs[209]);
    assign layer0_outputs[2789] = (inputs[30]) ^ (inputs[112]);
    assign layer0_outputs[2790] = inputs[51];
    assign layer0_outputs[2791] = (inputs[159]) | (inputs[128]);
    assign layer0_outputs[2792] = (inputs[147]) | (inputs[236]);
    assign layer0_outputs[2793] = 1'b1;
    assign layer0_outputs[2794] = inputs[18];
    assign layer0_outputs[2795] = ~((inputs[95]) | (inputs[29]));
    assign layer0_outputs[2796] = (inputs[77]) | (inputs[123]);
    assign layer0_outputs[2797] = 1'b0;
    assign layer0_outputs[2798] = inputs[190];
    assign layer0_outputs[2799] = (inputs[161]) ^ (inputs[230]);
    assign layer0_outputs[2800] = (inputs[58]) ^ (inputs[138]);
    assign layer0_outputs[2801] = (inputs[99]) ^ (inputs[71]);
    assign layer0_outputs[2802] = (inputs[14]) & ~(inputs[220]);
    assign layer0_outputs[2803] = ~((inputs[68]) ^ (inputs[159]));
    assign layer0_outputs[2804] = (inputs[210]) & (inputs[240]);
    assign layer0_outputs[2805] = (inputs[95]) ^ (inputs[41]);
    assign layer0_outputs[2806] = inputs[164];
    assign layer0_outputs[2807] = ~((inputs[22]) | (inputs[95]));
    assign layer0_outputs[2808] = 1'b0;
    assign layer0_outputs[2809] = inputs[57];
    assign layer0_outputs[2810] = ~(inputs[197]) | (inputs[47]);
    assign layer0_outputs[2811] = ~(inputs[119]) | (inputs[216]);
    assign layer0_outputs[2812] = 1'b0;
    assign layer0_outputs[2813] = inputs[17];
    assign layer0_outputs[2814] = 1'b0;
    assign layer0_outputs[2815] = ~(inputs[133]) | (inputs[222]);
    assign layer0_outputs[2816] = (inputs[203]) ^ (inputs[79]);
    assign layer0_outputs[2817] = inputs[147];
    assign layer0_outputs[2818] = (inputs[90]) & ~(inputs[233]);
    assign layer0_outputs[2819] = (inputs[189]) | (inputs[209]);
    assign layer0_outputs[2820] = (inputs[237]) & ~(inputs[88]);
    assign layer0_outputs[2821] = ~((inputs[216]) & (inputs[203]));
    assign layer0_outputs[2822] = ~((inputs[253]) & (inputs[44]));
    assign layer0_outputs[2823] = ~((inputs[77]) ^ (inputs[29]));
    assign layer0_outputs[2824] = inputs[55];
    assign layer0_outputs[2825] = ~(inputs[103]);
    assign layer0_outputs[2826] = ~(inputs[84]);
    assign layer0_outputs[2827] = (inputs[106]) | (inputs[101]);
    assign layer0_outputs[2828] = inputs[209];
    assign layer0_outputs[2829] = inputs[153];
    assign layer0_outputs[2830] = inputs[128];
    assign layer0_outputs[2831] = inputs[31];
    assign layer0_outputs[2832] = ~((inputs[174]) & (inputs[59]));
    assign layer0_outputs[2833] = ~((inputs[70]) | (inputs[147]));
    assign layer0_outputs[2834] = ~((inputs[72]) | (inputs[253]));
    assign layer0_outputs[2835] = inputs[151];
    assign layer0_outputs[2836] = ~(inputs[0]);
    assign layer0_outputs[2837] = ~(inputs[161]);
    assign layer0_outputs[2838] = ~(inputs[104]);
    assign layer0_outputs[2839] = ~(inputs[148]);
    assign layer0_outputs[2840] = ~(inputs[97]);
    assign layer0_outputs[2841] = ~(inputs[225]) | (inputs[67]);
    assign layer0_outputs[2842] = ~(inputs[202]);
    assign layer0_outputs[2843] = ~(inputs[207]) | (inputs[242]);
    assign layer0_outputs[2844] = (inputs[60]) | (inputs[123]);
    assign layer0_outputs[2845] = ~(inputs[180]);
    assign layer0_outputs[2846] = ~(inputs[7]) | (inputs[161]);
    assign layer0_outputs[2847] = ~(inputs[178]);
    assign layer0_outputs[2848] = (inputs[143]) | (inputs[4]);
    assign layer0_outputs[2849] = (inputs[136]) & ~(inputs[3]);
    assign layer0_outputs[2850] = ~((inputs[1]) ^ (inputs[54]));
    assign layer0_outputs[2851] = inputs[166];
    assign layer0_outputs[2852] = ~((inputs[128]) ^ (inputs[146]));
    assign layer0_outputs[2853] = (inputs[40]) & ~(inputs[149]);
    assign layer0_outputs[2854] = (inputs[29]) ^ (inputs[88]);
    assign layer0_outputs[2855] = ~((inputs[116]) | (inputs[223]));
    assign layer0_outputs[2856] = ~(inputs[183]);
    assign layer0_outputs[2857] = ~(inputs[69]);
    assign layer0_outputs[2858] = ~((inputs[84]) ^ (inputs[164]));
    assign layer0_outputs[2859] = ~(inputs[163]);
    assign layer0_outputs[2860] = (inputs[130]) | (inputs[199]);
    assign layer0_outputs[2861] = ~((inputs[62]) | (inputs[134]));
    assign layer0_outputs[2862] = inputs[169];
    assign layer0_outputs[2863] = (inputs[27]) | (inputs[172]);
    assign layer0_outputs[2864] = (inputs[54]) | (inputs[13]);
    assign layer0_outputs[2865] = (inputs[202]) | (inputs[176]);
    assign layer0_outputs[2866] = ~((inputs[172]) | (inputs[203]));
    assign layer0_outputs[2867] = ~(inputs[99]);
    assign layer0_outputs[2868] = inputs[10];
    assign layer0_outputs[2869] = inputs[161];
    assign layer0_outputs[2870] = (inputs[34]) | (inputs[6]);
    assign layer0_outputs[2871] = ~((inputs[63]) ^ (inputs[19]));
    assign layer0_outputs[2872] = ~((inputs[57]) | (inputs[160]));
    assign layer0_outputs[2873] = ~(inputs[148]);
    assign layer0_outputs[2874] = ~(inputs[28]);
    assign layer0_outputs[2875] = (inputs[147]) | (inputs[209]);
    assign layer0_outputs[2876] = inputs[165];
    assign layer0_outputs[2877] = ~(inputs[96]);
    assign layer0_outputs[2878] = 1'b1;
    assign layer0_outputs[2879] = (inputs[162]) | (inputs[198]);
    assign layer0_outputs[2880] = inputs[240];
    assign layer0_outputs[2881] = (inputs[167]) ^ (inputs[129]);
    assign layer0_outputs[2882] = inputs[128];
    assign layer0_outputs[2883] = ~((inputs[150]) | (inputs[198]));
    assign layer0_outputs[2884] = (inputs[45]) & ~(inputs[254]);
    assign layer0_outputs[2885] = ~((inputs[42]) ^ (inputs[15]));
    assign layer0_outputs[2886] = (inputs[5]) & ~(inputs[158]);
    assign layer0_outputs[2887] = (inputs[100]) ^ (inputs[69]);
    assign layer0_outputs[2888] = inputs[5];
    assign layer0_outputs[2889] = (inputs[159]) & (inputs[129]);
    assign layer0_outputs[2890] = ~(inputs[136]) | (inputs[185]);
    assign layer0_outputs[2891] = ~((inputs[143]) ^ (inputs[152]));
    assign layer0_outputs[2892] = (inputs[129]) & ~(inputs[254]);
    assign layer0_outputs[2893] = (inputs[25]) & ~(inputs[178]);
    assign layer0_outputs[2894] = ~((inputs[2]) & (inputs[162]));
    assign layer0_outputs[2895] = ~(inputs[73]);
    assign layer0_outputs[2896] = ~(inputs[114]);
    assign layer0_outputs[2897] = ~((inputs[139]) ^ (inputs[141]));
    assign layer0_outputs[2898] = inputs[27];
    assign layer0_outputs[2899] = (inputs[97]) ^ (inputs[187]);
    assign layer0_outputs[2900] = (inputs[223]) & (inputs[213]);
    assign layer0_outputs[2901] = (inputs[9]) & ~(inputs[190]);
    assign layer0_outputs[2902] = ~(inputs[221]);
    assign layer0_outputs[2903] = ~(inputs[13]);
    assign layer0_outputs[2904] = ~((inputs[159]) & (inputs[179]));
    assign layer0_outputs[2905] = ~(inputs[178]);
    assign layer0_outputs[2906] = ~((inputs[26]) | (inputs[226]));
    assign layer0_outputs[2907] = ~(inputs[14]);
    assign layer0_outputs[2908] = ~((inputs[27]) | (inputs[132]));
    assign layer0_outputs[2909] = 1'b0;
    assign layer0_outputs[2910] = ~(inputs[90]) | (inputs[112]);
    assign layer0_outputs[2911] = ~(inputs[34]);
    assign layer0_outputs[2912] = inputs[151];
    assign layer0_outputs[2913] = inputs[191];
    assign layer0_outputs[2914] = ~(inputs[214]) | (inputs[173]);
    assign layer0_outputs[2915] = 1'b0;
    assign layer0_outputs[2916] = ~((inputs[134]) ^ (inputs[248]));
    assign layer0_outputs[2917] = (inputs[147]) & ~(inputs[63]);
    assign layer0_outputs[2918] = ~((inputs[83]) ^ (inputs[0]));
    assign layer0_outputs[2919] = inputs[211];
    assign layer0_outputs[2920] = (inputs[23]) & (inputs[26]);
    assign layer0_outputs[2921] = (inputs[194]) | (inputs[221]);
    assign layer0_outputs[2922] = ~((inputs[96]) | (inputs[70]));
    assign layer0_outputs[2923] = ~(inputs[86]);
    assign layer0_outputs[2924] = inputs[195];
    assign layer0_outputs[2925] = ~((inputs[198]) ^ (inputs[77]));
    assign layer0_outputs[2926] = inputs[150];
    assign layer0_outputs[2927] = ~(inputs[201]);
    assign layer0_outputs[2928] = ~((inputs[249]) & (inputs[244]));
    assign layer0_outputs[2929] = ~(inputs[183]) | (inputs[216]);
    assign layer0_outputs[2930] = inputs[236];
    assign layer0_outputs[2931] = (inputs[230]) & ~(inputs[35]);
    assign layer0_outputs[2932] = ~(inputs[135]);
    assign layer0_outputs[2933] = ~((inputs[159]) & (inputs[243]));
    assign layer0_outputs[2934] = ~((inputs[223]) | (inputs[152]));
    assign layer0_outputs[2935] = (inputs[178]) ^ (inputs[180]);
    assign layer0_outputs[2936] = ~(inputs[170]) | (inputs[85]);
    assign layer0_outputs[2937] = ~((inputs[55]) ^ (inputs[55]));
    assign layer0_outputs[2938] = (inputs[234]) ^ (inputs[86]);
    assign layer0_outputs[2939] = inputs[211];
    assign layer0_outputs[2940] = (inputs[27]) & ~(inputs[140]);
    assign layer0_outputs[2941] = (inputs[173]) & ~(inputs[3]);
    assign layer0_outputs[2942] = (inputs[22]) & (inputs[41]);
    assign layer0_outputs[2943] = (inputs[10]) & ~(inputs[246]);
    assign layer0_outputs[2944] = ~((inputs[49]) | (inputs[29]));
    assign layer0_outputs[2945] = inputs[220];
    assign layer0_outputs[2946] = (inputs[221]) & ~(inputs[177]);
    assign layer0_outputs[2947] = (inputs[212]) | (inputs[127]);
    assign layer0_outputs[2948] = (inputs[206]) | (inputs[217]);
    assign layer0_outputs[2949] = ~(inputs[72]);
    assign layer0_outputs[2950] = (inputs[54]) | (inputs[101]);
    assign layer0_outputs[2951] = inputs[75];
    assign layer0_outputs[2952] = (inputs[221]) & ~(inputs[41]);
    assign layer0_outputs[2953] = ~((inputs[233]) | (inputs[200]));
    assign layer0_outputs[2954] = inputs[192];
    assign layer0_outputs[2955] = ~((inputs[193]) | (inputs[133]));
    assign layer0_outputs[2956] = inputs[207];
    assign layer0_outputs[2957] = (inputs[61]) | (inputs[181]);
    assign layer0_outputs[2958] = ~(inputs[48]);
    assign layer0_outputs[2959] = (inputs[245]) | (inputs[177]);
    assign layer0_outputs[2960] = ~((inputs[251]) ^ (inputs[164]));
    assign layer0_outputs[2961] = (inputs[148]) ^ (inputs[3]);
    assign layer0_outputs[2962] = inputs[4];
    assign layer0_outputs[2963] = (inputs[70]) & (inputs[127]);
    assign layer0_outputs[2964] = inputs[169];
    assign layer0_outputs[2965] = inputs[71];
    assign layer0_outputs[2966] = (inputs[206]) | (inputs[238]);
    assign layer0_outputs[2967] = ~((inputs[53]) ^ (inputs[221]));
    assign layer0_outputs[2968] = ~((inputs[90]) ^ (inputs[162]));
    assign layer0_outputs[2969] = inputs[90];
    assign layer0_outputs[2970] = ~(inputs[137]);
    assign layer0_outputs[2971] = 1'b0;
    assign layer0_outputs[2972] = ~(inputs[196]);
    assign layer0_outputs[2973] = ~(inputs[106]) | (inputs[46]);
    assign layer0_outputs[2974] = (inputs[176]) | (inputs[233]);
    assign layer0_outputs[2975] = (inputs[109]) | (inputs[95]);
    assign layer0_outputs[2976] = ~((inputs[225]) | (inputs[242]));
    assign layer0_outputs[2977] = ~((inputs[82]) | (inputs[215]));
    assign layer0_outputs[2978] = inputs[31];
    assign layer0_outputs[2979] = ~(inputs[72]);
    assign layer0_outputs[2980] = ~((inputs[19]) & (inputs[46]));
    assign layer0_outputs[2981] = (inputs[235]) ^ (inputs[116]);
    assign layer0_outputs[2982] = inputs[109];
    assign layer0_outputs[2983] = (inputs[191]) | (inputs[49]);
    assign layer0_outputs[2984] = ~((inputs[227]) | (inputs[209]));
    assign layer0_outputs[2985] = ~(inputs[151]) | (inputs[210]);
    assign layer0_outputs[2986] = ~(inputs[73]) | (inputs[55]);
    assign layer0_outputs[2987] = ~((inputs[222]) ^ (inputs[60]));
    assign layer0_outputs[2988] = (inputs[37]) & ~(inputs[18]);
    assign layer0_outputs[2989] = 1'b0;
    assign layer0_outputs[2990] = ~(inputs[71]);
    assign layer0_outputs[2991] = ~(inputs[130]);
    assign layer0_outputs[2992] = (inputs[81]) ^ (inputs[147]);
    assign layer0_outputs[2993] = ~(inputs[211]);
    assign layer0_outputs[2994] = ~((inputs[101]) ^ (inputs[112]));
    assign layer0_outputs[2995] = ~((inputs[224]) | (inputs[31]));
    assign layer0_outputs[2996] = 1'b0;
    assign layer0_outputs[2997] = inputs[87];
    assign layer0_outputs[2998] = (inputs[104]) & (inputs[188]);
    assign layer0_outputs[2999] = ~(inputs[0]);
    assign layer0_outputs[3000] = inputs[62];
    assign layer0_outputs[3001] = ~((inputs[62]) ^ (inputs[17]));
    assign layer0_outputs[3002] = ~(inputs[99]) | (inputs[3]);
    assign layer0_outputs[3003] = (inputs[188]) & ~(inputs[102]);
    assign layer0_outputs[3004] = (inputs[50]) & ~(inputs[122]);
    assign layer0_outputs[3005] = (inputs[63]) & ~(inputs[161]);
    assign layer0_outputs[3006] = inputs[197];
    assign layer0_outputs[3007] = ~((inputs[162]) | (inputs[52]));
    assign layer0_outputs[3008] = ~((inputs[3]) | (inputs[189]));
    assign layer0_outputs[3009] = (inputs[81]) | (inputs[139]);
    assign layer0_outputs[3010] = ~((inputs[230]) | (inputs[113]));
    assign layer0_outputs[3011] = ~(inputs[176]) | (inputs[250]);
    assign layer0_outputs[3012] = ~((inputs[188]) & (inputs[179]));
    assign layer0_outputs[3013] = 1'b0;
    assign layer0_outputs[3014] = (inputs[194]) & ~(inputs[18]);
    assign layer0_outputs[3015] = ~(inputs[105]) | (inputs[145]);
    assign layer0_outputs[3016] = 1'b0;
    assign layer0_outputs[3017] = inputs[223];
    assign layer0_outputs[3018] = 1'b0;
    assign layer0_outputs[3019] = (inputs[195]) ^ (inputs[244]);
    assign layer0_outputs[3020] = 1'b0;
    assign layer0_outputs[3021] = (inputs[6]) | (inputs[210]);
    assign layer0_outputs[3022] = inputs[158];
    assign layer0_outputs[3023] = inputs[129];
    assign layer0_outputs[3024] = ~((inputs[95]) ^ (inputs[167]));
    assign layer0_outputs[3025] = inputs[78];
    assign layer0_outputs[3026] = inputs[217];
    assign layer0_outputs[3027] = 1'b1;
    assign layer0_outputs[3028] = ~(inputs[97]);
    assign layer0_outputs[3029] = ~(inputs[99]);
    assign layer0_outputs[3030] = ~((inputs[177]) ^ (inputs[198]));
    assign layer0_outputs[3031] = (inputs[50]) | (inputs[248]);
    assign layer0_outputs[3032] = (inputs[28]) | (inputs[34]);
    assign layer0_outputs[3033] = (inputs[49]) ^ (inputs[139]);
    assign layer0_outputs[3034] = ~((inputs[59]) ^ (inputs[172]));
    assign layer0_outputs[3035] = (inputs[107]) & ~(inputs[82]);
    assign layer0_outputs[3036] = 1'b0;
    assign layer0_outputs[3037] = (inputs[71]) & ~(inputs[22]);
    assign layer0_outputs[3038] = ~((inputs[31]) | (inputs[219]));
    assign layer0_outputs[3039] = (inputs[53]) ^ (inputs[132]);
    assign layer0_outputs[3040] = (inputs[238]) | (inputs[88]);
    assign layer0_outputs[3041] = ~(inputs[34]);
    assign layer0_outputs[3042] = ~(inputs[109]);
    assign layer0_outputs[3043] = 1'b0;
    assign layer0_outputs[3044] = inputs[115];
    assign layer0_outputs[3045] = ~(inputs[81]) | (inputs[170]);
    assign layer0_outputs[3046] = ~(inputs[24]) | (inputs[118]);
    assign layer0_outputs[3047] = inputs[136];
    assign layer0_outputs[3048] = (inputs[77]) ^ (inputs[237]);
    assign layer0_outputs[3049] = inputs[157];
    assign layer0_outputs[3050] = (inputs[119]) & ~(inputs[31]);
    assign layer0_outputs[3051] = inputs[229];
    assign layer0_outputs[3052] = ~((inputs[236]) & (inputs[25]));
    assign layer0_outputs[3053] = inputs[36];
    assign layer0_outputs[3054] = ~((inputs[238]) | (inputs[99]));
    assign layer0_outputs[3055] = (inputs[234]) & (inputs[11]);
    assign layer0_outputs[3056] = (inputs[40]) & (inputs[250]);
    assign layer0_outputs[3057] = ~(inputs[219]);
    assign layer0_outputs[3058] = ~(inputs[168]);
    assign layer0_outputs[3059] = ~(inputs[60]) | (inputs[164]);
    assign layer0_outputs[3060] = ~((inputs[254]) | (inputs[179]));
    assign layer0_outputs[3061] = ~(inputs[123]) | (inputs[161]);
    assign layer0_outputs[3062] = ~((inputs[184]) | (inputs[185]));
    assign layer0_outputs[3063] = ~(inputs[235]) | (inputs[112]);
    assign layer0_outputs[3064] = ~((inputs[204]) | (inputs[120]));
    assign layer0_outputs[3065] = ~((inputs[41]) | (inputs[49]));
    assign layer0_outputs[3066] = ~((inputs[134]) ^ (inputs[114]));
    assign layer0_outputs[3067] = inputs[182];
    assign layer0_outputs[3068] = ~((inputs[229]) | (inputs[177]));
    assign layer0_outputs[3069] = (inputs[58]) & ~(inputs[178]);
    assign layer0_outputs[3070] = (inputs[50]) | (inputs[89]);
    assign layer0_outputs[3071] = ~(inputs[101]);
    assign layer0_outputs[3072] = (inputs[248]) & ~(inputs[121]);
    assign layer0_outputs[3073] = 1'b0;
    assign layer0_outputs[3074] = ~((inputs[92]) | (inputs[60]));
    assign layer0_outputs[3075] = (inputs[170]) ^ (inputs[67]);
    assign layer0_outputs[3076] = (inputs[142]) ^ (inputs[198]);
    assign layer0_outputs[3077] = 1'b0;
    assign layer0_outputs[3078] = ~((inputs[49]) & (inputs[230]));
    assign layer0_outputs[3079] = ~(inputs[219]);
    assign layer0_outputs[3080] = inputs[58];
    assign layer0_outputs[3081] = inputs[241];
    assign layer0_outputs[3082] = inputs[35];
    assign layer0_outputs[3083] = inputs[222];
    assign layer0_outputs[3084] = inputs[75];
    assign layer0_outputs[3085] = ~(inputs[100]) | (inputs[109]);
    assign layer0_outputs[3086] = ~((inputs[29]) | (inputs[131]));
    assign layer0_outputs[3087] = ~((inputs[201]) | (inputs[188]));
    assign layer0_outputs[3088] = ~((inputs[180]) | (inputs[153]));
    assign layer0_outputs[3089] = inputs[185];
    assign layer0_outputs[3090] = inputs[67];
    assign layer0_outputs[3091] = (inputs[34]) & ~(inputs[11]);
    assign layer0_outputs[3092] = (inputs[137]) & ~(inputs[32]);
    assign layer0_outputs[3093] = ~((inputs[227]) | (inputs[34]));
    assign layer0_outputs[3094] = (inputs[12]) | (inputs[115]);
    assign layer0_outputs[3095] = ~((inputs[139]) ^ (inputs[175]));
    assign layer0_outputs[3096] = (inputs[20]) ^ (inputs[169]);
    assign layer0_outputs[3097] = ~(inputs[23]) | (inputs[143]);
    assign layer0_outputs[3098] = inputs[87];
    assign layer0_outputs[3099] = ~((inputs[50]) & (inputs[184]));
    assign layer0_outputs[3100] = ~(inputs[172]);
    assign layer0_outputs[3101] = (inputs[30]) & ~(inputs[155]);
    assign layer0_outputs[3102] = (inputs[187]) | (inputs[13]);
    assign layer0_outputs[3103] = ~((inputs[243]) | (inputs[134]));
    assign layer0_outputs[3104] = (inputs[255]) & ~(inputs[251]);
    assign layer0_outputs[3105] = ~(inputs[138]);
    assign layer0_outputs[3106] = (inputs[224]) & ~(inputs[131]);
    assign layer0_outputs[3107] = inputs[46];
    assign layer0_outputs[3108] = inputs[24];
    assign layer0_outputs[3109] = ~(inputs[104]);
    assign layer0_outputs[3110] = ~(inputs[189]) | (inputs[228]);
    assign layer0_outputs[3111] = ~((inputs[163]) ^ (inputs[182]));
    assign layer0_outputs[3112] = ~(inputs[64]) | (inputs[43]);
    assign layer0_outputs[3113] = ~(inputs[66]) | (inputs[157]);
    assign layer0_outputs[3114] = inputs[24];
    assign layer0_outputs[3115] = ~(inputs[91]) | (inputs[214]);
    assign layer0_outputs[3116] = (inputs[232]) & ~(inputs[56]);
    assign layer0_outputs[3117] = inputs[94];
    assign layer0_outputs[3118] = ~((inputs[21]) ^ (inputs[45]));
    assign layer0_outputs[3119] = ~((inputs[182]) | (inputs[35]));
    assign layer0_outputs[3120] = (inputs[34]) | (inputs[9]);
    assign layer0_outputs[3121] = ~(inputs[119]);
    assign layer0_outputs[3122] = inputs[211];
    assign layer0_outputs[3123] = ~(inputs[30]) | (inputs[127]);
    assign layer0_outputs[3124] = 1'b0;
    assign layer0_outputs[3125] = (inputs[228]) | (inputs[194]);
    assign layer0_outputs[3126] = (inputs[218]) & ~(inputs[115]);
    assign layer0_outputs[3127] = inputs[62];
    assign layer0_outputs[3128] = 1'b1;
    assign layer0_outputs[3129] = inputs[40];
    assign layer0_outputs[3130] = inputs[119];
    assign layer0_outputs[3131] = ~(inputs[43]);
    assign layer0_outputs[3132] = (inputs[118]) | (inputs[211]);
    assign layer0_outputs[3133] = ~((inputs[155]) | (inputs[255]));
    assign layer0_outputs[3134] = inputs[73];
    assign layer0_outputs[3135] = ~(inputs[209]);
    assign layer0_outputs[3136] = ~((inputs[6]) | (inputs[192]));
    assign layer0_outputs[3137] = (inputs[57]) & ~(inputs[50]);
    assign layer0_outputs[3138] = ~(inputs[72]);
    assign layer0_outputs[3139] = ~(inputs[57]);
    assign layer0_outputs[3140] = ~((inputs[146]) | (inputs[95]));
    assign layer0_outputs[3141] = (inputs[221]) & (inputs[123]);
    assign layer0_outputs[3142] = ~((inputs[210]) | (inputs[144]));
    assign layer0_outputs[3143] = inputs[69];
    assign layer0_outputs[3144] = (inputs[78]) | (inputs[223]);
    assign layer0_outputs[3145] = ~((inputs[51]) ^ (inputs[46]));
    assign layer0_outputs[3146] = inputs[115];
    assign layer0_outputs[3147] = inputs[166];
    assign layer0_outputs[3148] = ~(inputs[91]) | (inputs[146]);
    assign layer0_outputs[3149] = (inputs[26]) & ~(inputs[252]);
    assign layer0_outputs[3150] = ~((inputs[18]) | (inputs[118]));
    assign layer0_outputs[3151] = inputs[148];
    assign layer0_outputs[3152] = ~((inputs[23]) ^ (inputs[124]));
    assign layer0_outputs[3153] = ~(inputs[30]);
    assign layer0_outputs[3154] = 1'b0;
    assign layer0_outputs[3155] = ~(inputs[129]) | (inputs[220]);
    assign layer0_outputs[3156] = ~(inputs[45]) | (inputs[173]);
    assign layer0_outputs[3157] = ~((inputs[132]) ^ (inputs[255]));
    assign layer0_outputs[3158] = (inputs[220]) & ~(inputs[1]);
    assign layer0_outputs[3159] = ~(inputs[98]);
    assign layer0_outputs[3160] = ~(inputs[12]);
    assign layer0_outputs[3161] = (inputs[180]) ^ (inputs[25]);
    assign layer0_outputs[3162] = ~((inputs[129]) | (inputs[99]));
    assign layer0_outputs[3163] = (inputs[76]) | (inputs[141]);
    assign layer0_outputs[3164] = (inputs[14]) | (inputs[120]);
    assign layer0_outputs[3165] = ~((inputs[163]) | (inputs[85]));
    assign layer0_outputs[3166] = ~(inputs[235]) | (inputs[47]);
    assign layer0_outputs[3167] = inputs[208];
    assign layer0_outputs[3168] = (inputs[35]) & ~(inputs[251]);
    assign layer0_outputs[3169] = ~((inputs[142]) & (inputs[120]));
    assign layer0_outputs[3170] = inputs[103];
    assign layer0_outputs[3171] = ~(inputs[165]);
    assign layer0_outputs[3172] = inputs[86];
    assign layer0_outputs[3173] = (inputs[35]) | (inputs[174]);
    assign layer0_outputs[3174] = ~((inputs[253]) & (inputs[5]));
    assign layer0_outputs[3175] = inputs[216];
    assign layer0_outputs[3176] = (inputs[40]) & ~(inputs[108]);
    assign layer0_outputs[3177] = (inputs[220]) | (inputs[175]);
    assign layer0_outputs[3178] = (inputs[34]) & ~(inputs[128]);
    assign layer0_outputs[3179] = ~(inputs[215]) | (inputs[60]);
    assign layer0_outputs[3180] = (inputs[96]) | (inputs[98]);
    assign layer0_outputs[3181] = ~(inputs[221]) | (inputs[7]);
    assign layer0_outputs[3182] = 1'b0;
    assign layer0_outputs[3183] = (inputs[57]) & (inputs[212]);
    assign layer0_outputs[3184] = inputs[88];
    assign layer0_outputs[3185] = (inputs[52]) & ~(inputs[134]);
    assign layer0_outputs[3186] = ~(inputs[149]);
    assign layer0_outputs[3187] = (inputs[248]) | (inputs[231]);
    assign layer0_outputs[3188] = ~((inputs[148]) & (inputs[142]));
    assign layer0_outputs[3189] = ~((inputs[203]) | (inputs[4]));
    assign layer0_outputs[3190] = ~((inputs[164]) & (inputs[140]));
    assign layer0_outputs[3191] = 1'b1;
    assign layer0_outputs[3192] = ~(inputs[204]);
    assign layer0_outputs[3193] = (inputs[8]) & ~(inputs[14]);
    assign layer0_outputs[3194] = (inputs[102]) & ~(inputs[131]);
    assign layer0_outputs[3195] = ~(inputs[37]);
    assign layer0_outputs[3196] = (inputs[240]) ^ (inputs[118]);
    assign layer0_outputs[3197] = ~((inputs[50]) ^ (inputs[60]));
    assign layer0_outputs[3198] = ~((inputs[73]) ^ (inputs[171]));
    assign layer0_outputs[3199] = ~(inputs[172]) | (inputs[147]);
    assign layer0_outputs[3200] = inputs[45];
    assign layer0_outputs[3201] = (inputs[81]) & ~(inputs[190]);
    assign layer0_outputs[3202] = ~((inputs[195]) | (inputs[225]));
    assign layer0_outputs[3203] = ~((inputs[149]) | (inputs[134]));
    assign layer0_outputs[3204] = ~((inputs[177]) | (inputs[83]));
    assign layer0_outputs[3205] = ~(inputs[98]) | (inputs[111]);
    assign layer0_outputs[3206] = ~(inputs[102]);
    assign layer0_outputs[3207] = (inputs[248]) & (inputs[111]);
    assign layer0_outputs[3208] = ~(inputs[9]);
    assign layer0_outputs[3209] = ~((inputs[204]) | (inputs[235]));
    assign layer0_outputs[3210] = ~((inputs[97]) ^ (inputs[145]));
    assign layer0_outputs[3211] = ~((inputs[236]) | (inputs[32]));
    assign layer0_outputs[3212] = (inputs[22]) ^ (inputs[48]);
    assign layer0_outputs[3213] = (inputs[32]) ^ (inputs[70]);
    assign layer0_outputs[3214] = inputs[151];
    assign layer0_outputs[3215] = ~(inputs[212]);
    assign layer0_outputs[3216] = (inputs[42]) & ~(inputs[103]);
    assign layer0_outputs[3217] = ~((inputs[68]) ^ (inputs[35]));
    assign layer0_outputs[3218] = ~(inputs[192]);
    assign layer0_outputs[3219] = (inputs[58]) & ~(inputs[48]);
    assign layer0_outputs[3220] = ~(inputs[124]) | (inputs[157]);
    assign layer0_outputs[3221] = ~((inputs[105]) ^ (inputs[171]));
    assign layer0_outputs[3222] = inputs[129];
    assign layer0_outputs[3223] = (inputs[151]) | (inputs[239]);
    assign layer0_outputs[3224] = ~(inputs[117]);
    assign layer0_outputs[3225] = (inputs[245]) & ~(inputs[14]);
    assign layer0_outputs[3226] = ~(inputs[222]) | (inputs[36]);
    assign layer0_outputs[3227] = ~(inputs[93]);
    assign layer0_outputs[3228] = (inputs[251]) ^ (inputs[151]);
    assign layer0_outputs[3229] = (inputs[130]) | (inputs[152]);
    assign layer0_outputs[3230] = ~((inputs[157]) ^ (inputs[109]));
    assign layer0_outputs[3231] = (inputs[146]) ^ (inputs[229]);
    assign layer0_outputs[3232] = (inputs[236]) ^ (inputs[17]);
    assign layer0_outputs[3233] = (inputs[251]) | (inputs[153]);
    assign layer0_outputs[3234] = ~(inputs[131]) | (inputs[73]);
    assign layer0_outputs[3235] = (inputs[112]) & (inputs[196]);
    assign layer0_outputs[3236] = (inputs[130]) | (inputs[134]);
    assign layer0_outputs[3237] = ~(inputs[249]);
    assign layer0_outputs[3238] = ~(inputs[85]);
    assign layer0_outputs[3239] = (inputs[186]) & ~(inputs[98]);
    assign layer0_outputs[3240] = 1'b1;
    assign layer0_outputs[3241] = (inputs[90]) & ~(inputs[238]);
    assign layer0_outputs[3242] = (inputs[206]) ^ (inputs[107]);
    assign layer0_outputs[3243] = inputs[229];
    assign layer0_outputs[3244] = ~(inputs[202]);
    assign layer0_outputs[3245] = ~((inputs[26]) ^ (inputs[159]));
    assign layer0_outputs[3246] = ~(inputs[156]);
    assign layer0_outputs[3247] = ~((inputs[15]) | (inputs[254]));
    assign layer0_outputs[3248] = (inputs[203]) ^ (inputs[140]);
    assign layer0_outputs[3249] = ~(inputs[93]);
    assign layer0_outputs[3250] = (inputs[146]) | (inputs[110]);
    assign layer0_outputs[3251] = (inputs[237]) ^ (inputs[207]);
    assign layer0_outputs[3252] = ~(inputs[224]);
    assign layer0_outputs[3253] = inputs[120];
    assign layer0_outputs[3254] = ~((inputs[229]) | (inputs[244]));
    assign layer0_outputs[3255] = 1'b1;
    assign layer0_outputs[3256] = ~(inputs[58]);
    assign layer0_outputs[3257] = (inputs[36]) ^ (inputs[210]);
    assign layer0_outputs[3258] = (inputs[199]) & ~(inputs[135]);
    assign layer0_outputs[3259] = ~(inputs[188]) | (inputs[112]);
    assign layer0_outputs[3260] = (inputs[100]) | (inputs[253]);
    assign layer0_outputs[3261] = ~((inputs[10]) | (inputs[4]));
    assign layer0_outputs[3262] = (inputs[235]) & ~(inputs[119]);
    assign layer0_outputs[3263] = (inputs[137]) & ~(inputs[54]);
    assign layer0_outputs[3264] = ~(inputs[10]);
    assign layer0_outputs[3265] = (inputs[39]) | (inputs[97]);
    assign layer0_outputs[3266] = ~((inputs[109]) & (inputs[194]));
    assign layer0_outputs[3267] = inputs[228];
    assign layer0_outputs[3268] = ~(inputs[112]) | (inputs[127]);
    assign layer0_outputs[3269] = ~(inputs[18]) | (inputs[13]);
    assign layer0_outputs[3270] = inputs[73];
    assign layer0_outputs[3271] = ~(inputs[166]);
    assign layer0_outputs[3272] = ~((inputs[147]) ^ (inputs[97]));
    assign layer0_outputs[3273] = ~((inputs[114]) | (inputs[148]));
    assign layer0_outputs[3274] = inputs[175];
    assign layer0_outputs[3275] = (inputs[176]) | (inputs[99]);
    assign layer0_outputs[3276] = ~(inputs[90]);
    assign layer0_outputs[3277] = ~((inputs[182]) & (inputs[18]));
    assign layer0_outputs[3278] = inputs[121];
    assign layer0_outputs[3279] = (inputs[145]) & ~(inputs[59]);
    assign layer0_outputs[3280] = 1'b1;
    assign layer0_outputs[3281] = ~((inputs[4]) ^ (inputs[16]));
    assign layer0_outputs[3282] = ~(inputs[137]);
    assign layer0_outputs[3283] = (inputs[40]) & ~(inputs[129]);
    assign layer0_outputs[3284] = ~(inputs[164]);
    assign layer0_outputs[3285] = (inputs[40]) | (inputs[20]);
    assign layer0_outputs[3286] = inputs[199];
    assign layer0_outputs[3287] = inputs[250];
    assign layer0_outputs[3288] = (inputs[110]) & (inputs[63]);
    assign layer0_outputs[3289] = ~(inputs[8]);
    assign layer0_outputs[3290] = (inputs[156]) & (inputs[217]);
    assign layer0_outputs[3291] = (inputs[143]) | (inputs[231]);
    assign layer0_outputs[3292] = inputs[158];
    assign layer0_outputs[3293] = ~(inputs[173]);
    assign layer0_outputs[3294] = (inputs[226]) | (inputs[223]);
    assign layer0_outputs[3295] = (inputs[201]) ^ (inputs[233]);
    assign layer0_outputs[3296] = ~((inputs[172]) & (inputs[245]));
    assign layer0_outputs[3297] = ~(inputs[11]);
    assign layer0_outputs[3298] = inputs[217];
    assign layer0_outputs[3299] = ~(inputs[42]);
    assign layer0_outputs[3300] = ~(inputs[76]);
    assign layer0_outputs[3301] = (inputs[248]) & ~(inputs[106]);
    assign layer0_outputs[3302] = (inputs[1]) & (inputs[82]);
    assign layer0_outputs[3303] = ~(inputs[100]);
    assign layer0_outputs[3304] = ~(inputs[72]) | (inputs[82]);
    assign layer0_outputs[3305] = ~((inputs[221]) & (inputs[221]));
    assign layer0_outputs[3306] = ~(inputs[217]);
    assign layer0_outputs[3307] = ~((inputs[242]) | (inputs[127]));
    assign layer0_outputs[3308] = (inputs[248]) & ~(inputs[75]);
    assign layer0_outputs[3309] = inputs[232];
    assign layer0_outputs[3310] = (inputs[242]) & ~(inputs[98]);
    assign layer0_outputs[3311] = ~((inputs[116]) | (inputs[254]));
    assign layer0_outputs[3312] = (inputs[29]) & (inputs[145]);
    assign layer0_outputs[3313] = (inputs[128]) ^ (inputs[164]);
    assign layer0_outputs[3314] = ~(inputs[43]) | (inputs[239]);
    assign layer0_outputs[3315] = inputs[65];
    assign layer0_outputs[3316] = ~(inputs[166]) | (inputs[62]);
    assign layer0_outputs[3317] = (inputs[170]) & ~(inputs[226]);
    assign layer0_outputs[3318] = ~(inputs[20]) | (inputs[192]);
    assign layer0_outputs[3319] = ~((inputs[1]) | (inputs[238]));
    assign layer0_outputs[3320] = inputs[123];
    assign layer0_outputs[3321] = (inputs[15]) & ~(inputs[53]);
    assign layer0_outputs[3322] = (inputs[245]) ^ (inputs[214]);
    assign layer0_outputs[3323] = ~((inputs[1]) | (inputs[35]));
    assign layer0_outputs[3324] = ~(inputs[59]) | (inputs[16]);
    assign layer0_outputs[3325] = ~(inputs[70]) | (inputs[145]);
    assign layer0_outputs[3326] = 1'b1;
    assign layer0_outputs[3327] = ~((inputs[85]) ^ (inputs[229]));
    assign layer0_outputs[3328] = inputs[53];
    assign layer0_outputs[3329] = ~((inputs[191]) | (inputs[78]));
    assign layer0_outputs[3330] = ~(inputs[188]);
    assign layer0_outputs[3331] = (inputs[122]) & ~(inputs[164]);
    assign layer0_outputs[3332] = (inputs[208]) ^ (inputs[222]);
    assign layer0_outputs[3333] = ~((inputs[48]) | (inputs[119]));
    assign layer0_outputs[3334] = ~((inputs[60]) ^ (inputs[186]));
    assign layer0_outputs[3335] = ~((inputs[133]) & (inputs[136]));
    assign layer0_outputs[3336] = 1'b1;
    assign layer0_outputs[3337] = ~(inputs[251]) | (inputs[55]);
    assign layer0_outputs[3338] = ~((inputs[120]) & (inputs[72]));
    assign layer0_outputs[3339] = ~(inputs[237]);
    assign layer0_outputs[3340] = (inputs[218]) ^ (inputs[186]);
    assign layer0_outputs[3341] = ~(inputs[7]);
    assign layer0_outputs[3342] = (inputs[64]) | (inputs[2]);
    assign layer0_outputs[3343] = (inputs[158]) ^ (inputs[78]);
    assign layer0_outputs[3344] = ~((inputs[20]) ^ (inputs[237]));
    assign layer0_outputs[3345] = (inputs[214]) | (inputs[95]);
    assign layer0_outputs[3346] = ~(inputs[117]) | (inputs[94]);
    assign layer0_outputs[3347] = ~(inputs[178]);
    assign layer0_outputs[3348] = ~((inputs[236]) | (inputs[215]));
    assign layer0_outputs[3349] = ~((inputs[15]) ^ (inputs[145]));
    assign layer0_outputs[3350] = ~((inputs[181]) | (inputs[194]));
    assign layer0_outputs[3351] = (inputs[199]) | (inputs[234]);
    assign layer0_outputs[3352] = ~((inputs[68]) | (inputs[198]));
    assign layer0_outputs[3353] = ~((inputs[222]) | (inputs[216]));
    assign layer0_outputs[3354] = ~((inputs[133]) ^ (inputs[86]));
    assign layer0_outputs[3355] = ~((inputs[25]) | (inputs[143]));
    assign layer0_outputs[3356] = ~(inputs[19]);
    assign layer0_outputs[3357] = 1'b0;
    assign layer0_outputs[3358] = (inputs[222]) | (inputs[198]);
    assign layer0_outputs[3359] = inputs[101];
    assign layer0_outputs[3360] = ~((inputs[210]) ^ (inputs[219]));
    assign layer0_outputs[3361] = ~(inputs[77]);
    assign layer0_outputs[3362] = ~(inputs[44]);
    assign layer0_outputs[3363] = (inputs[183]) ^ (inputs[238]);
    assign layer0_outputs[3364] = inputs[229];
    assign layer0_outputs[3365] = ~(inputs[212]) | (inputs[130]);
    assign layer0_outputs[3366] = ~(inputs[166]);
    assign layer0_outputs[3367] = (inputs[40]) & (inputs[38]);
    assign layer0_outputs[3368] = inputs[91];
    assign layer0_outputs[3369] = ~(inputs[91]) | (inputs[240]);
    assign layer0_outputs[3370] = ~(inputs[179]);
    assign layer0_outputs[3371] = 1'b0;
    assign layer0_outputs[3372] = (inputs[205]) & ~(inputs[77]);
    assign layer0_outputs[3373] = ~(inputs[58]);
    assign layer0_outputs[3374] = (inputs[173]) ^ (inputs[111]);
    assign layer0_outputs[3375] = ~(inputs[148]);
    assign layer0_outputs[3376] = inputs[42];
    assign layer0_outputs[3377] = (inputs[81]) ^ (inputs[68]);
    assign layer0_outputs[3378] = inputs[221];
    assign layer0_outputs[3379] = ~((inputs[213]) | (inputs[234]));
    assign layer0_outputs[3380] = ~(inputs[210]);
    assign layer0_outputs[3381] = (inputs[38]) & ~(inputs[163]);
    assign layer0_outputs[3382] = ~((inputs[225]) | (inputs[21]));
    assign layer0_outputs[3383] = ~(inputs[110]);
    assign layer0_outputs[3384] = ~(inputs[156]);
    assign layer0_outputs[3385] = inputs[154];
    assign layer0_outputs[3386] = ~(inputs[147]);
    assign layer0_outputs[3387] = 1'b1;
    assign layer0_outputs[3388] = 1'b0;
    assign layer0_outputs[3389] = 1'b1;
    assign layer0_outputs[3390] = ~((inputs[161]) | (inputs[162]));
    assign layer0_outputs[3391] = ~(inputs[129]);
    assign layer0_outputs[3392] = (inputs[173]) ^ (inputs[237]);
    assign layer0_outputs[3393] = 1'b0;
    assign layer0_outputs[3394] = (inputs[69]) | (inputs[25]);
    assign layer0_outputs[3395] = ~((inputs[100]) & (inputs[140]));
    assign layer0_outputs[3396] = ~((inputs[42]) ^ (inputs[13]));
    assign layer0_outputs[3397] = inputs[231];
    assign layer0_outputs[3398] = ~(inputs[183]);
    assign layer0_outputs[3399] = ~(inputs[230]) | (inputs[59]);
    assign layer0_outputs[3400] = ~((inputs[93]) & (inputs[79]));
    assign layer0_outputs[3401] = ~((inputs[8]) | (inputs[128]));
    assign layer0_outputs[3402] = (inputs[57]) & ~(inputs[102]);
    assign layer0_outputs[3403] = ~((inputs[96]) ^ (inputs[210]));
    assign layer0_outputs[3404] = ~((inputs[230]) | (inputs[82]));
    assign layer0_outputs[3405] = (inputs[163]) | (inputs[181]);
    assign layer0_outputs[3406] = ~((inputs[224]) & (inputs[217]));
    assign layer0_outputs[3407] = (inputs[171]) & ~(inputs[49]);
    assign layer0_outputs[3408] = (inputs[18]) ^ (inputs[0]);
    assign layer0_outputs[3409] = (inputs[228]) & ~(inputs[174]);
    assign layer0_outputs[3410] = (inputs[185]) | (inputs[181]);
    assign layer0_outputs[3411] = ~((inputs[86]) & (inputs[230]));
    assign layer0_outputs[3412] = (inputs[52]) & (inputs[23]);
    assign layer0_outputs[3413] = ~((inputs[28]) | (inputs[248]));
    assign layer0_outputs[3414] = 1'b0;
    assign layer0_outputs[3415] = (inputs[101]) | (inputs[197]);
    assign layer0_outputs[3416] = inputs[133];
    assign layer0_outputs[3417] = (inputs[110]) ^ (inputs[92]);
    assign layer0_outputs[3418] = (inputs[179]) | (inputs[6]);
    assign layer0_outputs[3419] = ~((inputs[217]) | (inputs[185]));
    assign layer0_outputs[3420] = (inputs[231]) & ~(inputs[92]);
    assign layer0_outputs[3421] = (inputs[208]) | (inputs[250]);
    assign layer0_outputs[3422] = (inputs[207]) | (inputs[238]);
    assign layer0_outputs[3423] = ~(inputs[85]) | (inputs[32]);
    assign layer0_outputs[3424] = inputs[77];
    assign layer0_outputs[3425] = (inputs[197]) ^ (inputs[39]);
    assign layer0_outputs[3426] = ~(inputs[48]) | (inputs[249]);
    assign layer0_outputs[3427] = (inputs[182]) & ~(inputs[77]);
    assign layer0_outputs[3428] = ~((inputs[228]) ^ (inputs[40]));
    assign layer0_outputs[3429] = ~((inputs[106]) | (inputs[180]));
    assign layer0_outputs[3430] = (inputs[217]) | (inputs[201]);
    assign layer0_outputs[3431] = inputs[13];
    assign layer0_outputs[3432] = ~(inputs[20]);
    assign layer0_outputs[3433] = ~(inputs[132]);
    assign layer0_outputs[3434] = ~(inputs[36]) | (inputs[226]);
    assign layer0_outputs[3435] = (inputs[179]) & ~(inputs[112]);
    assign layer0_outputs[3436] = (inputs[144]) ^ (inputs[230]);
    assign layer0_outputs[3437] = inputs[136];
    assign layer0_outputs[3438] = (inputs[80]) | (inputs[25]);
    assign layer0_outputs[3439] = inputs[19];
    assign layer0_outputs[3440] = 1'b1;
    assign layer0_outputs[3441] = ~(inputs[201]) | (inputs[115]);
    assign layer0_outputs[3442] = ~(inputs[7]);
    assign layer0_outputs[3443] = ~((inputs[64]) ^ (inputs[6]));
    assign layer0_outputs[3444] = ~(inputs[172]) | (inputs[2]);
    assign layer0_outputs[3445] = 1'b0;
    assign layer0_outputs[3446] = ~(inputs[7]) | (inputs[168]);
    assign layer0_outputs[3447] = (inputs[184]) | (inputs[97]);
    assign layer0_outputs[3448] = inputs[146];
    assign layer0_outputs[3449] = ~(inputs[167]) | (inputs[41]);
    assign layer0_outputs[3450] = (inputs[91]) | (inputs[77]);
    assign layer0_outputs[3451] = ~(inputs[34]);
    assign layer0_outputs[3452] = 1'b0;
    assign layer0_outputs[3453] = (inputs[40]) | (inputs[55]);
    assign layer0_outputs[3454] = inputs[139];
    assign layer0_outputs[3455] = (inputs[160]) & (inputs[82]);
    assign layer0_outputs[3456] = ~(inputs[254]);
    assign layer0_outputs[3457] = (inputs[165]) ^ (inputs[77]);
    assign layer0_outputs[3458] = (inputs[180]) & (inputs[184]);
    assign layer0_outputs[3459] = ~((inputs[134]) | (inputs[199]));
    assign layer0_outputs[3460] = (inputs[134]) & ~(inputs[113]);
    assign layer0_outputs[3461] = ~((inputs[52]) | (inputs[10]));
    assign layer0_outputs[3462] = (inputs[155]) | (inputs[233]);
    assign layer0_outputs[3463] = (inputs[19]) ^ (inputs[250]);
    assign layer0_outputs[3464] = (inputs[90]) & ~(inputs[174]);
    assign layer0_outputs[3465] = ~((inputs[117]) | (inputs[208]));
    assign layer0_outputs[3466] = ~(inputs[255]);
    assign layer0_outputs[3467] = (inputs[146]) & ~(inputs[31]);
    assign layer0_outputs[3468] = (inputs[226]) ^ (inputs[213]);
    assign layer0_outputs[3469] = (inputs[154]) & ~(inputs[25]);
    assign layer0_outputs[3470] = ~((inputs[29]) ^ (inputs[76]));
    assign layer0_outputs[3471] = inputs[113];
    assign layer0_outputs[3472] = 1'b1;
    assign layer0_outputs[3473] = (inputs[61]) | (inputs[39]);
    assign layer0_outputs[3474] = ~(inputs[219]) | (inputs[123]);
    assign layer0_outputs[3475] = ~(inputs[89]) | (inputs[135]);
    assign layer0_outputs[3476] = (inputs[10]) | (inputs[82]);
    assign layer0_outputs[3477] = ~((inputs[16]) | (inputs[3]));
    assign layer0_outputs[3478] = 1'b1;
    assign layer0_outputs[3479] = ~((inputs[84]) | (inputs[52]));
    assign layer0_outputs[3480] = ~((inputs[74]) ^ (inputs[222]));
    assign layer0_outputs[3481] = ~((inputs[73]) ^ (inputs[135]));
    assign layer0_outputs[3482] = ~(inputs[22]);
    assign layer0_outputs[3483] = (inputs[167]) & ~(inputs[189]);
    assign layer0_outputs[3484] = 1'b0;
    assign layer0_outputs[3485] = ~(inputs[120]);
    assign layer0_outputs[3486] = ~(inputs[195]) | (inputs[253]);
    assign layer0_outputs[3487] = ~(inputs[188]);
    assign layer0_outputs[3488] = (inputs[5]) ^ (inputs[125]);
    assign layer0_outputs[3489] = ~(inputs[228]);
    assign layer0_outputs[3490] = (inputs[167]) | (inputs[249]);
    assign layer0_outputs[3491] = ~(inputs[122]);
    assign layer0_outputs[3492] = (inputs[85]) ^ (inputs[23]);
    assign layer0_outputs[3493] = ~(inputs[72]) | (inputs[1]);
    assign layer0_outputs[3494] = 1'b0;
    assign layer0_outputs[3495] = ~(inputs[74]);
    assign layer0_outputs[3496] = (inputs[76]) | (inputs[94]);
    assign layer0_outputs[3497] = inputs[76];
    assign layer0_outputs[3498] = (inputs[197]) & (inputs[167]);
    assign layer0_outputs[3499] = ~((inputs[174]) | (inputs[99]));
    assign layer0_outputs[3500] = 1'b0;
    assign layer0_outputs[3501] = (inputs[130]) | (inputs[192]);
    assign layer0_outputs[3502] = ~((inputs[75]) | (inputs[9]));
    assign layer0_outputs[3503] = ~(inputs[189]);
    assign layer0_outputs[3504] = ~(inputs[130]) | (inputs[208]);
    assign layer0_outputs[3505] = ~(inputs[97]);
    assign layer0_outputs[3506] = ~(inputs[170]);
    assign layer0_outputs[3507] = ~((inputs[52]) & (inputs[110]));
    assign layer0_outputs[3508] = (inputs[136]) ^ (inputs[254]);
    assign layer0_outputs[3509] = ~(inputs[20]) | (inputs[99]);
    assign layer0_outputs[3510] = ~((inputs[130]) | (inputs[11]));
    assign layer0_outputs[3511] = (inputs[141]) & (inputs[20]);
    assign layer0_outputs[3512] = (inputs[54]) & ~(inputs[110]);
    assign layer0_outputs[3513] = ~(inputs[218]);
    assign layer0_outputs[3514] = ~(inputs[117]);
    assign layer0_outputs[3515] = ~(inputs[74]);
    assign layer0_outputs[3516] = 1'b0;
    assign layer0_outputs[3517] = (inputs[31]) & (inputs[27]);
    assign layer0_outputs[3518] = ~(inputs[40]);
    assign layer0_outputs[3519] = ~(inputs[72]) | (inputs[50]);
    assign layer0_outputs[3520] = ~((inputs[104]) ^ (inputs[62]));
    assign layer0_outputs[3521] = ~(inputs[6]) | (inputs[97]);
    assign layer0_outputs[3522] = ~(inputs[211]) | (inputs[1]);
    assign layer0_outputs[3523] = ~((inputs[48]) & (inputs[75]));
    assign layer0_outputs[3524] = inputs[98];
    assign layer0_outputs[3525] = (inputs[144]) ^ (inputs[204]);
    assign layer0_outputs[3526] = 1'b1;
    assign layer0_outputs[3527] = (inputs[117]) & ~(inputs[126]);
    assign layer0_outputs[3528] = (inputs[72]) & ~(inputs[13]);
    assign layer0_outputs[3529] = (inputs[16]) ^ (inputs[7]);
    assign layer0_outputs[3530] = (inputs[168]) ^ (inputs[15]);
    assign layer0_outputs[3531] = (inputs[245]) & (inputs[249]);
    assign layer0_outputs[3532] = (inputs[60]) & ~(inputs[38]);
    assign layer0_outputs[3533] = (inputs[55]) | (inputs[131]);
    assign layer0_outputs[3534] = inputs[89];
    assign layer0_outputs[3535] = ~((inputs[208]) | (inputs[24]));
    assign layer0_outputs[3536] = ~((inputs[51]) ^ (inputs[19]));
    assign layer0_outputs[3537] = (inputs[183]) & ~(inputs[186]);
    assign layer0_outputs[3538] = (inputs[5]) ^ (inputs[215]);
    assign layer0_outputs[3539] = inputs[78];
    assign layer0_outputs[3540] = ~((inputs[24]) | (inputs[8]));
    assign layer0_outputs[3541] = ~((inputs[88]) | (inputs[39]));
    assign layer0_outputs[3542] = ~((inputs[47]) | (inputs[22]));
    assign layer0_outputs[3543] = (inputs[214]) & ~(inputs[50]);
    assign layer0_outputs[3544] = (inputs[0]) ^ (inputs[145]);
    assign layer0_outputs[3545] = ~((inputs[193]) ^ (inputs[254]));
    assign layer0_outputs[3546] = (inputs[201]) ^ (inputs[191]);
    assign layer0_outputs[3547] = ~((inputs[33]) | (inputs[18]));
    assign layer0_outputs[3548] = ~(inputs[204]) | (inputs[154]);
    assign layer0_outputs[3549] = ~(inputs[103]);
    assign layer0_outputs[3550] = ~((inputs[53]) ^ (inputs[21]));
    assign layer0_outputs[3551] = ~(inputs[255]) | (inputs[59]);
    assign layer0_outputs[3552] = (inputs[34]) ^ (inputs[3]);
    assign layer0_outputs[3553] = (inputs[35]) & ~(inputs[59]);
    assign layer0_outputs[3554] = (inputs[21]) ^ (inputs[108]);
    assign layer0_outputs[3555] = (inputs[113]) ^ (inputs[5]);
    assign layer0_outputs[3556] = inputs[26];
    assign layer0_outputs[3557] = (inputs[151]) | (inputs[118]);
    assign layer0_outputs[3558] = (inputs[90]) & (inputs[115]);
    assign layer0_outputs[3559] = ~(inputs[52]) | (inputs[195]);
    assign layer0_outputs[3560] = (inputs[96]) | (inputs[94]);
    assign layer0_outputs[3561] = ~(inputs[117]);
    assign layer0_outputs[3562] = ~(inputs[93]);
    assign layer0_outputs[3563] = ~((inputs[180]) | (inputs[197]));
    assign layer0_outputs[3564] = ~((inputs[206]) ^ (inputs[114]));
    assign layer0_outputs[3565] = (inputs[238]) & (inputs[158]);
    assign layer0_outputs[3566] = ~((inputs[168]) | (inputs[170]));
    assign layer0_outputs[3567] = ~(inputs[23]);
    assign layer0_outputs[3568] = (inputs[29]) | (inputs[17]);
    assign layer0_outputs[3569] = ~(inputs[147]);
    assign layer0_outputs[3570] = inputs[49];
    assign layer0_outputs[3571] = (inputs[240]) & ~(inputs[29]);
    assign layer0_outputs[3572] = inputs[198];
    assign layer0_outputs[3573] = ~((inputs[146]) ^ (inputs[246]));
    assign layer0_outputs[3574] = (inputs[28]) | (inputs[5]);
    assign layer0_outputs[3575] = ~(inputs[41]) | (inputs[167]);
    assign layer0_outputs[3576] = 1'b0;
    assign layer0_outputs[3577] = inputs[188];
    assign layer0_outputs[3578] = ~(inputs[41]);
    assign layer0_outputs[3579] = (inputs[234]) | (inputs[168]);
    assign layer0_outputs[3580] = ~((inputs[204]) | (inputs[177]));
    assign layer0_outputs[3581] = (inputs[76]) & (inputs[9]);
    assign layer0_outputs[3582] = inputs[193];
    assign layer0_outputs[3583] = ~((inputs[52]) ^ (inputs[21]));
    assign layer0_outputs[3584] = ~(inputs[181]);
    assign layer0_outputs[3585] = ~(inputs[112]) | (inputs[111]);
    assign layer0_outputs[3586] = (inputs[70]) | (inputs[119]);
    assign layer0_outputs[3587] = inputs[21];
    assign layer0_outputs[3588] = (inputs[92]) & ~(inputs[207]);
    assign layer0_outputs[3589] = 1'b1;
    assign layer0_outputs[3590] = ~(inputs[154]);
    assign layer0_outputs[3591] = ~((inputs[63]) | (inputs[37]));
    assign layer0_outputs[3592] = ~((inputs[81]) & (inputs[138]));
    assign layer0_outputs[3593] = (inputs[176]) ^ (inputs[253]);
    assign layer0_outputs[3594] = inputs[30];
    assign layer0_outputs[3595] = ~((inputs[144]) | (inputs[170]));
    assign layer0_outputs[3596] = ~(inputs[41]) | (inputs[168]);
    assign layer0_outputs[3597] = ~(inputs[108]);
    assign layer0_outputs[3598] = 1'b0;
    assign layer0_outputs[3599] = (inputs[239]) | (inputs[36]);
    assign layer0_outputs[3600] = (inputs[167]) & (inputs[24]);
    assign layer0_outputs[3601] = inputs[27];
    assign layer0_outputs[3602] = inputs[63];
    assign layer0_outputs[3603] = (inputs[159]) | (inputs[232]);
    assign layer0_outputs[3604] = ~(inputs[125]) | (inputs[225]);
    assign layer0_outputs[3605] = (inputs[24]) | (inputs[250]);
    assign layer0_outputs[3606] = (inputs[104]) | (inputs[83]);
    assign layer0_outputs[3607] = inputs[237];
    assign layer0_outputs[3608] = ~(inputs[183]) | (inputs[113]);
    assign layer0_outputs[3609] = ~(inputs[20]);
    assign layer0_outputs[3610] = ~(inputs[11]);
    assign layer0_outputs[3611] = inputs[146];
    assign layer0_outputs[3612] = ~((inputs[146]) | (inputs[46]));
    assign layer0_outputs[3613] = (inputs[128]) & ~(inputs[171]);
    assign layer0_outputs[3614] = ~(inputs[253]) | (inputs[17]);
    assign layer0_outputs[3615] = (inputs[157]) | (inputs[236]);
    assign layer0_outputs[3616] = ~((inputs[142]) & (inputs[133]));
    assign layer0_outputs[3617] = inputs[15];
    assign layer0_outputs[3618] = ~((inputs[104]) & (inputs[46]));
    assign layer0_outputs[3619] = ~((inputs[89]) | (inputs[104]));
    assign layer0_outputs[3620] = ~((inputs[133]) & (inputs[232]));
    assign layer0_outputs[3621] = (inputs[139]) ^ (inputs[27]);
    assign layer0_outputs[3622] = ~((inputs[23]) & (inputs[230]));
    assign layer0_outputs[3623] = ~((inputs[150]) | (inputs[80]));
    assign layer0_outputs[3624] = ~(inputs[125]);
    assign layer0_outputs[3625] = inputs[144];
    assign layer0_outputs[3626] = (inputs[29]) | (inputs[156]);
    assign layer0_outputs[3627] = 1'b0;
    assign layer0_outputs[3628] = inputs[135];
    assign layer0_outputs[3629] = ~(inputs[9]);
    assign layer0_outputs[3630] = (inputs[120]) ^ (inputs[154]);
    assign layer0_outputs[3631] = ~((inputs[163]) | (inputs[140]));
    assign layer0_outputs[3632] = ~((inputs[71]) ^ (inputs[35]));
    assign layer0_outputs[3633] = ~((inputs[197]) | (inputs[213]));
    assign layer0_outputs[3634] = inputs[99];
    assign layer0_outputs[3635] = ~(inputs[228]) | (inputs[38]);
    assign layer0_outputs[3636] = (inputs[130]) | (inputs[50]);
    assign layer0_outputs[3637] = ~(inputs[80]);
    assign layer0_outputs[3638] = ~((inputs[13]) & (inputs[16]));
    assign layer0_outputs[3639] = (inputs[214]) | (inputs[158]);
    assign layer0_outputs[3640] = (inputs[153]) | (inputs[18]);
    assign layer0_outputs[3641] = (inputs[37]) & (inputs[44]);
    assign layer0_outputs[3642] = ~(inputs[56]);
    assign layer0_outputs[3643] = (inputs[83]) ^ (inputs[127]);
    assign layer0_outputs[3644] = inputs[231];
    assign layer0_outputs[3645] = ~(inputs[130]) | (inputs[154]);
    assign layer0_outputs[3646] = inputs[216];
    assign layer0_outputs[3647] = (inputs[155]) | (inputs[13]);
    assign layer0_outputs[3648] = ~((inputs[69]) | (inputs[60]));
    assign layer0_outputs[3649] = ~((inputs[124]) & (inputs[165]));
    assign layer0_outputs[3650] = ~((inputs[222]) | (inputs[182]));
    assign layer0_outputs[3651] = inputs[148];
    assign layer0_outputs[3652] = inputs[91];
    assign layer0_outputs[3653] = (inputs[236]) | (inputs[88]);
    assign layer0_outputs[3654] = ~(inputs[172]) | (inputs[66]);
    assign layer0_outputs[3655] = (inputs[51]) & ~(inputs[41]);
    assign layer0_outputs[3656] = ~(inputs[112]) | (inputs[252]);
    assign layer0_outputs[3657] = inputs[193];
    assign layer0_outputs[3658] = (inputs[243]) | (inputs[71]);
    assign layer0_outputs[3659] = ~(inputs[131]);
    assign layer0_outputs[3660] = inputs[138];
    assign layer0_outputs[3661] = (inputs[211]) ^ (inputs[47]);
    assign layer0_outputs[3662] = ~((inputs[120]) | (inputs[118]));
    assign layer0_outputs[3663] = (inputs[17]) | (inputs[172]);
    assign layer0_outputs[3664] = inputs[204];
    assign layer0_outputs[3665] = ~(inputs[136]);
    assign layer0_outputs[3666] = ~(inputs[15]);
    assign layer0_outputs[3667] = (inputs[145]) | (inputs[222]);
    assign layer0_outputs[3668] = ~(inputs[38]) | (inputs[130]);
    assign layer0_outputs[3669] = ~(inputs[137]) | (inputs[10]);
    assign layer0_outputs[3670] = (inputs[20]) | (inputs[220]);
    assign layer0_outputs[3671] = ~(inputs[147]);
    assign layer0_outputs[3672] = ~(inputs[162]) | (inputs[33]);
    assign layer0_outputs[3673] = (inputs[49]) & (inputs[80]);
    assign layer0_outputs[3674] = ~(inputs[227]);
    assign layer0_outputs[3675] = (inputs[70]) & (inputs[71]);
    assign layer0_outputs[3676] = 1'b1;
    assign layer0_outputs[3677] = 1'b0;
    assign layer0_outputs[3678] = ~(inputs[155]) | (inputs[167]);
    assign layer0_outputs[3679] = inputs[103];
    assign layer0_outputs[3680] = ~(inputs[13]) | (inputs[233]);
    assign layer0_outputs[3681] = ~(inputs[135]);
    assign layer0_outputs[3682] = ~(inputs[38]) | (inputs[46]);
    assign layer0_outputs[3683] = inputs[74];
    assign layer0_outputs[3684] = (inputs[74]) & ~(inputs[53]);
    assign layer0_outputs[3685] = inputs[98];
    assign layer0_outputs[3686] = ~(inputs[240]);
    assign layer0_outputs[3687] = ~((inputs[6]) & (inputs[73]));
    assign layer0_outputs[3688] = ~(inputs[43]) | (inputs[167]);
    assign layer0_outputs[3689] = (inputs[61]) & ~(inputs[96]);
    assign layer0_outputs[3690] = inputs[238];
    assign layer0_outputs[3691] = (inputs[226]) & ~(inputs[86]);
    assign layer0_outputs[3692] = 1'b1;
    assign layer0_outputs[3693] = inputs[123];
    assign layer0_outputs[3694] = ~((inputs[193]) | (inputs[249]));
    assign layer0_outputs[3695] = (inputs[82]) | (inputs[116]);
    assign layer0_outputs[3696] = (inputs[195]) & ~(inputs[33]);
    assign layer0_outputs[3697] = inputs[66];
    assign layer0_outputs[3698] = inputs[193];
    assign layer0_outputs[3699] = ~((inputs[37]) ^ (inputs[28]));
    assign layer0_outputs[3700] = inputs[136];
    assign layer0_outputs[3701] = 1'b1;
    assign layer0_outputs[3702] = ~((inputs[244]) ^ (inputs[182]));
    assign layer0_outputs[3703] = ~((inputs[175]) | (inputs[184]));
    assign layer0_outputs[3704] = (inputs[151]) | (inputs[71]);
    assign layer0_outputs[3705] = (inputs[33]) & ~(inputs[110]);
    assign layer0_outputs[3706] = (inputs[49]) ^ (inputs[18]);
    assign layer0_outputs[3707] = inputs[137];
    assign layer0_outputs[3708] = (inputs[203]) & ~(inputs[29]);
    assign layer0_outputs[3709] = ~((inputs[238]) | (inputs[91]));
    assign layer0_outputs[3710] = ~((inputs[211]) & (inputs[211]));
    assign layer0_outputs[3711] = (inputs[11]) & ~(inputs[172]);
    assign layer0_outputs[3712] = (inputs[138]) & ~(inputs[192]);
    assign layer0_outputs[3713] = ~((inputs[142]) & (inputs[250]));
    assign layer0_outputs[3714] = ~(inputs[152]);
    assign layer0_outputs[3715] = 1'b1;
    assign layer0_outputs[3716] = (inputs[149]) & ~(inputs[41]);
    assign layer0_outputs[3717] = (inputs[61]) & ~(inputs[113]);
    assign layer0_outputs[3718] = 1'b1;
    assign layer0_outputs[3719] = ~(inputs[40]) | (inputs[178]);
    assign layer0_outputs[3720] = ~(inputs[250]) | (inputs[140]);
    assign layer0_outputs[3721] = ~(inputs[154]);
    assign layer0_outputs[3722] = inputs[82];
    assign layer0_outputs[3723] = (inputs[176]) ^ (inputs[83]);
    assign layer0_outputs[3724] = (inputs[80]) | (inputs[165]);
    assign layer0_outputs[3725] = (inputs[177]) & ~(inputs[51]);
    assign layer0_outputs[3726] = ~(inputs[177]);
    assign layer0_outputs[3727] = ~(inputs[148]);
    assign layer0_outputs[3728] = ~((inputs[32]) ^ (inputs[51]));
    assign layer0_outputs[3729] = (inputs[249]) & ~(inputs[20]);
    assign layer0_outputs[3730] = inputs[121];
    assign layer0_outputs[3731] = ~((inputs[20]) & (inputs[185]));
    assign layer0_outputs[3732] = (inputs[28]) & (inputs[111]);
    assign layer0_outputs[3733] = ~((inputs[202]) & (inputs[215]));
    assign layer0_outputs[3734] = ~((inputs[43]) ^ (inputs[70]));
    assign layer0_outputs[3735] = 1'b0;
    assign layer0_outputs[3736] = (inputs[163]) & (inputs[131]);
    assign layer0_outputs[3737] = (inputs[135]) & ~(inputs[195]);
    assign layer0_outputs[3738] = (inputs[165]) & (inputs[6]);
    assign layer0_outputs[3739] = (inputs[64]) | (inputs[241]);
    assign layer0_outputs[3740] = ~(inputs[28]);
    assign layer0_outputs[3741] = ~(inputs[112]);
    assign layer0_outputs[3742] = 1'b1;
    assign layer0_outputs[3743] = ~((inputs[25]) ^ (inputs[73]));
    assign layer0_outputs[3744] = ~((inputs[171]) & (inputs[132]));
    assign layer0_outputs[3745] = ~(inputs[167]);
    assign layer0_outputs[3746] = ~(inputs[26]) | (inputs[254]);
    assign layer0_outputs[3747] = inputs[75];
    assign layer0_outputs[3748] = ~(inputs[197]);
    assign layer0_outputs[3749] = (inputs[60]) & ~(inputs[222]);
    assign layer0_outputs[3750] = ~((inputs[161]) | (inputs[79]));
    assign layer0_outputs[3751] = (inputs[25]) ^ (inputs[231]);
    assign layer0_outputs[3752] = ~((inputs[156]) | (inputs[220]));
    assign layer0_outputs[3753] = ~(inputs[180]);
    assign layer0_outputs[3754] = (inputs[113]) | (inputs[200]);
    assign layer0_outputs[3755] = (inputs[76]) | (inputs[147]);
    assign layer0_outputs[3756] = (inputs[42]) | (inputs[158]);
    assign layer0_outputs[3757] = (inputs[179]) & ~(inputs[123]);
    assign layer0_outputs[3758] = (inputs[155]) & (inputs[154]);
    assign layer0_outputs[3759] = ~(inputs[253]);
    assign layer0_outputs[3760] = ~((inputs[238]) | (inputs[169]));
    assign layer0_outputs[3761] = 1'b1;
    assign layer0_outputs[3762] = ~(inputs[63]) | (inputs[180]);
    assign layer0_outputs[3763] = ~(inputs[188]) | (inputs[223]);
    assign layer0_outputs[3764] = ~((inputs[184]) | (inputs[2]));
    assign layer0_outputs[3765] = ~(inputs[22]);
    assign layer0_outputs[3766] = (inputs[122]) & ~(inputs[227]);
    assign layer0_outputs[3767] = inputs[123];
    assign layer0_outputs[3768] = inputs[211];
    assign layer0_outputs[3769] = inputs[167];
    assign layer0_outputs[3770] = ~(inputs[193]) | (inputs[93]);
    assign layer0_outputs[3771] = inputs[104];
    assign layer0_outputs[3772] = ~((inputs[6]) ^ (inputs[34]));
    assign layer0_outputs[3773] = ~(inputs[61]) | (inputs[144]);
    assign layer0_outputs[3774] = (inputs[18]) | (inputs[38]);
    assign layer0_outputs[3775] = (inputs[222]) & ~(inputs[38]);
    assign layer0_outputs[3776] = (inputs[144]) | (inputs[87]);
    assign layer0_outputs[3777] = ~(inputs[80]);
    assign layer0_outputs[3778] = inputs[124];
    assign layer0_outputs[3779] = ~(inputs[174]);
    assign layer0_outputs[3780] = (inputs[163]) ^ (inputs[145]);
    assign layer0_outputs[3781] = inputs[118];
    assign layer0_outputs[3782] = inputs[204];
    assign layer0_outputs[3783] = (inputs[8]) & ~(inputs[99]);
    assign layer0_outputs[3784] = (inputs[49]) ^ (inputs[152]);
    assign layer0_outputs[3785] = ~(inputs[39]) | (inputs[29]);
    assign layer0_outputs[3786] = 1'b0;
    assign layer0_outputs[3787] = ~(inputs[114]);
    assign layer0_outputs[3788] = ~((inputs[99]) ^ (inputs[62]));
    assign layer0_outputs[3789] = ~(inputs[245]) | (inputs[167]);
    assign layer0_outputs[3790] = inputs[145];
    assign layer0_outputs[3791] = (inputs[101]) & (inputs[49]);
    assign layer0_outputs[3792] = ~((inputs[50]) | (inputs[87]));
    assign layer0_outputs[3793] = (inputs[195]) & ~(inputs[63]);
    assign layer0_outputs[3794] = ~((inputs[150]) & (inputs[67]));
    assign layer0_outputs[3795] = ~((inputs[125]) | (inputs[139]));
    assign layer0_outputs[3796] = (inputs[230]) | (inputs[245]);
    assign layer0_outputs[3797] = ~((inputs[190]) ^ (inputs[107]));
    assign layer0_outputs[3798] = ~(inputs[176]);
    assign layer0_outputs[3799] = (inputs[170]) & ~(inputs[113]);
    assign layer0_outputs[3800] = ~(inputs[189]) | (inputs[216]);
    assign layer0_outputs[3801] = ~(inputs[101]) | (inputs[194]);
    assign layer0_outputs[3802] = ~(inputs[239]) | (inputs[160]);
    assign layer0_outputs[3803] = ~((inputs[144]) | (inputs[186]));
    assign layer0_outputs[3804] = (inputs[85]) & ~(inputs[1]);
    assign layer0_outputs[3805] = ~(inputs[83]);
    assign layer0_outputs[3806] = ~((inputs[156]) ^ (inputs[29]));
    assign layer0_outputs[3807] = inputs[105];
    assign layer0_outputs[3808] = (inputs[161]) & ~(inputs[44]);
    assign layer0_outputs[3809] = ~(inputs[251]) | (inputs[49]);
    assign layer0_outputs[3810] = ~(inputs[101]) | (inputs[172]);
    assign layer0_outputs[3811] = ~((inputs[33]) | (inputs[122]));
    assign layer0_outputs[3812] = ~((inputs[28]) & (inputs[69]));
    assign layer0_outputs[3813] = 1'b1;
    assign layer0_outputs[3814] = ~((inputs[199]) ^ (inputs[8]));
    assign layer0_outputs[3815] = ~(inputs[90]);
    assign layer0_outputs[3816] = (inputs[89]) | (inputs[211]);
    assign layer0_outputs[3817] = ~((inputs[15]) | (inputs[249]));
    assign layer0_outputs[3818] = ~((inputs[96]) ^ (inputs[86]));
    assign layer0_outputs[3819] = ~((inputs[29]) | (inputs[44]));
    assign layer0_outputs[3820] = ~(inputs[198]);
    assign layer0_outputs[3821] = ~((inputs[181]) & (inputs[116]));
    assign layer0_outputs[3822] = inputs[34];
    assign layer0_outputs[3823] = (inputs[235]) ^ (inputs[209]);
    assign layer0_outputs[3824] = (inputs[42]) & (inputs[23]);
    assign layer0_outputs[3825] = (inputs[150]) & ~(inputs[234]);
    assign layer0_outputs[3826] = (inputs[214]) & ~(inputs[64]);
    assign layer0_outputs[3827] = (inputs[231]) & ~(inputs[90]);
    assign layer0_outputs[3828] = inputs[78];
    assign layer0_outputs[3829] = ~(inputs[21]) | (inputs[114]);
    assign layer0_outputs[3830] = ~((inputs[239]) & (inputs[207]));
    assign layer0_outputs[3831] = ~((inputs[248]) ^ (inputs[218]));
    assign layer0_outputs[3832] = inputs[155];
    assign layer0_outputs[3833] = (inputs[103]) & ~(inputs[63]);
    assign layer0_outputs[3834] = ~((inputs[56]) & (inputs[19]));
    assign layer0_outputs[3835] = 1'b1;
    assign layer0_outputs[3836] = (inputs[52]) & ~(inputs[219]);
    assign layer0_outputs[3837] = 1'b1;
    assign layer0_outputs[3838] = ~(inputs[150]) | (inputs[55]);
    assign layer0_outputs[3839] = ~(inputs[219]) | (inputs[29]);
    assign layer0_outputs[3840] = ~(inputs[110]);
    assign layer0_outputs[3841] = (inputs[153]) & ~(inputs[56]);
    assign layer0_outputs[3842] = ~(inputs[163]);
    assign layer0_outputs[3843] = inputs[67];
    assign layer0_outputs[3844] = inputs[131];
    assign layer0_outputs[3845] = (inputs[141]) | (inputs[122]);
    assign layer0_outputs[3846] = ~(inputs[207]) | (inputs[122]);
    assign layer0_outputs[3847] = (inputs[4]) | (inputs[31]);
    assign layer0_outputs[3848] = (inputs[228]) & ~(inputs[142]);
    assign layer0_outputs[3849] = (inputs[165]) & ~(inputs[165]);
    assign layer0_outputs[3850] = (inputs[203]) | (inputs[255]);
    assign layer0_outputs[3851] = 1'b1;
    assign layer0_outputs[3852] = ~(inputs[122]) | (inputs[56]);
    assign layer0_outputs[3853] = ~(inputs[183]);
    assign layer0_outputs[3854] = ~(inputs[119]);
    assign layer0_outputs[3855] = (inputs[154]) & ~(inputs[204]);
    assign layer0_outputs[3856] = ~(inputs[92]) | (inputs[40]);
    assign layer0_outputs[3857] = ~(inputs[164]);
    assign layer0_outputs[3858] = ~((inputs[35]) & (inputs[38]));
    assign layer0_outputs[3859] = ~(inputs[219]) | (inputs[237]);
    assign layer0_outputs[3860] = ~(inputs[164]) | (inputs[254]);
    assign layer0_outputs[3861] = ~((inputs[151]) | (inputs[15]));
    assign layer0_outputs[3862] = (inputs[130]) & ~(inputs[240]);
    assign layer0_outputs[3863] = inputs[237];
    assign layer0_outputs[3864] = (inputs[207]) & ~(inputs[32]);
    assign layer0_outputs[3865] = ~(inputs[47]) | (inputs[205]);
    assign layer0_outputs[3866] = ~(inputs[32]);
    assign layer0_outputs[3867] = inputs[60];
    assign layer0_outputs[3868] = inputs[194];
    assign layer0_outputs[3869] = ~(inputs[138]) | (inputs[31]);
    assign layer0_outputs[3870] = ~((inputs[170]) | (inputs[88]));
    assign layer0_outputs[3871] = (inputs[14]) & ~(inputs[239]);
    assign layer0_outputs[3872] = inputs[75];
    assign layer0_outputs[3873] = ~((inputs[80]) ^ (inputs[103]));
    assign layer0_outputs[3874] = ~(inputs[9]);
    assign layer0_outputs[3875] = inputs[25];
    assign layer0_outputs[3876] = 1'b1;
    assign layer0_outputs[3877] = ~(inputs[168]);
    assign layer0_outputs[3878] = (inputs[43]) & ~(inputs[101]);
    assign layer0_outputs[3879] = ~(inputs[45]);
    assign layer0_outputs[3880] = inputs[213];
    assign layer0_outputs[3881] = inputs[69];
    assign layer0_outputs[3882] = (inputs[151]) & ~(inputs[156]);
    assign layer0_outputs[3883] = ~(inputs[135]);
    assign layer0_outputs[3884] = (inputs[239]) ^ (inputs[89]);
    assign layer0_outputs[3885] = (inputs[22]) | (inputs[37]);
    assign layer0_outputs[3886] = ~((inputs[242]) | (inputs[2]));
    assign layer0_outputs[3887] = (inputs[9]) & ~(inputs[205]);
    assign layer0_outputs[3888] = ~((inputs[52]) | (inputs[26]));
    assign layer0_outputs[3889] = 1'b0;
    assign layer0_outputs[3890] = (inputs[40]) & ~(inputs[129]);
    assign layer0_outputs[3891] = ~(inputs[100]);
    assign layer0_outputs[3892] = ~(inputs[52]);
    assign layer0_outputs[3893] = ~((inputs[119]) ^ (inputs[89]));
    assign layer0_outputs[3894] = ~((inputs[187]) | (inputs[122]));
    assign layer0_outputs[3895] = ~(inputs[44]);
    assign layer0_outputs[3896] = (inputs[120]) & ~(inputs[19]);
    assign layer0_outputs[3897] = (inputs[248]) & (inputs[234]);
    assign layer0_outputs[3898] = ~(inputs[105]) | (inputs[8]);
    assign layer0_outputs[3899] = (inputs[132]) | (inputs[122]);
    assign layer0_outputs[3900] = ~(inputs[91]) | (inputs[87]);
    assign layer0_outputs[3901] = (inputs[240]) & (inputs[142]);
    assign layer0_outputs[3902] = inputs[36];
    assign layer0_outputs[3903] = (inputs[163]) & ~(inputs[142]);
    assign layer0_outputs[3904] = (inputs[196]) & (inputs[74]);
    assign layer0_outputs[3905] = ~(inputs[147]) | (inputs[109]);
    assign layer0_outputs[3906] = ~((inputs[118]) | (inputs[117]));
    assign layer0_outputs[3907] = ~(inputs[17]);
    assign layer0_outputs[3908] = (inputs[72]) & ~(inputs[186]);
    assign layer0_outputs[3909] = (inputs[129]) | (inputs[75]);
    assign layer0_outputs[3910] = ~(inputs[153]) | (inputs[40]);
    assign layer0_outputs[3911] = inputs[108];
    assign layer0_outputs[3912] = ~((inputs[175]) | (inputs[158]));
    assign layer0_outputs[3913] = ~((inputs[62]) | (inputs[192]));
    assign layer0_outputs[3914] = inputs[154];
    assign layer0_outputs[3915] = (inputs[37]) | (inputs[52]);
    assign layer0_outputs[3916] = (inputs[66]) | (inputs[210]);
    assign layer0_outputs[3917] = ~((inputs[37]) | (inputs[84]));
    assign layer0_outputs[3918] = ~(inputs[194]) | (inputs[96]);
    assign layer0_outputs[3919] = ~(inputs[177]);
    assign layer0_outputs[3920] = inputs[199];
    assign layer0_outputs[3921] = ~((inputs[93]) | (inputs[47]));
    assign layer0_outputs[3922] = (inputs[27]) | (inputs[12]);
    assign layer0_outputs[3923] = (inputs[36]) ^ (inputs[22]);
    assign layer0_outputs[3924] = 1'b1;
    assign layer0_outputs[3925] = (inputs[150]) | (inputs[250]);
    assign layer0_outputs[3926] = inputs[204];
    assign layer0_outputs[3927] = (inputs[47]) ^ (inputs[55]);
    assign layer0_outputs[3928] = (inputs[5]) & ~(inputs[159]);
    assign layer0_outputs[3929] = 1'b1;
    assign layer0_outputs[3930] = ~(inputs[101]);
    assign layer0_outputs[3931] = (inputs[204]) & ~(inputs[240]);
    assign layer0_outputs[3932] = (inputs[224]) & ~(inputs[238]);
    assign layer0_outputs[3933] = ~((inputs[176]) ^ (inputs[111]));
    assign layer0_outputs[3934] = ~(inputs[166]);
    assign layer0_outputs[3935] = inputs[43];
    assign layer0_outputs[3936] = ~(inputs[121]);
    assign layer0_outputs[3937] = (inputs[231]) ^ (inputs[199]);
    assign layer0_outputs[3938] = inputs[220];
    assign layer0_outputs[3939] = (inputs[130]) & ~(inputs[162]);
    assign layer0_outputs[3940] = ~(inputs[238]) | (inputs[15]);
    assign layer0_outputs[3941] = ~(inputs[117]);
    assign layer0_outputs[3942] = ~((inputs[195]) ^ (inputs[227]));
    assign layer0_outputs[3943] = 1'b1;
    assign layer0_outputs[3944] = inputs[69];
    assign layer0_outputs[3945] = ~(inputs[129]);
    assign layer0_outputs[3946] = ~((inputs[90]) | (inputs[80]));
    assign layer0_outputs[3947] = 1'b1;
    assign layer0_outputs[3948] = ~(inputs[37]);
    assign layer0_outputs[3949] = (inputs[115]) & ~(inputs[239]);
    assign layer0_outputs[3950] = ~(inputs[82]) | (inputs[82]);
    assign layer0_outputs[3951] = (inputs[219]) & ~(inputs[142]);
    assign layer0_outputs[3952] = 1'b1;
    assign layer0_outputs[3953] = ~(inputs[39]) | (inputs[241]);
    assign layer0_outputs[3954] = (inputs[107]) & (inputs[228]);
    assign layer0_outputs[3955] = (inputs[152]) | (inputs[245]);
    assign layer0_outputs[3956] = inputs[56];
    assign layer0_outputs[3957] = inputs[194];
    assign layer0_outputs[3958] = (inputs[9]) & ~(inputs[15]);
    assign layer0_outputs[3959] = (inputs[142]) & (inputs[186]);
    assign layer0_outputs[3960] = ~((inputs[231]) ^ (inputs[13]));
    assign layer0_outputs[3961] = inputs[175];
    assign layer0_outputs[3962] = (inputs[94]) ^ (inputs[178]);
    assign layer0_outputs[3963] = ~((inputs[176]) | (inputs[109]));
    assign layer0_outputs[3964] = ~((inputs[74]) & (inputs[69]));
    assign layer0_outputs[3965] = (inputs[232]) | (inputs[11]);
    assign layer0_outputs[3966] = ~(inputs[11]);
    assign layer0_outputs[3967] = ~((inputs[101]) | (inputs[235]));
    assign layer0_outputs[3968] = inputs[181];
    assign layer0_outputs[3969] = (inputs[115]) & ~(inputs[226]);
    assign layer0_outputs[3970] = ~(inputs[39]);
    assign layer0_outputs[3971] = (inputs[50]) | (inputs[187]);
    assign layer0_outputs[3972] = ~((inputs[252]) | (inputs[234]));
    assign layer0_outputs[3973] = ~(inputs[139]) | (inputs[13]);
    assign layer0_outputs[3974] = ~((inputs[39]) | (inputs[0]));
    assign layer0_outputs[3975] = ~((inputs[204]) ^ (inputs[241]));
    assign layer0_outputs[3976] = (inputs[87]) & ~(inputs[238]);
    assign layer0_outputs[3977] = inputs[83];
    assign layer0_outputs[3978] = ~((inputs[196]) | (inputs[167]));
    assign layer0_outputs[3979] = ~(inputs[181]);
    assign layer0_outputs[3980] = ~(inputs[220]);
    assign layer0_outputs[3981] = ~(inputs[69]);
    assign layer0_outputs[3982] = inputs[75];
    assign layer0_outputs[3983] = inputs[57];
    assign layer0_outputs[3984] = ~((inputs[241]) | (inputs[147]));
    assign layer0_outputs[3985] = inputs[79];
    assign layer0_outputs[3986] = ~(inputs[97]);
    assign layer0_outputs[3987] = (inputs[243]) | (inputs[159]);
    assign layer0_outputs[3988] = ~(inputs[208]);
    assign layer0_outputs[3989] = ~((inputs[201]) ^ (inputs[179]));
    assign layer0_outputs[3990] = ~(inputs[172]);
    assign layer0_outputs[3991] = 1'b1;
    assign layer0_outputs[3992] = 1'b0;
    assign layer0_outputs[3993] = (inputs[185]) & ~(inputs[225]);
    assign layer0_outputs[3994] = (inputs[128]) & ~(inputs[213]);
    assign layer0_outputs[3995] = ~((inputs[201]) & (inputs[215]));
    assign layer0_outputs[3996] = inputs[59];
    assign layer0_outputs[3997] = (inputs[179]) & ~(inputs[97]);
    assign layer0_outputs[3998] = ~((inputs[197]) | (inputs[249]));
    assign layer0_outputs[3999] = ~((inputs[208]) | (inputs[197]));
    assign layer0_outputs[4000] = (inputs[128]) | (inputs[37]);
    assign layer0_outputs[4001] = (inputs[116]) ^ (inputs[66]);
    assign layer0_outputs[4002] = (inputs[157]) & ~(inputs[58]);
    assign layer0_outputs[4003] = (inputs[229]) ^ (inputs[0]);
    assign layer0_outputs[4004] = ~(inputs[156]);
    assign layer0_outputs[4005] = (inputs[178]) | (inputs[198]);
    assign layer0_outputs[4006] = (inputs[253]) & ~(inputs[181]);
    assign layer0_outputs[4007] = (inputs[104]) & ~(inputs[160]);
    assign layer0_outputs[4008] = ~(inputs[7]) | (inputs[159]);
    assign layer0_outputs[4009] = ~(inputs[89]) | (inputs[239]);
    assign layer0_outputs[4010] = ~((inputs[21]) | (inputs[90]));
    assign layer0_outputs[4011] = ~((inputs[94]) ^ (inputs[175]));
    assign layer0_outputs[4012] = inputs[160];
    assign layer0_outputs[4013] = (inputs[205]) & (inputs[253]);
    assign layer0_outputs[4014] = (inputs[249]) ^ (inputs[247]);
    assign layer0_outputs[4015] = inputs[26];
    assign layer0_outputs[4016] = ~((inputs[213]) ^ (inputs[241]));
    assign layer0_outputs[4017] = ~((inputs[128]) ^ (inputs[171]));
    assign layer0_outputs[4018] = ~((inputs[102]) | (inputs[205]));
    assign layer0_outputs[4019] = ~((inputs[21]) ^ (inputs[229]));
    assign layer0_outputs[4020] = inputs[2];
    assign layer0_outputs[4021] = (inputs[128]) & (inputs[47]);
    assign layer0_outputs[4022] = ~(inputs[109]);
    assign layer0_outputs[4023] = (inputs[131]) ^ (inputs[131]);
    assign layer0_outputs[4024] = ~((inputs[229]) | (inputs[65]));
    assign layer0_outputs[4025] = ~((inputs[89]) | (inputs[136]));
    assign layer0_outputs[4026] = ~(inputs[160]);
    assign layer0_outputs[4027] = (inputs[6]) | (inputs[195]);
    assign layer0_outputs[4028] = (inputs[223]) & ~(inputs[143]);
    assign layer0_outputs[4029] = inputs[183];
    assign layer0_outputs[4030] = ~((inputs[217]) & (inputs[80]));
    assign layer0_outputs[4031] = ~((inputs[66]) | (inputs[153]));
    assign layer0_outputs[4032] = ~((inputs[112]) | (inputs[210]));
    assign layer0_outputs[4033] = ~((inputs[248]) ^ (inputs[216]));
    assign layer0_outputs[4034] = inputs[22];
    assign layer0_outputs[4035] = ~((inputs[49]) | (inputs[90]));
    assign layer0_outputs[4036] = 1'b1;
    assign layer0_outputs[4037] = inputs[51];
    assign layer0_outputs[4038] = ~(inputs[149]);
    assign layer0_outputs[4039] = ~(inputs[152]) | (inputs[130]);
    assign layer0_outputs[4040] = ~((inputs[149]) ^ (inputs[87]));
    assign layer0_outputs[4041] = ~((inputs[125]) & (inputs[152]));
    assign layer0_outputs[4042] = ~(inputs[119]);
    assign layer0_outputs[4043] = (inputs[66]) | (inputs[141]);
    assign layer0_outputs[4044] = ~(inputs[27]) | (inputs[221]);
    assign layer0_outputs[4045] = 1'b0;
    assign layer0_outputs[4046] = (inputs[208]) | (inputs[74]);
    assign layer0_outputs[4047] = (inputs[18]) & ~(inputs[103]);
    assign layer0_outputs[4048] = (inputs[102]) & (inputs[145]);
    assign layer0_outputs[4049] = (inputs[103]) & ~(inputs[68]);
    assign layer0_outputs[4050] = (inputs[23]) | (inputs[141]);
    assign layer0_outputs[4051] = (inputs[32]) & ~(inputs[29]);
    assign layer0_outputs[4052] = ~(inputs[183]) | (inputs[192]);
    assign layer0_outputs[4053] = ~(inputs[47]);
    assign layer0_outputs[4054] = ~(inputs[184]);
    assign layer0_outputs[4055] = 1'b1;
    assign layer0_outputs[4056] = inputs[195];
    assign layer0_outputs[4057] = ~(inputs[177]);
    assign layer0_outputs[4058] = ~((inputs[63]) | (inputs[51]));
    assign layer0_outputs[4059] = inputs[235];
    assign layer0_outputs[4060] = ~((inputs[195]) | (inputs[43]));
    assign layer0_outputs[4061] = ~(inputs[149]);
    assign layer0_outputs[4062] = (inputs[252]) | (inputs[148]);
    assign layer0_outputs[4063] = 1'b1;
    assign layer0_outputs[4064] = (inputs[33]) | (inputs[122]);
    assign layer0_outputs[4065] = ~(inputs[100]);
    assign layer0_outputs[4066] = ~(inputs[55]) | (inputs[73]);
    assign layer0_outputs[4067] = inputs[160];
    assign layer0_outputs[4068] = ~(inputs[178]) | (inputs[166]);
    assign layer0_outputs[4069] = ~(inputs[167]);
    assign layer0_outputs[4070] = ~(inputs[160]);
    assign layer0_outputs[4071] = 1'b0;
    assign layer0_outputs[4072] = ~(inputs[109]) | (inputs[33]);
    assign layer0_outputs[4073] = ~((inputs[137]) | (inputs[64]));
    assign layer0_outputs[4074] = inputs[10];
    assign layer0_outputs[4075] = ~(inputs[34]);
    assign layer0_outputs[4076] = ~(inputs[104]) | (inputs[58]);
    assign layer0_outputs[4077] = (inputs[246]) | (inputs[81]);
    assign layer0_outputs[4078] = inputs[33];
    assign layer0_outputs[4079] = ~(inputs[35]);
    assign layer0_outputs[4080] = (inputs[147]) & (inputs[163]);
    assign layer0_outputs[4081] = ~(inputs[247]);
    assign layer0_outputs[4082] = ~((inputs[142]) ^ (inputs[86]));
    assign layer0_outputs[4083] = inputs[217];
    assign layer0_outputs[4084] = (inputs[40]) & ~(inputs[242]);
    assign layer0_outputs[4085] = ~(inputs[210]);
    assign layer0_outputs[4086] = (inputs[105]) & ~(inputs[250]);
    assign layer0_outputs[4087] = (inputs[210]) | (inputs[217]);
    assign layer0_outputs[4088] = inputs[169];
    assign layer0_outputs[4089] = ~((inputs[74]) ^ (inputs[6]));
    assign layer0_outputs[4090] = ~(inputs[242]) | (inputs[94]);
    assign layer0_outputs[4091] = ~(inputs[205]) | (inputs[6]);
    assign layer0_outputs[4092] = (inputs[53]) & ~(inputs[227]);
    assign layer0_outputs[4093] = ~(inputs[44]);
    assign layer0_outputs[4094] = (inputs[194]) & ~(inputs[129]);
    assign layer0_outputs[4095] = ~((inputs[196]) | (inputs[71]));
    assign layer0_outputs[4096] = ~(inputs[131]);
    assign layer0_outputs[4097] = (inputs[154]) | (inputs[71]);
    assign layer0_outputs[4098] = (inputs[72]) | (inputs[204]);
    assign layer0_outputs[4099] = (inputs[245]) | (inputs[173]);
    assign layer0_outputs[4100] = ~(inputs[27]) | (inputs[119]);
    assign layer0_outputs[4101] = inputs[245];
    assign layer0_outputs[4102] = inputs[40];
    assign layer0_outputs[4103] = (inputs[20]) & ~(inputs[137]);
    assign layer0_outputs[4104] = ~((inputs[237]) ^ (inputs[69]));
    assign layer0_outputs[4105] = (inputs[35]) & (inputs[243]);
    assign layer0_outputs[4106] = (inputs[254]) | (inputs[8]);
    assign layer0_outputs[4107] = (inputs[175]) & ~(inputs[114]);
    assign layer0_outputs[4108] = (inputs[165]) | (inputs[17]);
    assign layer0_outputs[4109] = ~(inputs[44]);
    assign layer0_outputs[4110] = (inputs[154]) ^ (inputs[253]);
    assign layer0_outputs[4111] = ~(inputs[7]);
    assign layer0_outputs[4112] = (inputs[105]) | (inputs[128]);
    assign layer0_outputs[4113] = ~(inputs[59]);
    assign layer0_outputs[4114] = (inputs[45]) & ~(inputs[132]);
    assign layer0_outputs[4115] = (inputs[64]) | (inputs[149]);
    assign layer0_outputs[4116] = 1'b0;
    assign layer0_outputs[4117] = inputs[164];
    assign layer0_outputs[4118] = ~((inputs[118]) | (inputs[20]));
    assign layer0_outputs[4119] = (inputs[246]) & ~(inputs[125]);
    assign layer0_outputs[4120] = ~(inputs[10]);
    assign layer0_outputs[4121] = ~(inputs[145]) | (inputs[121]);
    assign layer0_outputs[4122] = (inputs[209]) ^ (inputs[217]);
    assign layer0_outputs[4123] = (inputs[204]) & (inputs[45]);
    assign layer0_outputs[4124] = (inputs[192]) | (inputs[179]);
    assign layer0_outputs[4125] = ~((inputs[133]) | (inputs[80]));
    assign layer0_outputs[4126] = ~((inputs[39]) ^ (inputs[8]));
    assign layer0_outputs[4127] = ~(inputs[149]) | (inputs[34]);
    assign layer0_outputs[4128] = 1'b0;
    assign layer0_outputs[4129] = inputs[216];
    assign layer0_outputs[4130] = (inputs[127]) & ~(inputs[48]);
    assign layer0_outputs[4131] = ~(inputs[219]);
    assign layer0_outputs[4132] = (inputs[104]) & ~(inputs[253]);
    assign layer0_outputs[4133] = ~(inputs[158]) | (inputs[204]);
    assign layer0_outputs[4134] = ~(inputs[42]) | (inputs[235]);
    assign layer0_outputs[4135] = ~(inputs[189]) | (inputs[66]);
    assign layer0_outputs[4136] = ~(inputs[104]) | (inputs[98]);
    assign layer0_outputs[4137] = (inputs[60]) ^ (inputs[223]);
    assign layer0_outputs[4138] = ~(inputs[102]);
    assign layer0_outputs[4139] = 1'b0;
    assign layer0_outputs[4140] = (inputs[218]) & (inputs[10]);
    assign layer0_outputs[4141] = inputs[248];
    assign layer0_outputs[4142] = ~(inputs[136]);
    assign layer0_outputs[4143] = ~(inputs[75]) | (inputs[103]);
    assign layer0_outputs[4144] = (inputs[113]) ^ (inputs[197]);
    assign layer0_outputs[4145] = ~((inputs[180]) ^ (inputs[135]));
    assign layer0_outputs[4146] = ~(inputs[40]);
    assign layer0_outputs[4147] = inputs[83];
    assign layer0_outputs[4148] = ~(inputs[22]);
    assign layer0_outputs[4149] = ~((inputs[146]) | (inputs[85]));
    assign layer0_outputs[4150] = (inputs[63]) & ~(inputs[254]);
    assign layer0_outputs[4151] = ~(inputs[7]);
    assign layer0_outputs[4152] = ~(inputs[167]);
    assign layer0_outputs[4153] = ~((inputs[136]) ^ (inputs[155]));
    assign layer0_outputs[4154] = (inputs[128]) | (inputs[33]);
    assign layer0_outputs[4155] = ~(inputs[155]);
    assign layer0_outputs[4156] = ~((inputs[6]) | (inputs[47]));
    assign layer0_outputs[4157] = ~((inputs[142]) | (inputs[88]));
    assign layer0_outputs[4158] = ~((inputs[22]) ^ (inputs[190]));
    assign layer0_outputs[4159] = ~(inputs[188]) | (inputs[207]);
    assign layer0_outputs[4160] = 1'b1;
    assign layer0_outputs[4161] = (inputs[157]) | (inputs[149]);
    assign layer0_outputs[4162] = ~(inputs[168]) | (inputs[34]);
    assign layer0_outputs[4163] = 1'b0;
    assign layer0_outputs[4164] = ~((inputs[63]) ^ (inputs[32]));
    assign layer0_outputs[4165] = (inputs[189]) & ~(inputs[211]);
    assign layer0_outputs[4166] = ~(inputs[166]);
    assign layer0_outputs[4167] = (inputs[122]) & ~(inputs[8]);
    assign layer0_outputs[4168] = ~(inputs[86]);
    assign layer0_outputs[4169] = ~((inputs[176]) | (inputs[138]));
    assign layer0_outputs[4170] = (inputs[35]) | (inputs[225]);
    assign layer0_outputs[4171] = ~(inputs[46]) | (inputs[139]);
    assign layer0_outputs[4172] = ~(inputs[224]) | (inputs[13]);
    assign layer0_outputs[4173] = (inputs[92]) ^ (inputs[19]);
    assign layer0_outputs[4174] = ~((inputs[130]) ^ (inputs[150]));
    assign layer0_outputs[4175] = ~((inputs[146]) | (inputs[76]));
    assign layer0_outputs[4176] = 1'b1;
    assign layer0_outputs[4177] = ~(inputs[163]);
    assign layer0_outputs[4178] = (inputs[215]) | (inputs[207]);
    assign layer0_outputs[4179] = inputs[124];
    assign layer0_outputs[4180] = (inputs[164]) & ~(inputs[112]);
    assign layer0_outputs[4181] = (inputs[56]) & ~(inputs[53]);
    assign layer0_outputs[4182] = inputs[209];
    assign layer0_outputs[4183] = ~(inputs[254]);
    assign layer0_outputs[4184] = ~((inputs[0]) & (inputs[223]));
    assign layer0_outputs[4185] = (inputs[154]) ^ (inputs[137]);
    assign layer0_outputs[4186] = inputs[123];
    assign layer0_outputs[4187] = ~(inputs[160]);
    assign layer0_outputs[4188] = inputs[3];
    assign layer0_outputs[4189] = ~((inputs[149]) | (inputs[117]));
    assign layer0_outputs[4190] = ~(inputs[56]);
    assign layer0_outputs[4191] = (inputs[55]) | (inputs[39]);
    assign layer0_outputs[4192] = (inputs[140]) ^ (inputs[127]);
    assign layer0_outputs[4193] = (inputs[202]) & ~(inputs[181]);
    assign layer0_outputs[4194] = (inputs[238]) | (inputs[20]);
    assign layer0_outputs[4195] = 1'b0;
    assign layer0_outputs[4196] = (inputs[40]) | (inputs[245]);
    assign layer0_outputs[4197] = ~(inputs[232]);
    assign layer0_outputs[4198] = (inputs[81]) & (inputs[73]);
    assign layer0_outputs[4199] = inputs[58];
    assign layer0_outputs[4200] = ~((inputs[72]) ^ (inputs[47]));
    assign layer0_outputs[4201] = (inputs[204]) | (inputs[32]);
    assign layer0_outputs[4202] = (inputs[165]) & ~(inputs[129]);
    assign layer0_outputs[4203] = (inputs[228]) & ~(inputs[88]);
    assign layer0_outputs[4204] = (inputs[203]) | (inputs[163]);
    assign layer0_outputs[4205] = inputs[194];
    assign layer0_outputs[4206] = (inputs[82]) | (inputs[196]);
    assign layer0_outputs[4207] = ~(inputs[2]);
    assign layer0_outputs[4208] = (inputs[224]) | (inputs[234]);
    assign layer0_outputs[4209] = ~(inputs[120]) | (inputs[123]);
    assign layer0_outputs[4210] = ~(inputs[243]);
    assign layer0_outputs[4211] = ~(inputs[52]) | (inputs[134]);
    assign layer0_outputs[4212] = ~(inputs[125]);
    assign layer0_outputs[4213] = 1'b0;
    assign layer0_outputs[4214] = inputs[229];
    assign layer0_outputs[4215] = 1'b0;
    assign layer0_outputs[4216] = ~((inputs[84]) ^ (inputs[205]));
    assign layer0_outputs[4217] = ~(inputs[163]);
    assign layer0_outputs[4218] = inputs[139];
    assign layer0_outputs[4219] = ~((inputs[189]) & (inputs[136]));
    assign layer0_outputs[4220] = (inputs[89]) ^ (inputs[223]);
    assign layer0_outputs[4221] = inputs[146];
    assign layer0_outputs[4222] = (inputs[212]) ^ (inputs[157]);
    assign layer0_outputs[4223] = ~((inputs[150]) | (inputs[45]));
    assign layer0_outputs[4224] = inputs[90];
    assign layer0_outputs[4225] = inputs[110];
    assign layer0_outputs[4226] = ~(inputs[44]);
    assign layer0_outputs[4227] = inputs[85];
    assign layer0_outputs[4228] = ~(inputs[245]) | (inputs[16]);
    assign layer0_outputs[4229] = ~(inputs[237]) | (inputs[157]);
    assign layer0_outputs[4230] = (inputs[189]) | (inputs[238]);
    assign layer0_outputs[4231] = ~((inputs[205]) & (inputs[202]));
    assign layer0_outputs[4232] = ~(inputs[99]);
    assign layer0_outputs[4233] = inputs[8];
    assign layer0_outputs[4234] = (inputs[100]) & ~(inputs[95]);
    assign layer0_outputs[4235] = ~(inputs[32]) | (inputs[219]);
    assign layer0_outputs[4236] = (inputs[114]) & ~(inputs[232]);
    assign layer0_outputs[4237] = inputs[76];
    assign layer0_outputs[4238] = inputs[183];
    assign layer0_outputs[4239] = (inputs[195]) | (inputs[194]);
    assign layer0_outputs[4240] = inputs[219];
    assign layer0_outputs[4241] = ~((inputs[190]) ^ (inputs[237]));
    assign layer0_outputs[4242] = ~(inputs[143]);
    assign layer0_outputs[4243] = ~(inputs[162]);
    assign layer0_outputs[4244] = (inputs[10]) & (inputs[24]);
    assign layer0_outputs[4245] = (inputs[167]) | (inputs[164]);
    assign layer0_outputs[4246] = ~(inputs[131]) | (inputs[220]);
    assign layer0_outputs[4247] = ~((inputs[185]) ^ (inputs[174]));
    assign layer0_outputs[4248] = (inputs[215]) | (inputs[202]);
    assign layer0_outputs[4249] = ~((inputs[217]) ^ (inputs[124]));
    assign layer0_outputs[4250] = inputs[120];
    assign layer0_outputs[4251] = ~((inputs[28]) ^ (inputs[49]));
    assign layer0_outputs[4252] = (inputs[55]) & ~(inputs[237]);
    assign layer0_outputs[4253] = ~(inputs[29]) | (inputs[158]);
    assign layer0_outputs[4254] = (inputs[83]) | (inputs[98]);
    assign layer0_outputs[4255] = (inputs[215]) & ~(inputs[158]);
    assign layer0_outputs[4256] = ~(inputs[183]) | (inputs[183]);
    assign layer0_outputs[4257] = inputs[163];
    assign layer0_outputs[4258] = 1'b1;
    assign layer0_outputs[4259] = (inputs[5]) & (inputs[66]);
    assign layer0_outputs[4260] = inputs[23];
    assign layer0_outputs[4261] = ~(inputs[28]);
    assign layer0_outputs[4262] = (inputs[34]) & ~(inputs[142]);
    assign layer0_outputs[4263] = ~(inputs[168]);
    assign layer0_outputs[4264] = inputs[84];
    assign layer0_outputs[4265] = (inputs[229]) ^ (inputs[161]);
    assign layer0_outputs[4266] = ~(inputs[102]) | (inputs[74]);
    assign layer0_outputs[4267] = inputs[139];
    assign layer0_outputs[4268] = ~(inputs[118]);
    assign layer0_outputs[4269] = ~((inputs[56]) | (inputs[113]));
    assign layer0_outputs[4270] = ~((inputs[221]) | (inputs[166]));
    assign layer0_outputs[4271] = ~((inputs[197]) ^ (inputs[150]));
    assign layer0_outputs[4272] = ~((inputs[63]) | (inputs[25]));
    assign layer0_outputs[4273] = ~(inputs[34]);
    assign layer0_outputs[4274] = inputs[253];
    assign layer0_outputs[4275] = inputs[153];
    assign layer0_outputs[4276] = ~(inputs[110]) | (inputs[118]);
    assign layer0_outputs[4277] = (inputs[230]) | (inputs[158]);
    assign layer0_outputs[4278] = (inputs[80]) | (inputs[180]);
    assign layer0_outputs[4279] = inputs[60];
    assign layer0_outputs[4280] = ~((inputs[209]) | (inputs[206]));
    assign layer0_outputs[4281] = 1'b0;
    assign layer0_outputs[4282] = (inputs[171]) & ~(inputs[174]);
    assign layer0_outputs[4283] = ~((inputs[105]) | (inputs[240]));
    assign layer0_outputs[4284] = (inputs[97]) | (inputs[128]);
    assign layer0_outputs[4285] = ~(inputs[170]);
    assign layer0_outputs[4286] = (inputs[69]) ^ (inputs[81]);
    assign layer0_outputs[4287] = inputs[76];
    assign layer0_outputs[4288] = inputs[149];
    assign layer0_outputs[4289] = ~(inputs[215]) | (inputs[107]);
    assign layer0_outputs[4290] = (inputs[215]) & (inputs[234]);
    assign layer0_outputs[4291] = (inputs[36]) ^ (inputs[118]);
    assign layer0_outputs[4292] = inputs[188];
    assign layer0_outputs[4293] = ~(inputs[12]) | (inputs[240]);
    assign layer0_outputs[4294] = (inputs[106]) & ~(inputs[126]);
    assign layer0_outputs[4295] = ~((inputs[9]) | (inputs[243]));
    assign layer0_outputs[4296] = ~(inputs[233]);
    assign layer0_outputs[4297] = ~((inputs[78]) ^ (inputs[92]));
    assign layer0_outputs[4298] = 1'b1;
    assign layer0_outputs[4299] = 1'b1;
    assign layer0_outputs[4300] = ~(inputs[238]) | (inputs[206]);
    assign layer0_outputs[4301] = ~((inputs[189]) | (inputs[209]));
    assign layer0_outputs[4302] = (inputs[207]) | (inputs[81]);
    assign layer0_outputs[4303] = (inputs[207]) & ~(inputs[125]);
    assign layer0_outputs[4304] = inputs[60];
    assign layer0_outputs[4305] = inputs[254];
    assign layer0_outputs[4306] = inputs[58];
    assign layer0_outputs[4307] = 1'b1;
    assign layer0_outputs[4308] = (inputs[64]) ^ (inputs[40]);
    assign layer0_outputs[4309] = (inputs[179]) | (inputs[111]);
    assign layer0_outputs[4310] = ~(inputs[205]);
    assign layer0_outputs[4311] = (inputs[186]) | (inputs[165]);
    assign layer0_outputs[4312] = ~(inputs[106]);
    assign layer0_outputs[4313] = (inputs[175]) | (inputs[228]);
    assign layer0_outputs[4314] = 1'b0;
    assign layer0_outputs[4315] = ~(inputs[13]) | (inputs[184]);
    assign layer0_outputs[4316] = ~(inputs[35]);
    assign layer0_outputs[4317] = inputs[21];
    assign layer0_outputs[4318] = ~((inputs[185]) & (inputs[166]));
    assign layer0_outputs[4319] = ~(inputs[194]) | (inputs[168]);
    assign layer0_outputs[4320] = ~(inputs[51]);
    assign layer0_outputs[4321] = ~(inputs[212]);
    assign layer0_outputs[4322] = ~(inputs[133]) | (inputs[49]);
    assign layer0_outputs[4323] = (inputs[132]) & (inputs[155]);
    assign layer0_outputs[4324] = ~(inputs[168]);
    assign layer0_outputs[4325] = inputs[72];
    assign layer0_outputs[4326] = ~(inputs[254]) | (inputs[178]);
    assign layer0_outputs[4327] = ~((inputs[105]) ^ (inputs[165]));
    assign layer0_outputs[4328] = ~(inputs[111]);
    assign layer0_outputs[4329] = ~((inputs[243]) | (inputs[33]));
    assign layer0_outputs[4330] = (inputs[106]) ^ (inputs[16]);
    assign layer0_outputs[4331] = ~((inputs[48]) | (inputs[235]));
    assign layer0_outputs[4332] = (inputs[201]) & ~(inputs[142]);
    assign layer0_outputs[4333] = (inputs[86]) | (inputs[3]);
    assign layer0_outputs[4334] = ~((inputs[80]) ^ (inputs[51]));
    assign layer0_outputs[4335] = (inputs[38]) ^ (inputs[71]);
    assign layer0_outputs[4336] = ~((inputs[178]) | (inputs[252]));
    assign layer0_outputs[4337] = ~((inputs[14]) | (inputs[41]));
    assign layer0_outputs[4338] = ~(inputs[178]);
    assign layer0_outputs[4339] = ~(inputs[33]);
    assign layer0_outputs[4340] = ~(inputs[45]) | (inputs[252]);
    assign layer0_outputs[4341] = (inputs[173]) ^ (inputs[19]);
    assign layer0_outputs[4342] = inputs[110];
    assign layer0_outputs[4343] = ~(inputs[245]);
    assign layer0_outputs[4344] = ~(inputs[192]);
    assign layer0_outputs[4345] = ~((inputs[162]) ^ (inputs[158]));
    assign layer0_outputs[4346] = ~((inputs[211]) | (inputs[198]));
    assign layer0_outputs[4347] = inputs[101];
    assign layer0_outputs[4348] = inputs[163];
    assign layer0_outputs[4349] = (inputs[49]) | (inputs[26]);
    assign layer0_outputs[4350] = inputs[215];
    assign layer0_outputs[4351] = (inputs[129]) ^ (inputs[109]);
    assign layer0_outputs[4352] = ~(inputs[25]);
    assign layer0_outputs[4353] = (inputs[84]) ^ (inputs[82]);
    assign layer0_outputs[4354] = ~((inputs[237]) & (inputs[58]));
    assign layer0_outputs[4355] = ~(inputs[66]) | (inputs[224]);
    assign layer0_outputs[4356] = ~((inputs[94]) ^ (inputs[89]));
    assign layer0_outputs[4357] = 1'b1;
    assign layer0_outputs[4358] = (inputs[121]) & ~(inputs[157]);
    assign layer0_outputs[4359] = ~(inputs[35]);
    assign layer0_outputs[4360] = inputs[88];
    assign layer0_outputs[4361] = (inputs[83]) & ~(inputs[2]);
    assign layer0_outputs[4362] = inputs[78];
    assign layer0_outputs[4363] = inputs[162];
    assign layer0_outputs[4364] = ~(inputs[124]) | (inputs[144]);
    assign layer0_outputs[4365] = inputs[189];
    assign layer0_outputs[4366] = 1'b0;
    assign layer0_outputs[4367] = 1'b1;
    assign layer0_outputs[4368] = ~(inputs[10]);
    assign layer0_outputs[4369] = ~(inputs[12]) | (inputs[80]);
    assign layer0_outputs[4370] = ~(inputs[121]);
    assign layer0_outputs[4371] = (inputs[149]) & ~(inputs[229]);
    assign layer0_outputs[4372] = (inputs[78]) | (inputs[155]);
    assign layer0_outputs[4373] = (inputs[66]) & ~(inputs[215]);
    assign layer0_outputs[4374] = inputs[180];
    assign layer0_outputs[4375] = ~((inputs[39]) | (inputs[22]));
    assign layer0_outputs[4376] = ~(inputs[59]);
    assign layer0_outputs[4377] = ~((inputs[144]) | (inputs[133]));
    assign layer0_outputs[4378] = ~(inputs[115]);
    assign layer0_outputs[4379] = (inputs[194]) & ~(inputs[188]);
    assign layer0_outputs[4380] = (inputs[168]) | (inputs[137]);
    assign layer0_outputs[4381] = ~(inputs[137]) | (inputs[142]);
    assign layer0_outputs[4382] = inputs[165];
    assign layer0_outputs[4383] = (inputs[206]) ^ (inputs[108]);
    assign layer0_outputs[4384] = (inputs[120]) | (inputs[84]);
    assign layer0_outputs[4385] = ~((inputs[129]) & (inputs[96]));
    assign layer0_outputs[4386] = (inputs[48]) | (inputs[52]);
    assign layer0_outputs[4387] = (inputs[255]) | (inputs[193]);
    assign layer0_outputs[4388] = ~(inputs[77]) | (inputs[178]);
    assign layer0_outputs[4389] = (inputs[175]) & ~(inputs[142]);
    assign layer0_outputs[4390] = ~((inputs[83]) | (inputs[177]));
    assign layer0_outputs[4391] = ~(inputs[172]) | (inputs[152]);
    assign layer0_outputs[4392] = (inputs[98]) & (inputs[42]);
    assign layer0_outputs[4393] = inputs[153];
    assign layer0_outputs[4394] = (inputs[117]) | (inputs[248]);
    assign layer0_outputs[4395] = (inputs[215]) & ~(inputs[71]);
    assign layer0_outputs[4396] = (inputs[54]) & ~(inputs[149]);
    assign layer0_outputs[4397] = ~((inputs[144]) ^ (inputs[132]));
    assign layer0_outputs[4398] = ~((inputs[59]) | (inputs[77]));
    assign layer0_outputs[4399] = ~((inputs[247]) ^ (inputs[143]));
    assign layer0_outputs[4400] = 1'b0;
    assign layer0_outputs[4401] = ~(inputs[1]);
    assign layer0_outputs[4402] = ~((inputs[20]) ^ (inputs[68]));
    assign layer0_outputs[4403] = (inputs[128]) & ~(inputs[70]);
    assign layer0_outputs[4404] = (inputs[138]) & ~(inputs[27]);
    assign layer0_outputs[4405] = inputs[211];
    assign layer0_outputs[4406] = 1'b1;
    assign layer0_outputs[4407] = ~(inputs[235]);
    assign layer0_outputs[4408] = (inputs[214]) & ~(inputs[73]);
    assign layer0_outputs[4409] = ~((inputs[26]) | (inputs[94]));
    assign layer0_outputs[4410] = (inputs[171]) & ~(inputs[14]);
    assign layer0_outputs[4411] = ~(inputs[16]);
    assign layer0_outputs[4412] = inputs[19];
    assign layer0_outputs[4413] = inputs[246];
    assign layer0_outputs[4414] = (inputs[85]) | (inputs[55]);
    assign layer0_outputs[4415] = (inputs[222]) & ~(inputs[108]);
    assign layer0_outputs[4416] = (inputs[234]) & ~(inputs[45]);
    assign layer0_outputs[4417] = inputs[109];
    assign layer0_outputs[4418] = ~((inputs[166]) ^ (inputs[247]));
    assign layer0_outputs[4419] = (inputs[33]) | (inputs[199]);
    assign layer0_outputs[4420] = inputs[215];
    assign layer0_outputs[4421] = (inputs[106]) | (inputs[60]);
    assign layer0_outputs[4422] = ~(inputs[242]) | (inputs[200]);
    assign layer0_outputs[4423] = (inputs[128]) & ~(inputs[112]);
    assign layer0_outputs[4424] = inputs[98];
    assign layer0_outputs[4425] = ~((inputs[134]) ^ (inputs[161]));
    assign layer0_outputs[4426] = inputs[6];
    assign layer0_outputs[4427] = ~((inputs[1]) | (inputs[65]));
    assign layer0_outputs[4428] = ~(inputs[40]);
    assign layer0_outputs[4429] = inputs[233];
    assign layer0_outputs[4430] = (inputs[75]) & (inputs[103]);
    assign layer0_outputs[4431] = ~((inputs[89]) ^ (inputs[42]));
    assign layer0_outputs[4432] = inputs[127];
    assign layer0_outputs[4433] = ~((inputs[217]) ^ (inputs[184]));
    assign layer0_outputs[4434] = ~(inputs[151]);
    assign layer0_outputs[4435] = (inputs[143]) | (inputs[89]);
    assign layer0_outputs[4436] = (inputs[5]) & ~(inputs[144]);
    assign layer0_outputs[4437] = ~(inputs[246]) | (inputs[178]);
    assign layer0_outputs[4438] = inputs[68];
    assign layer0_outputs[4439] = (inputs[221]) & (inputs[144]);
    assign layer0_outputs[4440] = inputs[92];
    assign layer0_outputs[4441] = ~((inputs[197]) ^ (inputs[191]));
    assign layer0_outputs[4442] = inputs[114];
    assign layer0_outputs[4443] = (inputs[148]) & ~(inputs[152]);
    assign layer0_outputs[4444] = ~((inputs[28]) ^ (inputs[176]));
    assign layer0_outputs[4445] = ~(inputs[64]);
    assign layer0_outputs[4446] = inputs[145];
    assign layer0_outputs[4447] = inputs[123];
    assign layer0_outputs[4448] = ~(inputs[131]);
    assign layer0_outputs[4449] = ~((inputs[136]) | (inputs[168]));
    assign layer0_outputs[4450] = (inputs[189]) & ~(inputs[33]);
    assign layer0_outputs[4451] = (inputs[213]) | (inputs[229]);
    assign layer0_outputs[4452] = ~((inputs[202]) | (inputs[174]));
    assign layer0_outputs[4453] = inputs[89];
    assign layer0_outputs[4454] = ~(inputs[176]) | (inputs[4]);
    assign layer0_outputs[4455] = (inputs[251]) | (inputs[198]);
    assign layer0_outputs[4456] = ~(inputs[135]) | (inputs[128]);
    assign layer0_outputs[4457] = ~(inputs[122]) | (inputs[253]);
    assign layer0_outputs[4458] = ~(inputs[116]);
    assign layer0_outputs[4459] = (inputs[24]) | (inputs[111]);
    assign layer0_outputs[4460] = (inputs[58]) ^ (inputs[40]);
    assign layer0_outputs[4461] = (inputs[158]) ^ (inputs[100]);
    assign layer0_outputs[4462] = ~((inputs[10]) | (inputs[97]));
    assign layer0_outputs[4463] = (inputs[7]) & ~(inputs[145]);
    assign layer0_outputs[4464] = (inputs[104]) ^ (inputs[123]);
    assign layer0_outputs[4465] = (inputs[58]) & ~(inputs[216]);
    assign layer0_outputs[4466] = inputs[122];
    assign layer0_outputs[4467] = ~(inputs[132]) | (inputs[48]);
    assign layer0_outputs[4468] = (inputs[8]) & (inputs[25]);
    assign layer0_outputs[4469] = ~(inputs[39]) | (inputs[241]);
    assign layer0_outputs[4470] = (inputs[129]) & ~(inputs[239]);
    assign layer0_outputs[4471] = (inputs[178]) ^ (inputs[112]);
    assign layer0_outputs[4472] = ~((inputs[130]) | (inputs[186]));
    assign layer0_outputs[4473] = ~(inputs[143]) | (inputs[171]);
    assign layer0_outputs[4474] = ~(inputs[232]) | (inputs[242]);
    assign layer0_outputs[4475] = ~((inputs[71]) ^ (inputs[203]));
    assign layer0_outputs[4476] = (inputs[132]) & ~(inputs[13]);
    assign layer0_outputs[4477] = ~(inputs[99]);
    assign layer0_outputs[4478] = ~((inputs[130]) | (inputs[132]));
    assign layer0_outputs[4479] = (inputs[232]) & ~(inputs[35]);
    assign layer0_outputs[4480] = ~(inputs[79]);
    assign layer0_outputs[4481] = (inputs[42]) & ~(inputs[170]);
    assign layer0_outputs[4482] = ~(inputs[167]) | (inputs[46]);
    assign layer0_outputs[4483] = ~(inputs[232]);
    assign layer0_outputs[4484] = ~(inputs[174]);
    assign layer0_outputs[4485] = ~(inputs[7]) | (inputs[0]);
    assign layer0_outputs[4486] = (inputs[118]) ^ (inputs[131]);
    assign layer0_outputs[4487] = inputs[10];
    assign layer0_outputs[4488] = ~(inputs[6]) | (inputs[221]);
    assign layer0_outputs[4489] = ~(inputs[20]) | (inputs[153]);
    assign layer0_outputs[4490] = (inputs[81]) ^ (inputs[79]);
    assign layer0_outputs[4491] = inputs[94];
    assign layer0_outputs[4492] = ~((inputs[162]) | (inputs[7]));
    assign layer0_outputs[4493] = ~((inputs[109]) | (inputs[23]));
    assign layer0_outputs[4494] = ~((inputs[64]) ^ (inputs[61]));
    assign layer0_outputs[4495] = (inputs[86]) & ~(inputs[249]);
    assign layer0_outputs[4496] = (inputs[216]) | (inputs[164]);
    assign layer0_outputs[4497] = (inputs[13]) | (inputs[96]);
    assign layer0_outputs[4498] = ~(inputs[165]) | (inputs[84]);
    assign layer0_outputs[4499] = ~(inputs[89]);
    assign layer0_outputs[4500] = ~(inputs[8]) | (inputs[1]);
    assign layer0_outputs[4501] = ~(inputs[63]);
    assign layer0_outputs[4502] = ~(inputs[88]) | (inputs[227]);
    assign layer0_outputs[4503] = ~((inputs[24]) | (inputs[1]));
    assign layer0_outputs[4504] = (inputs[181]) ^ (inputs[179]);
    assign layer0_outputs[4505] = ~((inputs[225]) & (inputs[179]));
    assign layer0_outputs[4506] = inputs[114];
    assign layer0_outputs[4507] = (inputs[24]) & ~(inputs[178]);
    assign layer0_outputs[4508] = ~(inputs[174]);
    assign layer0_outputs[4509] = 1'b0;
    assign layer0_outputs[4510] = ~(inputs[13]) | (inputs[151]);
    assign layer0_outputs[4511] = ~(inputs[132]) | (inputs[45]);
    assign layer0_outputs[4512] = ~(inputs[230]);
    assign layer0_outputs[4513] = ~(inputs[138]) | (inputs[140]);
    assign layer0_outputs[4514] = ~((inputs[68]) | (inputs[188]));
    assign layer0_outputs[4515] = (inputs[176]) | (inputs[14]);
    assign layer0_outputs[4516] = ~(inputs[148]);
    assign layer0_outputs[4517] = inputs[17];
    assign layer0_outputs[4518] = ~((inputs[255]) | (inputs[177]));
    assign layer0_outputs[4519] = ~(inputs[152]) | (inputs[203]);
    assign layer0_outputs[4520] = (inputs[202]) & ~(inputs[108]);
    assign layer0_outputs[4521] = ~((inputs[237]) | (inputs[164]));
    assign layer0_outputs[4522] = 1'b0;
    assign layer0_outputs[4523] = ~(inputs[124]);
    assign layer0_outputs[4524] = ~(inputs[234]);
    assign layer0_outputs[4525] = ~((inputs[126]) ^ (inputs[243]));
    assign layer0_outputs[4526] = ~((inputs[10]) | (inputs[91]));
    assign layer0_outputs[4527] = (inputs[24]) & ~(inputs[115]);
    assign layer0_outputs[4528] = (inputs[18]) ^ (inputs[91]);
    assign layer0_outputs[4529] = inputs[153];
    assign layer0_outputs[4530] = ~((inputs[168]) & (inputs[19]));
    assign layer0_outputs[4531] = inputs[20];
    assign layer0_outputs[4532] = ~((inputs[164]) | (inputs[201]));
    assign layer0_outputs[4533] = (inputs[184]) ^ (inputs[83]);
    assign layer0_outputs[4534] = (inputs[144]) | (inputs[142]);
    assign layer0_outputs[4535] = ~((inputs[194]) | (inputs[196]));
    assign layer0_outputs[4536] = (inputs[25]) ^ (inputs[71]);
    assign layer0_outputs[4537] = ~(inputs[60]);
    assign layer0_outputs[4538] = ~(inputs[12]) | (inputs[95]);
    assign layer0_outputs[4539] = ~((inputs[170]) | (inputs[206]));
    assign layer0_outputs[4540] = (inputs[204]) | (inputs[249]);
    assign layer0_outputs[4541] = ~(inputs[155]) | (inputs[109]);
    assign layer0_outputs[4542] = ~(inputs[122]);
    assign layer0_outputs[4543] = ~((inputs[203]) & (inputs[4]));
    assign layer0_outputs[4544] = (inputs[117]) | (inputs[148]);
    assign layer0_outputs[4545] = ~(inputs[50]);
    assign layer0_outputs[4546] = ~(inputs[209]);
    assign layer0_outputs[4547] = (inputs[50]) | (inputs[29]);
    assign layer0_outputs[4548] = 1'b1;
    assign layer0_outputs[4549] = ~(inputs[104]);
    assign layer0_outputs[4550] = ~((inputs[41]) & (inputs[228]));
    assign layer0_outputs[4551] = inputs[36];
    assign layer0_outputs[4552] = (inputs[104]) & ~(inputs[54]);
    assign layer0_outputs[4553] = 1'b0;
    assign layer0_outputs[4554] = inputs[111];
    assign layer0_outputs[4555] = ~((inputs[252]) ^ (inputs[142]));
    assign layer0_outputs[4556] = (inputs[252]) | (inputs[176]);
    assign layer0_outputs[4557] = (inputs[138]) | (inputs[77]);
    assign layer0_outputs[4558] = ~(inputs[122]);
    assign layer0_outputs[4559] = ~(inputs[86]);
    assign layer0_outputs[4560] = ~(inputs[40]);
    assign layer0_outputs[4561] = (inputs[83]) & (inputs[16]);
    assign layer0_outputs[4562] = (inputs[24]) & (inputs[26]);
    assign layer0_outputs[4563] = inputs[196];
    assign layer0_outputs[4564] = ~(inputs[148]);
    assign layer0_outputs[4565] = inputs[51];
    assign layer0_outputs[4566] = ~(inputs[229]);
    assign layer0_outputs[4567] = (inputs[214]) & ~(inputs[156]);
    assign layer0_outputs[4568] = ~(inputs[53]) | (inputs[192]);
    assign layer0_outputs[4569] = inputs[169];
    assign layer0_outputs[4570] = ~(inputs[187]);
    assign layer0_outputs[4571] = (inputs[156]) & ~(inputs[12]);
    assign layer0_outputs[4572] = (inputs[106]) | (inputs[205]);
    assign layer0_outputs[4573] = (inputs[246]) ^ (inputs[214]);
    assign layer0_outputs[4574] = ~(inputs[214]);
    assign layer0_outputs[4575] = ~(inputs[248]);
    assign layer0_outputs[4576] = (inputs[190]) & ~(inputs[225]);
    assign layer0_outputs[4577] = inputs[100];
    assign layer0_outputs[4578] = inputs[237];
    assign layer0_outputs[4579] = ~(inputs[122]);
    assign layer0_outputs[4580] = inputs[39];
    assign layer0_outputs[4581] = (inputs[171]) & ~(inputs[37]);
    assign layer0_outputs[4582] = (inputs[163]) | (inputs[178]);
    assign layer0_outputs[4583] = (inputs[143]) | (inputs[12]);
    assign layer0_outputs[4584] = ~(inputs[179]);
    assign layer0_outputs[4585] = (inputs[121]) | (inputs[91]);
    assign layer0_outputs[4586] = (inputs[125]) ^ (inputs[204]);
    assign layer0_outputs[4587] = (inputs[5]) | (inputs[41]);
    assign layer0_outputs[4588] = ~(inputs[175]);
    assign layer0_outputs[4589] = (inputs[127]) ^ (inputs[0]);
    assign layer0_outputs[4590] = (inputs[64]) | (inputs[75]);
    assign layer0_outputs[4591] = ~((inputs[236]) ^ (inputs[172]));
    assign layer0_outputs[4592] = ~(inputs[243]) | (inputs[56]);
    assign layer0_outputs[4593] = (inputs[220]) | (inputs[105]);
    assign layer0_outputs[4594] = inputs[21];
    assign layer0_outputs[4595] = inputs[75];
    assign layer0_outputs[4596] = ~((inputs[27]) | (inputs[208]));
    assign layer0_outputs[4597] = ~(inputs[59]) | (inputs[205]);
    assign layer0_outputs[4598] = (inputs[119]) | (inputs[71]);
    assign layer0_outputs[4599] = ~((inputs[162]) | (inputs[144]));
    assign layer0_outputs[4600] = ~(inputs[44]);
    assign layer0_outputs[4601] = ~(inputs[127]);
    assign layer0_outputs[4602] = ~((inputs[40]) | (inputs[175]));
    assign layer0_outputs[4603] = inputs[233];
    assign layer0_outputs[4604] = inputs[98];
    assign layer0_outputs[4605] = ~(inputs[24]) | (inputs[166]);
    assign layer0_outputs[4606] = ~(inputs[246]);
    assign layer0_outputs[4607] = inputs[188];
    assign layer0_outputs[4608] = 1'b1;
    assign layer0_outputs[4609] = ~(inputs[139]) | (inputs[243]);
    assign layer0_outputs[4610] = ~((inputs[211]) ^ (inputs[16]));
    assign layer0_outputs[4611] = ~((inputs[199]) | (inputs[215]));
    assign layer0_outputs[4612] = ~((inputs[109]) | (inputs[82]));
    assign layer0_outputs[4613] = ~((inputs[74]) | (inputs[33]));
    assign layer0_outputs[4614] = 1'b1;
    assign layer0_outputs[4615] = (inputs[181]) ^ (inputs[138]);
    assign layer0_outputs[4616] = (inputs[227]) ^ (inputs[134]);
    assign layer0_outputs[4617] = ~(inputs[112]) | (inputs[30]);
    assign layer0_outputs[4618] = (inputs[145]) | (inputs[248]);
    assign layer0_outputs[4619] = (inputs[177]) | (inputs[247]);
    assign layer0_outputs[4620] = (inputs[30]) | (inputs[56]);
    assign layer0_outputs[4621] = ~((inputs[161]) ^ (inputs[218]));
    assign layer0_outputs[4622] = 1'b1;
    assign layer0_outputs[4623] = (inputs[11]) | (inputs[13]);
    assign layer0_outputs[4624] = inputs[179];
    assign layer0_outputs[4625] = inputs[184];
    assign layer0_outputs[4626] = ~((inputs[3]) & (inputs[157]));
    assign layer0_outputs[4627] = ~(inputs[154]);
    assign layer0_outputs[4628] = ~(inputs[160]);
    assign layer0_outputs[4629] = ~((inputs[76]) | (inputs[97]));
    assign layer0_outputs[4630] = ~(inputs[247]) | (inputs[12]);
    assign layer0_outputs[4631] = inputs[46];
    assign layer0_outputs[4632] = (inputs[186]) & (inputs[179]);
    assign layer0_outputs[4633] = (inputs[158]) | (inputs[4]);
    assign layer0_outputs[4634] = (inputs[154]) & ~(inputs[248]);
    assign layer0_outputs[4635] = ~(inputs[102]);
    assign layer0_outputs[4636] = ~((inputs[16]) | (inputs[10]));
    assign layer0_outputs[4637] = ~(inputs[102]) | (inputs[17]);
    assign layer0_outputs[4638] = 1'b0;
    assign layer0_outputs[4639] = ~(inputs[220]) | (inputs[196]);
    assign layer0_outputs[4640] = ~(inputs[29]);
    assign layer0_outputs[4641] = ~(inputs[128]) | (inputs[3]);
    assign layer0_outputs[4642] = ~(inputs[115]) | (inputs[31]);
    assign layer0_outputs[4643] = (inputs[15]) & ~(inputs[20]);
    assign layer0_outputs[4644] = ~(inputs[54]) | (inputs[180]);
    assign layer0_outputs[4645] = inputs[91];
    assign layer0_outputs[4646] = inputs[121];
    assign layer0_outputs[4647] = ~((inputs[128]) ^ (inputs[82]));
    assign layer0_outputs[4648] = 1'b1;
    assign layer0_outputs[4649] = ~((inputs[207]) ^ (inputs[250]));
    assign layer0_outputs[4650] = (inputs[14]) ^ (inputs[47]);
    assign layer0_outputs[4651] = ~(inputs[82]);
    assign layer0_outputs[4652] = ~((inputs[246]) & (inputs[251]));
    assign layer0_outputs[4653] = ~(inputs[229]);
    assign layer0_outputs[4654] = inputs[5];
    assign layer0_outputs[4655] = (inputs[96]) & (inputs[166]);
    assign layer0_outputs[4656] = (inputs[71]) & ~(inputs[177]);
    assign layer0_outputs[4657] = ~(inputs[79]);
    assign layer0_outputs[4658] = inputs[162];
    assign layer0_outputs[4659] = ~(inputs[80]);
    assign layer0_outputs[4660] = ~(inputs[150]) | (inputs[47]);
    assign layer0_outputs[4661] = ~(inputs[181]);
    assign layer0_outputs[4662] = inputs[218];
    assign layer0_outputs[4663] = (inputs[103]) & ~(inputs[103]);
    assign layer0_outputs[4664] = ~((inputs[166]) & (inputs[43]));
    assign layer0_outputs[4665] = (inputs[8]) | (inputs[91]);
    assign layer0_outputs[4666] = 1'b1;
    assign layer0_outputs[4667] = ~((inputs[255]) ^ (inputs[117]));
    assign layer0_outputs[4668] = (inputs[100]) ^ (inputs[71]);
    assign layer0_outputs[4669] = ~(inputs[103]);
    assign layer0_outputs[4670] = (inputs[48]) & ~(inputs[242]);
    assign layer0_outputs[4671] = ~((inputs[200]) & (inputs[118]));
    assign layer0_outputs[4672] = ~((inputs[192]) | (inputs[200]));
    assign layer0_outputs[4673] = ~(inputs[142]) | (inputs[79]);
    assign layer0_outputs[4674] = ~(inputs[55]) | (inputs[130]);
    assign layer0_outputs[4675] = (inputs[231]) & (inputs[23]);
    assign layer0_outputs[4676] = (inputs[147]) | (inputs[212]);
    assign layer0_outputs[4677] = inputs[55];
    assign layer0_outputs[4678] = 1'b1;
    assign layer0_outputs[4679] = (inputs[57]) & ~(inputs[187]);
    assign layer0_outputs[4680] = ~(inputs[136]) | (inputs[99]);
    assign layer0_outputs[4681] = (inputs[252]) | (inputs[237]);
    assign layer0_outputs[4682] = (inputs[247]) ^ (inputs[67]);
    assign layer0_outputs[4683] = ~(inputs[92]);
    assign layer0_outputs[4684] = ~(inputs[121]) | (inputs[175]);
    assign layer0_outputs[4685] = ~((inputs[152]) ^ (inputs[49]));
    assign layer0_outputs[4686] = ~((inputs[126]) ^ (inputs[108]));
    assign layer0_outputs[4687] = inputs[93];
    assign layer0_outputs[4688] = ~((inputs[225]) & (inputs[16]));
    assign layer0_outputs[4689] = ~(inputs[163]) | (inputs[241]);
    assign layer0_outputs[4690] = 1'b0;
    assign layer0_outputs[4691] = (inputs[250]) | (inputs[139]);
    assign layer0_outputs[4692] = (inputs[121]) ^ (inputs[146]);
    assign layer0_outputs[4693] = ~(inputs[117]) | (inputs[146]);
    assign layer0_outputs[4694] = ~(inputs[60]);
    assign layer0_outputs[4695] = ~((inputs[226]) | (inputs[239]));
    assign layer0_outputs[4696] = (inputs[230]) | (inputs[32]);
    assign layer0_outputs[4697] = ~((inputs[25]) & (inputs[22]));
    assign layer0_outputs[4698] = ~(inputs[106]);
    assign layer0_outputs[4699] = inputs[199];
    assign layer0_outputs[4700] = (inputs[90]) | (inputs[74]);
    assign layer0_outputs[4701] = ~(inputs[246]);
    assign layer0_outputs[4702] = ~((inputs[215]) | (inputs[170]));
    assign layer0_outputs[4703] = ~(inputs[23]) | (inputs[160]);
    assign layer0_outputs[4704] = ~((inputs[192]) | (inputs[176]));
    assign layer0_outputs[4705] = ~(inputs[62]);
    assign layer0_outputs[4706] = (inputs[128]) & (inputs[40]);
    assign layer0_outputs[4707] = ~(inputs[167]);
    assign layer0_outputs[4708] = ~(inputs[131]) | (inputs[66]);
    assign layer0_outputs[4709] = ~(inputs[136]);
    assign layer0_outputs[4710] = inputs[216];
    assign layer0_outputs[4711] = inputs[231];
    assign layer0_outputs[4712] = (inputs[44]) & ~(inputs[91]);
    assign layer0_outputs[4713] = (inputs[72]) & ~(inputs[117]);
    assign layer0_outputs[4714] = (inputs[51]) | (inputs[170]);
    assign layer0_outputs[4715] = inputs[37];
    assign layer0_outputs[4716] = (inputs[233]) ^ (inputs[61]);
    assign layer0_outputs[4717] = (inputs[150]) & (inputs[219]);
    assign layer0_outputs[4718] = ~(inputs[54]);
    assign layer0_outputs[4719] = (inputs[186]) | (inputs[98]);
    assign layer0_outputs[4720] = ~((inputs[64]) ^ (inputs[69]));
    assign layer0_outputs[4721] = ~((inputs[242]) & (inputs[229]));
    assign layer0_outputs[4722] = (inputs[194]) & ~(inputs[94]);
    assign layer0_outputs[4723] = ~(inputs[109]) | (inputs[30]);
    assign layer0_outputs[4724] = ~(inputs[57]) | (inputs[102]);
    assign layer0_outputs[4725] = ~((inputs[97]) & (inputs[210]));
    assign layer0_outputs[4726] = 1'b1;
    assign layer0_outputs[4727] = ~((inputs[243]) ^ (inputs[243]));
    assign layer0_outputs[4728] = (inputs[40]) | (inputs[226]);
    assign layer0_outputs[4729] = inputs[204];
    assign layer0_outputs[4730] = ~(inputs[73]);
    assign layer0_outputs[4731] = ~(inputs[21]);
    assign layer0_outputs[4732] = (inputs[114]) ^ (inputs[47]);
    assign layer0_outputs[4733] = 1'b1;
    assign layer0_outputs[4734] = (inputs[40]) & ~(inputs[68]);
    assign layer0_outputs[4735] = inputs[59];
    assign layer0_outputs[4736] = ~(inputs[208]) | (inputs[13]);
    assign layer0_outputs[4737] = ~(inputs[87]);
    assign layer0_outputs[4738] = inputs[202];
    assign layer0_outputs[4739] = (inputs[252]) & ~(inputs[162]);
    assign layer0_outputs[4740] = (inputs[64]) & (inputs[3]);
    assign layer0_outputs[4741] = ~(inputs[220]);
    assign layer0_outputs[4742] = ~(inputs[148]);
    assign layer0_outputs[4743] = (inputs[221]) & ~(inputs[240]);
    assign layer0_outputs[4744] = ~((inputs[4]) ^ (inputs[125]));
    assign layer0_outputs[4745] = ~(inputs[247]);
    assign layer0_outputs[4746] = (inputs[203]) | (inputs[219]);
    assign layer0_outputs[4747] = ~((inputs[82]) | (inputs[111]));
    assign layer0_outputs[4748] = (inputs[158]) | (inputs[160]);
    assign layer0_outputs[4749] = ~(inputs[169]) | (inputs[154]);
    assign layer0_outputs[4750] = (inputs[84]) | (inputs[132]);
    assign layer0_outputs[4751] = ~(inputs[110]) | (inputs[239]);
    assign layer0_outputs[4752] = ~(inputs[37]) | (inputs[206]);
    assign layer0_outputs[4753] = inputs[7];
    assign layer0_outputs[4754] = ~((inputs[138]) | (inputs[87]));
    assign layer0_outputs[4755] = ~(inputs[131]);
    assign layer0_outputs[4756] = 1'b1;
    assign layer0_outputs[4757] = inputs[114];
    assign layer0_outputs[4758] = ~(inputs[109]) | (inputs[39]);
    assign layer0_outputs[4759] = inputs[8];
    assign layer0_outputs[4760] = ~(inputs[199]);
    assign layer0_outputs[4761] = (inputs[167]) ^ (inputs[11]);
    assign layer0_outputs[4762] = 1'b0;
    assign layer0_outputs[4763] = ~(inputs[250]) | (inputs[126]);
    assign layer0_outputs[4764] = ~(inputs[227]) | (inputs[77]);
    assign layer0_outputs[4765] = (inputs[2]) | (inputs[223]);
    assign layer0_outputs[4766] = inputs[3];
    assign layer0_outputs[4767] = (inputs[225]) & ~(inputs[239]);
    assign layer0_outputs[4768] = (inputs[48]) & ~(inputs[49]);
    assign layer0_outputs[4769] = (inputs[140]) | (inputs[162]);
    assign layer0_outputs[4770] = ~(inputs[73]);
    assign layer0_outputs[4771] = (inputs[116]) & ~(inputs[193]);
    assign layer0_outputs[4772] = ~(inputs[25]);
    assign layer0_outputs[4773] = ~(inputs[240]);
    assign layer0_outputs[4774] = (inputs[33]) & ~(inputs[161]);
    assign layer0_outputs[4775] = ~(inputs[173]);
    assign layer0_outputs[4776] = ~(inputs[98]);
    assign layer0_outputs[4777] = (inputs[26]) & ~(inputs[243]);
    assign layer0_outputs[4778] = ~((inputs[35]) | (inputs[236]));
    assign layer0_outputs[4779] = (inputs[27]) & (inputs[26]);
    assign layer0_outputs[4780] = 1'b0;
    assign layer0_outputs[4781] = ~((inputs[47]) | (inputs[104]));
    assign layer0_outputs[4782] = (inputs[190]) | (inputs[88]);
    assign layer0_outputs[4783] = 1'b1;
    assign layer0_outputs[4784] = (inputs[3]) ^ (inputs[63]);
    assign layer0_outputs[4785] = ~(inputs[185]) | (inputs[14]);
    assign layer0_outputs[4786] = 1'b0;
    assign layer0_outputs[4787] = 1'b1;
    assign layer0_outputs[4788] = (inputs[197]) | (inputs[156]);
    assign layer0_outputs[4789] = (inputs[245]) ^ (inputs[201]);
    assign layer0_outputs[4790] = inputs[96];
    assign layer0_outputs[4791] = ~(inputs[101]);
    assign layer0_outputs[4792] = ~((inputs[21]) & (inputs[25]));
    assign layer0_outputs[4793] = ~(inputs[69]);
    assign layer0_outputs[4794] = (inputs[191]) ^ (inputs[149]);
    assign layer0_outputs[4795] = inputs[103];
    assign layer0_outputs[4796] = (inputs[236]) | (inputs[109]);
    assign layer0_outputs[4797] = (inputs[146]) ^ (inputs[25]);
    assign layer0_outputs[4798] = (inputs[8]) & ~(inputs[164]);
    assign layer0_outputs[4799] = (inputs[159]) ^ (inputs[0]);
    assign layer0_outputs[4800] = (inputs[53]) & ~(inputs[118]);
    assign layer0_outputs[4801] = ~((inputs[104]) | (inputs[203]));
    assign layer0_outputs[4802] = ~(inputs[117]) | (inputs[237]);
    assign layer0_outputs[4803] = inputs[38];
    assign layer0_outputs[4804] = (inputs[217]) | (inputs[129]);
    assign layer0_outputs[4805] = ~(inputs[8]);
    assign layer0_outputs[4806] = (inputs[48]) & ~(inputs[255]);
    assign layer0_outputs[4807] = ~(inputs[147]);
    assign layer0_outputs[4808] = ~(inputs[38]);
    assign layer0_outputs[4809] = (inputs[184]) & ~(inputs[201]);
    assign layer0_outputs[4810] = ~(inputs[135]) | (inputs[1]);
    assign layer0_outputs[4811] = ~(inputs[166]);
    assign layer0_outputs[4812] = ~(inputs[110]);
    assign layer0_outputs[4813] = 1'b1;
    assign layer0_outputs[4814] = (inputs[61]) | (inputs[50]);
    assign layer0_outputs[4815] = (inputs[42]) & ~(inputs[3]);
    assign layer0_outputs[4816] = ~(inputs[191]);
    assign layer0_outputs[4817] = inputs[180];
    assign layer0_outputs[4818] = ~((inputs[185]) & (inputs[217]));
    assign layer0_outputs[4819] = (inputs[102]) & (inputs[157]);
    assign layer0_outputs[4820] = 1'b1;
    assign layer0_outputs[4821] = ~(inputs[234]);
    assign layer0_outputs[4822] = inputs[239];
    assign layer0_outputs[4823] = ~(inputs[132]) | (inputs[157]);
    assign layer0_outputs[4824] = (inputs[216]) & (inputs[199]);
    assign layer0_outputs[4825] = inputs[132];
    assign layer0_outputs[4826] = inputs[235];
    assign layer0_outputs[4827] = ~(inputs[237]) | (inputs[250]);
    assign layer0_outputs[4828] = (inputs[184]) & ~(inputs[67]);
    assign layer0_outputs[4829] = ~(inputs[206]) | (inputs[184]);
    assign layer0_outputs[4830] = (inputs[209]) & ~(inputs[65]);
    assign layer0_outputs[4831] = ~(inputs[105]);
    assign layer0_outputs[4832] = ~(inputs[147]) | (inputs[57]);
    assign layer0_outputs[4833] = ~(inputs[80]);
    assign layer0_outputs[4834] = (inputs[201]) | (inputs[37]);
    assign layer0_outputs[4835] = ~((inputs[67]) ^ (inputs[221]));
    assign layer0_outputs[4836] = ~((inputs[21]) ^ (inputs[229]));
    assign layer0_outputs[4837] = inputs[165];
    assign layer0_outputs[4838] = 1'b1;
    assign layer0_outputs[4839] = (inputs[179]) | (inputs[17]);
    assign layer0_outputs[4840] = inputs[105];
    assign layer0_outputs[4841] = ~((inputs[85]) | (inputs[147]));
    assign layer0_outputs[4842] = ~(inputs[157]);
    assign layer0_outputs[4843] = ~(inputs[47]);
    assign layer0_outputs[4844] = ~(inputs[80]);
    assign layer0_outputs[4845] = (inputs[11]) & ~(inputs[202]);
    assign layer0_outputs[4846] = 1'b1;
    assign layer0_outputs[4847] = inputs[4];
    assign layer0_outputs[4848] = 1'b1;
    assign layer0_outputs[4849] = ~((inputs[31]) ^ (inputs[159]));
    assign layer0_outputs[4850] = ~(inputs[83]) | (inputs[184]);
    assign layer0_outputs[4851] = (inputs[239]) ^ (inputs[144]);
    assign layer0_outputs[4852] = 1'b1;
    assign layer0_outputs[4853] = ~(inputs[183]) | (inputs[177]);
    assign layer0_outputs[4854] = (inputs[47]) | (inputs[224]);
    assign layer0_outputs[4855] = (inputs[49]) & (inputs[114]);
    assign layer0_outputs[4856] = ~((inputs[113]) | (inputs[114]));
    assign layer0_outputs[4857] = ~(inputs[74]);
    assign layer0_outputs[4858] = (inputs[7]) & ~(inputs[143]);
    assign layer0_outputs[4859] = ~((inputs[163]) | (inputs[223]));
    assign layer0_outputs[4860] = 1'b0;
    assign layer0_outputs[4861] = (inputs[109]) | (inputs[185]);
    assign layer0_outputs[4862] = ~(inputs[46]);
    assign layer0_outputs[4863] = ~(inputs[18]) | (inputs[96]);
    assign layer0_outputs[4864] = ~(inputs[134]);
    assign layer0_outputs[4865] = ~((inputs[106]) ^ (inputs[204]));
    assign layer0_outputs[4866] = ~((inputs[127]) ^ (inputs[193]));
    assign layer0_outputs[4867] = (inputs[179]) | (inputs[234]);
    assign layer0_outputs[4868] = ~((inputs[154]) & (inputs[66]));
    assign layer0_outputs[4869] = ~((inputs[143]) | (inputs[182]));
    assign layer0_outputs[4870] = ~((inputs[95]) | (inputs[224]));
    assign layer0_outputs[4871] = ~((inputs[213]) | (inputs[125]));
    assign layer0_outputs[4872] = (inputs[65]) | (inputs[82]);
    assign layer0_outputs[4873] = ~((inputs[33]) & (inputs[82]));
    assign layer0_outputs[4874] = ~(inputs[186]) | (inputs[6]);
    assign layer0_outputs[4875] = (inputs[39]) | (inputs[147]);
    assign layer0_outputs[4876] = (inputs[6]) | (inputs[111]);
    assign layer0_outputs[4877] = (inputs[185]) & ~(inputs[16]);
    assign layer0_outputs[4878] = inputs[234];
    assign layer0_outputs[4879] = (inputs[66]) ^ (inputs[168]);
    assign layer0_outputs[4880] = ~(inputs[30]) | (inputs[79]);
    assign layer0_outputs[4881] = inputs[37];
    assign layer0_outputs[4882] = ~(inputs[8]);
    assign layer0_outputs[4883] = ~(inputs[153]) | (inputs[34]);
    assign layer0_outputs[4884] = 1'b0;
    assign layer0_outputs[4885] = (inputs[44]) & ~(inputs[213]);
    assign layer0_outputs[4886] = (inputs[132]) & ~(inputs[94]);
    assign layer0_outputs[4887] = (inputs[129]) ^ (inputs[188]);
    assign layer0_outputs[4888] = ~((inputs[23]) & (inputs[182]));
    assign layer0_outputs[4889] = ~((inputs[126]) | (inputs[184]));
    assign layer0_outputs[4890] = ~(inputs[120]);
    assign layer0_outputs[4891] = ~(inputs[13]);
    assign layer0_outputs[4892] = (inputs[124]) | (inputs[101]);
    assign layer0_outputs[4893] = ~((inputs[219]) | (inputs[230]));
    assign layer0_outputs[4894] = (inputs[117]) & ~(inputs[4]);
    assign layer0_outputs[4895] = ~((inputs[244]) | (inputs[234]));
    assign layer0_outputs[4896] = ~(inputs[218]);
    assign layer0_outputs[4897] = 1'b0;
    assign layer0_outputs[4898] = (inputs[237]) | (inputs[109]);
    assign layer0_outputs[4899] = (inputs[139]) & ~(inputs[69]);
    assign layer0_outputs[4900] = ~((inputs[158]) ^ (inputs[84]));
    assign layer0_outputs[4901] = ~((inputs[167]) | (inputs[183]));
    assign layer0_outputs[4902] = inputs[71];
    assign layer0_outputs[4903] = inputs[124];
    assign layer0_outputs[4904] = ~(inputs[235]);
    assign layer0_outputs[4905] = ~(inputs[124]) | (inputs[238]);
    assign layer0_outputs[4906] = (inputs[12]) ^ (inputs[128]);
    assign layer0_outputs[4907] = ~(inputs[50]);
    assign layer0_outputs[4908] = ~((inputs[153]) | (inputs[47]));
    assign layer0_outputs[4909] = 1'b1;
    assign layer0_outputs[4910] = (inputs[134]) ^ (inputs[224]);
    assign layer0_outputs[4911] = ~(inputs[144]);
    assign layer0_outputs[4912] = inputs[182];
    assign layer0_outputs[4913] = 1'b1;
    assign layer0_outputs[4914] = (inputs[205]) | (inputs[206]);
    assign layer0_outputs[4915] = (inputs[200]) & ~(inputs[1]);
    assign layer0_outputs[4916] = inputs[168];
    assign layer0_outputs[4917] = inputs[139];
    assign layer0_outputs[4918] = ~(inputs[21]);
    assign layer0_outputs[4919] = (inputs[225]) | (inputs[89]);
    assign layer0_outputs[4920] = (inputs[162]) | (inputs[160]);
    assign layer0_outputs[4921] = ~(inputs[246]);
    assign layer0_outputs[4922] = (inputs[212]) & ~(inputs[233]);
    assign layer0_outputs[4923] = inputs[74];
    assign layer0_outputs[4924] = ~(inputs[8]);
    assign layer0_outputs[4925] = 1'b0;
    assign layer0_outputs[4926] = ~((inputs[38]) ^ (inputs[68]));
    assign layer0_outputs[4927] = (inputs[146]) | (inputs[93]);
    assign layer0_outputs[4928] = inputs[112];
    assign layer0_outputs[4929] = ~(inputs[5]) | (inputs[27]);
    assign layer0_outputs[4930] = inputs[218];
    assign layer0_outputs[4931] = ~((inputs[195]) | (inputs[192]));
    assign layer0_outputs[4932] = (inputs[142]) ^ (inputs[175]);
    assign layer0_outputs[4933] = (inputs[189]) & ~(inputs[26]);
    assign layer0_outputs[4934] = inputs[23];
    assign layer0_outputs[4935] = ~(inputs[31]) | (inputs[217]);
    assign layer0_outputs[4936] = ~((inputs[56]) ^ (inputs[43]));
    assign layer0_outputs[4937] = inputs[219];
    assign layer0_outputs[4938] = ~((inputs[6]) ^ (inputs[172]));
    assign layer0_outputs[4939] = ~(inputs[173]);
    assign layer0_outputs[4940] = inputs[183];
    assign layer0_outputs[4941] = inputs[144];
    assign layer0_outputs[4942] = ~((inputs[58]) & (inputs[95]));
    assign layer0_outputs[4943] = ~((inputs[27]) ^ (inputs[104]));
    assign layer0_outputs[4944] = (inputs[5]) & (inputs[204]);
    assign layer0_outputs[4945] = (inputs[145]) & ~(inputs[53]);
    assign layer0_outputs[4946] = inputs[38];
    assign layer0_outputs[4947] = (inputs[19]) & ~(inputs[255]);
    assign layer0_outputs[4948] = inputs[67];
    assign layer0_outputs[4949] = (inputs[74]) & ~(inputs[179]);
    assign layer0_outputs[4950] = ~((inputs[1]) & (inputs[215]));
    assign layer0_outputs[4951] = (inputs[153]) & ~(inputs[177]);
    assign layer0_outputs[4952] = ~((inputs[53]) ^ (inputs[20]));
    assign layer0_outputs[4953] = ~(inputs[245]);
    assign layer0_outputs[4954] = ~(inputs[179]) | (inputs[253]);
    assign layer0_outputs[4955] = ~(inputs[46]) | (inputs[9]);
    assign layer0_outputs[4956] = 1'b0;
    assign layer0_outputs[4957] = ~((inputs[2]) ^ (inputs[115]));
    assign layer0_outputs[4958] = ~((inputs[163]) | (inputs[239]));
    assign layer0_outputs[4959] = inputs[155];
    assign layer0_outputs[4960] = (inputs[125]) & ~(inputs[238]);
    assign layer0_outputs[4961] = inputs[184];
    assign layer0_outputs[4962] = inputs[25];
    assign layer0_outputs[4963] = ~((inputs[205]) | (inputs[57]));
    assign layer0_outputs[4964] = (inputs[12]) & ~(inputs[222]);
    assign layer0_outputs[4965] = (inputs[33]) ^ (inputs[189]);
    assign layer0_outputs[4966] = ~((inputs[69]) & (inputs[33]));
    assign layer0_outputs[4967] = ~((inputs[176]) ^ (inputs[33]));
    assign layer0_outputs[4968] = (inputs[112]) | (inputs[187]);
    assign layer0_outputs[4969] = inputs[102];
    assign layer0_outputs[4970] = ~(inputs[182]);
    assign layer0_outputs[4971] = inputs[246];
    assign layer0_outputs[4972] = ~((inputs[25]) ^ (inputs[3]));
    assign layer0_outputs[4973] = (inputs[220]) | (inputs[208]);
    assign layer0_outputs[4974] = ~(inputs[206]);
    assign layer0_outputs[4975] = inputs[100];
    assign layer0_outputs[4976] = ~((inputs[255]) | (inputs[123]));
    assign layer0_outputs[4977] = inputs[83];
    assign layer0_outputs[4978] = ~((inputs[139]) & (inputs[155]));
    assign layer0_outputs[4979] = ~(inputs[102]) | (inputs[117]);
    assign layer0_outputs[4980] = (inputs[33]) | (inputs[252]);
    assign layer0_outputs[4981] = inputs[176];
    assign layer0_outputs[4982] = ~(inputs[153]);
    assign layer0_outputs[4983] = (inputs[233]) & (inputs[15]);
    assign layer0_outputs[4984] = ~((inputs[158]) ^ (inputs[255]));
    assign layer0_outputs[4985] = inputs[0];
    assign layer0_outputs[4986] = ~((inputs[112]) ^ (inputs[232]));
    assign layer0_outputs[4987] = ~((inputs[212]) & (inputs[234]));
    assign layer0_outputs[4988] = inputs[50];
    assign layer0_outputs[4989] = inputs[141];
    assign layer0_outputs[4990] = inputs[162];
    assign layer0_outputs[4991] = ~(inputs[78]);
    assign layer0_outputs[4992] = inputs[175];
    assign layer0_outputs[4993] = inputs[132];
    assign layer0_outputs[4994] = ~((inputs[12]) ^ (inputs[22]));
    assign layer0_outputs[4995] = (inputs[114]) & ~(inputs[207]);
    assign layer0_outputs[4996] = ~(inputs[113]);
    assign layer0_outputs[4997] = (inputs[24]) & ~(inputs[142]);
    assign layer0_outputs[4998] = ~((inputs[198]) ^ (inputs[61]));
    assign layer0_outputs[4999] = ~((inputs[80]) | (inputs[251]));
    assign layer0_outputs[5000] = ~((inputs[213]) | (inputs[243]));
    assign layer0_outputs[5001] = ~(inputs[86]) | (inputs[70]);
    assign layer0_outputs[5002] = (inputs[116]) & ~(inputs[34]);
    assign layer0_outputs[5003] = ~((inputs[89]) ^ (inputs[228]));
    assign layer0_outputs[5004] = inputs[86];
    assign layer0_outputs[5005] = 1'b1;
    assign layer0_outputs[5006] = ~(inputs[52]);
    assign layer0_outputs[5007] = (inputs[55]) & (inputs[40]);
    assign layer0_outputs[5008] = (inputs[173]) ^ (inputs[19]);
    assign layer0_outputs[5009] = (inputs[234]) | (inputs[3]);
    assign layer0_outputs[5010] = (inputs[198]) & (inputs[95]);
    assign layer0_outputs[5011] = inputs[109];
    assign layer0_outputs[5012] = ~((inputs[125]) ^ (inputs[125]));
    assign layer0_outputs[5013] = inputs[165];
    assign layer0_outputs[5014] = inputs[199];
    assign layer0_outputs[5015] = inputs[105];
    assign layer0_outputs[5016] = ~(inputs[61]);
    assign layer0_outputs[5017] = ~((inputs[220]) & (inputs[30]));
    assign layer0_outputs[5018] = ~((inputs[23]) ^ (inputs[85]));
    assign layer0_outputs[5019] = 1'b0;
    assign layer0_outputs[5020] = (inputs[116]) | (inputs[249]);
    assign layer0_outputs[5021] = 1'b0;
    assign layer0_outputs[5022] = inputs[54];
    assign layer0_outputs[5023] = inputs[35];
    assign layer0_outputs[5024] = ~(inputs[75]) | (inputs[227]);
    assign layer0_outputs[5025] = ~((inputs[77]) ^ (inputs[17]));
    assign layer0_outputs[5026] = ~((inputs[8]) & (inputs[132]));
    assign layer0_outputs[5027] = inputs[157];
    assign layer0_outputs[5028] = ~(inputs[7]) | (inputs[8]);
    assign layer0_outputs[5029] = ~(inputs[148]);
    assign layer0_outputs[5030] = ~(inputs[90]) | (inputs[221]);
    assign layer0_outputs[5031] = ~(inputs[161]);
    assign layer0_outputs[5032] = (inputs[133]) | (inputs[14]);
    assign layer0_outputs[5033] = ~((inputs[168]) | (inputs[111]));
    assign layer0_outputs[5034] = ~((inputs[165]) & (inputs[245]));
    assign layer0_outputs[5035] = ~(inputs[124]);
    assign layer0_outputs[5036] = inputs[23];
    assign layer0_outputs[5037] = ~((inputs[189]) | (inputs[249]));
    assign layer0_outputs[5038] = ~((inputs[72]) | (inputs[206]));
    assign layer0_outputs[5039] = (inputs[100]) | (inputs[195]);
    assign layer0_outputs[5040] = ~(inputs[59]) | (inputs[205]);
    assign layer0_outputs[5041] = inputs[184];
    assign layer0_outputs[5042] = ~((inputs[144]) ^ (inputs[65]));
    assign layer0_outputs[5043] = ~(inputs[202]);
    assign layer0_outputs[5044] = inputs[23];
    assign layer0_outputs[5045] = ~(inputs[138]);
    assign layer0_outputs[5046] = (inputs[107]) & ~(inputs[133]);
    assign layer0_outputs[5047] = ~((inputs[41]) & (inputs[45]));
    assign layer0_outputs[5048] = (inputs[13]) & ~(inputs[245]);
    assign layer0_outputs[5049] = ~(inputs[87]) | (inputs[37]);
    assign layer0_outputs[5050] = (inputs[106]) & ~(inputs[47]);
    assign layer0_outputs[5051] = (inputs[26]) | (inputs[9]);
    assign layer0_outputs[5052] = ~(inputs[18]) | (inputs[141]);
    assign layer0_outputs[5053] = ~((inputs[115]) & (inputs[131]));
    assign layer0_outputs[5054] = ~((inputs[90]) | (inputs[146]));
    assign layer0_outputs[5055] = ~(inputs[219]);
    assign layer0_outputs[5056] = ~(inputs[88]) | (inputs[80]);
    assign layer0_outputs[5057] = ~(inputs[148]);
    assign layer0_outputs[5058] = (inputs[163]) ^ (inputs[95]);
    assign layer0_outputs[5059] = (inputs[90]) & ~(inputs[162]);
    assign layer0_outputs[5060] = (inputs[117]) & (inputs[255]);
    assign layer0_outputs[5061] = (inputs[36]) | (inputs[51]);
    assign layer0_outputs[5062] = (inputs[208]) | (inputs[205]);
    assign layer0_outputs[5063] = ~(inputs[23]);
    assign layer0_outputs[5064] = (inputs[119]) & ~(inputs[170]);
    assign layer0_outputs[5065] = inputs[77];
    assign layer0_outputs[5066] = ~(inputs[180]) | (inputs[89]);
    assign layer0_outputs[5067] = (inputs[1]) | (inputs[151]);
    assign layer0_outputs[5068] = inputs[35];
    assign layer0_outputs[5069] = (inputs[202]) & ~(inputs[97]);
    assign layer0_outputs[5070] = ~(inputs[232]);
    assign layer0_outputs[5071] = (inputs[210]) & ~(inputs[80]);
    assign layer0_outputs[5072] = (inputs[152]) ^ (inputs[255]);
    assign layer0_outputs[5073] = ~(inputs[151]);
    assign layer0_outputs[5074] = ~((inputs[150]) | (inputs[137]));
    assign layer0_outputs[5075] = (inputs[12]) ^ (inputs[21]);
    assign layer0_outputs[5076] = ~((inputs[175]) ^ (inputs[246]));
    assign layer0_outputs[5077] = inputs[215];
    assign layer0_outputs[5078] = ~(inputs[131]);
    assign layer0_outputs[5079] = (inputs[148]) & ~(inputs[145]);
    assign layer0_outputs[5080] = (inputs[167]) ^ (inputs[152]);
    assign layer0_outputs[5081] = inputs[124];
    assign layer0_outputs[5082] = ~((inputs[102]) & (inputs[232]));
    assign layer0_outputs[5083] = ~((inputs[33]) | (inputs[211]));
    assign layer0_outputs[5084] = (inputs[186]) | (inputs[31]);
    assign layer0_outputs[5085] = (inputs[83]) & ~(inputs[117]);
    assign layer0_outputs[5086] = ~(inputs[58]) | (inputs[32]);
    assign layer0_outputs[5087] = ~((inputs[94]) | (inputs[44]));
    assign layer0_outputs[5088] = (inputs[173]) & ~(inputs[255]);
    assign layer0_outputs[5089] = ~(inputs[224]) | (inputs[15]);
    assign layer0_outputs[5090] = inputs[12];
    assign layer0_outputs[5091] = ~((inputs[66]) ^ (inputs[226]));
    assign layer0_outputs[5092] = (inputs[59]) & ~(inputs[175]);
    assign layer0_outputs[5093] = (inputs[12]) | (inputs[185]);
    assign layer0_outputs[5094] = ~((inputs[217]) ^ (inputs[238]));
    assign layer0_outputs[5095] = ~(inputs[105]);
    assign layer0_outputs[5096] = (inputs[172]) ^ (inputs[36]);
    assign layer0_outputs[5097] = 1'b0;
    assign layer0_outputs[5098] = (inputs[81]) & (inputs[35]);
    assign layer0_outputs[5099] = inputs[157];
    assign layer0_outputs[5100] = (inputs[146]) & ~(inputs[63]);
    assign layer0_outputs[5101] = ~(inputs[19]);
    assign layer0_outputs[5102] = ~(inputs[129]);
    assign layer0_outputs[5103] = (inputs[52]) | (inputs[221]);
    assign layer0_outputs[5104] = ~(inputs[12]) | (inputs[193]);
    assign layer0_outputs[5105] = inputs[93];
    assign layer0_outputs[5106] = (inputs[40]) & ~(inputs[134]);
    assign layer0_outputs[5107] = ~(inputs[45]);
    assign layer0_outputs[5108] = ~(inputs[30]) | (inputs[246]);
    assign layer0_outputs[5109] = (inputs[70]) & (inputs[41]);
    assign layer0_outputs[5110] = ~((inputs[232]) | (inputs[157]));
    assign layer0_outputs[5111] = ~((inputs[78]) | (inputs[98]));
    assign layer0_outputs[5112] = ~(inputs[198]);
    assign layer0_outputs[5113] = ~((inputs[154]) | (inputs[221]));
    assign layer0_outputs[5114] = (inputs[42]) | (inputs[108]);
    assign layer0_outputs[5115] = inputs[195];
    assign layer0_outputs[5116] = ~(inputs[239]);
    assign layer0_outputs[5117] = ~((inputs[241]) | (inputs[171]));
    assign layer0_outputs[5118] = (inputs[65]) & (inputs[4]);
    assign layer0_outputs[5119] = inputs[239];
    assign layer0_outputs[5120] = inputs[24];
    assign layer0_outputs[5121] = (inputs[65]) ^ (inputs[74]);
    assign layer0_outputs[5122] = (inputs[161]) & ~(inputs[124]);
    assign layer0_outputs[5123] = ~(inputs[231]);
    assign layer0_outputs[5124] = inputs[107];
    assign layer0_outputs[5125] = ~(inputs[166]) | (inputs[91]);
    assign layer0_outputs[5126] = ~(inputs[118]) | (inputs[24]);
    assign layer0_outputs[5127] = (inputs[33]) & (inputs[105]);
    assign layer0_outputs[5128] = ~(inputs[204]) | (inputs[168]);
    assign layer0_outputs[5129] = ~(inputs[7]);
    assign layer0_outputs[5130] = ~((inputs[84]) ^ (inputs[132]));
    assign layer0_outputs[5131] = ~(inputs[105]);
    assign layer0_outputs[5132] = ~((inputs[85]) | (inputs[144]));
    assign layer0_outputs[5133] = (inputs[229]) ^ (inputs[197]);
    assign layer0_outputs[5134] = ~(inputs[63]);
    assign layer0_outputs[5135] = (inputs[86]) & ~(inputs[2]);
    assign layer0_outputs[5136] = (inputs[142]) | (inputs[147]);
    assign layer0_outputs[5137] = (inputs[198]) & ~(inputs[87]);
    assign layer0_outputs[5138] = ~((inputs[134]) | (inputs[81]));
    assign layer0_outputs[5139] = ~(inputs[229]);
    assign layer0_outputs[5140] = ~(inputs[127]);
    assign layer0_outputs[5141] = ~((inputs[176]) ^ (inputs[93]));
    assign layer0_outputs[5142] = ~(inputs[133]) | (inputs[224]);
    assign layer0_outputs[5143] = ~((inputs[47]) | (inputs[169]));
    assign layer0_outputs[5144] = ~(inputs[45]) | (inputs[48]);
    assign layer0_outputs[5145] = ~(inputs[48]) | (inputs[24]);
    assign layer0_outputs[5146] = (inputs[8]) | (inputs[204]);
    assign layer0_outputs[5147] = (inputs[235]) | (inputs[171]);
    assign layer0_outputs[5148] = inputs[243];
    assign layer0_outputs[5149] = (inputs[104]) ^ (inputs[18]);
    assign layer0_outputs[5150] = 1'b1;
    assign layer0_outputs[5151] = (inputs[54]) & ~(inputs[192]);
    assign layer0_outputs[5152] = (inputs[135]) & ~(inputs[154]);
    assign layer0_outputs[5153] = ~(inputs[255]) | (inputs[31]);
    assign layer0_outputs[5154] = ~(inputs[82]);
    assign layer0_outputs[5155] = (inputs[182]) & ~(inputs[91]);
    assign layer0_outputs[5156] = inputs[243];
    assign layer0_outputs[5157] = 1'b0;
    assign layer0_outputs[5158] = ~(inputs[171]);
    assign layer0_outputs[5159] = inputs[75];
    assign layer0_outputs[5160] = (inputs[247]) & ~(inputs[68]);
    assign layer0_outputs[5161] = ~(inputs[107]);
    assign layer0_outputs[5162] = ~((inputs[210]) | (inputs[223]));
    assign layer0_outputs[5163] = ~(inputs[39]);
    assign layer0_outputs[5164] = inputs[202];
    assign layer0_outputs[5165] = inputs[83];
    assign layer0_outputs[5166] = (inputs[246]) & ~(inputs[91]);
    assign layer0_outputs[5167] = (inputs[223]) & ~(inputs[221]);
    assign layer0_outputs[5168] = (inputs[85]) & ~(inputs[243]);
    assign layer0_outputs[5169] = inputs[123];
    assign layer0_outputs[5170] = (inputs[200]) & ~(inputs[88]);
    assign layer0_outputs[5171] = inputs[100];
    assign layer0_outputs[5172] = 1'b0;
    assign layer0_outputs[5173] = ~(inputs[227]) | (inputs[133]);
    assign layer0_outputs[5174] = (inputs[68]) | (inputs[75]);
    assign layer0_outputs[5175] = inputs[86];
    assign layer0_outputs[5176] = ~(inputs[170]) | (inputs[65]);
    assign layer0_outputs[5177] = ~(inputs[45]) | (inputs[169]);
    assign layer0_outputs[5178] = ~(inputs[227]);
    assign layer0_outputs[5179] = ~((inputs[95]) | (inputs[11]));
    assign layer0_outputs[5180] = ~((inputs[33]) | (inputs[35]));
    assign layer0_outputs[5181] = ~(inputs[70]) | (inputs[119]);
    assign layer0_outputs[5182] = ~(inputs[24]);
    assign layer0_outputs[5183] = ~(inputs[180]);
    assign layer0_outputs[5184] = ~(inputs[102]);
    assign layer0_outputs[5185] = inputs[152];
    assign layer0_outputs[5186] = ~((inputs[111]) ^ (inputs[31]));
    assign layer0_outputs[5187] = (inputs[254]) | (inputs[222]);
    assign layer0_outputs[5188] = ~((inputs[121]) | (inputs[166]));
    assign layer0_outputs[5189] = ~(inputs[100]);
    assign layer0_outputs[5190] = ~((inputs[17]) | (inputs[88]));
    assign layer0_outputs[5191] = 1'b0;
    assign layer0_outputs[5192] = (inputs[98]) | (inputs[168]);
    assign layer0_outputs[5193] = (inputs[81]) ^ (inputs[19]);
    assign layer0_outputs[5194] = (inputs[208]) ^ (inputs[29]);
    assign layer0_outputs[5195] = inputs[134];
    assign layer0_outputs[5196] = ~(inputs[116]);
    assign layer0_outputs[5197] = (inputs[181]) | (inputs[102]);
    assign layer0_outputs[5198] = ~((inputs[194]) | (inputs[125]));
    assign layer0_outputs[5199] = ~((inputs[21]) | (inputs[124]));
    assign layer0_outputs[5200] = (inputs[253]) | (inputs[205]);
    assign layer0_outputs[5201] = ~(inputs[108]) | (inputs[175]);
    assign layer0_outputs[5202] = ~(inputs[6]) | (inputs[13]);
    assign layer0_outputs[5203] = ~((inputs[223]) | (inputs[159]));
    assign layer0_outputs[5204] = ~(inputs[36]);
    assign layer0_outputs[5205] = inputs[78];
    assign layer0_outputs[5206] = ~(inputs[153]);
    assign layer0_outputs[5207] = (inputs[53]) | (inputs[55]);
    assign layer0_outputs[5208] = (inputs[63]) & ~(inputs[45]);
    assign layer0_outputs[5209] = (inputs[66]) | (inputs[48]);
    assign layer0_outputs[5210] = (inputs[116]) ^ (inputs[98]);
    assign layer0_outputs[5211] = ~(inputs[200]);
    assign layer0_outputs[5212] = ~((inputs[81]) | (inputs[103]));
    assign layer0_outputs[5213] = ~(inputs[169]) | (inputs[72]);
    assign layer0_outputs[5214] = ~(inputs[186]) | (inputs[8]);
    assign layer0_outputs[5215] = (inputs[159]) & ~(inputs[155]);
    assign layer0_outputs[5216] = inputs[213];
    assign layer0_outputs[5217] = ~(inputs[90]) | (inputs[168]);
    assign layer0_outputs[5218] = inputs[55];
    assign layer0_outputs[5219] = ~(inputs[13]);
    assign layer0_outputs[5220] = ~(inputs[216]);
    assign layer0_outputs[5221] = ~(inputs[50]) | (inputs[199]);
    assign layer0_outputs[5222] = ~(inputs[224]);
    assign layer0_outputs[5223] = ~(inputs[144]);
    assign layer0_outputs[5224] = (inputs[80]) | (inputs[124]);
    assign layer0_outputs[5225] = (inputs[92]) & ~(inputs[221]);
    assign layer0_outputs[5226] = ~(inputs[190]);
    assign layer0_outputs[5227] = ~(inputs[93]);
    assign layer0_outputs[5228] = 1'b1;
    assign layer0_outputs[5229] = inputs[227];
    assign layer0_outputs[5230] = ~(inputs[214]);
    assign layer0_outputs[5231] = 1'b1;
    assign layer0_outputs[5232] = (inputs[68]) ^ (inputs[51]);
    assign layer0_outputs[5233] = ~((inputs[156]) | (inputs[116]));
    assign layer0_outputs[5234] = ~(inputs[243]) | (inputs[57]);
    assign layer0_outputs[5235] = inputs[162];
    assign layer0_outputs[5236] = (inputs[24]) & ~(inputs[14]);
    assign layer0_outputs[5237] = 1'b1;
    assign layer0_outputs[5238] = ~(inputs[38]) | (inputs[210]);
    assign layer0_outputs[5239] = inputs[24];
    assign layer0_outputs[5240] = (inputs[95]) ^ (inputs[225]);
    assign layer0_outputs[5241] = (inputs[183]) & ~(inputs[155]);
    assign layer0_outputs[5242] = ~((inputs[145]) ^ (inputs[118]));
    assign layer0_outputs[5243] = 1'b1;
    assign layer0_outputs[5244] = (inputs[190]) ^ (inputs[13]);
    assign layer0_outputs[5245] = ~((inputs[102]) ^ (inputs[182]));
    assign layer0_outputs[5246] = (inputs[81]) | (inputs[82]);
    assign layer0_outputs[5247] = ~((inputs[81]) & (inputs[207]));
    assign layer0_outputs[5248] = ~((inputs[37]) ^ (inputs[64]));
    assign layer0_outputs[5249] = ~(inputs[206]);
    assign layer0_outputs[5250] = ~((inputs[37]) ^ (inputs[146]));
    assign layer0_outputs[5251] = ~(inputs[83]) | (inputs[174]);
    assign layer0_outputs[5252] = ~(inputs[156]);
    assign layer0_outputs[5253] = ~((inputs[86]) ^ (inputs[126]));
    assign layer0_outputs[5254] = inputs[56];
    assign layer0_outputs[5255] = ~(inputs[136]) | (inputs[202]);
    assign layer0_outputs[5256] = 1'b1;
    assign layer0_outputs[5257] = inputs[224];
    assign layer0_outputs[5258] = ~((inputs[84]) | (inputs[148]));
    assign layer0_outputs[5259] = ~((inputs[115]) | (inputs[131]));
    assign layer0_outputs[5260] = (inputs[151]) & ~(inputs[140]);
    assign layer0_outputs[5261] = ~(inputs[80]);
    assign layer0_outputs[5262] = ~(inputs[32]) | (inputs[32]);
    assign layer0_outputs[5263] = (inputs[60]) | (inputs[79]);
    assign layer0_outputs[5264] = (inputs[68]) & (inputs[24]);
    assign layer0_outputs[5265] = (inputs[232]) | (inputs[67]);
    assign layer0_outputs[5266] = (inputs[80]) ^ (inputs[110]);
    assign layer0_outputs[5267] = ~(inputs[174]) | (inputs[186]);
    assign layer0_outputs[5268] = ~((inputs[106]) & (inputs[137]));
    assign layer0_outputs[5269] = (inputs[238]) | (inputs[238]);
    assign layer0_outputs[5270] = (inputs[226]) & ~(inputs[217]);
    assign layer0_outputs[5271] = ~(inputs[201]) | (inputs[207]);
    assign layer0_outputs[5272] = inputs[225];
    assign layer0_outputs[5273] = ~((inputs[238]) | (inputs[106]));
    assign layer0_outputs[5274] = (inputs[136]) | (inputs[122]);
    assign layer0_outputs[5275] = ~(inputs[103]);
    assign layer0_outputs[5276] = (inputs[10]) & ~(inputs[31]);
    assign layer0_outputs[5277] = ~(inputs[221]);
    assign layer0_outputs[5278] = ~(inputs[237]);
    assign layer0_outputs[5279] = inputs[121];
    assign layer0_outputs[5280] = (inputs[129]) ^ (inputs[127]);
    assign layer0_outputs[5281] = (inputs[21]) & ~(inputs[205]);
    assign layer0_outputs[5282] = (inputs[167]) & ~(inputs[128]);
    assign layer0_outputs[5283] = ~(inputs[177]);
    assign layer0_outputs[5284] = ~(inputs[32]) | (inputs[38]);
    assign layer0_outputs[5285] = inputs[51];
    assign layer0_outputs[5286] = ~((inputs[235]) ^ (inputs[186]));
    assign layer0_outputs[5287] = ~(inputs[247]);
    assign layer0_outputs[5288] = (inputs[95]) | (inputs[102]);
    assign layer0_outputs[5289] = ~((inputs[124]) ^ (inputs[7]));
    assign layer0_outputs[5290] = ~(inputs[58]) | (inputs[13]);
    assign layer0_outputs[5291] = inputs[83];
    assign layer0_outputs[5292] = ~(inputs[110]);
    assign layer0_outputs[5293] = (inputs[168]) | (inputs[126]);
    assign layer0_outputs[5294] = ~(inputs[56]);
    assign layer0_outputs[5295] = ~(inputs[216]) | (inputs[145]);
    assign layer0_outputs[5296] = ~((inputs[38]) & (inputs[198]));
    assign layer0_outputs[5297] = 1'b0;
    assign layer0_outputs[5298] = inputs[60];
    assign layer0_outputs[5299] = ~(inputs[14]) | (inputs[127]);
    assign layer0_outputs[5300] = inputs[50];
    assign layer0_outputs[5301] = ~(inputs[123]);
    assign layer0_outputs[5302] = ~(inputs[211]) | (inputs[205]);
    assign layer0_outputs[5303] = ~((inputs[232]) ^ (inputs[16]));
    assign layer0_outputs[5304] = ~((inputs[168]) | (inputs[97]));
    assign layer0_outputs[5305] = ~(inputs[156]) | (inputs[9]);
    assign layer0_outputs[5306] = (inputs[124]) & ~(inputs[112]);
    assign layer0_outputs[5307] = (inputs[148]) ^ (inputs[2]);
    assign layer0_outputs[5308] = (inputs[157]) & ~(inputs[102]);
    assign layer0_outputs[5309] = ~((inputs[32]) ^ (inputs[76]));
    assign layer0_outputs[5310] = ~(inputs[83]) | (inputs[161]);
    assign layer0_outputs[5311] = ~(inputs[122]) | (inputs[223]);
    assign layer0_outputs[5312] = (inputs[87]) & ~(inputs[48]);
    assign layer0_outputs[5313] = ~(inputs[41]) | (inputs[60]);
    assign layer0_outputs[5314] = inputs[39];
    assign layer0_outputs[5315] = ~((inputs[161]) | (inputs[243]));
    assign layer0_outputs[5316] = (inputs[208]) & ~(inputs[176]);
    assign layer0_outputs[5317] = (inputs[5]) & ~(inputs[153]);
    assign layer0_outputs[5318] = inputs[40];
    assign layer0_outputs[5319] = ~(inputs[151]);
    assign layer0_outputs[5320] = (inputs[69]) & ~(inputs[172]);
    assign layer0_outputs[5321] = (inputs[255]) & ~(inputs[148]);
    assign layer0_outputs[5322] = ~((inputs[155]) ^ (inputs[190]));
    assign layer0_outputs[5323] = ~((inputs[223]) ^ (inputs[237]));
    assign layer0_outputs[5324] = inputs[166];
    assign layer0_outputs[5325] = (inputs[97]) | (inputs[185]);
    assign layer0_outputs[5326] = ~(inputs[38]) | (inputs[13]);
    assign layer0_outputs[5327] = inputs[123];
    assign layer0_outputs[5328] = ~((inputs[236]) & (inputs[241]));
    assign layer0_outputs[5329] = ~(inputs[176]) | (inputs[146]);
    assign layer0_outputs[5330] = inputs[167];
    assign layer0_outputs[5331] = ~(inputs[24]);
    assign layer0_outputs[5332] = (inputs[185]) ^ (inputs[136]);
    assign layer0_outputs[5333] = ~(inputs[183]);
    assign layer0_outputs[5334] = (inputs[19]) & (inputs[99]);
    assign layer0_outputs[5335] = ~((inputs[92]) ^ (inputs[33]));
    assign layer0_outputs[5336] = ~(inputs[193]);
    assign layer0_outputs[5337] = (inputs[127]) & ~(inputs[228]);
    assign layer0_outputs[5338] = inputs[84];
    assign layer0_outputs[5339] = ~(inputs[9]);
    assign layer0_outputs[5340] = ~((inputs[75]) | (inputs[28]));
    assign layer0_outputs[5341] = ~((inputs[224]) | (inputs[4]));
    assign layer0_outputs[5342] = ~((inputs[160]) ^ (inputs[100]));
    assign layer0_outputs[5343] = ~(inputs[6]) | (inputs[96]);
    assign layer0_outputs[5344] = (inputs[224]) & ~(inputs[210]);
    assign layer0_outputs[5345] = ~((inputs[235]) | (inputs[97]));
    assign layer0_outputs[5346] = ~((inputs[60]) | (inputs[46]));
    assign layer0_outputs[5347] = (inputs[161]) | (inputs[217]);
    assign layer0_outputs[5348] = (inputs[23]) & ~(inputs[59]);
    assign layer0_outputs[5349] = inputs[129];
    assign layer0_outputs[5350] = ~((inputs[94]) ^ (inputs[197]));
    assign layer0_outputs[5351] = (inputs[35]) ^ (inputs[131]);
    assign layer0_outputs[5352] = (inputs[18]) ^ (inputs[70]);
    assign layer0_outputs[5353] = (inputs[60]) & ~(inputs[238]);
    assign layer0_outputs[5354] = (inputs[245]) ^ (inputs[161]);
    assign layer0_outputs[5355] = ~(inputs[170]) | (inputs[69]);
    assign layer0_outputs[5356] = ~(inputs[194]);
    assign layer0_outputs[5357] = (inputs[19]) | (inputs[8]);
    assign layer0_outputs[5358] = ~((inputs[28]) | (inputs[177]));
    assign layer0_outputs[5359] = (inputs[243]) & ~(inputs[142]);
    assign layer0_outputs[5360] = ~(inputs[115]) | (inputs[109]);
    assign layer0_outputs[5361] = ~((inputs[225]) | (inputs[211]));
    assign layer0_outputs[5362] = ~((inputs[151]) | (inputs[207]));
    assign layer0_outputs[5363] = (inputs[1]) | (inputs[197]);
    assign layer0_outputs[5364] = ~((inputs[173]) | (inputs[53]));
    assign layer0_outputs[5365] = (inputs[231]) ^ (inputs[255]);
    assign layer0_outputs[5366] = ~(inputs[125]);
    assign layer0_outputs[5367] = (inputs[67]) & (inputs[153]);
    assign layer0_outputs[5368] = ~(inputs[160]);
    assign layer0_outputs[5369] = (inputs[144]) ^ (inputs[84]);
    assign layer0_outputs[5370] = inputs[234];
    assign layer0_outputs[5371] = (inputs[162]) & ~(inputs[251]);
    assign layer0_outputs[5372] = 1'b1;
    assign layer0_outputs[5373] = (inputs[116]) ^ (inputs[128]);
    assign layer0_outputs[5374] = ~(inputs[245]);
    assign layer0_outputs[5375] = (inputs[174]) & ~(inputs[117]);
    assign layer0_outputs[5376] = inputs[212];
    assign layer0_outputs[5377] = (inputs[217]) ^ (inputs[210]);
    assign layer0_outputs[5378] = (inputs[69]) | (inputs[62]);
    assign layer0_outputs[5379] = ~(inputs[214]) | (inputs[13]);
    assign layer0_outputs[5380] = ~(inputs[223]) | (inputs[195]);
    assign layer0_outputs[5381] = inputs[41];
    assign layer0_outputs[5382] = ~(inputs[69]) | (inputs[101]);
    assign layer0_outputs[5383] = ~((inputs[219]) & (inputs[114]));
    assign layer0_outputs[5384] = inputs[76];
    assign layer0_outputs[5385] = ~(inputs[93]);
    assign layer0_outputs[5386] = ~(inputs[166]);
    assign layer0_outputs[5387] = (inputs[200]) | (inputs[99]);
    assign layer0_outputs[5388] = 1'b0;
    assign layer0_outputs[5389] = ~((inputs[63]) ^ (inputs[90]));
    assign layer0_outputs[5390] = (inputs[226]) & ~(inputs[45]);
    assign layer0_outputs[5391] = ~((inputs[90]) | (inputs[136]));
    assign layer0_outputs[5392] = (inputs[204]) | (inputs[66]);
    assign layer0_outputs[5393] = ~((inputs[188]) | (inputs[228]));
    assign layer0_outputs[5394] = ~((inputs[96]) & (inputs[74]));
    assign layer0_outputs[5395] = ~(inputs[253]);
    assign layer0_outputs[5396] = ~(inputs[246]) | (inputs[119]);
    assign layer0_outputs[5397] = (inputs[65]) & ~(inputs[108]);
    assign layer0_outputs[5398] = (inputs[66]) & ~(inputs[79]);
    assign layer0_outputs[5399] = (inputs[179]) & ~(inputs[160]);
    assign layer0_outputs[5400] = (inputs[95]) ^ (inputs[19]);
    assign layer0_outputs[5401] = ~((inputs[50]) | (inputs[86]));
    assign layer0_outputs[5402] = (inputs[77]) & ~(inputs[254]);
    assign layer0_outputs[5403] = ~(inputs[225]);
    assign layer0_outputs[5404] = ~((inputs[80]) | (inputs[196]));
    assign layer0_outputs[5405] = ~(inputs[211]) | (inputs[8]);
    assign layer0_outputs[5406] = ~(inputs[251]) | (inputs[246]);
    assign layer0_outputs[5407] = ~((inputs[210]) & (inputs[199]));
    assign layer0_outputs[5408] = (inputs[97]) & (inputs[97]);
    assign layer0_outputs[5409] = ~((inputs[189]) | (inputs[7]));
    assign layer0_outputs[5410] = (inputs[112]) ^ (inputs[99]);
    assign layer0_outputs[5411] = 1'b1;
    assign layer0_outputs[5412] = (inputs[9]) & ~(inputs[191]);
    assign layer0_outputs[5413] = ~(inputs[234]);
    assign layer0_outputs[5414] = (inputs[144]) & ~(inputs[223]);
    assign layer0_outputs[5415] = ~((inputs[214]) & (inputs[148]));
    assign layer0_outputs[5416] = ~(inputs[17]) | (inputs[222]);
    assign layer0_outputs[5417] = ~(inputs[184]);
    assign layer0_outputs[5418] = inputs[151];
    assign layer0_outputs[5419] = ~(inputs[196]) | (inputs[113]);
    assign layer0_outputs[5420] = (inputs[105]) & ~(inputs[161]);
    assign layer0_outputs[5421] = (inputs[48]) ^ (inputs[17]);
    assign layer0_outputs[5422] = ~(inputs[13]);
    assign layer0_outputs[5423] = ~((inputs[72]) ^ (inputs[12]));
    assign layer0_outputs[5424] = ~(inputs[188]) | (inputs[244]);
    assign layer0_outputs[5425] = inputs[190];
    assign layer0_outputs[5426] = ~((inputs[118]) ^ (inputs[150]));
    assign layer0_outputs[5427] = ~((inputs[105]) & (inputs[179]));
    assign layer0_outputs[5428] = (inputs[202]) & ~(inputs[198]);
    assign layer0_outputs[5429] = ~((inputs[134]) | (inputs[134]));
    assign layer0_outputs[5430] = ~(inputs[195]) | (inputs[57]);
    assign layer0_outputs[5431] = (inputs[46]) & ~(inputs[191]);
    assign layer0_outputs[5432] = 1'b0;
    assign layer0_outputs[5433] = 1'b1;
    assign layer0_outputs[5434] = ~(inputs[75]);
    assign layer0_outputs[5435] = ~((inputs[164]) | (inputs[163]));
    assign layer0_outputs[5436] = inputs[69];
    assign layer0_outputs[5437] = (inputs[76]) & ~(inputs[121]);
    assign layer0_outputs[5438] = inputs[103];
    assign layer0_outputs[5439] = inputs[188];
    assign layer0_outputs[5440] = (inputs[158]) & (inputs[212]);
    assign layer0_outputs[5441] = (inputs[192]) | (inputs[6]);
    assign layer0_outputs[5442] = ~((inputs[163]) & (inputs[100]));
    assign layer0_outputs[5443] = ~((inputs[227]) ^ (inputs[248]));
    assign layer0_outputs[5444] = inputs[136];
    assign layer0_outputs[5445] = (inputs[246]) & (inputs[6]);
    assign layer0_outputs[5446] = ~((inputs[149]) & (inputs[141]));
    assign layer0_outputs[5447] = ~(inputs[42]) | (inputs[143]);
    assign layer0_outputs[5448] = inputs[73];
    assign layer0_outputs[5449] = (inputs[205]) & (inputs[154]);
    assign layer0_outputs[5450] = inputs[56];
    assign layer0_outputs[5451] = (inputs[72]) & ~(inputs[58]);
    assign layer0_outputs[5452] = 1'b1;
    assign layer0_outputs[5453] = ~((inputs[184]) ^ (inputs[246]));
    assign layer0_outputs[5454] = 1'b0;
    assign layer0_outputs[5455] = (inputs[198]) & ~(inputs[236]);
    assign layer0_outputs[5456] = ~(inputs[244]);
    assign layer0_outputs[5457] = ~(inputs[55]) | (inputs[112]);
    assign layer0_outputs[5458] = (inputs[76]) ^ (inputs[73]);
    assign layer0_outputs[5459] = ~(inputs[148]) | (inputs[247]);
    assign layer0_outputs[5460] = ~((inputs[107]) ^ (inputs[0]));
    assign layer0_outputs[5461] = (inputs[116]) ^ (inputs[145]);
    assign layer0_outputs[5462] = ~((inputs[149]) | (inputs[188]));
    assign layer0_outputs[5463] = ~(inputs[247]) | (inputs[223]);
    assign layer0_outputs[5464] = inputs[17];
    assign layer0_outputs[5465] = inputs[162];
    assign layer0_outputs[5466] = ~((inputs[106]) ^ (inputs[142]));
    assign layer0_outputs[5467] = (inputs[157]) & ~(inputs[239]);
    assign layer0_outputs[5468] = 1'b0;
    assign layer0_outputs[5469] = ~(inputs[125]);
    assign layer0_outputs[5470] = 1'b1;
    assign layer0_outputs[5471] = (inputs[149]) ^ (inputs[194]);
    assign layer0_outputs[5472] = (inputs[164]) ^ (inputs[250]);
    assign layer0_outputs[5473] = ~(inputs[222]);
    assign layer0_outputs[5474] = (inputs[199]) & ~(inputs[16]);
    assign layer0_outputs[5475] = (inputs[56]) ^ (inputs[13]);
    assign layer0_outputs[5476] = 1'b0;
    assign layer0_outputs[5477] = ~(inputs[97]);
    assign layer0_outputs[5478] = (inputs[211]) & ~(inputs[93]);
    assign layer0_outputs[5479] = (inputs[48]) & (inputs[94]);
    assign layer0_outputs[5480] = ~(inputs[73]);
    assign layer0_outputs[5481] = (inputs[49]) & (inputs[111]);
    assign layer0_outputs[5482] = ~((inputs[213]) | (inputs[14]));
    assign layer0_outputs[5483] = ~(inputs[61]);
    assign layer0_outputs[5484] = inputs[143];
    assign layer0_outputs[5485] = 1'b0;
    assign layer0_outputs[5486] = ~(inputs[152]) | (inputs[111]);
    assign layer0_outputs[5487] = 1'b0;
    assign layer0_outputs[5488] = ~(inputs[147]);
    assign layer0_outputs[5489] = ~(inputs[225]);
    assign layer0_outputs[5490] = ~(inputs[134]);
    assign layer0_outputs[5491] = ~(inputs[106]) | (inputs[83]);
    assign layer0_outputs[5492] = (inputs[156]) & ~(inputs[211]);
    assign layer0_outputs[5493] = ~(inputs[5]) | (inputs[11]);
    assign layer0_outputs[5494] = (inputs[246]) | (inputs[159]);
    assign layer0_outputs[5495] = ~((inputs[184]) & (inputs[186]));
    assign layer0_outputs[5496] = inputs[134];
    assign layer0_outputs[5497] = ~((inputs[14]) | (inputs[119]));
    assign layer0_outputs[5498] = inputs[214];
    assign layer0_outputs[5499] = inputs[145];
    assign layer0_outputs[5500] = ~(inputs[89]) | (inputs[238]);
    assign layer0_outputs[5501] = ~((inputs[134]) | (inputs[143]));
    assign layer0_outputs[5502] = (inputs[175]) ^ (inputs[35]);
    assign layer0_outputs[5503] = ~(inputs[182]) | (inputs[215]);
    assign layer0_outputs[5504] = (inputs[107]) ^ (inputs[35]);
    assign layer0_outputs[5505] = (inputs[253]) & ~(inputs[237]);
    assign layer0_outputs[5506] = 1'b1;
    assign layer0_outputs[5507] = inputs[119];
    assign layer0_outputs[5508] = ~(inputs[233]);
    assign layer0_outputs[5509] = (inputs[165]) & ~(inputs[144]);
    assign layer0_outputs[5510] = ~((inputs[24]) & (inputs[27]));
    assign layer0_outputs[5511] = (inputs[186]) | (inputs[117]);
    assign layer0_outputs[5512] = ~(inputs[43]) | (inputs[100]);
    assign layer0_outputs[5513] = (inputs[14]) & ~(inputs[42]);
    assign layer0_outputs[5514] = inputs[213];
    assign layer0_outputs[5515] = ~((inputs[139]) | (inputs[147]));
    assign layer0_outputs[5516] = (inputs[134]) | (inputs[204]);
    assign layer0_outputs[5517] = ~(inputs[46]) | (inputs[42]);
    assign layer0_outputs[5518] = inputs[118];
    assign layer0_outputs[5519] = (inputs[175]) | (inputs[186]);
    assign layer0_outputs[5520] = ~(inputs[213]) | (inputs[201]);
    assign layer0_outputs[5521] = inputs[162];
    assign layer0_outputs[5522] = ~(inputs[243]) | (inputs[161]);
    assign layer0_outputs[5523] = inputs[85];
    assign layer0_outputs[5524] = ~(inputs[185]);
    assign layer0_outputs[5525] = 1'b0;
    assign layer0_outputs[5526] = (inputs[226]) ^ (inputs[155]);
    assign layer0_outputs[5527] = (inputs[30]) & (inputs[34]);
    assign layer0_outputs[5528] = (inputs[92]) & (inputs[68]);
    assign layer0_outputs[5529] = (inputs[129]) | (inputs[189]);
    assign layer0_outputs[5530] = (inputs[89]) & ~(inputs[191]);
    assign layer0_outputs[5531] = (inputs[172]) | (inputs[112]);
    assign layer0_outputs[5532] = (inputs[48]) & ~(inputs[39]);
    assign layer0_outputs[5533] = ~((inputs[231]) ^ (inputs[226]));
    assign layer0_outputs[5534] = ~(inputs[23]) | (inputs[162]);
    assign layer0_outputs[5535] = (inputs[11]) & ~(inputs[157]);
    assign layer0_outputs[5536] = ~(inputs[140]) | (inputs[218]);
    assign layer0_outputs[5537] = inputs[85];
    assign layer0_outputs[5538] = ~((inputs[79]) & (inputs[192]));
    assign layer0_outputs[5539] = inputs[186];
    assign layer0_outputs[5540] = (inputs[154]) & ~(inputs[15]);
    assign layer0_outputs[5541] = inputs[29];
    assign layer0_outputs[5542] = ~((inputs[95]) ^ (inputs[60]));
    assign layer0_outputs[5543] = ~(inputs[199]) | (inputs[119]);
    assign layer0_outputs[5544] = inputs[214];
    assign layer0_outputs[5545] = 1'b1;
    assign layer0_outputs[5546] = (inputs[230]) & (inputs[104]);
    assign layer0_outputs[5547] = (inputs[33]) | (inputs[51]);
    assign layer0_outputs[5548] = inputs[77];
    assign layer0_outputs[5549] = ~(inputs[171]);
    assign layer0_outputs[5550] = ~((inputs[2]) | (inputs[21]));
    assign layer0_outputs[5551] = inputs[77];
    assign layer0_outputs[5552] = 1'b0;
    assign layer0_outputs[5553] = ~((inputs[246]) | (inputs[226]));
    assign layer0_outputs[5554] = ~(inputs[101]);
    assign layer0_outputs[5555] = ~(inputs[67]);
    assign layer0_outputs[5556] = ~(inputs[129]);
    assign layer0_outputs[5557] = (inputs[46]) ^ (inputs[32]);
    assign layer0_outputs[5558] = ~(inputs[80]);
    assign layer0_outputs[5559] = (inputs[45]) ^ (inputs[241]);
    assign layer0_outputs[5560] = ~((inputs[95]) | (inputs[185]));
    assign layer0_outputs[5561] = (inputs[229]) & ~(inputs[94]);
    assign layer0_outputs[5562] = (inputs[210]) | (inputs[238]);
    assign layer0_outputs[5563] = ~((inputs[202]) | (inputs[189]));
    assign layer0_outputs[5564] = inputs[228];
    assign layer0_outputs[5565] = ~(inputs[33]) | (inputs[31]);
    assign layer0_outputs[5566] = inputs[230];
    assign layer0_outputs[5567] = (inputs[120]) & ~(inputs[157]);
    assign layer0_outputs[5568] = ~(inputs[255]) | (inputs[227]);
    assign layer0_outputs[5569] = ~(inputs[49]);
    assign layer0_outputs[5570] = ~((inputs[149]) | (inputs[137]));
    assign layer0_outputs[5571] = (inputs[103]) | (inputs[68]);
    assign layer0_outputs[5572] = inputs[186];
    assign layer0_outputs[5573] = (inputs[31]) | (inputs[10]);
    assign layer0_outputs[5574] = (inputs[142]) ^ (inputs[118]);
    assign layer0_outputs[5575] = (inputs[219]) | (inputs[212]);
    assign layer0_outputs[5576] = ~(inputs[240]) | (inputs[28]);
    assign layer0_outputs[5577] = (inputs[139]) | (inputs[187]);
    assign layer0_outputs[5578] = inputs[136];
    assign layer0_outputs[5579] = inputs[96];
    assign layer0_outputs[5580] = inputs[7];
    assign layer0_outputs[5581] = (inputs[130]) & ~(inputs[213]);
    assign layer0_outputs[5582] = inputs[61];
    assign layer0_outputs[5583] = ~(inputs[28]) | (inputs[255]);
    assign layer0_outputs[5584] = ~((inputs[84]) & (inputs[83]));
    assign layer0_outputs[5585] = (inputs[250]) | (inputs[14]);
    assign layer0_outputs[5586] = (inputs[65]) & ~(inputs[244]);
    assign layer0_outputs[5587] = ~((inputs[20]) ^ (inputs[188]));
    assign layer0_outputs[5588] = ~(inputs[40]);
    assign layer0_outputs[5589] = inputs[27];
    assign layer0_outputs[5590] = (inputs[28]) & (inputs[85]);
    assign layer0_outputs[5591] = ~(inputs[78]);
    assign layer0_outputs[5592] = ~((inputs[216]) ^ (inputs[234]));
    assign layer0_outputs[5593] = (inputs[207]) & ~(inputs[178]);
    assign layer0_outputs[5594] = inputs[156];
    assign layer0_outputs[5595] = inputs[57];
    assign layer0_outputs[5596] = (inputs[25]) ^ (inputs[231]);
    assign layer0_outputs[5597] = ~(inputs[121]) | (inputs[144]);
    assign layer0_outputs[5598] = (inputs[61]) & ~(inputs[170]);
    assign layer0_outputs[5599] = (inputs[232]) | (inputs[113]);
    assign layer0_outputs[5600] = (inputs[194]) ^ (inputs[220]);
    assign layer0_outputs[5601] = ~(inputs[213]);
    assign layer0_outputs[5602] = (inputs[160]) | (inputs[245]);
    assign layer0_outputs[5603] = ~((inputs[132]) & (inputs[157]));
    assign layer0_outputs[5604] = ~((inputs[180]) ^ (inputs[160]));
    assign layer0_outputs[5605] = (inputs[134]) | (inputs[166]);
    assign layer0_outputs[5606] = (inputs[114]) & (inputs[25]);
    assign layer0_outputs[5607] = ~((inputs[213]) & (inputs[246]));
    assign layer0_outputs[5608] = ~(inputs[249]);
    assign layer0_outputs[5609] = ~((inputs[150]) | (inputs[22]));
    assign layer0_outputs[5610] = inputs[14];
    assign layer0_outputs[5611] = ~((inputs[11]) ^ (inputs[207]));
    assign layer0_outputs[5612] = inputs[10];
    assign layer0_outputs[5613] = inputs[97];
    assign layer0_outputs[5614] = ~((inputs[160]) | (inputs[32]));
    assign layer0_outputs[5615] = ~(inputs[190]);
    assign layer0_outputs[5616] = ~(inputs[34]) | (inputs[191]);
    assign layer0_outputs[5617] = ~(inputs[194]);
    assign layer0_outputs[5618] = (inputs[231]) & (inputs[253]);
    assign layer0_outputs[5619] = (inputs[19]) & ~(inputs[187]);
    assign layer0_outputs[5620] = inputs[162];
    assign layer0_outputs[5621] = ~(inputs[242]);
    assign layer0_outputs[5622] = ~((inputs[44]) | (inputs[63]));
    assign layer0_outputs[5623] = ~((inputs[255]) | (inputs[240]));
    assign layer0_outputs[5624] = ~((inputs[83]) | (inputs[221]));
    assign layer0_outputs[5625] = ~(inputs[40]);
    assign layer0_outputs[5626] = ~((inputs[130]) ^ (inputs[206]));
    assign layer0_outputs[5627] = inputs[235];
    assign layer0_outputs[5628] = ~(inputs[24]);
    assign layer0_outputs[5629] = (inputs[250]) & (inputs[182]);
    assign layer0_outputs[5630] = ~(inputs[27]) | (inputs[103]);
    assign layer0_outputs[5631] = ~((inputs[230]) | (inputs[65]));
    assign layer0_outputs[5632] = inputs[50];
    assign layer0_outputs[5633] = 1'b1;
    assign layer0_outputs[5634] = ~((inputs[197]) | (inputs[78]));
    assign layer0_outputs[5635] = ~((inputs[18]) & (inputs[235]));
    assign layer0_outputs[5636] = (inputs[113]) | (inputs[181]);
    assign layer0_outputs[5637] = ~(inputs[90]) | (inputs[224]);
    assign layer0_outputs[5638] = ~((inputs[145]) ^ (inputs[130]));
    assign layer0_outputs[5639] = inputs[195];
    assign layer0_outputs[5640] = inputs[19];
    assign layer0_outputs[5641] = ~(inputs[29]);
    assign layer0_outputs[5642] = (inputs[73]) & (inputs[5]);
    assign layer0_outputs[5643] = inputs[34];
    assign layer0_outputs[5644] = inputs[7];
    assign layer0_outputs[5645] = ~(inputs[62]) | (inputs[50]);
    assign layer0_outputs[5646] = ~(inputs[104]);
    assign layer0_outputs[5647] = ~(inputs[124]);
    assign layer0_outputs[5648] = (inputs[34]) ^ (inputs[212]);
    assign layer0_outputs[5649] = ~(inputs[167]) | (inputs[82]);
    assign layer0_outputs[5650] = ~(inputs[78]);
    assign layer0_outputs[5651] = 1'b0;
    assign layer0_outputs[5652] = ~(inputs[124]);
    assign layer0_outputs[5653] = ~(inputs[23]);
    assign layer0_outputs[5654] = ~(inputs[209]) | (inputs[107]);
    assign layer0_outputs[5655] = (inputs[150]) | (inputs[183]);
    assign layer0_outputs[5656] = ~(inputs[57]);
    assign layer0_outputs[5657] = ~(inputs[119]);
    assign layer0_outputs[5658] = (inputs[242]) | (inputs[75]);
    assign layer0_outputs[5659] = (inputs[156]) | (inputs[162]);
    assign layer0_outputs[5660] = (inputs[244]) & ~(inputs[121]);
    assign layer0_outputs[5661] = ~((inputs[103]) | (inputs[167]));
    assign layer0_outputs[5662] = 1'b1;
    assign layer0_outputs[5663] = (inputs[182]) | (inputs[160]);
    assign layer0_outputs[5664] = ~(inputs[235]);
    assign layer0_outputs[5665] = 1'b0;
    assign layer0_outputs[5666] = ~(inputs[60]) | (inputs[129]);
    assign layer0_outputs[5667] = ~((inputs[224]) | (inputs[25]));
    assign layer0_outputs[5668] = (inputs[128]) ^ (inputs[18]);
    assign layer0_outputs[5669] = (inputs[229]) & ~(inputs[137]);
    assign layer0_outputs[5670] = (inputs[238]) & (inputs[25]);
    assign layer0_outputs[5671] = (inputs[230]) | (inputs[247]);
    assign layer0_outputs[5672] = ~(inputs[28]) | (inputs[176]);
    assign layer0_outputs[5673] = inputs[99];
    assign layer0_outputs[5674] = ~((inputs[187]) ^ (inputs[158]));
    assign layer0_outputs[5675] = ~(inputs[243]);
    assign layer0_outputs[5676] = (inputs[13]) | (inputs[100]);
    assign layer0_outputs[5677] = ~((inputs[37]) & (inputs[19]));
    assign layer0_outputs[5678] = ~(inputs[232]);
    assign layer0_outputs[5679] = 1'b1;
    assign layer0_outputs[5680] = (inputs[94]) | (inputs[67]);
    assign layer0_outputs[5681] = ~((inputs[49]) ^ (inputs[16]));
    assign layer0_outputs[5682] = ~(inputs[25]);
    assign layer0_outputs[5683] = (inputs[145]) | (inputs[233]);
    assign layer0_outputs[5684] = ~(inputs[47]);
    assign layer0_outputs[5685] = (inputs[192]) & ~(inputs[94]);
    assign layer0_outputs[5686] = (inputs[104]) & ~(inputs[254]);
    assign layer0_outputs[5687] = inputs[193];
    assign layer0_outputs[5688] = ~(inputs[56]);
    assign layer0_outputs[5689] = ~((inputs[205]) | (inputs[53]));
    assign layer0_outputs[5690] = ~((inputs[123]) | (inputs[49]));
    assign layer0_outputs[5691] = (inputs[235]) ^ (inputs[238]);
    assign layer0_outputs[5692] = (inputs[86]) | (inputs[117]);
    assign layer0_outputs[5693] = (inputs[50]) & ~(inputs[248]);
    assign layer0_outputs[5694] = (inputs[62]) ^ (inputs[219]);
    assign layer0_outputs[5695] = (inputs[185]) & (inputs[157]);
    assign layer0_outputs[5696] = (inputs[90]) & ~(inputs[20]);
    assign layer0_outputs[5697] = (inputs[118]) & (inputs[140]);
    assign layer0_outputs[5698] = 1'b0;
    assign layer0_outputs[5699] = 1'b0;
    assign layer0_outputs[5700] = inputs[8];
    assign layer0_outputs[5701] = ~((inputs[88]) | (inputs[53]));
    assign layer0_outputs[5702] = ~(inputs[58]);
    assign layer0_outputs[5703] = ~((inputs[35]) ^ (inputs[17]));
    assign layer0_outputs[5704] = ~(inputs[198]);
    assign layer0_outputs[5705] = ~(inputs[131]);
    assign layer0_outputs[5706] = (inputs[50]) & (inputs[88]);
    assign layer0_outputs[5707] = inputs[241];
    assign layer0_outputs[5708] = inputs[231];
    assign layer0_outputs[5709] = ~(inputs[135]);
    assign layer0_outputs[5710] = (inputs[10]) & ~(inputs[87]);
    assign layer0_outputs[5711] = (inputs[101]) | (inputs[227]);
    assign layer0_outputs[5712] = (inputs[157]) & ~(inputs[254]);
    assign layer0_outputs[5713] = (inputs[239]) & (inputs[6]);
    assign layer0_outputs[5714] = ~(inputs[230]) | (inputs[4]);
    assign layer0_outputs[5715] = (inputs[125]) | (inputs[248]);
    assign layer0_outputs[5716] = ~(inputs[145]) | (inputs[255]);
    assign layer0_outputs[5717] = (inputs[56]) ^ (inputs[6]);
    assign layer0_outputs[5718] = inputs[224];
    assign layer0_outputs[5719] = (inputs[160]) & ~(inputs[28]);
    assign layer0_outputs[5720] = (inputs[99]) ^ (inputs[15]);
    assign layer0_outputs[5721] = ~(inputs[194]);
    assign layer0_outputs[5722] = ~(inputs[84]);
    assign layer0_outputs[5723] = ~((inputs[117]) ^ (inputs[103]));
    assign layer0_outputs[5724] = (inputs[37]) & ~(inputs[102]);
    assign layer0_outputs[5725] = ~(inputs[253]);
    assign layer0_outputs[5726] = (inputs[154]) & ~(inputs[201]);
    assign layer0_outputs[5727] = 1'b1;
    assign layer0_outputs[5728] = inputs[245];
    assign layer0_outputs[5729] = ~(inputs[90]);
    assign layer0_outputs[5730] = ~(inputs[143]);
    assign layer0_outputs[5731] = ~((inputs[90]) & (inputs[120]));
    assign layer0_outputs[5732] = (inputs[75]) & ~(inputs[190]);
    assign layer0_outputs[5733] = ~(inputs[127]);
    assign layer0_outputs[5734] = ~(inputs[187]);
    assign layer0_outputs[5735] = inputs[179];
    assign layer0_outputs[5736] = ~(inputs[176]) | (inputs[129]);
    assign layer0_outputs[5737] = ~((inputs[179]) ^ (inputs[220]));
    assign layer0_outputs[5738] = 1'b0;
    assign layer0_outputs[5739] = ~(inputs[38]);
    assign layer0_outputs[5740] = inputs[237];
    assign layer0_outputs[5741] = (inputs[236]) ^ (inputs[182]);
    assign layer0_outputs[5742] = ~(inputs[105]);
    assign layer0_outputs[5743] = ~((inputs[136]) & (inputs[44]));
    assign layer0_outputs[5744] = (inputs[126]) & ~(inputs[220]);
    assign layer0_outputs[5745] = (inputs[86]) & ~(inputs[242]);
    assign layer0_outputs[5746] = inputs[222];
    assign layer0_outputs[5747] = (inputs[117]) & ~(inputs[33]);
    assign layer0_outputs[5748] = ~(inputs[242]);
    assign layer0_outputs[5749] = inputs[232];
    assign layer0_outputs[5750] = inputs[118];
    assign layer0_outputs[5751] = (inputs[103]) & ~(inputs[251]);
    assign layer0_outputs[5752] = (inputs[44]) & ~(inputs[187]);
    assign layer0_outputs[5753] = ~((inputs[93]) | (inputs[76]));
    assign layer0_outputs[5754] = (inputs[165]) & ~(inputs[96]);
    assign layer0_outputs[5755] = ~((inputs[231]) ^ (inputs[159]));
    assign layer0_outputs[5756] = inputs[96];
    assign layer0_outputs[5757] = 1'b0;
    assign layer0_outputs[5758] = (inputs[87]) & ~(inputs[179]);
    assign layer0_outputs[5759] = (inputs[148]) | (inputs[48]);
    assign layer0_outputs[5760] = (inputs[214]) ^ (inputs[108]);
    assign layer0_outputs[5761] = (inputs[187]) | (inputs[176]);
    assign layer0_outputs[5762] = inputs[52];
    assign layer0_outputs[5763] = ~((inputs[252]) ^ (inputs[190]));
    assign layer0_outputs[5764] = ~(inputs[140]);
    assign layer0_outputs[5765] = inputs[232];
    assign layer0_outputs[5766] = (inputs[126]) & ~(inputs[14]);
    assign layer0_outputs[5767] = ~(inputs[118]);
    assign layer0_outputs[5768] = (inputs[107]) ^ (inputs[77]);
    assign layer0_outputs[5769] = (inputs[247]) & (inputs[149]);
    assign layer0_outputs[5770] = ~(inputs[21]) | (inputs[224]);
    assign layer0_outputs[5771] = ~(inputs[214]) | (inputs[37]);
    assign layer0_outputs[5772] = ~((inputs[223]) | (inputs[227]));
    assign layer0_outputs[5773] = (inputs[109]) & ~(inputs[9]);
    assign layer0_outputs[5774] = inputs[145];
    assign layer0_outputs[5775] = ~(inputs[75]) | (inputs[124]);
    assign layer0_outputs[5776] = ~(inputs[115]);
    assign layer0_outputs[5777] = (inputs[144]) ^ (inputs[174]);
    assign layer0_outputs[5778] = (inputs[128]) | (inputs[23]);
    assign layer0_outputs[5779] = 1'b1;
    assign layer0_outputs[5780] = ~((inputs[117]) ^ (inputs[149]));
    assign layer0_outputs[5781] = ~(inputs[95]);
    assign layer0_outputs[5782] = ~(inputs[193]) | (inputs[65]);
    assign layer0_outputs[5783] = (inputs[187]) ^ (inputs[131]);
    assign layer0_outputs[5784] = (inputs[242]) ^ (inputs[244]);
    assign layer0_outputs[5785] = ~((inputs[158]) | (inputs[110]));
    assign layer0_outputs[5786] = inputs[167];
    assign layer0_outputs[5787] = ~((inputs[87]) ^ (inputs[42]));
    assign layer0_outputs[5788] = ~(inputs[150]) | (inputs[22]);
    assign layer0_outputs[5789] = ~(inputs[125]);
    assign layer0_outputs[5790] = 1'b0;
    assign layer0_outputs[5791] = ~(inputs[236]);
    assign layer0_outputs[5792] = (inputs[103]) | (inputs[241]);
    assign layer0_outputs[5793] = (inputs[172]) | (inputs[4]);
    assign layer0_outputs[5794] = 1'b1;
    assign layer0_outputs[5795] = 1'b1;
    assign layer0_outputs[5796] = ~((inputs[195]) & (inputs[141]));
    assign layer0_outputs[5797] = ~(inputs[38]) | (inputs[179]);
    assign layer0_outputs[5798] = (inputs[0]) & ~(inputs[28]);
    assign layer0_outputs[5799] = (inputs[124]) & ~(inputs[197]);
    assign layer0_outputs[5800] = (inputs[206]) & ~(inputs[43]);
    assign layer0_outputs[5801] = ~(inputs[249]);
    assign layer0_outputs[5802] = (inputs[1]) | (inputs[210]);
    assign layer0_outputs[5803] = 1'b1;
    assign layer0_outputs[5804] = (inputs[43]) | (inputs[14]);
    assign layer0_outputs[5805] = ~(inputs[212]);
    assign layer0_outputs[5806] = 1'b0;
    assign layer0_outputs[5807] = ~(inputs[155]);
    assign layer0_outputs[5808] = inputs[105];
    assign layer0_outputs[5809] = (inputs[30]) ^ (inputs[86]);
    assign layer0_outputs[5810] = (inputs[93]) & (inputs[127]);
    assign layer0_outputs[5811] = inputs[182];
    assign layer0_outputs[5812] = inputs[164];
    assign layer0_outputs[5813] = ~(inputs[239]) | (inputs[200]);
    assign layer0_outputs[5814] = inputs[134];
    assign layer0_outputs[5815] = inputs[163];
    assign layer0_outputs[5816] = (inputs[190]) | (inputs[96]);
    assign layer0_outputs[5817] = ~((inputs[150]) | (inputs[66]));
    assign layer0_outputs[5818] = ~(inputs[254]) | (inputs[251]);
    assign layer0_outputs[5819] = ~(inputs[165]);
    assign layer0_outputs[5820] = (inputs[236]) ^ (inputs[173]);
    assign layer0_outputs[5821] = ~(inputs[117]);
    assign layer0_outputs[5822] = (inputs[119]) ^ (inputs[74]);
    assign layer0_outputs[5823] = ~(inputs[158]) | (inputs[28]);
    assign layer0_outputs[5824] = (inputs[157]) ^ (inputs[226]);
    assign layer0_outputs[5825] = (inputs[62]) & ~(inputs[14]);
    assign layer0_outputs[5826] = inputs[152];
    assign layer0_outputs[5827] = 1'b1;
    assign layer0_outputs[5828] = ~(inputs[245]) | (inputs[79]);
    assign layer0_outputs[5829] = (inputs[79]) | (inputs[125]);
    assign layer0_outputs[5830] = ~(inputs[118]);
    assign layer0_outputs[5831] = ~(inputs[58]) | (inputs[207]);
    assign layer0_outputs[5832] = ~(inputs[85]) | (inputs[240]);
    assign layer0_outputs[5833] = (inputs[6]) ^ (inputs[133]);
    assign layer0_outputs[5834] = ~((inputs[89]) | (inputs[11]));
    assign layer0_outputs[5835] = (inputs[190]) & ~(inputs[254]);
    assign layer0_outputs[5836] = ~(inputs[27]);
    assign layer0_outputs[5837] = 1'b0;
    assign layer0_outputs[5838] = (inputs[33]) & ~(inputs[184]);
    assign layer0_outputs[5839] = ~(inputs[169]);
    assign layer0_outputs[5840] = (inputs[56]) & ~(inputs[35]);
    assign layer0_outputs[5841] = ~((inputs[0]) | (inputs[68]));
    assign layer0_outputs[5842] = inputs[48];
    assign layer0_outputs[5843] = ~(inputs[220]);
    assign layer0_outputs[5844] = (inputs[73]) & (inputs[196]);
    assign layer0_outputs[5845] = ~((inputs[144]) | (inputs[88]));
    assign layer0_outputs[5846] = ~(inputs[234]);
    assign layer0_outputs[5847] = (inputs[28]) & ~(inputs[243]);
    assign layer0_outputs[5848] = ~(inputs[228]);
    assign layer0_outputs[5849] = ~((inputs[70]) | (inputs[97]));
    assign layer0_outputs[5850] = ~(inputs[119]);
    assign layer0_outputs[5851] = ~(inputs[62]);
    assign layer0_outputs[5852] = (inputs[232]) & ~(inputs[36]);
    assign layer0_outputs[5853] = ~((inputs[119]) & (inputs[71]));
    assign layer0_outputs[5854] = inputs[77];
    assign layer0_outputs[5855] = inputs[164];
    assign layer0_outputs[5856] = inputs[167];
    assign layer0_outputs[5857] = inputs[247];
    assign layer0_outputs[5858] = inputs[63];
    assign layer0_outputs[5859] = (inputs[98]) ^ (inputs[235]);
    assign layer0_outputs[5860] = ~(inputs[120]) | (inputs[149]);
    assign layer0_outputs[5861] = ~(inputs[114]) | (inputs[134]);
    assign layer0_outputs[5862] = ~((inputs[19]) ^ (inputs[38]));
    assign layer0_outputs[5863] = ~(inputs[44]) | (inputs[117]);
    assign layer0_outputs[5864] = (inputs[36]) & ~(inputs[231]);
    assign layer0_outputs[5865] = inputs[55];
    assign layer0_outputs[5866] = ~(inputs[79]) | (inputs[15]);
    assign layer0_outputs[5867] = ~(inputs[178]);
    assign layer0_outputs[5868] = (inputs[188]) | (inputs[247]);
    assign layer0_outputs[5869] = inputs[159];
    assign layer0_outputs[5870] = ~(inputs[54]) | (inputs[92]);
    assign layer0_outputs[5871] = inputs[237];
    assign layer0_outputs[5872] = ~(inputs[249]) | (inputs[231]);
    assign layer0_outputs[5873] = ~(inputs[171]) | (inputs[167]);
    assign layer0_outputs[5874] = inputs[123];
    assign layer0_outputs[5875] = (inputs[192]) & ~(inputs[208]);
    assign layer0_outputs[5876] = 1'b1;
    assign layer0_outputs[5877] = (inputs[253]) ^ (inputs[179]);
    assign layer0_outputs[5878] = ~(inputs[210]);
    assign layer0_outputs[5879] = (inputs[181]) | (inputs[180]);
    assign layer0_outputs[5880] = ~((inputs[199]) | (inputs[3]));
    assign layer0_outputs[5881] = (inputs[7]) & ~(inputs[30]);
    assign layer0_outputs[5882] = ~((inputs[220]) | (inputs[180]));
    assign layer0_outputs[5883] = 1'b0;
    assign layer0_outputs[5884] = ~(inputs[78]) | (inputs[234]);
    assign layer0_outputs[5885] = ~(inputs[0]) | (inputs[237]);
    assign layer0_outputs[5886] = ~(inputs[104]) | (inputs[111]);
    assign layer0_outputs[5887] = (inputs[113]) | (inputs[240]);
    assign layer0_outputs[5888] = inputs[82];
    assign layer0_outputs[5889] = ~(inputs[120]);
    assign layer0_outputs[5890] = ~(inputs[85]);
    assign layer0_outputs[5891] = ~((inputs[232]) | (inputs[234]));
    assign layer0_outputs[5892] = inputs[35];
    assign layer0_outputs[5893] = inputs[54];
    assign layer0_outputs[5894] = inputs[180];
    assign layer0_outputs[5895] = (inputs[120]) ^ (inputs[213]);
    assign layer0_outputs[5896] = ~((inputs[101]) | (inputs[86]));
    assign layer0_outputs[5897] = inputs[171];
    assign layer0_outputs[5898] = (inputs[168]) & ~(inputs[53]);
    assign layer0_outputs[5899] = ~((inputs[177]) | (inputs[116]));
    assign layer0_outputs[5900] = inputs[101];
    assign layer0_outputs[5901] = inputs[238];
    assign layer0_outputs[5902] = (inputs[98]) | (inputs[223]);
    assign layer0_outputs[5903] = ~(inputs[129]);
    assign layer0_outputs[5904] = ~((inputs[86]) ^ (inputs[149]));
    assign layer0_outputs[5905] = ~((inputs[107]) ^ (inputs[144]));
    assign layer0_outputs[5906] = ~(inputs[7]) | (inputs[249]);
    assign layer0_outputs[5907] = inputs[217];
    assign layer0_outputs[5908] = ~((inputs[163]) ^ (inputs[174]));
    assign layer0_outputs[5909] = ~((inputs[236]) ^ (inputs[255]));
    assign layer0_outputs[5910] = 1'b1;
    assign layer0_outputs[5911] = inputs[162];
    assign layer0_outputs[5912] = (inputs[124]) | (inputs[234]);
    assign layer0_outputs[5913] = inputs[2];
    assign layer0_outputs[5914] = ~((inputs[86]) ^ (inputs[55]));
    assign layer0_outputs[5915] = 1'b0;
    assign layer0_outputs[5916] = ~(inputs[246]);
    assign layer0_outputs[5917] = (inputs[140]) | (inputs[174]);
    assign layer0_outputs[5918] = inputs[80];
    assign layer0_outputs[5919] = inputs[148];
    assign layer0_outputs[5920] = inputs[45];
    assign layer0_outputs[5921] = ~((inputs[35]) & (inputs[20]));
    assign layer0_outputs[5922] = (inputs[201]) & (inputs[202]);
    assign layer0_outputs[5923] = (inputs[139]) | (inputs[77]);
    assign layer0_outputs[5924] = ~(inputs[10]) | (inputs[15]);
    assign layer0_outputs[5925] = ~((inputs[235]) | (inputs[2]));
    assign layer0_outputs[5926] = (inputs[237]) ^ (inputs[179]);
    assign layer0_outputs[5927] = ~(inputs[165]);
    assign layer0_outputs[5928] = (inputs[117]) & ~(inputs[3]);
    assign layer0_outputs[5929] = 1'b1;
    assign layer0_outputs[5930] = ~((inputs[60]) | (inputs[176]));
    assign layer0_outputs[5931] = (inputs[178]) & ~(inputs[128]);
    assign layer0_outputs[5932] = (inputs[121]) & ~(inputs[33]);
    assign layer0_outputs[5933] = inputs[117];
    assign layer0_outputs[5934] = ~(inputs[228]) | (inputs[0]);
    assign layer0_outputs[5935] = (inputs[204]) | (inputs[132]);
    assign layer0_outputs[5936] = inputs[82];
    assign layer0_outputs[5937] = (inputs[69]) | (inputs[15]);
    assign layer0_outputs[5938] = ~((inputs[15]) ^ (inputs[168]));
    assign layer0_outputs[5939] = ~(inputs[60]);
    assign layer0_outputs[5940] = inputs[98];
    assign layer0_outputs[5941] = inputs[197];
    assign layer0_outputs[5942] = ~(inputs[184]);
    assign layer0_outputs[5943] = ~(inputs[181]);
    assign layer0_outputs[5944] = inputs[203];
    assign layer0_outputs[5945] = inputs[158];
    assign layer0_outputs[5946] = (inputs[14]) | (inputs[183]);
    assign layer0_outputs[5947] = ~(inputs[92]);
    assign layer0_outputs[5948] = ~((inputs[246]) | (inputs[66]));
    assign layer0_outputs[5949] = ~(inputs[211]) | (inputs[166]);
    assign layer0_outputs[5950] = ~((inputs[84]) ^ (inputs[113]));
    assign layer0_outputs[5951] = ~(inputs[39]);
    assign layer0_outputs[5952] = ~(inputs[201]) | (inputs[47]);
    assign layer0_outputs[5953] = ~((inputs[56]) & (inputs[206]));
    assign layer0_outputs[5954] = (inputs[177]) | (inputs[162]);
    assign layer0_outputs[5955] = inputs[228];
    assign layer0_outputs[5956] = ~(inputs[94]);
    assign layer0_outputs[5957] = inputs[160];
    assign layer0_outputs[5958] = inputs[135];
    assign layer0_outputs[5959] = ~((inputs[80]) ^ (inputs[230]));
    assign layer0_outputs[5960] = ~(inputs[120]) | (inputs[65]);
    assign layer0_outputs[5961] = (inputs[91]) & (inputs[40]);
    assign layer0_outputs[5962] = ~(inputs[121]) | (inputs[56]);
    assign layer0_outputs[5963] = ~((inputs[159]) | (inputs[127]));
    assign layer0_outputs[5964] = ~((inputs[236]) ^ (inputs[12]));
    assign layer0_outputs[5965] = (inputs[224]) ^ (inputs[251]);
    assign layer0_outputs[5966] = (inputs[42]) & ~(inputs[203]);
    assign layer0_outputs[5967] = inputs[124];
    assign layer0_outputs[5968] = ~((inputs[177]) ^ (inputs[197]));
    assign layer0_outputs[5969] = inputs[75];
    assign layer0_outputs[5970] = ~((inputs[168]) ^ (inputs[180]));
    assign layer0_outputs[5971] = (inputs[164]) & ~(inputs[23]);
    assign layer0_outputs[5972] = ~(inputs[129]);
    assign layer0_outputs[5973] = inputs[125];
    assign layer0_outputs[5974] = ~(inputs[23]);
    assign layer0_outputs[5975] = ~((inputs[116]) | (inputs[89]));
    assign layer0_outputs[5976] = ~(inputs[0]) | (inputs[190]);
    assign layer0_outputs[5977] = (inputs[115]) ^ (inputs[50]);
    assign layer0_outputs[5978] = (inputs[61]) | (inputs[233]);
    assign layer0_outputs[5979] = (inputs[124]) | (inputs[44]);
    assign layer0_outputs[5980] = (inputs[51]) | (inputs[69]);
    assign layer0_outputs[5981] = ~((inputs[37]) | (inputs[123]));
    assign layer0_outputs[5982] = (inputs[3]) ^ (inputs[134]);
    assign layer0_outputs[5983] = (inputs[181]) ^ (inputs[95]);
    assign layer0_outputs[5984] = (inputs[103]) & (inputs[135]);
    assign layer0_outputs[5985] = inputs[212];
    assign layer0_outputs[5986] = (inputs[192]) | (inputs[202]);
    assign layer0_outputs[5987] = inputs[239];
    assign layer0_outputs[5988] = inputs[139];
    assign layer0_outputs[5989] = ~(inputs[232]);
    assign layer0_outputs[5990] = ~((inputs[234]) | (inputs[61]));
    assign layer0_outputs[5991] = ~((inputs[18]) | (inputs[197]));
    assign layer0_outputs[5992] = (inputs[122]) | (inputs[110]);
    assign layer0_outputs[5993] = (inputs[87]) & ~(inputs[215]);
    assign layer0_outputs[5994] = ~(inputs[240]);
    assign layer0_outputs[5995] = (inputs[196]) & ~(inputs[222]);
    assign layer0_outputs[5996] = ~(inputs[199]) | (inputs[152]);
    assign layer0_outputs[5997] = ~((inputs[38]) | (inputs[55]));
    assign layer0_outputs[5998] = (inputs[32]) | (inputs[125]);
    assign layer0_outputs[5999] = ~(inputs[89]) | (inputs[121]);
    assign layer0_outputs[6000] = inputs[233];
    assign layer0_outputs[6001] = ~(inputs[183]);
    assign layer0_outputs[6002] = ~((inputs[159]) | (inputs[113]));
    assign layer0_outputs[6003] = 1'b0;
    assign layer0_outputs[6004] = ~((inputs[85]) ^ (inputs[19]));
    assign layer0_outputs[6005] = inputs[70];
    assign layer0_outputs[6006] = inputs[120];
    assign layer0_outputs[6007] = (inputs[189]) | (inputs[160]);
    assign layer0_outputs[6008] = ~(inputs[87]);
    assign layer0_outputs[6009] = ~(inputs[215]);
    assign layer0_outputs[6010] = ~((inputs[239]) ^ (inputs[137]));
    assign layer0_outputs[6011] = (inputs[128]) & ~(inputs[109]);
    assign layer0_outputs[6012] = ~(inputs[232]) | (inputs[52]);
    assign layer0_outputs[6013] = inputs[238];
    assign layer0_outputs[6014] = (inputs[18]) | (inputs[244]);
    assign layer0_outputs[6015] = ~(inputs[178]) | (inputs[62]);
    assign layer0_outputs[6016] = ~((inputs[125]) | (inputs[180]));
    assign layer0_outputs[6017] = ~((inputs[158]) & (inputs[60]));
    assign layer0_outputs[6018] = ~((inputs[246]) | (inputs[130]));
    assign layer0_outputs[6019] = (inputs[164]) ^ (inputs[233]);
    assign layer0_outputs[6020] = ~(inputs[84]);
    assign layer0_outputs[6021] = ~(inputs[155]) | (inputs[250]);
    assign layer0_outputs[6022] = ~(inputs[111]) | (inputs[46]);
    assign layer0_outputs[6023] = (inputs[79]) | (inputs[187]);
    assign layer0_outputs[6024] = inputs[197];
    assign layer0_outputs[6025] = ~((inputs[165]) | (inputs[48]));
    assign layer0_outputs[6026] = (inputs[206]) & ~(inputs[201]);
    assign layer0_outputs[6027] = ~(inputs[148]);
    assign layer0_outputs[6028] = ~(inputs[86]) | (inputs[33]);
    assign layer0_outputs[6029] = (inputs[197]) | (inputs[221]);
    assign layer0_outputs[6030] = (inputs[143]) & ~(inputs[153]);
    assign layer0_outputs[6031] = inputs[131];
    assign layer0_outputs[6032] = ~(inputs[93]);
    assign layer0_outputs[6033] = ~(inputs[206]) | (inputs[116]);
    assign layer0_outputs[6034] = inputs[114];
    assign layer0_outputs[6035] = inputs[56];
    assign layer0_outputs[6036] = inputs[65];
    assign layer0_outputs[6037] = inputs[94];
    assign layer0_outputs[6038] = inputs[251];
    assign layer0_outputs[6039] = ~((inputs[62]) | (inputs[0]));
    assign layer0_outputs[6040] = ~((inputs[108]) ^ (inputs[210]));
    assign layer0_outputs[6041] = (inputs[167]) ^ (inputs[43]);
    assign layer0_outputs[6042] = ~((inputs[168]) ^ (inputs[209]));
    assign layer0_outputs[6043] = (inputs[243]) & ~(inputs[145]);
    assign layer0_outputs[6044] = ~((inputs[180]) | (inputs[31]));
    assign layer0_outputs[6045] = ~(inputs[80]);
    assign layer0_outputs[6046] = ~((inputs[153]) ^ (inputs[107]));
    assign layer0_outputs[6047] = ~(inputs[195]) | (inputs[94]);
    assign layer0_outputs[6048] = ~(inputs[4]);
    assign layer0_outputs[6049] = (inputs[125]) | (inputs[212]);
    assign layer0_outputs[6050] = ~((inputs[196]) ^ (inputs[145]));
    assign layer0_outputs[6051] = ~(inputs[47]);
    assign layer0_outputs[6052] = (inputs[6]) ^ (inputs[176]);
    assign layer0_outputs[6053] = ~((inputs[2]) ^ (inputs[224]));
    assign layer0_outputs[6054] = ~((inputs[166]) ^ (inputs[202]));
    assign layer0_outputs[6055] = ~(inputs[89]) | (inputs[203]);
    assign layer0_outputs[6056] = ~(inputs[96]);
    assign layer0_outputs[6057] = (inputs[226]) | (inputs[56]);
    assign layer0_outputs[6058] = inputs[136];
    assign layer0_outputs[6059] = ~(inputs[57]) | (inputs[151]);
    assign layer0_outputs[6060] = (inputs[200]) & ~(inputs[35]);
    assign layer0_outputs[6061] = inputs[39];
    assign layer0_outputs[6062] = 1'b0;
    assign layer0_outputs[6063] = inputs[253];
    assign layer0_outputs[6064] = ~(inputs[231]);
    assign layer0_outputs[6065] = ~(inputs[28]);
    assign layer0_outputs[6066] = (inputs[96]) | (inputs[98]);
    assign layer0_outputs[6067] = (inputs[179]) & ~(inputs[125]);
    assign layer0_outputs[6068] = ~((inputs[33]) ^ (inputs[67]));
    assign layer0_outputs[6069] = ~((inputs[169]) | (inputs[161]));
    assign layer0_outputs[6070] = ~(inputs[79]) | (inputs[1]);
    assign layer0_outputs[6071] = (inputs[240]) & (inputs[51]);
    assign layer0_outputs[6072] = ~(inputs[133]);
    assign layer0_outputs[6073] = ~((inputs[58]) ^ (inputs[23]));
    assign layer0_outputs[6074] = (inputs[131]) & ~(inputs[85]);
    assign layer0_outputs[6075] = inputs[88];
    assign layer0_outputs[6076] = ~((inputs[143]) | (inputs[196]));
    assign layer0_outputs[6077] = (inputs[187]) ^ (inputs[239]);
    assign layer0_outputs[6078] = ~((inputs[135]) ^ (inputs[72]));
    assign layer0_outputs[6079] = ~(inputs[167]);
    assign layer0_outputs[6080] = ~(inputs[143]);
    assign layer0_outputs[6081] = inputs[57];
    assign layer0_outputs[6082] = inputs[98];
    assign layer0_outputs[6083] = (inputs[8]) | (inputs[205]);
    assign layer0_outputs[6084] = 1'b0;
    assign layer0_outputs[6085] = ~(inputs[167]);
    assign layer0_outputs[6086] = (inputs[220]) ^ (inputs[128]);
    assign layer0_outputs[6087] = inputs[167];
    assign layer0_outputs[6088] = ~(inputs[117]) | (inputs[9]);
    assign layer0_outputs[6089] = ~(inputs[198]);
    assign layer0_outputs[6090] = 1'b0;
    assign layer0_outputs[6091] = inputs[98];
    assign layer0_outputs[6092] = (inputs[8]) & (inputs[90]);
    assign layer0_outputs[6093] = ~((inputs[89]) ^ (inputs[8]));
    assign layer0_outputs[6094] = ~((inputs[60]) | (inputs[125]));
    assign layer0_outputs[6095] = (inputs[165]) & ~(inputs[200]);
    assign layer0_outputs[6096] = (inputs[107]) & ~(inputs[234]);
    assign layer0_outputs[6097] = ~(inputs[42]) | (inputs[230]);
    assign layer0_outputs[6098] = ~(inputs[100]);
    assign layer0_outputs[6099] = (inputs[57]) | (inputs[134]);
    assign layer0_outputs[6100] = inputs[100];
    assign layer0_outputs[6101] = (inputs[53]) | (inputs[86]);
    assign layer0_outputs[6102] = ~(inputs[204]) | (inputs[49]);
    assign layer0_outputs[6103] = ~(inputs[93]) | (inputs[217]);
    assign layer0_outputs[6104] = ~((inputs[89]) ^ (inputs[42]));
    assign layer0_outputs[6105] = ~(inputs[119]) | (inputs[190]);
    assign layer0_outputs[6106] = inputs[74];
    assign layer0_outputs[6107] = (inputs[90]) & (inputs[76]);
    assign layer0_outputs[6108] = ~(inputs[118]);
    assign layer0_outputs[6109] = (inputs[43]) & ~(inputs[175]);
    assign layer0_outputs[6110] = (inputs[237]) | (inputs[102]);
    assign layer0_outputs[6111] = ~(inputs[90]);
    assign layer0_outputs[6112] = (inputs[236]) | (inputs[126]);
    assign layer0_outputs[6113] = (inputs[178]) | (inputs[48]);
    assign layer0_outputs[6114] = ~((inputs[153]) | (inputs[185]));
    assign layer0_outputs[6115] = (inputs[231]) ^ (inputs[197]);
    assign layer0_outputs[6116] = ~(inputs[233]) | (inputs[208]);
    assign layer0_outputs[6117] = ~((inputs[99]) | (inputs[100]));
    assign layer0_outputs[6118] = ~((inputs[208]) | (inputs[188]));
    assign layer0_outputs[6119] = ~(inputs[155]);
    assign layer0_outputs[6120] = inputs[46];
    assign layer0_outputs[6121] = inputs[194];
    assign layer0_outputs[6122] = ~(inputs[107]);
    assign layer0_outputs[6123] = ~((inputs[140]) ^ (inputs[112]));
    assign layer0_outputs[6124] = inputs[137];
    assign layer0_outputs[6125] = (inputs[46]) | (inputs[14]);
    assign layer0_outputs[6126] = ~((inputs[152]) & (inputs[101]));
    assign layer0_outputs[6127] = ~(inputs[98]);
    assign layer0_outputs[6128] = (inputs[90]) ^ (inputs[95]);
    assign layer0_outputs[6129] = (inputs[88]) & ~(inputs[187]);
    assign layer0_outputs[6130] = inputs[250];
    assign layer0_outputs[6131] = inputs[49];
    assign layer0_outputs[6132] = (inputs[30]) ^ (inputs[157]);
    assign layer0_outputs[6133] = ~((inputs[24]) ^ (inputs[206]));
    assign layer0_outputs[6134] = inputs[184];
    assign layer0_outputs[6135] = ~(inputs[69]) | (inputs[123]);
    assign layer0_outputs[6136] = inputs[32];
    assign layer0_outputs[6137] = (inputs[95]) ^ (inputs[92]);
    assign layer0_outputs[6138] = ~(inputs[126]);
    assign layer0_outputs[6139] = ~(inputs[191]);
    assign layer0_outputs[6140] = ~(inputs[57]);
    assign layer0_outputs[6141] = ~((inputs[214]) & (inputs[126]));
    assign layer0_outputs[6142] = (inputs[142]) | (inputs[137]);
    assign layer0_outputs[6143] = ~(inputs[91]);
    assign layer0_outputs[6144] = ~((inputs[209]) | (inputs[46]));
    assign layer0_outputs[6145] = (inputs[232]) ^ (inputs[248]);
    assign layer0_outputs[6146] = (inputs[205]) ^ (inputs[87]);
    assign layer0_outputs[6147] = inputs[206];
    assign layer0_outputs[6148] = ~((inputs[198]) & (inputs[19]));
    assign layer0_outputs[6149] = ~(inputs[220]) | (inputs[128]);
    assign layer0_outputs[6150] = ~((inputs[124]) ^ (inputs[225]));
    assign layer0_outputs[6151] = ~(inputs[31]);
    assign layer0_outputs[6152] = inputs[23];
    assign layer0_outputs[6153] = (inputs[163]) | (inputs[93]);
    assign layer0_outputs[6154] = ~(inputs[169]);
    assign layer0_outputs[6155] = ~(inputs[238]) | (inputs[31]);
    assign layer0_outputs[6156] = ~(inputs[233]) | (inputs[139]);
    assign layer0_outputs[6157] = (inputs[96]) | (inputs[145]);
    assign layer0_outputs[6158] = inputs[247];
    assign layer0_outputs[6159] = ~((inputs[150]) | (inputs[183]));
    assign layer0_outputs[6160] = ~(inputs[142]);
    assign layer0_outputs[6161] = (inputs[182]) ^ (inputs[61]);
    assign layer0_outputs[6162] = ~((inputs[214]) & (inputs[16]));
    assign layer0_outputs[6163] = ~(inputs[4]) | (inputs[94]);
    assign layer0_outputs[6164] = ~((inputs[129]) ^ (inputs[132]));
    assign layer0_outputs[6165] = ~(inputs[23]) | (inputs[246]);
    assign layer0_outputs[6166] = ~(inputs[59]) | (inputs[254]);
    assign layer0_outputs[6167] = (inputs[123]) & (inputs[63]);
    assign layer0_outputs[6168] = inputs[158];
    assign layer0_outputs[6169] = (inputs[222]) | (inputs[6]);
    assign layer0_outputs[6170] = ~((inputs[126]) | (inputs[60]));
    assign layer0_outputs[6171] = inputs[166];
    assign layer0_outputs[6172] = (inputs[65]) | (inputs[139]);
    assign layer0_outputs[6173] = (inputs[35]) ^ (inputs[112]);
    assign layer0_outputs[6174] = (inputs[54]) | (inputs[209]);
    assign layer0_outputs[6175] = ~(inputs[116]);
    assign layer0_outputs[6176] = (inputs[255]) ^ (inputs[121]);
    assign layer0_outputs[6177] = ~(inputs[204]);
    assign layer0_outputs[6178] = 1'b1;
    assign layer0_outputs[6179] = ~((inputs[138]) & (inputs[134]));
    assign layer0_outputs[6180] = inputs[184];
    assign layer0_outputs[6181] = ~((inputs[128]) | (inputs[83]));
    assign layer0_outputs[6182] = inputs[6];
    assign layer0_outputs[6183] = inputs[185];
    assign layer0_outputs[6184] = 1'b0;
    assign layer0_outputs[6185] = inputs[86];
    assign layer0_outputs[6186] = (inputs[150]) | (inputs[167]);
    assign layer0_outputs[6187] = ~((inputs[20]) & (inputs[10]));
    assign layer0_outputs[6188] = inputs[134];
    assign layer0_outputs[6189] = ~(inputs[192]) | (inputs[180]);
    assign layer0_outputs[6190] = (inputs[100]) & ~(inputs[93]);
    assign layer0_outputs[6191] = (inputs[112]) & ~(inputs[127]);
    assign layer0_outputs[6192] = inputs[128];
    assign layer0_outputs[6193] = ~(inputs[14]);
    assign layer0_outputs[6194] = 1'b0;
    assign layer0_outputs[6195] = ~((inputs[66]) | (inputs[38]));
    assign layer0_outputs[6196] = ~((inputs[74]) ^ (inputs[223]));
    assign layer0_outputs[6197] = ~((inputs[210]) | (inputs[36]));
    assign layer0_outputs[6198] = ~((inputs[244]) & (inputs[199]));
    assign layer0_outputs[6199] = ~((inputs[192]) & (inputs[189]));
    assign layer0_outputs[6200] = (inputs[137]) & ~(inputs[21]);
    assign layer0_outputs[6201] = inputs[231];
    assign layer0_outputs[6202] = (inputs[55]) | (inputs[207]);
    assign layer0_outputs[6203] = ~((inputs[125]) | (inputs[141]));
    assign layer0_outputs[6204] = inputs[65];
    assign layer0_outputs[6205] = ~(inputs[70]) | (inputs[239]);
    assign layer0_outputs[6206] = inputs[200];
    assign layer0_outputs[6207] = ~((inputs[131]) | (inputs[71]));
    assign layer0_outputs[6208] = inputs[88];
    assign layer0_outputs[6209] = inputs[83];
    assign layer0_outputs[6210] = ~(inputs[45]);
    assign layer0_outputs[6211] = ~((inputs[231]) | (inputs[230]));
    assign layer0_outputs[6212] = ~((inputs[66]) & (inputs[126]));
    assign layer0_outputs[6213] = (inputs[19]) ^ (inputs[238]);
    assign layer0_outputs[6214] = ~(inputs[95]) | (inputs[34]);
    assign layer0_outputs[6215] = 1'b0;
    assign layer0_outputs[6216] = (inputs[135]) & ~(inputs[67]);
    assign layer0_outputs[6217] = (inputs[106]) | (inputs[13]);
    assign layer0_outputs[6218] = (inputs[202]) & ~(inputs[18]);
    assign layer0_outputs[6219] = ~(inputs[181]);
    assign layer0_outputs[6220] = ~((inputs[208]) & (inputs[201]));
    assign layer0_outputs[6221] = ~((inputs[76]) & (inputs[92]));
    assign layer0_outputs[6222] = (inputs[115]) ^ (inputs[30]);
    assign layer0_outputs[6223] = (inputs[30]) | (inputs[141]);
    assign layer0_outputs[6224] = ~(inputs[83]);
    assign layer0_outputs[6225] = (inputs[30]) | (inputs[19]);
    assign layer0_outputs[6226] = ~(inputs[182]) | (inputs[50]);
    assign layer0_outputs[6227] = (inputs[37]) | (inputs[9]);
    assign layer0_outputs[6228] = ~(inputs[221]);
    assign layer0_outputs[6229] = ~(inputs[157]) | (inputs[212]);
    assign layer0_outputs[6230] = (inputs[72]) & ~(inputs[154]);
    assign layer0_outputs[6231] = (inputs[222]) & ~(inputs[66]);
    assign layer0_outputs[6232] = ~((inputs[167]) | (inputs[65]));
    assign layer0_outputs[6233] = ~(inputs[32]);
    assign layer0_outputs[6234] = (inputs[22]) & ~(inputs[121]);
    assign layer0_outputs[6235] = ~((inputs[23]) & (inputs[0]));
    assign layer0_outputs[6236] = ~((inputs[224]) | (inputs[108]));
    assign layer0_outputs[6237] = ~(inputs[227]);
    assign layer0_outputs[6238] = inputs[88];
    assign layer0_outputs[6239] = ~((inputs[230]) ^ (inputs[207]));
    assign layer0_outputs[6240] = ~(inputs[133]) | (inputs[172]);
    assign layer0_outputs[6241] = (inputs[190]) & ~(inputs[233]);
    assign layer0_outputs[6242] = ~((inputs[64]) | (inputs[149]));
    assign layer0_outputs[6243] = ~((inputs[124]) ^ (inputs[205]));
    assign layer0_outputs[6244] = ~((inputs[24]) | (inputs[28]));
    assign layer0_outputs[6245] = ~(inputs[253]);
    assign layer0_outputs[6246] = 1'b1;
    assign layer0_outputs[6247] = (inputs[18]) | (inputs[247]);
    assign layer0_outputs[6248] = ~(inputs[210]) | (inputs[113]);
    assign layer0_outputs[6249] = inputs[166];
    assign layer0_outputs[6250] = inputs[77];
    assign layer0_outputs[6251] = (inputs[167]) | (inputs[138]);
    assign layer0_outputs[6252] = ~(inputs[101]) | (inputs[63]);
    assign layer0_outputs[6253] = inputs[104];
    assign layer0_outputs[6254] = (inputs[132]) ^ (inputs[129]);
    assign layer0_outputs[6255] = ~(inputs[213]);
    assign layer0_outputs[6256] = inputs[232];
    assign layer0_outputs[6257] = ~(inputs[10]) | (inputs[174]);
    assign layer0_outputs[6258] = (inputs[125]) | (inputs[206]);
    assign layer0_outputs[6259] = ~(inputs[145]);
    assign layer0_outputs[6260] = (inputs[159]) & (inputs[190]);
    assign layer0_outputs[6261] = 1'b0;
    assign layer0_outputs[6262] = inputs[225];
    assign layer0_outputs[6263] = ~((inputs[70]) | (inputs[205]));
    assign layer0_outputs[6264] = ~((inputs[123]) & (inputs[242]));
    assign layer0_outputs[6265] = ~((inputs[77]) & (inputs[164]));
    assign layer0_outputs[6266] = ~(inputs[251]);
    assign layer0_outputs[6267] = inputs[114];
    assign layer0_outputs[6268] = 1'b1;
    assign layer0_outputs[6269] = ~(inputs[52]) | (inputs[234]);
    assign layer0_outputs[6270] = (inputs[159]) & ~(inputs[253]);
    assign layer0_outputs[6271] = ~(inputs[104]) | (inputs[239]);
    assign layer0_outputs[6272] = (inputs[140]) & ~(inputs[202]);
    assign layer0_outputs[6273] = ~((inputs[173]) ^ (inputs[212]));
    assign layer0_outputs[6274] = (inputs[52]) & (inputs[143]);
    assign layer0_outputs[6275] = ~(inputs[126]);
    assign layer0_outputs[6276] = (inputs[91]) & ~(inputs[65]);
    assign layer0_outputs[6277] = ~((inputs[151]) | (inputs[252]));
    assign layer0_outputs[6278] = ~(inputs[159]);
    assign layer0_outputs[6279] = ~(inputs[169]);
    assign layer0_outputs[6280] = ~((inputs[158]) ^ (inputs[85]));
    assign layer0_outputs[6281] = ~((inputs[207]) ^ (inputs[219]));
    assign layer0_outputs[6282] = ~((inputs[179]) ^ (inputs[210]));
    assign layer0_outputs[6283] = ~(inputs[33]) | (inputs[82]);
    assign layer0_outputs[6284] = ~(inputs[35]) | (inputs[216]);
    assign layer0_outputs[6285] = 1'b0;
    assign layer0_outputs[6286] = ~(inputs[153]) | (inputs[91]);
    assign layer0_outputs[6287] = ~((inputs[75]) ^ (inputs[87]));
    assign layer0_outputs[6288] = inputs[112];
    assign layer0_outputs[6289] = (inputs[121]) ^ (inputs[186]);
    assign layer0_outputs[6290] = inputs[36];
    assign layer0_outputs[6291] = ~((inputs[175]) ^ (inputs[111]));
    assign layer0_outputs[6292] = ~((inputs[118]) ^ (inputs[197]));
    assign layer0_outputs[6293] = 1'b1;
    assign layer0_outputs[6294] = (inputs[105]) & ~(inputs[111]);
    assign layer0_outputs[6295] = ~(inputs[225]) | (inputs[143]);
    assign layer0_outputs[6296] = ~((inputs[150]) | (inputs[210]));
    assign layer0_outputs[6297] = inputs[134];
    assign layer0_outputs[6298] = ~(inputs[79]);
    assign layer0_outputs[6299] = ~(inputs[182]) | (inputs[91]);
    assign layer0_outputs[6300] = ~(inputs[122]) | (inputs[102]);
    assign layer0_outputs[6301] = 1'b1;
    assign layer0_outputs[6302] = (inputs[240]) | (inputs[125]);
    assign layer0_outputs[6303] = ~(inputs[35]);
    assign layer0_outputs[6304] = (inputs[233]) ^ (inputs[127]);
    assign layer0_outputs[6305] = inputs[150];
    assign layer0_outputs[6306] = (inputs[247]) & ~(inputs[224]);
    assign layer0_outputs[6307] = (inputs[68]) ^ (inputs[147]);
    assign layer0_outputs[6308] = ~(inputs[42]) | (inputs[234]);
    assign layer0_outputs[6309] = ~(inputs[38]) | (inputs[147]);
    assign layer0_outputs[6310] = ~((inputs[255]) | (inputs[127]));
    assign layer0_outputs[6311] = ~((inputs[121]) | (inputs[44]));
    assign layer0_outputs[6312] = inputs[226];
    assign layer0_outputs[6313] = (inputs[85]) ^ (inputs[207]);
    assign layer0_outputs[6314] = ~(inputs[196]);
    assign layer0_outputs[6315] = (inputs[199]) & (inputs[23]);
    assign layer0_outputs[6316] = ~((inputs[245]) | (inputs[49]));
    assign layer0_outputs[6317] = inputs[23];
    assign layer0_outputs[6318] = ~(inputs[9]);
    assign layer0_outputs[6319] = 1'b1;
    assign layer0_outputs[6320] = ~((inputs[246]) | (inputs[143]));
    assign layer0_outputs[6321] = ~(inputs[67]) | (inputs[251]);
    assign layer0_outputs[6322] = ~(inputs[231]);
    assign layer0_outputs[6323] = ~(inputs[193]);
    assign layer0_outputs[6324] = ~(inputs[114]);
    assign layer0_outputs[6325] = ~((inputs[41]) ^ (inputs[101]));
    assign layer0_outputs[6326] = ~((inputs[108]) ^ (inputs[63]));
    assign layer0_outputs[6327] = 1'b1;
    assign layer0_outputs[6328] = (inputs[25]) & (inputs[80]);
    assign layer0_outputs[6329] = (inputs[219]) | (inputs[158]);
    assign layer0_outputs[6330] = (inputs[169]) & ~(inputs[120]);
    assign layer0_outputs[6331] = ~((inputs[91]) | (inputs[2]));
    assign layer0_outputs[6332] = ~((inputs[219]) | (inputs[64]));
    assign layer0_outputs[6333] = ~(inputs[200]) | (inputs[131]);
    assign layer0_outputs[6334] = inputs[23];
    assign layer0_outputs[6335] = (inputs[188]) & ~(inputs[179]);
    assign layer0_outputs[6336] = ~((inputs[128]) ^ (inputs[151]));
    assign layer0_outputs[6337] = ~(inputs[160]) | (inputs[140]);
    assign layer0_outputs[6338] = (inputs[55]) ^ (inputs[84]);
    assign layer0_outputs[6339] = ~((inputs[105]) ^ (inputs[124]));
    assign layer0_outputs[6340] = inputs[70];
    assign layer0_outputs[6341] = ~(inputs[230]) | (inputs[106]);
    assign layer0_outputs[6342] = (inputs[13]) | (inputs[86]);
    assign layer0_outputs[6343] = (inputs[117]) & ~(inputs[222]);
    assign layer0_outputs[6344] = ~(inputs[107]);
    assign layer0_outputs[6345] = (inputs[61]) & ~(inputs[48]);
    assign layer0_outputs[6346] = inputs[94];
    assign layer0_outputs[6347] = (inputs[82]) & ~(inputs[55]);
    assign layer0_outputs[6348] = (inputs[234]) ^ (inputs[204]);
    assign layer0_outputs[6349] = ~(inputs[176]);
    assign layer0_outputs[6350] = inputs[156];
    assign layer0_outputs[6351] = 1'b0;
    assign layer0_outputs[6352] = ~(inputs[138]);
    assign layer0_outputs[6353] = inputs[10];
    assign layer0_outputs[6354] = (inputs[79]) | (inputs[50]);
    assign layer0_outputs[6355] = (inputs[74]) & ~(inputs[144]);
    assign layer0_outputs[6356] = 1'b1;
    assign layer0_outputs[6357] = inputs[73];
    assign layer0_outputs[6358] = ~(inputs[172]) | (inputs[50]);
    assign layer0_outputs[6359] = ~(inputs[134]) | (inputs[141]);
    assign layer0_outputs[6360] = inputs[39];
    assign layer0_outputs[6361] = inputs[148];
    assign layer0_outputs[6362] = ~(inputs[37]);
    assign layer0_outputs[6363] = (inputs[81]) ^ (inputs[86]);
    assign layer0_outputs[6364] = inputs[178];
    assign layer0_outputs[6365] = inputs[116];
    assign layer0_outputs[6366] = inputs[204];
    assign layer0_outputs[6367] = inputs[21];
    assign layer0_outputs[6368] = inputs[49];
    assign layer0_outputs[6369] = ~(inputs[100]);
    assign layer0_outputs[6370] = ~(inputs[164]);
    assign layer0_outputs[6371] = ~(inputs[109]);
    assign layer0_outputs[6372] = 1'b1;
    assign layer0_outputs[6373] = ~(inputs[84]);
    assign layer0_outputs[6374] = (inputs[64]) & ~(inputs[68]);
    assign layer0_outputs[6375] = (inputs[144]) | (inputs[84]);
    assign layer0_outputs[6376] = inputs[209];
    assign layer0_outputs[6377] = (inputs[221]) & ~(inputs[141]);
    assign layer0_outputs[6378] = (inputs[26]) & ~(inputs[178]);
    assign layer0_outputs[6379] = ~((inputs[5]) | (inputs[20]));
    assign layer0_outputs[6380] = (inputs[140]) ^ (inputs[5]);
    assign layer0_outputs[6381] = (inputs[54]) & ~(inputs[255]);
    assign layer0_outputs[6382] = (inputs[43]) ^ (inputs[65]);
    assign layer0_outputs[6383] = (inputs[134]) | (inputs[172]);
    assign layer0_outputs[6384] = ~(inputs[152]);
    assign layer0_outputs[6385] = ~((inputs[204]) | (inputs[205]));
    assign layer0_outputs[6386] = ~(inputs[56]) | (inputs[143]);
    assign layer0_outputs[6387] = ~((inputs[5]) ^ (inputs[81]));
    assign layer0_outputs[6388] = inputs[62];
    assign layer0_outputs[6389] = ~(inputs[4]) | (inputs[80]);
    assign layer0_outputs[6390] = (inputs[37]) & ~(inputs[113]);
    assign layer0_outputs[6391] = (inputs[126]) ^ (inputs[27]);
    assign layer0_outputs[6392] = ~(inputs[62]) | (inputs[173]);
    assign layer0_outputs[6393] = ~(inputs[230]);
    assign layer0_outputs[6394] = (inputs[64]) | (inputs[209]);
    assign layer0_outputs[6395] = ~((inputs[157]) ^ (inputs[94]));
    assign layer0_outputs[6396] = ~((inputs[164]) | (inputs[83]));
    assign layer0_outputs[6397] = ~((inputs[0]) | (inputs[73]));
    assign layer0_outputs[6398] = ~(inputs[39]);
    assign layer0_outputs[6399] = (inputs[29]) ^ (inputs[192]);
    assign layer0_outputs[6400] = ~((inputs[238]) | (inputs[30]));
    assign layer0_outputs[6401] = ~((inputs[5]) | (inputs[89]));
    assign layer0_outputs[6402] = (inputs[171]) & ~(inputs[169]);
    assign layer0_outputs[6403] = ~((inputs[79]) ^ (inputs[92]));
    assign layer0_outputs[6404] = (inputs[29]) & ~(inputs[55]);
    assign layer0_outputs[6405] = (inputs[175]) & ~(inputs[14]);
    assign layer0_outputs[6406] = inputs[169];
    assign layer0_outputs[6407] = ~(inputs[172]) | (inputs[30]);
    assign layer0_outputs[6408] = ~((inputs[221]) | (inputs[17]));
    assign layer0_outputs[6409] = inputs[25];
    assign layer0_outputs[6410] = inputs[183];
    assign layer0_outputs[6411] = ~(inputs[184]) | (inputs[18]);
    assign layer0_outputs[6412] = ~(inputs[11]);
    assign layer0_outputs[6413] = inputs[163];
    assign layer0_outputs[6414] = ~(inputs[68]);
    assign layer0_outputs[6415] = inputs[113];
    assign layer0_outputs[6416] = (inputs[187]) & ~(inputs[33]);
    assign layer0_outputs[6417] = ~((inputs[85]) ^ (inputs[223]));
    assign layer0_outputs[6418] = (inputs[233]) | (inputs[223]);
    assign layer0_outputs[6419] = inputs[24];
    assign layer0_outputs[6420] = inputs[117];
    assign layer0_outputs[6421] = (inputs[216]) & ~(inputs[98]);
    assign layer0_outputs[6422] = (inputs[235]) | (inputs[185]);
    assign layer0_outputs[6423] = (inputs[234]) & ~(inputs[79]);
    assign layer0_outputs[6424] = (inputs[148]) | (inputs[5]);
    assign layer0_outputs[6425] = ~(inputs[161]);
    assign layer0_outputs[6426] = 1'b1;
    assign layer0_outputs[6427] = inputs[64];
    assign layer0_outputs[6428] = ~(inputs[128]);
    assign layer0_outputs[6429] = (inputs[221]) | (inputs[92]);
    assign layer0_outputs[6430] = 1'b1;
    assign layer0_outputs[6431] = (inputs[117]) & ~(inputs[47]);
    assign layer0_outputs[6432] = (inputs[148]) & ~(inputs[91]);
    assign layer0_outputs[6433] = (inputs[89]) & ~(inputs[219]);
    assign layer0_outputs[6434] = ~(inputs[140]) | (inputs[36]);
    assign layer0_outputs[6435] = (inputs[234]) & ~(inputs[114]);
    assign layer0_outputs[6436] = ~(inputs[63]);
    assign layer0_outputs[6437] = (inputs[101]) & ~(inputs[127]);
    assign layer0_outputs[6438] = inputs[26];
    assign layer0_outputs[6439] = ~(inputs[220]) | (inputs[66]);
    assign layer0_outputs[6440] = ~(inputs[54]) | (inputs[126]);
    assign layer0_outputs[6441] = ~(inputs[163]) | (inputs[81]);
    assign layer0_outputs[6442] = inputs[248];
    assign layer0_outputs[6443] = inputs[138];
    assign layer0_outputs[6444] = ~(inputs[68]) | (inputs[48]);
    assign layer0_outputs[6445] = ~(inputs[241]);
    assign layer0_outputs[6446] = (inputs[31]) | (inputs[164]);
    assign layer0_outputs[6447] = ~(inputs[160]);
    assign layer0_outputs[6448] = ~(inputs[196]);
    assign layer0_outputs[6449] = 1'b0;
    assign layer0_outputs[6450] = ~(inputs[116]) | (inputs[237]);
    assign layer0_outputs[6451] = ~((inputs[184]) | (inputs[131]));
    assign layer0_outputs[6452] = ~((inputs[251]) | (inputs[243]));
    assign layer0_outputs[6453] = ~(inputs[218]) | (inputs[110]);
    assign layer0_outputs[6454] = (inputs[63]) | (inputs[2]);
    assign layer0_outputs[6455] = ~((inputs[80]) | (inputs[221]));
    assign layer0_outputs[6456] = (inputs[138]) & ~(inputs[10]);
    assign layer0_outputs[6457] = ~(inputs[127]) | (inputs[29]);
    assign layer0_outputs[6458] = (inputs[253]) ^ (inputs[19]);
    assign layer0_outputs[6459] = ~(inputs[115]);
    assign layer0_outputs[6460] = ~((inputs[188]) ^ (inputs[219]));
    assign layer0_outputs[6461] = inputs[80];
    assign layer0_outputs[6462] = inputs[83];
    assign layer0_outputs[6463] = inputs[27];
    assign layer0_outputs[6464] = inputs[8];
    assign layer0_outputs[6465] = ~((inputs[236]) ^ (inputs[178]));
    assign layer0_outputs[6466] = ~((inputs[88]) | (inputs[59]));
    assign layer0_outputs[6467] = ~(inputs[25]);
    assign layer0_outputs[6468] = (inputs[144]) ^ (inputs[205]);
    assign layer0_outputs[6469] = ~(inputs[142]) | (inputs[153]);
    assign layer0_outputs[6470] = ~((inputs[28]) | (inputs[21]));
    assign layer0_outputs[6471] = inputs[126];
    assign layer0_outputs[6472] = ~((inputs[202]) ^ (inputs[220]));
    assign layer0_outputs[6473] = ~((inputs[228]) | (inputs[99]));
    assign layer0_outputs[6474] = (inputs[138]) ^ (inputs[139]);
    assign layer0_outputs[6475] = (inputs[243]) ^ (inputs[212]);
    assign layer0_outputs[6476] = (inputs[224]) ^ (inputs[172]);
    assign layer0_outputs[6477] = (inputs[172]) | (inputs[31]);
    assign layer0_outputs[6478] = (inputs[157]) & ~(inputs[131]);
    assign layer0_outputs[6479] = inputs[32];
    assign layer0_outputs[6480] = ~(inputs[54]);
    assign layer0_outputs[6481] = ~(inputs[165]) | (inputs[242]);
    assign layer0_outputs[6482] = inputs[43];
    assign layer0_outputs[6483] = ~((inputs[25]) ^ (inputs[49]));
    assign layer0_outputs[6484] = ~(inputs[1]) | (inputs[169]);
    assign layer0_outputs[6485] = (inputs[213]) | (inputs[250]);
    assign layer0_outputs[6486] = ~((inputs[115]) & (inputs[212]));
    assign layer0_outputs[6487] = (inputs[246]) & ~(inputs[107]);
    assign layer0_outputs[6488] = (inputs[87]) | (inputs[86]);
    assign layer0_outputs[6489] = (inputs[74]) ^ (inputs[171]);
    assign layer0_outputs[6490] = (inputs[125]) | (inputs[92]);
    assign layer0_outputs[6491] = (inputs[231]) ^ (inputs[125]);
    assign layer0_outputs[6492] = (inputs[11]) | (inputs[51]);
    assign layer0_outputs[6493] = inputs[223];
    assign layer0_outputs[6494] = inputs[169];
    assign layer0_outputs[6495] = (inputs[22]) ^ (inputs[64]);
    assign layer0_outputs[6496] = inputs[174];
    assign layer0_outputs[6497] = 1'b0;
    assign layer0_outputs[6498] = inputs[214];
    assign layer0_outputs[6499] = (inputs[161]) ^ (inputs[231]);
    assign layer0_outputs[6500] = ~((inputs[176]) ^ (inputs[227]));
    assign layer0_outputs[6501] = ~((inputs[53]) ^ (inputs[7]));
    assign layer0_outputs[6502] = ~(inputs[28]);
    assign layer0_outputs[6503] = ~(inputs[207]) | (inputs[133]);
    assign layer0_outputs[6504] = (inputs[236]) | (inputs[118]);
    assign layer0_outputs[6505] = (inputs[68]) | (inputs[13]);
    assign layer0_outputs[6506] = (inputs[119]) | (inputs[167]);
    assign layer0_outputs[6507] = ~((inputs[253]) & (inputs[128]));
    assign layer0_outputs[6508] = (inputs[44]) | (inputs[169]);
    assign layer0_outputs[6509] = ~((inputs[213]) | (inputs[191]));
    assign layer0_outputs[6510] = (inputs[127]) & ~(inputs[191]);
    assign layer0_outputs[6511] = ~((inputs[90]) | (inputs[16]));
    assign layer0_outputs[6512] = ~((inputs[207]) | (inputs[204]));
    assign layer0_outputs[6513] = inputs[142];
    assign layer0_outputs[6514] = inputs[42];
    assign layer0_outputs[6515] = (inputs[205]) | (inputs[217]);
    assign layer0_outputs[6516] = ~((inputs[243]) | (inputs[109]));
    assign layer0_outputs[6517] = inputs[91];
    assign layer0_outputs[6518] = 1'b1;
    assign layer0_outputs[6519] = (inputs[180]) ^ (inputs[182]);
    assign layer0_outputs[6520] = (inputs[53]) ^ (inputs[38]);
    assign layer0_outputs[6521] = ~((inputs[91]) & (inputs[140]));
    assign layer0_outputs[6522] = 1'b1;
    assign layer0_outputs[6523] = (inputs[36]) & ~(inputs[252]);
    assign layer0_outputs[6524] = inputs[75];
    assign layer0_outputs[6525] = inputs[94];
    assign layer0_outputs[6526] = inputs[58];
    assign layer0_outputs[6527] = ~(inputs[165]) | (inputs[191]);
    assign layer0_outputs[6528] = ~((inputs[185]) | (inputs[252]));
    assign layer0_outputs[6529] = (inputs[126]) | (inputs[81]);
    assign layer0_outputs[6530] = ~((inputs[99]) | (inputs[98]));
    assign layer0_outputs[6531] = 1'b0;
    assign layer0_outputs[6532] = inputs[101];
    assign layer0_outputs[6533] = ~((inputs[18]) ^ (inputs[105]));
    assign layer0_outputs[6534] = ~(inputs[66]);
    assign layer0_outputs[6535] = (inputs[189]) & ~(inputs[204]);
    assign layer0_outputs[6536] = ~(inputs[249]);
    assign layer0_outputs[6537] = ~(inputs[72]);
    assign layer0_outputs[6538] = ~(inputs[178]);
    assign layer0_outputs[6539] = inputs[20];
    assign layer0_outputs[6540] = (inputs[255]) ^ (inputs[102]);
    assign layer0_outputs[6541] = ~(inputs[213]) | (inputs[31]);
    assign layer0_outputs[6542] = (inputs[39]) ^ (inputs[116]);
    assign layer0_outputs[6543] = (inputs[44]) & ~(inputs[11]);
    assign layer0_outputs[6544] = ~(inputs[77]);
    assign layer0_outputs[6545] = ~((inputs[33]) | (inputs[45]));
    assign layer0_outputs[6546] = ~(inputs[245]) | (inputs[53]);
    assign layer0_outputs[6547] = (inputs[102]) & ~(inputs[254]);
    assign layer0_outputs[6548] = ~(inputs[43]);
    assign layer0_outputs[6549] = ~(inputs[253]);
    assign layer0_outputs[6550] = inputs[213];
    assign layer0_outputs[6551] = ~(inputs[212]);
    assign layer0_outputs[6552] = ~((inputs[244]) | (inputs[187]));
    assign layer0_outputs[6553] = ~(inputs[120]) | (inputs[178]);
    assign layer0_outputs[6554] = (inputs[227]) & ~(inputs[107]);
    assign layer0_outputs[6555] = 1'b0;
    assign layer0_outputs[6556] = (inputs[169]) ^ (inputs[106]);
    assign layer0_outputs[6557] = ~((inputs[201]) | (inputs[97]));
    assign layer0_outputs[6558] = ~((inputs[65]) | (inputs[166]));
    assign layer0_outputs[6559] = inputs[72];
    assign layer0_outputs[6560] = ~(inputs[7]) | (inputs[239]);
    assign layer0_outputs[6561] = inputs[219];
    assign layer0_outputs[6562] = ~((inputs[17]) | (inputs[187]));
    assign layer0_outputs[6563] = ~(inputs[143]);
    assign layer0_outputs[6564] = ~(inputs[23]) | (inputs[20]);
    assign layer0_outputs[6565] = (inputs[107]) ^ (inputs[105]);
    assign layer0_outputs[6566] = 1'b1;
    assign layer0_outputs[6567] = (inputs[41]) | (inputs[145]);
    assign layer0_outputs[6568] = inputs[193];
    assign layer0_outputs[6569] = (inputs[51]) | (inputs[165]);
    assign layer0_outputs[6570] = (inputs[226]) & (inputs[200]);
    assign layer0_outputs[6571] = inputs[199];
    assign layer0_outputs[6572] = ~(inputs[100]);
    assign layer0_outputs[6573] = inputs[119];
    assign layer0_outputs[6574] = ~(inputs[105]);
    assign layer0_outputs[6575] = inputs[112];
    assign layer0_outputs[6576] = inputs[76];
    assign layer0_outputs[6577] = ~((inputs[61]) ^ (inputs[254]));
    assign layer0_outputs[6578] = ~((inputs[57]) | (inputs[157]));
    assign layer0_outputs[6579] = ~(inputs[127]);
    assign layer0_outputs[6580] = ~((inputs[83]) | (inputs[63]));
    assign layer0_outputs[6581] = inputs[60];
    assign layer0_outputs[6582] = (inputs[179]) | (inputs[157]);
    assign layer0_outputs[6583] = ~(inputs[76]) | (inputs[229]);
    assign layer0_outputs[6584] = ~((inputs[198]) ^ (inputs[228]));
    assign layer0_outputs[6585] = inputs[0];
    assign layer0_outputs[6586] = (inputs[248]) & ~(inputs[43]);
    assign layer0_outputs[6587] = (inputs[24]) & ~(inputs[113]);
    assign layer0_outputs[6588] = inputs[181];
    assign layer0_outputs[6589] = ~(inputs[84]);
    assign layer0_outputs[6590] = ~(inputs[130]);
    assign layer0_outputs[6591] = (inputs[52]) & (inputs[139]);
    assign layer0_outputs[6592] = ~(inputs[101]);
    assign layer0_outputs[6593] = ~(inputs[6]) | (inputs[80]);
    assign layer0_outputs[6594] = 1'b1;
    assign layer0_outputs[6595] = ~(inputs[18]) | (inputs[95]);
    assign layer0_outputs[6596] = (inputs[74]) | (inputs[142]);
    assign layer0_outputs[6597] = (inputs[177]) ^ (inputs[246]);
    assign layer0_outputs[6598] = (inputs[121]) & ~(inputs[239]);
    assign layer0_outputs[6599] = inputs[195];
    assign layer0_outputs[6600] = ~(inputs[218]);
    assign layer0_outputs[6601] = ~(inputs[9]);
    assign layer0_outputs[6602] = inputs[213];
    assign layer0_outputs[6603] = ~(inputs[54]) | (inputs[106]);
    assign layer0_outputs[6604] = ~(inputs[135]) | (inputs[195]);
    assign layer0_outputs[6605] = (inputs[112]) & ~(inputs[47]);
    assign layer0_outputs[6606] = ~(inputs[242]) | (inputs[43]);
    assign layer0_outputs[6607] = (inputs[162]) & ~(inputs[63]);
    assign layer0_outputs[6608] = ~((inputs[194]) & (inputs[120]));
    assign layer0_outputs[6609] = 1'b0;
    assign layer0_outputs[6610] = (inputs[71]) & (inputs[19]);
    assign layer0_outputs[6611] = ~((inputs[147]) | (inputs[219]));
    assign layer0_outputs[6612] = ~((inputs[90]) | (inputs[75]));
    assign layer0_outputs[6613] = (inputs[179]) | (inputs[43]);
    assign layer0_outputs[6614] = (inputs[111]) ^ (inputs[26]);
    assign layer0_outputs[6615] = 1'b1;
    assign layer0_outputs[6616] = ~(inputs[226]) | (inputs[139]);
    assign layer0_outputs[6617] = ~(inputs[137]) | (inputs[93]);
    assign layer0_outputs[6618] = (inputs[219]) & (inputs[239]);
    assign layer0_outputs[6619] = ~(inputs[43]);
    assign layer0_outputs[6620] = ~((inputs[170]) | (inputs[131]));
    assign layer0_outputs[6621] = ~(inputs[40]);
    assign layer0_outputs[6622] = inputs[114];
    assign layer0_outputs[6623] = (inputs[0]) ^ (inputs[247]);
    assign layer0_outputs[6624] = ~((inputs[160]) ^ (inputs[92]));
    assign layer0_outputs[6625] = ~((inputs[171]) ^ (inputs[155]));
    assign layer0_outputs[6626] = (inputs[190]) & ~(inputs[66]);
    assign layer0_outputs[6627] = ~((inputs[52]) | (inputs[228]));
    assign layer0_outputs[6628] = (inputs[18]) ^ (inputs[202]);
    assign layer0_outputs[6629] = ~((inputs[232]) | (inputs[51]));
    assign layer0_outputs[6630] = ~(inputs[178]);
    assign layer0_outputs[6631] = inputs[102];
    assign layer0_outputs[6632] = ~(inputs[173]);
    assign layer0_outputs[6633] = ~(inputs[103]);
    assign layer0_outputs[6634] = ~((inputs[93]) | (inputs[218]));
    assign layer0_outputs[6635] = (inputs[137]) & (inputs[10]);
    assign layer0_outputs[6636] = inputs[122];
    assign layer0_outputs[6637] = ~((inputs[221]) ^ (inputs[157]));
    assign layer0_outputs[6638] = (inputs[86]) ^ (inputs[144]);
    assign layer0_outputs[6639] = (inputs[106]) & ~(inputs[182]);
    assign layer0_outputs[6640] = (inputs[162]) ^ (inputs[245]);
    assign layer0_outputs[6641] = (inputs[227]) & ~(inputs[150]);
    assign layer0_outputs[6642] = ~((inputs[53]) | (inputs[65]));
    assign layer0_outputs[6643] = inputs[168];
    assign layer0_outputs[6644] = ~((inputs[250]) & (inputs[189]));
    assign layer0_outputs[6645] = (inputs[14]) & ~(inputs[199]);
    assign layer0_outputs[6646] = ~((inputs[72]) & (inputs[108]));
    assign layer0_outputs[6647] = ~((inputs[162]) | (inputs[92]));
    assign layer0_outputs[6648] = ~(inputs[58]);
    assign layer0_outputs[6649] = inputs[122];
    assign layer0_outputs[6650] = (inputs[22]) ^ (inputs[101]);
    assign layer0_outputs[6651] = inputs[129];
    assign layer0_outputs[6652] = ~(inputs[85]);
    assign layer0_outputs[6653] = ~(inputs[181]);
    assign layer0_outputs[6654] = inputs[231];
    assign layer0_outputs[6655] = ~(inputs[56]);
    assign layer0_outputs[6656] = ~(inputs[130]);
    assign layer0_outputs[6657] = ~(inputs[127]);
    assign layer0_outputs[6658] = (inputs[94]) & (inputs[52]);
    assign layer0_outputs[6659] = ~(inputs[181]);
    assign layer0_outputs[6660] = (inputs[254]) & ~(inputs[56]);
    assign layer0_outputs[6661] = ~(inputs[67]);
    assign layer0_outputs[6662] = ~(inputs[124]);
    assign layer0_outputs[6663] = inputs[132];
    assign layer0_outputs[6664] = inputs[228];
    assign layer0_outputs[6665] = ~(inputs[20]);
    assign layer0_outputs[6666] = inputs[137];
    assign layer0_outputs[6667] = ~(inputs[7]);
    assign layer0_outputs[6668] = (inputs[75]) & ~(inputs[136]);
    assign layer0_outputs[6669] = ~((inputs[202]) | (inputs[110]));
    assign layer0_outputs[6670] = ~((inputs[146]) | (inputs[30]));
    assign layer0_outputs[6671] = inputs[108];
    assign layer0_outputs[6672] = inputs[208];
    assign layer0_outputs[6673] = inputs[121];
    assign layer0_outputs[6674] = (inputs[105]) | (inputs[155]);
    assign layer0_outputs[6675] = ~((inputs[74]) | (inputs[80]));
    assign layer0_outputs[6676] = ~(inputs[129]);
    assign layer0_outputs[6677] = (inputs[174]) & ~(inputs[46]);
    assign layer0_outputs[6678] = ~((inputs[211]) | (inputs[57]));
    assign layer0_outputs[6679] = inputs[55];
    assign layer0_outputs[6680] = 1'b1;
    assign layer0_outputs[6681] = ~(inputs[64]);
    assign layer0_outputs[6682] = inputs[20];
    assign layer0_outputs[6683] = ~((inputs[3]) | (inputs[154]));
    assign layer0_outputs[6684] = ~(inputs[245]);
    assign layer0_outputs[6685] = (inputs[172]) | (inputs[238]);
    assign layer0_outputs[6686] = ~((inputs[109]) ^ (inputs[34]));
    assign layer0_outputs[6687] = ~((inputs[18]) ^ (inputs[26]));
    assign layer0_outputs[6688] = ~((inputs[97]) ^ (inputs[102]));
    assign layer0_outputs[6689] = (inputs[188]) | (inputs[144]);
    assign layer0_outputs[6690] = (inputs[188]) ^ (inputs[189]);
    assign layer0_outputs[6691] = (inputs[79]) ^ (inputs[2]);
    assign layer0_outputs[6692] = ~((inputs[150]) | (inputs[52]));
    assign layer0_outputs[6693] = (inputs[206]) | (inputs[230]);
    assign layer0_outputs[6694] = 1'b0;
    assign layer0_outputs[6695] = inputs[218];
    assign layer0_outputs[6696] = ~((inputs[37]) | (inputs[77]));
    assign layer0_outputs[6697] = ~(inputs[24]);
    assign layer0_outputs[6698] = inputs[84];
    assign layer0_outputs[6699] = ~((inputs[90]) ^ (inputs[242]));
    assign layer0_outputs[6700] = (inputs[225]) | (inputs[205]);
    assign layer0_outputs[6701] = ~(inputs[52]) | (inputs[83]);
    assign layer0_outputs[6702] = inputs[172];
    assign layer0_outputs[6703] = ~(inputs[2]);
    assign layer0_outputs[6704] = ~(inputs[193]);
    assign layer0_outputs[6705] = ~((inputs[188]) | (inputs[210]));
    assign layer0_outputs[6706] = ~(inputs[9]);
    assign layer0_outputs[6707] = (inputs[162]) | (inputs[152]);
    assign layer0_outputs[6708] = (inputs[115]) | (inputs[117]);
    assign layer0_outputs[6709] = ~((inputs[0]) ^ (inputs[118]));
    assign layer0_outputs[6710] = (inputs[230]) ^ (inputs[168]);
    assign layer0_outputs[6711] = (inputs[252]) | (inputs[116]);
    assign layer0_outputs[6712] = (inputs[70]) | (inputs[172]);
    assign layer0_outputs[6713] = (inputs[120]) | (inputs[30]);
    assign layer0_outputs[6714] = 1'b0;
    assign layer0_outputs[6715] = inputs[22];
    assign layer0_outputs[6716] = ~(inputs[62]);
    assign layer0_outputs[6717] = ~(inputs[107]) | (inputs[127]);
    assign layer0_outputs[6718] = (inputs[198]) & ~(inputs[63]);
    assign layer0_outputs[6719] = inputs[23];
    assign layer0_outputs[6720] = ~(inputs[109]);
    assign layer0_outputs[6721] = (inputs[83]) | (inputs[38]);
    assign layer0_outputs[6722] = (inputs[77]) ^ (inputs[228]);
    assign layer0_outputs[6723] = (inputs[0]) & ~(inputs[6]);
    assign layer0_outputs[6724] = inputs[194];
    assign layer0_outputs[6725] = (inputs[249]) | (inputs[56]);
    assign layer0_outputs[6726] = inputs[83];
    assign layer0_outputs[6727] = ~(inputs[187]);
    assign layer0_outputs[6728] = inputs[173];
    assign layer0_outputs[6729] = ~(inputs[118]) | (inputs[6]);
    assign layer0_outputs[6730] = ~((inputs[42]) ^ (inputs[11]));
    assign layer0_outputs[6731] = ~((inputs[239]) | (inputs[70]));
    assign layer0_outputs[6732] = inputs[140];
    assign layer0_outputs[6733] = (inputs[20]) & ~(inputs[224]);
    assign layer0_outputs[6734] = ~((inputs[9]) ^ (inputs[111]));
    assign layer0_outputs[6735] = ~((inputs[38]) ^ (inputs[160]));
    assign layer0_outputs[6736] = (inputs[243]) ^ (inputs[169]);
    assign layer0_outputs[6737] = inputs[163];
    assign layer0_outputs[6738] = ~(inputs[187]) | (inputs[0]);
    assign layer0_outputs[6739] = inputs[214];
    assign layer0_outputs[6740] = ~((inputs[177]) ^ (inputs[22]));
    assign layer0_outputs[6741] = ~(inputs[54]);
    assign layer0_outputs[6742] = ~((inputs[0]) & (inputs[159]));
    assign layer0_outputs[6743] = ~(inputs[61]);
    assign layer0_outputs[6744] = (inputs[120]) & ~(inputs[1]);
    assign layer0_outputs[6745] = ~((inputs[252]) ^ (inputs[89]));
    assign layer0_outputs[6746] = (inputs[24]) & ~(inputs[222]);
    assign layer0_outputs[6747] = ~(inputs[200]) | (inputs[46]);
    assign layer0_outputs[6748] = 1'b0;
    assign layer0_outputs[6749] = (inputs[90]) | (inputs[73]);
    assign layer0_outputs[6750] = (inputs[171]) & (inputs[181]);
    assign layer0_outputs[6751] = (inputs[108]) & ~(inputs[47]);
    assign layer0_outputs[6752] = inputs[200];
    assign layer0_outputs[6753] = (inputs[97]) ^ (inputs[71]);
    assign layer0_outputs[6754] = (inputs[44]) | (inputs[15]);
    assign layer0_outputs[6755] = (inputs[95]) | (inputs[193]);
    assign layer0_outputs[6756] = ~((inputs[228]) ^ (inputs[155]));
    assign layer0_outputs[6757] = ~((inputs[147]) | (inputs[20]));
    assign layer0_outputs[6758] = inputs[94];
    assign layer0_outputs[6759] = ~((inputs[110]) & (inputs[139]));
    assign layer0_outputs[6760] = ~(inputs[151]);
    assign layer0_outputs[6761] = (inputs[123]) & (inputs[18]);
    assign layer0_outputs[6762] = (inputs[101]) & (inputs[171]);
    assign layer0_outputs[6763] = ~(inputs[36]) | (inputs[0]);
    assign layer0_outputs[6764] = (inputs[23]) ^ (inputs[51]);
    assign layer0_outputs[6765] = ~(inputs[179]) | (inputs[135]);
    assign layer0_outputs[6766] = ~(inputs[207]) | (inputs[201]);
    assign layer0_outputs[6767] = (inputs[36]) & ~(inputs[216]);
    assign layer0_outputs[6768] = ~(inputs[90]) | (inputs[161]);
    assign layer0_outputs[6769] = (inputs[88]) & (inputs[240]);
    assign layer0_outputs[6770] = ~(inputs[211]);
    assign layer0_outputs[6771] = ~(inputs[253]);
    assign layer0_outputs[6772] = (inputs[57]) & (inputs[126]);
    assign layer0_outputs[6773] = inputs[170];
    assign layer0_outputs[6774] = ~(inputs[162]);
    assign layer0_outputs[6775] = (inputs[6]) & (inputs[71]);
    assign layer0_outputs[6776] = (inputs[178]) & (inputs[139]);
    assign layer0_outputs[6777] = (inputs[244]) | (inputs[11]);
    assign layer0_outputs[6778] = inputs[51];
    assign layer0_outputs[6779] = inputs[108];
    assign layer0_outputs[6780] = ~((inputs[5]) | (inputs[78]));
    assign layer0_outputs[6781] = ~(inputs[99]);
    assign layer0_outputs[6782] = ~((inputs[247]) ^ (inputs[237]));
    assign layer0_outputs[6783] = (inputs[25]) | (inputs[35]);
    assign layer0_outputs[6784] = (inputs[156]) & ~(inputs[135]);
    assign layer0_outputs[6785] = ~((inputs[2]) | (inputs[29]));
    assign layer0_outputs[6786] = ~((inputs[90]) | (inputs[4]));
    assign layer0_outputs[6787] = ~((inputs[105]) | (inputs[153]));
    assign layer0_outputs[6788] = (inputs[23]) & ~(inputs[96]);
    assign layer0_outputs[6789] = (inputs[196]) & ~(inputs[78]);
    assign layer0_outputs[6790] = ~((inputs[95]) & (inputs[139]));
    assign layer0_outputs[6791] = 1'b1;
    assign layer0_outputs[6792] = ~(inputs[125]);
    assign layer0_outputs[6793] = (inputs[178]) & ~(inputs[18]);
    assign layer0_outputs[6794] = ~(inputs[29]);
    assign layer0_outputs[6795] = inputs[223];
    assign layer0_outputs[6796] = (inputs[172]) & (inputs[248]);
    assign layer0_outputs[6797] = (inputs[104]) ^ (inputs[89]);
    assign layer0_outputs[6798] = ~(inputs[65]);
    assign layer0_outputs[6799] = ~(inputs[169]);
    assign layer0_outputs[6800] = ~(inputs[107]);
    assign layer0_outputs[6801] = (inputs[137]) & (inputs[68]);
    assign layer0_outputs[6802] = (inputs[61]) | (inputs[39]);
    assign layer0_outputs[6803] = (inputs[247]) ^ (inputs[18]);
    assign layer0_outputs[6804] = inputs[108];
    assign layer0_outputs[6805] = inputs[182];
    assign layer0_outputs[6806] = ~(inputs[39]);
    assign layer0_outputs[6807] = 1'b1;
    assign layer0_outputs[6808] = ~(inputs[133]) | (inputs[70]);
    assign layer0_outputs[6809] = (inputs[157]) | (inputs[205]);
    assign layer0_outputs[6810] = (inputs[99]) | (inputs[96]);
    assign layer0_outputs[6811] = ~(inputs[36]);
    assign layer0_outputs[6812] = (inputs[163]) & ~(inputs[107]);
    assign layer0_outputs[6813] = (inputs[193]) | (inputs[194]);
    assign layer0_outputs[6814] = ~((inputs[253]) ^ (inputs[144]));
    assign layer0_outputs[6815] = (inputs[193]) ^ (inputs[229]);
    assign layer0_outputs[6816] = ~((inputs[12]) | (inputs[163]));
    assign layer0_outputs[6817] = ~(inputs[114]);
    assign layer0_outputs[6818] = inputs[82];
    assign layer0_outputs[6819] = (inputs[18]) | (inputs[199]);
    assign layer0_outputs[6820] = (inputs[186]) & ~(inputs[16]);
    assign layer0_outputs[6821] = ~((inputs[182]) | (inputs[66]));
    assign layer0_outputs[6822] = ~((inputs[23]) | (inputs[94]));
    assign layer0_outputs[6823] = ~((inputs[80]) ^ (inputs[9]));
    assign layer0_outputs[6824] = ~(inputs[44]);
    assign layer0_outputs[6825] = ~((inputs[203]) & (inputs[90]));
    assign layer0_outputs[6826] = inputs[94];
    assign layer0_outputs[6827] = ~((inputs[217]) | (inputs[116]));
    assign layer0_outputs[6828] = ~((inputs[67]) ^ (inputs[69]));
    assign layer0_outputs[6829] = ~(inputs[189]);
    assign layer0_outputs[6830] = (inputs[194]) & ~(inputs[21]);
    assign layer0_outputs[6831] = inputs[194];
    assign layer0_outputs[6832] = inputs[247];
    assign layer0_outputs[6833] = (inputs[187]) ^ (inputs[161]);
    assign layer0_outputs[6834] = (inputs[17]) | (inputs[71]);
    assign layer0_outputs[6835] = (inputs[167]) & (inputs[41]);
    assign layer0_outputs[6836] = ~(inputs[191]);
    assign layer0_outputs[6837] = ~((inputs[218]) ^ (inputs[15]));
    assign layer0_outputs[6838] = ~((inputs[197]) ^ (inputs[229]));
    assign layer0_outputs[6839] = 1'b0;
    assign layer0_outputs[6840] = ~((inputs[182]) ^ (inputs[162]));
    assign layer0_outputs[6841] = ~(inputs[50]) | (inputs[217]);
    assign layer0_outputs[6842] = ~(inputs[95]);
    assign layer0_outputs[6843] = (inputs[60]) ^ (inputs[22]);
    assign layer0_outputs[6844] = ~(inputs[45]);
    assign layer0_outputs[6845] = ~(inputs[35]);
    assign layer0_outputs[6846] = (inputs[129]) ^ (inputs[74]);
    assign layer0_outputs[6847] = inputs[92];
    assign layer0_outputs[6848] = ~(inputs[75]);
    assign layer0_outputs[6849] = 1'b1;
    assign layer0_outputs[6850] = ~(inputs[1]);
    assign layer0_outputs[6851] = ~((inputs[208]) ^ (inputs[189]));
    assign layer0_outputs[6852] = ~((inputs[227]) ^ (inputs[96]));
    assign layer0_outputs[6853] = ~(inputs[169]);
    assign layer0_outputs[6854] = ~(inputs[248]);
    assign layer0_outputs[6855] = (inputs[238]) | (inputs[253]);
    assign layer0_outputs[6856] = ~((inputs[203]) | (inputs[228]));
    assign layer0_outputs[6857] = (inputs[198]) & ~(inputs[116]);
    assign layer0_outputs[6858] = (inputs[22]) ^ (inputs[83]);
    assign layer0_outputs[6859] = ~((inputs[29]) | (inputs[228]));
    assign layer0_outputs[6860] = ~(inputs[67]);
    assign layer0_outputs[6861] = ~(inputs[158]) | (inputs[157]);
    assign layer0_outputs[6862] = ~(inputs[158]);
    assign layer0_outputs[6863] = ~((inputs[13]) | (inputs[4]));
    assign layer0_outputs[6864] = (inputs[238]) & ~(inputs[157]);
    assign layer0_outputs[6865] = (inputs[68]) ^ (inputs[195]);
    assign layer0_outputs[6866] = (inputs[204]) & ~(inputs[200]);
    assign layer0_outputs[6867] = (inputs[173]) & ~(inputs[199]);
    assign layer0_outputs[6868] = (inputs[95]) | (inputs[177]);
    assign layer0_outputs[6869] = inputs[1];
    assign layer0_outputs[6870] = (inputs[210]) | (inputs[51]);
    assign layer0_outputs[6871] = ~(inputs[136]) | (inputs[147]);
    assign layer0_outputs[6872] = ~((inputs[234]) | (inputs[160]));
    assign layer0_outputs[6873] = ~((inputs[18]) | (inputs[36]));
    assign layer0_outputs[6874] = ~((inputs[19]) | (inputs[51]));
    assign layer0_outputs[6875] = inputs[238];
    assign layer0_outputs[6876] = ~((inputs[46]) | (inputs[205]));
    assign layer0_outputs[6877] = (inputs[182]) & ~(inputs[40]);
    assign layer0_outputs[6878] = ~(inputs[57]);
    assign layer0_outputs[6879] = ~(inputs[216]);
    assign layer0_outputs[6880] = 1'b1;
    assign layer0_outputs[6881] = ~((inputs[94]) | (inputs[41]));
    assign layer0_outputs[6882] = inputs[84];
    assign layer0_outputs[6883] = (inputs[134]) & ~(inputs[140]);
    assign layer0_outputs[6884] = (inputs[209]) & ~(inputs[119]);
    assign layer0_outputs[6885] = ~((inputs[25]) ^ (inputs[55]));
    assign layer0_outputs[6886] = (inputs[159]) & (inputs[159]);
    assign layer0_outputs[6887] = 1'b0;
    assign layer0_outputs[6888] = ~(inputs[123]) | (inputs[46]);
    assign layer0_outputs[6889] = 1'b1;
    assign layer0_outputs[6890] = ~(inputs[91]);
    assign layer0_outputs[6891] = 1'b1;
    assign layer0_outputs[6892] = ~(inputs[217]);
    assign layer0_outputs[6893] = ~(inputs[78]) | (inputs[236]);
    assign layer0_outputs[6894] = inputs[215];
    assign layer0_outputs[6895] = (inputs[132]) & ~(inputs[172]);
    assign layer0_outputs[6896] = ~((inputs[107]) | (inputs[60]));
    assign layer0_outputs[6897] = (inputs[150]) | (inputs[70]);
    assign layer0_outputs[6898] = ~(inputs[249]);
    assign layer0_outputs[6899] = ~((inputs[224]) | (inputs[136]));
    assign layer0_outputs[6900] = ~(inputs[3]) | (inputs[233]);
    assign layer0_outputs[6901] = ~(inputs[101]) | (inputs[191]);
    assign layer0_outputs[6902] = (inputs[19]) & ~(inputs[254]);
    assign layer0_outputs[6903] = ~((inputs[100]) | (inputs[56]));
    assign layer0_outputs[6904] = (inputs[79]) | (inputs[211]);
    assign layer0_outputs[6905] = (inputs[229]) ^ (inputs[167]);
    assign layer0_outputs[6906] = ~(inputs[243]);
    assign layer0_outputs[6907] = (inputs[107]) & (inputs[92]);
    assign layer0_outputs[6908] = (inputs[23]) | (inputs[109]);
    assign layer0_outputs[6909] = inputs[197];
    assign layer0_outputs[6910] = 1'b0;
    assign layer0_outputs[6911] = ~((inputs[233]) | (inputs[226]));
    assign layer0_outputs[6912] = 1'b1;
    assign layer0_outputs[6913] = ~(inputs[55]);
    assign layer0_outputs[6914] = (inputs[179]) | (inputs[34]);
    assign layer0_outputs[6915] = ~(inputs[114]) | (inputs[74]);
    assign layer0_outputs[6916] = (inputs[176]) | (inputs[103]);
    assign layer0_outputs[6917] = ~(inputs[94]);
    assign layer0_outputs[6918] = ~(inputs[228]);
    assign layer0_outputs[6919] = ~((inputs[201]) ^ (inputs[191]));
    assign layer0_outputs[6920] = ~((inputs[202]) | (inputs[178]));
    assign layer0_outputs[6921] = (inputs[22]) & ~(inputs[158]);
    assign layer0_outputs[6922] = ~(inputs[79]);
    assign layer0_outputs[6923] = ~(inputs[28]);
    assign layer0_outputs[6924] = 1'b1;
    assign layer0_outputs[6925] = (inputs[100]) | (inputs[187]);
    assign layer0_outputs[6926] = ~(inputs[41]) | (inputs[93]);
    assign layer0_outputs[6927] = (inputs[80]) ^ (inputs[193]);
    assign layer0_outputs[6928] = ~((inputs[42]) | (inputs[27]));
    assign layer0_outputs[6929] = (inputs[134]) & (inputs[104]);
    assign layer0_outputs[6930] = ~((inputs[240]) ^ (inputs[127]));
    assign layer0_outputs[6931] = ~(inputs[129]);
    assign layer0_outputs[6932] = ~((inputs[23]) & (inputs[158]));
    assign layer0_outputs[6933] = 1'b0;
    assign layer0_outputs[6934] = (inputs[18]) | (inputs[181]);
    assign layer0_outputs[6935] = inputs[125];
    assign layer0_outputs[6936] = (inputs[69]) | (inputs[56]);
    assign layer0_outputs[6937] = ~(inputs[116]) | (inputs[245]);
    assign layer0_outputs[6938] = inputs[255];
    assign layer0_outputs[6939] = inputs[129];
    assign layer0_outputs[6940] = ~(inputs[145]);
    assign layer0_outputs[6941] = 1'b0;
    assign layer0_outputs[6942] = inputs[27];
    assign layer0_outputs[6943] = (inputs[14]) & ~(inputs[211]);
    assign layer0_outputs[6944] = ~((inputs[162]) ^ (inputs[215]));
    assign layer0_outputs[6945] = ~(inputs[54]);
    assign layer0_outputs[6946] = (inputs[207]) | (inputs[227]);
    assign layer0_outputs[6947] = ~(inputs[118]);
    assign layer0_outputs[6948] = ~(inputs[121]);
    assign layer0_outputs[6949] = (inputs[231]) & (inputs[224]);
    assign layer0_outputs[6950] = (inputs[254]) ^ (inputs[93]);
    assign layer0_outputs[6951] = ~(inputs[234]);
    assign layer0_outputs[6952] = ~(inputs[220]);
    assign layer0_outputs[6953] = (inputs[47]) | (inputs[4]);
    assign layer0_outputs[6954] = inputs[216];
    assign layer0_outputs[6955] = (inputs[34]) | (inputs[151]);
    assign layer0_outputs[6956] = (inputs[159]) | (inputs[197]);
    assign layer0_outputs[6957] = inputs[203];
    assign layer0_outputs[6958] = (inputs[210]) & ~(inputs[40]);
    assign layer0_outputs[6959] = ~(inputs[239]);
    assign layer0_outputs[6960] = ~(inputs[232]) | (inputs[6]);
    assign layer0_outputs[6961] = ~(inputs[168]);
    assign layer0_outputs[6962] = 1'b1;
    assign layer0_outputs[6963] = ~((inputs[56]) ^ (inputs[4]));
    assign layer0_outputs[6964] = ~(inputs[14]);
    assign layer0_outputs[6965] = (inputs[111]) & (inputs[55]);
    assign layer0_outputs[6966] = ~((inputs[139]) ^ (inputs[120]));
    assign layer0_outputs[6967] = ~(inputs[200]);
    assign layer0_outputs[6968] = inputs[73];
    assign layer0_outputs[6969] = ~((inputs[175]) | (inputs[204]));
    assign layer0_outputs[6970] = inputs[144];
    assign layer0_outputs[6971] = ~(inputs[196]);
    assign layer0_outputs[6972] = ~(inputs[218]);
    assign layer0_outputs[6973] = ~(inputs[151]) | (inputs[139]);
    assign layer0_outputs[6974] = ~(inputs[100]) | (inputs[88]);
    assign layer0_outputs[6975] = ~(inputs[56]) | (inputs[237]);
    assign layer0_outputs[6976] = (inputs[230]) & ~(inputs[224]);
    assign layer0_outputs[6977] = ~((inputs[236]) | (inputs[104]));
    assign layer0_outputs[6978] = (inputs[116]) & ~(inputs[169]);
    assign layer0_outputs[6979] = (inputs[101]) & (inputs[92]);
    assign layer0_outputs[6980] = ~((inputs[142]) | (inputs[85]));
    assign layer0_outputs[6981] = inputs[92];
    assign layer0_outputs[6982] = ~(inputs[39]) | (inputs[127]);
    assign layer0_outputs[6983] = (inputs[107]) ^ (inputs[73]);
    assign layer0_outputs[6984] = ~(inputs[11]) | (inputs[72]);
    assign layer0_outputs[6985] = (inputs[177]) ^ (inputs[8]);
    assign layer0_outputs[6986] = ~(inputs[213]) | (inputs[13]);
    assign layer0_outputs[6987] = ~(inputs[153]);
    assign layer0_outputs[6988] = (inputs[10]) | (inputs[97]);
    assign layer0_outputs[6989] = inputs[21];
    assign layer0_outputs[6990] = (inputs[213]) | (inputs[135]);
    assign layer0_outputs[6991] = inputs[143];
    assign layer0_outputs[6992] = (inputs[26]) ^ (inputs[32]);
    assign layer0_outputs[6993] = ~(inputs[38]);
    assign layer0_outputs[6994] = (inputs[70]) | (inputs[111]);
    assign layer0_outputs[6995] = ~((inputs[204]) | (inputs[112]));
    assign layer0_outputs[6996] = ~(inputs[231]);
    assign layer0_outputs[6997] = (inputs[211]) & ~(inputs[60]);
    assign layer0_outputs[6998] = inputs[122];
    assign layer0_outputs[6999] = (inputs[44]) ^ (inputs[196]);
    assign layer0_outputs[7000] = ~(inputs[155]);
    assign layer0_outputs[7001] = (inputs[177]) & ~(inputs[150]);
    assign layer0_outputs[7002] = ~(inputs[243]) | (inputs[107]);
    assign layer0_outputs[7003] = (inputs[208]) & ~(inputs[64]);
    assign layer0_outputs[7004] = ~((inputs[163]) ^ (inputs[196]));
    assign layer0_outputs[7005] = ~(inputs[184]);
    assign layer0_outputs[7006] = ~((inputs[244]) & (inputs[189]));
    assign layer0_outputs[7007] = ~(inputs[4]) | (inputs[65]);
    assign layer0_outputs[7008] = ~(inputs[164]);
    assign layer0_outputs[7009] = ~(inputs[107]) | (inputs[193]);
    assign layer0_outputs[7010] = ~((inputs[204]) ^ (inputs[65]));
    assign layer0_outputs[7011] = ~(inputs[47]);
    assign layer0_outputs[7012] = ~(inputs[195]) | (inputs[121]);
    assign layer0_outputs[7013] = ~(inputs[244]) | (inputs[158]);
    assign layer0_outputs[7014] = (inputs[231]) & ~(inputs[119]);
    assign layer0_outputs[7015] = inputs[253];
    assign layer0_outputs[7016] = ~((inputs[64]) & (inputs[255]));
    assign layer0_outputs[7017] = ~((inputs[194]) | (inputs[129]));
    assign layer0_outputs[7018] = ~((inputs[207]) | (inputs[187]));
    assign layer0_outputs[7019] = (inputs[50]) | (inputs[105]);
    assign layer0_outputs[7020] = ~(inputs[65]) | (inputs[245]);
    assign layer0_outputs[7021] = inputs[101];
    assign layer0_outputs[7022] = ~(inputs[125]) | (inputs[231]);
    assign layer0_outputs[7023] = 1'b1;
    assign layer0_outputs[7024] = ~(inputs[135]) | (inputs[238]);
    assign layer0_outputs[7025] = (inputs[253]) | (inputs[1]);
    assign layer0_outputs[7026] = ~(inputs[241]) | (inputs[211]);
    assign layer0_outputs[7027] = ~(inputs[106]);
    assign layer0_outputs[7028] = ~(inputs[172]);
    assign layer0_outputs[7029] = ~(inputs[76]);
    assign layer0_outputs[7030] = ~(inputs[6]) | (inputs[218]);
    assign layer0_outputs[7031] = ~(inputs[198]) | (inputs[98]);
    assign layer0_outputs[7032] = ~(inputs[188]);
    assign layer0_outputs[7033] = ~((inputs[48]) & (inputs[12]));
    assign layer0_outputs[7034] = (inputs[25]) | (inputs[225]);
    assign layer0_outputs[7035] = (inputs[116]) & ~(inputs[34]);
    assign layer0_outputs[7036] = ~(inputs[152]);
    assign layer0_outputs[7037] = (inputs[125]) & ~(inputs[110]);
    assign layer0_outputs[7038] = (inputs[15]) & (inputs[185]);
    assign layer0_outputs[7039] = inputs[93];
    assign layer0_outputs[7040] = inputs[86];
    assign layer0_outputs[7041] = ~((inputs[251]) & (inputs[19]));
    assign layer0_outputs[7042] = ~((inputs[50]) | (inputs[195]));
    assign layer0_outputs[7043] = ~(inputs[116]);
    assign layer0_outputs[7044] = ~((inputs[51]) ^ (inputs[23]));
    assign layer0_outputs[7045] = ~((inputs[87]) | (inputs[101]));
    assign layer0_outputs[7046] = (inputs[35]) ^ (inputs[147]);
    assign layer0_outputs[7047] = ~((inputs[212]) | (inputs[46]));
    assign layer0_outputs[7048] = ~(inputs[113]) | (inputs[235]);
    assign layer0_outputs[7049] = ~(inputs[241]);
    assign layer0_outputs[7050] = ~((inputs[68]) | (inputs[78]));
    assign layer0_outputs[7051] = inputs[54];
    assign layer0_outputs[7052] = (inputs[52]) | (inputs[52]);
    assign layer0_outputs[7053] = inputs[50];
    assign layer0_outputs[7054] = ~(inputs[196]) | (inputs[78]);
    assign layer0_outputs[7055] = inputs[208];
    assign layer0_outputs[7056] = (inputs[187]) & (inputs[54]);
    assign layer0_outputs[7057] = (inputs[184]) & ~(inputs[42]);
    assign layer0_outputs[7058] = (inputs[27]) ^ (inputs[168]);
    assign layer0_outputs[7059] = (inputs[65]) & (inputs[39]);
    assign layer0_outputs[7060] = (inputs[28]) & (inputs[149]);
    assign layer0_outputs[7061] = ~(inputs[148]);
    assign layer0_outputs[7062] = (inputs[97]) | (inputs[10]);
    assign layer0_outputs[7063] = (inputs[34]) & ~(inputs[196]);
    assign layer0_outputs[7064] = (inputs[27]) & ~(inputs[195]);
    assign layer0_outputs[7065] = ~(inputs[180]) | (inputs[14]);
    assign layer0_outputs[7066] = ~(inputs[229]) | (inputs[163]);
    assign layer0_outputs[7067] = ~(inputs[141]) | (inputs[50]);
    assign layer0_outputs[7068] = (inputs[166]) | (inputs[178]);
    assign layer0_outputs[7069] = ~(inputs[210]);
    assign layer0_outputs[7070] = ~(inputs[190]) | (inputs[12]);
    assign layer0_outputs[7071] = inputs[183];
    assign layer0_outputs[7072] = ~(inputs[244]) | (inputs[15]);
    assign layer0_outputs[7073] = ~(inputs[14]);
    assign layer0_outputs[7074] = ~((inputs[48]) ^ (inputs[69]));
    assign layer0_outputs[7075] = ~(inputs[119]);
    assign layer0_outputs[7076] = (inputs[140]) & ~(inputs[175]);
    assign layer0_outputs[7077] = ~(inputs[151]);
    assign layer0_outputs[7078] = (inputs[177]) & ~(inputs[239]);
    assign layer0_outputs[7079] = ~(inputs[83]);
    assign layer0_outputs[7080] = (inputs[249]) | (inputs[229]);
    assign layer0_outputs[7081] = ~((inputs[192]) ^ (inputs[206]));
    assign layer0_outputs[7082] = ~((inputs[43]) ^ (inputs[71]));
    assign layer0_outputs[7083] = (inputs[36]) | (inputs[247]);
    assign layer0_outputs[7084] = ~(inputs[224]);
    assign layer0_outputs[7085] = (inputs[3]) & ~(inputs[142]);
    assign layer0_outputs[7086] = (inputs[41]) & (inputs[60]);
    assign layer0_outputs[7087] = ~((inputs[75]) | (inputs[7]));
    assign layer0_outputs[7088] = ~(inputs[169]);
    assign layer0_outputs[7089] = (inputs[76]) ^ (inputs[159]);
    assign layer0_outputs[7090] = ~(inputs[194]);
    assign layer0_outputs[7091] = ~((inputs[97]) ^ (inputs[129]));
    assign layer0_outputs[7092] = ~((inputs[73]) | (inputs[74]));
    assign layer0_outputs[7093] = ~((inputs[87]) ^ (inputs[43]));
    assign layer0_outputs[7094] = ~((inputs[66]) | (inputs[67]));
    assign layer0_outputs[7095] = 1'b1;
    assign layer0_outputs[7096] = (inputs[47]) ^ (inputs[5]);
    assign layer0_outputs[7097] = (inputs[250]) | (inputs[144]);
    assign layer0_outputs[7098] = (inputs[43]) & ~(inputs[159]);
    assign layer0_outputs[7099] = ~(inputs[213]);
    assign layer0_outputs[7100] = inputs[170];
    assign layer0_outputs[7101] = (inputs[139]) & (inputs[45]);
    assign layer0_outputs[7102] = ~(inputs[12]);
    assign layer0_outputs[7103] = inputs[202];
    assign layer0_outputs[7104] = ~(inputs[89]);
    assign layer0_outputs[7105] = ~((inputs[145]) | (inputs[191]));
    assign layer0_outputs[7106] = ~(inputs[47]);
    assign layer0_outputs[7107] = ~((inputs[116]) | (inputs[77]));
    assign layer0_outputs[7108] = ~((inputs[70]) | (inputs[93]));
    assign layer0_outputs[7109] = ~((inputs[123]) & (inputs[251]));
    assign layer0_outputs[7110] = ~(inputs[20]);
    assign layer0_outputs[7111] = (inputs[130]) | (inputs[34]);
    assign layer0_outputs[7112] = (inputs[1]) | (inputs[116]);
    assign layer0_outputs[7113] = ~((inputs[124]) | (inputs[130]));
    assign layer0_outputs[7114] = (inputs[136]) & ~(inputs[203]);
    assign layer0_outputs[7115] = (inputs[12]) | (inputs[79]);
    assign layer0_outputs[7116] = (inputs[100]) & (inputs[116]);
    assign layer0_outputs[7117] = ~((inputs[59]) & (inputs[82]));
    assign layer0_outputs[7118] = (inputs[11]) & (inputs[5]);
    assign layer0_outputs[7119] = ~(inputs[3]);
    assign layer0_outputs[7120] = inputs[190];
    assign layer0_outputs[7121] = ~((inputs[164]) ^ (inputs[222]));
    assign layer0_outputs[7122] = (inputs[80]) & ~(inputs[212]);
    assign layer0_outputs[7123] = (inputs[12]) & ~(inputs[162]);
    assign layer0_outputs[7124] = ~(inputs[18]) | (inputs[127]);
    assign layer0_outputs[7125] = (inputs[176]) & ~(inputs[226]);
    assign layer0_outputs[7126] = ~(inputs[61]) | (inputs[16]);
    assign layer0_outputs[7127] = ~(inputs[130]);
    assign layer0_outputs[7128] = (inputs[74]) & (inputs[236]);
    assign layer0_outputs[7129] = inputs[221];
    assign layer0_outputs[7130] = ~(inputs[27]) | (inputs[200]);
    assign layer0_outputs[7131] = inputs[92];
    assign layer0_outputs[7132] = ~(inputs[145]) | (inputs[235]);
    assign layer0_outputs[7133] = (inputs[9]) ^ (inputs[219]);
    assign layer0_outputs[7134] = ~(inputs[226]);
    assign layer0_outputs[7135] = inputs[249];
    assign layer0_outputs[7136] = ~((inputs[22]) ^ (inputs[68]));
    assign layer0_outputs[7137] = (inputs[21]) | (inputs[171]);
    assign layer0_outputs[7138] = ~(inputs[157]);
    assign layer0_outputs[7139] = (inputs[85]) | (inputs[35]);
    assign layer0_outputs[7140] = ~(inputs[86]);
    assign layer0_outputs[7141] = ~(inputs[206]);
    assign layer0_outputs[7142] = ~(inputs[172]);
    assign layer0_outputs[7143] = (inputs[193]) & ~(inputs[216]);
    assign layer0_outputs[7144] = (inputs[97]) & (inputs[5]);
    assign layer0_outputs[7145] = (inputs[109]) & ~(inputs[151]);
    assign layer0_outputs[7146] = inputs[158];
    assign layer0_outputs[7147] = ~(inputs[199]);
    assign layer0_outputs[7148] = (inputs[124]) & (inputs[48]);
    assign layer0_outputs[7149] = (inputs[207]) | (inputs[232]);
    assign layer0_outputs[7150] = inputs[4];
    assign layer0_outputs[7151] = ~(inputs[202]) | (inputs[94]);
    assign layer0_outputs[7152] = ~(inputs[138]);
    assign layer0_outputs[7153] = (inputs[219]) & (inputs[201]);
    assign layer0_outputs[7154] = inputs[134];
    assign layer0_outputs[7155] = (inputs[254]) ^ (inputs[35]);
    assign layer0_outputs[7156] = ~(inputs[67]);
    assign layer0_outputs[7157] = (inputs[188]) ^ (inputs[252]);
    assign layer0_outputs[7158] = 1'b1;
    assign layer0_outputs[7159] = ~((inputs[186]) & (inputs[167]));
    assign layer0_outputs[7160] = ~((inputs[157]) | (inputs[156]));
    assign layer0_outputs[7161] = inputs[0];
    assign layer0_outputs[7162] = ~(inputs[150]) | (inputs[76]);
    assign layer0_outputs[7163] = ~(inputs[182]) | (inputs[132]);
    assign layer0_outputs[7164] = inputs[194];
    assign layer0_outputs[7165] = inputs[85];
    assign layer0_outputs[7166] = (inputs[41]) ^ (inputs[165]);
    assign layer0_outputs[7167] = (inputs[42]) & ~(inputs[24]);
    assign layer0_outputs[7168] = ~(inputs[179]);
    assign layer0_outputs[7169] = ~(inputs[206]) | (inputs[49]);
    assign layer0_outputs[7170] = (inputs[69]) & ~(inputs[32]);
    assign layer0_outputs[7171] = ~(inputs[175]);
    assign layer0_outputs[7172] = (inputs[71]) & ~(inputs[51]);
    assign layer0_outputs[7173] = ~(inputs[197]) | (inputs[31]);
    assign layer0_outputs[7174] = ~(inputs[141]) | (inputs[33]);
    assign layer0_outputs[7175] = (inputs[244]) ^ (inputs[212]);
    assign layer0_outputs[7176] = 1'b0;
    assign layer0_outputs[7177] = ~((inputs[217]) & (inputs[39]));
    assign layer0_outputs[7178] = 1'b0;
    assign layer0_outputs[7179] = inputs[54];
    assign layer0_outputs[7180] = (inputs[220]) ^ (inputs[174]);
    assign layer0_outputs[7181] = ~(inputs[187]) | (inputs[10]);
    assign layer0_outputs[7182] = ~(inputs[140]) | (inputs[108]);
    assign layer0_outputs[7183] = inputs[62];
    assign layer0_outputs[7184] = ~(inputs[123]);
    assign layer0_outputs[7185] = (inputs[131]) | (inputs[206]);
    assign layer0_outputs[7186] = (inputs[245]) ^ (inputs[143]);
    assign layer0_outputs[7187] = ~(inputs[187]);
    assign layer0_outputs[7188] = inputs[196];
    assign layer0_outputs[7189] = ~((inputs[49]) | (inputs[43]));
    assign layer0_outputs[7190] = ~(inputs[240]) | (inputs[166]);
    assign layer0_outputs[7191] = inputs[209];
    assign layer0_outputs[7192] = ~(inputs[86]);
    assign layer0_outputs[7193] = (inputs[51]) & ~(inputs[240]);
    assign layer0_outputs[7194] = ~(inputs[37]) | (inputs[194]);
    assign layer0_outputs[7195] = ~((inputs[44]) | (inputs[92]));
    assign layer0_outputs[7196] = inputs[170];
    assign layer0_outputs[7197] = (inputs[126]) ^ (inputs[123]);
    assign layer0_outputs[7198] = inputs[140];
    assign layer0_outputs[7199] = inputs[184];
    assign layer0_outputs[7200] = ~((inputs[154]) | (inputs[103]));
    assign layer0_outputs[7201] = (inputs[36]) | (inputs[79]);
    assign layer0_outputs[7202] = ~((inputs[205]) & (inputs[170]));
    assign layer0_outputs[7203] = ~(inputs[185]);
    assign layer0_outputs[7204] = (inputs[9]) & ~(inputs[197]);
    assign layer0_outputs[7205] = (inputs[231]) & (inputs[227]);
    assign layer0_outputs[7206] = (inputs[93]) | (inputs[27]);
    assign layer0_outputs[7207] = (inputs[251]) & ~(inputs[72]);
    assign layer0_outputs[7208] = ~(inputs[196]) | (inputs[161]);
    assign layer0_outputs[7209] = ~(inputs[136]) | (inputs[172]);
    assign layer0_outputs[7210] = (inputs[55]) | (inputs[109]);
    assign layer0_outputs[7211] = (inputs[148]) | (inputs[15]);
    assign layer0_outputs[7212] = 1'b0;
    assign layer0_outputs[7213] = ~(inputs[171]);
    assign layer0_outputs[7214] = ~(inputs[53]);
    assign layer0_outputs[7215] = ~((inputs[189]) ^ (inputs[187]));
    assign layer0_outputs[7216] = (inputs[4]) ^ (inputs[79]);
    assign layer0_outputs[7217] = inputs[59];
    assign layer0_outputs[7218] = ~(inputs[101]);
    assign layer0_outputs[7219] = ~(inputs[224]) | (inputs[169]);
    assign layer0_outputs[7220] = ~((inputs[65]) ^ (inputs[141]));
    assign layer0_outputs[7221] = (inputs[11]) | (inputs[12]);
    assign layer0_outputs[7222] = (inputs[148]) | (inputs[216]);
    assign layer0_outputs[7223] = ~(inputs[81]) | (inputs[139]);
    assign layer0_outputs[7224] = ~((inputs[45]) & (inputs[210]));
    assign layer0_outputs[7225] = ~((inputs[24]) ^ (inputs[147]));
    assign layer0_outputs[7226] = ~(inputs[54]);
    assign layer0_outputs[7227] = (inputs[242]) & ~(inputs[215]);
    assign layer0_outputs[7228] = ~(inputs[129]) | (inputs[140]);
    assign layer0_outputs[7229] = ~(inputs[28]) | (inputs[184]);
    assign layer0_outputs[7230] = inputs[200];
    assign layer0_outputs[7231] = (inputs[132]) ^ (inputs[51]);
    assign layer0_outputs[7232] = ~(inputs[250]);
    assign layer0_outputs[7233] = ~(inputs[109]) | (inputs[83]);
    assign layer0_outputs[7234] = ~((inputs[110]) | (inputs[33]));
    assign layer0_outputs[7235] = (inputs[17]) | (inputs[100]);
    assign layer0_outputs[7236] = (inputs[212]) & ~(inputs[221]);
    assign layer0_outputs[7237] = ~(inputs[165]);
    assign layer0_outputs[7238] = ~(inputs[172]);
    assign layer0_outputs[7239] = ~(inputs[101]) | (inputs[63]);
    assign layer0_outputs[7240] = ~((inputs[197]) ^ (inputs[213]));
    assign layer0_outputs[7241] = ~((inputs[63]) & (inputs[3]));
    assign layer0_outputs[7242] = ~(inputs[109]);
    assign layer0_outputs[7243] = ~(inputs[45]);
    assign layer0_outputs[7244] = ~(inputs[180]);
    assign layer0_outputs[7245] = ~(inputs[64]);
    assign layer0_outputs[7246] = (inputs[152]) | (inputs[175]);
    assign layer0_outputs[7247] = (inputs[88]) ^ (inputs[119]);
    assign layer0_outputs[7248] = inputs[171];
    assign layer0_outputs[7249] = (inputs[204]) & (inputs[219]);
    assign layer0_outputs[7250] = (inputs[8]) | (inputs[154]);
    assign layer0_outputs[7251] = ~((inputs[168]) ^ (inputs[62]));
    assign layer0_outputs[7252] = ~((inputs[48]) & (inputs[0]));
    assign layer0_outputs[7253] = ~(inputs[25]);
    assign layer0_outputs[7254] = ~(inputs[26]) | (inputs[17]);
    assign layer0_outputs[7255] = (inputs[183]) & ~(inputs[172]);
    assign layer0_outputs[7256] = ~(inputs[135]) | (inputs[76]);
    assign layer0_outputs[7257] = (inputs[71]) | (inputs[223]);
    assign layer0_outputs[7258] = (inputs[18]) | (inputs[16]);
    assign layer0_outputs[7259] = ~(inputs[121]) | (inputs[20]);
    assign layer0_outputs[7260] = (inputs[190]) ^ (inputs[209]);
    assign layer0_outputs[7261] = inputs[106];
    assign layer0_outputs[7262] = ~(inputs[12]) | (inputs[176]);
    assign layer0_outputs[7263] = (inputs[2]) & (inputs[254]);
    assign layer0_outputs[7264] = (inputs[137]) & ~(inputs[95]);
    assign layer0_outputs[7265] = inputs[0];
    assign layer0_outputs[7266] = ~(inputs[67]);
    assign layer0_outputs[7267] = (inputs[7]) & ~(inputs[217]);
    assign layer0_outputs[7268] = inputs[118];
    assign layer0_outputs[7269] = ~(inputs[162]);
    assign layer0_outputs[7270] = ~(inputs[68]);
    assign layer0_outputs[7271] = (inputs[81]) | (inputs[143]);
    assign layer0_outputs[7272] = ~(inputs[102]) | (inputs[176]);
    assign layer0_outputs[7273] = inputs[110];
    assign layer0_outputs[7274] = inputs[22];
    assign layer0_outputs[7275] = (inputs[19]) & ~(inputs[211]);
    assign layer0_outputs[7276] = (inputs[96]) ^ (inputs[53]);
    assign layer0_outputs[7277] = (inputs[92]) | (inputs[53]);
    assign layer0_outputs[7278] = 1'b1;
    assign layer0_outputs[7279] = (inputs[161]) ^ (inputs[8]);
    assign layer0_outputs[7280] = (inputs[27]) & ~(inputs[61]);
    assign layer0_outputs[7281] = (inputs[250]) & ~(inputs[238]);
    assign layer0_outputs[7282] = ~(inputs[132]);
    assign layer0_outputs[7283] = ~(inputs[196]) | (inputs[3]);
    assign layer0_outputs[7284] = ~(inputs[147]) | (inputs[66]);
    assign layer0_outputs[7285] = ~((inputs[223]) ^ (inputs[123]));
    assign layer0_outputs[7286] = ~(inputs[184]);
    assign layer0_outputs[7287] = ~((inputs[199]) & (inputs[201]));
    assign layer0_outputs[7288] = ~(inputs[91]) | (inputs[160]);
    assign layer0_outputs[7289] = ~(inputs[11]) | (inputs[117]);
    assign layer0_outputs[7290] = ~(inputs[193]);
    assign layer0_outputs[7291] = ~((inputs[48]) | (inputs[14]));
    assign layer0_outputs[7292] = ~(inputs[18]);
    assign layer0_outputs[7293] = (inputs[96]) | (inputs[168]);
    assign layer0_outputs[7294] = ~((inputs[122]) | (inputs[137]));
    assign layer0_outputs[7295] = inputs[138];
    assign layer0_outputs[7296] = inputs[211];
    assign layer0_outputs[7297] = ~(inputs[135]) | (inputs[108]);
    assign layer0_outputs[7298] = (inputs[254]) & ~(inputs[36]);
    assign layer0_outputs[7299] = inputs[106];
    assign layer0_outputs[7300] = ~((inputs[110]) & (inputs[203]));
    assign layer0_outputs[7301] = (inputs[72]) & ~(inputs[93]);
    assign layer0_outputs[7302] = (inputs[8]) & ~(inputs[3]);
    assign layer0_outputs[7303] = (inputs[142]) ^ (inputs[19]);
    assign layer0_outputs[7304] = ~((inputs[216]) ^ (inputs[248]));
    assign layer0_outputs[7305] = 1'b0;
    assign layer0_outputs[7306] = ~(inputs[92]);
    assign layer0_outputs[7307] = (inputs[128]) | (inputs[53]);
    assign layer0_outputs[7308] = ~((inputs[14]) & (inputs[199]));
    assign layer0_outputs[7309] = ~(inputs[228]);
    assign layer0_outputs[7310] = ~(inputs[214]);
    assign layer0_outputs[7311] = inputs[71];
    assign layer0_outputs[7312] = ~((inputs[14]) | (inputs[102]));
    assign layer0_outputs[7313] = ~((inputs[34]) ^ (inputs[19]));
    assign layer0_outputs[7314] = ~(inputs[91]) | (inputs[160]);
    assign layer0_outputs[7315] = inputs[162];
    assign layer0_outputs[7316] = (inputs[182]) & ~(inputs[133]);
    assign layer0_outputs[7317] = (inputs[79]) ^ (inputs[174]);
    assign layer0_outputs[7318] = (inputs[39]) ^ (inputs[28]);
    assign layer0_outputs[7319] = ~(inputs[158]);
    assign layer0_outputs[7320] = inputs[206];
    assign layer0_outputs[7321] = ~(inputs[244]) | (inputs[95]);
    assign layer0_outputs[7322] = ~((inputs[59]) | (inputs[145]));
    assign layer0_outputs[7323] = ~((inputs[61]) | (inputs[60]));
    assign layer0_outputs[7324] = inputs[86];
    assign layer0_outputs[7325] = ~(inputs[70]);
    assign layer0_outputs[7326] = (inputs[199]) & ~(inputs[46]);
    assign layer0_outputs[7327] = 1'b0;
    assign layer0_outputs[7328] = inputs[195];
    assign layer0_outputs[7329] = (inputs[91]) | (inputs[89]);
    assign layer0_outputs[7330] = (inputs[66]) & ~(inputs[54]);
    assign layer0_outputs[7331] = inputs[165];
    assign layer0_outputs[7332] = ~(inputs[141]) | (inputs[255]);
    assign layer0_outputs[7333] = ~(inputs[244]);
    assign layer0_outputs[7334] = ~(inputs[107]);
    assign layer0_outputs[7335] = (inputs[164]) ^ (inputs[228]);
    assign layer0_outputs[7336] = inputs[248];
    assign layer0_outputs[7337] = ~(inputs[37]) | (inputs[54]);
    assign layer0_outputs[7338] = (inputs[172]) ^ (inputs[5]);
    assign layer0_outputs[7339] = ~(inputs[21]) | (inputs[85]);
    assign layer0_outputs[7340] = inputs[233];
    assign layer0_outputs[7341] = ~((inputs[0]) | (inputs[22]));
    assign layer0_outputs[7342] = inputs[108];
    assign layer0_outputs[7343] = ~((inputs[245]) | (inputs[29]));
    assign layer0_outputs[7344] = (inputs[153]) & ~(inputs[58]);
    assign layer0_outputs[7345] = 1'b0;
    assign layer0_outputs[7346] = ~((inputs[88]) | (inputs[152]));
    assign layer0_outputs[7347] = ~(inputs[12]) | (inputs[223]);
    assign layer0_outputs[7348] = (inputs[68]) ^ (inputs[65]);
    assign layer0_outputs[7349] = inputs[72];
    assign layer0_outputs[7350] = ~(inputs[40]);
    assign layer0_outputs[7351] = ~(inputs[188]);
    assign layer0_outputs[7352] = ~((inputs[209]) | (inputs[149]));
    assign layer0_outputs[7353] = ~(inputs[5]) | (inputs[54]);
    assign layer0_outputs[7354] = ~(inputs[179]) | (inputs[35]);
    assign layer0_outputs[7355] = ~(inputs[162]);
    assign layer0_outputs[7356] = (inputs[193]) & ~(inputs[112]);
    assign layer0_outputs[7357] = ~((inputs[44]) & (inputs[39]));
    assign layer0_outputs[7358] = (inputs[161]) ^ (inputs[141]);
    assign layer0_outputs[7359] = ~((inputs[8]) | (inputs[154]));
    assign layer0_outputs[7360] = (inputs[14]) & ~(inputs[78]);
    assign layer0_outputs[7361] = ~((inputs[155]) ^ (inputs[146]));
    assign layer0_outputs[7362] = ~((inputs[69]) & (inputs[5]));
    assign layer0_outputs[7363] = ~((inputs[17]) | (inputs[230]));
    assign layer0_outputs[7364] = inputs[138];
    assign layer0_outputs[7365] = (inputs[105]) | (inputs[97]);
    assign layer0_outputs[7366] = ~((inputs[99]) & (inputs[193]));
    assign layer0_outputs[7367] = ~(inputs[152]) | (inputs[247]);
    assign layer0_outputs[7368] = (inputs[147]) & ~(inputs[217]);
    assign layer0_outputs[7369] = (inputs[121]) & ~(inputs[132]);
    assign layer0_outputs[7370] = ~((inputs[132]) ^ (inputs[98]));
    assign layer0_outputs[7371] = ~((inputs[214]) ^ (inputs[206]));
    assign layer0_outputs[7372] = ~(inputs[182]) | (inputs[63]);
    assign layer0_outputs[7373] = ~((inputs[12]) ^ (inputs[17]));
    assign layer0_outputs[7374] = inputs[144];
    assign layer0_outputs[7375] = 1'b1;
    assign layer0_outputs[7376] = (inputs[171]) | (inputs[186]);
    assign layer0_outputs[7377] = ~(inputs[164]);
    assign layer0_outputs[7378] = (inputs[236]) | (inputs[243]);
    assign layer0_outputs[7379] = inputs[22];
    assign layer0_outputs[7380] = ~((inputs[181]) | (inputs[148]));
    assign layer0_outputs[7381] = ~(inputs[142]);
    assign layer0_outputs[7382] = inputs[112];
    assign layer0_outputs[7383] = ~((inputs[99]) | (inputs[187]));
    assign layer0_outputs[7384] = (inputs[30]) & (inputs[132]);
    assign layer0_outputs[7385] = inputs[179];
    assign layer0_outputs[7386] = ~((inputs[222]) ^ (inputs[235]));
    assign layer0_outputs[7387] = (inputs[76]) & (inputs[190]);
    assign layer0_outputs[7388] = (inputs[21]) & ~(inputs[77]);
    assign layer0_outputs[7389] = ~(inputs[152]) | (inputs[45]);
    assign layer0_outputs[7390] = (inputs[248]) & ~(inputs[30]);
    assign layer0_outputs[7391] = ~(inputs[121]) | (inputs[149]);
    assign layer0_outputs[7392] = (inputs[74]) ^ (inputs[24]);
    assign layer0_outputs[7393] = (inputs[142]) | (inputs[249]);
    assign layer0_outputs[7394] = ~(inputs[223]);
    assign layer0_outputs[7395] = ~(inputs[42]) | (inputs[98]);
    assign layer0_outputs[7396] = 1'b1;
    assign layer0_outputs[7397] = inputs[52];
    assign layer0_outputs[7398] = ~((inputs[119]) ^ (inputs[160]));
    assign layer0_outputs[7399] = ~((inputs[8]) | (inputs[66]));
    assign layer0_outputs[7400] = inputs[113];
    assign layer0_outputs[7401] = inputs[215];
    assign layer0_outputs[7402] = (inputs[53]) & ~(inputs[241]);
    assign layer0_outputs[7403] = ~(inputs[3]) | (inputs[32]);
    assign layer0_outputs[7404] = ~((inputs[111]) | (inputs[124]));
    assign layer0_outputs[7405] = 1'b0;
    assign layer0_outputs[7406] = (inputs[230]) | (inputs[51]);
    assign layer0_outputs[7407] = ~((inputs[115]) | (inputs[43]));
    assign layer0_outputs[7408] = ~(inputs[103]) | (inputs[181]);
    assign layer0_outputs[7409] = inputs[113];
    assign layer0_outputs[7410] = ~(inputs[119]) | (inputs[230]);
    assign layer0_outputs[7411] = inputs[54];
    assign layer0_outputs[7412] = 1'b0;
    assign layer0_outputs[7413] = inputs[72];
    assign layer0_outputs[7414] = inputs[21];
    assign layer0_outputs[7415] = ~((inputs[171]) & (inputs[255]));
    assign layer0_outputs[7416] = ~(inputs[115]) | (inputs[104]);
    assign layer0_outputs[7417] = ~(inputs[228]);
    assign layer0_outputs[7418] = ~((inputs[211]) ^ (inputs[115]));
    assign layer0_outputs[7419] = (inputs[99]) & ~(inputs[201]);
    assign layer0_outputs[7420] = inputs[105];
    assign layer0_outputs[7421] = ~((inputs[146]) | (inputs[2]));
    assign layer0_outputs[7422] = inputs[181];
    assign layer0_outputs[7423] = inputs[62];
    assign layer0_outputs[7424] = ~(inputs[11]);
    assign layer0_outputs[7425] = ~(inputs[24]);
    assign layer0_outputs[7426] = (inputs[130]) | (inputs[30]);
    assign layer0_outputs[7427] = ~((inputs[234]) | (inputs[104]));
    assign layer0_outputs[7428] = ~(inputs[70]) | (inputs[240]);
    assign layer0_outputs[7429] = inputs[134];
    assign layer0_outputs[7430] = ~((inputs[208]) | (inputs[172]));
    assign layer0_outputs[7431] = ~(inputs[86]);
    assign layer0_outputs[7432] = ~(inputs[249]) | (inputs[84]);
    assign layer0_outputs[7433] = ~(inputs[253]);
    assign layer0_outputs[7434] = 1'b1;
    assign layer0_outputs[7435] = ~(inputs[57]);
    assign layer0_outputs[7436] = (inputs[69]) | (inputs[181]);
    assign layer0_outputs[7437] = inputs[42];
    assign layer0_outputs[7438] = (inputs[182]) & ~(inputs[168]);
    assign layer0_outputs[7439] = ~((inputs[105]) ^ (inputs[167]));
    assign layer0_outputs[7440] = ~(inputs[237]);
    assign layer0_outputs[7441] = 1'b1;
    assign layer0_outputs[7442] = (inputs[57]) ^ (inputs[252]);
    assign layer0_outputs[7443] = inputs[210];
    assign layer0_outputs[7444] = 1'b1;
    assign layer0_outputs[7445] = ~(inputs[235]) | (inputs[114]);
    assign layer0_outputs[7446] = ~((inputs[180]) | (inputs[170]));
    assign layer0_outputs[7447] = ~(inputs[99]);
    assign layer0_outputs[7448] = (inputs[184]) | (inputs[84]);
    assign layer0_outputs[7449] = inputs[45];
    assign layer0_outputs[7450] = (inputs[207]) | (inputs[20]);
    assign layer0_outputs[7451] = inputs[247];
    assign layer0_outputs[7452] = inputs[171];
    assign layer0_outputs[7453] = (inputs[180]) ^ (inputs[182]);
    assign layer0_outputs[7454] = ~(inputs[121]);
    assign layer0_outputs[7455] = 1'b1;
    assign layer0_outputs[7456] = ~(inputs[247]) | (inputs[57]);
    assign layer0_outputs[7457] = (inputs[124]) & (inputs[92]);
    assign layer0_outputs[7458] = ~(inputs[200]) | (inputs[26]);
    assign layer0_outputs[7459] = (inputs[73]) ^ (inputs[45]);
    assign layer0_outputs[7460] = ~(inputs[79]) | (inputs[202]);
    assign layer0_outputs[7461] = ~((inputs[172]) | (inputs[217]));
    assign layer0_outputs[7462] = ~(inputs[152]);
    assign layer0_outputs[7463] = (inputs[227]) | (inputs[96]);
    assign layer0_outputs[7464] = ~((inputs[58]) | (inputs[153]));
    assign layer0_outputs[7465] = (inputs[91]) & ~(inputs[195]);
    assign layer0_outputs[7466] = ~(inputs[234]) | (inputs[112]);
    assign layer0_outputs[7467] = ~((inputs[206]) | (inputs[251]));
    assign layer0_outputs[7468] = ~(inputs[122]);
    assign layer0_outputs[7469] = inputs[58];
    assign layer0_outputs[7470] = (inputs[208]) & ~(inputs[113]);
    assign layer0_outputs[7471] = inputs[174];
    assign layer0_outputs[7472] = inputs[199];
    assign layer0_outputs[7473] = 1'b0;
    assign layer0_outputs[7474] = (inputs[191]) ^ (inputs[172]);
    assign layer0_outputs[7475] = ~(inputs[195]);
    assign layer0_outputs[7476] = (inputs[152]) & ~(inputs[234]);
    assign layer0_outputs[7477] = ~((inputs[227]) | (inputs[19]));
    assign layer0_outputs[7478] = ~((inputs[72]) | (inputs[143]));
    assign layer0_outputs[7479] = (inputs[124]) | (inputs[37]);
    assign layer0_outputs[7480] = (inputs[174]) ^ (inputs[126]);
    assign layer0_outputs[7481] = ~(inputs[35]);
    assign layer0_outputs[7482] = ~(inputs[112]) | (inputs[232]);
    assign layer0_outputs[7483] = (inputs[125]) | (inputs[156]);
    assign layer0_outputs[7484] = ~(inputs[189]);
    assign layer0_outputs[7485] = ~(inputs[197]);
    assign layer0_outputs[7486] = ~(inputs[27]);
    assign layer0_outputs[7487] = (inputs[60]) & ~(inputs[236]);
    assign layer0_outputs[7488] = (inputs[190]) | (inputs[141]);
    assign layer0_outputs[7489] = ~((inputs[209]) ^ (inputs[173]));
    assign layer0_outputs[7490] = (inputs[88]) & ~(inputs[3]);
    assign layer0_outputs[7491] = ~((inputs[225]) | (inputs[15]));
    assign layer0_outputs[7492] = (inputs[11]) & ~(inputs[239]);
    assign layer0_outputs[7493] = inputs[169];
    assign layer0_outputs[7494] = (inputs[229]) ^ (inputs[171]);
    assign layer0_outputs[7495] = 1'b0;
    assign layer0_outputs[7496] = ~((inputs[17]) | (inputs[196]));
    assign layer0_outputs[7497] = ~(inputs[127]);
    assign layer0_outputs[7498] = ~(inputs[126]);
    assign layer0_outputs[7499] = ~(inputs[246]);
    assign layer0_outputs[7500] = (inputs[189]) | (inputs[205]);
    assign layer0_outputs[7501] = (inputs[193]) & ~(inputs[169]);
    assign layer0_outputs[7502] = ~(inputs[74]);
    assign layer0_outputs[7503] = (inputs[230]) & ~(inputs[152]);
    assign layer0_outputs[7504] = ~((inputs[80]) ^ (inputs[70]));
    assign layer0_outputs[7505] = ~(inputs[245]);
    assign layer0_outputs[7506] = (inputs[171]) & (inputs[214]);
    assign layer0_outputs[7507] = ~((inputs[95]) ^ (inputs[104]));
    assign layer0_outputs[7508] = inputs[92];
    assign layer0_outputs[7509] = (inputs[126]) | (inputs[13]);
    assign layer0_outputs[7510] = ~(inputs[136]) | (inputs[64]);
    assign layer0_outputs[7511] = 1'b0;
    assign layer0_outputs[7512] = (inputs[133]) & ~(inputs[190]);
    assign layer0_outputs[7513] = ~((inputs[51]) ^ (inputs[199]));
    assign layer0_outputs[7514] = (inputs[83]) | (inputs[112]);
    assign layer0_outputs[7515] = (inputs[126]) | (inputs[181]);
    assign layer0_outputs[7516] = inputs[37];
    assign layer0_outputs[7517] = ~(inputs[95]);
    assign layer0_outputs[7518] = inputs[217];
    assign layer0_outputs[7519] = ~((inputs[74]) | (inputs[129]));
    assign layer0_outputs[7520] = ~((inputs[57]) & (inputs[53]));
    assign layer0_outputs[7521] = inputs[81];
    assign layer0_outputs[7522] = ~(inputs[183]) | (inputs[207]);
    assign layer0_outputs[7523] = ~(inputs[38]) | (inputs[201]);
    assign layer0_outputs[7524] = (inputs[100]) & ~(inputs[80]);
    assign layer0_outputs[7525] = (inputs[49]) & ~(inputs[209]);
    assign layer0_outputs[7526] = (inputs[178]) & ~(inputs[31]);
    assign layer0_outputs[7527] = ~(inputs[138]);
    assign layer0_outputs[7528] = (inputs[195]) ^ (inputs[0]);
    assign layer0_outputs[7529] = (inputs[255]) | (inputs[49]);
    assign layer0_outputs[7530] = ~(inputs[238]);
    assign layer0_outputs[7531] = ~((inputs[86]) ^ (inputs[19]));
    assign layer0_outputs[7532] = ~((inputs[26]) | (inputs[92]));
    assign layer0_outputs[7533] = ~(inputs[89]) | (inputs[248]);
    assign layer0_outputs[7534] = (inputs[188]) ^ (inputs[179]);
    assign layer0_outputs[7535] = ~((inputs[192]) | (inputs[95]));
    assign layer0_outputs[7536] = 1'b0;
    assign layer0_outputs[7537] = ~((inputs[50]) | (inputs[79]));
    assign layer0_outputs[7538] = (inputs[88]) & (inputs[61]);
    assign layer0_outputs[7539] = inputs[242];
    assign layer0_outputs[7540] = (inputs[141]) | (inputs[97]);
    assign layer0_outputs[7541] = inputs[218];
    assign layer0_outputs[7542] = inputs[85];
    assign layer0_outputs[7543] = ~((inputs[114]) | (inputs[102]));
    assign layer0_outputs[7544] = ~(inputs[191]);
    assign layer0_outputs[7545] = ~((inputs[192]) & (inputs[132]));
    assign layer0_outputs[7546] = (inputs[187]) & ~(inputs[14]);
    assign layer0_outputs[7547] = 1'b1;
    assign layer0_outputs[7548] = (inputs[112]) & ~(inputs[238]);
    assign layer0_outputs[7549] = ~(inputs[73]);
    assign layer0_outputs[7550] = ~((inputs[149]) ^ (inputs[221]));
    assign layer0_outputs[7551] = (inputs[139]) | (inputs[106]);
    assign layer0_outputs[7552] = (inputs[75]) & ~(inputs[81]);
    assign layer0_outputs[7553] = inputs[201];
    assign layer0_outputs[7554] = ~(inputs[87]) | (inputs[13]);
    assign layer0_outputs[7555] = (inputs[17]) & ~(inputs[3]);
    assign layer0_outputs[7556] = (inputs[158]) ^ (inputs[39]);
    assign layer0_outputs[7557] = (inputs[207]) ^ (inputs[255]);
    assign layer0_outputs[7558] = ~(inputs[9]);
    assign layer0_outputs[7559] = ~(inputs[107]) | (inputs[40]);
    assign layer0_outputs[7560] = (inputs[186]) & ~(inputs[102]);
    assign layer0_outputs[7561] = ~((inputs[214]) | (inputs[183]));
    assign layer0_outputs[7562] = ~(inputs[3]);
    assign layer0_outputs[7563] = (inputs[129]) | (inputs[156]);
    assign layer0_outputs[7564] = (inputs[161]) | (inputs[175]);
    assign layer0_outputs[7565] = ~((inputs[129]) | (inputs[149]));
    assign layer0_outputs[7566] = ~(inputs[76]);
    assign layer0_outputs[7567] = 1'b0;
    assign layer0_outputs[7568] = (inputs[251]) & (inputs[139]);
    assign layer0_outputs[7569] = ~(inputs[34]);
    assign layer0_outputs[7570] = (inputs[183]) ^ (inputs[230]);
    assign layer0_outputs[7571] = inputs[213];
    assign layer0_outputs[7572] = 1'b0;
    assign layer0_outputs[7573] = (inputs[19]) ^ (inputs[3]);
    assign layer0_outputs[7574] = ~((inputs[31]) | (inputs[122]));
    assign layer0_outputs[7575] = ~((inputs[66]) ^ (inputs[91]));
    assign layer0_outputs[7576] = ~(inputs[82]) | (inputs[240]);
    assign layer0_outputs[7577] = (inputs[202]) ^ (inputs[111]);
    assign layer0_outputs[7578] = ~(inputs[138]);
    assign layer0_outputs[7579] = (inputs[120]) & ~(inputs[155]);
    assign layer0_outputs[7580] = (inputs[99]) | (inputs[46]);
    assign layer0_outputs[7581] = ~((inputs[252]) ^ (inputs[129]));
    assign layer0_outputs[7582] = (inputs[253]) | (inputs[61]);
    assign layer0_outputs[7583] = inputs[38];
    assign layer0_outputs[7584] = (inputs[179]) | (inputs[111]);
    assign layer0_outputs[7585] = ~(inputs[71]) | (inputs[224]);
    assign layer0_outputs[7586] = inputs[177];
    assign layer0_outputs[7587] = ~(inputs[51]);
    assign layer0_outputs[7588] = ~((inputs[44]) | (inputs[84]));
    assign layer0_outputs[7589] = inputs[228];
    assign layer0_outputs[7590] = ~((inputs[138]) ^ (inputs[74]));
    assign layer0_outputs[7591] = (inputs[89]) ^ (inputs[112]);
    assign layer0_outputs[7592] = (inputs[32]) ^ (inputs[128]);
    assign layer0_outputs[7593] = ~(inputs[127]);
    assign layer0_outputs[7594] = (inputs[158]) & ~(inputs[126]);
    assign layer0_outputs[7595] = ~((inputs[167]) | (inputs[111]));
    assign layer0_outputs[7596] = ~((inputs[166]) | (inputs[33]));
    assign layer0_outputs[7597] = ~(inputs[132]) | (inputs[190]);
    assign layer0_outputs[7598] = ~(inputs[146]);
    assign layer0_outputs[7599] = ~((inputs[214]) | (inputs[19]));
    assign layer0_outputs[7600] = ~((inputs[128]) | (inputs[58]));
    assign layer0_outputs[7601] = (inputs[226]) ^ (inputs[232]);
    assign layer0_outputs[7602] = (inputs[233]) | (inputs[26]);
    assign layer0_outputs[7603] = (inputs[203]) & ~(inputs[42]);
    assign layer0_outputs[7604] = (inputs[107]) & ~(inputs[153]);
    assign layer0_outputs[7605] = (inputs[197]) | (inputs[76]);
    assign layer0_outputs[7606] = ~(inputs[101]) | (inputs[160]);
    assign layer0_outputs[7607] = (inputs[134]) & ~(inputs[7]);
    assign layer0_outputs[7608] = ~(inputs[105]);
    assign layer0_outputs[7609] = (inputs[235]) ^ (inputs[250]);
    assign layer0_outputs[7610] = ~(inputs[90]) | (inputs[188]);
    assign layer0_outputs[7611] = ~(inputs[156]) | (inputs[65]);
    assign layer0_outputs[7612] = ~((inputs[83]) ^ (inputs[82]));
    assign layer0_outputs[7613] = ~(inputs[29]) | (inputs[50]);
    assign layer0_outputs[7614] = inputs[34];
    assign layer0_outputs[7615] = ~(inputs[8]);
    assign layer0_outputs[7616] = (inputs[158]) & (inputs[218]);
    assign layer0_outputs[7617] = ~(inputs[107]);
    assign layer0_outputs[7618] = (inputs[107]) | (inputs[74]);
    assign layer0_outputs[7619] = 1'b1;
    assign layer0_outputs[7620] = ~(inputs[70]);
    assign layer0_outputs[7621] = ~(inputs[178]);
    assign layer0_outputs[7622] = (inputs[43]) | (inputs[218]);
    assign layer0_outputs[7623] = ~((inputs[242]) & (inputs[235]));
    assign layer0_outputs[7624] = inputs[202];
    assign layer0_outputs[7625] = ~((inputs[65]) ^ (inputs[104]));
    assign layer0_outputs[7626] = ~(inputs[19]) | (inputs[178]);
    assign layer0_outputs[7627] = inputs[202];
    assign layer0_outputs[7628] = 1'b0;
    assign layer0_outputs[7629] = (inputs[240]) & ~(inputs[177]);
    assign layer0_outputs[7630] = inputs[85];
    assign layer0_outputs[7631] = ~((inputs[118]) | (inputs[164]));
    assign layer0_outputs[7632] = ~(inputs[74]) | (inputs[167]);
    assign layer0_outputs[7633] = ~(inputs[68]);
    assign layer0_outputs[7634] = ~((inputs[156]) ^ (inputs[122]));
    assign layer0_outputs[7635] = ~(inputs[60]);
    assign layer0_outputs[7636] = (inputs[236]) | (inputs[161]);
    assign layer0_outputs[7637] = (inputs[172]) | (inputs[217]);
    assign layer0_outputs[7638] = ~(inputs[121]);
    assign layer0_outputs[7639] = (inputs[12]) & ~(inputs[61]);
    assign layer0_outputs[7640] = 1'b1;
    assign layer0_outputs[7641] = ~((inputs[43]) | (inputs[106]));
    assign layer0_outputs[7642] = 1'b1;
    assign layer0_outputs[7643] = ~(inputs[134]);
    assign layer0_outputs[7644] = (inputs[224]) | (inputs[89]);
    assign layer0_outputs[7645] = (inputs[21]) & ~(inputs[68]);
    assign layer0_outputs[7646] = (inputs[124]) ^ (inputs[35]);
    assign layer0_outputs[7647] = ~((inputs[8]) ^ (inputs[0]));
    assign layer0_outputs[7648] = ~((inputs[124]) | (inputs[101]));
    assign layer0_outputs[7649] = (inputs[9]) & (inputs[75]);
    assign layer0_outputs[7650] = ~(inputs[68]) | (inputs[231]);
    assign layer0_outputs[7651] = (inputs[82]) & ~(inputs[233]);
    assign layer0_outputs[7652] = ~((inputs[254]) | (inputs[190]));
    assign layer0_outputs[7653] = inputs[85];
    assign layer0_outputs[7654] = ~(inputs[68]);
    assign layer0_outputs[7655] = (inputs[133]) & ~(inputs[188]);
    assign layer0_outputs[7656] = 1'b0;
    assign layer0_outputs[7657] = ~((inputs[141]) | (inputs[147]));
    assign layer0_outputs[7658] = (inputs[180]) | (inputs[224]);
    assign layer0_outputs[7659] = inputs[63];
    assign layer0_outputs[7660] = ~((inputs[1]) ^ (inputs[224]));
    assign layer0_outputs[7661] = ~((inputs[247]) | (inputs[87]));
    assign layer0_outputs[7662] = ~((inputs[77]) ^ (inputs[28]));
    assign layer0_outputs[7663] = (inputs[57]) ^ (inputs[0]);
    assign layer0_outputs[7664] = (inputs[153]) & (inputs[135]);
    assign layer0_outputs[7665] = ~(inputs[142]);
    assign layer0_outputs[7666] = ~(inputs[250]);
    assign layer0_outputs[7667] = ~(inputs[177]);
    assign layer0_outputs[7668] = ~(inputs[120]) | (inputs[28]);
    assign layer0_outputs[7669] = 1'b0;
    assign layer0_outputs[7670] = (inputs[118]) & ~(inputs[178]);
    assign layer0_outputs[7671] = (inputs[253]) | (inputs[225]);
    assign layer0_outputs[7672] = ~((inputs[180]) ^ (inputs[15]));
    assign layer0_outputs[7673] = inputs[10];
    assign layer0_outputs[7674] = (inputs[126]) & ~(inputs[147]);
    assign layer0_outputs[7675] = inputs[152];
    assign layer0_outputs[7676] = ~(inputs[96]);
    assign layer0_outputs[7677] = (inputs[60]) | (inputs[129]);
    assign layer0_outputs[7678] = ~((inputs[138]) ^ (inputs[109]));
    assign layer0_outputs[7679] = inputs[120];
    assign layer0_outputs[7680] = ~(inputs[220]);
    assign layer0_outputs[7681] = ~((inputs[171]) & (inputs[164]));
    assign layer0_outputs[7682] = (inputs[174]) | (inputs[160]);
    assign layer0_outputs[7683] = ~(inputs[52]) | (inputs[33]);
    assign layer0_outputs[7684] = (inputs[36]) & ~(inputs[1]);
    assign layer0_outputs[7685] = inputs[138];
    assign layer0_outputs[7686] = inputs[23];
    assign layer0_outputs[7687] = ~(inputs[205]) | (inputs[250]);
    assign layer0_outputs[7688] = (inputs[137]) & (inputs[97]);
    assign layer0_outputs[7689] = (inputs[231]) & (inputs[27]);
    assign layer0_outputs[7690] = ~(inputs[106]) | (inputs[58]);
    assign layer0_outputs[7691] = inputs[228];
    assign layer0_outputs[7692] = ~(inputs[38]);
    assign layer0_outputs[7693] = inputs[237];
    assign layer0_outputs[7694] = (inputs[117]) | (inputs[86]);
    assign layer0_outputs[7695] = (inputs[245]) & ~(inputs[34]);
    assign layer0_outputs[7696] = (inputs[48]) & ~(inputs[49]);
    assign layer0_outputs[7697] = inputs[230];
    assign layer0_outputs[7698] = ~(inputs[93]);
    assign layer0_outputs[7699] = (inputs[146]) & ~(inputs[3]);
    assign layer0_outputs[7700] = ~(inputs[90]);
    assign layer0_outputs[7701] = (inputs[138]) & ~(inputs[103]);
    assign layer0_outputs[7702] = (inputs[6]) & ~(inputs[143]);
    assign layer0_outputs[7703] = (inputs[219]) | (inputs[226]);
    assign layer0_outputs[7704] = ~((inputs[62]) & (inputs[62]));
    assign layer0_outputs[7705] = (inputs[196]) | (inputs[253]);
    assign layer0_outputs[7706] = (inputs[191]) | (inputs[166]);
    assign layer0_outputs[7707] = ~(inputs[155]);
    assign layer0_outputs[7708] = inputs[154];
    assign layer0_outputs[7709] = ~(inputs[24]);
    assign layer0_outputs[7710] = ~(inputs[88]) | (inputs[38]);
    assign layer0_outputs[7711] = ~(inputs[48]);
    assign layer0_outputs[7712] = ~((inputs[52]) ^ (inputs[176]));
    assign layer0_outputs[7713] = (inputs[235]) | (inputs[223]);
    assign layer0_outputs[7714] = ~((inputs[113]) ^ (inputs[57]));
    assign layer0_outputs[7715] = inputs[162];
    assign layer0_outputs[7716] = ~(inputs[112]);
    assign layer0_outputs[7717] = ~(inputs[126]);
    assign layer0_outputs[7718] = inputs[169];
    assign layer0_outputs[7719] = ~(inputs[231]);
    assign layer0_outputs[7720] = 1'b0;
    assign layer0_outputs[7721] = ~(inputs[64]);
    assign layer0_outputs[7722] = ~(inputs[251]);
    assign layer0_outputs[7723] = ~(inputs[127]);
    assign layer0_outputs[7724] = inputs[94];
    assign layer0_outputs[7725] = (inputs[103]) ^ (inputs[147]);
    assign layer0_outputs[7726] = ~((inputs[16]) | (inputs[60]));
    assign layer0_outputs[7727] = (inputs[16]) & ~(inputs[155]);
    assign layer0_outputs[7728] = ~(inputs[135]) | (inputs[160]);
    assign layer0_outputs[7729] = inputs[110];
    assign layer0_outputs[7730] = (inputs[61]) | (inputs[84]);
    assign layer0_outputs[7731] = (inputs[23]) ^ (inputs[232]);
    assign layer0_outputs[7732] = ~(inputs[168]);
    assign layer0_outputs[7733] = ~(inputs[78]);
    assign layer0_outputs[7734] = inputs[164];
    assign layer0_outputs[7735] = ~((inputs[81]) | (inputs[188]));
    assign layer0_outputs[7736] = ~(inputs[21]);
    assign layer0_outputs[7737] = ~((inputs[183]) & (inputs[32]));
    assign layer0_outputs[7738] = (inputs[97]) | (inputs[228]);
    assign layer0_outputs[7739] = ~((inputs[196]) | (inputs[65]));
    assign layer0_outputs[7740] = ~(inputs[152]);
    assign layer0_outputs[7741] = ~((inputs[74]) | (inputs[67]));
    assign layer0_outputs[7742] = ~(inputs[34]);
    assign layer0_outputs[7743] = (inputs[225]) | (inputs[78]);
    assign layer0_outputs[7744] = ~((inputs[241]) | (inputs[222]));
    assign layer0_outputs[7745] = ~(inputs[185]);
    assign layer0_outputs[7746] = ~((inputs[8]) | (inputs[121]));
    assign layer0_outputs[7747] = ~(inputs[136]);
    assign layer0_outputs[7748] = inputs[107];
    assign layer0_outputs[7749] = (inputs[180]) | (inputs[228]);
    assign layer0_outputs[7750] = (inputs[150]) ^ (inputs[153]);
    assign layer0_outputs[7751] = (inputs[29]) & (inputs[21]);
    assign layer0_outputs[7752] = (inputs[175]) & ~(inputs[57]);
    assign layer0_outputs[7753] = (inputs[186]) & ~(inputs[123]);
    assign layer0_outputs[7754] = 1'b0;
    assign layer0_outputs[7755] = (inputs[183]) & ~(inputs[10]);
    assign layer0_outputs[7756] = 1'b0;
    assign layer0_outputs[7757] = 1'b0;
    assign layer0_outputs[7758] = ~(inputs[144]) | (inputs[246]);
    assign layer0_outputs[7759] = 1'b0;
    assign layer0_outputs[7760] = ~(inputs[1]);
    assign layer0_outputs[7761] = inputs[62];
    assign layer0_outputs[7762] = inputs[36];
    assign layer0_outputs[7763] = ~(inputs[213]);
    assign layer0_outputs[7764] = (inputs[127]) | (inputs[38]);
    assign layer0_outputs[7765] = ~(inputs[203]) | (inputs[109]);
    assign layer0_outputs[7766] = ~(inputs[245]) | (inputs[77]);
    assign layer0_outputs[7767] = inputs[139];
    assign layer0_outputs[7768] = (inputs[194]) & ~(inputs[126]);
    assign layer0_outputs[7769] = (inputs[176]) & ~(inputs[82]);
    assign layer0_outputs[7770] = ~((inputs[125]) ^ (inputs[127]));
    assign layer0_outputs[7771] = ~(inputs[49]);
    assign layer0_outputs[7772] = ~(inputs[140]) | (inputs[69]);
    assign layer0_outputs[7773] = ~(inputs[225]);
    assign layer0_outputs[7774] = (inputs[181]) & ~(inputs[99]);
    assign layer0_outputs[7775] = inputs[146];
    assign layer0_outputs[7776] = ~(inputs[181]);
    assign layer0_outputs[7777] = inputs[156];
    assign layer0_outputs[7778] = ~(inputs[46]) | (inputs[236]);
    assign layer0_outputs[7779] = inputs[43];
    assign layer0_outputs[7780] = ~((inputs[180]) | (inputs[2]));
    assign layer0_outputs[7781] = ~(inputs[99]) | (inputs[11]);
    assign layer0_outputs[7782] = ~((inputs[65]) | (inputs[51]));
    assign layer0_outputs[7783] = ~(inputs[150]);
    assign layer0_outputs[7784] = (inputs[32]) & ~(inputs[220]);
    assign layer0_outputs[7785] = (inputs[216]) | (inputs[215]);
    assign layer0_outputs[7786] = ~(inputs[53]);
    assign layer0_outputs[7787] = 1'b1;
    assign layer0_outputs[7788] = ~(inputs[22]) | (inputs[174]);
    assign layer0_outputs[7789] = (inputs[250]) ^ (inputs[209]);
    assign layer0_outputs[7790] = inputs[144];
    assign layer0_outputs[7791] = (inputs[230]) | (inputs[219]);
    assign layer0_outputs[7792] = ~((inputs[163]) & (inputs[112]));
    assign layer0_outputs[7793] = ~(inputs[231]);
    assign layer0_outputs[7794] = (inputs[91]) & ~(inputs[190]);
    assign layer0_outputs[7795] = (inputs[20]) | (inputs[148]);
    assign layer0_outputs[7796] = (inputs[145]) | (inputs[185]);
    assign layer0_outputs[7797] = ~((inputs[76]) | (inputs[23]));
    assign layer0_outputs[7798] = inputs[154];
    assign layer0_outputs[7799] = ~((inputs[30]) & (inputs[108]));
    assign layer0_outputs[7800] = (inputs[187]) | (inputs[108]);
    assign layer0_outputs[7801] = ~((inputs[9]) | (inputs[62]));
    assign layer0_outputs[7802] = ~(inputs[116]) | (inputs[169]);
    assign layer0_outputs[7803] = (inputs[220]) | (inputs[239]);
    assign layer0_outputs[7804] = ~((inputs[46]) & (inputs[236]));
    assign layer0_outputs[7805] = inputs[101];
    assign layer0_outputs[7806] = ~(inputs[198]);
    assign layer0_outputs[7807] = 1'b0;
    assign layer0_outputs[7808] = (inputs[78]) & ~(inputs[19]);
    assign layer0_outputs[7809] = ~(inputs[146]);
    assign layer0_outputs[7810] = (inputs[23]) & ~(inputs[118]);
    assign layer0_outputs[7811] = ~((inputs[192]) & (inputs[69]));
    assign layer0_outputs[7812] = ~(inputs[91]);
    assign layer0_outputs[7813] = inputs[255];
    assign layer0_outputs[7814] = inputs[7];
    assign layer0_outputs[7815] = ~((inputs[165]) | (inputs[143]));
    assign layer0_outputs[7816] = 1'b1;
    assign layer0_outputs[7817] = inputs[93];
    assign layer0_outputs[7818] = ~((inputs[221]) ^ (inputs[253]));
    assign layer0_outputs[7819] = inputs[58];
    assign layer0_outputs[7820] = (inputs[150]) & ~(inputs[220]);
    assign layer0_outputs[7821] = ~(inputs[41]) | (inputs[77]);
    assign layer0_outputs[7822] = 1'b1;
    assign layer0_outputs[7823] = ~(inputs[87]) | (inputs[214]);
    assign layer0_outputs[7824] = (inputs[140]) & (inputs[222]);
    assign layer0_outputs[7825] = inputs[5];
    assign layer0_outputs[7826] = ~((inputs[37]) ^ (inputs[254]));
    assign layer0_outputs[7827] = ~((inputs[49]) | (inputs[195]));
    assign layer0_outputs[7828] = ~((inputs[14]) | (inputs[54]));
    assign layer0_outputs[7829] = inputs[40];
    assign layer0_outputs[7830] = inputs[120];
    assign layer0_outputs[7831] = ~(inputs[218]) | (inputs[133]);
    assign layer0_outputs[7832] = (inputs[53]) | (inputs[161]);
    assign layer0_outputs[7833] = ~(inputs[132]);
    assign layer0_outputs[7834] = 1'b1;
    assign layer0_outputs[7835] = (inputs[69]) ^ (inputs[164]);
    assign layer0_outputs[7836] = ~(inputs[142]) | (inputs[126]);
    assign layer0_outputs[7837] = (inputs[67]) & ~(inputs[161]);
    assign layer0_outputs[7838] = ~(inputs[4]) | (inputs[90]);
    assign layer0_outputs[7839] = (inputs[95]) & ~(inputs[51]);
    assign layer0_outputs[7840] = (inputs[164]) & (inputs[35]);
    assign layer0_outputs[7841] = ~(inputs[133]) | (inputs[254]);
    assign layer0_outputs[7842] = ~((inputs[43]) | (inputs[196]));
    assign layer0_outputs[7843] = ~(inputs[42]);
    assign layer0_outputs[7844] = ~(inputs[99]) | (inputs[174]);
    assign layer0_outputs[7845] = (inputs[99]) | (inputs[23]);
    assign layer0_outputs[7846] = (inputs[85]) | (inputs[147]);
    assign layer0_outputs[7847] = ~((inputs[83]) & (inputs[80]));
    assign layer0_outputs[7848] = 1'b0;
    assign layer0_outputs[7849] = (inputs[89]) | (inputs[65]);
    assign layer0_outputs[7850] = ~(inputs[179]);
    assign layer0_outputs[7851] = inputs[202];
    assign layer0_outputs[7852] = (inputs[135]) | (inputs[107]);
    assign layer0_outputs[7853] = 1'b1;
    assign layer0_outputs[7854] = ~((inputs[253]) | (inputs[185]));
    assign layer0_outputs[7855] = ~(inputs[43]);
    assign layer0_outputs[7856] = ~(inputs[78]) | (inputs[26]);
    assign layer0_outputs[7857] = (inputs[106]) | (inputs[187]);
    assign layer0_outputs[7858] = ~((inputs[250]) | (inputs[145]));
    assign layer0_outputs[7859] = ~(inputs[111]);
    assign layer0_outputs[7860] = (inputs[222]) | (inputs[111]);
    assign layer0_outputs[7861] = ~(inputs[130]);
    assign layer0_outputs[7862] = (inputs[218]) & ~(inputs[109]);
    assign layer0_outputs[7863] = inputs[91];
    assign layer0_outputs[7864] = ~(inputs[133]);
    assign layer0_outputs[7865] = ~(inputs[84]);
    assign layer0_outputs[7866] = ~((inputs[54]) | (inputs[226]));
    assign layer0_outputs[7867] = (inputs[116]) | (inputs[112]);
    assign layer0_outputs[7868] = inputs[119];
    assign layer0_outputs[7869] = ~(inputs[2]);
    assign layer0_outputs[7870] = ~((inputs[232]) ^ (inputs[242]));
    assign layer0_outputs[7871] = ~(inputs[184]);
    assign layer0_outputs[7872] = ~(inputs[233]) | (inputs[211]);
    assign layer0_outputs[7873] = ~(inputs[249]) | (inputs[18]);
    assign layer0_outputs[7874] = ~((inputs[125]) | (inputs[94]));
    assign layer0_outputs[7875] = inputs[106];
    assign layer0_outputs[7876] = inputs[200];
    assign layer0_outputs[7877] = inputs[133];
    assign layer0_outputs[7878] = (inputs[78]) | (inputs[79]);
    assign layer0_outputs[7879] = inputs[48];
    assign layer0_outputs[7880] = ~(inputs[8]);
    assign layer0_outputs[7881] = inputs[223];
    assign layer0_outputs[7882] = ~((inputs[222]) & (inputs[7]));
    assign layer0_outputs[7883] = ~(inputs[154]);
    assign layer0_outputs[7884] = (inputs[90]) & ~(inputs[219]);
    assign layer0_outputs[7885] = inputs[107];
    assign layer0_outputs[7886] = (inputs[75]) & ~(inputs[235]);
    assign layer0_outputs[7887] = ~(inputs[115]);
    assign layer0_outputs[7888] = (inputs[81]) ^ (inputs[42]);
    assign layer0_outputs[7889] = (inputs[198]) ^ (inputs[75]);
    assign layer0_outputs[7890] = ~(inputs[166]) | (inputs[222]);
    assign layer0_outputs[7891] = ~(inputs[103]);
    assign layer0_outputs[7892] = ~((inputs[71]) ^ (inputs[74]));
    assign layer0_outputs[7893] = (inputs[200]) ^ (inputs[201]);
    assign layer0_outputs[7894] = ~(inputs[159]) | (inputs[151]);
    assign layer0_outputs[7895] = (inputs[228]) & ~(inputs[132]);
    assign layer0_outputs[7896] = inputs[0];
    assign layer0_outputs[7897] = (inputs[92]) & ~(inputs[12]);
    assign layer0_outputs[7898] = inputs[161];
    assign layer0_outputs[7899] = inputs[180];
    assign layer0_outputs[7900] = (inputs[118]) ^ (inputs[103]);
    assign layer0_outputs[7901] = inputs[168];
    assign layer0_outputs[7902] = (inputs[134]) & ~(inputs[105]);
    assign layer0_outputs[7903] = ~(inputs[103]);
    assign layer0_outputs[7904] = inputs[100];
    assign layer0_outputs[7905] = ~(inputs[103]) | (inputs[1]);
    assign layer0_outputs[7906] = 1'b1;
    assign layer0_outputs[7907] = (inputs[193]) | (inputs[5]);
    assign layer0_outputs[7908] = ~(inputs[194]) | (inputs[5]);
    assign layer0_outputs[7909] = inputs[196];
    assign layer0_outputs[7910] = ~(inputs[93]);
    assign layer0_outputs[7911] = ~((inputs[152]) | (inputs[182]));
    assign layer0_outputs[7912] = ~((inputs[44]) ^ (inputs[74]));
    assign layer0_outputs[7913] = ~((inputs[148]) | (inputs[148]));
    assign layer0_outputs[7914] = 1'b1;
    assign layer0_outputs[7915] = inputs[141];
    assign layer0_outputs[7916] = ~(inputs[8]);
    assign layer0_outputs[7917] = inputs[24];
    assign layer0_outputs[7918] = (inputs[177]) ^ (inputs[234]);
    assign layer0_outputs[7919] = ~((inputs[246]) | (inputs[207]));
    assign layer0_outputs[7920] = (inputs[221]) ^ (inputs[189]);
    assign layer0_outputs[7921] = (inputs[234]) | (inputs[207]);
    assign layer0_outputs[7922] = ~(inputs[122]);
    assign layer0_outputs[7923] = (inputs[123]) ^ (inputs[170]);
    assign layer0_outputs[7924] = ~((inputs[204]) & (inputs[139]));
    assign layer0_outputs[7925] = (inputs[243]) ^ (inputs[210]);
    assign layer0_outputs[7926] = 1'b1;
    assign layer0_outputs[7927] = ~((inputs[86]) ^ (inputs[80]));
    assign layer0_outputs[7928] = inputs[70];
    assign layer0_outputs[7929] = ~((inputs[155]) ^ (inputs[51]));
    assign layer0_outputs[7930] = ~(inputs[57]) | (inputs[20]);
    assign layer0_outputs[7931] = inputs[44];
    assign layer0_outputs[7932] = ~((inputs[33]) | (inputs[236]));
    assign layer0_outputs[7933] = inputs[143];
    assign layer0_outputs[7934] = (inputs[151]) & ~(inputs[73]);
    assign layer0_outputs[7935] = ~(inputs[56]);
    assign layer0_outputs[7936] = ~(inputs[194]);
    assign layer0_outputs[7937] = ~(inputs[118]);
    assign layer0_outputs[7938] = ~((inputs[168]) & (inputs[77]));
    assign layer0_outputs[7939] = (inputs[229]) & ~(inputs[104]);
    assign layer0_outputs[7940] = inputs[104];
    assign layer0_outputs[7941] = (inputs[212]) | (inputs[6]);
    assign layer0_outputs[7942] = ~((inputs[91]) & (inputs[163]));
    assign layer0_outputs[7943] = ~((inputs[0]) & (inputs[40]));
    assign layer0_outputs[7944] = inputs[36];
    assign layer0_outputs[7945] = ~((inputs[51]) & (inputs[169]));
    assign layer0_outputs[7946] = ~((inputs[4]) ^ (inputs[11]));
    assign layer0_outputs[7947] = ~((inputs[141]) | (inputs[132]));
    assign layer0_outputs[7948] = (inputs[219]) & ~(inputs[142]);
    assign layer0_outputs[7949] = (inputs[62]) ^ (inputs[218]);
    assign layer0_outputs[7950] = ~((inputs[220]) | (inputs[109]));
    assign layer0_outputs[7951] = inputs[148];
    assign layer0_outputs[7952] = ~(inputs[223]) | (inputs[96]);
    assign layer0_outputs[7953] = ~(inputs[187]);
    assign layer0_outputs[7954] = (inputs[101]) & ~(inputs[115]);
    assign layer0_outputs[7955] = (inputs[216]) | (inputs[9]);
    assign layer0_outputs[7956] = (inputs[166]) ^ (inputs[108]);
    assign layer0_outputs[7957] = inputs[108];
    assign layer0_outputs[7958] = (inputs[62]) ^ (inputs[247]);
    assign layer0_outputs[7959] = (inputs[212]) & ~(inputs[111]);
    assign layer0_outputs[7960] = (inputs[223]) & (inputs[128]);
    assign layer0_outputs[7961] = ~(inputs[59]);
    assign layer0_outputs[7962] = ~(inputs[165]) | (inputs[47]);
    assign layer0_outputs[7963] = (inputs[210]) & ~(inputs[27]);
    assign layer0_outputs[7964] = ~(inputs[41]);
    assign layer0_outputs[7965] = (inputs[143]) & ~(inputs[248]);
    assign layer0_outputs[7966] = inputs[169];
    assign layer0_outputs[7967] = (inputs[89]) & ~(inputs[224]);
    assign layer0_outputs[7968] = inputs[136];
    assign layer0_outputs[7969] = (inputs[212]) | (inputs[212]);
    assign layer0_outputs[7970] = ~(inputs[133]) | (inputs[137]);
    assign layer0_outputs[7971] = 1'b1;
    assign layer0_outputs[7972] = inputs[46];
    assign layer0_outputs[7973] = ~(inputs[65]) | (inputs[145]);
    assign layer0_outputs[7974] = inputs[2];
    assign layer0_outputs[7975] = inputs[20];
    assign layer0_outputs[7976] = 1'b1;
    assign layer0_outputs[7977] = (inputs[217]) & ~(inputs[123]);
    assign layer0_outputs[7978] = ~(inputs[214]);
    assign layer0_outputs[7979] = inputs[98];
    assign layer0_outputs[7980] = ~(inputs[110]);
    assign layer0_outputs[7981] = ~(inputs[87]) | (inputs[73]);
    assign layer0_outputs[7982] = (inputs[93]) | (inputs[93]);
    assign layer0_outputs[7983] = inputs[111];
    assign layer0_outputs[7984] = (inputs[97]) | (inputs[99]);
    assign layer0_outputs[7985] = 1'b0;
    assign layer0_outputs[7986] = (inputs[209]) ^ (inputs[251]);
    assign layer0_outputs[7987] = (inputs[153]) ^ (inputs[42]);
    assign layer0_outputs[7988] = ~((inputs[55]) ^ (inputs[6]));
    assign layer0_outputs[7989] = (inputs[65]) ^ (inputs[35]);
    assign layer0_outputs[7990] = ~((inputs[156]) | (inputs[163]));
    assign layer0_outputs[7991] = ~((inputs[208]) ^ (inputs[38]));
    assign layer0_outputs[7992] = ~(inputs[80]) | (inputs[198]);
    assign layer0_outputs[7993] = (inputs[190]) ^ (inputs[180]);
    assign layer0_outputs[7994] = ~((inputs[63]) ^ (inputs[204]));
    assign layer0_outputs[7995] = ~(inputs[99]);
    assign layer0_outputs[7996] = ~(inputs[233]);
    assign layer0_outputs[7997] = ~(inputs[247]) | (inputs[163]);
    assign layer0_outputs[7998] = ~(inputs[3]) | (inputs[206]);
    assign layer0_outputs[7999] = inputs[36];
    assign layer0_outputs[8000] = (inputs[203]) ^ (inputs[135]);
    assign layer0_outputs[8001] = ~(inputs[92]) | (inputs[235]);
    assign layer0_outputs[8002] = (inputs[32]) ^ (inputs[63]);
    assign layer0_outputs[8003] = ~((inputs[112]) | (inputs[160]));
    assign layer0_outputs[8004] = ~((inputs[238]) | (inputs[191]));
    assign layer0_outputs[8005] = (inputs[213]) & ~(inputs[49]);
    assign layer0_outputs[8006] = inputs[85];
    assign layer0_outputs[8007] = (inputs[92]) & ~(inputs[83]);
    assign layer0_outputs[8008] = ~((inputs[201]) | (inputs[151]));
    assign layer0_outputs[8009] = ~((inputs[195]) | (inputs[233]));
    assign layer0_outputs[8010] = inputs[41];
    assign layer0_outputs[8011] = (inputs[23]) & ~(inputs[188]);
    assign layer0_outputs[8012] = (inputs[93]) ^ (inputs[160]);
    assign layer0_outputs[8013] = inputs[92];
    assign layer0_outputs[8014] = (inputs[46]) & ~(inputs[8]);
    assign layer0_outputs[8015] = (inputs[65]) | (inputs[116]);
    assign layer0_outputs[8016] = (inputs[31]) ^ (inputs[39]);
    assign layer0_outputs[8017] = (inputs[199]) & ~(inputs[147]);
    assign layer0_outputs[8018] = inputs[194];
    assign layer0_outputs[8019] = (inputs[16]) & ~(inputs[160]);
    assign layer0_outputs[8020] = ~(inputs[10]);
    assign layer0_outputs[8021] = (inputs[187]) | (inputs[49]);
    assign layer0_outputs[8022] = ~((inputs[178]) | (inputs[245]));
    assign layer0_outputs[8023] = ~(inputs[149]) | (inputs[124]);
    assign layer0_outputs[8024] = (inputs[13]) | (inputs[2]);
    assign layer0_outputs[8025] = (inputs[176]) | (inputs[181]);
    assign layer0_outputs[8026] = ~(inputs[221]);
    assign layer0_outputs[8027] = ~(inputs[144]) | (inputs[0]);
    assign layer0_outputs[8028] = ~(inputs[203]) | (inputs[117]);
    assign layer0_outputs[8029] = (inputs[115]) & ~(inputs[19]);
    assign layer0_outputs[8030] = ~((inputs[247]) & (inputs[172]));
    assign layer0_outputs[8031] = ~(inputs[146]);
    assign layer0_outputs[8032] = ~(inputs[178]) | (inputs[179]);
    assign layer0_outputs[8033] = (inputs[50]) | (inputs[33]);
    assign layer0_outputs[8034] = (inputs[119]) | (inputs[237]);
    assign layer0_outputs[8035] = (inputs[96]) & ~(inputs[77]);
    assign layer0_outputs[8036] = (inputs[200]) | (inputs[124]);
    assign layer0_outputs[8037] = ~((inputs[115]) ^ (inputs[173]));
    assign layer0_outputs[8038] = (inputs[102]) & ~(inputs[4]);
    assign layer0_outputs[8039] = (inputs[189]) & ~(inputs[154]);
    assign layer0_outputs[8040] = ~((inputs[229]) | (inputs[224]));
    assign layer0_outputs[8041] = (inputs[175]) | (inputs[146]);
    assign layer0_outputs[8042] = (inputs[36]) | (inputs[2]);
    assign layer0_outputs[8043] = ~(inputs[192]);
    assign layer0_outputs[8044] = (inputs[205]) | (inputs[133]);
    assign layer0_outputs[8045] = (inputs[161]) & (inputs[158]);
    assign layer0_outputs[8046] = ~(inputs[170]);
    assign layer0_outputs[8047] = (inputs[53]) & ~(inputs[144]);
    assign layer0_outputs[8048] = ~((inputs[67]) | (inputs[230]));
    assign layer0_outputs[8049] = (inputs[210]) & ~(inputs[142]);
    assign layer0_outputs[8050] = (inputs[97]) & ~(inputs[121]);
    assign layer0_outputs[8051] = ~(inputs[54]);
    assign layer0_outputs[8052] = inputs[140];
    assign layer0_outputs[8053] = ~((inputs[82]) ^ (inputs[111]));
    assign layer0_outputs[8054] = (inputs[58]) ^ (inputs[43]);
    assign layer0_outputs[8055] = ~(inputs[113]) | (inputs[72]);
    assign layer0_outputs[8056] = ~(inputs[186]) | (inputs[106]);
    assign layer0_outputs[8057] = ~(inputs[146]);
    assign layer0_outputs[8058] = (inputs[242]) | (inputs[39]);
    assign layer0_outputs[8059] = inputs[16];
    assign layer0_outputs[8060] = (inputs[143]) ^ (inputs[204]);
    assign layer0_outputs[8061] = ~((inputs[174]) | (inputs[199]));
    assign layer0_outputs[8062] = inputs[119];
    assign layer0_outputs[8063] = ~((inputs[100]) | (inputs[141]));
    assign layer0_outputs[8064] = (inputs[201]) & ~(inputs[40]);
    assign layer0_outputs[8065] = (inputs[230]) | (inputs[176]);
    assign layer0_outputs[8066] = ~(inputs[157]);
    assign layer0_outputs[8067] = ~(inputs[187]);
    assign layer0_outputs[8068] = (inputs[60]) & ~(inputs[231]);
    assign layer0_outputs[8069] = ~(inputs[225]);
    assign layer0_outputs[8070] = ~((inputs[254]) & (inputs[12]));
    assign layer0_outputs[8071] = ~(inputs[224]) | (inputs[109]);
    assign layer0_outputs[8072] = (inputs[144]) | (inputs[34]);
    assign layer0_outputs[8073] = inputs[7];
    assign layer0_outputs[8074] = (inputs[123]) & ~(inputs[194]);
    assign layer0_outputs[8075] = ~(inputs[158]);
    assign layer0_outputs[8076] = (inputs[240]) | (inputs[64]);
    assign layer0_outputs[8077] = ~(inputs[58]);
    assign layer0_outputs[8078] = (inputs[59]) | (inputs[75]);
    assign layer0_outputs[8079] = (inputs[150]) & ~(inputs[233]);
    assign layer0_outputs[8080] = ~((inputs[204]) | (inputs[11]));
    assign layer0_outputs[8081] = ~((inputs[87]) & (inputs[143]));
    assign layer0_outputs[8082] = (inputs[112]) & ~(inputs[87]);
    assign layer0_outputs[8083] = (inputs[191]) & ~(inputs[104]);
    assign layer0_outputs[8084] = inputs[188];
    assign layer0_outputs[8085] = (inputs[212]) & ~(inputs[53]);
    assign layer0_outputs[8086] = ~((inputs[205]) | (inputs[23]));
    assign layer0_outputs[8087] = ~(inputs[96]) | (inputs[1]);
    assign layer0_outputs[8088] = ~((inputs[99]) | (inputs[140]));
    assign layer0_outputs[8089] = ~(inputs[187]) | (inputs[184]);
    assign layer0_outputs[8090] = inputs[120];
    assign layer0_outputs[8091] = (inputs[188]) & ~(inputs[110]);
    assign layer0_outputs[8092] = (inputs[195]) & ~(inputs[2]);
    assign layer0_outputs[8093] = ~((inputs[2]) | (inputs[200]));
    assign layer0_outputs[8094] = ~((inputs[159]) & (inputs[2]));
    assign layer0_outputs[8095] = ~((inputs[144]) ^ (inputs[163]));
    assign layer0_outputs[8096] = inputs[149];
    assign layer0_outputs[8097] = (inputs[241]) | (inputs[202]);
    assign layer0_outputs[8098] = (inputs[251]) | (inputs[163]);
    assign layer0_outputs[8099] = ~((inputs[185]) & (inputs[224]));
    assign layer0_outputs[8100] = ~(inputs[178]);
    assign layer0_outputs[8101] = ~(inputs[127]);
    assign layer0_outputs[8102] = (inputs[253]) | (inputs[41]);
    assign layer0_outputs[8103] = ~((inputs[189]) | (inputs[239]));
    assign layer0_outputs[8104] = ~(inputs[6]);
    assign layer0_outputs[8105] = 1'b1;
    assign layer0_outputs[8106] = ~((inputs[35]) | (inputs[206]));
    assign layer0_outputs[8107] = ~(inputs[151]) | (inputs[185]);
    assign layer0_outputs[8108] = ~((inputs[239]) | (inputs[246]));
    assign layer0_outputs[8109] = ~(inputs[229]);
    assign layer0_outputs[8110] = ~(inputs[152]);
    assign layer0_outputs[8111] = inputs[154];
    assign layer0_outputs[8112] = ~((inputs[107]) | (inputs[15]));
    assign layer0_outputs[8113] = ~((inputs[200]) | (inputs[206]));
    assign layer0_outputs[8114] = ~((inputs[162]) | (inputs[161]));
    assign layer0_outputs[8115] = ~((inputs[67]) ^ (inputs[128]));
    assign layer0_outputs[8116] = ~(inputs[61]);
    assign layer0_outputs[8117] = ~(inputs[240]);
    assign layer0_outputs[8118] = inputs[35];
    assign layer0_outputs[8119] = ~(inputs[122]) | (inputs[181]);
    assign layer0_outputs[8120] = (inputs[199]) ^ (inputs[89]);
    assign layer0_outputs[8121] = (inputs[89]) & ~(inputs[81]);
    assign layer0_outputs[8122] = (inputs[17]) | (inputs[155]);
    assign layer0_outputs[8123] = ~(inputs[22]);
    assign layer0_outputs[8124] = (inputs[235]) | (inputs[206]);
    assign layer0_outputs[8125] = inputs[209];
    assign layer0_outputs[8126] = (inputs[34]) | (inputs[21]);
    assign layer0_outputs[8127] = inputs[125];
    assign layer0_outputs[8128] = ~(inputs[86]);
    assign layer0_outputs[8129] = ~((inputs[56]) & (inputs[195]));
    assign layer0_outputs[8130] = ~((inputs[179]) | (inputs[11]));
    assign layer0_outputs[8131] = (inputs[244]) & (inputs[226]);
    assign layer0_outputs[8132] = ~((inputs[190]) | (inputs[117]));
    assign layer0_outputs[8133] = ~((inputs[124]) ^ (inputs[92]));
    assign layer0_outputs[8134] = ~(inputs[215]);
    assign layer0_outputs[8135] = (inputs[177]) | (inputs[117]);
    assign layer0_outputs[8136] = ~(inputs[133]) | (inputs[177]);
    assign layer0_outputs[8137] = ~((inputs[151]) | (inputs[221]));
    assign layer0_outputs[8138] = (inputs[24]) ^ (inputs[72]);
    assign layer0_outputs[8139] = (inputs[100]) & (inputs[22]);
    assign layer0_outputs[8140] = ~(inputs[206]);
    assign layer0_outputs[8141] = ~(inputs[41]);
    assign layer0_outputs[8142] = ~((inputs[171]) ^ (inputs[236]));
    assign layer0_outputs[8143] = ~((inputs[125]) ^ (inputs[19]));
    assign layer0_outputs[8144] = ~(inputs[160]);
    assign layer0_outputs[8145] = ~(inputs[57]);
    assign layer0_outputs[8146] = ~(inputs[137]);
    assign layer0_outputs[8147] = inputs[250];
    assign layer0_outputs[8148] = ~((inputs[87]) & (inputs[244]));
    assign layer0_outputs[8149] = ~(inputs[18]);
    assign layer0_outputs[8150] = ~((inputs[169]) | (inputs[63]));
    assign layer0_outputs[8151] = ~(inputs[91]);
    assign layer0_outputs[8152] = inputs[221];
    assign layer0_outputs[8153] = ~(inputs[188]) | (inputs[32]);
    assign layer0_outputs[8154] = ~((inputs[143]) | (inputs[12]));
    assign layer0_outputs[8155] = ~((inputs[10]) ^ (inputs[43]));
    assign layer0_outputs[8156] = ~((inputs[35]) | (inputs[17]));
    assign layer0_outputs[8157] = (inputs[209]) & ~(inputs[1]);
    assign layer0_outputs[8158] = ~((inputs[255]) & (inputs[15]));
    assign layer0_outputs[8159] = ~(inputs[214]);
    assign layer0_outputs[8160] = inputs[67];
    assign layer0_outputs[8161] = inputs[174];
    assign layer0_outputs[8162] = ~(inputs[116]) | (inputs[2]);
    assign layer0_outputs[8163] = (inputs[138]) | (inputs[149]);
    assign layer0_outputs[8164] = ~(inputs[46]);
    assign layer0_outputs[8165] = ~(inputs[68]);
    assign layer0_outputs[8166] = ~(inputs[201]) | (inputs[203]);
    assign layer0_outputs[8167] = inputs[151];
    assign layer0_outputs[8168] = ~((inputs[242]) ^ (inputs[64]));
    assign layer0_outputs[8169] = ~((inputs[79]) ^ (inputs[141]));
    assign layer0_outputs[8170] = (inputs[83]) | (inputs[88]);
    assign layer0_outputs[8171] = ~((inputs[199]) & (inputs[210]));
    assign layer0_outputs[8172] = (inputs[165]) & ~(inputs[166]);
    assign layer0_outputs[8173] = ~(inputs[98]) | (inputs[238]);
    assign layer0_outputs[8174] = (inputs[197]) & ~(inputs[101]);
    assign layer0_outputs[8175] = ~((inputs[206]) ^ (inputs[85]));
    assign layer0_outputs[8176] = inputs[100];
    assign layer0_outputs[8177] = (inputs[169]) ^ (inputs[171]);
    assign layer0_outputs[8178] = (inputs[115]) | (inputs[130]);
    assign layer0_outputs[8179] = (inputs[89]) ^ (inputs[188]);
    assign layer0_outputs[8180] = inputs[189];
    assign layer0_outputs[8181] = (inputs[222]) & ~(inputs[200]);
    assign layer0_outputs[8182] = inputs[133];
    assign layer0_outputs[8183] = (inputs[246]) ^ (inputs[198]);
    assign layer0_outputs[8184] = ~(inputs[237]);
    assign layer0_outputs[8185] = ~((inputs[131]) ^ (inputs[101]));
    assign layer0_outputs[8186] = (inputs[57]) ^ (inputs[88]);
    assign layer0_outputs[8187] = ~((inputs[126]) | (inputs[0]));
    assign layer0_outputs[8188] = (inputs[72]) & ~(inputs[41]);
    assign layer0_outputs[8189] = ~(inputs[232]) | (inputs[185]);
    assign layer0_outputs[8190] = (inputs[37]) | (inputs[5]);
    assign layer0_outputs[8191] = ~(inputs[230]);
    assign layer0_outputs[8192] = (inputs[195]) & ~(inputs[239]);
    assign layer0_outputs[8193] = (inputs[71]) & ~(inputs[120]);
    assign layer0_outputs[8194] = (inputs[230]) & ~(inputs[20]);
    assign layer0_outputs[8195] = (inputs[183]) ^ (inputs[125]);
    assign layer0_outputs[8196] = inputs[131];
    assign layer0_outputs[8197] = ~((inputs[200]) & (inputs[218]));
    assign layer0_outputs[8198] = ~((inputs[161]) | (inputs[218]));
    assign layer0_outputs[8199] = ~(inputs[71]);
    assign layer0_outputs[8200] = 1'b1;
    assign layer0_outputs[8201] = (inputs[238]) ^ (inputs[143]);
    assign layer0_outputs[8202] = inputs[235];
    assign layer0_outputs[8203] = ~(inputs[45]);
    assign layer0_outputs[8204] = (inputs[234]) | (inputs[224]);
    assign layer0_outputs[8205] = (inputs[208]) | (inputs[32]);
    assign layer0_outputs[8206] = inputs[167];
    assign layer0_outputs[8207] = (inputs[135]) & ~(inputs[133]);
    assign layer0_outputs[8208] = (inputs[76]) & ~(inputs[253]);
    assign layer0_outputs[8209] = (inputs[10]) | (inputs[247]);
    assign layer0_outputs[8210] = (inputs[195]) & ~(inputs[19]);
    assign layer0_outputs[8211] = ~(inputs[187]) | (inputs[5]);
    assign layer0_outputs[8212] = ~(inputs[147]);
    assign layer0_outputs[8213] = inputs[111];
    assign layer0_outputs[8214] = (inputs[172]) & ~(inputs[63]);
    assign layer0_outputs[8215] = (inputs[235]) & ~(inputs[97]);
    assign layer0_outputs[8216] = 1'b0;
    assign layer0_outputs[8217] = ~(inputs[167]);
    assign layer0_outputs[8218] = ~(inputs[166]) | (inputs[198]);
    assign layer0_outputs[8219] = (inputs[79]) ^ (inputs[226]);
    assign layer0_outputs[8220] = (inputs[133]) ^ (inputs[152]);
    assign layer0_outputs[8221] = ~(inputs[164]);
    assign layer0_outputs[8222] = (inputs[65]) | (inputs[103]);
    assign layer0_outputs[8223] = ~(inputs[98]);
    assign layer0_outputs[8224] = (inputs[43]) & ~(inputs[234]);
    assign layer0_outputs[8225] = (inputs[244]) & ~(inputs[120]);
    assign layer0_outputs[8226] = inputs[130];
    assign layer0_outputs[8227] = ~((inputs[241]) | (inputs[15]));
    assign layer0_outputs[8228] = ~(inputs[85]) | (inputs[164]);
    assign layer0_outputs[8229] = (inputs[211]) & (inputs[129]);
    assign layer0_outputs[8230] = inputs[201];
    assign layer0_outputs[8231] = ~((inputs[80]) | (inputs[5]));
    assign layer0_outputs[8232] = inputs[21];
    assign layer0_outputs[8233] = (inputs[22]) & ~(inputs[18]);
    assign layer0_outputs[8234] = (inputs[58]) & ~(inputs[176]);
    assign layer0_outputs[8235] = ~(inputs[40]) | (inputs[113]);
    assign layer0_outputs[8236] = ~(inputs[104]) | (inputs[102]);
    assign layer0_outputs[8237] = (inputs[137]) & ~(inputs[178]);
    assign layer0_outputs[8238] = (inputs[29]) & ~(inputs[142]);
    assign layer0_outputs[8239] = inputs[85];
    assign layer0_outputs[8240] = ~(inputs[255]);
    assign layer0_outputs[8241] = ~(inputs[68]);
    assign layer0_outputs[8242] = inputs[233];
    assign layer0_outputs[8243] = ~((inputs[107]) & (inputs[23]));
    assign layer0_outputs[8244] = ~((inputs[120]) & (inputs[120]));
    assign layer0_outputs[8245] = ~(inputs[150]);
    assign layer0_outputs[8246] = ~(inputs[149]) | (inputs[44]);
    assign layer0_outputs[8247] = ~(inputs[68]);
    assign layer0_outputs[8248] = inputs[94];
    assign layer0_outputs[8249] = (inputs[37]) ^ (inputs[254]);
    assign layer0_outputs[8250] = ~(inputs[90]) | (inputs[192]);
    assign layer0_outputs[8251] = ~(inputs[111]);
    assign layer0_outputs[8252] = inputs[98];
    assign layer0_outputs[8253] = ~(inputs[173]);
    assign layer0_outputs[8254] = ~(inputs[224]) | (inputs[181]);
    assign layer0_outputs[8255] = 1'b0;
    assign layer0_outputs[8256] = ~(inputs[204]) | (inputs[32]);
    assign layer0_outputs[8257] = (inputs[236]) & ~(inputs[156]);
    assign layer0_outputs[8258] = inputs[144];
    assign layer0_outputs[8259] = 1'b0;
    assign layer0_outputs[8260] = (inputs[133]) & ~(inputs[34]);
    assign layer0_outputs[8261] = ~((inputs[133]) & (inputs[233]));
    assign layer0_outputs[8262] = ~((inputs[47]) | (inputs[52]));
    assign layer0_outputs[8263] = ~((inputs[114]) ^ (inputs[156]));
    assign layer0_outputs[8264] = 1'b1;
    assign layer0_outputs[8265] = ~(inputs[45]);
    assign layer0_outputs[8266] = ~((inputs[72]) | (inputs[235]));
    assign layer0_outputs[8267] = ~(inputs[232]);
    assign layer0_outputs[8268] = (inputs[176]) | (inputs[217]);
    assign layer0_outputs[8269] = inputs[29];
    assign layer0_outputs[8270] = inputs[64];
    assign layer0_outputs[8271] = ~((inputs[231]) & (inputs[101]));
    assign layer0_outputs[8272] = (inputs[181]) | (inputs[254]);
    assign layer0_outputs[8273] = (inputs[88]) & ~(inputs[233]);
    assign layer0_outputs[8274] = ~((inputs[181]) | (inputs[125]));
    assign layer0_outputs[8275] = ~(inputs[135]);
    assign layer0_outputs[8276] = ~(inputs[244]) | (inputs[86]);
    assign layer0_outputs[8277] = (inputs[35]) | (inputs[253]);
    assign layer0_outputs[8278] = ~(inputs[90]) | (inputs[221]);
    assign layer0_outputs[8279] = ~(inputs[31]);
    assign layer0_outputs[8280] = ~(inputs[8]);
    assign layer0_outputs[8281] = ~((inputs[11]) | (inputs[66]));
    assign layer0_outputs[8282] = 1'b0;
    assign layer0_outputs[8283] = ~(inputs[82]) | (inputs[189]);
    assign layer0_outputs[8284] = ~(inputs[118]);
    assign layer0_outputs[8285] = ~(inputs[86]);
    assign layer0_outputs[8286] = inputs[245];
    assign layer0_outputs[8287] = ~(inputs[105]);
    assign layer0_outputs[8288] = ~((inputs[149]) | (inputs[48]));
    assign layer0_outputs[8289] = ~(inputs[231]) | (inputs[216]);
    assign layer0_outputs[8290] = ~(inputs[193]) | (inputs[48]);
    assign layer0_outputs[8291] = ~(inputs[124]);
    assign layer0_outputs[8292] = 1'b0;
    assign layer0_outputs[8293] = inputs[40];
    assign layer0_outputs[8294] = ~(inputs[71]);
    assign layer0_outputs[8295] = inputs[110];
    assign layer0_outputs[8296] = ~((inputs[67]) ^ (inputs[20]));
    assign layer0_outputs[8297] = (inputs[65]) | (inputs[29]);
    assign layer0_outputs[8298] = inputs[49];
    assign layer0_outputs[8299] = ~((inputs[162]) | (inputs[203]));
    assign layer0_outputs[8300] = ~((inputs[149]) | (inputs[116]));
    assign layer0_outputs[8301] = ~((inputs[151]) | (inputs[227]));
    assign layer0_outputs[8302] = ~(inputs[91]);
    assign layer0_outputs[8303] = ~((inputs[200]) & (inputs[166]));
    assign layer0_outputs[8304] = ~((inputs[110]) | (inputs[182]));
    assign layer0_outputs[8305] = ~((inputs[174]) | (inputs[179]));
    assign layer0_outputs[8306] = ~(inputs[173]);
    assign layer0_outputs[8307] = ~(inputs[56]);
    assign layer0_outputs[8308] = inputs[133];
    assign layer0_outputs[8309] = (inputs[182]) & ~(inputs[70]);
    assign layer0_outputs[8310] = ~(inputs[199]) | (inputs[175]);
    assign layer0_outputs[8311] = ~(inputs[234]);
    assign layer0_outputs[8312] = ~((inputs[248]) | (inputs[160]));
    assign layer0_outputs[8313] = (inputs[196]) & ~(inputs[132]);
    assign layer0_outputs[8314] = inputs[126];
    assign layer0_outputs[8315] = ~(inputs[161]);
    assign layer0_outputs[8316] = ~(inputs[1]);
    assign layer0_outputs[8317] = (inputs[43]) & ~(inputs[16]);
    assign layer0_outputs[8318] = 1'b0;
    assign layer0_outputs[8319] = ~((inputs[160]) ^ (inputs[228]));
    assign layer0_outputs[8320] = ~((inputs[193]) & (inputs[1]));
    assign layer0_outputs[8321] = (inputs[131]) ^ (inputs[64]);
    assign layer0_outputs[8322] = ~((inputs[220]) | (inputs[107]));
    assign layer0_outputs[8323] = (inputs[1]) ^ (inputs[151]);
    assign layer0_outputs[8324] = (inputs[198]) & (inputs[203]);
    assign layer0_outputs[8325] = (inputs[73]) | (inputs[90]);
    assign layer0_outputs[8326] = ~(inputs[79]) | (inputs[207]);
    assign layer0_outputs[8327] = ~(inputs[4]) | (inputs[190]);
    assign layer0_outputs[8328] = inputs[202];
    assign layer0_outputs[8329] = ~((inputs[69]) | (inputs[185]));
    assign layer0_outputs[8330] = ~((inputs[195]) ^ (inputs[59]));
    assign layer0_outputs[8331] = inputs[146];
    assign layer0_outputs[8332] = inputs[172];
    assign layer0_outputs[8333] = ~((inputs[80]) | (inputs[167]));
    assign layer0_outputs[8334] = (inputs[50]) & (inputs[243]);
    assign layer0_outputs[8335] = ~(inputs[55]);
    assign layer0_outputs[8336] = ~((inputs[5]) | (inputs[180]));
    assign layer0_outputs[8337] = ~((inputs[243]) ^ (inputs[12]));
    assign layer0_outputs[8338] = ~(inputs[83]);
    assign layer0_outputs[8339] = ~(inputs[155]) | (inputs[15]);
    assign layer0_outputs[8340] = 1'b1;
    assign layer0_outputs[8341] = inputs[59];
    assign layer0_outputs[8342] = (inputs[130]) | (inputs[242]);
    assign layer0_outputs[8343] = inputs[130];
    assign layer0_outputs[8344] = (inputs[163]) | (inputs[49]);
    assign layer0_outputs[8345] = ~((inputs[162]) | (inputs[87]));
    assign layer0_outputs[8346] = ~((inputs[176]) | (inputs[48]));
    assign layer0_outputs[8347] = ~(inputs[183]);
    assign layer0_outputs[8348] = ~((inputs[241]) ^ (inputs[165]));
    assign layer0_outputs[8349] = ~(inputs[1]);
    assign layer0_outputs[8350] = (inputs[60]) ^ (inputs[43]);
    assign layer0_outputs[8351] = ~(inputs[127]) | (inputs[13]);
    assign layer0_outputs[8352] = inputs[113];
    assign layer0_outputs[8353] = ~((inputs[145]) | (inputs[14]));
    assign layer0_outputs[8354] = (inputs[5]) | (inputs[246]);
    assign layer0_outputs[8355] = ~((inputs[2]) ^ (inputs[175]));
    assign layer0_outputs[8356] = ~(inputs[184]) | (inputs[7]);
    assign layer0_outputs[8357] = (inputs[49]) | (inputs[190]);
    assign layer0_outputs[8358] = (inputs[113]) & ~(inputs[28]);
    assign layer0_outputs[8359] = (inputs[243]) ^ (inputs[95]);
    assign layer0_outputs[8360] = inputs[162];
    assign layer0_outputs[8361] = inputs[57];
    assign layer0_outputs[8362] = ~(inputs[232]) | (inputs[126]);
    assign layer0_outputs[8363] = ~((inputs[56]) | (inputs[5]));
    assign layer0_outputs[8364] = ~(inputs[49]);
    assign layer0_outputs[8365] = ~(inputs[144]) | (inputs[143]);
    assign layer0_outputs[8366] = ~((inputs[111]) ^ (inputs[9]));
    assign layer0_outputs[8367] = 1'b0;
    assign layer0_outputs[8368] = ~(inputs[135]) | (inputs[92]);
    assign layer0_outputs[8369] = inputs[187];
    assign layer0_outputs[8370] = ~(inputs[42]) | (inputs[99]);
    assign layer0_outputs[8371] = ~(inputs[69]);
    assign layer0_outputs[8372] = (inputs[176]) ^ (inputs[88]);
    assign layer0_outputs[8373] = ~((inputs[190]) ^ (inputs[139]));
    assign layer0_outputs[8374] = ~(inputs[140]) | (inputs[185]);
    assign layer0_outputs[8375] = ~((inputs[205]) | (inputs[167]));
    assign layer0_outputs[8376] = ~(inputs[109]);
    assign layer0_outputs[8377] = 1'b1;
    assign layer0_outputs[8378] = (inputs[218]) | (inputs[77]);
    assign layer0_outputs[8379] = (inputs[200]) | (inputs[255]);
    assign layer0_outputs[8380] = (inputs[11]) | (inputs[169]);
    assign layer0_outputs[8381] = inputs[21];
    assign layer0_outputs[8382] = 1'b0;
    assign layer0_outputs[8383] = ~(inputs[88]);
    assign layer0_outputs[8384] = (inputs[37]) ^ (inputs[247]);
    assign layer0_outputs[8385] = ~(inputs[221]);
    assign layer0_outputs[8386] = (inputs[8]) & ~(inputs[15]);
    assign layer0_outputs[8387] = inputs[198];
    assign layer0_outputs[8388] = ~((inputs[175]) | (inputs[209]));
    assign layer0_outputs[8389] = ~(inputs[136]) | (inputs[252]);
    assign layer0_outputs[8390] = ~((inputs[204]) & (inputs[182]));
    assign layer0_outputs[8391] = ~((inputs[226]) | (inputs[193]));
    assign layer0_outputs[8392] = inputs[47];
    assign layer0_outputs[8393] = ~((inputs[187]) ^ (inputs[37]));
    assign layer0_outputs[8394] = inputs[56];
    assign layer0_outputs[8395] = inputs[92];
    assign layer0_outputs[8396] = inputs[178];
    assign layer0_outputs[8397] = inputs[121];
    assign layer0_outputs[8398] = ~(inputs[119]) | (inputs[10]);
    assign layer0_outputs[8399] = ~((inputs[250]) ^ (inputs[227]));
    assign layer0_outputs[8400] = ~(inputs[187]) | (inputs[126]);
    assign layer0_outputs[8401] = inputs[149];
    assign layer0_outputs[8402] = 1'b0;
    assign layer0_outputs[8403] = ~(inputs[134]);
    assign layer0_outputs[8404] = ~((inputs[181]) ^ (inputs[39]));
    assign layer0_outputs[8405] = (inputs[205]) & ~(inputs[145]);
    assign layer0_outputs[8406] = ~((inputs[161]) ^ (inputs[16]));
    assign layer0_outputs[8407] = ~((inputs[138]) ^ (inputs[61]));
    assign layer0_outputs[8408] = ~((inputs[186]) ^ (inputs[147]));
    assign layer0_outputs[8409] = ~(inputs[94]) | (inputs[237]);
    assign layer0_outputs[8410] = ~((inputs[117]) | (inputs[205]));
    assign layer0_outputs[8411] = ~((inputs[106]) ^ (inputs[48]));
    assign layer0_outputs[8412] = ~(inputs[36]) | (inputs[144]);
    assign layer0_outputs[8413] = ~(inputs[213]);
    assign layer0_outputs[8414] = (inputs[2]) | (inputs[61]);
    assign layer0_outputs[8415] = inputs[99];
    assign layer0_outputs[8416] = (inputs[170]) ^ (inputs[162]);
    assign layer0_outputs[8417] = ~((inputs[135]) | (inputs[7]));
    assign layer0_outputs[8418] = (inputs[46]) | (inputs[16]);
    assign layer0_outputs[8419] = inputs[185];
    assign layer0_outputs[8420] = (inputs[246]) | (inputs[95]);
    assign layer0_outputs[8421] = inputs[212];
    assign layer0_outputs[8422] = ~(inputs[212]) | (inputs[111]);
    assign layer0_outputs[8423] = ~(inputs[102]);
    assign layer0_outputs[8424] = (inputs[240]) & ~(inputs[42]);
    assign layer0_outputs[8425] = ~(inputs[203]) | (inputs[15]);
    assign layer0_outputs[8426] = ~(inputs[241]) | (inputs[100]);
    assign layer0_outputs[8427] = ~((inputs[143]) | (inputs[2]));
    assign layer0_outputs[8428] = (inputs[181]) & ~(inputs[148]);
    assign layer0_outputs[8429] = inputs[146];
    assign layer0_outputs[8430] = (inputs[101]) & ~(inputs[108]);
    assign layer0_outputs[8431] = ~(inputs[145]);
    assign layer0_outputs[8432] = ~(inputs[166]) | (inputs[191]);
    assign layer0_outputs[8433] = ~(inputs[86]);
    assign layer0_outputs[8434] = ~(inputs[235]);
    assign layer0_outputs[8435] = ~((inputs[73]) ^ (inputs[62]));
    assign layer0_outputs[8436] = (inputs[81]) & ~(inputs[204]);
    assign layer0_outputs[8437] = ~(inputs[212]) | (inputs[47]);
    assign layer0_outputs[8438] = (inputs[117]) & (inputs[75]);
    assign layer0_outputs[8439] = (inputs[164]) & ~(inputs[58]);
    assign layer0_outputs[8440] = ~(inputs[131]);
    assign layer0_outputs[8441] = ~(inputs[174]);
    assign layer0_outputs[8442] = inputs[139];
    assign layer0_outputs[8443] = 1'b1;
    assign layer0_outputs[8444] = ~((inputs[90]) ^ (inputs[87]));
    assign layer0_outputs[8445] = inputs[17];
    assign layer0_outputs[8446] = ~((inputs[198]) | (inputs[182]));
    assign layer0_outputs[8447] = ~((inputs[205]) & (inputs[52]));
    assign layer0_outputs[8448] = ~(inputs[36]);
    assign layer0_outputs[8449] = ~(inputs[203]) | (inputs[164]);
    assign layer0_outputs[8450] = ~((inputs[232]) & (inputs[147]));
    assign layer0_outputs[8451] = (inputs[245]) & ~(inputs[61]);
    assign layer0_outputs[8452] = ~(inputs[245]) | (inputs[5]);
    assign layer0_outputs[8453] = ~((inputs[53]) ^ (inputs[9]));
    assign layer0_outputs[8454] = ~(inputs[222]);
    assign layer0_outputs[8455] = (inputs[58]) & (inputs[74]);
    assign layer0_outputs[8456] = 1'b1;
    assign layer0_outputs[8457] = ~(inputs[128]);
    assign layer0_outputs[8458] = ~((inputs[126]) | (inputs[127]));
    assign layer0_outputs[8459] = inputs[118];
    assign layer0_outputs[8460] = ~(inputs[157]) | (inputs[29]);
    assign layer0_outputs[8461] = ~(inputs[57]) | (inputs[161]);
    assign layer0_outputs[8462] = inputs[100];
    assign layer0_outputs[8463] = inputs[165];
    assign layer0_outputs[8464] = ~(inputs[137]);
    assign layer0_outputs[8465] = (inputs[251]) ^ (inputs[187]);
    assign layer0_outputs[8466] = inputs[54];
    assign layer0_outputs[8467] = inputs[214];
    assign layer0_outputs[8468] = (inputs[132]) & ~(inputs[251]);
    assign layer0_outputs[8469] = (inputs[134]) & ~(inputs[123]);
    assign layer0_outputs[8470] = (inputs[23]) | (inputs[129]);
    assign layer0_outputs[8471] = ~((inputs[64]) | (inputs[53]));
    assign layer0_outputs[8472] = (inputs[178]) & (inputs[131]);
    assign layer0_outputs[8473] = (inputs[158]) ^ (inputs[235]);
    assign layer0_outputs[8474] = ~((inputs[114]) | (inputs[115]));
    assign layer0_outputs[8475] = inputs[96];
    assign layer0_outputs[8476] = 1'b0;
    assign layer0_outputs[8477] = ~((inputs[221]) | (inputs[119]));
    assign layer0_outputs[8478] = inputs[202];
    assign layer0_outputs[8479] = (inputs[151]) & ~(inputs[115]);
    assign layer0_outputs[8480] = ~(inputs[147]) | (inputs[14]);
    assign layer0_outputs[8481] = ~((inputs[3]) | (inputs[180]));
    assign layer0_outputs[8482] = (inputs[107]) & ~(inputs[191]);
    assign layer0_outputs[8483] = (inputs[166]) | (inputs[24]);
    assign layer0_outputs[8484] = (inputs[197]) & ~(inputs[141]);
    assign layer0_outputs[8485] = (inputs[64]) & ~(inputs[242]);
    assign layer0_outputs[8486] = (inputs[21]) | (inputs[25]);
    assign layer0_outputs[8487] = ~(inputs[5]) | (inputs[172]);
    assign layer0_outputs[8488] = ~(inputs[176]);
    assign layer0_outputs[8489] = ~(inputs[230]) | (inputs[61]);
    assign layer0_outputs[8490] = ~(inputs[8]) | (inputs[223]);
    assign layer0_outputs[8491] = (inputs[64]) | (inputs[38]);
    assign layer0_outputs[8492] = ~(inputs[154]) | (inputs[101]);
    assign layer0_outputs[8493] = ~((inputs[27]) ^ (inputs[238]));
    assign layer0_outputs[8494] = inputs[50];
    assign layer0_outputs[8495] = ~((inputs[166]) | (inputs[30]));
    assign layer0_outputs[8496] = (inputs[252]) ^ (inputs[8]);
    assign layer0_outputs[8497] = (inputs[44]) & (inputs[117]);
    assign layer0_outputs[8498] = (inputs[136]) | (inputs[117]);
    assign layer0_outputs[8499] = inputs[155];
    assign layer0_outputs[8500] = (inputs[30]) | (inputs[27]);
    assign layer0_outputs[8501] = ~(inputs[120]);
    assign layer0_outputs[8502] = (inputs[28]) | (inputs[111]);
    assign layer0_outputs[8503] = (inputs[171]) ^ (inputs[133]);
    assign layer0_outputs[8504] = (inputs[187]) | (inputs[46]);
    assign layer0_outputs[8505] = ~(inputs[111]) | (inputs[220]);
    assign layer0_outputs[8506] = (inputs[212]) | (inputs[194]);
    assign layer0_outputs[8507] = inputs[118];
    assign layer0_outputs[8508] = ~(inputs[248]);
    assign layer0_outputs[8509] = (inputs[166]) & ~(inputs[160]);
    assign layer0_outputs[8510] = inputs[37];
    assign layer0_outputs[8511] = (inputs[186]) & ~(inputs[105]);
    assign layer0_outputs[8512] = (inputs[8]) & ~(inputs[241]);
    assign layer0_outputs[8513] = inputs[166];
    assign layer0_outputs[8514] = ~((inputs[119]) ^ (inputs[184]));
    assign layer0_outputs[8515] = inputs[181];
    assign layer0_outputs[8516] = ~(inputs[207]) | (inputs[15]);
    assign layer0_outputs[8517] = ~((inputs[38]) | (inputs[16]));
    assign layer0_outputs[8518] = inputs[141];
    assign layer0_outputs[8519] = (inputs[147]) & ~(inputs[107]);
    assign layer0_outputs[8520] = inputs[4];
    assign layer0_outputs[8521] = inputs[201];
    assign layer0_outputs[8522] = ~((inputs[169]) | (inputs[138]));
    assign layer0_outputs[8523] = inputs[91];
    assign layer0_outputs[8524] = 1'b1;
    assign layer0_outputs[8525] = (inputs[150]) | (inputs[238]);
    assign layer0_outputs[8526] = ~((inputs[42]) | (inputs[79]));
    assign layer0_outputs[8527] = ~((inputs[241]) | (inputs[175]));
    assign layer0_outputs[8528] = ~((inputs[87]) & (inputs[221]));
    assign layer0_outputs[8529] = (inputs[165]) & ~(inputs[16]);
    assign layer0_outputs[8530] = ~(inputs[235]);
    assign layer0_outputs[8531] = ~(inputs[219]);
    assign layer0_outputs[8532] = ~((inputs[83]) | (inputs[10]));
    assign layer0_outputs[8533] = inputs[188];
    assign layer0_outputs[8534] = inputs[54];
    assign layer0_outputs[8535] = ~(inputs[77]) | (inputs[220]);
    assign layer0_outputs[8536] = (inputs[45]) | (inputs[69]);
    assign layer0_outputs[8537] = ~(inputs[238]);
    assign layer0_outputs[8538] = (inputs[24]) & (inputs[248]);
    assign layer0_outputs[8539] = (inputs[255]) | (inputs[230]);
    assign layer0_outputs[8540] = ~(inputs[121]) | (inputs[163]);
    assign layer0_outputs[8541] = ~(inputs[1]);
    assign layer0_outputs[8542] = ~(inputs[7]);
    assign layer0_outputs[8543] = ~(inputs[135]);
    assign layer0_outputs[8544] = (inputs[189]) & ~(inputs[242]);
    assign layer0_outputs[8545] = ~((inputs[120]) ^ (inputs[121]));
    assign layer0_outputs[8546] = inputs[41];
    assign layer0_outputs[8547] = (inputs[101]) & ~(inputs[244]);
    assign layer0_outputs[8548] = ~(inputs[198]);
    assign layer0_outputs[8549] = ~(inputs[24]) | (inputs[115]);
    assign layer0_outputs[8550] = ~((inputs[69]) ^ (inputs[20]));
    assign layer0_outputs[8551] = ~(inputs[42]) | (inputs[221]);
    assign layer0_outputs[8552] = ~(inputs[22]);
    assign layer0_outputs[8553] = (inputs[146]) & ~(inputs[235]);
    assign layer0_outputs[8554] = inputs[24];
    assign layer0_outputs[8555] = ~(inputs[106]) | (inputs[193]);
    assign layer0_outputs[8556] = (inputs[227]) & ~(inputs[155]);
    assign layer0_outputs[8557] = ~(inputs[108]);
    assign layer0_outputs[8558] = (inputs[54]) | (inputs[226]);
    assign layer0_outputs[8559] = inputs[36];
    assign layer0_outputs[8560] = ~(inputs[197]);
    assign layer0_outputs[8561] = ~(inputs[142]) | (inputs[93]);
    assign layer0_outputs[8562] = inputs[234];
    assign layer0_outputs[8563] = (inputs[208]) ^ (inputs[98]);
    assign layer0_outputs[8564] = (inputs[108]) & ~(inputs[248]);
    assign layer0_outputs[8565] = ~(inputs[113]) | (inputs[64]);
    assign layer0_outputs[8566] = ~(inputs[74]);
    assign layer0_outputs[8567] = inputs[148];
    assign layer0_outputs[8568] = inputs[222];
    assign layer0_outputs[8569] = (inputs[193]) & ~(inputs[73]);
    assign layer0_outputs[8570] = inputs[221];
    assign layer0_outputs[8571] = ~((inputs[102]) ^ (inputs[165]));
    assign layer0_outputs[8572] = (inputs[194]) & ~(inputs[100]);
    assign layer0_outputs[8573] = inputs[39];
    assign layer0_outputs[8574] = ~((inputs[204]) ^ (inputs[16]));
    assign layer0_outputs[8575] = ~(inputs[151]);
    assign layer0_outputs[8576] = (inputs[103]) ^ (inputs[135]);
    assign layer0_outputs[8577] = (inputs[215]) & (inputs[215]);
    assign layer0_outputs[8578] = 1'b1;
    assign layer0_outputs[8579] = ~((inputs[253]) | (inputs[236]));
    assign layer0_outputs[8580] = inputs[52];
    assign layer0_outputs[8581] = (inputs[236]) | (inputs[244]);
    assign layer0_outputs[8582] = ~((inputs[199]) | (inputs[183]));
    assign layer0_outputs[8583] = inputs[190];
    assign layer0_outputs[8584] = inputs[211];
    assign layer0_outputs[8585] = (inputs[227]) & ~(inputs[17]);
    assign layer0_outputs[8586] = (inputs[180]) & ~(inputs[29]);
    assign layer0_outputs[8587] = inputs[114];
    assign layer0_outputs[8588] = ~((inputs[7]) ^ (inputs[214]));
    assign layer0_outputs[8589] = ~(inputs[118]);
    assign layer0_outputs[8590] = ~(inputs[121]);
    assign layer0_outputs[8591] = (inputs[156]) | (inputs[205]);
    assign layer0_outputs[8592] = (inputs[157]) | (inputs[86]);
    assign layer0_outputs[8593] = inputs[131];
    assign layer0_outputs[8594] = ~((inputs[170]) ^ (inputs[94]));
    assign layer0_outputs[8595] = (inputs[131]) & (inputs[196]);
    assign layer0_outputs[8596] = (inputs[101]) ^ (inputs[71]);
    assign layer0_outputs[8597] = ~(inputs[189]);
    assign layer0_outputs[8598] = ~(inputs[220]) | (inputs[59]);
    assign layer0_outputs[8599] = 1'b1;
    assign layer0_outputs[8600] = ~((inputs[174]) ^ (inputs[123]));
    assign layer0_outputs[8601] = ~((inputs[99]) ^ (inputs[71]));
    assign layer0_outputs[8602] = ~(inputs[111]);
    assign layer0_outputs[8603] = ~(inputs[254]);
    assign layer0_outputs[8604] = (inputs[119]) & ~(inputs[235]);
    assign layer0_outputs[8605] = ~((inputs[244]) & (inputs[12]));
    assign layer0_outputs[8606] = (inputs[47]) & ~(inputs[16]);
    assign layer0_outputs[8607] = inputs[77];
    assign layer0_outputs[8608] = ~((inputs[184]) ^ (inputs[158]));
    assign layer0_outputs[8609] = ~(inputs[39]);
    assign layer0_outputs[8610] = ~(inputs[43]) | (inputs[254]);
    assign layer0_outputs[8611] = ~(inputs[85]);
    assign layer0_outputs[8612] = inputs[230];
    assign layer0_outputs[8613] = ~((inputs[89]) | (inputs[45]));
    assign layer0_outputs[8614] = ~((inputs[8]) | (inputs[231]));
    assign layer0_outputs[8615] = ~(inputs[136]);
    assign layer0_outputs[8616] = (inputs[19]) & ~(inputs[140]);
    assign layer0_outputs[8617] = (inputs[179]) & ~(inputs[4]);
    assign layer0_outputs[8618] = (inputs[233]) & (inputs[135]);
    assign layer0_outputs[8619] = (inputs[11]) | (inputs[12]);
    assign layer0_outputs[8620] = inputs[214];
    assign layer0_outputs[8621] = ~(inputs[117]);
    assign layer0_outputs[8622] = (inputs[185]) & ~(inputs[126]);
    assign layer0_outputs[8623] = inputs[198];
    assign layer0_outputs[8624] = 1'b0;
    assign layer0_outputs[8625] = (inputs[43]) | (inputs[114]);
    assign layer0_outputs[8626] = inputs[132];
    assign layer0_outputs[8627] = ~((inputs[102]) | (inputs[244]));
    assign layer0_outputs[8628] = inputs[21];
    assign layer0_outputs[8629] = ~(inputs[78]);
    assign layer0_outputs[8630] = (inputs[173]) ^ (inputs[71]);
    assign layer0_outputs[8631] = ~((inputs[11]) & (inputs[173]));
    assign layer0_outputs[8632] = ~(inputs[140]) | (inputs[191]);
    assign layer0_outputs[8633] = ~((inputs[165]) | (inputs[90]));
    assign layer0_outputs[8634] = (inputs[52]) | (inputs[6]);
    assign layer0_outputs[8635] = ~(inputs[230]) | (inputs[238]);
    assign layer0_outputs[8636] = ~((inputs[91]) & (inputs[8]));
    assign layer0_outputs[8637] = ~(inputs[222]);
    assign layer0_outputs[8638] = (inputs[88]) & (inputs[14]);
    assign layer0_outputs[8639] = (inputs[106]) | (inputs[123]);
    assign layer0_outputs[8640] = (inputs[214]) | (inputs[139]);
    assign layer0_outputs[8641] = ~(inputs[160]);
    assign layer0_outputs[8642] = (inputs[66]) | (inputs[30]);
    assign layer0_outputs[8643] = (inputs[151]) | (inputs[206]);
    assign layer0_outputs[8644] = (inputs[177]) & (inputs[151]);
    assign layer0_outputs[8645] = (inputs[50]) ^ (inputs[75]);
    assign layer0_outputs[8646] = (inputs[53]) | (inputs[7]);
    assign layer0_outputs[8647] = (inputs[178]) ^ (inputs[58]);
    assign layer0_outputs[8648] = (inputs[189]) & (inputs[219]);
    assign layer0_outputs[8649] = ~(inputs[59]);
    assign layer0_outputs[8650] = ~(inputs[155]);
    assign layer0_outputs[8651] = ~(inputs[99]) | (inputs[41]);
    assign layer0_outputs[8652] = (inputs[169]) & ~(inputs[39]);
    assign layer0_outputs[8653] = inputs[213];
    assign layer0_outputs[8654] = ~((inputs[70]) ^ (inputs[177]));
    assign layer0_outputs[8655] = ~(inputs[45]);
    assign layer0_outputs[8656] = ~((inputs[193]) | (inputs[63]));
    assign layer0_outputs[8657] = ~(inputs[200]) | (inputs[31]);
    assign layer0_outputs[8658] = (inputs[23]) & (inputs[25]);
    assign layer0_outputs[8659] = ~((inputs[5]) | (inputs[1]));
    assign layer0_outputs[8660] = ~(inputs[134]);
    assign layer0_outputs[8661] = ~((inputs[107]) ^ (inputs[86]));
    assign layer0_outputs[8662] = (inputs[86]) ^ (inputs[107]);
    assign layer0_outputs[8663] = inputs[172];
    assign layer0_outputs[8664] = ~(inputs[202]) | (inputs[32]);
    assign layer0_outputs[8665] = (inputs[147]) & ~(inputs[46]);
    assign layer0_outputs[8666] = ~((inputs[17]) | (inputs[227]));
    assign layer0_outputs[8667] = (inputs[128]) | (inputs[99]);
    assign layer0_outputs[8668] = 1'b1;
    assign layer0_outputs[8669] = ~(inputs[190]);
    assign layer0_outputs[8670] = ~(inputs[245]) | (inputs[68]);
    assign layer0_outputs[8671] = (inputs[105]) & ~(inputs[20]);
    assign layer0_outputs[8672] = inputs[115];
    assign layer0_outputs[8673] = inputs[127];
    assign layer0_outputs[8674] = ~(inputs[156]);
    assign layer0_outputs[8675] = inputs[9];
    assign layer0_outputs[8676] = (inputs[47]) & ~(inputs[207]);
    assign layer0_outputs[8677] = (inputs[250]) & (inputs[146]);
    assign layer0_outputs[8678] = inputs[197];
    assign layer0_outputs[8679] = inputs[182];
    assign layer0_outputs[8680] = (inputs[99]) & ~(inputs[54]);
    assign layer0_outputs[8681] = (inputs[18]) | (inputs[74]);
    assign layer0_outputs[8682] = inputs[102];
    assign layer0_outputs[8683] = ~(inputs[73]) | (inputs[156]);
    assign layer0_outputs[8684] = inputs[130];
    assign layer0_outputs[8685] = ~(inputs[71]) | (inputs[246]);
    assign layer0_outputs[8686] = 1'b0;
    assign layer0_outputs[8687] = (inputs[247]) | (inputs[111]);
    assign layer0_outputs[8688] = ~(inputs[44]) | (inputs[8]);
    assign layer0_outputs[8689] = ~(inputs[38]) | (inputs[223]);
    assign layer0_outputs[8690] = (inputs[135]) & ~(inputs[191]);
    assign layer0_outputs[8691] = inputs[49];
    assign layer0_outputs[8692] = (inputs[70]) & ~(inputs[246]);
    assign layer0_outputs[8693] = (inputs[130]) & (inputs[70]);
    assign layer0_outputs[8694] = (inputs[211]) & ~(inputs[236]);
    assign layer0_outputs[8695] = inputs[149];
    assign layer0_outputs[8696] = inputs[131];
    assign layer0_outputs[8697] = ~((inputs[232]) | (inputs[2]));
    assign layer0_outputs[8698] = (inputs[112]) & ~(inputs[126]);
    assign layer0_outputs[8699] = (inputs[80]) & ~(inputs[218]);
    assign layer0_outputs[8700] = ~((inputs[167]) & (inputs[44]));
    assign layer0_outputs[8701] = (inputs[221]) & ~(inputs[158]);
    assign layer0_outputs[8702] = 1'b0;
    assign layer0_outputs[8703] = ~((inputs[148]) | (inputs[22]));
    assign layer0_outputs[8704] = inputs[56];
    assign layer0_outputs[8705] = inputs[102];
    assign layer0_outputs[8706] = ~(inputs[135]);
    assign layer0_outputs[8707] = inputs[192];
    assign layer0_outputs[8708] = (inputs[238]) & (inputs[61]);
    assign layer0_outputs[8709] = ~(inputs[77]);
    assign layer0_outputs[8710] = (inputs[204]) ^ (inputs[101]);
    assign layer0_outputs[8711] = ~(inputs[249]);
    assign layer0_outputs[8712] = (inputs[46]) | (inputs[128]);
    assign layer0_outputs[8713] = (inputs[93]) & ~(inputs[194]);
    assign layer0_outputs[8714] = inputs[109];
    assign layer0_outputs[8715] = ~((inputs[153]) | (inputs[148]));
    assign layer0_outputs[8716] = 1'b1;
    assign layer0_outputs[8717] = ~((inputs[0]) & (inputs[146]));
    assign layer0_outputs[8718] = ~(inputs[214]);
    assign layer0_outputs[8719] = inputs[141];
    assign layer0_outputs[8720] = (inputs[231]) & ~(inputs[237]);
    assign layer0_outputs[8721] = ~(inputs[65]) | (inputs[184]);
    assign layer0_outputs[8722] = ~(inputs[103]);
    assign layer0_outputs[8723] = ~(inputs[124]);
    assign layer0_outputs[8724] = ~((inputs[220]) ^ (inputs[4]));
    assign layer0_outputs[8725] = (inputs[22]) & ~(inputs[146]);
    assign layer0_outputs[8726] = (inputs[164]) ^ (inputs[147]);
    assign layer0_outputs[8727] = ~((inputs[107]) | (inputs[61]));
    assign layer0_outputs[8728] = ~(inputs[236]);
    assign layer0_outputs[8729] = 1'b0;
    assign layer0_outputs[8730] = ~(inputs[72]);
    assign layer0_outputs[8731] = ~(inputs[93]);
    assign layer0_outputs[8732] = ~(inputs[11]);
    assign layer0_outputs[8733] = (inputs[51]) ^ (inputs[147]);
    assign layer0_outputs[8734] = inputs[245];
    assign layer0_outputs[8735] = (inputs[250]) | (inputs[55]);
    assign layer0_outputs[8736] = ~((inputs[147]) | (inputs[144]));
    assign layer0_outputs[8737] = ~((inputs[240]) & (inputs[18]));
    assign layer0_outputs[8738] = ~(inputs[173]);
    assign layer0_outputs[8739] = ~(inputs[133]) | (inputs[34]);
    assign layer0_outputs[8740] = (inputs[46]) | (inputs[114]);
    assign layer0_outputs[8741] = ~(inputs[75]);
    assign layer0_outputs[8742] = ~(inputs[23]);
    assign layer0_outputs[8743] = ~((inputs[251]) | (inputs[218]));
    assign layer0_outputs[8744] = (inputs[80]) | (inputs[196]);
    assign layer0_outputs[8745] = ~((inputs[106]) & (inputs[198]));
    assign layer0_outputs[8746] = ~(inputs[235]) | (inputs[78]);
    assign layer0_outputs[8747] = ~(inputs[159]);
    assign layer0_outputs[8748] = ~(inputs[251]) | (inputs[38]);
    assign layer0_outputs[8749] = inputs[62];
    assign layer0_outputs[8750] = (inputs[204]) | (inputs[37]);
    assign layer0_outputs[8751] = 1'b0;
    assign layer0_outputs[8752] = ~(inputs[119]);
    assign layer0_outputs[8753] = ~(inputs[214]);
    assign layer0_outputs[8754] = (inputs[6]) | (inputs[242]);
    assign layer0_outputs[8755] = (inputs[216]) | (inputs[55]);
    assign layer0_outputs[8756] = ~((inputs[110]) ^ (inputs[21]));
    assign layer0_outputs[8757] = ~(inputs[67]) | (inputs[225]);
    assign layer0_outputs[8758] = inputs[42];
    assign layer0_outputs[8759] = (inputs[197]) & ~(inputs[1]);
    assign layer0_outputs[8760] = ~(inputs[99]);
    assign layer0_outputs[8761] = (inputs[23]) ^ (inputs[106]);
    assign layer0_outputs[8762] = ~(inputs[26]);
    assign layer0_outputs[8763] = ~((inputs[225]) | (inputs[18]));
    assign layer0_outputs[8764] = (inputs[202]) & (inputs[78]);
    assign layer0_outputs[8765] = (inputs[254]) & ~(inputs[52]);
    assign layer0_outputs[8766] = (inputs[166]) & ~(inputs[188]);
    assign layer0_outputs[8767] = inputs[164];
    assign layer0_outputs[8768] = (inputs[215]) | (inputs[119]);
    assign layer0_outputs[8769] = ~(inputs[22]);
    assign layer0_outputs[8770] = ~((inputs[123]) | (inputs[73]));
    assign layer0_outputs[8771] = ~((inputs[213]) & (inputs[190]));
    assign layer0_outputs[8772] = ~((inputs[235]) | (inputs[210]));
    assign layer0_outputs[8773] = inputs[121];
    assign layer0_outputs[8774] = ~(inputs[248]) | (inputs[20]);
    assign layer0_outputs[8775] = (inputs[141]) & ~(inputs[154]);
    assign layer0_outputs[8776] = (inputs[201]) & ~(inputs[196]);
    assign layer0_outputs[8777] = inputs[231];
    assign layer0_outputs[8778] = (inputs[64]) ^ (inputs[114]);
    assign layer0_outputs[8779] = ~(inputs[126]);
    assign layer0_outputs[8780] = ~((inputs[49]) & (inputs[118]));
    assign layer0_outputs[8781] = (inputs[170]) | (inputs[185]);
    assign layer0_outputs[8782] = ~(inputs[22]) | (inputs[196]);
    assign layer0_outputs[8783] = ~(inputs[151]);
    assign layer0_outputs[8784] = ~(inputs[95]) | (inputs[250]);
    assign layer0_outputs[8785] = (inputs[18]) & ~(inputs[66]);
    assign layer0_outputs[8786] = inputs[78];
    assign layer0_outputs[8787] = (inputs[81]) | (inputs[114]);
    assign layer0_outputs[8788] = (inputs[100]) | (inputs[189]);
    assign layer0_outputs[8789] = (inputs[47]) | (inputs[27]);
    assign layer0_outputs[8790] = (inputs[114]) | (inputs[238]);
    assign layer0_outputs[8791] = ~((inputs[53]) ^ (inputs[22]));
    assign layer0_outputs[8792] = ~(inputs[162]);
    assign layer0_outputs[8793] = ~(inputs[138]) | (inputs[93]);
    assign layer0_outputs[8794] = ~((inputs[83]) | (inputs[219]));
    assign layer0_outputs[8795] = ~((inputs[210]) ^ (inputs[180]));
    assign layer0_outputs[8796] = ~(inputs[104]);
    assign layer0_outputs[8797] = (inputs[238]) | (inputs[72]);
    assign layer0_outputs[8798] = ~((inputs[161]) | (inputs[126]));
    assign layer0_outputs[8799] = (inputs[146]) | (inputs[68]);
    assign layer0_outputs[8800] = (inputs[255]) | (inputs[18]);
    assign layer0_outputs[8801] = (inputs[183]) & ~(inputs[173]);
    assign layer0_outputs[8802] = (inputs[20]) & ~(inputs[176]);
    assign layer0_outputs[8803] = (inputs[68]) & ~(inputs[3]);
    assign layer0_outputs[8804] = (inputs[199]) & (inputs[201]);
    assign layer0_outputs[8805] = (inputs[129]) | (inputs[34]);
    assign layer0_outputs[8806] = inputs[237];
    assign layer0_outputs[8807] = ~((inputs[20]) ^ (inputs[81]));
    assign layer0_outputs[8808] = inputs[106];
    assign layer0_outputs[8809] = ~((inputs[62]) ^ (inputs[44]));
    assign layer0_outputs[8810] = inputs[251];
    assign layer0_outputs[8811] = inputs[12];
    assign layer0_outputs[8812] = (inputs[194]) & ~(inputs[136]);
    assign layer0_outputs[8813] = ~(inputs[217]);
    assign layer0_outputs[8814] = ~(inputs[82]);
    assign layer0_outputs[8815] = ~(inputs[24]);
    assign layer0_outputs[8816] = ~((inputs[14]) & (inputs[117]));
    assign layer0_outputs[8817] = ~((inputs[231]) ^ (inputs[21]));
    assign layer0_outputs[8818] = (inputs[30]) | (inputs[69]);
    assign layer0_outputs[8819] = (inputs[133]) & (inputs[65]);
    assign layer0_outputs[8820] = inputs[57];
    assign layer0_outputs[8821] = ~(inputs[11]);
    assign layer0_outputs[8822] = ~((inputs[84]) ^ (inputs[218]));
    assign layer0_outputs[8823] = inputs[159];
    assign layer0_outputs[8824] = 1'b1;
    assign layer0_outputs[8825] = ~(inputs[133]);
    assign layer0_outputs[8826] = ~((inputs[34]) ^ (inputs[125]));
    assign layer0_outputs[8827] = (inputs[78]) ^ (inputs[6]);
    assign layer0_outputs[8828] = (inputs[3]) | (inputs[57]);
    assign layer0_outputs[8829] = ~(inputs[164]);
    assign layer0_outputs[8830] = ~((inputs[232]) ^ (inputs[246]));
    assign layer0_outputs[8831] = ~(inputs[54]);
    assign layer0_outputs[8832] = (inputs[144]) ^ (inputs[194]);
    assign layer0_outputs[8833] = ~(inputs[132]);
    assign layer0_outputs[8834] = ~(inputs[133]) | (inputs[29]);
    assign layer0_outputs[8835] = ~((inputs[170]) ^ (inputs[238]));
    assign layer0_outputs[8836] = ~(inputs[171]);
    assign layer0_outputs[8837] = 1'b1;
    assign layer0_outputs[8838] = ~((inputs[157]) ^ (inputs[119]));
    assign layer0_outputs[8839] = inputs[6];
    assign layer0_outputs[8840] = inputs[210];
    assign layer0_outputs[8841] = inputs[93];
    assign layer0_outputs[8842] = ~(inputs[171]) | (inputs[31]);
    assign layer0_outputs[8843] = (inputs[106]) & ~(inputs[153]);
    assign layer0_outputs[8844] = ~(inputs[28]) | (inputs[125]);
    assign layer0_outputs[8845] = 1'b0;
    assign layer0_outputs[8846] = ~((inputs[241]) ^ (inputs[156]));
    assign layer0_outputs[8847] = ~(inputs[169]);
    assign layer0_outputs[8848] = ~((inputs[31]) | (inputs[108]));
    assign layer0_outputs[8849] = inputs[9];
    assign layer0_outputs[8850] = 1'b1;
    assign layer0_outputs[8851] = ~(inputs[201]);
    assign layer0_outputs[8852] = ~(inputs[210]) | (inputs[146]);
    assign layer0_outputs[8853] = (inputs[17]) & (inputs[227]);
    assign layer0_outputs[8854] = ~((inputs[174]) | (inputs[193]));
    assign layer0_outputs[8855] = ~(inputs[233]) | (inputs[127]);
    assign layer0_outputs[8856] = ~(inputs[195]) | (inputs[113]);
    assign layer0_outputs[8857] = inputs[43];
    assign layer0_outputs[8858] = (inputs[106]) & ~(inputs[184]);
    assign layer0_outputs[8859] = inputs[122];
    assign layer0_outputs[8860] = (inputs[158]) ^ (inputs[185]);
    assign layer0_outputs[8861] = (inputs[205]) & ~(inputs[243]);
    assign layer0_outputs[8862] = ~((inputs[115]) ^ (inputs[128]));
    assign layer0_outputs[8863] = ~((inputs[192]) | (inputs[133]));
    assign layer0_outputs[8864] = (inputs[229]) & ~(inputs[223]);
    assign layer0_outputs[8865] = inputs[249];
    assign layer0_outputs[8866] = ~(inputs[176]) | (inputs[36]);
    assign layer0_outputs[8867] = (inputs[217]) | (inputs[67]);
    assign layer0_outputs[8868] = (inputs[98]) & ~(inputs[110]);
    assign layer0_outputs[8869] = inputs[242];
    assign layer0_outputs[8870] = ~((inputs[136]) | (inputs[225]));
    assign layer0_outputs[8871] = ~((inputs[9]) ^ (inputs[207]));
    assign layer0_outputs[8872] = (inputs[50]) & (inputs[62]);
    assign layer0_outputs[8873] = inputs[202];
    assign layer0_outputs[8874] = (inputs[75]) & (inputs[106]);
    assign layer0_outputs[8875] = inputs[76];
    assign layer0_outputs[8876] = (inputs[183]) & ~(inputs[83]);
    assign layer0_outputs[8877] = ~((inputs[197]) ^ (inputs[10]));
    assign layer0_outputs[8878] = ~((inputs[214]) | (inputs[181]));
    assign layer0_outputs[8879] = ~(inputs[185]);
    assign layer0_outputs[8880] = (inputs[241]) & ~(inputs[214]);
    assign layer0_outputs[8881] = ~(inputs[193]);
    assign layer0_outputs[8882] = ~((inputs[242]) & (inputs[55]));
    assign layer0_outputs[8883] = (inputs[89]) | (inputs[4]);
    assign layer0_outputs[8884] = ~(inputs[210]);
    assign layer0_outputs[8885] = ~(inputs[13]) | (inputs[90]);
    assign layer0_outputs[8886] = ~(inputs[47]);
    assign layer0_outputs[8887] = ~((inputs[37]) ^ (inputs[43]));
    assign layer0_outputs[8888] = ~(inputs[233]);
    assign layer0_outputs[8889] = ~((inputs[118]) ^ (inputs[116]));
    assign layer0_outputs[8890] = (inputs[233]) & ~(inputs[150]);
    assign layer0_outputs[8891] = 1'b1;
    assign layer0_outputs[8892] = 1'b1;
    assign layer0_outputs[8893] = ~(inputs[222]);
    assign layer0_outputs[8894] = ~(inputs[33]) | (inputs[65]);
    assign layer0_outputs[8895] = inputs[165];
    assign layer0_outputs[8896] = ~((inputs[139]) ^ (inputs[101]));
    assign layer0_outputs[8897] = (inputs[4]) | (inputs[64]);
    assign layer0_outputs[8898] = ~(inputs[100]);
    assign layer0_outputs[8899] = (inputs[149]) & ~(inputs[38]);
    assign layer0_outputs[8900] = inputs[150];
    assign layer0_outputs[8901] = ~(inputs[78]);
    assign layer0_outputs[8902] = inputs[107];
    assign layer0_outputs[8903] = 1'b0;
    assign layer0_outputs[8904] = (inputs[45]) & ~(inputs[137]);
    assign layer0_outputs[8905] = (inputs[219]) & (inputs[182]);
    assign layer0_outputs[8906] = ~(inputs[174]) | (inputs[153]);
    assign layer0_outputs[8907] = ~((inputs[253]) | (inputs[134]));
    assign layer0_outputs[8908] = ~((inputs[247]) & (inputs[227]));
    assign layer0_outputs[8909] = ~(inputs[24]);
    assign layer0_outputs[8910] = 1'b1;
    assign layer0_outputs[8911] = (inputs[159]) & ~(inputs[215]);
    assign layer0_outputs[8912] = ~((inputs[249]) | (inputs[254]));
    assign layer0_outputs[8913] = ~(inputs[45]);
    assign layer0_outputs[8914] = 1'b0;
    assign layer0_outputs[8915] = ~((inputs[232]) | (inputs[190]));
    assign layer0_outputs[8916] = ~(inputs[181]);
    assign layer0_outputs[8917] = inputs[119];
    assign layer0_outputs[8918] = ~(inputs[197]);
    assign layer0_outputs[8919] = 1'b1;
    assign layer0_outputs[8920] = (inputs[146]) | (inputs[50]);
    assign layer0_outputs[8921] = ~(inputs[37]);
    assign layer0_outputs[8922] = inputs[140];
    assign layer0_outputs[8923] = ~(inputs[193]) | (inputs[39]);
    assign layer0_outputs[8924] = ~(inputs[28]) | (inputs[253]);
    assign layer0_outputs[8925] = (inputs[154]) & ~(inputs[3]);
    assign layer0_outputs[8926] = (inputs[121]) & ~(inputs[93]);
    assign layer0_outputs[8927] = ~(inputs[229]);
    assign layer0_outputs[8928] = inputs[58];
    assign layer0_outputs[8929] = ~((inputs[39]) | (inputs[47]));
    assign layer0_outputs[8930] = (inputs[254]) & ~(inputs[220]);
    assign layer0_outputs[8931] = ~(inputs[136]);
    assign layer0_outputs[8932] = (inputs[148]) | (inputs[87]);
    assign layer0_outputs[8933] = ~(inputs[123]) | (inputs[59]);
    assign layer0_outputs[8934] = ~(inputs[207]);
    assign layer0_outputs[8935] = inputs[25];
    assign layer0_outputs[8936] = inputs[100];
    assign layer0_outputs[8937] = ~((inputs[159]) | (inputs[32]));
    assign layer0_outputs[8938] = (inputs[109]) & ~(inputs[239]);
    assign layer0_outputs[8939] = ~((inputs[53]) & (inputs[59]));
    assign layer0_outputs[8940] = (inputs[197]) & ~(inputs[190]);
    assign layer0_outputs[8941] = ~(inputs[35]);
    assign layer0_outputs[8942] = inputs[98];
    assign layer0_outputs[8943] = inputs[219];
    assign layer0_outputs[8944] = inputs[114];
    assign layer0_outputs[8945] = ~(inputs[252]);
    assign layer0_outputs[8946] = inputs[245];
    assign layer0_outputs[8947] = ~(inputs[88]) | (inputs[34]);
    assign layer0_outputs[8948] = ~(inputs[24]) | (inputs[97]);
    assign layer0_outputs[8949] = ~(inputs[129]);
    assign layer0_outputs[8950] = inputs[250];
    assign layer0_outputs[8951] = ~((inputs[145]) ^ (inputs[132]));
    assign layer0_outputs[8952] = inputs[247];
    assign layer0_outputs[8953] = ~((inputs[85]) & (inputs[85]));
    assign layer0_outputs[8954] = (inputs[85]) & (inputs[84]);
    assign layer0_outputs[8955] = ~(inputs[49]);
    assign layer0_outputs[8956] = (inputs[253]) | (inputs[254]);
    assign layer0_outputs[8957] = inputs[115];
    assign layer0_outputs[8958] = (inputs[91]) & ~(inputs[57]);
    assign layer0_outputs[8959] = (inputs[191]) ^ (inputs[108]);
    assign layer0_outputs[8960] = 1'b1;
    assign layer0_outputs[8961] = inputs[58];
    assign layer0_outputs[8962] = ~(inputs[93]);
    assign layer0_outputs[8963] = inputs[247];
    assign layer0_outputs[8964] = ~((inputs[170]) & (inputs[76]));
    assign layer0_outputs[8965] = ~(inputs[186]);
    assign layer0_outputs[8966] = ~((inputs[225]) | (inputs[63]));
    assign layer0_outputs[8967] = inputs[90];
    assign layer0_outputs[8968] = inputs[73];
    assign layer0_outputs[8969] = (inputs[70]) & ~(inputs[191]);
    assign layer0_outputs[8970] = (inputs[78]) | (inputs[45]);
    assign layer0_outputs[8971] = ~(inputs[212]);
    assign layer0_outputs[8972] = 1'b0;
    assign layer0_outputs[8973] = ~(inputs[171]);
    assign layer0_outputs[8974] = (inputs[79]) ^ (inputs[222]);
    assign layer0_outputs[8975] = ~(inputs[61]);
    assign layer0_outputs[8976] = ~(inputs[146]);
    assign layer0_outputs[8977] = ~(inputs[160]);
    assign layer0_outputs[8978] = inputs[167];
    assign layer0_outputs[8979] = ~(inputs[29]);
    assign layer0_outputs[8980] = ~(inputs[120]);
    assign layer0_outputs[8981] = (inputs[161]) | (inputs[222]);
    assign layer0_outputs[8982] = ~((inputs[88]) ^ (inputs[93]));
    assign layer0_outputs[8983] = ~(inputs[147]);
    assign layer0_outputs[8984] = ~(inputs[102]);
    assign layer0_outputs[8985] = (inputs[191]) & (inputs[32]);
    assign layer0_outputs[8986] = 1'b1;
    assign layer0_outputs[8987] = (inputs[186]) ^ (inputs[177]);
    assign layer0_outputs[8988] = ~((inputs[164]) ^ (inputs[176]));
    assign layer0_outputs[8989] = inputs[123];
    assign layer0_outputs[8990] = (inputs[22]) & ~(inputs[115]);
    assign layer0_outputs[8991] = ~(inputs[146]) | (inputs[220]);
    assign layer0_outputs[8992] = inputs[28];
    assign layer0_outputs[8993] = 1'b0;
    assign layer0_outputs[8994] = ~(inputs[11]) | (inputs[18]);
    assign layer0_outputs[8995] = inputs[117];
    assign layer0_outputs[8996] = ~((inputs[122]) ^ (inputs[110]));
    assign layer0_outputs[8997] = (inputs[85]) | (inputs[100]);
    assign layer0_outputs[8998] = (inputs[42]) & (inputs[66]);
    assign layer0_outputs[8999] = (inputs[91]) ^ (inputs[65]);
    assign layer0_outputs[9000] = (inputs[47]) ^ (inputs[105]);
    assign layer0_outputs[9001] = inputs[231];
    assign layer0_outputs[9002] = (inputs[13]) | (inputs[30]);
    assign layer0_outputs[9003] = (inputs[49]) ^ (inputs[123]);
    assign layer0_outputs[9004] = inputs[121];
    assign layer0_outputs[9005] = (inputs[236]) ^ (inputs[207]);
    assign layer0_outputs[9006] = ~((inputs[42]) | (inputs[79]));
    assign layer0_outputs[9007] = ~(inputs[243]) | (inputs[135]);
    assign layer0_outputs[9008] = ~((inputs[78]) & (inputs[88]));
    assign layer0_outputs[9009] = inputs[73];
    assign layer0_outputs[9010] = (inputs[158]) | (inputs[146]);
    assign layer0_outputs[9011] = ~((inputs[2]) | (inputs[183]));
    assign layer0_outputs[9012] = (inputs[203]) & (inputs[0]);
    assign layer0_outputs[9013] = ~(inputs[16]);
    assign layer0_outputs[9014] = (inputs[174]) | (inputs[160]);
    assign layer0_outputs[9015] = inputs[155];
    assign layer0_outputs[9016] = (inputs[41]) & ~(inputs[238]);
    assign layer0_outputs[9017] = (inputs[211]) & ~(inputs[88]);
    assign layer0_outputs[9018] = ~(inputs[121]);
    assign layer0_outputs[9019] = (inputs[64]) ^ (inputs[5]);
    assign layer0_outputs[9020] = (inputs[147]) | (inputs[124]);
    assign layer0_outputs[9021] = (inputs[228]) & ~(inputs[30]);
    assign layer0_outputs[9022] = ~((inputs[42]) | (inputs[6]));
    assign layer0_outputs[9023] = (inputs[76]) & ~(inputs[195]);
    assign layer0_outputs[9024] = inputs[176];
    assign layer0_outputs[9025] = (inputs[131]) | (inputs[53]);
    assign layer0_outputs[9026] = ~(inputs[110]);
    assign layer0_outputs[9027] = inputs[184];
    assign layer0_outputs[9028] = (inputs[128]) ^ (inputs[31]);
    assign layer0_outputs[9029] = 1'b1;
    assign layer0_outputs[9030] = ~(inputs[211]) | (inputs[95]);
    assign layer0_outputs[9031] = ~(inputs[166]);
    assign layer0_outputs[9032] = ~((inputs[48]) | (inputs[106]));
    assign layer0_outputs[9033] = (inputs[159]) & ~(inputs[145]);
    assign layer0_outputs[9034] = ~((inputs[178]) | (inputs[125]));
    assign layer0_outputs[9035] = ~(inputs[102]);
    assign layer0_outputs[9036] = 1'b1;
    assign layer0_outputs[9037] = inputs[74];
    assign layer0_outputs[9038] = (inputs[37]) ^ (inputs[252]);
    assign layer0_outputs[9039] = (inputs[26]) | (inputs[3]);
    assign layer0_outputs[9040] = ~(inputs[232]);
    assign layer0_outputs[9041] = ~((inputs[159]) & (inputs[40]));
    assign layer0_outputs[9042] = inputs[92];
    assign layer0_outputs[9043] = inputs[193];
    assign layer0_outputs[9044] = ~(inputs[130]);
    assign layer0_outputs[9045] = (inputs[141]) & ~(inputs[19]);
    assign layer0_outputs[9046] = inputs[193];
    assign layer0_outputs[9047] = (inputs[178]) ^ (inputs[219]);
    assign layer0_outputs[9048] = ~(inputs[13]) | (inputs[245]);
    assign layer0_outputs[9049] = (inputs[21]) & ~(inputs[207]);
    assign layer0_outputs[9050] = inputs[117];
    assign layer0_outputs[9051] = ~((inputs[108]) | (inputs[130]));
    assign layer0_outputs[9052] = (inputs[131]) & ~(inputs[241]);
    assign layer0_outputs[9053] = inputs[97];
    assign layer0_outputs[9054] = ~(inputs[146]);
    assign layer0_outputs[9055] = ~(inputs[148]);
    assign layer0_outputs[9056] = (inputs[229]) & ~(inputs[222]);
    assign layer0_outputs[9057] = ~(inputs[160]);
    assign layer0_outputs[9058] = ~((inputs[137]) | (inputs[59]));
    assign layer0_outputs[9059] = (inputs[141]) & (inputs[146]);
    assign layer0_outputs[9060] = inputs[68];
    assign layer0_outputs[9061] = ~((inputs[153]) ^ (inputs[94]));
    assign layer0_outputs[9062] = inputs[158];
    assign layer0_outputs[9063] = (inputs[176]) | (inputs[50]);
    assign layer0_outputs[9064] = ~((inputs[125]) | (inputs[49]));
    assign layer0_outputs[9065] = 1'b0;
    assign layer0_outputs[9066] = ~((inputs[229]) & (inputs[232]));
    assign layer0_outputs[9067] = ~((inputs[170]) | (inputs[236]));
    assign layer0_outputs[9068] = (inputs[88]) ^ (inputs[49]);
    assign layer0_outputs[9069] = (inputs[46]) | (inputs[66]);
    assign layer0_outputs[9070] = ~(inputs[23]) | (inputs[240]);
    assign layer0_outputs[9071] = inputs[203];
    assign layer0_outputs[9072] = ~(inputs[223]) | (inputs[36]);
    assign layer0_outputs[9073] = ~(inputs[70]);
    assign layer0_outputs[9074] = ~(inputs[177]) | (inputs[42]);
    assign layer0_outputs[9075] = ~((inputs[82]) | (inputs[54]));
    assign layer0_outputs[9076] = ~((inputs[49]) ^ (inputs[6]));
    assign layer0_outputs[9077] = (inputs[134]) & ~(inputs[237]);
    assign layer0_outputs[9078] = 1'b1;
    assign layer0_outputs[9079] = ~(inputs[212]) | (inputs[98]);
    assign layer0_outputs[9080] = ~(inputs[112]) | (inputs[31]);
    assign layer0_outputs[9081] = (inputs[59]) & (inputs[62]);
    assign layer0_outputs[9082] = ~((inputs[41]) | (inputs[190]));
    assign layer0_outputs[9083] = ~((inputs[175]) | (inputs[177]));
    assign layer0_outputs[9084] = ~((inputs[20]) | (inputs[89]));
    assign layer0_outputs[9085] = (inputs[206]) & ~(inputs[131]);
    assign layer0_outputs[9086] = inputs[127];
    assign layer0_outputs[9087] = 1'b0;
    assign layer0_outputs[9088] = ~(inputs[71]);
    assign layer0_outputs[9089] = inputs[248];
    assign layer0_outputs[9090] = ~(inputs[21]);
    assign layer0_outputs[9091] = ~(inputs[174]);
    assign layer0_outputs[9092] = (inputs[0]) ^ (inputs[62]);
    assign layer0_outputs[9093] = inputs[179];
    assign layer0_outputs[9094] = (inputs[188]) ^ (inputs[242]);
    assign layer0_outputs[9095] = (inputs[11]) & ~(inputs[201]);
    assign layer0_outputs[9096] = ~((inputs[201]) | (inputs[34]));
    assign layer0_outputs[9097] = inputs[169];
    assign layer0_outputs[9098] = (inputs[226]) & (inputs[44]);
    assign layer0_outputs[9099] = ~((inputs[249]) ^ (inputs[99]));
    assign layer0_outputs[9100] = ~(inputs[163]) | (inputs[31]);
    assign layer0_outputs[9101] = (inputs[241]) | (inputs[66]);
    assign layer0_outputs[9102] = ~(inputs[37]) | (inputs[153]);
    assign layer0_outputs[9103] = ~((inputs[62]) | (inputs[32]));
    assign layer0_outputs[9104] = ~(inputs[19]);
    assign layer0_outputs[9105] = ~(inputs[121]);
    assign layer0_outputs[9106] = (inputs[126]) & ~(inputs[154]);
    assign layer0_outputs[9107] = inputs[42];
    assign layer0_outputs[9108] = ~(inputs[105]);
    assign layer0_outputs[9109] = ~(inputs[233]) | (inputs[105]);
    assign layer0_outputs[9110] = ~(inputs[63]) | (inputs[16]);
    assign layer0_outputs[9111] = (inputs[180]) & ~(inputs[6]);
    assign layer0_outputs[9112] = inputs[128];
    assign layer0_outputs[9113] = (inputs[158]) | (inputs[176]);
    assign layer0_outputs[9114] = (inputs[108]) & (inputs[159]);
    assign layer0_outputs[9115] = ~(inputs[81]);
    assign layer0_outputs[9116] = inputs[117];
    assign layer0_outputs[9117] = (inputs[217]) ^ (inputs[192]);
    assign layer0_outputs[9118] = ~(inputs[118]);
    assign layer0_outputs[9119] = (inputs[22]) & ~(inputs[73]);
    assign layer0_outputs[9120] = (inputs[40]) & ~(inputs[217]);
    assign layer0_outputs[9121] = ~(inputs[73]) | (inputs[210]);
    assign layer0_outputs[9122] = (inputs[35]) & ~(inputs[125]);
    assign layer0_outputs[9123] = ~((inputs[145]) | (inputs[30]));
    assign layer0_outputs[9124] = (inputs[247]) | (inputs[228]);
    assign layer0_outputs[9125] = inputs[76];
    assign layer0_outputs[9126] = ~(inputs[127]);
    assign layer0_outputs[9127] = ~(inputs[190]);
    assign layer0_outputs[9128] = inputs[230];
    assign layer0_outputs[9129] = ~(inputs[13]) | (inputs[80]);
    assign layer0_outputs[9130] = ~(inputs[171]);
    assign layer0_outputs[9131] = ~((inputs[47]) | (inputs[32]));
    assign layer0_outputs[9132] = ~((inputs[211]) ^ (inputs[14]));
    assign layer0_outputs[9133] = ~((inputs[4]) | (inputs[35]));
    assign layer0_outputs[9134] = ~(inputs[234]);
    assign layer0_outputs[9135] = (inputs[39]) & ~(inputs[132]);
    assign layer0_outputs[9136] = (inputs[107]) | (inputs[30]);
    assign layer0_outputs[9137] = inputs[147];
    assign layer0_outputs[9138] = ~(inputs[84]);
    assign layer0_outputs[9139] = 1'b1;
    assign layer0_outputs[9140] = ~(inputs[82]);
    assign layer0_outputs[9141] = ~((inputs[187]) ^ (inputs[251]));
    assign layer0_outputs[9142] = (inputs[171]) | (inputs[97]);
    assign layer0_outputs[9143] = inputs[133];
    assign layer0_outputs[9144] = ~((inputs[132]) | (inputs[61]));
    assign layer0_outputs[9145] = 1'b0;
    assign layer0_outputs[9146] = ~(inputs[42]) | (inputs[135]);
    assign layer0_outputs[9147] = (inputs[65]) & (inputs[70]);
    assign layer0_outputs[9148] = inputs[247];
    assign layer0_outputs[9149] = (inputs[36]) ^ (inputs[254]);
    assign layer0_outputs[9150] = (inputs[195]) & ~(inputs[85]);
    assign layer0_outputs[9151] = 1'b0;
    assign layer0_outputs[9152] = inputs[83];
    assign layer0_outputs[9153] = ~(inputs[138]) | (inputs[60]);
    assign layer0_outputs[9154] = ~((inputs[199]) | (inputs[59]));
    assign layer0_outputs[9155] = (inputs[216]) & (inputs[209]);
    assign layer0_outputs[9156] = ~((inputs[113]) ^ (inputs[138]));
    assign layer0_outputs[9157] = ~((inputs[155]) | (inputs[35]));
    assign layer0_outputs[9158] = inputs[244];
    assign layer0_outputs[9159] = inputs[153];
    assign layer0_outputs[9160] = ~((inputs[98]) | (inputs[37]));
    assign layer0_outputs[9161] = (inputs[132]) & ~(inputs[252]);
    assign layer0_outputs[9162] = (inputs[152]) | (inputs[255]);
    assign layer0_outputs[9163] = ~(inputs[101]);
    assign layer0_outputs[9164] = inputs[47];
    assign layer0_outputs[9165] = inputs[128];
    assign layer0_outputs[9166] = (inputs[162]) & ~(inputs[243]);
    assign layer0_outputs[9167] = (inputs[239]) & ~(inputs[214]);
    assign layer0_outputs[9168] = (inputs[83]) | (inputs[201]);
    assign layer0_outputs[9169] = ~(inputs[228]);
    assign layer0_outputs[9170] = inputs[57];
    assign layer0_outputs[9171] = ~(inputs[78]);
    assign layer0_outputs[9172] = 1'b1;
    assign layer0_outputs[9173] = ~((inputs[145]) | (inputs[90]));
    assign layer0_outputs[9174] = ~(inputs[121]) | (inputs[229]);
    assign layer0_outputs[9175] = ~(inputs[107]);
    assign layer0_outputs[9176] = ~(inputs[104]);
    assign layer0_outputs[9177] = (inputs[222]) & ~(inputs[210]);
    assign layer0_outputs[9178] = (inputs[43]) | (inputs[75]);
    assign layer0_outputs[9179] = ~(inputs[229]);
    assign layer0_outputs[9180] = (inputs[82]) & ~(inputs[229]);
    assign layer0_outputs[9181] = inputs[149];
    assign layer0_outputs[9182] = ~(inputs[212]);
    assign layer0_outputs[9183] = ~((inputs[154]) ^ (inputs[236]));
    assign layer0_outputs[9184] = 1'b1;
    assign layer0_outputs[9185] = ~(inputs[73]) | (inputs[34]);
    assign layer0_outputs[9186] = ~((inputs[46]) | (inputs[101]));
    assign layer0_outputs[9187] = ~(inputs[44]);
    assign layer0_outputs[9188] = ~(inputs[209]) | (inputs[15]);
    assign layer0_outputs[9189] = (inputs[157]) | (inputs[172]);
    assign layer0_outputs[9190] = (inputs[226]) & (inputs[200]);
    assign layer0_outputs[9191] = ~((inputs[78]) & (inputs[63]));
    assign layer0_outputs[9192] = ~(inputs[85]);
    assign layer0_outputs[9193] = 1'b1;
    assign layer0_outputs[9194] = ~((inputs[142]) | (inputs[20]));
    assign layer0_outputs[9195] = ~(inputs[101]);
    assign layer0_outputs[9196] = ~(inputs[169]) | (inputs[82]);
    assign layer0_outputs[9197] = inputs[167];
    assign layer0_outputs[9198] = ~(inputs[115]) | (inputs[192]);
    assign layer0_outputs[9199] = ~(inputs[120]) | (inputs[55]);
    assign layer0_outputs[9200] = ~((inputs[241]) ^ (inputs[44]));
    assign layer0_outputs[9201] = ~((inputs[116]) | (inputs[87]));
    assign layer0_outputs[9202] = ~((inputs[238]) | (inputs[120]));
    assign layer0_outputs[9203] = 1'b0;
    assign layer0_outputs[9204] = ~((inputs[206]) ^ (inputs[20]));
    assign layer0_outputs[9205] = inputs[89];
    assign layer0_outputs[9206] = ~(inputs[145]) | (inputs[66]);
    assign layer0_outputs[9207] = ~((inputs[29]) | (inputs[53]));
    assign layer0_outputs[9208] = inputs[235];
    assign layer0_outputs[9209] = inputs[121];
    assign layer0_outputs[9210] = ~(inputs[101]) | (inputs[91]);
    assign layer0_outputs[9211] = ~(inputs[149]);
    assign layer0_outputs[9212] = ~(inputs[202]);
    assign layer0_outputs[9213] = ~((inputs[222]) ^ (inputs[211]));
    assign layer0_outputs[9214] = ~((inputs[186]) ^ (inputs[187]));
    assign layer0_outputs[9215] = ~((inputs[79]) | (inputs[25]));
    assign layer0_outputs[9216] = (inputs[99]) & ~(inputs[195]);
    assign layer0_outputs[9217] = (inputs[210]) & ~(inputs[64]);
    assign layer0_outputs[9218] = inputs[145];
    assign layer0_outputs[9219] = (inputs[101]) ^ (inputs[109]);
    assign layer0_outputs[9220] = (inputs[90]) | (inputs[181]);
    assign layer0_outputs[9221] = ~(inputs[90]);
    assign layer0_outputs[9222] = (inputs[37]) | (inputs[250]);
    assign layer0_outputs[9223] = ~((inputs[250]) | (inputs[223]));
    assign layer0_outputs[9224] = (inputs[225]) ^ (inputs[189]);
    assign layer0_outputs[9225] = (inputs[234]) & ~(inputs[175]);
    assign layer0_outputs[9226] = ~(inputs[31]);
    assign layer0_outputs[9227] = ~(inputs[193]);
    assign layer0_outputs[9228] = ~((inputs[34]) | (inputs[246]));
    assign layer0_outputs[9229] = inputs[156];
    assign layer0_outputs[9230] = ~((inputs[6]) | (inputs[131]));
    assign layer0_outputs[9231] = ~(inputs[156]);
    assign layer0_outputs[9232] = ~((inputs[144]) & (inputs[101]));
    assign layer0_outputs[9233] = inputs[82];
    assign layer0_outputs[9234] = 1'b0;
    assign layer0_outputs[9235] = (inputs[242]) | (inputs[246]);
    assign layer0_outputs[9236] = (inputs[66]) & ~(inputs[249]);
    assign layer0_outputs[9237] = ~((inputs[128]) ^ (inputs[130]));
    assign layer0_outputs[9238] = ~((inputs[243]) | (inputs[46]));
    assign layer0_outputs[9239] = 1'b0;
    assign layer0_outputs[9240] = inputs[121];
    assign layer0_outputs[9241] = (inputs[196]) ^ (inputs[148]);
    assign layer0_outputs[9242] = ~(inputs[37]);
    assign layer0_outputs[9243] = inputs[229];
    assign layer0_outputs[9244] = (inputs[167]) & ~(inputs[88]);
    assign layer0_outputs[9245] = ~((inputs[191]) & (inputs[31]));
    assign layer0_outputs[9246] = inputs[171];
    assign layer0_outputs[9247] = (inputs[205]) | (inputs[211]);
    assign layer0_outputs[9248] = inputs[18];
    assign layer0_outputs[9249] = ~(inputs[219]) | (inputs[29]);
    assign layer0_outputs[9250] = ~(inputs[126]);
    assign layer0_outputs[9251] = inputs[115];
    assign layer0_outputs[9252] = 1'b0;
    assign layer0_outputs[9253] = ~(inputs[203]);
    assign layer0_outputs[9254] = (inputs[222]) | (inputs[233]);
    assign layer0_outputs[9255] = inputs[163];
    assign layer0_outputs[9256] = ~(inputs[249]) | (inputs[0]);
    assign layer0_outputs[9257] = ~(inputs[196]);
    assign layer0_outputs[9258] = ~(inputs[50]);
    assign layer0_outputs[9259] = (inputs[19]) | (inputs[251]);
    assign layer0_outputs[9260] = inputs[45];
    assign layer0_outputs[9261] = (inputs[103]) & ~(inputs[2]);
    assign layer0_outputs[9262] = ~(inputs[28]);
    assign layer0_outputs[9263] = 1'b0;
    assign layer0_outputs[9264] = (inputs[216]) & ~(inputs[169]);
    assign layer0_outputs[9265] = ~(inputs[93]);
    assign layer0_outputs[9266] = ~(inputs[246]);
    assign layer0_outputs[9267] = ~(inputs[51]);
    assign layer0_outputs[9268] = (inputs[80]) & ~(inputs[99]);
    assign layer0_outputs[9269] = ~(inputs[50]);
    assign layer0_outputs[9270] = (inputs[176]) & ~(inputs[140]);
    assign layer0_outputs[9271] = inputs[87];
    assign layer0_outputs[9272] = inputs[67];
    assign layer0_outputs[9273] = (inputs[16]) ^ (inputs[204]);
    assign layer0_outputs[9274] = ~((inputs[142]) | (inputs[215]));
    assign layer0_outputs[9275] = 1'b1;
    assign layer0_outputs[9276] = (inputs[230]) & ~(inputs[28]);
    assign layer0_outputs[9277] = (inputs[100]) ^ (inputs[189]);
    assign layer0_outputs[9278] = ~((inputs[75]) & (inputs[9]));
    assign layer0_outputs[9279] = ~((inputs[16]) ^ (inputs[243]));
    assign layer0_outputs[9280] = ~((inputs[196]) | (inputs[155]));
    assign layer0_outputs[9281] = ~(inputs[151]);
    assign layer0_outputs[9282] = (inputs[172]) & ~(inputs[49]);
    assign layer0_outputs[9283] = ~(inputs[134]);
    assign layer0_outputs[9284] = (inputs[50]) | (inputs[181]);
    assign layer0_outputs[9285] = ~((inputs[223]) | (inputs[214]));
    assign layer0_outputs[9286] = ~((inputs[50]) | (inputs[196]));
    assign layer0_outputs[9287] = ~((inputs[146]) ^ (inputs[248]));
    assign layer0_outputs[9288] = ~((inputs[112]) ^ (inputs[85]));
    assign layer0_outputs[9289] = inputs[165];
    assign layer0_outputs[9290] = (inputs[5]) ^ (inputs[34]);
    assign layer0_outputs[9291] = ~(inputs[150]);
    assign layer0_outputs[9292] = inputs[94];
    assign layer0_outputs[9293] = inputs[133];
    assign layer0_outputs[9294] = inputs[145];
    assign layer0_outputs[9295] = ~((inputs[135]) | (inputs[151]));
    assign layer0_outputs[9296] = inputs[108];
    assign layer0_outputs[9297] = (inputs[107]) & ~(inputs[129]);
    assign layer0_outputs[9298] = (inputs[247]) ^ (inputs[114]);
    assign layer0_outputs[9299] = (inputs[165]) & ~(inputs[53]);
    assign layer0_outputs[9300] = 1'b1;
    assign layer0_outputs[9301] = (inputs[166]) | (inputs[185]);
    assign layer0_outputs[9302] = ~(inputs[221]);
    assign layer0_outputs[9303] = ~((inputs[174]) ^ (inputs[175]));
    assign layer0_outputs[9304] = inputs[108];
    assign layer0_outputs[9305] = ~(inputs[204]);
    assign layer0_outputs[9306] = (inputs[79]) ^ (inputs[2]);
    assign layer0_outputs[9307] = ~(inputs[60]);
    assign layer0_outputs[9308] = (inputs[34]) ^ (inputs[124]);
    assign layer0_outputs[9309] = ~(inputs[24]) | (inputs[235]);
    assign layer0_outputs[9310] = inputs[8];
    assign layer0_outputs[9311] = inputs[244];
    assign layer0_outputs[9312] = (inputs[217]) ^ (inputs[101]);
    assign layer0_outputs[9313] = inputs[226];
    assign layer0_outputs[9314] = ~(inputs[171]);
    assign layer0_outputs[9315] = inputs[113];
    assign layer0_outputs[9316] = ~((inputs[231]) ^ (inputs[236]));
    assign layer0_outputs[9317] = ~(inputs[76]) | (inputs[146]);
    assign layer0_outputs[9318] = ~((inputs[12]) | (inputs[22]));
    assign layer0_outputs[9319] = inputs[178];
    assign layer0_outputs[9320] = (inputs[75]) | (inputs[162]);
    assign layer0_outputs[9321] = (inputs[211]) & ~(inputs[164]);
    assign layer0_outputs[9322] = inputs[154];
    assign layer0_outputs[9323] = inputs[89];
    assign layer0_outputs[9324] = ~(inputs[29]);
    assign layer0_outputs[9325] = (inputs[176]) & ~(inputs[78]);
    assign layer0_outputs[9326] = ~(inputs[66]);
    assign layer0_outputs[9327] = (inputs[140]) & ~(inputs[197]);
    assign layer0_outputs[9328] = ~(inputs[199]);
    assign layer0_outputs[9329] = (inputs[163]) & ~(inputs[61]);
    assign layer0_outputs[9330] = 1'b1;
    assign layer0_outputs[9331] = ~((inputs[90]) | (inputs[173]));
    assign layer0_outputs[9332] = inputs[102];
    assign layer0_outputs[9333] = ~((inputs[155]) | (inputs[238]));
    assign layer0_outputs[9334] = (inputs[9]) & ~(inputs[240]);
    assign layer0_outputs[9335] = inputs[125];
    assign layer0_outputs[9336] = ~(inputs[173]);
    assign layer0_outputs[9337] = ~((inputs[249]) | (inputs[171]));
    assign layer0_outputs[9338] = inputs[108];
    assign layer0_outputs[9339] = ~(inputs[244]) | (inputs[219]);
    assign layer0_outputs[9340] = inputs[95];
    assign layer0_outputs[9341] = ~((inputs[19]) ^ (inputs[222]));
    assign layer0_outputs[9342] = ~(inputs[208]) | (inputs[67]);
    assign layer0_outputs[9343] = ~((inputs[101]) | (inputs[172]));
    assign layer0_outputs[9344] = inputs[46];
    assign layer0_outputs[9345] = ~(inputs[95]);
    assign layer0_outputs[9346] = (inputs[17]) & ~(inputs[118]);
    assign layer0_outputs[9347] = ~(inputs[126]);
    assign layer0_outputs[9348] = ~(inputs[153]);
    assign layer0_outputs[9349] = inputs[226];
    assign layer0_outputs[9350] = ~(inputs[252]) | (inputs[189]);
    assign layer0_outputs[9351] = (inputs[139]) | (inputs[144]);
    assign layer0_outputs[9352] = inputs[241];
    assign layer0_outputs[9353] = ~((inputs[108]) | (inputs[114]));
    assign layer0_outputs[9354] = 1'b0;
    assign layer0_outputs[9355] = ~(inputs[39]) | (inputs[63]);
    assign layer0_outputs[9356] = ~(inputs[66]);
    assign layer0_outputs[9357] = ~(inputs[92]);
    assign layer0_outputs[9358] = (inputs[231]) & ~(inputs[125]);
    assign layer0_outputs[9359] = ~((inputs[175]) | (inputs[196]));
    assign layer0_outputs[9360] = (inputs[19]) & ~(inputs[96]);
    assign layer0_outputs[9361] = 1'b1;
    assign layer0_outputs[9362] = (inputs[4]) | (inputs[103]);
    assign layer0_outputs[9363] = inputs[100];
    assign layer0_outputs[9364] = ~((inputs[40]) ^ (inputs[175]));
    assign layer0_outputs[9365] = ~((inputs[191]) ^ (inputs[236]));
    assign layer0_outputs[9366] = ~(inputs[106]);
    assign layer0_outputs[9367] = ~((inputs[15]) | (inputs[201]));
    assign layer0_outputs[9368] = ~(inputs[136]);
    assign layer0_outputs[9369] = ~(inputs[223]);
    assign layer0_outputs[9370] = (inputs[14]) & ~(inputs[76]);
    assign layer0_outputs[9371] = inputs[176];
    assign layer0_outputs[9372] = (inputs[42]) & (inputs[108]);
    assign layer0_outputs[9373] = (inputs[183]) & (inputs[36]);
    assign layer0_outputs[9374] = (inputs[73]) & ~(inputs[64]);
    assign layer0_outputs[9375] = ~((inputs[40]) ^ (inputs[60]));
    assign layer0_outputs[9376] = (inputs[2]) | (inputs[22]);
    assign layer0_outputs[9377] = (inputs[39]) & (inputs[237]);
    assign layer0_outputs[9378] = (inputs[30]) ^ (inputs[208]);
    assign layer0_outputs[9379] = ~((inputs[149]) ^ (inputs[176]));
    assign layer0_outputs[9380] = inputs[203];
    assign layer0_outputs[9381] = ~((inputs[177]) ^ (inputs[225]));
    assign layer0_outputs[9382] = (inputs[78]) ^ (inputs[133]);
    assign layer0_outputs[9383] = (inputs[91]) & ~(inputs[226]);
    assign layer0_outputs[9384] = (inputs[159]) & ~(inputs[190]);
    assign layer0_outputs[9385] = ~((inputs[35]) ^ (inputs[62]));
    assign layer0_outputs[9386] = ~(inputs[134]);
    assign layer0_outputs[9387] = (inputs[106]) & ~(inputs[89]);
    assign layer0_outputs[9388] = inputs[150];
    assign layer0_outputs[9389] = (inputs[196]) & ~(inputs[3]);
    assign layer0_outputs[9390] = ~(inputs[70]);
    assign layer0_outputs[9391] = ~(inputs[127]);
    assign layer0_outputs[9392] = inputs[148];
    assign layer0_outputs[9393] = ~((inputs[55]) ^ (inputs[49]));
    assign layer0_outputs[9394] = (inputs[248]) & ~(inputs[232]);
    assign layer0_outputs[9395] = ~(inputs[117]);
    assign layer0_outputs[9396] = ~(inputs[188]);
    assign layer0_outputs[9397] = ~((inputs[217]) | (inputs[187]));
    assign layer0_outputs[9398] = (inputs[85]) & ~(inputs[26]);
    assign layer0_outputs[9399] = ~((inputs[31]) | (inputs[3]));
    assign layer0_outputs[9400] = ~(inputs[23]) | (inputs[191]);
    assign layer0_outputs[9401] = ~(inputs[246]) | (inputs[240]);
    assign layer0_outputs[9402] = (inputs[61]) | (inputs[43]);
    assign layer0_outputs[9403] = (inputs[110]) ^ (inputs[163]);
    assign layer0_outputs[9404] = (inputs[120]) | (inputs[142]);
    assign layer0_outputs[9405] = 1'b1;
    assign layer0_outputs[9406] = (inputs[173]) & ~(inputs[65]);
    assign layer0_outputs[9407] = ~(inputs[81]) | (inputs[189]);
    assign layer0_outputs[9408] = inputs[125];
    assign layer0_outputs[9409] = ~((inputs[217]) | (inputs[132]));
    assign layer0_outputs[9410] = (inputs[117]) & ~(inputs[224]);
    assign layer0_outputs[9411] = ~(inputs[146]);
    assign layer0_outputs[9412] = ~(inputs[59]);
    assign layer0_outputs[9413] = ~(inputs[108]) | (inputs[133]);
    assign layer0_outputs[9414] = ~((inputs[178]) & (inputs[20]));
    assign layer0_outputs[9415] = inputs[162];
    assign layer0_outputs[9416] = ~((inputs[248]) & (inputs[138]));
    assign layer0_outputs[9417] = ~(inputs[125]);
    assign layer0_outputs[9418] = ~(inputs[211]);
    assign layer0_outputs[9419] = ~(inputs[93]);
    assign layer0_outputs[9420] = (inputs[75]) & ~(inputs[220]);
    assign layer0_outputs[9421] = inputs[75];
    assign layer0_outputs[9422] = ~((inputs[122]) ^ (inputs[92]));
    assign layer0_outputs[9423] = ~(inputs[23]) | (inputs[249]);
    assign layer0_outputs[9424] = ~((inputs[47]) & (inputs[229]));
    assign layer0_outputs[9425] = 1'b1;
    assign layer0_outputs[9426] = (inputs[61]) ^ (inputs[199]);
    assign layer0_outputs[9427] = ~(inputs[53]) | (inputs[207]);
    assign layer0_outputs[9428] = (inputs[139]) & (inputs[20]);
    assign layer0_outputs[9429] = ~((inputs[192]) | (inputs[226]));
    assign layer0_outputs[9430] = ~(inputs[233]) | (inputs[95]);
    assign layer0_outputs[9431] = ~(inputs[116]);
    assign layer0_outputs[9432] = (inputs[52]) ^ (inputs[226]);
    assign layer0_outputs[9433] = ~(inputs[146]);
    assign layer0_outputs[9434] = 1'b1;
    assign layer0_outputs[9435] = inputs[169];
    assign layer0_outputs[9436] = (inputs[141]) | (inputs[178]);
    assign layer0_outputs[9437] = (inputs[223]) ^ (inputs[130]);
    assign layer0_outputs[9438] = ~((inputs[251]) ^ (inputs[255]));
    assign layer0_outputs[9439] = ~(inputs[127]) | (inputs[10]);
    assign layer0_outputs[9440] = ~((inputs[130]) ^ (inputs[249]));
    assign layer0_outputs[9441] = ~((inputs[4]) | (inputs[209]));
    assign layer0_outputs[9442] = inputs[232];
    assign layer0_outputs[9443] = 1'b0;
    assign layer0_outputs[9444] = ~(inputs[247]);
    assign layer0_outputs[9445] = ~(inputs[6]) | (inputs[235]);
    assign layer0_outputs[9446] = 1'b0;
    assign layer0_outputs[9447] = ~(inputs[126]) | (inputs[245]);
    assign layer0_outputs[9448] = (inputs[165]) | (inputs[206]);
    assign layer0_outputs[9449] = ~(inputs[84]) | (inputs[24]);
    assign layer0_outputs[9450] = ~(inputs[98]);
    assign layer0_outputs[9451] = ~(inputs[88]);
    assign layer0_outputs[9452] = ~((inputs[187]) & (inputs[144]));
    assign layer0_outputs[9453] = ~(inputs[120]) | (inputs[113]);
    assign layer0_outputs[9454] = ~(inputs[73]);
    assign layer0_outputs[9455] = ~(inputs[176]);
    assign layer0_outputs[9456] = ~(inputs[136]);
    assign layer0_outputs[9457] = ~((inputs[235]) ^ (inputs[208]));
    assign layer0_outputs[9458] = ~(inputs[22]);
    assign layer0_outputs[9459] = (inputs[63]) | (inputs[243]);
    assign layer0_outputs[9460] = (inputs[62]) ^ (inputs[108]);
    assign layer0_outputs[9461] = 1'b0;
    assign layer0_outputs[9462] = ~(inputs[91]) | (inputs[97]);
    assign layer0_outputs[9463] = ~((inputs[109]) | (inputs[233]));
    assign layer0_outputs[9464] = (inputs[112]) & ~(inputs[73]);
    assign layer0_outputs[9465] = ~(inputs[198]);
    assign layer0_outputs[9466] = ~((inputs[0]) & (inputs[175]));
    assign layer0_outputs[9467] = ~((inputs[20]) | (inputs[242]));
    assign layer0_outputs[9468] = inputs[214];
    assign layer0_outputs[9469] = ~((inputs[77]) | (inputs[123]));
    assign layer0_outputs[9470] = ~(inputs[159]);
    assign layer0_outputs[9471] = (inputs[123]) ^ (inputs[45]);
    assign layer0_outputs[9472] = ~(inputs[199]) | (inputs[191]);
    assign layer0_outputs[9473] = inputs[80];
    assign layer0_outputs[9474] = 1'b1;
    assign layer0_outputs[9475] = ~(inputs[160]) | (inputs[253]);
    assign layer0_outputs[9476] = ~((inputs[119]) | (inputs[195]));
    assign layer0_outputs[9477] = (inputs[66]) | (inputs[244]);
    assign layer0_outputs[9478] = 1'b0;
    assign layer0_outputs[9479] = ~((inputs[72]) ^ (inputs[123]));
    assign layer0_outputs[9480] = (inputs[145]) & ~(inputs[168]);
    assign layer0_outputs[9481] = 1'b0;
    assign layer0_outputs[9482] = 1'b0;
    assign layer0_outputs[9483] = (inputs[163]) | (inputs[220]);
    assign layer0_outputs[9484] = inputs[2];
    assign layer0_outputs[9485] = ~((inputs[48]) ^ (inputs[252]));
    assign layer0_outputs[9486] = 1'b1;
    assign layer0_outputs[9487] = ~(inputs[231]);
    assign layer0_outputs[9488] = ~((inputs[242]) & (inputs[144]));
    assign layer0_outputs[9489] = ~((inputs[92]) | (inputs[237]));
    assign layer0_outputs[9490] = 1'b1;
    assign layer0_outputs[9491] = (inputs[194]) & ~(inputs[81]);
    assign layer0_outputs[9492] = ~((inputs[93]) ^ (inputs[91]));
    assign layer0_outputs[9493] = inputs[110];
    assign layer0_outputs[9494] = (inputs[141]) | (inputs[79]);
    assign layer0_outputs[9495] = (inputs[8]) ^ (inputs[191]);
    assign layer0_outputs[9496] = ~(inputs[182]);
    assign layer0_outputs[9497] = (inputs[173]) ^ (inputs[5]);
    assign layer0_outputs[9498] = ~(inputs[195]);
    assign layer0_outputs[9499] = (inputs[93]) | (inputs[38]);
    assign layer0_outputs[9500] = ~(inputs[108]);
    assign layer0_outputs[9501] = (inputs[243]) & ~(inputs[224]);
    assign layer0_outputs[9502] = inputs[216];
    assign layer0_outputs[9503] = (inputs[34]) & ~(inputs[187]);
    assign layer0_outputs[9504] = ~((inputs[186]) | (inputs[141]));
    assign layer0_outputs[9505] = ~(inputs[179]);
    assign layer0_outputs[9506] = ~((inputs[11]) | (inputs[196]));
    assign layer0_outputs[9507] = inputs[150];
    assign layer0_outputs[9508] = inputs[0];
    assign layer0_outputs[9509] = (inputs[117]) & ~(inputs[93]);
    assign layer0_outputs[9510] = ~((inputs[15]) & (inputs[190]));
    assign layer0_outputs[9511] = (inputs[213]) | (inputs[73]);
    assign layer0_outputs[9512] = ~(inputs[182]);
    assign layer0_outputs[9513] = inputs[70];
    assign layer0_outputs[9514] = ~((inputs[91]) ^ (inputs[142]));
    assign layer0_outputs[9515] = inputs[76];
    assign layer0_outputs[9516] = 1'b1;
    assign layer0_outputs[9517] = 1'b1;
    assign layer0_outputs[9518] = inputs[6];
    assign layer0_outputs[9519] = ~(inputs[244]);
    assign layer0_outputs[9520] = ~(inputs[68]) | (inputs[222]);
    assign layer0_outputs[9521] = ~(inputs[120]);
    assign layer0_outputs[9522] = ~(inputs[84]);
    assign layer0_outputs[9523] = inputs[124];
    assign layer0_outputs[9524] = (inputs[195]) & ~(inputs[45]);
    assign layer0_outputs[9525] = (inputs[146]) ^ (inputs[176]);
    assign layer0_outputs[9526] = (inputs[203]) | (inputs[146]);
    assign layer0_outputs[9527] = (inputs[53]) | (inputs[69]);
    assign layer0_outputs[9528] = (inputs[17]) | (inputs[240]);
    assign layer0_outputs[9529] = (inputs[145]) & ~(inputs[10]);
    assign layer0_outputs[9530] = ~(inputs[122]) | (inputs[129]);
    assign layer0_outputs[9531] = inputs[55];
    assign layer0_outputs[9532] = (inputs[156]) ^ (inputs[190]);
    assign layer0_outputs[9533] = inputs[161];
    assign layer0_outputs[9534] = ~((inputs[236]) ^ (inputs[172]));
    assign layer0_outputs[9535] = (inputs[243]) | (inputs[115]);
    assign layer0_outputs[9536] = ~(inputs[209]) | (inputs[198]);
    assign layer0_outputs[9537] = ~(inputs[228]) | (inputs[1]);
    assign layer0_outputs[9538] = ~((inputs[189]) ^ (inputs[249]));
    assign layer0_outputs[9539] = (inputs[47]) | (inputs[151]);
    assign layer0_outputs[9540] = ~(inputs[33]);
    assign layer0_outputs[9541] = 1'b0;
    assign layer0_outputs[9542] = ~(inputs[180]) | (inputs[173]);
    assign layer0_outputs[9543] = ~(inputs[220]) | (inputs[22]);
    assign layer0_outputs[9544] = ~(inputs[148]) | (inputs[105]);
    assign layer0_outputs[9545] = (inputs[213]) & ~(inputs[47]);
    assign layer0_outputs[9546] = ~(inputs[179]);
    assign layer0_outputs[9547] = (inputs[212]) & (inputs[29]);
    assign layer0_outputs[9548] = ~(inputs[146]);
    assign layer0_outputs[9549] = ~(inputs[222]);
    assign layer0_outputs[9550] = inputs[228];
    assign layer0_outputs[9551] = ~(inputs[203]);
    assign layer0_outputs[9552] = (inputs[154]) & ~(inputs[245]);
    assign layer0_outputs[9553] = 1'b0;
    assign layer0_outputs[9554] = ~((inputs[122]) | (inputs[229]));
    assign layer0_outputs[9555] = inputs[247];
    assign layer0_outputs[9556] = ~((inputs[20]) | (inputs[61]));
    assign layer0_outputs[9557] = ~((inputs[44]) | (inputs[188]));
    assign layer0_outputs[9558] = (inputs[96]) | (inputs[130]);
    assign layer0_outputs[9559] = (inputs[18]) & ~(inputs[209]);
    assign layer0_outputs[9560] = (inputs[232]) & (inputs[166]);
    assign layer0_outputs[9561] = 1'b0;
    assign layer0_outputs[9562] = ~(inputs[180]) | (inputs[46]);
    assign layer0_outputs[9563] = ~(inputs[170]);
    assign layer0_outputs[9564] = ~((inputs[167]) ^ (inputs[216]));
    assign layer0_outputs[9565] = (inputs[52]) ^ (inputs[255]);
    assign layer0_outputs[9566] = ~((inputs[95]) ^ (inputs[189]));
    assign layer0_outputs[9567] = inputs[193];
    assign layer0_outputs[9568] = ~(inputs[246]) | (inputs[113]);
    assign layer0_outputs[9569] = ~((inputs[112]) ^ (inputs[50]));
    assign layer0_outputs[9570] = ~((inputs[32]) ^ (inputs[170]));
    assign layer0_outputs[9571] = (inputs[99]) ^ (inputs[102]);
    assign layer0_outputs[9572] = ~((inputs[22]) ^ (inputs[85]));
    assign layer0_outputs[9573] = ~(inputs[209]);
    assign layer0_outputs[9574] = ~(inputs[255]);
    assign layer0_outputs[9575] = ~(inputs[156]);
    assign layer0_outputs[9576] = (inputs[134]) | (inputs[26]);
    assign layer0_outputs[9577] = 1'b0;
    assign layer0_outputs[9578] = (inputs[66]) | (inputs[65]);
    assign layer0_outputs[9579] = ~(inputs[142]) | (inputs[12]);
    assign layer0_outputs[9580] = inputs[188];
    assign layer0_outputs[9581] = inputs[24];
    assign layer0_outputs[9582] = ~((inputs[112]) ^ (inputs[116]));
    assign layer0_outputs[9583] = ~(inputs[147]);
    assign layer0_outputs[9584] = (inputs[201]) ^ (inputs[203]);
    assign layer0_outputs[9585] = (inputs[143]) | (inputs[47]);
    assign layer0_outputs[9586] = ~((inputs[209]) ^ (inputs[246]));
    assign layer0_outputs[9587] = (inputs[217]) & ~(inputs[74]);
    assign layer0_outputs[9588] = ~((inputs[156]) ^ (inputs[159]));
    assign layer0_outputs[9589] = (inputs[75]) ^ (inputs[1]);
    assign layer0_outputs[9590] = (inputs[79]) & (inputs[18]);
    assign layer0_outputs[9591] = (inputs[223]) ^ (inputs[79]);
    assign layer0_outputs[9592] = ~(inputs[207]);
    assign layer0_outputs[9593] = inputs[129];
    assign layer0_outputs[9594] = (inputs[82]) ^ (inputs[168]);
    assign layer0_outputs[9595] = ~((inputs[213]) | (inputs[144]));
    assign layer0_outputs[9596] = ~((inputs[12]) | (inputs[98]));
    assign layer0_outputs[9597] = ~(inputs[115]);
    assign layer0_outputs[9598] = ~(inputs[115]) | (inputs[13]);
    assign layer0_outputs[9599] = ~(inputs[133]);
    assign layer0_outputs[9600] = ~(inputs[238]) | (inputs[35]);
    assign layer0_outputs[9601] = ~(inputs[157]);
    assign layer0_outputs[9602] = (inputs[196]) & ~(inputs[31]);
    assign layer0_outputs[9603] = (inputs[118]) & ~(inputs[119]);
    assign layer0_outputs[9604] = inputs[229];
    assign layer0_outputs[9605] = ~((inputs[181]) & (inputs[24]));
    assign layer0_outputs[9606] = ~(inputs[126]);
    assign layer0_outputs[9607] = inputs[59];
    assign layer0_outputs[9608] = ~((inputs[179]) | (inputs[195]));
    assign layer0_outputs[9609] = ~(inputs[97]);
    assign layer0_outputs[9610] = ~(inputs[69]);
    assign layer0_outputs[9611] = 1'b0;
    assign layer0_outputs[9612] = ~((inputs[106]) | (inputs[171]));
    assign layer0_outputs[9613] = ~(inputs[7]);
    assign layer0_outputs[9614] = inputs[53];
    assign layer0_outputs[9615] = ~(inputs[190]);
    assign layer0_outputs[9616] = ~(inputs[44]) | (inputs[146]);
    assign layer0_outputs[9617] = ~(inputs[186]) | (inputs[165]);
    assign layer0_outputs[9618] = (inputs[200]) ^ (inputs[231]);
    assign layer0_outputs[9619] = ~(inputs[232]) | (inputs[225]);
    assign layer0_outputs[9620] = (inputs[197]) | (inputs[130]);
    assign layer0_outputs[9621] = inputs[24];
    assign layer0_outputs[9622] = inputs[120];
    assign layer0_outputs[9623] = ~((inputs[72]) | (inputs[83]));
    assign layer0_outputs[9624] = (inputs[24]) & ~(inputs[179]);
    assign layer0_outputs[9625] = ~(inputs[125]);
    assign layer0_outputs[9626] = inputs[11];
    assign layer0_outputs[9627] = (inputs[23]) & ~(inputs[192]);
    assign layer0_outputs[9628] = ~(inputs[38]) | (inputs[157]);
    assign layer0_outputs[9629] = ~(inputs[232]) | (inputs[223]);
    assign layer0_outputs[9630] = (inputs[178]) & ~(inputs[18]);
    assign layer0_outputs[9631] = inputs[175];
    assign layer0_outputs[9632] = inputs[24];
    assign layer0_outputs[9633] = ~((inputs[66]) | (inputs[154]));
    assign layer0_outputs[9634] = ~((inputs[175]) | (inputs[200]));
    assign layer0_outputs[9635] = (inputs[213]) & (inputs[120]);
    assign layer0_outputs[9636] = ~((inputs[171]) | (inputs[200]));
    assign layer0_outputs[9637] = ~(inputs[65]);
    assign layer0_outputs[9638] = ~((inputs[73]) & (inputs[185]));
    assign layer0_outputs[9639] = inputs[100];
    assign layer0_outputs[9640] = (inputs[89]) & ~(inputs[207]);
    assign layer0_outputs[9641] = (inputs[177]) | (inputs[211]);
    assign layer0_outputs[9642] = ~((inputs[26]) & (inputs[234]));
    assign layer0_outputs[9643] = (inputs[5]) | (inputs[158]);
    assign layer0_outputs[9644] = (inputs[100]) ^ (inputs[181]);
    assign layer0_outputs[9645] = (inputs[223]) & ~(inputs[156]);
    assign layer0_outputs[9646] = ~(inputs[151]) | (inputs[8]);
    assign layer0_outputs[9647] = inputs[114];
    assign layer0_outputs[9648] = ~((inputs[250]) ^ (inputs[81]));
    assign layer0_outputs[9649] = 1'b1;
    assign layer0_outputs[9650] = (inputs[26]) & ~(inputs[148]);
    assign layer0_outputs[9651] = ~((inputs[97]) & (inputs[222]));
    assign layer0_outputs[9652] = (inputs[255]) & ~(inputs[121]);
    assign layer0_outputs[9653] = inputs[150];
    assign layer0_outputs[9654] = ~((inputs[50]) ^ (inputs[69]));
    assign layer0_outputs[9655] = inputs[77];
    assign layer0_outputs[9656] = inputs[60];
    assign layer0_outputs[9657] = inputs[84];
    assign layer0_outputs[9658] = ~((inputs[215]) | (inputs[78]));
    assign layer0_outputs[9659] = ~(inputs[196]);
    assign layer0_outputs[9660] = inputs[53];
    assign layer0_outputs[9661] = ~(inputs[149]);
    assign layer0_outputs[9662] = ~((inputs[186]) | (inputs[51]));
    assign layer0_outputs[9663] = ~(inputs[198]);
    assign layer0_outputs[9664] = 1'b0;
    assign layer0_outputs[9665] = inputs[121];
    assign layer0_outputs[9666] = ~(inputs[229]) | (inputs[125]);
    assign layer0_outputs[9667] = ~((inputs[193]) | (inputs[62]));
    assign layer0_outputs[9668] = ~(inputs[173]) | (inputs[45]);
    assign layer0_outputs[9669] = ~(inputs[103]);
    assign layer0_outputs[9670] = ~((inputs[155]) | (inputs[177]));
    assign layer0_outputs[9671] = ~(inputs[173]);
    assign layer0_outputs[9672] = 1'b0;
    assign layer0_outputs[9673] = ~((inputs[75]) | (inputs[20]));
    assign layer0_outputs[9674] = ~((inputs[249]) | (inputs[11]));
    assign layer0_outputs[9675] = ~((inputs[18]) ^ (inputs[57]));
    assign layer0_outputs[9676] = ~(inputs[70]) | (inputs[173]);
    assign layer0_outputs[9677] = (inputs[229]) & (inputs[21]);
    assign layer0_outputs[9678] = ~(inputs[151]);
    assign layer0_outputs[9679] = ~((inputs[112]) ^ (inputs[87]));
    assign layer0_outputs[9680] = (inputs[25]) | (inputs[33]);
    assign layer0_outputs[9681] = 1'b0;
    assign layer0_outputs[9682] = inputs[100];
    assign layer0_outputs[9683] = ~(inputs[204]);
    assign layer0_outputs[9684] = (inputs[40]) ^ (inputs[191]);
    assign layer0_outputs[9685] = ~(inputs[59]) | (inputs[191]);
    assign layer0_outputs[9686] = inputs[218];
    assign layer0_outputs[9687] = 1'b0;
    assign layer0_outputs[9688] = ~(inputs[122]);
    assign layer0_outputs[9689] = inputs[123];
    assign layer0_outputs[9690] = ~((inputs[28]) & (inputs[138]));
    assign layer0_outputs[9691] = (inputs[99]) & ~(inputs[215]);
    assign layer0_outputs[9692] = ~(inputs[84]);
    assign layer0_outputs[9693] = ~(inputs[235]);
    assign layer0_outputs[9694] = 1'b1;
    assign layer0_outputs[9695] = (inputs[238]) & ~(inputs[17]);
    assign layer0_outputs[9696] = (inputs[28]) | (inputs[250]);
    assign layer0_outputs[9697] = inputs[224];
    assign layer0_outputs[9698] = ~(inputs[26]) | (inputs[198]);
    assign layer0_outputs[9699] = (inputs[177]) ^ (inputs[174]);
    assign layer0_outputs[9700] = ~((inputs[207]) | (inputs[94]));
    assign layer0_outputs[9701] = ~(inputs[140]) | (inputs[98]);
    assign layer0_outputs[9702] = ~((inputs[169]) & (inputs[197]));
    assign layer0_outputs[9703] = (inputs[58]) ^ (inputs[238]);
    assign layer0_outputs[9704] = ~(inputs[102]);
    assign layer0_outputs[9705] = ~(inputs[135]);
    assign layer0_outputs[9706] = ~((inputs[131]) | (inputs[226]));
    assign layer0_outputs[9707] = (inputs[118]) & ~(inputs[17]);
    assign layer0_outputs[9708] = (inputs[39]) & (inputs[57]);
    assign layer0_outputs[9709] = (inputs[91]) & ~(inputs[34]);
    assign layer0_outputs[9710] = (inputs[188]) | (inputs[13]);
    assign layer0_outputs[9711] = ~(inputs[248]);
    assign layer0_outputs[9712] = ~(inputs[41]);
    assign layer0_outputs[9713] = (inputs[100]) | (inputs[100]);
    assign layer0_outputs[9714] = (inputs[21]) ^ (inputs[255]);
    assign layer0_outputs[9715] = 1'b0;
    assign layer0_outputs[9716] = (inputs[126]) & ~(inputs[97]);
    assign layer0_outputs[9717] = (inputs[63]) | (inputs[36]);
    assign layer0_outputs[9718] = ~(inputs[229]);
    assign layer0_outputs[9719] = inputs[87];
    assign layer0_outputs[9720] = (inputs[207]) & ~(inputs[27]);
    assign layer0_outputs[9721] = ~(inputs[103]);
    assign layer0_outputs[9722] = (inputs[33]) & ~(inputs[174]);
    assign layer0_outputs[9723] = ~((inputs[187]) ^ (inputs[177]));
    assign layer0_outputs[9724] = (inputs[87]) ^ (inputs[129]);
    assign layer0_outputs[9725] = inputs[107];
    assign layer0_outputs[9726] = ~((inputs[81]) | (inputs[157]));
    assign layer0_outputs[9727] = ~(inputs[101]);
    assign layer0_outputs[9728] = 1'b1;
    assign layer0_outputs[9729] = inputs[33];
    assign layer0_outputs[9730] = (inputs[4]) | (inputs[123]);
    assign layer0_outputs[9731] = ~(inputs[49]);
    assign layer0_outputs[9732] = inputs[60];
    assign layer0_outputs[9733] = ~(inputs[36]) | (inputs[242]);
    assign layer0_outputs[9734] = ~(inputs[192]);
    assign layer0_outputs[9735] = ~(inputs[26]) | (inputs[54]);
    assign layer0_outputs[9736] = ~(inputs[183]);
    assign layer0_outputs[9737] = ~((inputs[210]) & (inputs[215]));
    assign layer0_outputs[9738] = (inputs[15]) & ~(inputs[217]);
    assign layer0_outputs[9739] = inputs[90];
    assign layer0_outputs[9740] = ~((inputs[132]) ^ (inputs[163]));
    assign layer0_outputs[9741] = ~(inputs[102]) | (inputs[126]);
    assign layer0_outputs[9742] = (inputs[17]) & ~(inputs[145]);
    assign layer0_outputs[9743] = ~(inputs[20]);
    assign layer0_outputs[9744] = (inputs[96]) ^ (inputs[114]);
    assign layer0_outputs[9745] = ~(inputs[101]);
    assign layer0_outputs[9746] = inputs[175];
    assign layer0_outputs[9747] = inputs[213];
    assign layer0_outputs[9748] = inputs[29];
    assign layer0_outputs[9749] = ~(inputs[98]) | (inputs[75]);
    assign layer0_outputs[9750] = (inputs[158]) | (inputs[219]);
    assign layer0_outputs[9751] = ~(inputs[99]) | (inputs[7]);
    assign layer0_outputs[9752] = ~(inputs[135]) | (inputs[217]);
    assign layer0_outputs[9753] = ~(inputs[32]);
    assign layer0_outputs[9754] = (inputs[172]) ^ (inputs[208]);
    assign layer0_outputs[9755] = (inputs[65]) ^ (inputs[53]);
    assign layer0_outputs[9756] = ~((inputs[250]) | (inputs[196]));
    assign layer0_outputs[9757] = inputs[159];
    assign layer0_outputs[9758] = ~((inputs[200]) ^ (inputs[176]));
    assign layer0_outputs[9759] = inputs[136];
    assign layer0_outputs[9760] = ~((inputs[235]) | (inputs[110]));
    assign layer0_outputs[9761] = ~(inputs[114]) | (inputs[114]);
    assign layer0_outputs[9762] = ~((inputs[200]) ^ (inputs[110]));
    assign layer0_outputs[9763] = (inputs[21]) & ~(inputs[179]);
    assign layer0_outputs[9764] = ~(inputs[211]) | (inputs[236]);
    assign layer0_outputs[9765] = ~(inputs[60]);
    assign layer0_outputs[9766] = ~(inputs[131]) | (inputs[209]);
    assign layer0_outputs[9767] = ~((inputs[70]) & (inputs[154]));
    assign layer0_outputs[9768] = ~(inputs[241]);
    assign layer0_outputs[9769] = (inputs[233]) ^ (inputs[238]);
    assign layer0_outputs[9770] = ~(inputs[85]);
    assign layer0_outputs[9771] = 1'b0;
    assign layer0_outputs[9772] = ~(inputs[28]);
    assign layer0_outputs[9773] = ~(inputs[57]);
    assign layer0_outputs[9774] = (inputs[135]) | (inputs[235]);
    assign layer0_outputs[9775] = (inputs[107]) & ~(inputs[104]);
    assign layer0_outputs[9776] = (inputs[217]) & ~(inputs[60]);
    assign layer0_outputs[9777] = (inputs[21]) | (inputs[26]);
    assign layer0_outputs[9778] = (inputs[79]) & ~(inputs[250]);
    assign layer0_outputs[9779] = ~(inputs[102]);
    assign layer0_outputs[9780] = ~(inputs[104]) | (inputs[84]);
    assign layer0_outputs[9781] = ~((inputs[40]) | (inputs[187]));
    assign layer0_outputs[9782] = ~((inputs[65]) & (inputs[191]));
    assign layer0_outputs[9783] = ~((inputs[1]) ^ (inputs[96]));
    assign layer0_outputs[9784] = ~((inputs[170]) ^ (inputs[65]));
    assign layer0_outputs[9785] = (inputs[41]) & ~(inputs[83]);
    assign layer0_outputs[9786] = inputs[22];
    assign layer0_outputs[9787] = (inputs[65]) | (inputs[91]);
    assign layer0_outputs[9788] = (inputs[221]) ^ (inputs[119]);
    assign layer0_outputs[9789] = (inputs[86]) & ~(inputs[34]);
    assign layer0_outputs[9790] = (inputs[153]) & (inputs[13]);
    assign layer0_outputs[9791] = ~(inputs[46]);
    assign layer0_outputs[9792] = (inputs[50]) ^ (inputs[12]);
    assign layer0_outputs[9793] = inputs[99];
    assign layer0_outputs[9794] = (inputs[227]) | (inputs[107]);
    assign layer0_outputs[9795] = ~(inputs[207]);
    assign layer0_outputs[9796] = 1'b1;
    assign layer0_outputs[9797] = ~(inputs[175]);
    assign layer0_outputs[9798] = ~(inputs[50]) | (inputs[12]);
    assign layer0_outputs[9799] = (inputs[162]) ^ (inputs[207]);
    assign layer0_outputs[9800] = ~(inputs[75]);
    assign layer0_outputs[9801] = (inputs[132]) & ~(inputs[160]);
    assign layer0_outputs[9802] = inputs[51];
    assign layer0_outputs[9803] = ~(inputs[22]);
    assign layer0_outputs[9804] = ~(inputs[42]);
    assign layer0_outputs[9805] = ~(inputs[42]) | (inputs[224]);
    assign layer0_outputs[9806] = (inputs[186]) ^ (inputs[80]);
    assign layer0_outputs[9807] = (inputs[70]) ^ (inputs[75]);
    assign layer0_outputs[9808] = ~(inputs[133]) | (inputs[41]);
    assign layer0_outputs[9809] = (inputs[146]) | (inputs[247]);
    assign layer0_outputs[9810] = ~(inputs[59]) | (inputs[173]);
    assign layer0_outputs[9811] = inputs[44];
    assign layer0_outputs[9812] = ~((inputs[71]) | (inputs[5]));
    assign layer0_outputs[9813] = inputs[27];
    assign layer0_outputs[9814] = inputs[110];
    assign layer0_outputs[9815] = (inputs[2]) & (inputs[230]);
    assign layer0_outputs[9816] = (inputs[37]) | (inputs[124]);
    assign layer0_outputs[9817] = inputs[161];
    assign layer0_outputs[9818] = ~(inputs[60]) | (inputs[207]);
    assign layer0_outputs[9819] = ~((inputs[2]) | (inputs[62]));
    assign layer0_outputs[9820] = (inputs[213]) | (inputs[118]);
    assign layer0_outputs[9821] = inputs[121];
    assign layer0_outputs[9822] = 1'b1;
    assign layer0_outputs[9823] = (inputs[142]) ^ (inputs[80]);
    assign layer0_outputs[9824] = ~((inputs[15]) | (inputs[74]));
    assign layer0_outputs[9825] = (inputs[62]) | (inputs[32]);
    assign layer0_outputs[9826] = ~(inputs[166]);
    assign layer0_outputs[9827] = inputs[131];
    assign layer0_outputs[9828] = (inputs[104]) | (inputs[29]);
    assign layer0_outputs[9829] = inputs[137];
    assign layer0_outputs[9830] = (inputs[209]) | (inputs[248]);
    assign layer0_outputs[9831] = ~(inputs[105]);
    assign layer0_outputs[9832] = ~(inputs[34]);
    assign layer0_outputs[9833] = ~(inputs[140]) | (inputs[135]);
    assign layer0_outputs[9834] = ~((inputs[165]) & (inputs[71]));
    assign layer0_outputs[9835] = ~(inputs[13]);
    assign layer0_outputs[9836] = (inputs[76]) ^ (inputs[211]);
    assign layer0_outputs[9837] = (inputs[93]) ^ (inputs[19]);
    assign layer0_outputs[9838] = ~(inputs[82]);
    assign layer0_outputs[9839] = ~(inputs[56]);
    assign layer0_outputs[9840] = (inputs[249]) & (inputs[189]);
    assign layer0_outputs[9841] = (inputs[167]) & ~(inputs[117]);
    assign layer0_outputs[9842] = ~((inputs[238]) & (inputs[17]));
    assign layer0_outputs[9843] = ~(inputs[108]);
    assign layer0_outputs[9844] = (inputs[245]) & (inputs[9]);
    assign layer0_outputs[9845] = (inputs[106]) ^ (inputs[175]);
    assign layer0_outputs[9846] = inputs[54];
    assign layer0_outputs[9847] = (inputs[111]) & ~(inputs[78]);
    assign layer0_outputs[9848] = (inputs[13]) & (inputs[27]);
    assign layer0_outputs[9849] = (inputs[25]) & ~(inputs[15]);
    assign layer0_outputs[9850] = ~(inputs[192]);
    assign layer0_outputs[9851] = 1'b1;
    assign layer0_outputs[9852] = ~(inputs[115]) | (inputs[29]);
    assign layer0_outputs[9853] = inputs[96];
    assign layer0_outputs[9854] = (inputs[188]) & ~(inputs[106]);
    assign layer0_outputs[9855] = ~(inputs[196]);
    assign layer0_outputs[9856] = ~(inputs[10]);
    assign layer0_outputs[9857] = inputs[51];
    assign layer0_outputs[9858] = (inputs[53]) & ~(inputs[190]);
    assign layer0_outputs[9859] = (inputs[239]) & (inputs[0]);
    assign layer0_outputs[9860] = ~((inputs[75]) | (inputs[106]));
    assign layer0_outputs[9861] = ~(inputs[62]);
    assign layer0_outputs[9862] = ~(inputs[42]) | (inputs[164]);
    assign layer0_outputs[9863] = ~(inputs[59]);
    assign layer0_outputs[9864] = (inputs[212]) ^ (inputs[244]);
    assign layer0_outputs[9865] = (inputs[150]) | (inputs[30]);
    assign layer0_outputs[9866] = ~(inputs[49]);
    assign layer0_outputs[9867] = (inputs[85]) & ~(inputs[143]);
    assign layer0_outputs[9868] = ~(inputs[120]);
    assign layer0_outputs[9869] = ~((inputs[177]) | (inputs[25]));
    assign layer0_outputs[9870] = inputs[130];
    assign layer0_outputs[9871] = ~(inputs[218]) | (inputs[253]);
    assign layer0_outputs[9872] = inputs[232];
    assign layer0_outputs[9873] = ~((inputs[16]) & (inputs[138]));
    assign layer0_outputs[9874] = inputs[253];
    assign layer0_outputs[9875] = inputs[34];
    assign layer0_outputs[9876] = ~(inputs[7]) | (inputs[220]);
    assign layer0_outputs[9877] = ~(inputs[232]) | (inputs[54]);
    assign layer0_outputs[9878] = (inputs[170]) ^ (inputs[83]);
    assign layer0_outputs[9879] = inputs[183];
    assign layer0_outputs[9880] = ~(inputs[23]);
    assign layer0_outputs[9881] = ~(inputs[243]);
    assign layer0_outputs[9882] = (inputs[127]) & ~(inputs[220]);
    assign layer0_outputs[9883] = (inputs[149]) & ~(inputs[123]);
    assign layer0_outputs[9884] = (inputs[87]) & ~(inputs[81]);
    assign layer0_outputs[9885] = ~(inputs[211]) | (inputs[73]);
    assign layer0_outputs[9886] = ~((inputs[8]) ^ (inputs[55]));
    assign layer0_outputs[9887] = 1'b0;
    assign layer0_outputs[9888] = ~(inputs[166]);
    assign layer0_outputs[9889] = (inputs[191]) & (inputs[6]);
    assign layer0_outputs[9890] = (inputs[177]) & ~(inputs[135]);
    assign layer0_outputs[9891] = inputs[137];
    assign layer0_outputs[9892] = 1'b0;
    assign layer0_outputs[9893] = ~((inputs[106]) & (inputs[46]));
    assign layer0_outputs[9894] = 1'b0;
    assign layer0_outputs[9895] = inputs[215];
    assign layer0_outputs[9896] = ~((inputs[255]) | (inputs[122]));
    assign layer0_outputs[9897] = inputs[228];
    assign layer0_outputs[9898] = (inputs[240]) | (inputs[156]);
    assign layer0_outputs[9899] = (inputs[212]) & (inputs[109]);
    assign layer0_outputs[9900] = inputs[98];
    assign layer0_outputs[9901] = (inputs[131]) & ~(inputs[33]);
    assign layer0_outputs[9902] = ~(inputs[58]);
    assign layer0_outputs[9903] = ~((inputs[83]) ^ (inputs[132]));
    assign layer0_outputs[9904] = ~(inputs[136]);
    assign layer0_outputs[9905] = 1'b1;
    assign layer0_outputs[9906] = ~(inputs[146]);
    assign layer0_outputs[9907] = ~(inputs[136]) | (inputs[244]);
    assign layer0_outputs[9908] = (inputs[172]) | (inputs[55]);
    assign layer0_outputs[9909] = inputs[244];
    assign layer0_outputs[9910] = (inputs[50]) | (inputs[60]);
    assign layer0_outputs[9911] = (inputs[10]) | (inputs[0]);
    assign layer0_outputs[9912] = ~((inputs[40]) | (inputs[25]));
    assign layer0_outputs[9913] = ~((inputs[127]) & (inputs[141]));
    assign layer0_outputs[9914] = (inputs[190]) | (inputs[123]);
    assign layer0_outputs[9915] = ~((inputs[228]) | (inputs[187]));
    assign layer0_outputs[9916] = inputs[33];
    assign layer0_outputs[9917] = ~(inputs[54]);
    assign layer0_outputs[9918] = ~((inputs[128]) & (inputs[143]));
    assign layer0_outputs[9919] = inputs[181];
    assign layer0_outputs[9920] = inputs[231];
    assign layer0_outputs[9921] = ~(inputs[22]) | (inputs[240]);
    assign layer0_outputs[9922] = ~(inputs[100]);
    assign layer0_outputs[9923] = ~(inputs[81]);
    assign layer0_outputs[9924] = (inputs[153]) | (inputs[67]);
    assign layer0_outputs[9925] = ~(inputs[16]) | (inputs[173]);
    assign layer0_outputs[9926] = ~(inputs[56]);
    assign layer0_outputs[9927] = inputs[140];
    assign layer0_outputs[9928] = (inputs[38]) | (inputs[131]);
    assign layer0_outputs[9929] = ~(inputs[132]);
    assign layer0_outputs[9930] = (inputs[188]) | (inputs[202]);
    assign layer0_outputs[9931] = (inputs[205]) | (inputs[118]);
    assign layer0_outputs[9932] = inputs[60];
    assign layer0_outputs[9933] = ~(inputs[30]) | (inputs[127]);
    assign layer0_outputs[9934] = (inputs[71]) ^ (inputs[229]);
    assign layer0_outputs[9935] = inputs[194];
    assign layer0_outputs[9936] = ~((inputs[199]) | (inputs[23]));
    assign layer0_outputs[9937] = (inputs[85]) & ~(inputs[140]);
    assign layer0_outputs[9938] = 1'b1;
    assign layer0_outputs[9939] = (inputs[144]) | (inputs[132]);
    assign layer0_outputs[9940] = ~((inputs[52]) ^ (inputs[39]));
    assign layer0_outputs[9941] = 1'b1;
    assign layer0_outputs[9942] = (inputs[81]) | (inputs[215]);
    assign layer0_outputs[9943] = (inputs[62]) | (inputs[250]);
    assign layer0_outputs[9944] = (inputs[191]) | (inputs[179]);
    assign layer0_outputs[9945] = ~((inputs[57]) ^ (inputs[12]));
    assign layer0_outputs[9946] = inputs[254];
    assign layer0_outputs[9947] = 1'b1;
    assign layer0_outputs[9948] = (inputs[167]) & ~(inputs[26]);
    assign layer0_outputs[9949] = inputs[165];
    assign layer0_outputs[9950] = (inputs[149]) & ~(inputs[0]);
    assign layer0_outputs[9951] = ~(inputs[100]);
    assign layer0_outputs[9952] = ~(inputs[163]) | (inputs[97]);
    assign layer0_outputs[9953] = inputs[25];
    assign layer0_outputs[9954] = ~(inputs[238]);
    assign layer0_outputs[9955] = (inputs[119]) & (inputs[149]);
    assign layer0_outputs[9956] = (inputs[245]) | (inputs[79]);
    assign layer0_outputs[9957] = ~(inputs[25]);
    assign layer0_outputs[9958] = (inputs[103]) & ~(inputs[127]);
    assign layer0_outputs[9959] = ~((inputs[105]) | (inputs[66]));
    assign layer0_outputs[9960] = ~((inputs[223]) | (inputs[126]));
    assign layer0_outputs[9961] = (inputs[190]) & ~(inputs[242]);
    assign layer0_outputs[9962] = ~((inputs[119]) ^ (inputs[113]));
    assign layer0_outputs[9963] = (inputs[52]) | (inputs[89]);
    assign layer0_outputs[9964] = (inputs[76]) & ~(inputs[178]);
    assign layer0_outputs[9965] = (inputs[106]) | (inputs[239]);
    assign layer0_outputs[9966] = (inputs[46]) | (inputs[237]);
    assign layer0_outputs[9967] = (inputs[34]) & ~(inputs[191]);
    assign layer0_outputs[9968] = ~(inputs[48]) | (inputs[22]);
    assign layer0_outputs[9969] = ~((inputs[192]) ^ (inputs[243]));
    assign layer0_outputs[9970] = (inputs[152]) & (inputs[189]);
    assign layer0_outputs[9971] = ~((inputs[161]) ^ (inputs[114]));
    assign layer0_outputs[9972] = (inputs[138]) | (inputs[251]);
    assign layer0_outputs[9973] = inputs[94];
    assign layer0_outputs[9974] = inputs[12];
    assign layer0_outputs[9975] = inputs[59];
    assign layer0_outputs[9976] = ~((inputs[9]) ^ (inputs[5]));
    assign layer0_outputs[9977] = (inputs[197]) | (inputs[53]);
    assign layer0_outputs[9978] = (inputs[67]) ^ (inputs[61]);
    assign layer0_outputs[9979] = (inputs[17]) & ~(inputs[63]);
    assign layer0_outputs[9980] = inputs[213];
    assign layer0_outputs[9981] = ~(inputs[111]) | (inputs[244]);
    assign layer0_outputs[9982] = (inputs[216]) ^ (inputs[161]);
    assign layer0_outputs[9983] = ~(inputs[84]);
    assign layer0_outputs[9984] = ~((inputs[128]) | (inputs[61]));
    assign layer0_outputs[9985] = ~(inputs[214]) | (inputs[125]);
    assign layer0_outputs[9986] = (inputs[229]) & ~(inputs[95]);
    assign layer0_outputs[9987] = inputs[76];
    assign layer0_outputs[9988] = ~(inputs[11]) | (inputs[67]);
    assign layer0_outputs[9989] = 1'b1;
    assign layer0_outputs[9990] = inputs[205];
    assign layer0_outputs[9991] = inputs[90];
    assign layer0_outputs[9992] = ~(inputs[191]) | (inputs[235]);
    assign layer0_outputs[9993] = ~(inputs[160]);
    assign layer0_outputs[9994] = ~(inputs[38]) | (inputs[112]);
    assign layer0_outputs[9995] = (inputs[164]) | (inputs[140]);
    assign layer0_outputs[9996] = ~(inputs[126]) | (inputs[244]);
    assign layer0_outputs[9997] = ~(inputs[91]) | (inputs[128]);
    assign layer0_outputs[9998] = (inputs[1]) | (inputs[165]);
    assign layer0_outputs[9999] = ~(inputs[11]) | (inputs[200]);
    assign layer0_outputs[10000] = (inputs[251]) & (inputs[184]);
    assign layer0_outputs[10001] = ~(inputs[7]) | (inputs[53]);
    assign layer0_outputs[10002] = (inputs[222]) | (inputs[246]);
    assign layer0_outputs[10003] = (inputs[141]) | (inputs[122]);
    assign layer0_outputs[10004] = ~(inputs[102]);
    assign layer0_outputs[10005] = 1'b0;
    assign layer0_outputs[10006] = 1'b1;
    assign layer0_outputs[10007] = (inputs[67]) & (inputs[132]);
    assign layer0_outputs[10008] = ~((inputs[25]) | (inputs[189]));
    assign layer0_outputs[10009] = ~((inputs[30]) & (inputs[45]));
    assign layer0_outputs[10010] = inputs[123];
    assign layer0_outputs[10011] = (inputs[188]) & ~(inputs[153]);
    assign layer0_outputs[10012] = (inputs[91]) & ~(inputs[235]);
    assign layer0_outputs[10013] = inputs[127];
    assign layer0_outputs[10014] = (inputs[17]) | (inputs[154]);
    assign layer0_outputs[10015] = ~(inputs[101]) | (inputs[126]);
    assign layer0_outputs[10016] = ~(inputs[119]);
    assign layer0_outputs[10017] = (inputs[43]) | (inputs[46]);
    assign layer0_outputs[10018] = ~(inputs[195]) | (inputs[44]);
    assign layer0_outputs[10019] = (inputs[95]) | (inputs[25]);
    assign layer0_outputs[10020] = ~((inputs[251]) | (inputs[156]));
    assign layer0_outputs[10021] = (inputs[29]) | (inputs[92]);
    assign layer0_outputs[10022] = 1'b1;
    assign layer0_outputs[10023] = (inputs[246]) & ~(inputs[236]);
    assign layer0_outputs[10024] = ~((inputs[174]) ^ (inputs[62]));
    assign layer0_outputs[10025] = (inputs[228]) ^ (inputs[176]);
    assign layer0_outputs[10026] = inputs[149];
    assign layer0_outputs[10027] = (inputs[248]) & ~(inputs[7]);
    assign layer0_outputs[10028] = ~((inputs[31]) ^ (inputs[177]));
    assign layer0_outputs[10029] = (inputs[76]) & (inputs[236]);
    assign layer0_outputs[10030] = ~((inputs[152]) | (inputs[221]));
    assign layer0_outputs[10031] = (inputs[177]) & ~(inputs[96]);
    assign layer0_outputs[10032] = inputs[85];
    assign layer0_outputs[10033] = (inputs[107]) & ~(inputs[194]);
    assign layer0_outputs[10034] = ~(inputs[24]);
    assign layer0_outputs[10035] = ~(inputs[76]);
    assign layer0_outputs[10036] = ~(inputs[172]) | (inputs[61]);
    assign layer0_outputs[10037] = inputs[130];
    assign layer0_outputs[10038] = ~(inputs[252]);
    assign layer0_outputs[10039] = ~((inputs[237]) ^ (inputs[93]));
    assign layer0_outputs[10040] = ~(inputs[246]);
    assign layer0_outputs[10041] = ~((inputs[235]) & (inputs[246]));
    assign layer0_outputs[10042] = ~(inputs[209]);
    assign layer0_outputs[10043] = inputs[213];
    assign layer0_outputs[10044] = ~((inputs[155]) ^ (inputs[197]));
    assign layer0_outputs[10045] = ~((inputs[191]) ^ (inputs[100]));
    assign layer0_outputs[10046] = ~((inputs[206]) | (inputs[20]));
    assign layer0_outputs[10047] = ~((inputs[168]) | (inputs[60]));
    assign layer0_outputs[10048] = (inputs[146]) & ~(inputs[120]);
    assign layer0_outputs[10049] = inputs[211];
    assign layer0_outputs[10050] = (inputs[222]) ^ (inputs[78]);
    assign layer0_outputs[10051] = (inputs[50]) ^ (inputs[155]);
    assign layer0_outputs[10052] = (inputs[195]) & ~(inputs[110]);
    assign layer0_outputs[10053] = (inputs[46]) | (inputs[44]);
    assign layer0_outputs[10054] = ~(inputs[254]) | (inputs[71]);
    assign layer0_outputs[10055] = inputs[197];
    assign layer0_outputs[10056] = (inputs[213]) & ~(inputs[14]);
    assign layer0_outputs[10057] = ~(inputs[112]);
    assign layer0_outputs[10058] = ~((inputs[192]) | (inputs[123]));
    assign layer0_outputs[10059] = (inputs[131]) & (inputs[146]);
    assign layer0_outputs[10060] = ~((inputs[217]) | (inputs[130]));
    assign layer0_outputs[10061] = (inputs[190]) | (inputs[149]);
    assign layer0_outputs[10062] = inputs[86];
    assign layer0_outputs[10063] = ~(inputs[143]);
    assign layer0_outputs[10064] = ~(inputs[155]);
    assign layer0_outputs[10065] = (inputs[113]) | (inputs[167]);
    assign layer0_outputs[10066] = ~(inputs[190]) | (inputs[52]);
    assign layer0_outputs[10067] = (inputs[62]) | (inputs[160]);
    assign layer0_outputs[10068] = ~(inputs[56]);
    assign layer0_outputs[10069] = ~(inputs[218]) | (inputs[93]);
    assign layer0_outputs[10070] = ~((inputs[154]) ^ (inputs[4]));
    assign layer0_outputs[10071] = inputs[180];
    assign layer0_outputs[10072] = ~((inputs[147]) ^ (inputs[223]));
    assign layer0_outputs[10073] = inputs[16];
    assign layer0_outputs[10074] = ~((inputs[206]) | (inputs[152]));
    assign layer0_outputs[10075] = ~(inputs[81]) | (inputs[30]);
    assign layer0_outputs[10076] = 1'b0;
    assign layer0_outputs[10077] = ~(inputs[95]) | (inputs[172]);
    assign layer0_outputs[10078] = inputs[191];
    assign layer0_outputs[10079] = inputs[124];
    assign layer0_outputs[10080] = ~((inputs[211]) | (inputs[145]));
    assign layer0_outputs[10081] = (inputs[103]) ^ (inputs[81]);
    assign layer0_outputs[10082] = inputs[97];
    assign layer0_outputs[10083] = ~((inputs[21]) | (inputs[31]));
    assign layer0_outputs[10084] = ~((inputs[25]) & (inputs[58]));
    assign layer0_outputs[10085] = (inputs[227]) | (inputs[99]);
    assign layer0_outputs[10086] = ~(inputs[196]);
    assign layer0_outputs[10087] = ~(inputs[144]);
    assign layer0_outputs[10088] = inputs[29];
    assign layer0_outputs[10089] = ~((inputs[109]) ^ (inputs[190]));
    assign layer0_outputs[10090] = inputs[82];
    assign layer0_outputs[10091] = ~(inputs[31]) | (inputs[240]);
    assign layer0_outputs[10092] = inputs[73];
    assign layer0_outputs[10093] = inputs[83];
    assign layer0_outputs[10094] = ~((inputs[47]) | (inputs[203]));
    assign layer0_outputs[10095] = inputs[228];
    assign layer0_outputs[10096] = ~((inputs[135]) & (inputs[69]));
    assign layer0_outputs[10097] = ~(inputs[95]) | (inputs[65]);
    assign layer0_outputs[10098] = ~((inputs[165]) | (inputs[249]));
    assign layer0_outputs[10099] = (inputs[220]) | (inputs[207]);
    assign layer0_outputs[10100] = ~(inputs[210]);
    assign layer0_outputs[10101] = inputs[223];
    assign layer0_outputs[10102] = (inputs[97]) & ~(inputs[151]);
    assign layer0_outputs[10103] = ~(inputs[37]);
    assign layer0_outputs[10104] = ~(inputs[179]) | (inputs[62]);
    assign layer0_outputs[10105] = (inputs[1]) & ~(inputs[119]);
    assign layer0_outputs[10106] = (inputs[62]) & ~(inputs[155]);
    assign layer0_outputs[10107] = ~((inputs[141]) | (inputs[37]));
    assign layer0_outputs[10108] = inputs[163];
    assign layer0_outputs[10109] = ~(inputs[124]) | (inputs[169]);
    assign layer0_outputs[10110] = ~((inputs[98]) ^ (inputs[21]));
    assign layer0_outputs[10111] = inputs[63];
    assign layer0_outputs[10112] = ~(inputs[71]);
    assign layer0_outputs[10113] = ~(inputs[214]) | (inputs[57]);
    assign layer0_outputs[10114] = (inputs[183]) & ~(inputs[175]);
    assign layer0_outputs[10115] = (inputs[143]) | (inputs[149]);
    assign layer0_outputs[10116] = (inputs[245]) & ~(inputs[113]);
    assign layer0_outputs[10117] = inputs[76];
    assign layer0_outputs[10118] = (inputs[218]) & ~(inputs[239]);
    assign layer0_outputs[10119] = (inputs[217]) | (inputs[252]);
    assign layer0_outputs[10120] = ~(inputs[96]);
    assign layer0_outputs[10121] = ~(inputs[36]) | (inputs[99]);
    assign layer0_outputs[10122] = ~((inputs[96]) & (inputs[109]));
    assign layer0_outputs[10123] = ~(inputs[240]);
    assign layer0_outputs[10124] = ~((inputs[179]) ^ (inputs[247]));
    assign layer0_outputs[10125] = inputs[243];
    assign layer0_outputs[10126] = ~((inputs[253]) ^ (inputs[145]));
    assign layer0_outputs[10127] = (inputs[86]) & ~(inputs[170]);
    assign layer0_outputs[10128] = (inputs[178]) ^ (inputs[247]);
    assign layer0_outputs[10129] = (inputs[211]) ^ (inputs[15]);
    assign layer0_outputs[10130] = ~((inputs[202]) ^ (inputs[234]));
    assign layer0_outputs[10131] = (inputs[157]) ^ (inputs[8]);
    assign layer0_outputs[10132] = (inputs[121]) | (inputs[91]);
    assign layer0_outputs[10133] = ~((inputs[113]) | (inputs[122]));
    assign layer0_outputs[10134] = ~(inputs[76]);
    assign layer0_outputs[10135] = ~((inputs[204]) ^ (inputs[144]));
    assign layer0_outputs[10136] = 1'b1;
    assign layer0_outputs[10137] = (inputs[226]) | (inputs[5]);
    assign layer0_outputs[10138] = 1'b1;
    assign layer0_outputs[10139] = ~((inputs[71]) ^ (inputs[84]));
    assign layer0_outputs[10140] = (inputs[47]) & ~(inputs[184]);
    assign layer0_outputs[10141] = (inputs[11]) & ~(inputs[68]);
    assign layer0_outputs[10142] = inputs[31];
    assign layer0_outputs[10143] = (inputs[158]) & ~(inputs[47]);
    assign layer0_outputs[10144] = (inputs[160]) ^ (inputs[39]);
    assign layer0_outputs[10145] = (inputs[234]) & ~(inputs[0]);
    assign layer0_outputs[10146] = ~((inputs[164]) ^ (inputs[135]));
    assign layer0_outputs[10147] = inputs[83];
    assign layer0_outputs[10148] = ~(inputs[42]) | (inputs[106]);
    assign layer0_outputs[10149] = ~((inputs[47]) | (inputs[13]));
    assign layer0_outputs[10150] = inputs[191];
    assign layer0_outputs[10151] = ~(inputs[122]) | (inputs[174]);
    assign layer0_outputs[10152] = ~((inputs[242]) & (inputs[186]));
    assign layer0_outputs[10153] = inputs[92];
    assign layer0_outputs[10154] = ~((inputs[171]) | (inputs[221]));
    assign layer0_outputs[10155] = ~(inputs[142]);
    assign layer0_outputs[10156] = ~(inputs[177]) | (inputs[10]);
    assign layer0_outputs[10157] = (inputs[75]) ^ (inputs[175]);
    assign layer0_outputs[10158] = (inputs[31]) ^ (inputs[156]);
    assign layer0_outputs[10159] = ~((inputs[133]) | (inputs[30]));
    assign layer0_outputs[10160] = inputs[137];
    assign layer0_outputs[10161] = inputs[246];
    assign layer0_outputs[10162] = (inputs[116]) & ~(inputs[55]);
    assign layer0_outputs[10163] = ~(inputs[114]);
    assign layer0_outputs[10164] = (inputs[145]) | (inputs[89]);
    assign layer0_outputs[10165] = ~(inputs[33]) | (inputs[253]);
    assign layer0_outputs[10166] = ~(inputs[103]);
    assign layer0_outputs[10167] = inputs[161];
    assign layer0_outputs[10168] = ~(inputs[155]);
    assign layer0_outputs[10169] = (inputs[180]) | (inputs[114]);
    assign layer0_outputs[10170] = ~(inputs[149]);
    assign layer0_outputs[10171] = inputs[102];
    assign layer0_outputs[10172] = (inputs[74]) & ~(inputs[141]);
    assign layer0_outputs[10173] = (inputs[219]) | (inputs[251]);
    assign layer0_outputs[10174] = ~((inputs[203]) ^ (inputs[252]));
    assign layer0_outputs[10175] = ~((inputs[233]) | (inputs[39]));
    assign layer0_outputs[10176] = ~(inputs[179]);
    assign layer0_outputs[10177] = (inputs[22]) & ~(inputs[160]);
    assign layer0_outputs[10178] = ~(inputs[149]);
    assign layer0_outputs[10179] = (inputs[186]) & ~(inputs[69]);
    assign layer0_outputs[10180] = ~((inputs[52]) ^ (inputs[117]));
    assign layer0_outputs[10181] = ~(inputs[24]);
    assign layer0_outputs[10182] = inputs[113];
    assign layer0_outputs[10183] = ~((inputs[182]) | (inputs[146]));
    assign layer0_outputs[10184] = ~(inputs[58]) | (inputs[210]);
    assign layer0_outputs[10185] = ~((inputs[164]) | (inputs[56]));
    assign layer0_outputs[10186] = (inputs[215]) ^ (inputs[246]);
    assign layer0_outputs[10187] = ~((inputs[128]) | (inputs[27]));
    assign layer0_outputs[10188] = (inputs[100]) & (inputs[122]);
    assign layer0_outputs[10189] = (inputs[209]) & ~(inputs[15]);
    assign layer0_outputs[10190] = (inputs[33]) & (inputs[48]);
    assign layer0_outputs[10191] = ~((inputs[67]) ^ (inputs[124]));
    assign layer0_outputs[10192] = ~(inputs[57]) | (inputs[183]);
    assign layer0_outputs[10193] = ~(inputs[89]);
    assign layer0_outputs[10194] = inputs[165];
    assign layer0_outputs[10195] = 1'b1;
    assign layer0_outputs[10196] = ~((inputs[232]) | (inputs[211]));
    assign layer0_outputs[10197] = ~((inputs[117]) & (inputs[170]));
    assign layer0_outputs[10198] = ~((inputs[26]) | (inputs[7]));
    assign layer0_outputs[10199] = inputs[68];
    assign layer0_outputs[10200] = inputs[24];
    assign layer0_outputs[10201] = (inputs[165]) & ~(inputs[62]);
    assign layer0_outputs[10202] = ~((inputs[58]) | (inputs[124]));
    assign layer0_outputs[10203] = (inputs[35]) | (inputs[37]);
    assign layer0_outputs[10204] = ~(inputs[176]) | (inputs[48]);
    assign layer0_outputs[10205] = ~(inputs[207]);
    assign layer0_outputs[10206] = 1'b1;
    assign layer0_outputs[10207] = ~((inputs[50]) | (inputs[172]));
    assign layer0_outputs[10208] = ~(inputs[77]) | (inputs[15]);
    assign layer0_outputs[10209] = inputs[0];
    assign layer0_outputs[10210] = ~((inputs[185]) ^ (inputs[198]));
    assign layer0_outputs[10211] = ~(inputs[237]);
    assign layer0_outputs[10212] = ~((inputs[160]) | (inputs[221]));
    assign layer0_outputs[10213] = (inputs[30]) | (inputs[207]);
    assign layer0_outputs[10214] = ~((inputs[126]) ^ (inputs[89]));
    assign layer0_outputs[10215] = inputs[224];
    assign layer0_outputs[10216] = inputs[1];
    assign layer0_outputs[10217] = ~((inputs[225]) ^ (inputs[248]));
    assign layer0_outputs[10218] = ~(inputs[255]);
    assign layer0_outputs[10219] = ~(inputs[166]);
    assign layer0_outputs[10220] = ~(inputs[43]) | (inputs[193]);
    assign layer0_outputs[10221] = inputs[209];
    assign layer0_outputs[10222] = ~(inputs[62]);
    assign layer0_outputs[10223] = ~(inputs[116]);
    assign layer0_outputs[10224] = ~(inputs[222]) | (inputs[116]);
    assign layer0_outputs[10225] = (inputs[217]) & (inputs[207]);
    assign layer0_outputs[10226] = ~(inputs[119]);
    assign layer0_outputs[10227] = ~(inputs[82]);
    assign layer0_outputs[10228] = ~((inputs[194]) & (inputs[231]));
    assign layer0_outputs[10229] = (inputs[126]) & ~(inputs[12]);
    assign layer0_outputs[10230] = 1'b0;
    assign layer0_outputs[10231] = (inputs[93]) | (inputs[171]);
    assign layer0_outputs[10232] = inputs[179];
    assign layer0_outputs[10233] = ~(inputs[10]) | (inputs[152]);
    assign layer0_outputs[10234] = inputs[94];
    assign layer0_outputs[10235] = 1'b1;
    assign layer0_outputs[10236] = ~((inputs[148]) ^ (inputs[68]));
    assign layer0_outputs[10237] = (inputs[215]) & ~(inputs[84]);
    assign layer0_outputs[10238] = inputs[197];
    assign layer0_outputs[10239] = ~(inputs[82]);
    assign layer0_outputs[10240] = (inputs[117]) ^ (inputs[87]);
    assign layer0_outputs[10241] = (inputs[247]) | (inputs[91]);
    assign layer0_outputs[10242] = ~(inputs[93]);
    assign layer0_outputs[10243] = inputs[216];
    assign layer0_outputs[10244] = ~(inputs[217]) | (inputs[141]);
    assign layer0_outputs[10245] = inputs[162];
    assign layer0_outputs[10246] = ~(inputs[99]) | (inputs[191]);
    assign layer0_outputs[10247] = inputs[93];
    assign layer0_outputs[10248] = ~(inputs[4]);
    assign layer0_outputs[10249] = ~(inputs[212]);
    assign layer0_outputs[10250] = ~((inputs[161]) | (inputs[172]));
    assign layer0_outputs[10251] = inputs[194];
    assign layer0_outputs[10252] = (inputs[203]) | (inputs[212]);
    assign layer0_outputs[10253] = inputs[76];
    assign layer0_outputs[10254] = 1'b0;
    assign layer0_outputs[10255] = ~((inputs[121]) | (inputs[165]));
    assign layer0_outputs[10256] = (inputs[146]) & ~(inputs[85]);
    assign layer0_outputs[10257] = (inputs[175]) ^ (inputs[54]);
    assign layer0_outputs[10258] = ~(inputs[26]) | (inputs[248]);
    assign layer0_outputs[10259] = inputs[67];
    assign layer0_outputs[10260] = (inputs[212]) & ~(inputs[9]);
    assign layer0_outputs[10261] = ~(inputs[96]);
    assign layer0_outputs[10262] = 1'b0;
    assign layer0_outputs[10263] = ~(inputs[26]) | (inputs[237]);
    assign layer0_outputs[10264] = inputs[122];
    assign layer0_outputs[10265] = ~(inputs[115]) | (inputs[233]);
    assign layer0_outputs[10266] = ~((inputs[65]) ^ (inputs[37]));
    assign layer0_outputs[10267] = (inputs[9]) & (inputs[26]);
    assign layer0_outputs[10268] = ~(inputs[78]);
    assign layer0_outputs[10269] = ~(inputs[195]) | (inputs[159]);
    assign layer0_outputs[10270] = (inputs[196]) ^ (inputs[2]);
    assign layer0_outputs[10271] = (inputs[19]) | (inputs[207]);
    assign layer0_outputs[10272] = ~((inputs[42]) | (inputs[63]));
    assign layer0_outputs[10273] = (inputs[44]) ^ (inputs[63]);
    assign layer0_outputs[10274] = (inputs[172]) & ~(inputs[13]);
    assign layer0_outputs[10275] = inputs[64];
    assign layer0_outputs[10276] = ~((inputs[49]) | (inputs[84]));
    assign layer0_outputs[10277] = (inputs[132]) & ~(inputs[185]);
    assign layer0_outputs[10278] = 1'b0;
    assign layer0_outputs[10279] = ~(inputs[162]) | (inputs[93]);
    assign layer0_outputs[10280] = inputs[69];
    assign layer0_outputs[10281] = (inputs[198]) ^ (inputs[137]);
    assign layer0_outputs[10282] = ~(inputs[203]);
    assign layer0_outputs[10283] = ~((inputs[130]) | (inputs[161]));
    assign layer0_outputs[10284] = ~(inputs[113]);
    assign layer0_outputs[10285] = (inputs[22]) & ~(inputs[222]);
    assign layer0_outputs[10286] = ~(inputs[246]);
    assign layer0_outputs[10287] = inputs[125];
    assign layer0_outputs[10288] = (inputs[20]) & ~(inputs[28]);
    assign layer0_outputs[10289] = 1'b1;
    assign layer0_outputs[10290] = ~((inputs[253]) | (inputs[107]));
    assign layer0_outputs[10291] = (inputs[243]) ^ (inputs[212]);
    assign layer0_outputs[10292] = ~((inputs[253]) | (inputs[32]));
    assign layer0_outputs[10293] = ~(inputs[159]);
    assign layer0_outputs[10294] = (inputs[5]) | (inputs[166]);
    assign layer0_outputs[10295] = ~((inputs[87]) & (inputs[124]));
    assign layer0_outputs[10296] = (inputs[89]) & ~(inputs[53]);
    assign layer0_outputs[10297] = inputs[77];
    assign layer0_outputs[10298] = ~((inputs[135]) | (inputs[71]));
    assign layer0_outputs[10299] = (inputs[96]) | (inputs[66]);
    assign layer0_outputs[10300] = ~((inputs[94]) ^ (inputs[197]));
    assign layer0_outputs[10301] = ~(inputs[234]);
    assign layer0_outputs[10302] = ~((inputs[142]) | (inputs[85]));
    assign layer0_outputs[10303] = 1'b0;
    assign layer0_outputs[10304] = (inputs[69]) & ~(inputs[145]);
    assign layer0_outputs[10305] = (inputs[26]) | (inputs[16]);
    assign layer0_outputs[10306] = inputs[156];
    assign layer0_outputs[10307] = ~((inputs[170]) ^ (inputs[109]));
    assign layer0_outputs[10308] = (inputs[231]) & (inputs[189]);
    assign layer0_outputs[10309] = ~((inputs[172]) ^ (inputs[48]));
    assign layer0_outputs[10310] = ~(inputs[74]);
    assign layer0_outputs[10311] = ~(inputs[168]);
    assign layer0_outputs[10312] = ~((inputs[182]) | (inputs[99]));
    assign layer0_outputs[10313] = ~((inputs[117]) ^ (inputs[217]));
    assign layer0_outputs[10314] = inputs[154];
    assign layer0_outputs[10315] = ~((inputs[35]) | (inputs[102]));
    assign layer0_outputs[10316] = (inputs[108]) & (inputs[200]);
    assign layer0_outputs[10317] = (inputs[228]) | (inputs[197]);
    assign layer0_outputs[10318] = inputs[180];
    assign layer0_outputs[10319] = inputs[202];
    assign layer0_outputs[10320] = ~(inputs[219]) | (inputs[69]);
    assign layer0_outputs[10321] = ~(inputs[124]);
    assign layer0_outputs[10322] = inputs[31];
    assign layer0_outputs[10323] = (inputs[125]) | (inputs[106]);
    assign layer0_outputs[10324] = ~((inputs[130]) | (inputs[175]));
    assign layer0_outputs[10325] = ~(inputs[126]);
    assign layer0_outputs[10326] = ~(inputs[221]);
    assign layer0_outputs[10327] = ~(inputs[133]);
    assign layer0_outputs[10328] = ~(inputs[83]) | (inputs[169]);
    assign layer0_outputs[10329] = (inputs[19]) | (inputs[32]);
    assign layer0_outputs[10330] = (inputs[216]) & ~(inputs[60]);
    assign layer0_outputs[10331] = (inputs[217]) | (inputs[63]);
    assign layer0_outputs[10332] = inputs[173];
    assign layer0_outputs[10333] = ~((inputs[159]) ^ (inputs[161]));
    assign layer0_outputs[10334] = ~((inputs[170]) | (inputs[203]));
    assign layer0_outputs[10335] = ~(inputs[157]) | (inputs[26]);
    assign layer0_outputs[10336] = ~((inputs[3]) ^ (inputs[209]));
    assign layer0_outputs[10337] = ~(inputs[173]);
    assign layer0_outputs[10338] = ~(inputs[109]) | (inputs[52]);
    assign layer0_outputs[10339] = ~(inputs[183]) | (inputs[68]);
    assign layer0_outputs[10340] = ~((inputs[78]) | (inputs[119]));
    assign layer0_outputs[10341] = (inputs[104]) | (inputs[87]);
    assign layer0_outputs[10342] = ~((inputs[52]) & (inputs[154]));
    assign layer0_outputs[10343] = ~((inputs[61]) | (inputs[142]));
    assign layer0_outputs[10344] = ~(inputs[132]) | (inputs[3]);
    assign layer0_outputs[10345] = (inputs[193]) & ~(inputs[91]);
    assign layer0_outputs[10346] = ~(inputs[45]);
    assign layer0_outputs[10347] = inputs[5];
    assign layer0_outputs[10348] = ~(inputs[138]) | (inputs[65]);
    assign layer0_outputs[10349] = ~((inputs[204]) ^ (inputs[79]));
    assign layer0_outputs[10350] = inputs[135];
    assign layer0_outputs[10351] = inputs[60];
    assign layer0_outputs[10352] = ~((inputs[107]) & (inputs[133]));
    assign layer0_outputs[10353] = ~(inputs[255]) | (inputs[113]);
    assign layer0_outputs[10354] = inputs[233];
    assign layer0_outputs[10355] = (inputs[10]) & ~(inputs[119]);
    assign layer0_outputs[10356] = (inputs[59]) & ~(inputs[236]);
    assign layer0_outputs[10357] = ~((inputs[105]) & (inputs[122]));
    assign layer0_outputs[10358] = (inputs[226]) | (inputs[17]);
    assign layer0_outputs[10359] = ~((inputs[204]) & (inputs[56]));
    assign layer0_outputs[10360] = ~(inputs[133]) | (inputs[4]);
    assign layer0_outputs[10361] = (inputs[162]) & ~(inputs[76]);
    assign layer0_outputs[10362] = ~(inputs[115]);
    assign layer0_outputs[10363] = inputs[92];
    assign layer0_outputs[10364] = ~((inputs[7]) & (inputs[228]));
    assign layer0_outputs[10365] = (inputs[223]) ^ (inputs[51]);
    assign layer0_outputs[10366] = (inputs[91]) & ~(inputs[116]);
    assign layer0_outputs[10367] = ~((inputs[229]) | (inputs[225]));
    assign layer0_outputs[10368] = ~(inputs[175]);
    assign layer0_outputs[10369] = 1'b1;
    assign layer0_outputs[10370] = (inputs[98]) & ~(inputs[87]);
    assign layer0_outputs[10371] = (inputs[90]) | (inputs[115]);
    assign layer0_outputs[10372] = ~(inputs[251]) | (inputs[172]);
    assign layer0_outputs[10373] = ~(inputs[182]) | (inputs[67]);
    assign layer0_outputs[10374] = ~(inputs[167]);
    assign layer0_outputs[10375] = ~(inputs[202]);
    assign layer0_outputs[10376] = ~((inputs[105]) | (inputs[160]));
    assign layer0_outputs[10377] = (inputs[163]) & ~(inputs[224]);
    assign layer0_outputs[10378] = ~((inputs[17]) | (inputs[143]));
    assign layer0_outputs[10379] = 1'b1;
    assign layer0_outputs[10380] = (inputs[230]) & (inputs[165]);
    assign layer0_outputs[10381] = inputs[226];
    assign layer0_outputs[10382] = inputs[96];
    assign layer0_outputs[10383] = ~(inputs[63]) | (inputs[254]);
    assign layer0_outputs[10384] = ~(inputs[3]);
    assign layer0_outputs[10385] = inputs[120];
    assign layer0_outputs[10386] = ~(inputs[215]);
    assign layer0_outputs[10387] = ~(inputs[118]) | (inputs[85]);
    assign layer0_outputs[10388] = ~((inputs[48]) | (inputs[174]));
    assign layer0_outputs[10389] = (inputs[73]) | (inputs[3]);
    assign layer0_outputs[10390] = (inputs[28]) & ~(inputs[241]);
    assign layer0_outputs[10391] = ~(inputs[26]);
    assign layer0_outputs[10392] = (inputs[192]) | (inputs[4]);
    assign layer0_outputs[10393] = (inputs[246]) | (inputs[154]);
    assign layer0_outputs[10394] = (inputs[227]) & (inputs[180]);
    assign layer0_outputs[10395] = (inputs[136]) & ~(inputs[63]);
    assign layer0_outputs[10396] = (inputs[192]) ^ (inputs[250]);
    assign layer0_outputs[10397] = ~((inputs[55]) | (inputs[95]));
    assign layer0_outputs[10398] = (inputs[148]) & ~(inputs[137]);
    assign layer0_outputs[10399] = ~((inputs[13]) | (inputs[52]));
    assign layer0_outputs[10400] = (inputs[131]) & ~(inputs[120]);
    assign layer0_outputs[10401] = ~((inputs[129]) ^ (inputs[103]));
    assign layer0_outputs[10402] = (inputs[251]) ^ (inputs[107]);
    assign layer0_outputs[10403] = 1'b1;
    assign layer0_outputs[10404] = ~(inputs[198]);
    assign layer0_outputs[10405] = (inputs[170]) & ~(inputs[87]);
    assign layer0_outputs[10406] = (inputs[218]) & ~(inputs[18]);
    assign layer0_outputs[10407] = ~(inputs[251]) | (inputs[242]);
    assign layer0_outputs[10408] = (inputs[213]) & ~(inputs[158]);
    assign layer0_outputs[10409] = ~(inputs[88]);
    assign layer0_outputs[10410] = ~(inputs[42]) | (inputs[190]);
    assign layer0_outputs[10411] = (inputs[138]) ^ (inputs[135]);
    assign layer0_outputs[10412] = inputs[248];
    assign layer0_outputs[10413] = (inputs[224]) | (inputs[2]);
    assign layer0_outputs[10414] = 1'b1;
    assign layer0_outputs[10415] = ~((inputs[40]) | (inputs[1]));
    assign layer0_outputs[10416] = inputs[163];
    assign layer0_outputs[10417] = ~(inputs[86]);
    assign layer0_outputs[10418] = 1'b0;
    assign layer0_outputs[10419] = ~((inputs[23]) | (inputs[36]));
    assign layer0_outputs[10420] = (inputs[94]) & (inputs[136]);
    assign layer0_outputs[10421] = ~(inputs[195]) | (inputs[136]);
    assign layer0_outputs[10422] = inputs[19];
    assign layer0_outputs[10423] = ~((inputs[40]) & (inputs[71]));
    assign layer0_outputs[10424] = ~((inputs[63]) ^ (inputs[29]));
    assign layer0_outputs[10425] = inputs[238];
    assign layer0_outputs[10426] = (inputs[122]) & ~(inputs[1]);
    assign layer0_outputs[10427] = ~(inputs[37]) | (inputs[254]);
    assign layer0_outputs[10428] = (inputs[45]) | (inputs[208]);
    assign layer0_outputs[10429] = ~(inputs[183]);
    assign layer0_outputs[10430] = ~(inputs[216]);
    assign layer0_outputs[10431] = (inputs[202]) ^ (inputs[185]);
    assign layer0_outputs[10432] = ~((inputs[87]) ^ (inputs[162]));
    assign layer0_outputs[10433] = inputs[94];
    assign layer0_outputs[10434] = ~((inputs[158]) ^ (inputs[116]));
    assign layer0_outputs[10435] = (inputs[59]) | (inputs[123]);
    assign layer0_outputs[10436] = (inputs[36]) & ~(inputs[103]);
    assign layer0_outputs[10437] = ~((inputs[193]) | (inputs[22]));
    assign layer0_outputs[10438] = inputs[105];
    assign layer0_outputs[10439] = (inputs[168]) | (inputs[72]);
    assign layer0_outputs[10440] = ~((inputs[63]) | (inputs[70]));
    assign layer0_outputs[10441] = ~(inputs[44]) | (inputs[238]);
    assign layer0_outputs[10442] = ~(inputs[240]) | (inputs[175]);
    assign layer0_outputs[10443] = ~((inputs[221]) & (inputs[249]));
    assign layer0_outputs[10444] = ~((inputs[5]) ^ (inputs[45]));
    assign layer0_outputs[10445] = (inputs[153]) & ~(inputs[24]);
    assign layer0_outputs[10446] = (inputs[252]) | (inputs[150]);
    assign layer0_outputs[10447] = ~((inputs[205]) | (inputs[175]));
    assign layer0_outputs[10448] = (inputs[219]) & ~(inputs[120]);
    assign layer0_outputs[10449] = inputs[212];
    assign layer0_outputs[10450] = ~((inputs[1]) ^ (inputs[140]));
    assign layer0_outputs[10451] = inputs[163];
    assign layer0_outputs[10452] = (inputs[250]) ^ (inputs[162]);
    assign layer0_outputs[10453] = (inputs[234]) ^ (inputs[74]);
    assign layer0_outputs[10454] = (inputs[242]) | (inputs[167]);
    assign layer0_outputs[10455] = ~(inputs[43]) | (inputs[200]);
    assign layer0_outputs[10456] = inputs[173];
    assign layer0_outputs[10457] = ~(inputs[229]) | (inputs[106]);
    assign layer0_outputs[10458] = (inputs[125]) & ~(inputs[200]);
    assign layer0_outputs[10459] = (inputs[227]) & ~(inputs[81]);
    assign layer0_outputs[10460] = (inputs[137]) ^ (inputs[101]);
    assign layer0_outputs[10461] = (inputs[207]) | (inputs[7]);
    assign layer0_outputs[10462] = 1'b1;
    assign layer0_outputs[10463] = (inputs[183]) & ~(inputs[13]);
    assign layer0_outputs[10464] = ~(inputs[52]) | (inputs[71]);
    assign layer0_outputs[10465] = inputs[64];
    assign layer0_outputs[10466] = (inputs[70]) | (inputs[58]);
    assign layer0_outputs[10467] = ~((inputs[239]) | (inputs[159]));
    assign layer0_outputs[10468] = ~((inputs[193]) & (inputs[200]));
    assign layer0_outputs[10469] = 1'b1;
    assign layer0_outputs[10470] = (inputs[108]) & ~(inputs[48]);
    assign layer0_outputs[10471] = ~(inputs[104]);
    assign layer0_outputs[10472] = ~(inputs[139]) | (inputs[8]);
    assign layer0_outputs[10473] = inputs[76];
    assign layer0_outputs[10474] = (inputs[49]) ^ (inputs[22]);
    assign layer0_outputs[10475] = (inputs[244]) | (inputs[164]);
    assign layer0_outputs[10476] = 1'b1;
    assign layer0_outputs[10477] = ~((inputs[9]) | (inputs[12]));
    assign layer0_outputs[10478] = ~((inputs[212]) | (inputs[192]));
    assign layer0_outputs[10479] = ~(inputs[58]);
    assign layer0_outputs[10480] = (inputs[103]) & ~(inputs[42]);
    assign layer0_outputs[10481] = ~((inputs[209]) ^ (inputs[254]));
    assign layer0_outputs[10482] = ~(inputs[113]);
    assign layer0_outputs[10483] = ~(inputs[155]) | (inputs[31]);
    assign layer0_outputs[10484] = ~(inputs[225]);
    assign layer0_outputs[10485] = ~((inputs[125]) ^ (inputs[189]));
    assign layer0_outputs[10486] = (inputs[141]) | (inputs[218]);
    assign layer0_outputs[10487] = (inputs[122]) & ~(inputs[32]);
    assign layer0_outputs[10488] = (inputs[178]) | (inputs[241]);
    assign layer0_outputs[10489] = (inputs[40]) & (inputs[218]);
    assign layer0_outputs[10490] = ~((inputs[129]) ^ (inputs[223]));
    assign layer0_outputs[10491] = (inputs[249]) & ~(inputs[111]);
    assign layer0_outputs[10492] = (inputs[153]) & ~(inputs[72]);
    assign layer0_outputs[10493] = ~(inputs[235]) | (inputs[7]);
    assign layer0_outputs[10494] = ~(inputs[210]);
    assign layer0_outputs[10495] = ~((inputs[116]) | (inputs[6]));
    assign layer0_outputs[10496] = (inputs[178]) & ~(inputs[46]);
    assign layer0_outputs[10497] = ~(inputs[173]) | (inputs[42]);
    assign layer0_outputs[10498] = ~(inputs[119]);
    assign layer0_outputs[10499] = ~(inputs[108]) | (inputs[151]);
    assign layer0_outputs[10500] = ~((inputs[39]) | (inputs[5]));
    assign layer0_outputs[10501] = ~(inputs[4]);
    assign layer0_outputs[10502] = (inputs[166]) & ~(inputs[157]);
    assign layer0_outputs[10503] = inputs[77];
    assign layer0_outputs[10504] = ~(inputs[189]);
    assign layer0_outputs[10505] = 1'b1;
    assign layer0_outputs[10506] = ~((inputs[17]) & (inputs[117]));
    assign layer0_outputs[10507] = ~(inputs[219]) | (inputs[26]);
    assign layer0_outputs[10508] = ~((inputs[246]) | (inputs[144]));
    assign layer0_outputs[10509] = (inputs[21]) ^ (inputs[37]);
    assign layer0_outputs[10510] = (inputs[174]) ^ (inputs[179]);
    assign layer0_outputs[10511] = inputs[105];
    assign layer0_outputs[10512] = (inputs[131]) & ~(inputs[153]);
    assign layer0_outputs[10513] = ~(inputs[14]);
    assign layer0_outputs[10514] = ~((inputs[67]) | (inputs[146]));
    assign layer0_outputs[10515] = ~((inputs[237]) | (inputs[50]));
    assign layer0_outputs[10516] = (inputs[194]) ^ (inputs[219]);
    assign layer0_outputs[10517] = ~(inputs[153]) | (inputs[108]);
    assign layer0_outputs[10518] = ~(inputs[61]);
    assign layer0_outputs[10519] = inputs[24];
    assign layer0_outputs[10520] = ~(inputs[109]);
    assign layer0_outputs[10521] = 1'b0;
    assign layer0_outputs[10522] = (inputs[229]) | (inputs[191]);
    assign layer0_outputs[10523] = (inputs[204]) ^ (inputs[224]);
    assign layer0_outputs[10524] = ~(inputs[144]) | (inputs[255]);
    assign layer0_outputs[10525] = ~(inputs[16]);
    assign layer0_outputs[10526] = ~((inputs[96]) ^ (inputs[139]));
    assign layer0_outputs[10527] = ~((inputs[30]) | (inputs[33]));
    assign layer0_outputs[10528] = inputs[106];
    assign layer0_outputs[10529] = (inputs[85]) & ~(inputs[77]);
    assign layer0_outputs[10530] = ~((inputs[75]) ^ (inputs[19]));
    assign layer0_outputs[10531] = (inputs[83]) | (inputs[233]);
    assign layer0_outputs[10532] = ~((inputs[91]) | (inputs[111]));
    assign layer0_outputs[10533] = 1'b1;
    assign layer0_outputs[10534] = ~((inputs[131]) ^ (inputs[145]));
    assign layer0_outputs[10535] = inputs[29];
    assign layer0_outputs[10536] = ~((inputs[137]) & (inputs[174]));
    assign layer0_outputs[10537] = (inputs[107]) ^ (inputs[75]);
    assign layer0_outputs[10538] = ~((inputs[169]) ^ (inputs[123]));
    assign layer0_outputs[10539] = (inputs[159]) & ~(inputs[252]);
    assign layer0_outputs[10540] = (inputs[178]) ^ (inputs[244]);
    assign layer0_outputs[10541] = ~(inputs[7]);
    assign layer0_outputs[10542] = ~(inputs[114]);
    assign layer0_outputs[10543] = ~(inputs[204]);
    assign layer0_outputs[10544] = ~(inputs[232]) | (inputs[97]);
    assign layer0_outputs[10545] = ~((inputs[112]) ^ (inputs[119]));
    assign layer0_outputs[10546] = ~(inputs[18]);
    assign layer0_outputs[10547] = ~((inputs[174]) ^ (inputs[17]));
    assign layer0_outputs[10548] = ~(inputs[198]);
    assign layer0_outputs[10549] = (inputs[140]) | (inputs[73]);
    assign layer0_outputs[10550] = inputs[152];
    assign layer0_outputs[10551] = ~((inputs[221]) | (inputs[13]));
    assign layer0_outputs[10552] = ~(inputs[56]);
    assign layer0_outputs[10553] = (inputs[28]) ^ (inputs[154]);
    assign layer0_outputs[10554] = (inputs[79]) ^ (inputs[206]);
    assign layer0_outputs[10555] = ~((inputs[27]) | (inputs[107]));
    assign layer0_outputs[10556] = ~(inputs[2]) | (inputs[159]);
    assign layer0_outputs[10557] = (inputs[21]) | (inputs[253]);
    assign layer0_outputs[10558] = (inputs[99]) & (inputs[152]);
    assign layer0_outputs[10559] = (inputs[181]) & ~(inputs[36]);
    assign layer0_outputs[10560] = ~(inputs[216]);
    assign layer0_outputs[10561] = ~(inputs[169]) | (inputs[4]);
    assign layer0_outputs[10562] = ~((inputs[116]) ^ (inputs[160]));
    assign layer0_outputs[10563] = ~(inputs[56]) | (inputs[18]);
    assign layer0_outputs[10564] = (inputs[71]) ^ (inputs[188]);
    assign layer0_outputs[10565] = ~((inputs[175]) ^ (inputs[36]));
    assign layer0_outputs[10566] = ~((inputs[125]) ^ (inputs[153]));
    assign layer0_outputs[10567] = ~((inputs[76]) & (inputs[90]));
    assign layer0_outputs[10568] = ~(inputs[30]);
    assign layer0_outputs[10569] = ~((inputs[92]) & (inputs[138]));
    assign layer0_outputs[10570] = (inputs[15]) & ~(inputs[201]);
    assign layer0_outputs[10571] = ~(inputs[208]) | (inputs[226]);
    assign layer0_outputs[10572] = ~((inputs[100]) ^ (inputs[118]));
    assign layer0_outputs[10573] = (inputs[94]) ^ (inputs[66]);
    assign layer0_outputs[10574] = (inputs[199]) & ~(inputs[113]);
    assign layer0_outputs[10575] = ~((inputs[103]) | (inputs[36]));
    assign layer0_outputs[10576] = (inputs[166]) & ~(inputs[18]);
    assign layer0_outputs[10577] = inputs[129];
    assign layer0_outputs[10578] = ~(inputs[51]) | (inputs[147]);
    assign layer0_outputs[10579] = ~(inputs[51]) | (inputs[198]);
    assign layer0_outputs[10580] = (inputs[104]) | (inputs[67]);
    assign layer0_outputs[10581] = (inputs[254]) ^ (inputs[181]);
    assign layer0_outputs[10582] = ~(inputs[136]);
    assign layer0_outputs[10583] = (inputs[184]) & (inputs[210]);
    assign layer0_outputs[10584] = ~(inputs[199]) | (inputs[139]);
    assign layer0_outputs[10585] = ~(inputs[72]) | (inputs[1]);
    assign layer0_outputs[10586] = (inputs[231]) & (inputs[188]);
    assign layer0_outputs[10587] = (inputs[251]) ^ (inputs[166]);
    assign layer0_outputs[10588] = ~(inputs[129]);
    assign layer0_outputs[10589] = ~(inputs[133]) | (inputs[18]);
    assign layer0_outputs[10590] = 1'b0;
    assign layer0_outputs[10591] = (inputs[130]) & ~(inputs[195]);
    assign layer0_outputs[10592] = 1'b1;
    assign layer0_outputs[10593] = inputs[237];
    assign layer0_outputs[10594] = 1'b0;
    assign layer0_outputs[10595] = inputs[19];
    assign layer0_outputs[10596] = (inputs[33]) | (inputs[208]);
    assign layer0_outputs[10597] = ~(inputs[119]);
    assign layer0_outputs[10598] = ~((inputs[146]) ^ (inputs[165]));
    assign layer0_outputs[10599] = 1'b1;
    assign layer0_outputs[10600] = ~((inputs[158]) | (inputs[235]));
    assign layer0_outputs[10601] = (inputs[113]) & (inputs[217]);
    assign layer0_outputs[10602] = inputs[136];
    assign layer0_outputs[10603] = (inputs[216]) | (inputs[171]);
    assign layer0_outputs[10604] = 1'b1;
    assign layer0_outputs[10605] = ~(inputs[78]) | (inputs[112]);
    assign layer0_outputs[10606] = (inputs[158]) & ~(inputs[205]);
    assign layer0_outputs[10607] = inputs[8];
    assign layer0_outputs[10608] = ~(inputs[107]) | (inputs[14]);
    assign layer0_outputs[10609] = inputs[209];
    assign layer0_outputs[10610] = inputs[133];
    assign layer0_outputs[10611] = (inputs[80]) | (inputs[189]);
    assign layer0_outputs[10612] = ~(inputs[30]) | (inputs[187]);
    assign layer0_outputs[10613] = ~(inputs[3]);
    assign layer0_outputs[10614] = ~((inputs[182]) ^ (inputs[81]));
    assign layer0_outputs[10615] = ~(inputs[92]) | (inputs[252]);
    assign layer0_outputs[10616] = inputs[43];
    assign layer0_outputs[10617] = (inputs[174]) | (inputs[206]);
    assign layer0_outputs[10618] = inputs[76];
    assign layer0_outputs[10619] = inputs[84];
    assign layer0_outputs[10620] = (inputs[241]) & (inputs[224]);
    assign layer0_outputs[10621] = ~((inputs[206]) | (inputs[221]));
    assign layer0_outputs[10622] = (inputs[34]) | (inputs[47]);
    assign layer0_outputs[10623] = ~(inputs[108]);
    assign layer0_outputs[10624] = inputs[138];
    assign layer0_outputs[10625] = ~((inputs[214]) | (inputs[105]));
    assign layer0_outputs[10626] = (inputs[106]) | (inputs[73]);
    assign layer0_outputs[10627] = (inputs[51]) & (inputs[59]);
    assign layer0_outputs[10628] = ~((inputs[211]) | (inputs[237]));
    assign layer0_outputs[10629] = ~((inputs[68]) | (inputs[220]));
    assign layer0_outputs[10630] = ~((inputs[133]) & (inputs[162]));
    assign layer0_outputs[10631] = (inputs[188]) | (inputs[187]);
    assign layer0_outputs[10632] = ~(inputs[53]);
    assign layer0_outputs[10633] = (inputs[111]) | (inputs[41]);
    assign layer0_outputs[10634] = (inputs[102]) & ~(inputs[0]);
    assign layer0_outputs[10635] = (inputs[211]) ^ (inputs[181]);
    assign layer0_outputs[10636] = inputs[11];
    assign layer0_outputs[10637] = ~((inputs[89]) | (inputs[221]));
    assign layer0_outputs[10638] = inputs[209];
    assign layer0_outputs[10639] = 1'b1;
    assign layer0_outputs[10640] = ~(inputs[91]);
    assign layer0_outputs[10641] = ~((inputs[118]) ^ (inputs[79]));
    assign layer0_outputs[10642] = (inputs[188]) & ~(inputs[242]);
    assign layer0_outputs[10643] = inputs[166];
    assign layer0_outputs[10644] = (inputs[57]) & (inputs[4]);
    assign layer0_outputs[10645] = ~(inputs[2]) | (inputs[80]);
    assign layer0_outputs[10646] = inputs[218];
    assign layer0_outputs[10647] = ~((inputs[255]) | (inputs[102]));
    assign layer0_outputs[10648] = (inputs[25]) | (inputs[25]);
    assign layer0_outputs[10649] = inputs[38];
    assign layer0_outputs[10650] = ~(inputs[198]) | (inputs[239]);
    assign layer0_outputs[10651] = (inputs[9]) | (inputs[203]);
    assign layer0_outputs[10652] = ~((inputs[79]) ^ (inputs[28]));
    assign layer0_outputs[10653] = inputs[166];
    assign layer0_outputs[10654] = ~((inputs[164]) | (inputs[29]));
    assign layer0_outputs[10655] = ~((inputs[97]) | (inputs[82]));
    assign layer0_outputs[10656] = ~(inputs[197]) | (inputs[201]);
    assign layer0_outputs[10657] = ~(inputs[58]);
    assign layer0_outputs[10658] = (inputs[177]) | (inputs[35]);
    assign layer0_outputs[10659] = inputs[72];
    assign layer0_outputs[10660] = 1'b0;
    assign layer0_outputs[10661] = (inputs[215]) ^ (inputs[171]);
    assign layer0_outputs[10662] = (inputs[210]) ^ (inputs[104]);
    assign layer0_outputs[10663] = (inputs[139]) ^ (inputs[219]);
    assign layer0_outputs[10664] = 1'b1;
    assign layer0_outputs[10665] = (inputs[104]) & ~(inputs[225]);
    assign layer0_outputs[10666] = ~(inputs[92]);
    assign layer0_outputs[10667] = (inputs[152]) & (inputs[40]);
    assign layer0_outputs[10668] = (inputs[241]) & (inputs[189]);
    assign layer0_outputs[10669] = ~(inputs[215]) | (inputs[241]);
    assign layer0_outputs[10670] = ~(inputs[231]);
    assign layer0_outputs[10671] = ~(inputs[229]);
    assign layer0_outputs[10672] = (inputs[163]) & ~(inputs[63]);
    assign layer0_outputs[10673] = ~(inputs[197]);
    assign layer0_outputs[10674] = ~((inputs[50]) ^ (inputs[5]));
    assign layer0_outputs[10675] = ~(inputs[138]);
    assign layer0_outputs[10676] = 1'b0;
    assign layer0_outputs[10677] = ~((inputs[81]) ^ (inputs[147]));
    assign layer0_outputs[10678] = ~((inputs[171]) | (inputs[86]));
    assign layer0_outputs[10679] = (inputs[15]) & ~(inputs[143]);
    assign layer0_outputs[10680] = ~(inputs[246]);
    assign layer0_outputs[10681] = ~(inputs[104]);
    assign layer0_outputs[10682] = ~(inputs[156]) | (inputs[254]);
    assign layer0_outputs[10683] = inputs[21];
    assign layer0_outputs[10684] = (inputs[133]) | (inputs[6]);
    assign layer0_outputs[10685] = (inputs[128]) & ~(inputs[82]);
    assign layer0_outputs[10686] = ~(inputs[196]);
    assign layer0_outputs[10687] = inputs[183];
    assign layer0_outputs[10688] = ~((inputs[194]) & (inputs[119]));
    assign layer0_outputs[10689] = inputs[37];
    assign layer0_outputs[10690] = (inputs[227]) | (inputs[52]);
    assign layer0_outputs[10691] = (inputs[99]) & ~(inputs[188]);
    assign layer0_outputs[10692] = (inputs[72]) ^ (inputs[103]);
    assign layer0_outputs[10693] = (inputs[136]) ^ (inputs[252]);
    assign layer0_outputs[10694] = ~(inputs[94]);
    assign layer0_outputs[10695] = inputs[188];
    assign layer0_outputs[10696] = ~((inputs[28]) | (inputs[98]));
    assign layer0_outputs[10697] = (inputs[212]) | (inputs[73]);
    assign layer0_outputs[10698] = ~(inputs[162]);
    assign layer0_outputs[10699] = ~(inputs[82]) | (inputs[192]);
    assign layer0_outputs[10700] = ~(inputs[149]);
    assign layer0_outputs[10701] = ~((inputs[227]) | (inputs[251]));
    assign layer0_outputs[10702] = ~(inputs[56]);
    assign layer0_outputs[10703] = ~((inputs[199]) | (inputs[97]));
    assign layer0_outputs[10704] = (inputs[66]) | (inputs[35]);
    assign layer0_outputs[10705] = (inputs[85]) & ~(inputs[191]);
    assign layer0_outputs[10706] = (inputs[196]) ^ (inputs[222]);
    assign layer0_outputs[10707] = inputs[134];
    assign layer0_outputs[10708] = (inputs[64]) | (inputs[173]);
    assign layer0_outputs[10709] = (inputs[52]) & ~(inputs[130]);
    assign layer0_outputs[10710] = ~((inputs[147]) & (inputs[86]));
    assign layer0_outputs[10711] = (inputs[251]) & ~(inputs[168]);
    assign layer0_outputs[10712] = 1'b1;
    assign layer0_outputs[10713] = (inputs[26]) & ~(inputs[253]);
    assign layer0_outputs[10714] = inputs[188];
    assign layer0_outputs[10715] = ~(inputs[180]);
    assign layer0_outputs[10716] = ~((inputs[179]) | (inputs[215]));
    assign layer0_outputs[10717] = inputs[70];
    assign layer0_outputs[10718] = (inputs[162]) | (inputs[130]);
    assign layer0_outputs[10719] = 1'b0;
    assign layer0_outputs[10720] = ~(inputs[129]);
    assign layer0_outputs[10721] = ~(inputs[54]);
    assign layer0_outputs[10722] = (inputs[188]) | (inputs[152]);
    assign layer0_outputs[10723] = (inputs[58]) & (inputs[109]);
    assign layer0_outputs[10724] = (inputs[42]) | (inputs[54]);
    assign layer0_outputs[10725] = 1'b0;
    assign layer0_outputs[10726] = (inputs[156]) & ~(inputs[37]);
    assign layer0_outputs[10727] = (inputs[32]) ^ (inputs[164]);
    assign layer0_outputs[10728] = inputs[155];
    assign layer0_outputs[10729] = ~(inputs[0]);
    assign layer0_outputs[10730] = (inputs[193]) | (inputs[81]);
    assign layer0_outputs[10731] = ~(inputs[227]) | (inputs[102]);
    assign layer0_outputs[10732] = (inputs[207]) ^ (inputs[69]);
    assign layer0_outputs[10733] = ~(inputs[242]);
    assign layer0_outputs[10734] = ~(inputs[56]);
    assign layer0_outputs[10735] = (inputs[170]) & (inputs[161]);
    assign layer0_outputs[10736] = (inputs[101]) | (inputs[103]);
    assign layer0_outputs[10737] = ~((inputs[58]) ^ (inputs[242]));
    assign layer0_outputs[10738] = inputs[233];
    assign layer0_outputs[10739] = inputs[204];
    assign layer0_outputs[10740] = (inputs[148]) & ~(inputs[252]);
    assign layer0_outputs[10741] = inputs[253];
    assign layer0_outputs[10742] = ~(inputs[173]);
    assign layer0_outputs[10743] = (inputs[27]) & ~(inputs[88]);
    assign layer0_outputs[10744] = inputs[113];
    assign layer0_outputs[10745] = inputs[103];
    assign layer0_outputs[10746] = (inputs[197]) | (inputs[168]);
    assign layer0_outputs[10747] = inputs[92];
    assign layer0_outputs[10748] = ~(inputs[56]);
    assign layer0_outputs[10749] = ~((inputs[81]) ^ (inputs[74]));
    assign layer0_outputs[10750] = (inputs[124]) & ~(inputs[253]);
    assign layer0_outputs[10751] = (inputs[32]) ^ (inputs[95]);
    assign layer0_outputs[10752] = ~((inputs[84]) | (inputs[173]));
    assign layer0_outputs[10753] = ~(inputs[142]) | (inputs[88]);
    assign layer0_outputs[10754] = (inputs[42]) & ~(inputs[83]);
    assign layer0_outputs[10755] = (inputs[24]) ^ (inputs[226]);
    assign layer0_outputs[10756] = (inputs[192]) & (inputs[135]);
    assign layer0_outputs[10757] = ~((inputs[194]) | (inputs[153]));
    assign layer0_outputs[10758] = (inputs[195]) & (inputs[43]);
    assign layer0_outputs[10759] = ~(inputs[151]);
    assign layer0_outputs[10760] = ~(inputs[100]);
    assign layer0_outputs[10761] = ~(inputs[229]);
    assign layer0_outputs[10762] = ~((inputs[126]) ^ (inputs[107]));
    assign layer0_outputs[10763] = (inputs[26]) | (inputs[205]);
    assign layer0_outputs[10764] = 1'b0;
    assign layer0_outputs[10765] = ~(inputs[204]);
    assign layer0_outputs[10766] = inputs[88];
    assign layer0_outputs[10767] = (inputs[121]) & ~(inputs[243]);
    assign layer0_outputs[10768] = inputs[74];
    assign layer0_outputs[10769] = ~(inputs[187]);
    assign layer0_outputs[10770] = (inputs[182]) & (inputs[106]);
    assign layer0_outputs[10771] = 1'b1;
    assign layer0_outputs[10772] = ~(inputs[102]) | (inputs[254]);
    assign layer0_outputs[10773] = (inputs[48]) ^ (inputs[211]);
    assign layer0_outputs[10774] = (inputs[180]) & ~(inputs[165]);
    assign layer0_outputs[10775] = inputs[93];
    assign layer0_outputs[10776] = (inputs[28]) | (inputs[75]);
    assign layer0_outputs[10777] = ~(inputs[167]);
    assign layer0_outputs[10778] = inputs[149];
    assign layer0_outputs[10779] = ~(inputs[146]) | (inputs[45]);
    assign layer0_outputs[10780] = inputs[27];
    assign layer0_outputs[10781] = ~(inputs[61]) | (inputs[72]);
    assign layer0_outputs[10782] = inputs[233];
    assign layer0_outputs[10783] = ~(inputs[226]) | (inputs[47]);
    assign layer0_outputs[10784] = ~(inputs[231]);
    assign layer0_outputs[10785] = ~(inputs[72]) | (inputs[44]);
    assign layer0_outputs[10786] = ~((inputs[84]) ^ (inputs[71]));
    assign layer0_outputs[10787] = (inputs[248]) & ~(inputs[20]);
    assign layer0_outputs[10788] = ~(inputs[89]);
    assign layer0_outputs[10789] = inputs[134];
    assign layer0_outputs[10790] = ~(inputs[178]);
    assign layer0_outputs[10791] = (inputs[84]) ^ (inputs[134]);
    assign layer0_outputs[10792] = (inputs[150]) & ~(inputs[209]);
    assign layer0_outputs[10793] = ~((inputs[69]) | (inputs[113]));
    assign layer0_outputs[10794] = ~(inputs[199]) | (inputs[2]);
    assign layer0_outputs[10795] = ~(inputs[188]) | (inputs[68]);
    assign layer0_outputs[10796] = ~(inputs[45]);
    assign layer0_outputs[10797] = ~((inputs[165]) ^ (inputs[205]));
    assign layer0_outputs[10798] = inputs[178];
    assign layer0_outputs[10799] = (inputs[74]) | (inputs[19]);
    assign layer0_outputs[10800] = ~((inputs[89]) & (inputs[54]));
    assign layer0_outputs[10801] = ~(inputs[119]);
    assign layer0_outputs[10802] = (inputs[177]) & (inputs[224]);
    assign layer0_outputs[10803] = ~((inputs[1]) ^ (inputs[63]));
    assign layer0_outputs[10804] = inputs[165];
    assign layer0_outputs[10805] = ~((inputs[90]) ^ (inputs[181]));
    assign layer0_outputs[10806] = (inputs[112]) | (inputs[193]);
    assign layer0_outputs[10807] = ~((inputs[124]) | (inputs[255]));
    assign layer0_outputs[10808] = ~((inputs[234]) | (inputs[195]));
    assign layer0_outputs[10809] = (inputs[78]) & ~(inputs[142]);
    assign layer0_outputs[10810] = ~((inputs[90]) ^ (inputs[72]));
    assign layer0_outputs[10811] = inputs[138];
    assign layer0_outputs[10812] = ~((inputs[7]) | (inputs[110]));
    assign layer0_outputs[10813] = ~(inputs[2]) | (inputs[223]);
    assign layer0_outputs[10814] = ~(inputs[231]) | (inputs[69]);
    assign layer0_outputs[10815] = ~((inputs[222]) & (inputs[45]));
    assign layer0_outputs[10816] = (inputs[213]) | (inputs[210]);
    assign layer0_outputs[10817] = inputs[219];
    assign layer0_outputs[10818] = ~(inputs[208]) | (inputs[36]);
    assign layer0_outputs[10819] = (inputs[175]) | (inputs[118]);
    assign layer0_outputs[10820] = inputs[214];
    assign layer0_outputs[10821] = ~((inputs[132]) & (inputs[124]));
    assign layer0_outputs[10822] = ~((inputs[32]) ^ (inputs[154]));
    assign layer0_outputs[10823] = 1'b1;
    assign layer0_outputs[10824] = inputs[161];
    assign layer0_outputs[10825] = inputs[87];
    assign layer0_outputs[10826] = ~((inputs[227]) | (inputs[171]));
    assign layer0_outputs[10827] = ~((inputs[112]) | (inputs[113]));
    assign layer0_outputs[10828] = (inputs[198]) ^ (inputs[36]);
    assign layer0_outputs[10829] = (inputs[142]) | (inputs[1]);
    assign layer0_outputs[10830] = (inputs[248]) & ~(inputs[45]);
    assign layer0_outputs[10831] = inputs[50];
    assign layer0_outputs[10832] = inputs[183];
    assign layer0_outputs[10833] = ~(inputs[87]);
    assign layer0_outputs[10834] = (inputs[222]) | (inputs[250]);
    assign layer0_outputs[10835] = ~(inputs[150]) | (inputs[141]);
    assign layer0_outputs[10836] = inputs[205];
    assign layer0_outputs[10837] = ~(inputs[222]) | (inputs[133]);
    assign layer0_outputs[10838] = (inputs[29]) | (inputs[170]);
    assign layer0_outputs[10839] = (inputs[98]) | (inputs[80]);
    assign layer0_outputs[10840] = ~(inputs[223]);
    assign layer0_outputs[10841] = ~(inputs[176]) | (inputs[143]);
    assign layer0_outputs[10842] = ~(inputs[25]) | (inputs[193]);
    assign layer0_outputs[10843] = (inputs[54]) | (inputs[109]);
    assign layer0_outputs[10844] = (inputs[191]) | (inputs[4]);
    assign layer0_outputs[10845] = (inputs[128]) ^ (inputs[112]);
    assign layer0_outputs[10846] = ~(inputs[83]);
    assign layer0_outputs[10847] = ~(inputs[118]) | (inputs[217]);
    assign layer0_outputs[10848] = ~(inputs[78]);
    assign layer0_outputs[10849] = ~(inputs[145]) | (inputs[14]);
    assign layer0_outputs[10850] = inputs[229];
    assign layer0_outputs[10851] = ~(inputs[73]) | (inputs[226]);
    assign layer0_outputs[10852] = 1'b0;
    assign layer0_outputs[10853] = ~((inputs[34]) | (inputs[116]));
    assign layer0_outputs[10854] = (inputs[87]) & (inputs[203]);
    assign layer0_outputs[10855] = (inputs[19]) | (inputs[111]);
    assign layer0_outputs[10856] = inputs[105];
    assign layer0_outputs[10857] = (inputs[224]) & (inputs[203]);
    assign layer0_outputs[10858] = ~((inputs[24]) ^ (inputs[81]));
    assign layer0_outputs[10859] = (inputs[201]) & ~(inputs[106]);
    assign layer0_outputs[10860] = ~(inputs[91]) | (inputs[193]);
    assign layer0_outputs[10861] = inputs[234];
    assign layer0_outputs[10862] = inputs[105];
    assign layer0_outputs[10863] = (inputs[23]) & ~(inputs[72]);
    assign layer0_outputs[10864] = (inputs[185]) | (inputs[19]);
    assign layer0_outputs[10865] = 1'b0;
    assign layer0_outputs[10866] = inputs[117];
    assign layer0_outputs[10867] = ~((inputs[104]) | (inputs[119]));
    assign layer0_outputs[10868] = ~((inputs[73]) & (inputs[145]));
    assign layer0_outputs[10869] = ~((inputs[43]) ^ (inputs[197]));
    assign layer0_outputs[10870] = ~(inputs[203]);
    assign layer0_outputs[10871] = (inputs[228]) & ~(inputs[119]);
    assign layer0_outputs[10872] = (inputs[57]) & (inputs[155]);
    assign layer0_outputs[10873] = inputs[182];
    assign layer0_outputs[10874] = ~(inputs[162]);
    assign layer0_outputs[10875] = ~((inputs[14]) ^ (inputs[124]));
    assign layer0_outputs[10876] = inputs[23];
    assign layer0_outputs[10877] = ~(inputs[59]);
    assign layer0_outputs[10878] = ~(inputs[89]) | (inputs[92]);
    assign layer0_outputs[10879] = ~((inputs[105]) & (inputs[217]));
    assign layer0_outputs[10880] = ~(inputs[242]);
    assign layer0_outputs[10881] = ~(inputs[127]) | (inputs[21]);
    assign layer0_outputs[10882] = (inputs[42]) & ~(inputs[210]);
    assign layer0_outputs[10883] = ~(inputs[164]) | (inputs[48]);
    assign layer0_outputs[10884] = inputs[54];
    assign layer0_outputs[10885] = 1'b0;
    assign layer0_outputs[10886] = inputs[245];
    assign layer0_outputs[10887] = ~((inputs[212]) | (inputs[250]));
    assign layer0_outputs[10888] = inputs[23];
    assign layer0_outputs[10889] = (inputs[141]) ^ (inputs[90]);
    assign layer0_outputs[10890] = ~(inputs[152]) | (inputs[120]);
    assign layer0_outputs[10891] = (inputs[148]) & (inputs[97]);
    assign layer0_outputs[10892] = ~(inputs[116]);
    assign layer0_outputs[10893] = ~(inputs[103]) | (inputs[20]);
    assign layer0_outputs[10894] = inputs[89];
    assign layer0_outputs[10895] = 1'b1;
    assign layer0_outputs[10896] = ~(inputs[11]) | (inputs[2]);
    assign layer0_outputs[10897] = ~(inputs[235]) | (inputs[199]);
    assign layer0_outputs[10898] = ~(inputs[164]);
    assign layer0_outputs[10899] = ~(inputs[141]) | (inputs[167]);
    assign layer0_outputs[10900] = (inputs[61]) & ~(inputs[201]);
    assign layer0_outputs[10901] = (inputs[121]) | (inputs[137]);
    assign layer0_outputs[10902] = (inputs[27]) & ~(inputs[150]);
    assign layer0_outputs[10903] = (inputs[126]) & ~(inputs[50]);
    assign layer0_outputs[10904] = 1'b0;
    assign layer0_outputs[10905] = inputs[180];
    assign layer0_outputs[10906] = inputs[194];
    assign layer0_outputs[10907] = ~(inputs[139]);
    assign layer0_outputs[10908] = ~(inputs[171]) | (inputs[104]);
    assign layer0_outputs[10909] = inputs[223];
    assign layer0_outputs[10910] = inputs[48];
    assign layer0_outputs[10911] = 1'b1;
    assign layer0_outputs[10912] = (inputs[170]) ^ (inputs[135]);
    assign layer0_outputs[10913] = ~(inputs[89]) | (inputs[62]);
    assign layer0_outputs[10914] = ~((inputs[138]) | (inputs[123]));
    assign layer0_outputs[10915] = (inputs[89]) | (inputs[31]);
    assign layer0_outputs[10916] = ~(inputs[86]);
    assign layer0_outputs[10917] = (inputs[254]) | (inputs[155]);
    assign layer0_outputs[10918] = ~(inputs[240]) | (inputs[100]);
    assign layer0_outputs[10919] = ~((inputs[189]) | (inputs[192]));
    assign layer0_outputs[10920] = ~((inputs[233]) | (inputs[245]));
    assign layer0_outputs[10921] = (inputs[230]) ^ (inputs[199]);
    assign layer0_outputs[10922] = ~((inputs[138]) | (inputs[252]));
    assign layer0_outputs[10923] = (inputs[239]) | (inputs[69]);
    assign layer0_outputs[10924] = (inputs[199]) | (inputs[213]);
    assign layer0_outputs[10925] = ~((inputs[127]) | (inputs[166]));
    assign layer0_outputs[10926] = ~(inputs[236]);
    assign layer0_outputs[10927] = (inputs[104]) ^ (inputs[174]);
    assign layer0_outputs[10928] = (inputs[105]) & ~(inputs[69]);
    assign layer0_outputs[10929] = (inputs[64]) & ~(inputs[107]);
    assign layer0_outputs[10930] = inputs[81];
    assign layer0_outputs[10931] = (inputs[127]) | (inputs[46]);
    assign layer0_outputs[10932] = (inputs[32]) & ~(inputs[79]);
    assign layer0_outputs[10933] = ~(inputs[34]) | (inputs[6]);
    assign layer0_outputs[10934] = (inputs[39]) & ~(inputs[120]);
    assign layer0_outputs[10935] = (inputs[205]) ^ (inputs[126]);
    assign layer0_outputs[10936] = (inputs[208]) | (inputs[170]);
    assign layer0_outputs[10937] = ~(inputs[127]) | (inputs[223]);
    assign layer0_outputs[10938] = ~((inputs[222]) ^ (inputs[22]));
    assign layer0_outputs[10939] = inputs[125];
    assign layer0_outputs[10940] = inputs[200];
    assign layer0_outputs[10941] = 1'b1;
    assign layer0_outputs[10942] = ~(inputs[255]);
    assign layer0_outputs[10943] = (inputs[8]) ^ (inputs[144]);
    assign layer0_outputs[10944] = ~((inputs[224]) | (inputs[40]));
    assign layer0_outputs[10945] = (inputs[156]) ^ (inputs[65]);
    assign layer0_outputs[10946] = (inputs[48]) ^ (inputs[204]);
    assign layer0_outputs[10947] = ~((inputs[34]) ^ (inputs[196]));
    assign layer0_outputs[10948] = (inputs[184]) & ~(inputs[195]);
    assign layer0_outputs[10949] = ~((inputs[252]) | (inputs[160]));
    assign layer0_outputs[10950] = inputs[247];
    assign layer0_outputs[10951] = inputs[231];
    assign layer0_outputs[10952] = ~(inputs[183]) | (inputs[228]);
    assign layer0_outputs[10953] = 1'b1;
    assign layer0_outputs[10954] = ~((inputs[67]) ^ (inputs[102]));
    assign layer0_outputs[10955] = (inputs[83]) | (inputs[182]);
    assign layer0_outputs[10956] = (inputs[223]) ^ (inputs[17]);
    assign layer0_outputs[10957] = 1'b1;
    assign layer0_outputs[10958] = ~((inputs[1]) | (inputs[109]));
    assign layer0_outputs[10959] = inputs[129];
    assign layer0_outputs[10960] = ~(inputs[148]) | (inputs[89]);
    assign layer0_outputs[10961] = (inputs[162]) | (inputs[113]);
    assign layer0_outputs[10962] = ~((inputs[94]) | (inputs[117]));
    assign layer0_outputs[10963] = inputs[246];
    assign layer0_outputs[10964] = inputs[60];
    assign layer0_outputs[10965] = (inputs[68]) & ~(inputs[39]);
    assign layer0_outputs[10966] = ~(inputs[161]);
    assign layer0_outputs[10967] = ~((inputs[181]) | (inputs[75]));
    assign layer0_outputs[10968] = ~(inputs[135]) | (inputs[47]);
    assign layer0_outputs[10969] = (inputs[184]) | (inputs[178]);
    assign layer0_outputs[10970] = ~(inputs[62]) | (inputs[76]);
    assign layer0_outputs[10971] = ~((inputs[15]) | (inputs[199]));
    assign layer0_outputs[10972] = (inputs[20]) ^ (inputs[140]);
    assign layer0_outputs[10973] = ~((inputs[7]) | (inputs[224]));
    assign layer0_outputs[10974] = ~(inputs[167]) | (inputs[154]);
    assign layer0_outputs[10975] = ~(inputs[80]) | (inputs[2]);
    assign layer0_outputs[10976] = (inputs[165]) ^ (inputs[148]);
    assign layer0_outputs[10977] = inputs[137];
    assign layer0_outputs[10978] = ~(inputs[176]);
    assign layer0_outputs[10979] = ~(inputs[168]);
    assign layer0_outputs[10980] = inputs[164];
    assign layer0_outputs[10981] = (inputs[15]) | (inputs[141]);
    assign layer0_outputs[10982] = inputs[190];
    assign layer0_outputs[10983] = ~(inputs[179]);
    assign layer0_outputs[10984] = ~((inputs[157]) ^ (inputs[25]));
    assign layer0_outputs[10985] = ~((inputs[80]) | (inputs[192]));
    assign layer0_outputs[10986] = ~(inputs[56]) | (inputs[26]);
    assign layer0_outputs[10987] = ~(inputs[128]);
    assign layer0_outputs[10988] = ~(inputs[168]) | (inputs[108]);
    assign layer0_outputs[10989] = ~((inputs[233]) ^ (inputs[14]));
    assign layer0_outputs[10990] = (inputs[208]) ^ (inputs[188]);
    assign layer0_outputs[10991] = ~(inputs[254]) | (inputs[40]);
    assign layer0_outputs[10992] = inputs[37];
    assign layer0_outputs[10993] = ~((inputs[122]) ^ (inputs[153]));
    assign layer0_outputs[10994] = inputs[182];
    assign layer0_outputs[10995] = (inputs[166]) & (inputs[115]);
    assign layer0_outputs[10996] = ~(inputs[149]) | (inputs[224]);
    assign layer0_outputs[10997] = (inputs[203]) & ~(inputs[158]);
    assign layer0_outputs[10998] = inputs[26];
    assign layer0_outputs[10999] = ~(inputs[8]) | (inputs[213]);
    assign layer0_outputs[11000] = ~(inputs[43]) | (inputs[105]);
    assign layer0_outputs[11001] = (inputs[46]) & (inputs[159]);
    assign layer0_outputs[11002] = (inputs[111]) & ~(inputs[2]);
    assign layer0_outputs[11003] = (inputs[6]) ^ (inputs[53]);
    assign layer0_outputs[11004] = ~(inputs[52]);
    assign layer0_outputs[11005] = ~((inputs[134]) | (inputs[151]));
    assign layer0_outputs[11006] = ~(inputs[77]) | (inputs[255]);
    assign layer0_outputs[11007] = ~(inputs[71]);
    assign layer0_outputs[11008] = ~(inputs[17]) | (inputs[83]);
    assign layer0_outputs[11009] = ~(inputs[59]);
    assign layer0_outputs[11010] = ~(inputs[10]) | (inputs[237]);
    assign layer0_outputs[11011] = (inputs[136]) & ~(inputs[30]);
    assign layer0_outputs[11012] = ~(inputs[145]);
    assign layer0_outputs[11013] = inputs[232];
    assign layer0_outputs[11014] = ~(inputs[227]);
    assign layer0_outputs[11015] = (inputs[195]) & ~(inputs[137]);
    assign layer0_outputs[11016] = ~(inputs[129]);
    assign layer0_outputs[11017] = ~(inputs[214]);
    assign layer0_outputs[11018] = ~(inputs[232]);
    assign layer0_outputs[11019] = ~((inputs[141]) ^ (inputs[250]));
    assign layer0_outputs[11020] = inputs[74];
    assign layer0_outputs[11021] = ~((inputs[158]) | (inputs[156]));
    assign layer0_outputs[11022] = ~((inputs[66]) | (inputs[79]));
    assign layer0_outputs[11023] = (inputs[236]) ^ (inputs[181]);
    assign layer0_outputs[11024] = (inputs[12]) | (inputs[6]);
    assign layer0_outputs[11025] = ~(inputs[190]);
    assign layer0_outputs[11026] = ~(inputs[67]);
    assign layer0_outputs[11027] = ~(inputs[218]) | (inputs[110]);
    assign layer0_outputs[11028] = (inputs[45]) & ~(inputs[251]);
    assign layer0_outputs[11029] = ~((inputs[182]) & (inputs[29]));
    assign layer0_outputs[11030] = ~((inputs[163]) ^ (inputs[117]));
    assign layer0_outputs[11031] = (inputs[219]) ^ (inputs[211]);
    assign layer0_outputs[11032] = inputs[24];
    assign layer0_outputs[11033] = (inputs[104]) & ~(inputs[124]);
    assign layer0_outputs[11034] = (inputs[208]) ^ (inputs[176]);
    assign layer0_outputs[11035] = ~((inputs[47]) | (inputs[250]));
    assign layer0_outputs[11036] = 1'b1;
    assign layer0_outputs[11037] = inputs[82];
    assign layer0_outputs[11038] = ~((inputs[124]) ^ (inputs[52]));
    assign layer0_outputs[11039] = ~(inputs[151]) | (inputs[115]);
    assign layer0_outputs[11040] = ~((inputs[81]) ^ (inputs[26]));
    assign layer0_outputs[11041] = ~(inputs[44]);
    assign layer0_outputs[11042] = (inputs[151]) & ~(inputs[44]);
    assign layer0_outputs[11043] = inputs[246];
    assign layer0_outputs[11044] = (inputs[223]) | (inputs[15]);
    assign layer0_outputs[11045] = (inputs[4]) ^ (inputs[222]);
    assign layer0_outputs[11046] = inputs[87];
    assign layer0_outputs[11047] = ~(inputs[103]);
    assign layer0_outputs[11048] = ~(inputs[218]) | (inputs[58]);
    assign layer0_outputs[11049] = (inputs[85]) | (inputs[15]);
    assign layer0_outputs[11050] = (inputs[26]) & (inputs[31]);
    assign layer0_outputs[11051] = ~(inputs[104]);
    assign layer0_outputs[11052] = ~((inputs[143]) ^ (inputs[73]));
    assign layer0_outputs[11053] = ~((inputs[84]) ^ (inputs[30]));
    assign layer0_outputs[11054] = (inputs[197]) & ~(inputs[82]);
    assign layer0_outputs[11055] = (inputs[202]) ^ (inputs[218]);
    assign layer0_outputs[11056] = (inputs[98]) & (inputs[107]);
    assign layer0_outputs[11057] = ~((inputs[70]) & (inputs[117]));
    assign layer0_outputs[11058] = ~((inputs[94]) ^ (inputs[27]));
    assign layer0_outputs[11059] = (inputs[212]) | (inputs[97]);
    assign layer0_outputs[11060] = (inputs[230]) ^ (inputs[52]);
    assign layer0_outputs[11061] = ~(inputs[209]) | (inputs[100]);
    assign layer0_outputs[11062] = ~(inputs[198]) | (inputs[164]);
    assign layer0_outputs[11063] = 1'b0;
    assign layer0_outputs[11064] = inputs[18];
    assign layer0_outputs[11065] = ~(inputs[169]) | (inputs[244]);
    assign layer0_outputs[11066] = ~(inputs[90]);
    assign layer0_outputs[11067] = ~((inputs[153]) & (inputs[231]));
    assign layer0_outputs[11068] = ~(inputs[228]);
    assign layer0_outputs[11069] = (inputs[44]) | (inputs[52]);
    assign layer0_outputs[11070] = ~(inputs[136]) | (inputs[60]);
    assign layer0_outputs[11071] = ~(inputs[25]);
    assign layer0_outputs[11072] = inputs[42];
    assign layer0_outputs[11073] = (inputs[120]) & ~(inputs[129]);
    assign layer0_outputs[11074] = (inputs[63]) & ~(inputs[241]);
    assign layer0_outputs[11075] = (inputs[40]) & ~(inputs[160]);
    assign layer0_outputs[11076] = (inputs[127]) | (inputs[97]);
    assign layer0_outputs[11077] = (inputs[143]) ^ (inputs[247]);
    assign layer0_outputs[11078] = inputs[53];
    assign layer0_outputs[11079] = (inputs[164]) & ~(inputs[170]);
    assign layer0_outputs[11080] = (inputs[249]) & ~(inputs[40]);
    assign layer0_outputs[11081] = inputs[241];
    assign layer0_outputs[11082] = inputs[108];
    assign layer0_outputs[11083] = (inputs[153]) & ~(inputs[27]);
    assign layer0_outputs[11084] = ~(inputs[231]);
    assign layer0_outputs[11085] = ~(inputs[142]);
    assign layer0_outputs[11086] = ~(inputs[87]);
    assign layer0_outputs[11087] = ~(inputs[173]) | (inputs[32]);
    assign layer0_outputs[11088] = inputs[176];
    assign layer0_outputs[11089] = ~((inputs[50]) | (inputs[148]));
    assign layer0_outputs[11090] = ~(inputs[151]);
    assign layer0_outputs[11091] = (inputs[38]) & ~(inputs[241]);
    assign layer0_outputs[11092] = ~((inputs[102]) & (inputs[79]));
    assign layer0_outputs[11093] = (inputs[65]) & (inputs[10]);
    assign layer0_outputs[11094] = ~(inputs[207]);
    assign layer0_outputs[11095] = ~((inputs[163]) | (inputs[218]));
    assign layer0_outputs[11096] = ~(inputs[37]);
    assign layer0_outputs[11097] = ~(inputs[35]);
    assign layer0_outputs[11098] = ~(inputs[147]);
    assign layer0_outputs[11099] = inputs[170];
    assign layer0_outputs[11100] = ~((inputs[5]) ^ (inputs[236]));
    assign layer0_outputs[11101] = ~((inputs[171]) ^ (inputs[132]));
    assign layer0_outputs[11102] = ~(inputs[115]) | (inputs[109]);
    assign layer0_outputs[11103] = inputs[59];
    assign layer0_outputs[11104] = ~((inputs[209]) & (inputs[34]));
    assign layer0_outputs[11105] = (inputs[16]) ^ (inputs[143]);
    assign layer0_outputs[11106] = (inputs[17]) & ~(inputs[119]);
    assign layer0_outputs[11107] = ~((inputs[185]) ^ (inputs[101]));
    assign layer0_outputs[11108] = ~(inputs[100]) | (inputs[191]);
    assign layer0_outputs[11109] = inputs[198];
    assign layer0_outputs[11110] = (inputs[110]) & ~(inputs[106]);
    assign layer0_outputs[11111] = (inputs[181]) & ~(inputs[226]);
    assign layer0_outputs[11112] = inputs[151];
    assign layer0_outputs[11113] = inputs[120];
    assign layer0_outputs[11114] = ~(inputs[152]);
    assign layer0_outputs[11115] = ~(inputs[1]) | (inputs[242]);
    assign layer0_outputs[11116] = inputs[36];
    assign layer0_outputs[11117] = 1'b0;
    assign layer0_outputs[11118] = 1'b1;
    assign layer0_outputs[11119] = ~(inputs[2]) | (inputs[239]);
    assign layer0_outputs[11120] = ~((inputs[221]) & (inputs[197]));
    assign layer0_outputs[11121] = ~(inputs[88]);
    assign layer0_outputs[11122] = ~(inputs[153]);
    assign layer0_outputs[11123] = ~(inputs[35]) | (inputs[104]);
    assign layer0_outputs[11124] = (inputs[103]) & ~(inputs[34]);
    assign layer0_outputs[11125] = inputs[51];
    assign layer0_outputs[11126] = 1'b1;
    assign layer0_outputs[11127] = ~(inputs[90]);
    assign layer0_outputs[11128] = (inputs[178]) | (inputs[136]);
    assign layer0_outputs[11129] = 1'b0;
    assign layer0_outputs[11130] = ~(inputs[33]);
    assign layer0_outputs[11131] = ~((inputs[107]) ^ (inputs[177]));
    assign layer0_outputs[11132] = (inputs[96]) & ~(inputs[178]);
    assign layer0_outputs[11133] = ~(inputs[190]) | (inputs[111]);
    assign layer0_outputs[11134] = ~((inputs[111]) | (inputs[157]));
    assign layer0_outputs[11135] = ~(inputs[60]) | (inputs[210]);
    assign layer0_outputs[11136] = ~(inputs[229]);
    assign layer0_outputs[11137] = ~((inputs[221]) ^ (inputs[106]));
    assign layer0_outputs[11138] = inputs[203];
    assign layer0_outputs[11139] = ~(inputs[25]);
    assign layer0_outputs[11140] = inputs[105];
    assign layer0_outputs[11141] = inputs[0];
    assign layer0_outputs[11142] = ~((inputs[66]) | (inputs[201]));
    assign layer0_outputs[11143] = ~((inputs[135]) ^ (inputs[134]));
    assign layer0_outputs[11144] = inputs[114];
    assign layer0_outputs[11145] = ~(inputs[25]) | (inputs[181]);
    assign layer0_outputs[11146] = ~(inputs[154]) | (inputs[195]);
    assign layer0_outputs[11147] = (inputs[120]) & ~(inputs[30]);
    assign layer0_outputs[11148] = ~((inputs[135]) ^ (inputs[138]));
    assign layer0_outputs[11149] = ~((inputs[67]) | (inputs[18]));
    assign layer0_outputs[11150] = ~(inputs[183]) | (inputs[96]);
    assign layer0_outputs[11151] = ~((inputs[128]) ^ (inputs[160]));
    assign layer0_outputs[11152] = (inputs[10]) ^ (inputs[55]);
    assign layer0_outputs[11153] = (inputs[29]) & ~(inputs[193]);
    assign layer0_outputs[11154] = (inputs[51]) | (inputs[220]);
    assign layer0_outputs[11155] = ~(inputs[173]) | (inputs[207]);
    assign layer0_outputs[11156] = (inputs[83]) | (inputs[9]);
    assign layer0_outputs[11157] = (inputs[186]) & ~(inputs[18]);
    assign layer0_outputs[11158] = inputs[46];
    assign layer0_outputs[11159] = ~(inputs[118]);
    assign layer0_outputs[11160] = ~(inputs[105]) | (inputs[108]);
    assign layer0_outputs[11161] = (inputs[30]) & ~(inputs[153]);
    assign layer0_outputs[11162] = (inputs[126]) & ~(inputs[156]);
    assign layer0_outputs[11163] = ~(inputs[245]);
    assign layer0_outputs[11164] = (inputs[13]) ^ (inputs[12]);
    assign layer0_outputs[11165] = ~((inputs[111]) | (inputs[176]));
    assign layer0_outputs[11166] = ~(inputs[198]) | (inputs[113]);
    assign layer0_outputs[11167] = ~(inputs[29]);
    assign layer0_outputs[11168] = ~((inputs[148]) | (inputs[38]));
    assign layer0_outputs[11169] = ~((inputs[170]) | (inputs[138]));
    assign layer0_outputs[11170] = (inputs[85]) & ~(inputs[191]);
    assign layer0_outputs[11171] = (inputs[130]) | (inputs[195]);
    assign layer0_outputs[11172] = inputs[56];
    assign layer0_outputs[11173] = ~((inputs[132]) | (inputs[94]));
    assign layer0_outputs[11174] = inputs[149];
    assign layer0_outputs[11175] = 1'b1;
    assign layer0_outputs[11176] = (inputs[183]) | (inputs[176]);
    assign layer0_outputs[11177] = (inputs[165]) | (inputs[116]);
    assign layer0_outputs[11178] = ~((inputs[163]) ^ (inputs[242]));
    assign layer0_outputs[11179] = ~((inputs[68]) | (inputs[174]));
    assign layer0_outputs[11180] = inputs[104];
    assign layer0_outputs[11181] = ~(inputs[196]) | (inputs[55]);
    assign layer0_outputs[11182] = ~(inputs[115]) | (inputs[79]);
    assign layer0_outputs[11183] = (inputs[184]) | (inputs[255]);
    assign layer0_outputs[11184] = (inputs[88]) ^ (inputs[161]);
    assign layer0_outputs[11185] = inputs[115];
    assign layer0_outputs[11186] = ~(inputs[198]) | (inputs[1]);
    assign layer0_outputs[11187] = ~((inputs[219]) ^ (inputs[143]));
    assign layer0_outputs[11188] = (inputs[119]) ^ (inputs[212]);
    assign layer0_outputs[11189] = 1'b0;
    assign layer0_outputs[11190] = (inputs[87]) & ~(inputs[183]);
    assign layer0_outputs[11191] = ~((inputs[178]) ^ (inputs[82]));
    assign layer0_outputs[11192] = inputs[110];
    assign layer0_outputs[11193] = ~((inputs[195]) ^ (inputs[234]));
    assign layer0_outputs[11194] = ~(inputs[22]) | (inputs[147]);
    assign layer0_outputs[11195] = ~(inputs[43]) | (inputs[48]);
    assign layer0_outputs[11196] = (inputs[170]) | (inputs[201]);
    assign layer0_outputs[11197] = inputs[89];
    assign layer0_outputs[11198] = ~(inputs[27]) | (inputs[195]);
    assign layer0_outputs[11199] = ~((inputs[232]) & (inputs[235]));
    assign layer0_outputs[11200] = ~(inputs[186]);
    assign layer0_outputs[11201] = ~(inputs[118]);
    assign layer0_outputs[11202] = ~((inputs[219]) | (inputs[252]));
    assign layer0_outputs[11203] = ~(inputs[132]);
    assign layer0_outputs[11204] = 1'b0;
    assign layer0_outputs[11205] = ~(inputs[53]);
    assign layer0_outputs[11206] = inputs[199];
    assign layer0_outputs[11207] = ~((inputs[96]) | (inputs[192]));
    assign layer0_outputs[11208] = inputs[147];
    assign layer0_outputs[11209] = 1'b0;
    assign layer0_outputs[11210] = ~(inputs[181]) | (inputs[28]);
    assign layer0_outputs[11211] = ~(inputs[173]) | (inputs[41]);
    assign layer0_outputs[11212] = (inputs[230]) ^ (inputs[208]);
    assign layer0_outputs[11213] = ~((inputs[234]) & (inputs[252]));
    assign layer0_outputs[11214] = (inputs[85]) ^ (inputs[236]);
    assign layer0_outputs[11215] = inputs[173];
    assign layer0_outputs[11216] = ~((inputs[20]) | (inputs[63]));
    assign layer0_outputs[11217] = (inputs[152]) ^ (inputs[185]);
    assign layer0_outputs[11218] = inputs[221];
    assign layer0_outputs[11219] = ~(inputs[59]);
    assign layer0_outputs[11220] = inputs[139];
    assign layer0_outputs[11221] = (inputs[135]) & ~(inputs[161]);
    assign layer0_outputs[11222] = ~(inputs[151]) | (inputs[65]);
    assign layer0_outputs[11223] = ~(inputs[76]) | (inputs[0]);
    assign layer0_outputs[11224] = ~(inputs[193]);
    assign layer0_outputs[11225] = inputs[82];
    assign layer0_outputs[11226] = (inputs[245]) & (inputs[20]);
    assign layer0_outputs[11227] = ~(inputs[180]);
    assign layer0_outputs[11228] = ~(inputs[61]);
    assign layer0_outputs[11229] = inputs[150];
    assign layer0_outputs[11230] = 1'b1;
    assign layer0_outputs[11231] = ~(inputs[182]);
    assign layer0_outputs[11232] = ~(inputs[205]) | (inputs[200]);
    assign layer0_outputs[11233] = (inputs[139]) & ~(inputs[242]);
    assign layer0_outputs[11234] = ~((inputs[208]) ^ (inputs[43]));
    assign layer0_outputs[11235] = inputs[86];
    assign layer0_outputs[11236] = ~(inputs[39]) | (inputs[72]);
    assign layer0_outputs[11237] = (inputs[129]) & ~(inputs[13]);
    assign layer0_outputs[11238] = 1'b1;
    assign layer0_outputs[11239] = inputs[177];
    assign layer0_outputs[11240] = inputs[21];
    assign layer0_outputs[11241] = 1'b0;
    assign layer0_outputs[11242] = 1'b0;
    assign layer0_outputs[11243] = inputs[84];
    assign layer0_outputs[11244] = inputs[36];
    assign layer0_outputs[11245] = ~((inputs[115]) | (inputs[78]));
    assign layer0_outputs[11246] = ~((inputs[62]) | (inputs[146]));
    assign layer0_outputs[11247] = (inputs[158]) ^ (inputs[155]);
    assign layer0_outputs[11248] = (inputs[72]) & ~(inputs[110]);
    assign layer0_outputs[11249] = 1'b1;
    assign layer0_outputs[11250] = inputs[239];
    assign layer0_outputs[11251] = inputs[92];
    assign layer0_outputs[11252] = ~(inputs[97]);
    assign layer0_outputs[11253] = ~(inputs[71]) | (inputs[0]);
    assign layer0_outputs[11254] = ~(inputs[163]) | (inputs[45]);
    assign layer0_outputs[11255] = ~(inputs[79]) | (inputs[236]);
    assign layer0_outputs[11256] = (inputs[234]) & ~(inputs[128]);
    assign layer0_outputs[11257] = (inputs[100]) | (inputs[35]);
    assign layer0_outputs[11258] = (inputs[93]) | (inputs[27]);
    assign layer0_outputs[11259] = ~((inputs[236]) | (inputs[49]));
    assign layer0_outputs[11260] = inputs[185];
    assign layer0_outputs[11261] = ~(inputs[59]) | (inputs[209]);
    assign layer0_outputs[11262] = ~(inputs[216]) | (inputs[141]);
    assign layer0_outputs[11263] = (inputs[168]) & ~(inputs[88]);
    assign layer0_outputs[11264] = ~(inputs[231]) | (inputs[73]);
    assign layer0_outputs[11265] = inputs[115];
    assign layer0_outputs[11266] = ~((inputs[140]) ^ (inputs[156]));
    assign layer0_outputs[11267] = ~((inputs[134]) | (inputs[131]));
    assign layer0_outputs[11268] = ~((inputs[115]) & (inputs[0]));
    assign layer0_outputs[11269] = ~(inputs[58]);
    assign layer0_outputs[11270] = (inputs[11]) ^ (inputs[202]);
    assign layer0_outputs[11271] = (inputs[122]) & ~(inputs[54]);
    assign layer0_outputs[11272] = (inputs[172]) & ~(inputs[153]);
    assign layer0_outputs[11273] = ~(inputs[85]);
    assign layer0_outputs[11274] = (inputs[230]) | (inputs[65]);
    assign layer0_outputs[11275] = ~(inputs[255]);
    assign layer0_outputs[11276] = ~((inputs[221]) | (inputs[207]));
    assign layer0_outputs[11277] = ~((inputs[29]) | (inputs[69]));
    assign layer0_outputs[11278] = (inputs[232]) & ~(inputs[103]);
    assign layer0_outputs[11279] = (inputs[156]) & (inputs[185]);
    assign layer0_outputs[11280] = ~(inputs[48]);
    assign layer0_outputs[11281] = (inputs[204]) ^ (inputs[69]);
    assign layer0_outputs[11282] = ~((inputs[228]) & (inputs[210]));
    assign layer0_outputs[11283] = ~(inputs[87]);
    assign layer0_outputs[11284] = (inputs[218]) ^ (inputs[82]);
    assign layer0_outputs[11285] = inputs[216];
    assign layer0_outputs[11286] = ~(inputs[81]);
    assign layer0_outputs[11287] = ~(inputs[208]) | (inputs[1]);
    assign layer0_outputs[11288] = ~(inputs[111]);
    assign layer0_outputs[11289] = ~(inputs[181]);
    assign layer0_outputs[11290] = (inputs[123]) & ~(inputs[9]);
    assign layer0_outputs[11291] = ~(inputs[58]);
    assign layer0_outputs[11292] = 1'b1;
    assign layer0_outputs[11293] = (inputs[74]) & ~(inputs[251]);
    assign layer0_outputs[11294] = inputs[88];
    assign layer0_outputs[11295] = (inputs[179]) ^ (inputs[177]);
    assign layer0_outputs[11296] = inputs[25];
    assign layer0_outputs[11297] = ~(inputs[222]);
    assign layer0_outputs[11298] = ~((inputs[160]) | (inputs[140]));
    assign layer0_outputs[11299] = (inputs[219]) ^ (inputs[156]);
    assign layer0_outputs[11300] = ~(inputs[218]) | (inputs[27]);
    assign layer0_outputs[11301] = ~(inputs[158]) | (inputs[97]);
    assign layer0_outputs[11302] = (inputs[116]) & ~(inputs[221]);
    assign layer0_outputs[11303] = ~(inputs[28]) | (inputs[235]);
    assign layer0_outputs[11304] = ~((inputs[146]) | (inputs[127]));
    assign layer0_outputs[11305] = inputs[110];
    assign layer0_outputs[11306] = ~((inputs[69]) | (inputs[56]));
    assign layer0_outputs[11307] = (inputs[121]) ^ (inputs[11]);
    assign layer0_outputs[11308] = ~(inputs[134]);
    assign layer0_outputs[11309] = inputs[105];
    assign layer0_outputs[11310] = inputs[137];
    assign layer0_outputs[11311] = ~(inputs[94]) | (inputs[134]);
    assign layer0_outputs[11312] = (inputs[178]) ^ (inputs[22]);
    assign layer0_outputs[11313] = (inputs[157]) | (inputs[100]);
    assign layer0_outputs[11314] = ~(inputs[207]);
    assign layer0_outputs[11315] = (inputs[146]) | (inputs[145]);
    assign layer0_outputs[11316] = ~((inputs[248]) | (inputs[247]));
    assign layer0_outputs[11317] = inputs[120];
    assign layer0_outputs[11318] = (inputs[10]) ^ (inputs[100]);
    assign layer0_outputs[11319] = ~((inputs[65]) ^ (inputs[54]));
    assign layer0_outputs[11320] = ~(inputs[198]) | (inputs[214]);
    assign layer0_outputs[11321] = (inputs[105]) & ~(inputs[69]);
    assign layer0_outputs[11322] = ~(inputs[48]);
    assign layer0_outputs[11323] = ~(inputs[136]) | (inputs[190]);
    assign layer0_outputs[11324] = (inputs[42]) & ~(inputs[209]);
    assign layer0_outputs[11325] = (inputs[244]) & (inputs[155]);
    assign layer0_outputs[11326] = (inputs[132]) | (inputs[157]);
    assign layer0_outputs[11327] = inputs[71];
    assign layer0_outputs[11328] = inputs[182];
    assign layer0_outputs[11329] = (inputs[120]) & (inputs[188]);
    assign layer0_outputs[11330] = ~(inputs[127]) | (inputs[200]);
    assign layer0_outputs[11331] = ~((inputs[156]) & (inputs[11]));
    assign layer0_outputs[11332] = ~(inputs[158]) | (inputs[213]);
    assign layer0_outputs[11333] = (inputs[13]) ^ (inputs[90]);
    assign layer0_outputs[11334] = ~(inputs[64]);
    assign layer0_outputs[11335] = ~((inputs[107]) ^ (inputs[189]));
    assign layer0_outputs[11336] = 1'b1;
    assign layer0_outputs[11337] = (inputs[236]) | (inputs[103]);
    assign layer0_outputs[11338] = (inputs[144]) & ~(inputs[238]);
    assign layer0_outputs[11339] = (inputs[136]) | (inputs[42]);
    assign layer0_outputs[11340] = ~(inputs[155]) | (inputs[77]);
    assign layer0_outputs[11341] = (inputs[185]) ^ (inputs[142]);
    assign layer0_outputs[11342] = ~(inputs[99]);
    assign layer0_outputs[11343] = (inputs[174]) ^ (inputs[179]);
    assign layer0_outputs[11344] = ~(inputs[151]);
    assign layer0_outputs[11345] = ~((inputs[87]) ^ (inputs[101]));
    assign layer0_outputs[11346] = ~((inputs[185]) ^ (inputs[102]));
    assign layer0_outputs[11347] = ~(inputs[88]);
    assign layer0_outputs[11348] = inputs[189];
    assign layer0_outputs[11349] = (inputs[29]) & ~(inputs[0]);
    assign layer0_outputs[11350] = ~(inputs[82]);
    assign layer0_outputs[11351] = inputs[232];
    assign layer0_outputs[11352] = (inputs[233]) | (inputs[216]);
    assign layer0_outputs[11353] = 1'b0;
    assign layer0_outputs[11354] = ~((inputs[26]) ^ (inputs[57]));
    assign layer0_outputs[11355] = (inputs[222]) & ~(inputs[81]);
    assign layer0_outputs[11356] = (inputs[72]) ^ (inputs[22]);
    assign layer0_outputs[11357] = (inputs[89]) & ~(inputs[191]);
    assign layer0_outputs[11358] = inputs[50];
    assign layer0_outputs[11359] = (inputs[236]) & ~(inputs[87]);
    assign layer0_outputs[11360] = 1'b1;
    assign layer0_outputs[11361] = ~((inputs[236]) | (inputs[13]));
    assign layer0_outputs[11362] = (inputs[21]) & ~(inputs[153]);
    assign layer0_outputs[11363] = ~(inputs[247]);
    assign layer0_outputs[11364] = ~((inputs[214]) | (inputs[27]));
    assign layer0_outputs[11365] = ~((inputs[155]) | (inputs[101]));
    assign layer0_outputs[11366] = (inputs[97]) | (inputs[98]);
    assign layer0_outputs[11367] = (inputs[46]) & ~(inputs[149]);
    assign layer0_outputs[11368] = ~((inputs[81]) | (inputs[116]));
    assign layer0_outputs[11369] = inputs[178];
    assign layer0_outputs[11370] = (inputs[110]) ^ (inputs[90]);
    assign layer0_outputs[11371] = (inputs[243]) & ~(inputs[144]);
    assign layer0_outputs[11372] = inputs[214];
    assign layer0_outputs[11373] = 1'b0;
    assign layer0_outputs[11374] = (inputs[89]) & ~(inputs[67]);
    assign layer0_outputs[11375] = ~(inputs[69]);
    assign layer0_outputs[11376] = inputs[76];
    assign layer0_outputs[11377] = ~(inputs[110]);
    assign layer0_outputs[11378] = (inputs[207]) & ~(inputs[158]);
    assign layer0_outputs[11379] = inputs[18];
    assign layer0_outputs[11380] = (inputs[136]) ^ (inputs[137]);
    assign layer0_outputs[11381] = (inputs[86]) & ~(inputs[142]);
    assign layer0_outputs[11382] = inputs[130];
    assign layer0_outputs[11383] = ~(inputs[59]) | (inputs[254]);
    assign layer0_outputs[11384] = (inputs[80]) | (inputs[94]);
    assign layer0_outputs[11385] = (inputs[77]) | (inputs[139]);
    assign layer0_outputs[11386] = inputs[168];
    assign layer0_outputs[11387] = (inputs[157]) & ~(inputs[122]);
    assign layer0_outputs[11388] = (inputs[39]) | (inputs[94]);
    assign layer0_outputs[11389] = (inputs[38]) | (inputs[140]);
    assign layer0_outputs[11390] = ~((inputs[210]) | (inputs[69]));
    assign layer0_outputs[11391] = ~((inputs[43]) ^ (inputs[92]));
    assign layer0_outputs[11392] = ~(inputs[232]) | (inputs[6]);
    assign layer0_outputs[11393] = ~(inputs[138]);
    assign layer0_outputs[11394] = ~((inputs[72]) | (inputs[58]));
    assign layer0_outputs[11395] = ~(inputs[135]);
    assign layer0_outputs[11396] = ~(inputs[166]) | (inputs[223]);
    assign layer0_outputs[11397] = (inputs[133]) & (inputs[98]);
    assign layer0_outputs[11398] = (inputs[25]) | (inputs[24]);
    assign layer0_outputs[11399] = (inputs[143]) & (inputs[149]);
    assign layer0_outputs[11400] = (inputs[238]) ^ (inputs[169]);
    assign layer0_outputs[11401] = ~(inputs[15]);
    assign layer0_outputs[11402] = (inputs[29]) ^ (inputs[61]);
    assign layer0_outputs[11403] = ~(inputs[112]) | (inputs[224]);
    assign layer0_outputs[11404] = ~((inputs[119]) | (inputs[89]));
    assign layer0_outputs[11405] = (inputs[33]) & ~(inputs[255]);
    assign layer0_outputs[11406] = ~((inputs[30]) | (inputs[4]));
    assign layer0_outputs[11407] = (inputs[151]) & (inputs[197]);
    assign layer0_outputs[11408] = (inputs[181]) & ~(inputs[112]);
    assign layer0_outputs[11409] = ~((inputs[127]) ^ (inputs[110]));
    assign layer0_outputs[11410] = ~((inputs[121]) ^ (inputs[189]));
    assign layer0_outputs[11411] = (inputs[77]) & ~(inputs[253]);
    assign layer0_outputs[11412] = ~(inputs[33]);
    assign layer0_outputs[11413] = ~((inputs[109]) | (inputs[253]));
    assign layer0_outputs[11414] = ~(inputs[239]) | (inputs[14]);
    assign layer0_outputs[11415] = ~((inputs[237]) ^ (inputs[224]));
    assign layer0_outputs[11416] = 1'b0;
    assign layer0_outputs[11417] = inputs[167];
    assign layer0_outputs[11418] = ~(inputs[108]);
    assign layer0_outputs[11419] = (inputs[190]) & (inputs[153]);
    assign layer0_outputs[11420] = ~((inputs[206]) | (inputs[36]));
    assign layer0_outputs[11421] = ~(inputs[79]) | (inputs[65]);
    assign layer0_outputs[11422] = ~(inputs[79]);
    assign layer0_outputs[11423] = inputs[172];
    assign layer0_outputs[11424] = (inputs[58]) & ~(inputs[231]);
    assign layer0_outputs[11425] = ~(inputs[141]);
    assign layer0_outputs[11426] = ~(inputs[49]) | (inputs[207]);
    assign layer0_outputs[11427] = inputs[147];
    assign layer0_outputs[11428] = (inputs[177]) & ~(inputs[26]);
    assign layer0_outputs[11429] = (inputs[196]) & ~(inputs[77]);
    assign layer0_outputs[11430] = ~((inputs[222]) | (inputs[77]));
    assign layer0_outputs[11431] = ~(inputs[193]) | (inputs[157]);
    assign layer0_outputs[11432] = ~(inputs[11]);
    assign layer0_outputs[11433] = ~(inputs[64]) | (inputs[5]);
    assign layer0_outputs[11434] = (inputs[112]) & ~(inputs[65]);
    assign layer0_outputs[11435] = inputs[186];
    assign layer0_outputs[11436] = ~(inputs[238]);
    assign layer0_outputs[11437] = (inputs[31]) | (inputs[141]);
    assign layer0_outputs[11438] = (inputs[211]) ^ (inputs[226]);
    assign layer0_outputs[11439] = inputs[72];
    assign layer0_outputs[11440] = (inputs[125]) & ~(inputs[173]);
    assign layer0_outputs[11441] = (inputs[75]) ^ (inputs[159]);
    assign layer0_outputs[11442] = ~(inputs[41]);
    assign layer0_outputs[11443] = (inputs[29]) & ~(inputs[185]);
    assign layer0_outputs[11444] = ~(inputs[128]) | (inputs[64]);
    assign layer0_outputs[11445] = (inputs[147]) | (inputs[235]);
    assign layer0_outputs[11446] = (inputs[6]) & (inputs[227]);
    assign layer0_outputs[11447] = inputs[231];
    assign layer0_outputs[11448] = ~(inputs[201]);
    assign layer0_outputs[11449] = ~((inputs[134]) ^ (inputs[208]));
    assign layer0_outputs[11450] = ~(inputs[168]);
    assign layer0_outputs[11451] = (inputs[173]) & (inputs[198]);
    assign layer0_outputs[11452] = ~(inputs[184]);
    assign layer0_outputs[11453] = 1'b0;
    assign layer0_outputs[11454] = ~((inputs[176]) | (inputs[54]));
    assign layer0_outputs[11455] = (inputs[216]) | (inputs[1]);
    assign layer0_outputs[11456] = (inputs[90]) & ~(inputs[242]);
    assign layer0_outputs[11457] = inputs[97];
    assign layer0_outputs[11458] = ~((inputs[119]) ^ (inputs[73]));
    assign layer0_outputs[11459] = (inputs[227]) & ~(inputs[95]);
    assign layer0_outputs[11460] = (inputs[228]) & (inputs[84]);
    assign layer0_outputs[11461] = inputs[165];
    assign layer0_outputs[11462] = ~(inputs[254]);
    assign layer0_outputs[11463] = ~(inputs[14]);
    assign layer0_outputs[11464] = ~((inputs[216]) & (inputs[40]));
    assign layer0_outputs[11465] = inputs[227];
    assign layer0_outputs[11466] = (inputs[154]) | (inputs[29]);
    assign layer0_outputs[11467] = (inputs[212]) & ~(inputs[251]);
    assign layer0_outputs[11468] = ~(inputs[113]) | (inputs[244]);
    assign layer0_outputs[11469] = ~(inputs[166]);
    assign layer0_outputs[11470] = (inputs[111]) & ~(inputs[1]);
    assign layer0_outputs[11471] = 1'b0;
    assign layer0_outputs[11472] = ~((inputs[176]) | (inputs[249]));
    assign layer0_outputs[11473] = ~((inputs[114]) | (inputs[131]));
    assign layer0_outputs[11474] = ~(inputs[245]);
    assign layer0_outputs[11475] = ~((inputs[162]) | (inputs[114]));
    assign layer0_outputs[11476] = ~(inputs[10]);
    assign layer0_outputs[11477] = ~(inputs[220]);
    assign layer0_outputs[11478] = inputs[82];
    assign layer0_outputs[11479] = (inputs[70]) & ~(inputs[32]);
    assign layer0_outputs[11480] = (inputs[130]) | (inputs[31]);
    assign layer0_outputs[11481] = ~((inputs[153]) ^ (inputs[0]));
    assign layer0_outputs[11482] = ~(inputs[234]);
    assign layer0_outputs[11483] = (inputs[146]) ^ (inputs[192]);
    assign layer0_outputs[11484] = (inputs[227]) & ~(inputs[95]);
    assign layer0_outputs[11485] = inputs[42];
    assign layer0_outputs[11486] = ~((inputs[125]) | (inputs[93]));
    assign layer0_outputs[11487] = ~((inputs[136]) | (inputs[240]));
    assign layer0_outputs[11488] = (inputs[97]) | (inputs[4]);
    assign layer0_outputs[11489] = 1'b0;
    assign layer0_outputs[11490] = (inputs[130]) & ~(inputs[237]);
    assign layer0_outputs[11491] = (inputs[195]) & ~(inputs[44]);
    assign layer0_outputs[11492] = inputs[57];
    assign layer0_outputs[11493] = (inputs[106]) & (inputs[110]);
    assign layer0_outputs[11494] = 1'b1;
    assign layer0_outputs[11495] = ~(inputs[146]);
    assign layer0_outputs[11496] = ~((inputs[169]) | (inputs[239]));
    assign layer0_outputs[11497] = ~(inputs[122]) | (inputs[3]);
    assign layer0_outputs[11498] = inputs[139];
    assign layer0_outputs[11499] = ~(inputs[15]);
    assign layer0_outputs[11500] = (inputs[129]) | (inputs[122]);
    assign layer0_outputs[11501] = (inputs[60]) & ~(inputs[1]);
    assign layer0_outputs[11502] = ~(inputs[125]) | (inputs[64]);
    assign layer0_outputs[11503] = inputs[122];
    assign layer0_outputs[11504] = 1'b0;
    assign layer0_outputs[11505] = ~((inputs[99]) ^ (inputs[25]));
    assign layer0_outputs[11506] = ~((inputs[247]) ^ (inputs[249]));
    assign layer0_outputs[11507] = (inputs[150]) | (inputs[78]);
    assign layer0_outputs[11508] = ~(inputs[223]) | (inputs[229]);
    assign layer0_outputs[11509] = ~((inputs[51]) & (inputs[150]));
    assign layer0_outputs[11510] = ~(inputs[43]);
    assign layer0_outputs[11511] = inputs[70];
    assign layer0_outputs[11512] = (inputs[111]) | (inputs[176]);
    assign layer0_outputs[11513] = inputs[130];
    assign layer0_outputs[11514] = ~((inputs[235]) ^ (inputs[161]));
    assign layer0_outputs[11515] = ~(inputs[68]);
    assign layer0_outputs[11516] = 1'b1;
    assign layer0_outputs[11517] = (inputs[84]) & ~(inputs[172]);
    assign layer0_outputs[11518] = ~(inputs[177]) | (inputs[112]);
    assign layer0_outputs[11519] = 1'b1;
    assign layer0_outputs[11520] = ~((inputs[113]) ^ (inputs[70]));
    assign layer0_outputs[11521] = inputs[32];
    assign layer0_outputs[11522] = ~((inputs[19]) | (inputs[105]));
    assign layer0_outputs[11523] = ~(inputs[152]) | (inputs[23]);
    assign layer0_outputs[11524] = (inputs[243]) & (inputs[251]);
    assign layer0_outputs[11525] = (inputs[81]) | (inputs[175]);
    assign layer0_outputs[11526] = (inputs[39]) & ~(inputs[103]);
    assign layer0_outputs[11527] = inputs[140];
    assign layer0_outputs[11528] = ~(inputs[148]);
    assign layer0_outputs[11529] = ~(inputs[75]);
    assign layer0_outputs[11530] = ~(inputs[195]);
    assign layer0_outputs[11531] = ~((inputs[7]) | (inputs[22]));
    assign layer0_outputs[11532] = (inputs[207]) & (inputs[202]);
    assign layer0_outputs[11533] = inputs[39];
    assign layer0_outputs[11534] = ~(inputs[173]) | (inputs[185]);
    assign layer0_outputs[11535] = inputs[9];
    assign layer0_outputs[11536] = ~(inputs[23]);
    assign layer0_outputs[11537] = ~((inputs[202]) & (inputs[92]));
    assign layer0_outputs[11538] = (inputs[16]) | (inputs[166]);
    assign layer0_outputs[11539] = (inputs[160]) | (inputs[239]);
    assign layer0_outputs[11540] = ~(inputs[173]);
    assign layer0_outputs[11541] = (inputs[211]) ^ (inputs[197]);
    assign layer0_outputs[11542] = ~(inputs[199]) | (inputs[94]);
    assign layer0_outputs[11543] = 1'b1;
    assign layer0_outputs[11544] = (inputs[103]) ^ (inputs[26]);
    assign layer0_outputs[11545] = inputs[223];
    assign layer0_outputs[11546] = ~((inputs[252]) & (inputs[140]));
    assign layer0_outputs[11547] = inputs[33];
    assign layer0_outputs[11548] = ~(inputs[73]);
    assign layer0_outputs[11549] = ~((inputs[132]) & (inputs[100]));
    assign layer0_outputs[11550] = (inputs[181]) & ~(inputs[95]);
    assign layer0_outputs[11551] = ~((inputs[254]) | (inputs[119]));
    assign layer0_outputs[11552] = (inputs[220]) & ~(inputs[46]);
    assign layer0_outputs[11553] = ~(inputs[136]);
    assign layer0_outputs[11554] = (inputs[7]) ^ (inputs[31]);
    assign layer0_outputs[11555] = inputs[232];
    assign layer0_outputs[11556] = ~((inputs[168]) | (inputs[126]));
    assign layer0_outputs[11557] = ~(inputs[174]);
    assign layer0_outputs[11558] = inputs[83];
    assign layer0_outputs[11559] = inputs[61];
    assign layer0_outputs[11560] = ~((inputs[176]) ^ (inputs[25]));
    assign layer0_outputs[11561] = inputs[37];
    assign layer0_outputs[11562] = (inputs[73]) & (inputs[239]);
    assign layer0_outputs[11563] = (inputs[193]) & ~(inputs[139]);
    assign layer0_outputs[11564] = (inputs[194]) | (inputs[185]);
    assign layer0_outputs[11565] = 1'b0;
    assign layer0_outputs[11566] = 1'b0;
    assign layer0_outputs[11567] = ~((inputs[107]) | (inputs[74]));
    assign layer0_outputs[11568] = 1'b1;
    assign layer0_outputs[11569] = ~((inputs[119]) | (inputs[206]));
    assign layer0_outputs[11570] = ~((inputs[206]) | (inputs[204]));
    assign layer0_outputs[11571] = ~(inputs[53]) | (inputs[76]);
    assign layer0_outputs[11572] = ~((inputs[168]) | (inputs[225]));
    assign layer0_outputs[11573] = inputs[169];
    assign layer0_outputs[11574] = ~(inputs[78]);
    assign layer0_outputs[11575] = ~(inputs[202]) | (inputs[31]);
    assign layer0_outputs[11576] = ~(inputs[232]) | (inputs[60]);
    assign layer0_outputs[11577] = (inputs[69]) & ~(inputs[216]);
    assign layer0_outputs[11578] = ~((inputs[136]) ^ (inputs[134]));
    assign layer0_outputs[11579] = inputs[25];
    assign layer0_outputs[11580] = (inputs[21]) | (inputs[14]);
    assign layer0_outputs[11581] = inputs[138];
    assign layer0_outputs[11582] = (inputs[135]) | (inputs[150]);
    assign layer0_outputs[11583] = ~(inputs[9]);
    assign layer0_outputs[11584] = inputs[201];
    assign layer0_outputs[11585] = (inputs[86]) | (inputs[156]);
    assign layer0_outputs[11586] = ~(inputs[61]) | (inputs[38]);
    assign layer0_outputs[11587] = ~((inputs[35]) ^ (inputs[165]));
    assign layer0_outputs[11588] = (inputs[45]) & ~(inputs[51]);
    assign layer0_outputs[11589] = ~(inputs[122]);
    assign layer0_outputs[11590] = ~((inputs[179]) & (inputs[232]));
    assign layer0_outputs[11591] = ~(inputs[104]);
    assign layer0_outputs[11592] = ~(inputs[1]);
    assign layer0_outputs[11593] = (inputs[166]) ^ (inputs[148]);
    assign layer0_outputs[11594] = (inputs[206]) ^ (inputs[192]);
    assign layer0_outputs[11595] = ~((inputs[141]) ^ (inputs[206]));
    assign layer0_outputs[11596] = ~(inputs[103]);
    assign layer0_outputs[11597] = ~(inputs[51]) | (inputs[88]);
    assign layer0_outputs[11598] = inputs[113];
    assign layer0_outputs[11599] = ~(inputs[16]);
    assign layer0_outputs[11600] = (inputs[178]) ^ (inputs[16]);
    assign layer0_outputs[11601] = ~(inputs[245]);
    assign layer0_outputs[11602] = ~(inputs[153]) | (inputs[233]);
    assign layer0_outputs[11603] = ~(inputs[182]);
    assign layer0_outputs[11604] = (inputs[75]) & ~(inputs[243]);
    assign layer0_outputs[11605] = ~(inputs[126]);
    assign layer0_outputs[11606] = (inputs[30]) & ~(inputs[114]);
    assign layer0_outputs[11607] = inputs[228];
    assign layer0_outputs[11608] = ~((inputs[176]) | (inputs[47]));
    assign layer0_outputs[11609] = (inputs[130]) ^ (inputs[133]);
    assign layer0_outputs[11610] = (inputs[46]) ^ (inputs[72]);
    assign layer0_outputs[11611] = ~(inputs[157]);
    assign layer0_outputs[11612] = ~(inputs[34]) | (inputs[200]);
    assign layer0_outputs[11613] = ~(inputs[247]);
    assign layer0_outputs[11614] = (inputs[145]) ^ (inputs[32]);
    assign layer0_outputs[11615] = (inputs[212]) & ~(inputs[31]);
    assign layer0_outputs[11616] = inputs[92];
    assign layer0_outputs[11617] = (inputs[109]) ^ (inputs[52]);
    assign layer0_outputs[11618] = ~((inputs[6]) | (inputs[211]));
    assign layer0_outputs[11619] = ~(inputs[105]);
    assign layer0_outputs[11620] = (inputs[162]) | (inputs[68]);
    assign layer0_outputs[11621] = ~((inputs[134]) | (inputs[185]));
    assign layer0_outputs[11622] = ~(inputs[80]);
    assign layer0_outputs[11623] = (inputs[45]) & (inputs[87]);
    assign layer0_outputs[11624] = ~((inputs[104]) | (inputs[31]));
    assign layer0_outputs[11625] = ~((inputs[255]) | (inputs[168]));
    assign layer0_outputs[11626] = inputs[230];
    assign layer0_outputs[11627] = (inputs[212]) & ~(inputs[131]);
    assign layer0_outputs[11628] = 1'b0;
    assign layer0_outputs[11629] = inputs[88];
    assign layer0_outputs[11630] = ~((inputs[193]) | (inputs[216]));
    assign layer0_outputs[11631] = ~(inputs[39]);
    assign layer0_outputs[11632] = 1'b0;
    assign layer0_outputs[11633] = inputs[170];
    assign layer0_outputs[11634] = inputs[44];
    assign layer0_outputs[11635] = (inputs[156]) | (inputs[23]);
    assign layer0_outputs[11636] = ~(inputs[161]);
    assign layer0_outputs[11637] = (inputs[4]) & ~(inputs[239]);
    assign layer0_outputs[11638] = (inputs[235]) | (inputs[217]);
    assign layer0_outputs[11639] = ~(inputs[233]) | (inputs[209]);
    assign layer0_outputs[11640] = ~(inputs[147]);
    assign layer0_outputs[11641] = (inputs[202]) | (inputs[188]);
    assign layer0_outputs[11642] = ~(inputs[95]);
    assign layer0_outputs[11643] = (inputs[70]) & ~(inputs[71]);
    assign layer0_outputs[11644] = (inputs[217]) ^ (inputs[148]);
    assign layer0_outputs[11645] = (inputs[42]) & ~(inputs[17]);
    assign layer0_outputs[11646] = (inputs[25]) & ~(inputs[225]);
    assign layer0_outputs[11647] = ~((inputs[34]) | (inputs[184]));
    assign layer0_outputs[11648] = ~(inputs[193]) | (inputs[239]);
    assign layer0_outputs[11649] = (inputs[72]) | (inputs[211]);
    assign layer0_outputs[11650] = ~((inputs[141]) | (inputs[155]));
    assign layer0_outputs[11651] = ~((inputs[6]) | (inputs[91]));
    assign layer0_outputs[11652] = inputs[52];
    assign layer0_outputs[11653] = inputs[193];
    assign layer0_outputs[11654] = (inputs[29]) ^ (inputs[101]);
    assign layer0_outputs[11655] = ~(inputs[140]);
    assign layer0_outputs[11656] = ~(inputs[228]) | (inputs[27]);
    assign layer0_outputs[11657] = (inputs[26]) ^ (inputs[93]);
    assign layer0_outputs[11658] = ~(inputs[104]);
    assign layer0_outputs[11659] = 1'b1;
    assign layer0_outputs[11660] = ~((inputs[156]) & (inputs[121]));
    assign layer0_outputs[11661] = ~((inputs[131]) ^ (inputs[119]));
    assign layer0_outputs[11662] = ~(inputs[213]) | (inputs[56]);
    assign layer0_outputs[11663] = ~(inputs[18]);
    assign layer0_outputs[11664] = inputs[2];
    assign layer0_outputs[11665] = (inputs[38]) ^ (inputs[11]);
    assign layer0_outputs[11666] = inputs[196];
    assign layer0_outputs[11667] = (inputs[69]) ^ (inputs[100]);
    assign layer0_outputs[11668] = inputs[53];
    assign layer0_outputs[11669] = (inputs[68]) | (inputs[61]);
    assign layer0_outputs[11670] = ~(inputs[218]);
    assign layer0_outputs[11671] = ~(inputs[193]);
    assign layer0_outputs[11672] = ~(inputs[238]);
    assign layer0_outputs[11673] = (inputs[131]) & ~(inputs[32]);
    assign layer0_outputs[11674] = (inputs[6]) & ~(inputs[180]);
    assign layer0_outputs[11675] = inputs[102];
    assign layer0_outputs[11676] = (inputs[202]) | (inputs[112]);
    assign layer0_outputs[11677] = (inputs[237]) ^ (inputs[136]);
    assign layer0_outputs[11678] = ~(inputs[195]);
    assign layer0_outputs[11679] = ~(inputs[142]) | (inputs[183]);
    assign layer0_outputs[11680] = ~(inputs[41]);
    assign layer0_outputs[11681] = ~(inputs[92]);
    assign layer0_outputs[11682] = (inputs[34]) & ~(inputs[51]);
    assign layer0_outputs[11683] = (inputs[245]) | (inputs[89]);
    assign layer0_outputs[11684] = inputs[241];
    assign layer0_outputs[11685] = (inputs[192]) & ~(inputs[70]);
    assign layer0_outputs[11686] = (inputs[134]) & ~(inputs[186]);
    assign layer0_outputs[11687] = (inputs[225]) | (inputs[225]);
    assign layer0_outputs[11688] = ~(inputs[191]) | (inputs[113]);
    assign layer0_outputs[11689] = ~((inputs[88]) | (inputs[106]));
    assign layer0_outputs[11690] = 1'b0;
    assign layer0_outputs[11691] = ~(inputs[82]);
    assign layer0_outputs[11692] = (inputs[220]) | (inputs[216]);
    assign layer0_outputs[11693] = ~((inputs[246]) | (inputs[162]));
    assign layer0_outputs[11694] = ~((inputs[145]) | (inputs[55]));
    assign layer0_outputs[11695] = inputs[24];
    assign layer0_outputs[11696] = ~(inputs[232]);
    assign layer0_outputs[11697] = ~((inputs[47]) | (inputs[106]));
    assign layer0_outputs[11698] = (inputs[166]) & ~(inputs[21]);
    assign layer0_outputs[11699] = inputs[115];
    assign layer0_outputs[11700] = (inputs[209]) & ~(inputs[247]);
    assign layer0_outputs[11701] = inputs[51];
    assign layer0_outputs[11702] = 1'b1;
    assign layer0_outputs[11703] = inputs[118];
    assign layer0_outputs[11704] = inputs[66];
    assign layer0_outputs[11705] = ~(inputs[148]);
    assign layer0_outputs[11706] = (inputs[82]) | (inputs[108]);
    assign layer0_outputs[11707] = ~(inputs[167]);
    assign layer0_outputs[11708] = ~((inputs[48]) | (inputs[10]));
    assign layer0_outputs[11709] = ~(inputs[210]);
    assign layer0_outputs[11710] = (inputs[54]) & (inputs[207]);
    assign layer0_outputs[11711] = ~(inputs[233]) | (inputs[208]);
    assign layer0_outputs[11712] = inputs[105];
    assign layer0_outputs[11713] = ~(inputs[214]) | (inputs[36]);
    assign layer0_outputs[11714] = ~(inputs[228]);
    assign layer0_outputs[11715] = inputs[46];
    assign layer0_outputs[11716] = ~(inputs[97]);
    assign layer0_outputs[11717] = inputs[138];
    assign layer0_outputs[11718] = ~(inputs[246]);
    assign layer0_outputs[11719] = ~((inputs[135]) | (inputs[91]));
    assign layer0_outputs[11720] = inputs[31];
    assign layer0_outputs[11721] = inputs[129];
    assign layer0_outputs[11722] = ~(inputs[182]) | (inputs[174]);
    assign layer0_outputs[11723] = (inputs[127]) ^ (inputs[92]);
    assign layer0_outputs[11724] = inputs[86];
    assign layer0_outputs[11725] = ~((inputs[66]) ^ (inputs[156]));
    assign layer0_outputs[11726] = (inputs[195]) ^ (inputs[28]);
    assign layer0_outputs[11727] = ~(inputs[62]);
    assign layer0_outputs[11728] = inputs[63];
    assign layer0_outputs[11729] = ~(inputs[243]) | (inputs[3]);
    assign layer0_outputs[11730] = ~(inputs[6]) | (inputs[85]);
    assign layer0_outputs[11731] = (inputs[180]) & ~(inputs[142]);
    assign layer0_outputs[11732] = ~((inputs[131]) | (inputs[152]));
    assign layer0_outputs[11733] = inputs[100];
    assign layer0_outputs[11734] = ~(inputs[206]) | (inputs[142]);
    assign layer0_outputs[11735] = inputs[225];
    assign layer0_outputs[11736] = ~((inputs[182]) & (inputs[200]));
    assign layer0_outputs[11737] = ~((inputs[22]) ^ (inputs[27]));
    assign layer0_outputs[11738] = 1'b1;
    assign layer0_outputs[11739] = (inputs[99]) & ~(inputs[163]);
    assign layer0_outputs[11740] = inputs[38];
    assign layer0_outputs[11741] = ~(inputs[90]);
    assign layer0_outputs[11742] = 1'b0;
    assign layer0_outputs[11743] = (inputs[135]) & ~(inputs[187]);
    assign layer0_outputs[11744] = inputs[244];
    assign layer0_outputs[11745] = (inputs[210]) & (inputs[245]);
    assign layer0_outputs[11746] = (inputs[205]) | (inputs[18]);
    assign layer0_outputs[11747] = (inputs[192]) & ~(inputs[253]);
    assign layer0_outputs[11748] = (inputs[32]) & ~(inputs[241]);
    assign layer0_outputs[11749] = (inputs[113]) & ~(inputs[95]);
    assign layer0_outputs[11750] = ~(inputs[200]) | (inputs[244]);
    assign layer0_outputs[11751] = ~(inputs[218]);
    assign layer0_outputs[11752] = (inputs[181]) & ~(inputs[124]);
    assign layer0_outputs[11753] = ~((inputs[220]) & (inputs[218]));
    assign layer0_outputs[11754] = inputs[40];
    assign layer0_outputs[11755] = ~((inputs[203]) | (inputs[247]));
    assign layer0_outputs[11756] = inputs[27];
    assign layer0_outputs[11757] = ~(inputs[54]);
    assign layer0_outputs[11758] = ~((inputs[197]) | (inputs[113]));
    assign layer0_outputs[11759] = ~((inputs[126]) | (inputs[228]));
    assign layer0_outputs[11760] = (inputs[44]) & (inputs[39]);
    assign layer0_outputs[11761] = (inputs[54]) | (inputs[167]);
    assign layer0_outputs[11762] = (inputs[109]) | (inputs[237]);
    assign layer0_outputs[11763] = 1'b1;
    assign layer0_outputs[11764] = (inputs[84]) & ~(inputs[58]);
    assign layer0_outputs[11765] = ~(inputs[230]) | (inputs[14]);
    assign layer0_outputs[11766] = (inputs[148]) & ~(inputs[52]);
    assign layer0_outputs[11767] = 1'b1;
    assign layer0_outputs[11768] = (inputs[44]) | (inputs[22]);
    assign layer0_outputs[11769] = inputs[248];
    assign layer0_outputs[11770] = 1'b1;
    assign layer0_outputs[11771] = inputs[86];
    assign layer0_outputs[11772] = ~((inputs[163]) ^ (inputs[76]));
    assign layer0_outputs[11773] = (inputs[41]) ^ (inputs[86]);
    assign layer0_outputs[11774] = (inputs[26]) & (inputs[227]);
    assign layer0_outputs[11775] = (inputs[135]) ^ (inputs[95]);
    assign layer0_outputs[11776] = (inputs[203]) & (inputs[200]);
    assign layer0_outputs[11777] = inputs[165];
    assign layer0_outputs[11778] = inputs[231];
    assign layer0_outputs[11779] = inputs[198];
    assign layer0_outputs[11780] = ~((inputs[39]) | (inputs[64]));
    assign layer0_outputs[11781] = ~(inputs[194]);
    assign layer0_outputs[11782] = ~(inputs[29]);
    assign layer0_outputs[11783] = ~(inputs[69]);
    assign layer0_outputs[11784] = ~(inputs[77]) | (inputs[255]);
    assign layer0_outputs[11785] = ~((inputs[236]) | (inputs[176]));
    assign layer0_outputs[11786] = 1'b0;
    assign layer0_outputs[11787] = ~(inputs[26]);
    assign layer0_outputs[11788] = ~(inputs[134]);
    assign layer0_outputs[11789] = (inputs[213]) ^ (inputs[250]);
    assign layer0_outputs[11790] = inputs[203];
    assign layer0_outputs[11791] = inputs[103];
    assign layer0_outputs[11792] = (inputs[129]) ^ (inputs[92]);
    assign layer0_outputs[11793] = ~(inputs[227]) | (inputs[226]);
    assign layer0_outputs[11794] = inputs[231];
    assign layer0_outputs[11795] = ~(inputs[91]) | (inputs[192]);
    assign layer0_outputs[11796] = (inputs[30]) ^ (inputs[6]);
    assign layer0_outputs[11797] = (inputs[29]) & (inputs[200]);
    assign layer0_outputs[11798] = ~((inputs[240]) ^ (inputs[172]));
    assign layer0_outputs[11799] = inputs[113];
    assign layer0_outputs[11800] = inputs[103];
    assign layer0_outputs[11801] = 1'b0;
    assign layer0_outputs[11802] = ~(inputs[22]) | (inputs[146]);
    assign layer0_outputs[11803] = (inputs[33]) & ~(inputs[29]);
    assign layer0_outputs[11804] = (inputs[72]) ^ (inputs[239]);
    assign layer0_outputs[11805] = inputs[230];
    assign layer0_outputs[11806] = ~(inputs[96]) | (inputs[122]);
    assign layer0_outputs[11807] = ~(inputs[26]) | (inputs[205]);
    assign layer0_outputs[11808] = ~(inputs[88]);
    assign layer0_outputs[11809] = ~((inputs[97]) | (inputs[236]));
    assign layer0_outputs[11810] = ~(inputs[206]);
    assign layer0_outputs[11811] = (inputs[63]) | (inputs[176]);
    assign layer0_outputs[11812] = ~(inputs[31]);
    assign layer0_outputs[11813] = (inputs[83]) | (inputs[221]);
    assign layer0_outputs[11814] = (inputs[204]) ^ (inputs[207]);
    assign layer0_outputs[11815] = ~(inputs[62]);
    assign layer0_outputs[11816] = (inputs[54]) | (inputs[101]);
    assign layer0_outputs[11817] = (inputs[39]) & (inputs[152]);
    assign layer0_outputs[11818] = ~(inputs[219]) | (inputs[109]);
    assign layer0_outputs[11819] = (inputs[47]) ^ (inputs[203]);
    assign layer0_outputs[11820] = inputs[139];
    assign layer0_outputs[11821] = (inputs[218]) | (inputs[245]);
    assign layer0_outputs[11822] = inputs[212];
    assign layer0_outputs[11823] = inputs[83];
    assign layer0_outputs[11824] = 1'b1;
    assign layer0_outputs[11825] = ~((inputs[124]) | (inputs[19]));
    assign layer0_outputs[11826] = ~(inputs[116]);
    assign layer0_outputs[11827] = inputs[173];
    assign layer0_outputs[11828] = ~(inputs[184]);
    assign layer0_outputs[11829] = (inputs[149]) | (inputs[52]);
    assign layer0_outputs[11830] = ~(inputs[217]) | (inputs[5]);
    assign layer0_outputs[11831] = ~((inputs[173]) ^ (inputs[105]));
    assign layer0_outputs[11832] = (inputs[170]) | (inputs[171]);
    assign layer0_outputs[11833] = ~((inputs[105]) | (inputs[67]));
    assign layer0_outputs[11834] = inputs[30];
    assign layer0_outputs[11835] = inputs[216];
    assign layer0_outputs[11836] = (inputs[169]) & ~(inputs[62]);
    assign layer0_outputs[11837] = ~(inputs[183]);
    assign layer0_outputs[11838] = ~((inputs[43]) | (inputs[141]));
    assign layer0_outputs[11839] = (inputs[54]) ^ (inputs[41]);
    assign layer0_outputs[11840] = (inputs[184]) & ~(inputs[88]);
    assign layer0_outputs[11841] = 1'b0;
    assign layer0_outputs[11842] = (inputs[233]) & ~(inputs[146]);
    assign layer0_outputs[11843] = inputs[140];
    assign layer0_outputs[11844] = ~(inputs[211]) | (inputs[15]);
    assign layer0_outputs[11845] = ~(inputs[8]);
    assign layer0_outputs[11846] = (inputs[185]) & ~(inputs[252]);
    assign layer0_outputs[11847] = ~(inputs[219]);
    assign layer0_outputs[11848] = ~((inputs[16]) | (inputs[245]));
    assign layer0_outputs[11849] = ~(inputs[192]);
    assign layer0_outputs[11850] = inputs[115];
    assign layer0_outputs[11851] = ~((inputs[249]) | (inputs[105]));
    assign layer0_outputs[11852] = ~((inputs[44]) | (inputs[49]));
    assign layer0_outputs[11853] = ~(inputs[139]) | (inputs[98]);
    assign layer0_outputs[11854] = ~(inputs[223]);
    assign layer0_outputs[11855] = 1'b1;
    assign layer0_outputs[11856] = (inputs[44]) & ~(inputs[182]);
    assign layer0_outputs[11857] = ~(inputs[32]) | (inputs[10]);
    assign layer0_outputs[11858] = ~(inputs[78]);
    assign layer0_outputs[11859] = inputs[73];
    assign layer0_outputs[11860] = ~((inputs[144]) | (inputs[171]));
    assign layer0_outputs[11861] = ~(inputs[27]);
    assign layer0_outputs[11862] = (inputs[228]) & ~(inputs[58]);
    assign layer0_outputs[11863] = ~((inputs[191]) | (inputs[203]));
    assign layer0_outputs[11864] = ~(inputs[45]) | (inputs[37]);
    assign layer0_outputs[11865] = inputs[108];
    assign layer0_outputs[11866] = inputs[122];
    assign layer0_outputs[11867] = inputs[83];
    assign layer0_outputs[11868] = (inputs[25]) & ~(inputs[111]);
    assign layer0_outputs[11869] = ~((inputs[197]) | (inputs[68]));
    assign layer0_outputs[11870] = inputs[199];
    assign layer0_outputs[11871] = ~(inputs[104]);
    assign layer0_outputs[11872] = ~((inputs[64]) | (inputs[179]));
    assign layer0_outputs[11873] = ~((inputs[57]) & (inputs[117]));
    assign layer0_outputs[11874] = (inputs[9]) | (inputs[134]);
    assign layer0_outputs[11875] = inputs[83];
    assign layer0_outputs[11876] = inputs[23];
    assign layer0_outputs[11877] = (inputs[131]) & ~(inputs[224]);
    assign layer0_outputs[11878] = ~(inputs[101]);
    assign layer0_outputs[11879] = (inputs[31]) & (inputs[144]);
    assign layer0_outputs[11880] = ~(inputs[55]) | (inputs[185]);
    assign layer0_outputs[11881] = (inputs[235]) | (inputs[48]);
    assign layer0_outputs[11882] = ~(inputs[252]) | (inputs[19]);
    assign layer0_outputs[11883] = (inputs[135]) & ~(inputs[97]);
    assign layer0_outputs[11884] = 1'b0;
    assign layer0_outputs[11885] = ~(inputs[24]);
    assign layer0_outputs[11886] = ~((inputs[87]) | (inputs[102]));
    assign layer0_outputs[11887] = (inputs[63]) ^ (inputs[27]);
    assign layer0_outputs[11888] = ~(inputs[68]) | (inputs[170]);
    assign layer0_outputs[11889] = ~(inputs[110]);
    assign layer0_outputs[11890] = ~((inputs[117]) | (inputs[147]));
    assign layer0_outputs[11891] = inputs[246];
    assign layer0_outputs[11892] = (inputs[223]) ^ (inputs[193]);
    assign layer0_outputs[11893] = ~(inputs[105]) | (inputs[217]);
    assign layer0_outputs[11894] = ~(inputs[3]);
    assign layer0_outputs[11895] = (inputs[226]) & ~(inputs[238]);
    assign layer0_outputs[11896] = ~((inputs[17]) | (inputs[121]));
    assign layer0_outputs[11897] = 1'b1;
    assign layer0_outputs[11898] = inputs[17];
    assign layer0_outputs[11899] = (inputs[193]) ^ (inputs[255]);
    assign layer0_outputs[11900] = (inputs[68]) & (inputs[116]);
    assign layer0_outputs[11901] = ~(inputs[19]);
    assign layer0_outputs[11902] = 1'b1;
    assign layer0_outputs[11903] = inputs[131];
    assign layer0_outputs[11904] = (inputs[77]) & ~(inputs[154]);
    assign layer0_outputs[11905] = inputs[245];
    assign layer0_outputs[11906] = ~(inputs[36]);
    assign layer0_outputs[11907] = ~(inputs[164]);
    assign layer0_outputs[11908] = ~((inputs[86]) | (inputs[240]));
    assign layer0_outputs[11909] = inputs[242];
    assign layer0_outputs[11910] = inputs[200];
    assign layer0_outputs[11911] = ~(inputs[136]);
    assign layer0_outputs[11912] = ~((inputs[191]) ^ (inputs[1]));
    assign layer0_outputs[11913] = (inputs[161]) & ~(inputs[197]);
    assign layer0_outputs[11914] = (inputs[248]) & ~(inputs[231]);
    assign layer0_outputs[11915] = inputs[163];
    assign layer0_outputs[11916] = ~((inputs[95]) ^ (inputs[5]));
    assign layer0_outputs[11917] = (inputs[169]) | (inputs[233]);
    assign layer0_outputs[11918] = ~((inputs[175]) ^ (inputs[242]));
    assign layer0_outputs[11919] = (inputs[51]) & ~(inputs[177]);
    assign layer0_outputs[11920] = ~((inputs[246]) | (inputs[159]));
    assign layer0_outputs[11921] = ~(inputs[28]);
    assign layer0_outputs[11922] = ~(inputs[110]);
    assign layer0_outputs[11923] = inputs[214];
    assign layer0_outputs[11924] = (inputs[182]) ^ (inputs[46]);
    assign layer0_outputs[11925] = (inputs[86]) | (inputs[97]);
    assign layer0_outputs[11926] = ~(inputs[224]);
    assign layer0_outputs[11927] = ~(inputs[102]) | (inputs[159]);
    assign layer0_outputs[11928] = inputs[11];
    assign layer0_outputs[11929] = inputs[155];
    assign layer0_outputs[11930] = ~(inputs[92]) | (inputs[226]);
    assign layer0_outputs[11931] = inputs[228];
    assign layer0_outputs[11932] = ~(inputs[44]) | (inputs[198]);
    assign layer0_outputs[11933] = inputs[181];
    assign layer0_outputs[11934] = inputs[81];
    assign layer0_outputs[11935] = ~((inputs[73]) | (inputs[41]));
    assign layer0_outputs[11936] = ~(inputs[167]);
    assign layer0_outputs[11937] = ~(inputs[37]);
    assign layer0_outputs[11938] = (inputs[248]) | (inputs[213]);
    assign layer0_outputs[11939] = ~(inputs[7]) | (inputs[184]);
    assign layer0_outputs[11940] = ~(inputs[121]);
    assign layer0_outputs[11941] = inputs[216];
    assign layer0_outputs[11942] = (inputs[165]) | (inputs[222]);
    assign layer0_outputs[11943] = ~(inputs[85]);
    assign layer0_outputs[11944] = ~((inputs[138]) | (inputs[23]));
    assign layer0_outputs[11945] = inputs[180];
    assign layer0_outputs[11946] = inputs[245];
    assign layer0_outputs[11947] = ~((inputs[141]) & (inputs[54]));
    assign layer0_outputs[11948] = ~(inputs[202]);
    assign layer0_outputs[11949] = ~(inputs[128]);
    assign layer0_outputs[11950] = (inputs[199]) ^ (inputs[46]);
    assign layer0_outputs[11951] = (inputs[213]) | (inputs[167]);
    assign layer0_outputs[11952] = inputs[104];
    assign layer0_outputs[11953] = ~(inputs[145]);
    assign layer0_outputs[11954] = ~((inputs[45]) | (inputs[156]));
    assign layer0_outputs[11955] = ~(inputs[190]);
    assign layer0_outputs[11956] = ~((inputs[130]) | (inputs[155]));
    assign layer0_outputs[11957] = ~(inputs[129]);
    assign layer0_outputs[11958] = inputs[201];
    assign layer0_outputs[11959] = ~(inputs[181]);
    assign layer0_outputs[11960] = ~(inputs[74]);
    assign layer0_outputs[11961] = inputs[121];
    assign layer0_outputs[11962] = ~((inputs[116]) | (inputs[22]));
    assign layer0_outputs[11963] = 1'b0;
    assign layer0_outputs[11964] = ~((inputs[213]) | (inputs[192]));
    assign layer0_outputs[11965] = inputs[2];
    assign layer0_outputs[11966] = 1'b0;
    assign layer0_outputs[11967] = (inputs[113]) | (inputs[27]);
    assign layer0_outputs[11968] = ~((inputs[87]) ^ (inputs[99]));
    assign layer0_outputs[11969] = ~(inputs[212]) | (inputs[43]);
    assign layer0_outputs[11970] = ~(inputs[134]);
    assign layer0_outputs[11971] = (inputs[115]) & ~(inputs[192]);
    assign layer0_outputs[11972] = ~(inputs[194]);
    assign layer0_outputs[11973] = ~(inputs[58]) | (inputs[192]);
    assign layer0_outputs[11974] = (inputs[83]) & ~(inputs[144]);
    assign layer0_outputs[11975] = inputs[87];
    assign layer0_outputs[11976] = inputs[159];
    assign layer0_outputs[11977] = ~(inputs[132]);
    assign layer0_outputs[11978] = inputs[152];
    assign layer0_outputs[11979] = ~(inputs[166]) | (inputs[179]);
    assign layer0_outputs[11980] = (inputs[148]) | (inputs[182]);
    assign layer0_outputs[11981] = ~((inputs[80]) | (inputs[248]));
    assign layer0_outputs[11982] = ~((inputs[190]) | (inputs[190]));
    assign layer0_outputs[11983] = ~((inputs[2]) ^ (inputs[168]));
    assign layer0_outputs[11984] = ~(inputs[62]) | (inputs[19]);
    assign layer0_outputs[11985] = inputs[87];
    assign layer0_outputs[11986] = inputs[57];
    assign layer0_outputs[11987] = ~(inputs[108]) | (inputs[68]);
    assign layer0_outputs[11988] = ~((inputs[187]) ^ (inputs[236]));
    assign layer0_outputs[11989] = ~((inputs[58]) ^ (inputs[26]));
    assign layer0_outputs[11990] = (inputs[44]) & (inputs[50]);
    assign layer0_outputs[11991] = ~((inputs[172]) | (inputs[243]));
    assign layer0_outputs[11992] = ~((inputs[3]) | (inputs[10]));
    assign layer0_outputs[11993] = inputs[3];
    assign layer0_outputs[11994] = ~(inputs[113]);
    assign layer0_outputs[11995] = 1'b0;
    assign layer0_outputs[11996] = ~((inputs[105]) | (inputs[184]));
    assign layer0_outputs[11997] = inputs[187];
    assign layer0_outputs[11998] = ~(inputs[100]);
    assign layer0_outputs[11999] = (inputs[70]) & ~(inputs[225]);
    assign layer0_outputs[12000] = (inputs[198]) ^ (inputs[168]);
    assign layer0_outputs[12001] = (inputs[97]) & ~(inputs[51]);
    assign layer0_outputs[12002] = inputs[130];
    assign layer0_outputs[12003] = inputs[29];
    assign layer0_outputs[12004] = (inputs[193]) & ~(inputs[176]);
    assign layer0_outputs[12005] = (inputs[32]) | (inputs[42]);
    assign layer0_outputs[12006] = ~((inputs[67]) | (inputs[7]));
    assign layer0_outputs[12007] = ~((inputs[144]) | (inputs[247]));
    assign layer0_outputs[12008] = ~((inputs[94]) | (inputs[84]));
    assign layer0_outputs[12009] = inputs[54];
    assign layer0_outputs[12010] = ~(inputs[196]);
    assign layer0_outputs[12011] = ~((inputs[89]) ^ (inputs[103]));
    assign layer0_outputs[12012] = ~(inputs[84]);
    assign layer0_outputs[12013] = (inputs[85]) & ~(inputs[112]);
    assign layer0_outputs[12014] = inputs[41];
    assign layer0_outputs[12015] = ~((inputs[195]) | (inputs[62]));
    assign layer0_outputs[12016] = ~(inputs[194]);
    assign layer0_outputs[12017] = (inputs[113]) & ~(inputs[237]);
    assign layer0_outputs[12018] = ~(inputs[63]);
    assign layer0_outputs[12019] = inputs[32];
    assign layer0_outputs[12020] = ~((inputs[79]) & (inputs[168]));
    assign layer0_outputs[12021] = (inputs[5]) ^ (inputs[143]);
    assign layer0_outputs[12022] = (inputs[235]) & (inputs[13]);
    assign layer0_outputs[12023] = ~((inputs[193]) & (inputs[145]));
    assign layer0_outputs[12024] = (inputs[165]) | (inputs[70]);
    assign layer0_outputs[12025] = inputs[86];
    assign layer0_outputs[12026] = ~(inputs[55]);
    assign layer0_outputs[12027] = (inputs[159]) ^ (inputs[88]);
    assign layer0_outputs[12028] = inputs[194];
    assign layer0_outputs[12029] = ~(inputs[202]) | (inputs[0]);
    assign layer0_outputs[12030] = ~((inputs[219]) & (inputs[82]));
    assign layer0_outputs[12031] = inputs[151];
    assign layer0_outputs[12032] = inputs[152];
    assign layer0_outputs[12033] = ~(inputs[70]) | (inputs[252]);
    assign layer0_outputs[12034] = (inputs[202]) & ~(inputs[110]);
    assign layer0_outputs[12035] = inputs[237];
    assign layer0_outputs[12036] = ~(inputs[129]);
    assign layer0_outputs[12037] = (inputs[204]) | (inputs[201]);
    assign layer0_outputs[12038] = ~(inputs[133]) | (inputs[49]);
    assign layer0_outputs[12039] = (inputs[57]) ^ (inputs[45]);
    assign layer0_outputs[12040] = (inputs[132]) & ~(inputs[87]);
    assign layer0_outputs[12041] = (inputs[244]) & ~(inputs[191]);
    assign layer0_outputs[12042] = ~((inputs[100]) | (inputs[14]));
    assign layer0_outputs[12043] = (inputs[195]) ^ (inputs[152]);
    assign layer0_outputs[12044] = 1'b1;
    assign layer0_outputs[12045] = ~(inputs[59]);
    assign layer0_outputs[12046] = ~((inputs[222]) | (inputs[168]));
    assign layer0_outputs[12047] = (inputs[208]) & (inputs[50]);
    assign layer0_outputs[12048] = ~(inputs[210]) | (inputs[20]);
    assign layer0_outputs[12049] = ~(inputs[101]);
    assign layer0_outputs[12050] = inputs[92];
    assign layer0_outputs[12051] = 1'b0;
    assign layer0_outputs[12052] = (inputs[18]) & (inputs[81]);
    assign layer0_outputs[12053] = inputs[174];
    assign layer0_outputs[12054] = 1'b0;
    assign layer0_outputs[12055] = ~(inputs[121]);
    assign layer0_outputs[12056] = ~(inputs[135]);
    assign layer0_outputs[12057] = (inputs[201]) & ~(inputs[125]);
    assign layer0_outputs[12058] = (inputs[37]) & ~(inputs[95]);
    assign layer0_outputs[12059] = ~(inputs[97]) | (inputs[35]);
    assign layer0_outputs[12060] = ~((inputs[245]) | (inputs[64]));
    assign layer0_outputs[12061] = (inputs[213]) & ~(inputs[84]);
    assign layer0_outputs[12062] = ~(inputs[145]);
    assign layer0_outputs[12063] = (inputs[219]) & (inputs[238]);
    assign layer0_outputs[12064] = (inputs[101]) | (inputs[159]);
    assign layer0_outputs[12065] = ~(inputs[6]);
    assign layer0_outputs[12066] = inputs[105];
    assign layer0_outputs[12067] = ~(inputs[4]);
    assign layer0_outputs[12068] = inputs[231];
    assign layer0_outputs[12069] = 1'b0;
    assign layer0_outputs[12070] = inputs[217];
    assign layer0_outputs[12071] = ~(inputs[138]);
    assign layer0_outputs[12072] = ~(inputs[75]) | (inputs[54]);
    assign layer0_outputs[12073] = inputs[235];
    assign layer0_outputs[12074] = (inputs[97]) ^ (inputs[222]);
    assign layer0_outputs[12075] = ~(inputs[182]);
    assign layer0_outputs[12076] = (inputs[183]) & ~(inputs[93]);
    assign layer0_outputs[12077] = ~(inputs[213]);
    assign layer0_outputs[12078] = (inputs[52]) | (inputs[185]);
    assign layer0_outputs[12079] = ~(inputs[84]);
    assign layer0_outputs[12080] = ~(inputs[96]) | (inputs[119]);
    assign layer0_outputs[12081] = ~((inputs[111]) | (inputs[51]));
    assign layer0_outputs[12082] = ~(inputs[227]) | (inputs[142]);
    assign layer0_outputs[12083] = (inputs[78]) & (inputs[88]);
    assign layer0_outputs[12084] = ~(inputs[22]);
    assign layer0_outputs[12085] = inputs[78];
    assign layer0_outputs[12086] = inputs[98];
    assign layer0_outputs[12087] = (inputs[111]) ^ (inputs[222]);
    assign layer0_outputs[12088] = (inputs[71]) & (inputs[130]);
    assign layer0_outputs[12089] = ~(inputs[113]);
    assign layer0_outputs[12090] = ~((inputs[189]) ^ (inputs[214]));
    assign layer0_outputs[12091] = ~(inputs[51]) | (inputs[248]);
    assign layer0_outputs[12092] = ~(inputs[91]) | (inputs[132]);
    assign layer0_outputs[12093] = ~(inputs[149]);
    assign layer0_outputs[12094] = (inputs[206]) | (inputs[220]);
    assign layer0_outputs[12095] = ~(inputs[224]);
    assign layer0_outputs[12096] = ~((inputs[192]) ^ (inputs[147]));
    assign layer0_outputs[12097] = inputs[195];
    assign layer0_outputs[12098] = (inputs[193]) & (inputs[32]);
    assign layer0_outputs[12099] = ~(inputs[106]) | (inputs[206]);
    assign layer0_outputs[12100] = (inputs[244]) & ~(inputs[28]);
    assign layer0_outputs[12101] = ~(inputs[229]) | (inputs[105]);
    assign layer0_outputs[12102] = (inputs[180]) | (inputs[237]);
    assign layer0_outputs[12103] = (inputs[70]) & ~(inputs[194]);
    assign layer0_outputs[12104] = (inputs[57]) & ~(inputs[248]);
    assign layer0_outputs[12105] = (inputs[248]) & (inputs[10]);
    assign layer0_outputs[12106] = (inputs[86]) & ~(inputs[230]);
    assign layer0_outputs[12107] = ~((inputs[159]) ^ (inputs[11]));
    assign layer0_outputs[12108] = ~((inputs[208]) | (inputs[24]));
    assign layer0_outputs[12109] = 1'b1;
    assign layer0_outputs[12110] = ~(inputs[116]);
    assign layer0_outputs[12111] = inputs[130];
    assign layer0_outputs[12112] = ~(inputs[163]) | (inputs[67]);
    assign layer0_outputs[12113] = ~(inputs[230]) | (inputs[195]);
    assign layer0_outputs[12114] = ~((inputs[0]) | (inputs[61]));
    assign layer0_outputs[12115] = inputs[180];
    assign layer0_outputs[12116] = ~(inputs[131]);
    assign layer0_outputs[12117] = ~(inputs[108]) | (inputs[65]);
    assign layer0_outputs[12118] = ~((inputs[169]) ^ (inputs[137]));
    assign layer0_outputs[12119] = ~((inputs[100]) | (inputs[96]));
    assign layer0_outputs[12120] = (inputs[7]) & ~(inputs[118]);
    assign layer0_outputs[12121] = ~(inputs[146]);
    assign layer0_outputs[12122] = ~(inputs[122]) | (inputs[248]);
    assign layer0_outputs[12123] = ~((inputs[124]) | (inputs[249]));
    assign layer0_outputs[12124] = ~(inputs[204]) | (inputs[180]);
    assign layer0_outputs[12125] = ~(inputs[132]) | (inputs[224]);
    assign layer0_outputs[12126] = ~(inputs[179]);
    assign layer0_outputs[12127] = (inputs[99]) & ~(inputs[32]);
    assign layer0_outputs[12128] = ~(inputs[141]) | (inputs[222]);
    assign layer0_outputs[12129] = (inputs[139]) & ~(inputs[246]);
    assign layer0_outputs[12130] = ~(inputs[132]) | (inputs[104]);
    assign layer0_outputs[12131] = (inputs[46]) | (inputs[32]);
    assign layer0_outputs[12132] = ~(inputs[6]);
    assign layer0_outputs[12133] = ~(inputs[26]);
    assign layer0_outputs[12134] = (inputs[117]) ^ (inputs[234]);
    assign layer0_outputs[12135] = (inputs[252]) & (inputs[217]);
    assign layer0_outputs[12136] = (inputs[229]) | (inputs[5]);
    assign layer0_outputs[12137] = ~((inputs[187]) | (inputs[113]));
    assign layer0_outputs[12138] = (inputs[50]) | (inputs[221]);
    assign layer0_outputs[12139] = inputs[149];
    assign layer0_outputs[12140] = (inputs[140]) | (inputs[3]);
    assign layer0_outputs[12141] = inputs[85];
    assign layer0_outputs[12142] = 1'b1;
    assign layer0_outputs[12143] = ~((inputs[145]) | (inputs[108]));
    assign layer0_outputs[12144] = ~((inputs[216]) ^ (inputs[248]));
    assign layer0_outputs[12145] = ~(inputs[141]);
    assign layer0_outputs[12146] = ~(inputs[163]) | (inputs[253]);
    assign layer0_outputs[12147] = (inputs[113]) | (inputs[246]);
    assign layer0_outputs[12148] = ~((inputs[198]) ^ (inputs[242]));
    assign layer0_outputs[12149] = ~(inputs[53]) | (inputs[5]);
    assign layer0_outputs[12150] = inputs[162];
    assign layer0_outputs[12151] = (inputs[60]) & ~(inputs[119]);
    assign layer0_outputs[12152] = (inputs[156]) | (inputs[61]);
    assign layer0_outputs[12153] = ~(inputs[72]);
    assign layer0_outputs[12154] = (inputs[114]) | (inputs[78]);
    assign layer0_outputs[12155] = ~(inputs[65]);
    assign layer0_outputs[12156] = ~(inputs[49]);
    assign layer0_outputs[12157] = ~((inputs[246]) | (inputs[112]));
    assign layer0_outputs[12158] = 1'b1;
    assign layer0_outputs[12159] = ~(inputs[167]);
    assign layer0_outputs[12160] = (inputs[211]) | (inputs[205]);
    assign layer0_outputs[12161] = ~(inputs[23]);
    assign layer0_outputs[12162] = (inputs[45]) | (inputs[8]);
    assign layer0_outputs[12163] = inputs[246];
    assign layer0_outputs[12164] = (inputs[2]) & (inputs[216]);
    assign layer0_outputs[12165] = inputs[8];
    assign layer0_outputs[12166] = (inputs[227]) | (inputs[254]);
    assign layer0_outputs[12167] = ~(inputs[59]);
    assign layer0_outputs[12168] = ~(inputs[247]);
    assign layer0_outputs[12169] = ~(inputs[99]) | (inputs[18]);
    assign layer0_outputs[12170] = ~(inputs[40]);
    assign layer0_outputs[12171] = inputs[14];
    assign layer0_outputs[12172] = ~(inputs[232]);
    assign layer0_outputs[12173] = 1'b0;
    assign layer0_outputs[12174] = ~(inputs[255]);
    assign layer0_outputs[12175] = ~((inputs[173]) | (inputs[206]));
    assign layer0_outputs[12176] = (inputs[127]) | (inputs[76]);
    assign layer0_outputs[12177] = ~(inputs[203]) | (inputs[146]);
    assign layer0_outputs[12178] = (inputs[43]) & ~(inputs[251]);
    assign layer0_outputs[12179] = inputs[25];
    assign layer0_outputs[12180] = inputs[136];
    assign layer0_outputs[12181] = inputs[135];
    assign layer0_outputs[12182] = (inputs[127]) | (inputs[194]);
    assign layer0_outputs[12183] = ~(inputs[158]);
    assign layer0_outputs[12184] = ~(inputs[59]) | (inputs[19]);
    assign layer0_outputs[12185] = (inputs[51]) | (inputs[50]);
    assign layer0_outputs[12186] = (inputs[230]) & ~(inputs[43]);
    assign layer0_outputs[12187] = ~((inputs[79]) ^ (inputs[88]));
    assign layer0_outputs[12188] = ~(inputs[52]) | (inputs[145]);
    assign layer0_outputs[12189] = 1'b0;
    assign layer0_outputs[12190] = (inputs[184]) | (inputs[2]);
    assign layer0_outputs[12191] = (inputs[211]) & ~(inputs[99]);
    assign layer0_outputs[12192] = ~(inputs[169]);
    assign layer0_outputs[12193] = ~(inputs[200]);
    assign layer0_outputs[12194] = inputs[37];
    assign layer0_outputs[12195] = ~((inputs[145]) | (inputs[96]));
    assign layer0_outputs[12196] = inputs[209];
    assign layer0_outputs[12197] = ~(inputs[49]);
    assign layer0_outputs[12198] = (inputs[9]) & ~(inputs[238]);
    assign layer0_outputs[12199] = ~(inputs[76]);
    assign layer0_outputs[12200] = ~(inputs[46]);
    assign layer0_outputs[12201] = (inputs[118]) | (inputs[29]);
    assign layer0_outputs[12202] = 1'b0;
    assign layer0_outputs[12203] = ~((inputs[203]) & (inputs[115]));
    assign layer0_outputs[12204] = ~(inputs[128]);
    assign layer0_outputs[12205] = ~(inputs[118]);
    assign layer0_outputs[12206] = (inputs[192]) & ~(inputs[60]);
    assign layer0_outputs[12207] = ~(inputs[140]) | (inputs[50]);
    assign layer0_outputs[12208] = ~((inputs[78]) | (inputs[61]));
    assign layer0_outputs[12209] = inputs[81];
    assign layer0_outputs[12210] = (inputs[213]) & ~(inputs[14]);
    assign layer0_outputs[12211] = (inputs[151]) & ~(inputs[63]);
    assign layer0_outputs[12212] = (inputs[182]) | (inputs[3]);
    assign layer0_outputs[12213] = inputs[159];
    assign layer0_outputs[12214] = inputs[86];
    assign layer0_outputs[12215] = inputs[9];
    assign layer0_outputs[12216] = (inputs[102]) ^ (inputs[20]);
    assign layer0_outputs[12217] = ~(inputs[157]) | (inputs[238]);
    assign layer0_outputs[12218] = inputs[205];
    assign layer0_outputs[12219] = ~(inputs[166]) | (inputs[110]);
    assign layer0_outputs[12220] = ~((inputs[29]) & (inputs[42]));
    assign layer0_outputs[12221] = inputs[242];
    assign layer0_outputs[12222] = (inputs[90]) & ~(inputs[142]);
    assign layer0_outputs[12223] = (inputs[192]) & ~(inputs[251]);
    assign layer0_outputs[12224] = ~((inputs[252]) ^ (inputs[161]));
    assign layer0_outputs[12225] = (inputs[218]) | (inputs[205]);
    assign layer0_outputs[12226] = ~(inputs[122]);
    assign layer0_outputs[12227] = ~(inputs[7]);
    assign layer0_outputs[12228] = ~(inputs[136]);
    assign layer0_outputs[12229] = ~((inputs[242]) | (inputs[110]));
    assign layer0_outputs[12230] = ~((inputs[191]) & (inputs[57]));
    assign layer0_outputs[12231] = (inputs[188]) | (inputs[175]);
    assign layer0_outputs[12232] = ~((inputs[56]) | (inputs[223]));
    assign layer0_outputs[12233] = ~(inputs[116]);
    assign layer0_outputs[12234] = (inputs[119]) & ~(inputs[221]);
    assign layer0_outputs[12235] = (inputs[55]) | (inputs[0]);
    assign layer0_outputs[12236] = ~(inputs[47]) | (inputs[16]);
    assign layer0_outputs[12237] = ~(inputs[21]);
    assign layer0_outputs[12238] = ~(inputs[137]);
    assign layer0_outputs[12239] = ~((inputs[10]) | (inputs[153]));
    assign layer0_outputs[12240] = inputs[230];
    assign layer0_outputs[12241] = ~((inputs[16]) | (inputs[45]));
    assign layer0_outputs[12242] = (inputs[100]) & ~(inputs[143]);
    assign layer0_outputs[12243] = ~(inputs[229]);
    assign layer0_outputs[12244] = 1'b0;
    assign layer0_outputs[12245] = inputs[93];
    assign layer0_outputs[12246] = ~(inputs[229]) | (inputs[109]);
    assign layer0_outputs[12247] = ~(inputs[127]);
    assign layer0_outputs[12248] = ~(inputs[221]);
    assign layer0_outputs[12249] = inputs[166];
    assign layer0_outputs[12250] = (inputs[40]) & ~(inputs[142]);
    assign layer0_outputs[12251] = ~((inputs[41]) ^ (inputs[59]));
    assign layer0_outputs[12252] = ~(inputs[153]) | (inputs[197]);
    assign layer0_outputs[12253] = 1'b0;
    assign layer0_outputs[12254] = ~((inputs[211]) | (inputs[179]));
    assign layer0_outputs[12255] = ~(inputs[203]);
    assign layer0_outputs[12256] = (inputs[149]) ^ (inputs[114]);
    assign layer0_outputs[12257] = inputs[90];
    assign layer0_outputs[12258] = ~(inputs[170]);
    assign layer0_outputs[12259] = (inputs[172]) & ~(inputs[255]);
    assign layer0_outputs[12260] = (inputs[214]) | (inputs[67]);
    assign layer0_outputs[12261] = ~(inputs[194]) | (inputs[0]);
    assign layer0_outputs[12262] = inputs[152];
    assign layer0_outputs[12263] = (inputs[92]) & (inputs[148]);
    assign layer0_outputs[12264] = ~(inputs[138]) | (inputs[84]);
    assign layer0_outputs[12265] = ~((inputs[140]) | (inputs[206]));
    assign layer0_outputs[12266] = ~(inputs[167]);
    assign layer0_outputs[12267] = ~(inputs[57]);
    assign layer0_outputs[12268] = ~((inputs[24]) ^ (inputs[144]));
    assign layer0_outputs[12269] = inputs[134];
    assign layer0_outputs[12270] = ~((inputs[248]) ^ (inputs[235]));
    assign layer0_outputs[12271] = ~((inputs[57]) & (inputs[56]));
    assign layer0_outputs[12272] = (inputs[11]) ^ (inputs[111]);
    assign layer0_outputs[12273] = (inputs[76]) | (inputs[144]);
    assign layer0_outputs[12274] = ~((inputs[76]) ^ (inputs[3]));
    assign layer0_outputs[12275] = ~((inputs[95]) & (inputs[43]));
    assign layer0_outputs[12276] = ~((inputs[184]) | (inputs[82]));
    assign layer0_outputs[12277] = inputs[100];
    assign layer0_outputs[12278] = ~(inputs[75]);
    assign layer0_outputs[12279] = ~(inputs[70]) | (inputs[177]);
    assign layer0_outputs[12280] = ~((inputs[105]) | (inputs[104]));
    assign layer0_outputs[12281] = (inputs[153]) | (inputs[57]);
    assign layer0_outputs[12282] = ~((inputs[207]) | (inputs[25]));
    assign layer0_outputs[12283] = ~(inputs[100]);
    assign layer0_outputs[12284] = (inputs[44]) & ~(inputs[130]);
    assign layer0_outputs[12285] = ~((inputs[193]) | (inputs[207]));
    assign layer0_outputs[12286] = 1'b1;
    assign layer0_outputs[12287] = ~(inputs[78]) | (inputs[206]);
    assign layer0_outputs[12288] = 1'b1;
    assign layer0_outputs[12289] = (inputs[183]) ^ (inputs[218]);
    assign layer0_outputs[12290] = ~(inputs[14]);
    assign layer0_outputs[12291] = ~(inputs[231]);
    assign layer0_outputs[12292] = ~((inputs[148]) | (inputs[101]));
    assign layer0_outputs[12293] = (inputs[60]) | (inputs[9]);
    assign layer0_outputs[12294] = ~((inputs[66]) ^ (inputs[20]));
    assign layer0_outputs[12295] = ~(inputs[26]);
    assign layer0_outputs[12296] = (inputs[184]) ^ (inputs[216]);
    assign layer0_outputs[12297] = ~(inputs[234]);
    assign layer0_outputs[12298] = 1'b1;
    assign layer0_outputs[12299] = 1'b1;
    assign layer0_outputs[12300] = ~(inputs[122]);
    assign layer0_outputs[12301] = ~(inputs[43]) | (inputs[186]);
    assign layer0_outputs[12302] = inputs[214];
    assign layer0_outputs[12303] = ~((inputs[74]) ^ (inputs[94]));
    assign layer0_outputs[12304] = (inputs[224]) | (inputs[103]);
    assign layer0_outputs[12305] = ~(inputs[37]);
    assign layer0_outputs[12306] = inputs[218];
    assign layer0_outputs[12307] = ~((inputs[245]) | (inputs[212]));
    assign layer0_outputs[12308] = inputs[135];
    assign layer0_outputs[12309] = (inputs[210]) | (inputs[215]);
    assign layer0_outputs[12310] = ~((inputs[64]) | (inputs[233]));
    assign layer0_outputs[12311] = ~((inputs[102]) | (inputs[77]));
    assign layer0_outputs[12312] = ~(inputs[241]) | (inputs[195]);
    assign layer0_outputs[12313] = (inputs[211]) ^ (inputs[8]);
    assign layer0_outputs[12314] = (inputs[141]) | (inputs[232]);
    assign layer0_outputs[12315] = 1'b0;
    assign layer0_outputs[12316] = inputs[231];
    assign layer0_outputs[12317] = ~(inputs[194]);
    assign layer0_outputs[12318] = inputs[115];
    assign layer0_outputs[12319] = 1'b1;
    assign layer0_outputs[12320] = ~((inputs[168]) ^ (inputs[0]));
    assign layer0_outputs[12321] = (inputs[96]) & (inputs[118]);
    assign layer0_outputs[12322] = ~((inputs[216]) ^ (inputs[168]));
    assign layer0_outputs[12323] = ~(inputs[76]);
    assign layer0_outputs[12324] = (inputs[135]) & ~(inputs[178]);
    assign layer0_outputs[12325] = (inputs[211]) | (inputs[227]);
    assign layer0_outputs[12326] = inputs[94];
    assign layer0_outputs[12327] = ~(inputs[249]);
    assign layer0_outputs[12328] = (inputs[148]) | (inputs[177]);
    assign layer0_outputs[12329] = (inputs[65]) | (inputs[247]);
    assign layer0_outputs[12330] = inputs[180];
    assign layer0_outputs[12331] = ~(inputs[108]);
    assign layer0_outputs[12332] = ~((inputs[147]) | (inputs[85]));
    assign layer0_outputs[12333] = inputs[56];
    assign layer0_outputs[12334] = (inputs[155]) & (inputs[2]);
    assign layer0_outputs[12335] = ~(inputs[128]);
    assign layer0_outputs[12336] = ~((inputs[153]) & (inputs[140]));
    assign layer0_outputs[12337] = ~((inputs[202]) & (inputs[158]));
    assign layer0_outputs[12338] = ~(inputs[187]);
    assign layer0_outputs[12339] = ~(inputs[78]);
    assign layer0_outputs[12340] = ~((inputs[136]) | (inputs[66]));
    assign layer0_outputs[12341] = (inputs[35]) ^ (inputs[91]);
    assign layer0_outputs[12342] = inputs[96];
    assign layer0_outputs[12343] = (inputs[143]) | (inputs[127]);
    assign layer0_outputs[12344] = 1'b1;
    assign layer0_outputs[12345] = ~(inputs[145]);
    assign layer0_outputs[12346] = ~((inputs[94]) ^ (inputs[76]));
    assign layer0_outputs[12347] = (inputs[221]) & ~(inputs[143]);
    assign layer0_outputs[12348] = ~((inputs[190]) | (inputs[74]));
    assign layer0_outputs[12349] = ~(inputs[211]);
    assign layer0_outputs[12350] = ~((inputs[163]) | (inputs[188]));
    assign layer0_outputs[12351] = (inputs[24]) | (inputs[252]);
    assign layer0_outputs[12352] = inputs[169];
    assign layer0_outputs[12353] = ~(inputs[69]) | (inputs[214]);
    assign layer0_outputs[12354] = ~(inputs[215]);
    assign layer0_outputs[12355] = inputs[30];
    assign layer0_outputs[12356] = inputs[200];
    assign layer0_outputs[12357] = ~((inputs[201]) | (inputs[252]));
    assign layer0_outputs[12358] = ~((inputs[205]) | (inputs[188]));
    assign layer0_outputs[12359] = ~(inputs[104]);
    assign layer0_outputs[12360] = 1'b1;
    assign layer0_outputs[12361] = ~((inputs[125]) | (inputs[133]));
    assign layer0_outputs[12362] = ~((inputs[254]) | (inputs[82]));
    assign layer0_outputs[12363] = (inputs[222]) & ~(inputs[132]);
    assign layer0_outputs[12364] = ~((inputs[173]) | (inputs[106]));
    assign layer0_outputs[12365] = (inputs[70]) | (inputs[45]);
    assign layer0_outputs[12366] = ~(inputs[199]) | (inputs[14]);
    assign layer0_outputs[12367] = (inputs[48]) | (inputs[75]);
    assign layer0_outputs[12368] = ~((inputs[19]) ^ (inputs[156]));
    assign layer0_outputs[12369] = (inputs[195]) ^ (inputs[222]);
    assign layer0_outputs[12370] = ~((inputs[71]) | (inputs[28]));
    assign layer0_outputs[12371] = ~(inputs[233]);
    assign layer0_outputs[12372] = ~(inputs[100]) | (inputs[59]);
    assign layer0_outputs[12373] = (inputs[124]) & ~(inputs[62]);
    assign layer0_outputs[12374] = ~(inputs[60]);
    assign layer0_outputs[12375] = ~((inputs[97]) | (inputs[23]));
    assign layer0_outputs[12376] = ~(inputs[34]) | (inputs[17]);
    assign layer0_outputs[12377] = (inputs[15]) ^ (inputs[205]);
    assign layer0_outputs[12378] = ~(inputs[234]) | (inputs[82]);
    assign layer0_outputs[12379] = ~((inputs[111]) | (inputs[138]));
    assign layer0_outputs[12380] = inputs[24];
    assign layer0_outputs[12381] = ~(inputs[49]);
    assign layer0_outputs[12382] = ~((inputs[106]) ^ (inputs[109]));
    assign layer0_outputs[12383] = inputs[174];
    assign layer0_outputs[12384] = ~(inputs[211]);
    assign layer0_outputs[12385] = ~(inputs[57]) | (inputs[90]);
    assign layer0_outputs[12386] = ~((inputs[111]) | (inputs[182]));
    assign layer0_outputs[12387] = ~((inputs[51]) | (inputs[177]));
    assign layer0_outputs[12388] = ~(inputs[19]);
    assign layer0_outputs[12389] = ~(inputs[176]) | (inputs[212]);
    assign layer0_outputs[12390] = ~(inputs[214]);
    assign layer0_outputs[12391] = (inputs[160]) & ~(inputs[121]);
    assign layer0_outputs[12392] = (inputs[0]) & (inputs[249]);
    assign layer0_outputs[12393] = (inputs[179]) & ~(inputs[240]);
    assign layer0_outputs[12394] = (inputs[54]) & ~(inputs[205]);
    assign layer0_outputs[12395] = ~((inputs[66]) ^ (inputs[24]));
    assign layer0_outputs[12396] = (inputs[129]) | (inputs[2]);
    assign layer0_outputs[12397] = inputs[118];
    assign layer0_outputs[12398] = ~((inputs[189]) | (inputs[247]));
    assign layer0_outputs[12399] = ~(inputs[116]);
    assign layer0_outputs[12400] = (inputs[82]) ^ (inputs[163]);
    assign layer0_outputs[12401] = ~(inputs[225]);
    assign layer0_outputs[12402] = ~(inputs[69]) | (inputs[194]);
    assign layer0_outputs[12403] = (inputs[103]) & ~(inputs[48]);
    assign layer0_outputs[12404] = ~(inputs[251]);
    assign layer0_outputs[12405] = ~((inputs[23]) & (inputs[111]));
    assign layer0_outputs[12406] = inputs[70];
    assign layer0_outputs[12407] = (inputs[233]) ^ (inputs[112]);
    assign layer0_outputs[12408] = ~((inputs[184]) ^ (inputs[16]));
    assign layer0_outputs[12409] = ~(inputs[7]);
    assign layer0_outputs[12410] = (inputs[147]) | (inputs[168]);
    assign layer0_outputs[12411] = (inputs[177]) ^ (inputs[155]);
    assign layer0_outputs[12412] = ~((inputs[76]) | (inputs[95]));
    assign layer0_outputs[12413] = ~(inputs[72]);
    assign layer0_outputs[12414] = (inputs[47]) & ~(inputs[192]);
    assign layer0_outputs[12415] = ~((inputs[78]) | (inputs[35]));
    assign layer0_outputs[12416] = (inputs[232]) & ~(inputs[127]);
    assign layer0_outputs[12417] = ~((inputs[255]) ^ (inputs[227]));
    assign layer0_outputs[12418] = ~(inputs[187]) | (inputs[10]);
    assign layer0_outputs[12419] = inputs[39];
    assign layer0_outputs[12420] = ~(inputs[25]) | (inputs[155]);
    assign layer0_outputs[12421] = inputs[250];
    assign layer0_outputs[12422] = ~(inputs[133]);
    assign layer0_outputs[12423] = ~((inputs[9]) | (inputs[77]));
    assign layer0_outputs[12424] = ~((inputs[110]) | (inputs[121]));
    assign layer0_outputs[12425] = (inputs[163]) ^ (inputs[230]);
    assign layer0_outputs[12426] = ~((inputs[26]) ^ (inputs[98]));
    assign layer0_outputs[12427] = 1'b1;
    assign layer0_outputs[12428] = (inputs[69]) & ~(inputs[177]);
    assign layer0_outputs[12429] = ~((inputs[173]) & (inputs[187]));
    assign layer0_outputs[12430] = ~(inputs[167]);
    assign layer0_outputs[12431] = ~(inputs[162]);
    assign layer0_outputs[12432] = inputs[179];
    assign layer0_outputs[12433] = ~((inputs[63]) ^ (inputs[25]));
    assign layer0_outputs[12434] = (inputs[221]) & ~(inputs[142]);
    assign layer0_outputs[12435] = (inputs[210]) & (inputs[235]);
    assign layer0_outputs[12436] = inputs[25];
    assign layer0_outputs[12437] = ~((inputs[134]) & (inputs[129]));
    assign layer0_outputs[12438] = (inputs[237]) | (inputs[235]);
    assign layer0_outputs[12439] = ~((inputs[79]) ^ (inputs[29]));
    assign layer0_outputs[12440] = ~(inputs[183]) | (inputs[91]);
    assign layer0_outputs[12441] = ~(inputs[183]);
    assign layer0_outputs[12442] = ~((inputs[54]) | (inputs[204]));
    assign layer0_outputs[12443] = (inputs[4]) & ~(inputs[225]);
    assign layer0_outputs[12444] = ~((inputs[102]) ^ (inputs[54]));
    assign layer0_outputs[12445] = inputs[130];
    assign layer0_outputs[12446] = ~(inputs[163]) | (inputs[208]);
    assign layer0_outputs[12447] = ~((inputs[15]) | (inputs[159]));
    assign layer0_outputs[12448] = inputs[165];
    assign layer0_outputs[12449] = (inputs[249]) | (inputs[149]);
    assign layer0_outputs[12450] = ~((inputs[132]) ^ (inputs[191]));
    assign layer0_outputs[12451] = ~(inputs[108]) | (inputs[154]);
    assign layer0_outputs[12452] = ~(inputs[1]) | (inputs[38]);
    assign layer0_outputs[12453] = ~(inputs[107]) | (inputs[220]);
    assign layer0_outputs[12454] = ~((inputs[34]) & (inputs[205]));
    assign layer0_outputs[12455] = ~(inputs[144]);
    assign layer0_outputs[12456] = ~(inputs[52]);
    assign layer0_outputs[12457] = ~((inputs[133]) | (inputs[80]));
    assign layer0_outputs[12458] = ~((inputs[17]) & (inputs[171]));
    assign layer0_outputs[12459] = ~((inputs[88]) & (inputs[26]));
    assign layer0_outputs[12460] = ~((inputs[10]) | (inputs[52]));
    assign layer0_outputs[12461] = ~(inputs[115]);
    assign layer0_outputs[12462] = ~(inputs[234]) | (inputs[78]);
    assign layer0_outputs[12463] = ~((inputs[55]) ^ (inputs[5]));
    assign layer0_outputs[12464] = ~(inputs[177]);
    assign layer0_outputs[12465] = inputs[110];
    assign layer0_outputs[12466] = (inputs[125]) & ~(inputs[194]);
    assign layer0_outputs[12467] = ~(inputs[145]);
    assign layer0_outputs[12468] = (inputs[87]) ^ (inputs[100]);
    assign layer0_outputs[12469] = ~(inputs[68]);
    assign layer0_outputs[12470] = (inputs[179]) | (inputs[45]);
    assign layer0_outputs[12471] = (inputs[107]) | (inputs[54]);
    assign layer0_outputs[12472] = inputs[10];
    assign layer0_outputs[12473] = (inputs[165]) & (inputs[177]);
    assign layer0_outputs[12474] = ~((inputs[19]) | (inputs[62]));
    assign layer0_outputs[12475] = ~((inputs[209]) | (inputs[194]));
    assign layer0_outputs[12476] = ~((inputs[66]) ^ (inputs[234]));
    assign layer0_outputs[12477] = (inputs[253]) | (inputs[117]);
    assign layer0_outputs[12478] = ~((inputs[65]) ^ (inputs[6]));
    assign layer0_outputs[12479] = ~((inputs[105]) ^ (inputs[102]));
    assign layer0_outputs[12480] = 1'b1;
    assign layer0_outputs[12481] = (inputs[25]) & ~(inputs[208]);
    assign layer0_outputs[12482] = ~(inputs[216]);
    assign layer0_outputs[12483] = ~((inputs[127]) ^ (inputs[4]));
    assign layer0_outputs[12484] = 1'b1;
    assign layer0_outputs[12485] = ~(inputs[5]) | (inputs[175]);
    assign layer0_outputs[12486] = (inputs[90]) & ~(inputs[128]);
    assign layer0_outputs[12487] = ~((inputs[18]) ^ (inputs[118]));
    assign layer0_outputs[12488] = 1'b1;
    assign layer0_outputs[12489] = (inputs[36]) & ~(inputs[229]);
    assign layer0_outputs[12490] = ~((inputs[39]) | (inputs[111]));
    assign layer0_outputs[12491] = ~((inputs[228]) | (inputs[163]));
    assign layer0_outputs[12492] = ~(inputs[254]);
    assign layer0_outputs[12493] = (inputs[152]) ^ (inputs[149]);
    assign layer0_outputs[12494] = ~((inputs[235]) | (inputs[181]));
    assign layer0_outputs[12495] = ~(inputs[63]);
    assign layer0_outputs[12496] = ~(inputs[164]);
    assign layer0_outputs[12497] = (inputs[98]) ^ (inputs[149]);
    assign layer0_outputs[12498] = (inputs[21]) ^ (inputs[194]);
    assign layer0_outputs[12499] = inputs[79];
    assign layer0_outputs[12500] = ~(inputs[76]);
    assign layer0_outputs[12501] = ~((inputs[38]) & (inputs[81]));
    assign layer0_outputs[12502] = (inputs[122]) | (inputs[35]);
    assign layer0_outputs[12503] = (inputs[19]) | (inputs[251]);
    assign layer0_outputs[12504] = (inputs[87]) & (inputs[177]);
    assign layer0_outputs[12505] = ~(inputs[220]);
    assign layer0_outputs[12506] = (inputs[255]) & ~(inputs[149]);
    assign layer0_outputs[12507] = 1'b0;
    assign layer0_outputs[12508] = ~((inputs[194]) ^ (inputs[225]));
    assign layer0_outputs[12509] = ~((inputs[67]) | (inputs[174]));
    assign layer0_outputs[12510] = ~(inputs[92]) | (inputs[139]);
    assign layer0_outputs[12511] = inputs[255];
    assign layer0_outputs[12512] = ~(inputs[6]) | (inputs[28]);
    assign layer0_outputs[12513] = (inputs[189]) | (inputs[215]);
    assign layer0_outputs[12514] = ~((inputs[135]) | (inputs[252]));
    assign layer0_outputs[12515] = ~(inputs[167]) | (inputs[94]);
    assign layer0_outputs[12516] = (inputs[49]) & ~(inputs[36]);
    assign layer0_outputs[12517] = (inputs[150]) & (inputs[95]);
    assign layer0_outputs[12518] = inputs[195];
    assign layer0_outputs[12519] = ~((inputs[50]) ^ (inputs[141]));
    assign layer0_outputs[12520] = 1'b1;
    assign layer0_outputs[12521] = (inputs[117]) ^ (inputs[219]);
    assign layer0_outputs[12522] = inputs[211];
    assign layer0_outputs[12523] = ~((inputs[143]) ^ (inputs[75]));
    assign layer0_outputs[12524] = ~(inputs[23]) | (inputs[27]);
    assign layer0_outputs[12525] = ~(inputs[225]);
    assign layer0_outputs[12526] = 1'b0;
    assign layer0_outputs[12527] = ~(inputs[214]);
    assign layer0_outputs[12528] = (inputs[3]) | (inputs[30]);
    assign layer0_outputs[12529] = ~((inputs[196]) ^ (inputs[103]));
    assign layer0_outputs[12530] = inputs[21];
    assign layer0_outputs[12531] = inputs[121];
    assign layer0_outputs[12532] = ~((inputs[246]) | (inputs[210]));
    assign layer0_outputs[12533] = ~((inputs[28]) | (inputs[141]));
    assign layer0_outputs[12534] = 1'b1;
    assign layer0_outputs[12535] = (inputs[204]) | (inputs[235]);
    assign layer0_outputs[12536] = (inputs[129]) | (inputs[140]);
    assign layer0_outputs[12537] = 1'b1;
    assign layer0_outputs[12538] = ~((inputs[236]) | (inputs[230]));
    assign layer0_outputs[12539] = ~((inputs[29]) ^ (inputs[56]));
    assign layer0_outputs[12540] = (inputs[28]) ^ (inputs[176]);
    assign layer0_outputs[12541] = (inputs[3]) ^ (inputs[213]);
    assign layer0_outputs[12542] = inputs[36];
    assign layer0_outputs[12543] = (inputs[32]) ^ (inputs[93]);
    assign layer0_outputs[12544] = ~(inputs[88]) | (inputs[98]);
    assign layer0_outputs[12545] = inputs[227];
    assign layer0_outputs[12546] = ~(inputs[45]);
    assign layer0_outputs[12547] = (inputs[123]) & ~(inputs[149]);
    assign layer0_outputs[12548] = (inputs[236]) | (inputs[219]);
    assign layer0_outputs[12549] = (inputs[11]) & ~(inputs[51]);
    assign layer0_outputs[12550] = ~((inputs[246]) & (inputs[247]));
    assign layer0_outputs[12551] = ~(inputs[104]);
    assign layer0_outputs[12552] = inputs[28];
    assign layer0_outputs[12553] = (inputs[211]) ^ (inputs[165]);
    assign layer0_outputs[12554] = (inputs[175]) | (inputs[128]);
    assign layer0_outputs[12555] = (inputs[247]) & ~(inputs[3]);
    assign layer0_outputs[12556] = (inputs[108]) | (inputs[39]);
    assign layer0_outputs[12557] = (inputs[234]) & ~(inputs[20]);
    assign layer0_outputs[12558] = ~(inputs[68]);
    assign layer0_outputs[12559] = (inputs[206]) & ~(inputs[144]);
    assign layer0_outputs[12560] = (inputs[49]) | (inputs[41]);
    assign layer0_outputs[12561] = inputs[147];
    assign layer0_outputs[12562] = ~(inputs[67]) | (inputs[227]);
    assign layer0_outputs[12563] = (inputs[106]) & ~(inputs[13]);
    assign layer0_outputs[12564] = (inputs[110]) | (inputs[131]);
    assign layer0_outputs[12565] = (inputs[62]) ^ (inputs[71]);
    assign layer0_outputs[12566] = ~(inputs[68]);
    assign layer0_outputs[12567] = ~(inputs[93]);
    assign layer0_outputs[12568] = ~((inputs[189]) ^ (inputs[185]));
    assign layer0_outputs[12569] = (inputs[174]) & (inputs[129]);
    assign layer0_outputs[12570] = (inputs[206]) | (inputs[192]);
    assign layer0_outputs[12571] = (inputs[67]) & ~(inputs[139]);
    assign layer0_outputs[12572] = (inputs[137]) & ~(inputs[57]);
    assign layer0_outputs[12573] = ~((inputs[17]) | (inputs[237]));
    assign layer0_outputs[12574] = 1'b0;
    assign layer0_outputs[12575] = 1'b1;
    assign layer0_outputs[12576] = (inputs[198]) & (inputs[186]);
    assign layer0_outputs[12577] = ~((inputs[162]) ^ (inputs[235]));
    assign layer0_outputs[12578] = ~(inputs[44]);
    assign layer0_outputs[12579] = ~((inputs[233]) ^ (inputs[176]));
    assign layer0_outputs[12580] = inputs[114];
    assign layer0_outputs[12581] = (inputs[49]) | (inputs[85]);
    assign layer0_outputs[12582] = ~(inputs[161]) | (inputs[141]);
    assign layer0_outputs[12583] = ~(inputs[20]);
    assign layer0_outputs[12584] = ~((inputs[112]) ^ (inputs[220]));
    assign layer0_outputs[12585] = ~(inputs[84]) | (inputs[72]);
    assign layer0_outputs[12586] = ~((inputs[184]) & (inputs[210]));
    assign layer0_outputs[12587] = inputs[93];
    assign layer0_outputs[12588] = ~(inputs[219]) | (inputs[135]);
    assign layer0_outputs[12589] = (inputs[106]) & ~(inputs[179]);
    assign layer0_outputs[12590] = ~(inputs[103]) | (inputs[195]);
    assign layer0_outputs[12591] = (inputs[110]) & ~(inputs[78]);
    assign layer0_outputs[12592] = (inputs[208]) & ~(inputs[187]);
    assign layer0_outputs[12593] = ~((inputs[32]) ^ (inputs[126]));
    assign layer0_outputs[12594] = ~(inputs[73]) | (inputs[106]);
    assign layer0_outputs[12595] = inputs[88];
    assign layer0_outputs[12596] = ~((inputs[73]) ^ (inputs[78]));
    assign layer0_outputs[12597] = ~(inputs[124]);
    assign layer0_outputs[12598] = (inputs[205]) | (inputs[246]);
    assign layer0_outputs[12599] = (inputs[226]) & ~(inputs[91]);
    assign layer0_outputs[12600] = ~((inputs[166]) | (inputs[110]));
    assign layer0_outputs[12601] = ~(inputs[179]) | (inputs[61]);
    assign layer0_outputs[12602] = inputs[129];
    assign layer0_outputs[12603] = (inputs[165]) ^ (inputs[129]);
    assign layer0_outputs[12604] = ~((inputs[186]) | (inputs[252]));
    assign layer0_outputs[12605] = ~((inputs[128]) ^ (inputs[78]));
    assign layer0_outputs[12606] = ~(inputs[121]) | (inputs[65]);
    assign layer0_outputs[12607] = inputs[243];
    assign layer0_outputs[12608] = ~(inputs[176]);
    assign layer0_outputs[12609] = 1'b0;
    assign layer0_outputs[12610] = (inputs[47]) ^ (inputs[27]);
    assign layer0_outputs[12611] = inputs[32];
    assign layer0_outputs[12612] = ~((inputs[142]) ^ (inputs[108]));
    assign layer0_outputs[12613] = ~((inputs[58]) | (inputs[241]));
    assign layer0_outputs[12614] = ~(inputs[193]) | (inputs[192]);
    assign layer0_outputs[12615] = ~((inputs[184]) ^ (inputs[28]));
    assign layer0_outputs[12616] = (inputs[136]) & (inputs[139]);
    assign layer0_outputs[12617] = (inputs[49]) | (inputs[18]);
    assign layer0_outputs[12618] = (inputs[196]) | (inputs[217]);
    assign layer0_outputs[12619] = inputs[153];
    assign layer0_outputs[12620] = ~((inputs[29]) ^ (inputs[107]));
    assign layer0_outputs[12621] = inputs[183];
    assign layer0_outputs[12622] = inputs[130];
    assign layer0_outputs[12623] = inputs[141];
    assign layer0_outputs[12624] = ~(inputs[174]);
    assign layer0_outputs[12625] = ~(inputs[217]) | (inputs[121]);
    assign layer0_outputs[12626] = (inputs[81]) | (inputs[190]);
    assign layer0_outputs[12627] = inputs[21];
    assign layer0_outputs[12628] = ~(inputs[61]) | (inputs[238]);
    assign layer0_outputs[12629] = inputs[40];
    assign layer0_outputs[12630] = ~((inputs[40]) ^ (inputs[24]));
    assign layer0_outputs[12631] = (inputs[196]) | (inputs[155]);
    assign layer0_outputs[12632] = (inputs[197]) & ~(inputs[124]);
    assign layer0_outputs[12633] = (inputs[130]) & (inputs[188]);
    assign layer0_outputs[12634] = ~(inputs[33]) | (inputs[241]);
    assign layer0_outputs[12635] = ~(inputs[133]);
    assign layer0_outputs[12636] = ~(inputs[21]) | (inputs[241]);
    assign layer0_outputs[12637] = ~(inputs[215]);
    assign layer0_outputs[12638] = ~((inputs[211]) | (inputs[244]));
    assign layer0_outputs[12639] = (inputs[142]) & ~(inputs[107]);
    assign layer0_outputs[12640] = ~(inputs[161]);
    assign layer0_outputs[12641] = 1'b1;
    assign layer0_outputs[12642] = ~((inputs[91]) ^ (inputs[95]));
    assign layer0_outputs[12643] = (inputs[99]) & ~(inputs[209]);
    assign layer0_outputs[12644] = ~(inputs[15]) | (inputs[138]);
    assign layer0_outputs[12645] = (inputs[42]) & (inputs[86]);
    assign layer0_outputs[12646] = ~((inputs[0]) & (inputs[87]));
    assign layer0_outputs[12647] = (inputs[73]) | (inputs[30]);
    assign layer0_outputs[12648] = ~(inputs[146]);
    assign layer0_outputs[12649] = (inputs[247]) & ~(inputs[177]);
    assign layer0_outputs[12650] = (inputs[224]) & ~(inputs[74]);
    assign layer0_outputs[12651] = ~(inputs[99]);
    assign layer0_outputs[12652] = ~(inputs[161]);
    assign layer0_outputs[12653] = (inputs[119]) & ~(inputs[203]);
    assign layer0_outputs[12654] = ~(inputs[82]);
    assign layer0_outputs[12655] = (inputs[48]) | (inputs[217]);
    assign layer0_outputs[12656] = inputs[27];
    assign layer0_outputs[12657] = ~((inputs[161]) | (inputs[18]));
    assign layer0_outputs[12658] = ~(inputs[75]) | (inputs[206]);
    assign layer0_outputs[12659] = (inputs[47]) | (inputs[142]);
    assign layer0_outputs[12660] = inputs[76];
    assign layer0_outputs[12661] = ~(inputs[116]);
    assign layer0_outputs[12662] = inputs[147];
    assign layer0_outputs[12663] = inputs[125];
    assign layer0_outputs[12664] = inputs[128];
    assign layer0_outputs[12665] = ~(inputs[179]);
    assign layer0_outputs[12666] = inputs[244];
    assign layer0_outputs[12667] = ~(inputs[115]);
    assign layer0_outputs[12668] = ~(inputs[3]) | (inputs[20]);
    assign layer0_outputs[12669] = (inputs[61]) | (inputs[127]);
    assign layer0_outputs[12670] = ~(inputs[120]);
    assign layer0_outputs[12671] = ~((inputs[52]) ^ (inputs[118]));
    assign layer0_outputs[12672] = ~((inputs[84]) ^ (inputs[122]));
    assign layer0_outputs[12673] = ~((inputs[140]) ^ (inputs[204]));
    assign layer0_outputs[12674] = (inputs[137]) & ~(inputs[174]);
    assign layer0_outputs[12675] = ~(inputs[250]);
    assign layer0_outputs[12676] = ~((inputs[73]) | (inputs[199]));
    assign layer0_outputs[12677] = ~(inputs[152]) | (inputs[110]);
    assign layer0_outputs[12678] = ~((inputs[152]) ^ (inputs[250]));
    assign layer0_outputs[12679] = ~(inputs[89]);
    assign layer0_outputs[12680] = ~(inputs[3]) | (inputs[76]);
    assign layer0_outputs[12681] = inputs[84];
    assign layer0_outputs[12682] = ~(inputs[85]) | (inputs[173]);
    assign layer0_outputs[12683] = ~((inputs[191]) | (inputs[244]));
    assign layer0_outputs[12684] = inputs[251];
    assign layer0_outputs[12685] = (inputs[102]) | (inputs[191]);
    assign layer0_outputs[12686] = inputs[149];
    assign layer0_outputs[12687] = ~((inputs[54]) & (inputs[67]));
    assign layer0_outputs[12688] = ~((inputs[34]) ^ (inputs[136]));
    assign layer0_outputs[12689] = ~(inputs[133]);
    assign layer0_outputs[12690] = ~((inputs[68]) | (inputs[227]));
    assign layer0_outputs[12691] = inputs[120];
    assign layer0_outputs[12692] = ~(inputs[74]);
    assign layer0_outputs[12693] = ~((inputs[240]) & (inputs[14]));
    assign layer0_outputs[12694] = 1'b0;
    assign layer0_outputs[12695] = (inputs[252]) & (inputs[145]);
    assign layer0_outputs[12696] = 1'b1;
    assign layer0_outputs[12697] = ~((inputs[179]) | (inputs[75]));
    assign layer0_outputs[12698] = ~(inputs[74]);
    assign layer0_outputs[12699] = (inputs[194]) ^ (inputs[192]);
    assign layer0_outputs[12700] = ~((inputs[76]) ^ (inputs[247]));
    assign layer0_outputs[12701] = inputs[77];
    assign layer0_outputs[12702] = ~(inputs[56]);
    assign layer0_outputs[12703] = inputs[228];
    assign layer0_outputs[12704] = (inputs[0]) | (inputs[138]);
    assign layer0_outputs[12705] = ~(inputs[120]) | (inputs[69]);
    assign layer0_outputs[12706] = inputs[154];
    assign layer0_outputs[12707] = (inputs[30]) | (inputs[134]);
    assign layer0_outputs[12708] = (inputs[95]) | (inputs[59]);
    assign layer0_outputs[12709] = ~((inputs[241]) & (inputs[221]));
    assign layer0_outputs[12710] = 1'b1;
    assign layer0_outputs[12711] = inputs[163];
    assign layer0_outputs[12712] = ~((inputs[210]) ^ (inputs[206]));
    assign layer0_outputs[12713] = (inputs[231]) & ~(inputs[82]);
    assign layer0_outputs[12714] = (inputs[74]) & ~(inputs[27]);
    assign layer0_outputs[12715] = (inputs[118]) & ~(inputs[108]);
    assign layer0_outputs[12716] = ~(inputs[6]);
    assign layer0_outputs[12717] = ~((inputs[56]) | (inputs[105]));
    assign layer0_outputs[12718] = (inputs[30]) ^ (inputs[46]);
    assign layer0_outputs[12719] = ~(inputs[232]) | (inputs[222]);
    assign layer0_outputs[12720] = ~(inputs[248]) | (inputs[5]);
    assign layer0_outputs[12721] = (inputs[136]) | (inputs[4]);
    assign layer0_outputs[12722] = ~(inputs[97]) | (inputs[107]);
    assign layer0_outputs[12723] = 1'b1;
    assign layer0_outputs[12724] = (inputs[251]) & ~(inputs[249]);
    assign layer0_outputs[12725] = ~(inputs[244]);
    assign layer0_outputs[12726] = (inputs[149]) & (inputs[188]);
    assign layer0_outputs[12727] = (inputs[85]) | (inputs[72]);
    assign layer0_outputs[12728] = ~(inputs[76]) | (inputs[177]);
    assign layer0_outputs[12729] = ~(inputs[101]);
    assign layer0_outputs[12730] = (inputs[31]) ^ (inputs[92]);
    assign layer0_outputs[12731] = (inputs[196]) | (inputs[141]);
    assign layer0_outputs[12732] = ~((inputs[199]) & (inputs[253]));
    assign layer0_outputs[12733] = ~((inputs[86]) ^ (inputs[19]));
    assign layer0_outputs[12734] = ~(inputs[84]) | (inputs[18]);
    assign layer0_outputs[12735] = (inputs[43]) & ~(inputs[225]);
    assign layer0_outputs[12736] = ~((inputs[214]) ^ (inputs[2]));
    assign layer0_outputs[12737] = (inputs[154]) | (inputs[174]);
    assign layer0_outputs[12738] = ~((inputs[91]) ^ (inputs[78]));
    assign layer0_outputs[12739] = ~((inputs[165]) ^ (inputs[189]));
    assign layer0_outputs[12740] = (inputs[137]) & (inputs[0]);
    assign layer0_outputs[12741] = (inputs[53]) & ~(inputs[150]);
    assign layer0_outputs[12742] = inputs[186];
    assign layer0_outputs[12743] = 1'b1;
    assign layer0_outputs[12744] = ~(inputs[17]) | (inputs[143]);
    assign layer0_outputs[12745] = (inputs[64]) & (inputs[220]);
    assign layer0_outputs[12746] = ~(inputs[178]);
    assign layer0_outputs[12747] = (inputs[18]) ^ (inputs[223]);
    assign layer0_outputs[12748] = inputs[194];
    assign layer0_outputs[12749] = ~((inputs[61]) | (inputs[244]));
    assign layer0_outputs[12750] = inputs[113];
    assign layer0_outputs[12751] = (inputs[56]) & ~(inputs[206]);
    assign layer0_outputs[12752] = ~((inputs[3]) | (inputs[248]));
    assign layer0_outputs[12753] = ~((inputs[236]) ^ (inputs[230]));
    assign layer0_outputs[12754] = inputs[130];
    assign layer0_outputs[12755] = ~(inputs[84]);
    assign layer0_outputs[12756] = (inputs[142]) ^ (inputs[253]);
    assign layer0_outputs[12757] = inputs[73];
    assign layer0_outputs[12758] = (inputs[183]) & ~(inputs[81]);
    assign layer0_outputs[12759] = inputs[64];
    assign layer0_outputs[12760] = ~(inputs[167]) | (inputs[194]);
    assign layer0_outputs[12761] = ~((inputs[176]) | (inputs[254]));
    assign layer0_outputs[12762] = ~(inputs[252]);
    assign layer0_outputs[12763] = ~(inputs[182]) | (inputs[63]);
    assign layer0_outputs[12764] = ~(inputs[9]) | (inputs[131]);
    assign layer0_outputs[12765] = ~(inputs[207]);
    assign layer0_outputs[12766] = inputs[154];
    assign layer0_outputs[12767] = (inputs[140]) ^ (inputs[143]);
    assign layer0_outputs[12768] = ~(inputs[123]);
    assign layer0_outputs[12769] = (inputs[156]) | (inputs[194]);
    assign layer0_outputs[12770] = inputs[227];
    assign layer0_outputs[12771] = ~(inputs[141]);
    assign layer0_outputs[12772] = ~(inputs[188]);
    assign layer0_outputs[12773] = (inputs[38]) & ~(inputs[47]);
    assign layer0_outputs[12774] = inputs[193];
    assign layer0_outputs[12775] = inputs[59];
    assign layer0_outputs[12776] = ~(inputs[46]);
    assign layer0_outputs[12777] = (inputs[59]) & ~(inputs[142]);
    assign layer0_outputs[12778] = (inputs[186]) & ~(inputs[90]);
    assign layer0_outputs[12779] = inputs[68];
    assign layer0_outputs[12780] = ~((inputs[118]) ^ (inputs[72]));
    assign layer0_outputs[12781] = (inputs[89]) & ~(inputs[33]);
    assign layer0_outputs[12782] = (inputs[216]) & ~(inputs[246]);
    assign layer0_outputs[12783] = (inputs[145]) | (inputs[148]);
    assign layer0_outputs[12784] = ~(inputs[139]) | (inputs[94]);
    assign layer0_outputs[12785] = ~(inputs[8]);
    assign layer0_outputs[12786] = (inputs[78]) & ~(inputs[239]);
    assign layer0_outputs[12787] = inputs[178];
    assign layer0_outputs[12788] = ~(inputs[244]);
    assign layer0_outputs[12789] = ~(inputs[150]);
    assign layer0_outputs[12790] = ~((inputs[61]) | (inputs[75]));
    assign layer0_outputs[12791] = ~(inputs[91]);
    assign layer0_outputs[12792] = ~(inputs[116]) | (inputs[163]);
    assign layer0_outputs[12793] = inputs[1];
    assign layer0_outputs[12794] = 1'b0;
    assign layer0_outputs[12795] = inputs[208];
    assign layer0_outputs[12796] = ~(inputs[208]);
    assign layer0_outputs[12797] = (inputs[60]) ^ (inputs[14]);
    assign layer0_outputs[12798] = ~(inputs[64]) | (inputs[30]);
    assign layer0_outputs[12799] = ~((inputs[46]) | (inputs[123]));
    assign layer1_outputs[0] = (layer0_outputs[2066]) | (layer0_outputs[9142]);
    assign layer1_outputs[1] = ~(layer0_outputs[705]);
    assign layer1_outputs[2] = ~((layer0_outputs[1387]) | (layer0_outputs[10225]));
    assign layer1_outputs[3] = (layer0_outputs[5591]) ^ (layer0_outputs[9562]);
    assign layer1_outputs[4] = ~(layer0_outputs[8688]);
    assign layer1_outputs[5] = ~(layer0_outputs[3270]);
    assign layer1_outputs[6] = ~((layer0_outputs[2997]) & (layer0_outputs[1994]));
    assign layer1_outputs[7] = layer0_outputs[8907];
    assign layer1_outputs[8] = (layer0_outputs[5499]) ^ (layer0_outputs[10882]);
    assign layer1_outputs[9] = layer0_outputs[2817];
    assign layer1_outputs[10] = ~(layer0_outputs[1194]);
    assign layer1_outputs[11] = layer0_outputs[8832];
    assign layer1_outputs[12] = ~((layer0_outputs[8879]) ^ (layer0_outputs[3779]));
    assign layer1_outputs[13] = ~(layer0_outputs[2526]);
    assign layer1_outputs[14] = (layer0_outputs[9254]) & ~(layer0_outputs[5661]);
    assign layer1_outputs[15] = ~((layer0_outputs[7713]) & (layer0_outputs[2707]));
    assign layer1_outputs[16] = (layer0_outputs[1237]) | (layer0_outputs[12022]);
    assign layer1_outputs[17] = ~(layer0_outputs[2840]) | (layer0_outputs[1304]);
    assign layer1_outputs[18] = ~(layer0_outputs[12066]);
    assign layer1_outputs[19] = layer0_outputs[12780];
    assign layer1_outputs[20] = ~(layer0_outputs[2087]);
    assign layer1_outputs[21] = layer0_outputs[8733];
    assign layer1_outputs[22] = ~((layer0_outputs[890]) ^ (layer0_outputs[10289]));
    assign layer1_outputs[23] = ~((layer0_outputs[12769]) | (layer0_outputs[8946]));
    assign layer1_outputs[24] = layer0_outputs[12407];
    assign layer1_outputs[25] = layer0_outputs[1013];
    assign layer1_outputs[26] = (layer0_outputs[11276]) & (layer0_outputs[3567]);
    assign layer1_outputs[27] = ~(layer0_outputs[4802]) | (layer0_outputs[955]);
    assign layer1_outputs[28] = layer0_outputs[423];
    assign layer1_outputs[29] = ~(layer0_outputs[7466]) | (layer0_outputs[9592]);
    assign layer1_outputs[30] = ~((layer0_outputs[475]) & (layer0_outputs[945]));
    assign layer1_outputs[31] = ~(layer0_outputs[4034]);
    assign layer1_outputs[32] = (layer0_outputs[11518]) & ~(layer0_outputs[2425]);
    assign layer1_outputs[33] = layer0_outputs[6689];
    assign layer1_outputs[34] = ~((layer0_outputs[8750]) ^ (layer0_outputs[189]));
    assign layer1_outputs[35] = ~(layer0_outputs[998]) | (layer0_outputs[5567]);
    assign layer1_outputs[36] = ~((layer0_outputs[8689]) & (layer0_outputs[2292]));
    assign layer1_outputs[37] = layer0_outputs[1014];
    assign layer1_outputs[38] = ~((layer0_outputs[6853]) ^ (layer0_outputs[9665]));
    assign layer1_outputs[39] = ~((layer0_outputs[212]) & (layer0_outputs[5953]));
    assign layer1_outputs[40] = (layer0_outputs[1191]) & (layer0_outputs[4800]);
    assign layer1_outputs[41] = (layer0_outputs[3065]) | (layer0_outputs[12400]);
    assign layer1_outputs[42] = ~(layer0_outputs[11806]);
    assign layer1_outputs[43] = (layer0_outputs[3684]) | (layer0_outputs[1723]);
    assign layer1_outputs[44] = ~(layer0_outputs[8183]);
    assign layer1_outputs[45] = (layer0_outputs[10209]) & (layer0_outputs[2592]);
    assign layer1_outputs[46] = ~(layer0_outputs[10775]);
    assign layer1_outputs[47] = ~(layer0_outputs[6701]) | (layer0_outputs[4550]);
    assign layer1_outputs[48] = ~(layer0_outputs[11842]);
    assign layer1_outputs[49] = (layer0_outputs[2326]) & (layer0_outputs[1371]);
    assign layer1_outputs[50] = layer0_outputs[456];
    assign layer1_outputs[51] = ~(layer0_outputs[10358]);
    assign layer1_outputs[52] = ~(layer0_outputs[4381]);
    assign layer1_outputs[53] = ~(layer0_outputs[2252]);
    assign layer1_outputs[54] = (layer0_outputs[5988]) | (layer0_outputs[4610]);
    assign layer1_outputs[55] = ~((layer0_outputs[5960]) & (layer0_outputs[10623]));
    assign layer1_outputs[56] = ~(layer0_outputs[1042]) | (layer0_outputs[10528]);
    assign layer1_outputs[57] = layer0_outputs[6841];
    assign layer1_outputs[58] = ~((layer0_outputs[10878]) ^ (layer0_outputs[11074]));
    assign layer1_outputs[59] = 1'b0;
    assign layer1_outputs[60] = ~((layer0_outputs[7915]) | (layer0_outputs[10817]));
    assign layer1_outputs[61] = ~(layer0_outputs[7775]);
    assign layer1_outputs[62] = ~(layer0_outputs[11324]);
    assign layer1_outputs[63] = layer0_outputs[1489];
    assign layer1_outputs[64] = layer0_outputs[1845];
    assign layer1_outputs[65] = ~(layer0_outputs[2430]) | (layer0_outputs[2633]);
    assign layer1_outputs[66] = layer0_outputs[10127];
    assign layer1_outputs[67] = (layer0_outputs[8715]) & ~(layer0_outputs[6801]);
    assign layer1_outputs[68] = layer0_outputs[5514];
    assign layer1_outputs[69] = ~(layer0_outputs[7739]);
    assign layer1_outputs[70] = (layer0_outputs[12275]) ^ (layer0_outputs[3938]);
    assign layer1_outputs[71] = ~(layer0_outputs[5218]);
    assign layer1_outputs[72] = layer0_outputs[9787];
    assign layer1_outputs[73] = layer0_outputs[2995];
    assign layer1_outputs[74] = ~(layer0_outputs[9017]);
    assign layer1_outputs[75] = 1'b1;
    assign layer1_outputs[76] = (layer0_outputs[4841]) | (layer0_outputs[6755]);
    assign layer1_outputs[77] = ~((layer0_outputs[9333]) ^ (layer0_outputs[2163]));
    assign layer1_outputs[78] = layer0_outputs[7021];
    assign layer1_outputs[79] = ~(layer0_outputs[6674]);
    assign layer1_outputs[80] = layer0_outputs[4931];
    assign layer1_outputs[81] = layer0_outputs[10540];
    assign layer1_outputs[82] = ~(layer0_outputs[8770]);
    assign layer1_outputs[83] = layer0_outputs[9503];
    assign layer1_outputs[84] = ~(layer0_outputs[10436]) | (layer0_outputs[8280]);
    assign layer1_outputs[85] = (layer0_outputs[7944]) & (layer0_outputs[5314]);
    assign layer1_outputs[86] = (layer0_outputs[8094]) & ~(layer0_outputs[2361]);
    assign layer1_outputs[87] = ~(layer0_outputs[11629]) | (layer0_outputs[4983]);
    assign layer1_outputs[88] = ~(layer0_outputs[7799]);
    assign layer1_outputs[89] = ~(layer0_outputs[4778]) | (layer0_outputs[10708]);
    assign layer1_outputs[90] = (layer0_outputs[6645]) & ~(layer0_outputs[11251]);
    assign layer1_outputs[91] = (layer0_outputs[4653]) & ~(layer0_outputs[6602]);
    assign layer1_outputs[92] = (layer0_outputs[12388]) & ~(layer0_outputs[7776]);
    assign layer1_outputs[93] = ~((layer0_outputs[2784]) & (layer0_outputs[8239]));
    assign layer1_outputs[94] = ~((layer0_outputs[10645]) & (layer0_outputs[2180]));
    assign layer1_outputs[95] = 1'b1;
    assign layer1_outputs[96] = (layer0_outputs[7947]) ^ (layer0_outputs[3206]);
    assign layer1_outputs[97] = (layer0_outputs[3662]) & (layer0_outputs[10494]);
    assign layer1_outputs[98] = ~(layer0_outputs[6927]);
    assign layer1_outputs[99] = ~(layer0_outputs[12624]) | (layer0_outputs[12657]);
    assign layer1_outputs[100] = (layer0_outputs[6217]) & ~(layer0_outputs[5122]);
    assign layer1_outputs[101] = layer0_outputs[5948];
    assign layer1_outputs[102] = ~(layer0_outputs[2157]);
    assign layer1_outputs[103] = ~(layer0_outputs[4142]);
    assign layer1_outputs[104] = (layer0_outputs[7220]) & (layer0_outputs[3244]);
    assign layer1_outputs[105] = ~(layer0_outputs[8780]) | (layer0_outputs[4581]);
    assign layer1_outputs[106] = (layer0_outputs[11746]) & (layer0_outputs[12422]);
    assign layer1_outputs[107] = ~((layer0_outputs[5231]) & (layer0_outputs[4068]));
    assign layer1_outputs[108] = (layer0_outputs[9329]) & ~(layer0_outputs[8484]);
    assign layer1_outputs[109] = (layer0_outputs[7952]) & ~(layer0_outputs[9678]);
    assign layer1_outputs[110] = layer0_outputs[8199];
    assign layer1_outputs[111] = ~(layer0_outputs[12019]);
    assign layer1_outputs[112] = layer0_outputs[675];
    assign layer1_outputs[113] = (layer0_outputs[8926]) & (layer0_outputs[12146]);
    assign layer1_outputs[114] = (layer0_outputs[10112]) ^ (layer0_outputs[7155]);
    assign layer1_outputs[115] = (layer0_outputs[6344]) & ~(layer0_outputs[7240]);
    assign layer1_outputs[116] = ~((layer0_outputs[1083]) | (layer0_outputs[5652]));
    assign layer1_outputs[117] = ~(layer0_outputs[4734]) | (layer0_outputs[12227]);
    assign layer1_outputs[118] = ~(layer0_outputs[9647]);
    assign layer1_outputs[119] = ~(layer0_outputs[7997]);
    assign layer1_outputs[120] = ~(layer0_outputs[1719]) | (layer0_outputs[2083]);
    assign layer1_outputs[121] = ~((layer0_outputs[10020]) & (layer0_outputs[32]));
    assign layer1_outputs[122] = ~((layer0_outputs[9058]) | (layer0_outputs[4099]));
    assign layer1_outputs[123] = ~((layer0_outputs[9187]) & (layer0_outputs[8732]));
    assign layer1_outputs[124] = (layer0_outputs[1166]) & (layer0_outputs[4036]);
    assign layer1_outputs[125] = ~(layer0_outputs[3944]) | (layer0_outputs[7026]);
    assign layer1_outputs[126] = ~(layer0_outputs[6788]) | (layer0_outputs[5777]);
    assign layer1_outputs[127] = layer0_outputs[4253];
    assign layer1_outputs[128] = ~(layer0_outputs[5497]);
    assign layer1_outputs[129] = ~((layer0_outputs[6690]) | (layer0_outputs[1125]));
    assign layer1_outputs[130] = (layer0_outputs[1706]) ^ (layer0_outputs[9827]);
    assign layer1_outputs[131] = ~((layer0_outputs[5241]) ^ (layer0_outputs[5659]));
    assign layer1_outputs[132] = layer0_outputs[1769];
    assign layer1_outputs[133] = 1'b1;
    assign layer1_outputs[134] = ~((layer0_outputs[9457]) & (layer0_outputs[10544]));
    assign layer1_outputs[135] = (layer0_outputs[1578]) & ~(layer0_outputs[363]);
    assign layer1_outputs[136] = ~(layer0_outputs[5662]);
    assign layer1_outputs[137] = ~(layer0_outputs[9668]) | (layer0_outputs[4490]);
    assign layer1_outputs[138] = ~(layer0_outputs[4217]) | (layer0_outputs[9046]);
    assign layer1_outputs[139] = layer0_outputs[10472];
    assign layer1_outputs[140] = ~(layer0_outputs[1881]) | (layer0_outputs[3124]);
    assign layer1_outputs[141] = ~((layer0_outputs[7577]) ^ (layer0_outputs[6927]));
    assign layer1_outputs[142] = ~(layer0_outputs[2867]);
    assign layer1_outputs[143] = (layer0_outputs[63]) & ~(layer0_outputs[1828]);
    assign layer1_outputs[144] = ~((layer0_outputs[1230]) & (layer0_outputs[9646]));
    assign layer1_outputs[145] = layer0_outputs[2216];
    assign layer1_outputs[146] = ~(layer0_outputs[1433]) | (layer0_outputs[1428]);
    assign layer1_outputs[147] = ~(layer0_outputs[142]);
    assign layer1_outputs[148] = 1'b0;
    assign layer1_outputs[149] = ~((layer0_outputs[7066]) ^ (layer0_outputs[1458]));
    assign layer1_outputs[150] = (layer0_outputs[12200]) & ~(layer0_outputs[7999]);
    assign layer1_outputs[151] = layer0_outputs[4078];
    assign layer1_outputs[152] = (layer0_outputs[3620]) & ~(layer0_outputs[7933]);
    assign layer1_outputs[153] = ~((layer0_outputs[2142]) & (layer0_outputs[1594]));
    assign layer1_outputs[154] = 1'b0;
    assign layer1_outputs[155] = layer0_outputs[9949];
    assign layer1_outputs[156] = (layer0_outputs[6658]) | (layer0_outputs[4776]);
    assign layer1_outputs[157] = ~((layer0_outputs[9802]) | (layer0_outputs[3045]));
    assign layer1_outputs[158] = (layer0_outputs[6095]) & ~(layer0_outputs[2450]);
    assign layer1_outputs[159] = ~((layer0_outputs[727]) & (layer0_outputs[9499]));
    assign layer1_outputs[160] = (layer0_outputs[11583]) ^ (layer0_outputs[11423]);
    assign layer1_outputs[161] = (layer0_outputs[12155]) & (layer0_outputs[2583]);
    assign layer1_outputs[162] = ~(layer0_outputs[12350]) | (layer0_outputs[1233]);
    assign layer1_outputs[163] = ~(layer0_outputs[1375]);
    assign layer1_outputs[164] = ~((layer0_outputs[7764]) | (layer0_outputs[8777]));
    assign layer1_outputs[165] = (layer0_outputs[10011]) | (layer0_outputs[4675]);
    assign layer1_outputs[166] = (layer0_outputs[12082]) & ~(layer0_outputs[556]);
    assign layer1_outputs[167] = ~(layer0_outputs[4097]);
    assign layer1_outputs[168] = ~(layer0_outputs[7367]);
    assign layer1_outputs[169] = layer0_outputs[5948];
    assign layer1_outputs[170] = ~(layer0_outputs[5224]);
    assign layer1_outputs[171] = ~(layer0_outputs[1794]);
    assign layer1_outputs[172] = ~(layer0_outputs[6860]);
    assign layer1_outputs[173] = (layer0_outputs[5758]) & (layer0_outputs[2171]);
    assign layer1_outputs[174] = (layer0_outputs[857]) & (layer0_outputs[6814]);
    assign layer1_outputs[175] = ~(layer0_outputs[6515]);
    assign layer1_outputs[176] = (layer0_outputs[19]) ^ (layer0_outputs[1162]);
    assign layer1_outputs[177] = layer0_outputs[5621];
    assign layer1_outputs[178] = layer0_outputs[795];
    assign layer1_outputs[179] = ~(layer0_outputs[11137]) | (layer0_outputs[8809]);
    assign layer1_outputs[180] = (layer0_outputs[3016]) & ~(layer0_outputs[12180]);
    assign layer1_outputs[181] = ~((layer0_outputs[12472]) & (layer0_outputs[585]));
    assign layer1_outputs[182] = ~(layer0_outputs[10652]);
    assign layer1_outputs[183] = ~(layer0_outputs[3350]) | (layer0_outputs[6695]);
    assign layer1_outputs[184] = ~(layer0_outputs[949]) | (layer0_outputs[11490]);
    assign layer1_outputs[185] = ~(layer0_outputs[1914]);
    assign layer1_outputs[186] = 1'b1;
    assign layer1_outputs[187] = ~(layer0_outputs[12521]);
    assign layer1_outputs[188] = ~(layer0_outputs[5212]);
    assign layer1_outputs[189] = ~(layer0_outputs[8569]);
    assign layer1_outputs[190] = (layer0_outputs[12203]) | (layer0_outputs[2277]);
    assign layer1_outputs[191] = layer0_outputs[4136];
    assign layer1_outputs[192] = layer0_outputs[5582];
    assign layer1_outputs[193] = (layer0_outputs[389]) & (layer0_outputs[5807]);
    assign layer1_outputs[194] = (layer0_outputs[8132]) | (layer0_outputs[6600]);
    assign layer1_outputs[195] = (layer0_outputs[2561]) & ~(layer0_outputs[4950]);
    assign layer1_outputs[196] = ~((layer0_outputs[9697]) | (layer0_outputs[4271]));
    assign layer1_outputs[197] = ~(layer0_outputs[3386]) | (layer0_outputs[6581]);
    assign layer1_outputs[198] = (layer0_outputs[10606]) ^ (layer0_outputs[240]);
    assign layer1_outputs[199] = ~((layer0_outputs[144]) ^ (layer0_outputs[4869]));
    assign layer1_outputs[200] = ~(layer0_outputs[1246]);
    assign layer1_outputs[201] = ~(layer0_outputs[12113]);
    assign layer1_outputs[202] = ~(layer0_outputs[9521]);
    assign layer1_outputs[203] = ~(layer0_outputs[12352]);
    assign layer1_outputs[204] = ~((layer0_outputs[10318]) & (layer0_outputs[9007]));
    assign layer1_outputs[205] = ~(layer0_outputs[8817]) | (layer0_outputs[7965]);
    assign layer1_outputs[206] = (layer0_outputs[5153]) & ~(layer0_outputs[9432]);
    assign layer1_outputs[207] = layer0_outputs[12328];
    assign layer1_outputs[208] = ~((layer0_outputs[11745]) ^ (layer0_outputs[1715]));
    assign layer1_outputs[209] = (layer0_outputs[11131]) & ~(layer0_outputs[7898]);
    assign layer1_outputs[210] = ~((layer0_outputs[12506]) ^ (layer0_outputs[8214]));
    assign layer1_outputs[211] = layer0_outputs[7057];
    assign layer1_outputs[212] = (layer0_outputs[2107]) ^ (layer0_outputs[11208]);
    assign layer1_outputs[213] = ~((layer0_outputs[6294]) & (layer0_outputs[4999]));
    assign layer1_outputs[214] = (layer0_outputs[3444]) & (layer0_outputs[12653]);
    assign layer1_outputs[215] = ~(layer0_outputs[9690]);
    assign layer1_outputs[216] = ~((layer0_outputs[2614]) | (layer0_outputs[5573]));
    assign layer1_outputs[217] = (layer0_outputs[1657]) ^ (layer0_outputs[4166]);
    assign layer1_outputs[218] = ~((layer0_outputs[8325]) ^ (layer0_outputs[972]));
    assign layer1_outputs[219] = ~(layer0_outputs[12393]);
    assign layer1_outputs[220] = layer0_outputs[6117];
    assign layer1_outputs[221] = (layer0_outputs[8905]) & (layer0_outputs[9876]);
    assign layer1_outputs[222] = (layer0_outputs[2842]) | (layer0_outputs[7084]);
    assign layer1_outputs[223] = (layer0_outputs[11099]) | (layer0_outputs[6660]);
    assign layer1_outputs[224] = layer0_outputs[949];
    assign layer1_outputs[225] = ~(layer0_outputs[11783]);
    assign layer1_outputs[226] = (layer0_outputs[2858]) & (layer0_outputs[8535]);
    assign layer1_outputs[227] = layer0_outputs[3212];
    assign layer1_outputs[228] = (layer0_outputs[9614]) & ~(layer0_outputs[2540]);
    assign layer1_outputs[229] = ~((layer0_outputs[6032]) & (layer0_outputs[8250]));
    assign layer1_outputs[230] = layer0_outputs[151];
    assign layer1_outputs[231] = layer0_outputs[3905];
    assign layer1_outputs[232] = ~((layer0_outputs[4125]) & (layer0_outputs[12236]));
    assign layer1_outputs[233] = layer0_outputs[437];
    assign layer1_outputs[234] = (layer0_outputs[9969]) & (layer0_outputs[3841]);
    assign layer1_outputs[235] = layer0_outputs[12255];
    assign layer1_outputs[236] = (layer0_outputs[6563]) & ~(layer0_outputs[1463]);
    assign layer1_outputs[237] = ~(layer0_outputs[2968]);
    assign layer1_outputs[238] = layer0_outputs[6975];
    assign layer1_outputs[239] = layer0_outputs[6205];
    assign layer1_outputs[240] = (layer0_outputs[3589]) | (layer0_outputs[8845]);
    assign layer1_outputs[241] = (layer0_outputs[1720]) ^ (layer0_outputs[11090]);
    assign layer1_outputs[242] = (layer0_outputs[8873]) ^ (layer0_outputs[1328]);
    assign layer1_outputs[243] = (layer0_outputs[1677]) ^ (layer0_outputs[7462]);
    assign layer1_outputs[244] = (layer0_outputs[7007]) & (layer0_outputs[5034]);
    assign layer1_outputs[245] = (layer0_outputs[3529]) & ~(layer0_outputs[6034]);
    assign layer1_outputs[246] = ~((layer0_outputs[6858]) ^ (layer0_outputs[6681]));
    assign layer1_outputs[247] = ~(layer0_outputs[10846]) | (layer0_outputs[1054]);
    assign layer1_outputs[248] = ~((layer0_outputs[5050]) ^ (layer0_outputs[11680]));
    assign layer1_outputs[249] = ~(layer0_outputs[11097]);
    assign layer1_outputs[250] = ~(layer0_outputs[8803]);
    assign layer1_outputs[251] = ~(layer0_outputs[7642]);
    assign layer1_outputs[252] = layer0_outputs[8100];
    assign layer1_outputs[253] = ~((layer0_outputs[11749]) | (layer0_outputs[12536]));
    assign layer1_outputs[254] = ~(layer0_outputs[641]) | (layer0_outputs[786]);
    assign layer1_outputs[255] = ~(layer0_outputs[9222]);
    assign layer1_outputs[256] = ~((layer0_outputs[3944]) | (layer0_outputs[81]));
    assign layer1_outputs[257] = layer0_outputs[10876];
    assign layer1_outputs[258] = ~(layer0_outputs[10228]) | (layer0_outputs[2169]);
    assign layer1_outputs[259] = ~(layer0_outputs[4502]);
    assign layer1_outputs[260] = (layer0_outputs[242]) & (layer0_outputs[7126]);
    assign layer1_outputs[261] = ~((layer0_outputs[1446]) | (layer0_outputs[904]));
    assign layer1_outputs[262] = ~(layer0_outputs[9450]);
    assign layer1_outputs[263] = (layer0_outputs[1044]) & ~(layer0_outputs[4662]);
    assign layer1_outputs[264] = ~(layer0_outputs[7389]);
    assign layer1_outputs[265] = ~(layer0_outputs[12557]);
    assign layer1_outputs[266] = layer0_outputs[5792];
    assign layer1_outputs[267] = layer0_outputs[6538];
    assign layer1_outputs[268] = (layer0_outputs[4442]) & ~(layer0_outputs[8865]);
    assign layer1_outputs[269] = ~((layer0_outputs[6232]) ^ (layer0_outputs[5482]));
    assign layer1_outputs[270] = layer0_outputs[264];
    assign layer1_outputs[271] = (layer0_outputs[11]) ^ (layer0_outputs[6511]);
    assign layer1_outputs[272] = ~(layer0_outputs[9050]);
    assign layer1_outputs[273] = ~((layer0_outputs[11901]) | (layer0_outputs[3333]));
    assign layer1_outputs[274] = layer0_outputs[9441];
    assign layer1_outputs[275] = ~((layer0_outputs[10416]) | (layer0_outputs[7281]));
    assign layer1_outputs[276] = ~((layer0_outputs[1935]) & (layer0_outputs[9282]));
    assign layer1_outputs[277] = ~(layer0_outputs[7215]);
    assign layer1_outputs[278] = ~(layer0_outputs[2740]);
    assign layer1_outputs[279] = ~(layer0_outputs[1493]);
    assign layer1_outputs[280] = (layer0_outputs[9793]) ^ (layer0_outputs[7994]);
    assign layer1_outputs[281] = (layer0_outputs[3091]) ^ (layer0_outputs[10569]);
    assign layer1_outputs[282] = ~(layer0_outputs[1298]);
    assign layer1_outputs[283] = ~(layer0_outputs[9757]);
    assign layer1_outputs[284] = ~(layer0_outputs[8849]) | (layer0_outputs[11879]);
    assign layer1_outputs[285] = layer0_outputs[12223];
    assign layer1_outputs[286] = (layer0_outputs[8603]) & ~(layer0_outputs[7472]);
    assign layer1_outputs[287] = ~(layer0_outputs[10158]);
    assign layer1_outputs[288] = ~(layer0_outputs[4996]);
    assign layer1_outputs[289] = ~(layer0_outputs[10650]);
    assign layer1_outputs[290] = layer0_outputs[6913];
    assign layer1_outputs[291] = ~(layer0_outputs[7178]);
    assign layer1_outputs[292] = ~((layer0_outputs[6846]) | (layer0_outputs[12759]));
    assign layer1_outputs[293] = (layer0_outputs[2124]) | (layer0_outputs[1405]);
    assign layer1_outputs[294] = layer0_outputs[10394];
    assign layer1_outputs[295] = (layer0_outputs[11555]) & ~(layer0_outputs[4822]);
    assign layer1_outputs[296] = ~((layer0_outputs[10727]) & (layer0_outputs[473]));
    assign layer1_outputs[297] = ~(layer0_outputs[2902]);
    assign layer1_outputs[298] = (layer0_outputs[8700]) | (layer0_outputs[12791]);
    assign layer1_outputs[299] = layer0_outputs[12411];
    assign layer1_outputs[300] = ~(layer0_outputs[4350]) | (layer0_outputs[2040]);
    assign layer1_outputs[301] = layer0_outputs[6561];
    assign layer1_outputs[302] = layer0_outputs[3566];
    assign layer1_outputs[303] = ~(layer0_outputs[12387]) | (layer0_outputs[7237]);
    assign layer1_outputs[304] = layer0_outputs[398];
    assign layer1_outputs[305] = ~(layer0_outputs[6756]);
    assign layer1_outputs[306] = layer0_outputs[2807];
    assign layer1_outputs[307] = (layer0_outputs[7804]) & (layer0_outputs[2138]);
    assign layer1_outputs[308] = ~(layer0_outputs[55]) | (layer0_outputs[9987]);
    assign layer1_outputs[309] = (layer0_outputs[1636]) | (layer0_outputs[5931]);
    assign layer1_outputs[310] = 1'b0;
    assign layer1_outputs[311] = ~(layer0_outputs[12364]);
    assign layer1_outputs[312] = ~((layer0_outputs[1087]) & (layer0_outputs[5429]));
    assign layer1_outputs[313] = ~((layer0_outputs[4774]) | (layer0_outputs[1144]));
    assign layer1_outputs[314] = ~((layer0_outputs[11510]) ^ (layer0_outputs[1715]));
    assign layer1_outputs[315] = ~(layer0_outputs[4745]) | (layer0_outputs[7320]);
    assign layer1_outputs[316] = ~(layer0_outputs[11404]);
    assign layer1_outputs[317] = ~((layer0_outputs[6666]) | (layer0_outputs[11875]));
    assign layer1_outputs[318] = ~(layer0_outputs[10784]);
    assign layer1_outputs[319] = 1'b1;
    assign layer1_outputs[320] = ~(layer0_outputs[1045]);
    assign layer1_outputs[321] = ~(layer0_outputs[4605]) | (layer0_outputs[11366]);
    assign layer1_outputs[322] = layer0_outputs[921];
    assign layer1_outputs[323] = (layer0_outputs[10583]) | (layer0_outputs[12692]);
    assign layer1_outputs[324] = ~(layer0_outputs[12645]);
    assign layer1_outputs[325] = (layer0_outputs[10512]) | (layer0_outputs[5163]);
    assign layer1_outputs[326] = ~((layer0_outputs[1953]) ^ (layer0_outputs[3143]));
    assign layer1_outputs[327] = ~(layer0_outputs[4650]);
    assign layer1_outputs[328] = ~((layer0_outputs[2794]) | (layer0_outputs[7908]));
    assign layer1_outputs[329] = ~(layer0_outputs[6902]);
    assign layer1_outputs[330] = ~(layer0_outputs[5551]) | (layer0_outputs[8274]);
    assign layer1_outputs[331] = (layer0_outputs[3581]) & (layer0_outputs[1043]);
    assign layer1_outputs[332] = ~((layer0_outputs[8459]) ^ (layer0_outputs[8166]));
    assign layer1_outputs[333] = layer0_outputs[8016];
    assign layer1_outputs[334] = ~(layer0_outputs[5254]);
    assign layer1_outputs[335] = ~((layer0_outputs[12036]) | (layer0_outputs[134]));
    assign layer1_outputs[336] = layer0_outputs[1631];
    assign layer1_outputs[337] = layer0_outputs[1048];
    assign layer1_outputs[338] = layer0_outputs[7335];
    assign layer1_outputs[339] = (layer0_outputs[9416]) | (layer0_outputs[4641]);
    assign layer1_outputs[340] = ~(layer0_outputs[5679]) | (layer0_outputs[5503]);
    assign layer1_outputs[341] = (layer0_outputs[11730]) & (layer0_outputs[8668]);
    assign layer1_outputs[342] = ~((layer0_outputs[11257]) ^ (layer0_outputs[4446]));
    assign layer1_outputs[343] = (layer0_outputs[3798]) & ~(layer0_outputs[10909]);
    assign layer1_outputs[344] = layer0_outputs[581];
    assign layer1_outputs[345] = ~((layer0_outputs[10128]) ^ (layer0_outputs[8861]));
    assign layer1_outputs[346] = ~(layer0_outputs[3033]);
    assign layer1_outputs[347] = ~((layer0_outputs[7357]) & (layer0_outputs[2786]));
    assign layer1_outputs[348] = layer0_outputs[11839];
    assign layer1_outputs[349] = 1'b1;
    assign layer1_outputs[350] = ~(layer0_outputs[8577]);
    assign layer1_outputs[351] = (layer0_outputs[11867]) & ~(layer0_outputs[1594]);
    assign layer1_outputs[352] = ~(layer0_outputs[8238]);
    assign layer1_outputs[353] = ~(layer0_outputs[2163]) | (layer0_outputs[8871]);
    assign layer1_outputs[354] = (layer0_outputs[11289]) ^ (layer0_outputs[5570]);
    assign layer1_outputs[355] = (layer0_outputs[10685]) & (layer0_outputs[724]);
    assign layer1_outputs[356] = ~(layer0_outputs[660]);
    assign layer1_outputs[357] = (layer0_outputs[8800]) | (layer0_outputs[5112]);
    assign layer1_outputs[358] = ~(layer0_outputs[10459]) | (layer0_outputs[405]);
    assign layer1_outputs[359] = ~(layer0_outputs[11389]);
    assign layer1_outputs[360] = (layer0_outputs[4593]) | (layer0_outputs[642]);
    assign layer1_outputs[361] = ~(layer0_outputs[3375]);
    assign layer1_outputs[362] = ~((layer0_outputs[12568]) & (layer0_outputs[8151]));
    assign layer1_outputs[363] = ~((layer0_outputs[9330]) | (layer0_outputs[9407]));
    assign layer1_outputs[364] = ~(layer0_outputs[6419]) | (layer0_outputs[8527]);
    assign layer1_outputs[365] = ~(layer0_outputs[640]) | (layer0_outputs[1972]);
    assign layer1_outputs[366] = ~(layer0_outputs[6650]);
    assign layer1_outputs[367] = ~((layer0_outputs[2469]) ^ (layer0_outputs[10243]));
    assign layer1_outputs[368] = layer0_outputs[10129];
    assign layer1_outputs[369] = layer0_outputs[6401];
    assign layer1_outputs[370] = ~((layer0_outputs[7401]) & (layer0_outputs[11902]));
    assign layer1_outputs[371] = (layer0_outputs[1826]) & (layer0_outputs[2769]);
    assign layer1_outputs[372] = ~(layer0_outputs[4649]) | (layer0_outputs[6417]);
    assign layer1_outputs[373] = (layer0_outputs[8207]) & ~(layer0_outputs[9836]);
    assign layer1_outputs[374] = ~((layer0_outputs[1630]) ^ (layer0_outputs[6482]));
    assign layer1_outputs[375] = (layer0_outputs[2849]) & (layer0_outputs[10568]);
    assign layer1_outputs[376] = 1'b1;
    assign layer1_outputs[377] = ~((layer0_outputs[8827]) ^ (layer0_outputs[5398]));
    assign layer1_outputs[378] = ~(layer0_outputs[10101]) | (layer0_outputs[6297]);
    assign layer1_outputs[379] = ~(layer0_outputs[9931]);
    assign layer1_outputs[380] = ~((layer0_outputs[12432]) | (layer0_outputs[3622]));
    assign layer1_outputs[381] = ~(layer0_outputs[6252]) | (layer0_outputs[11712]);
    assign layer1_outputs[382] = layer0_outputs[6146];
    assign layer1_outputs[383] = 1'b1;
    assign layer1_outputs[384] = ~(layer0_outputs[7334]) | (layer0_outputs[8290]);
    assign layer1_outputs[385] = layer0_outputs[5783];
    assign layer1_outputs[386] = ~(layer0_outputs[7506]);
    assign layer1_outputs[387] = ~(layer0_outputs[5461]);
    assign layer1_outputs[388] = (layer0_outputs[9350]) & ~(layer0_outputs[1951]);
    assign layer1_outputs[389] = layer0_outputs[9468];
    assign layer1_outputs[390] = ~(layer0_outputs[12737]) | (layer0_outputs[7391]);
    assign layer1_outputs[391] = layer0_outputs[3776];
    assign layer1_outputs[392] = ~(layer0_outputs[3439]);
    assign layer1_outputs[393] = ~(layer0_outputs[175]) | (layer0_outputs[1346]);
    assign layer1_outputs[394] = (layer0_outputs[7227]) & ~(layer0_outputs[2358]);
    assign layer1_outputs[395] = (layer0_outputs[3035]) | (layer0_outputs[1948]);
    assign layer1_outputs[396] = ~((layer0_outputs[11049]) ^ (layer0_outputs[1075]));
    assign layer1_outputs[397] = (layer0_outputs[6907]) | (layer0_outputs[6974]);
    assign layer1_outputs[398] = ~(layer0_outputs[12370]);
    assign layer1_outputs[399] = layer0_outputs[294];
    assign layer1_outputs[400] = 1'b0;
    assign layer1_outputs[401] = ~(layer0_outputs[11084]);
    assign layer1_outputs[402] = layer0_outputs[4353];
    assign layer1_outputs[403] = (layer0_outputs[3732]) | (layer0_outputs[1124]);
    assign layer1_outputs[404] = ~(layer0_outputs[8968]);
    assign layer1_outputs[405] = ~((layer0_outputs[5006]) ^ (layer0_outputs[58]));
    assign layer1_outputs[406] = layer0_outputs[10201];
    assign layer1_outputs[407] = ~(layer0_outputs[1802]) | (layer0_outputs[2316]);
    assign layer1_outputs[408] = (layer0_outputs[11879]) & ~(layer0_outputs[10384]);
    assign layer1_outputs[409] = ~(layer0_outputs[10422]);
    assign layer1_outputs[410] = ~(layer0_outputs[5716]);
    assign layer1_outputs[411] = ~(layer0_outputs[825]);
    assign layer1_outputs[412] = layer0_outputs[5183];
    assign layer1_outputs[413] = layer0_outputs[11030];
    assign layer1_outputs[414] = ~(layer0_outputs[6686]) | (layer0_outputs[10253]);
    assign layer1_outputs[415] = ~((layer0_outputs[1438]) & (layer0_outputs[9762]));
    assign layer1_outputs[416] = ~(layer0_outputs[1058]);
    assign layer1_outputs[417] = ~(layer0_outputs[2949]);
    assign layer1_outputs[418] = ~((layer0_outputs[2299]) ^ (layer0_outputs[5475]));
    assign layer1_outputs[419] = layer0_outputs[10410];
    assign layer1_outputs[420] = ~(layer0_outputs[10347]);
    assign layer1_outputs[421] = layer0_outputs[3960];
    assign layer1_outputs[422] = layer0_outputs[8252];
    assign layer1_outputs[423] = ~(layer0_outputs[7476]) | (layer0_outputs[11668]);
    assign layer1_outputs[424] = layer0_outputs[2531];
    assign layer1_outputs[425] = ~(layer0_outputs[10743]) | (layer0_outputs[11146]);
    assign layer1_outputs[426] = layer0_outputs[2349];
    assign layer1_outputs[427] = layer0_outputs[11544];
    assign layer1_outputs[428] = ~(layer0_outputs[11720]);
    assign layer1_outputs[429] = ~(layer0_outputs[11176]);
    assign layer1_outputs[430] = ~((layer0_outputs[2879]) ^ (layer0_outputs[874]));
    assign layer1_outputs[431] = ~((layer0_outputs[9444]) ^ (layer0_outputs[2862]));
    assign layer1_outputs[432] = layer0_outputs[3719];
    assign layer1_outputs[433] = ~(layer0_outputs[12706]);
    assign layer1_outputs[434] = (layer0_outputs[6938]) ^ (layer0_outputs[7064]);
    assign layer1_outputs[435] = (layer0_outputs[1397]) & (layer0_outputs[10603]);
    assign layer1_outputs[436] = (layer0_outputs[10970]) & ~(layer0_outputs[5341]);
    assign layer1_outputs[437] = layer0_outputs[12372];
    assign layer1_outputs[438] = layer0_outputs[331];
    assign layer1_outputs[439] = layer0_outputs[8085];
    assign layer1_outputs[440] = layer0_outputs[8192];
    assign layer1_outputs[441] = layer0_outputs[1196];
    assign layer1_outputs[442] = ~(layer0_outputs[12621]);
    assign layer1_outputs[443] = ~((layer0_outputs[8283]) ^ (layer0_outputs[9911]));
    assign layer1_outputs[444] = ~((layer0_outputs[526]) ^ (layer0_outputs[11427]));
    assign layer1_outputs[445] = layer0_outputs[10490];
    assign layer1_outputs[446] = layer0_outputs[12587];
    assign layer1_outputs[447] = ~(layer0_outputs[2103]) | (layer0_outputs[10946]);
    assign layer1_outputs[448] = ~((layer0_outputs[4522]) | (layer0_outputs[1062]));
    assign layer1_outputs[449] = (layer0_outputs[11001]) | (layer0_outputs[9088]);
    assign layer1_outputs[450] = ~((layer0_outputs[4905]) & (layer0_outputs[12015]));
    assign layer1_outputs[451] = layer0_outputs[12560];
    assign layer1_outputs[452] = ~(layer0_outputs[11002]);
    assign layer1_outputs[453] = (layer0_outputs[1973]) ^ (layer0_outputs[8308]);
    assign layer1_outputs[454] = ~(layer0_outputs[5541]) | (layer0_outputs[214]);
    assign layer1_outputs[455] = layer0_outputs[12566];
    assign layer1_outputs[456] = ~(layer0_outputs[10277]);
    assign layer1_outputs[457] = ~((layer0_outputs[11497]) | (layer0_outputs[9593]));
    assign layer1_outputs[458] = layer0_outputs[3356];
    assign layer1_outputs[459] = (layer0_outputs[4424]) & (layer0_outputs[11120]);
    assign layer1_outputs[460] = (layer0_outputs[6243]) & (layer0_outputs[1343]);
    assign layer1_outputs[461] = (layer0_outputs[11969]) & ~(layer0_outputs[10147]);
    assign layer1_outputs[462] = ~(layer0_outputs[7259]) | (layer0_outputs[9973]);
    assign layer1_outputs[463] = (layer0_outputs[8412]) ^ (layer0_outputs[11193]);
    assign layer1_outputs[464] = ~(layer0_outputs[8626]);
    assign layer1_outputs[465] = (layer0_outputs[5578]) & ~(layer0_outputs[8146]);
    assign layer1_outputs[466] = layer0_outputs[3480];
    assign layer1_outputs[467] = ~(layer0_outputs[1479]);
    assign layer1_outputs[468] = layer0_outputs[85];
    assign layer1_outputs[469] = ~(layer0_outputs[8614]) | (layer0_outputs[9621]);
    assign layer1_outputs[470] = ~(layer0_outputs[4671]);
    assign layer1_outputs[471] = ~(layer0_outputs[429]);
    assign layer1_outputs[472] = (layer0_outputs[1038]) | (layer0_outputs[7271]);
    assign layer1_outputs[473] = (layer0_outputs[9705]) & ~(layer0_outputs[4854]);
    assign layer1_outputs[474] = ~(layer0_outputs[11058]);
    assign layer1_outputs[475] = (layer0_outputs[6314]) & ~(layer0_outputs[9656]);
    assign layer1_outputs[476] = (layer0_outputs[11385]) & (layer0_outputs[8999]);
    assign layer1_outputs[477] = ~(layer0_outputs[10108]);
    assign layer1_outputs[478] = (layer0_outputs[6769]) | (layer0_outputs[795]);
    assign layer1_outputs[479] = (layer0_outputs[5159]) ^ (layer0_outputs[1220]);
    assign layer1_outputs[480] = (layer0_outputs[11882]) & ~(layer0_outputs[3178]);
    assign layer1_outputs[481] = layer0_outputs[5914];
    assign layer1_outputs[482] = ~(layer0_outputs[9926]);
    assign layer1_outputs[483] = ~(layer0_outputs[5675]);
    assign layer1_outputs[484] = ~(layer0_outputs[7175]);
    assign layer1_outputs[485] = (layer0_outputs[8386]) ^ (layer0_outputs[12607]);
    assign layer1_outputs[486] = ~((layer0_outputs[6125]) ^ (layer0_outputs[7085]));
    assign layer1_outputs[487] = (layer0_outputs[2388]) | (layer0_outputs[281]);
    assign layer1_outputs[488] = ~(layer0_outputs[2288]);
    assign layer1_outputs[489] = ~(layer0_outputs[7225]);
    assign layer1_outputs[490] = (layer0_outputs[533]) & ~(layer0_outputs[4622]);
    assign layer1_outputs[491] = ~((layer0_outputs[3977]) ^ (layer0_outputs[3451]));
    assign layer1_outputs[492] = (layer0_outputs[10907]) & (layer0_outputs[6496]);
    assign layer1_outputs[493] = ~(layer0_outputs[10925]);
    assign layer1_outputs[494] = ~(layer0_outputs[217]);
    assign layer1_outputs[495] = (layer0_outputs[11361]) & ~(layer0_outputs[3217]);
    assign layer1_outputs[496] = ~(layer0_outputs[12153]);
    assign layer1_outputs[497] = ~(layer0_outputs[11106]);
    assign layer1_outputs[498] = ~(layer0_outputs[2364]);
    assign layer1_outputs[499] = ~(layer0_outputs[1296]);
    assign layer1_outputs[500] = 1'b1;
    assign layer1_outputs[501] = ~(layer0_outputs[2930]);
    assign layer1_outputs[502] = ~(layer0_outputs[7308]) | (layer0_outputs[615]);
    assign layer1_outputs[503] = layer0_outputs[3725];
    assign layer1_outputs[504] = ~(layer0_outputs[4444]);
    assign layer1_outputs[505] = (layer0_outputs[7498]) & ~(layer0_outputs[4120]);
    assign layer1_outputs[506] = layer0_outputs[2174];
    assign layer1_outputs[507] = layer0_outputs[10562];
    assign layer1_outputs[508] = ~((layer0_outputs[132]) & (layer0_outputs[2902]));
    assign layer1_outputs[509] = ~(layer0_outputs[9207]);
    assign layer1_outputs[510] = (layer0_outputs[9102]) ^ (layer0_outputs[5056]);
    assign layer1_outputs[511] = ~(layer0_outputs[7670]) | (layer0_outputs[3448]);
    assign layer1_outputs[512] = ~((layer0_outputs[10103]) | (layer0_outputs[4658]));
    assign layer1_outputs[513] = ~(layer0_outputs[12746]) | (layer0_outputs[8956]);
    assign layer1_outputs[514] = ~(layer0_outputs[2768]) | (layer0_outputs[203]);
    assign layer1_outputs[515] = layer0_outputs[10338];
    assign layer1_outputs[516] = (layer0_outputs[4427]) & ~(layer0_outputs[3994]);
    assign layer1_outputs[517] = layer0_outputs[1728];
    assign layer1_outputs[518] = ~(layer0_outputs[11686]);
    assign layer1_outputs[519] = ~((layer0_outputs[1445]) ^ (layer0_outputs[5168]));
    assign layer1_outputs[520] = (layer0_outputs[412]) & (layer0_outputs[10843]);
    assign layer1_outputs[521] = (layer0_outputs[1940]) ^ (layer0_outputs[3560]);
    assign layer1_outputs[522] = ~(layer0_outputs[9314]) | (layer0_outputs[6306]);
    assign layer1_outputs[523] = (layer0_outputs[7480]) ^ (layer0_outputs[11944]);
    assign layer1_outputs[524] = (layer0_outputs[6691]) ^ (layer0_outputs[9140]);
    assign layer1_outputs[525] = ~(layer0_outputs[7534]);
    assign layer1_outputs[526] = ~(layer0_outputs[6]);
    assign layer1_outputs[527] = ~((layer0_outputs[7526]) | (layer0_outputs[7104]));
    assign layer1_outputs[528] = 1'b1;
    assign layer1_outputs[529] = layer0_outputs[2459];
    assign layer1_outputs[530] = ~(layer0_outputs[5622]) | (layer0_outputs[5732]);
    assign layer1_outputs[531] = layer0_outputs[8311];
    assign layer1_outputs[532] = layer0_outputs[2882];
    assign layer1_outputs[533] = ~(layer0_outputs[8223]);
    assign layer1_outputs[534] = ~(layer0_outputs[1281]);
    assign layer1_outputs[535] = layer0_outputs[5389];
    assign layer1_outputs[536] = (layer0_outputs[8656]) ^ (layer0_outputs[3974]);
    assign layer1_outputs[537] = 1'b0;
    assign layer1_outputs[538] = ~(layer0_outputs[4319]);
    assign layer1_outputs[539] = ~((layer0_outputs[1821]) | (layer0_outputs[7378]));
    assign layer1_outputs[540] = layer0_outputs[3567];
    assign layer1_outputs[541] = ~((layer0_outputs[2626]) ^ (layer0_outputs[2272]));
    assign layer1_outputs[542] = (layer0_outputs[2688]) & ~(layer0_outputs[3096]);
    assign layer1_outputs[543] = layer0_outputs[9628];
    assign layer1_outputs[544] = ~(layer0_outputs[11967]);
    assign layer1_outputs[545] = ~(layer0_outputs[8929]);
    assign layer1_outputs[546] = 1'b1;
    assign layer1_outputs[547] = (layer0_outputs[943]) ^ (layer0_outputs[10067]);
    assign layer1_outputs[548] = (layer0_outputs[1502]) & ~(layer0_outputs[4964]);
    assign layer1_outputs[549] = ~(layer0_outputs[8170]) | (layer0_outputs[9752]);
    assign layer1_outputs[550] = (layer0_outputs[329]) ^ (layer0_outputs[12120]);
    assign layer1_outputs[551] = (layer0_outputs[1680]) & ~(layer0_outputs[1284]);
    assign layer1_outputs[552] = layer0_outputs[2578];
    assign layer1_outputs[553] = ~((layer0_outputs[3269]) ^ (layer0_outputs[5825]));
    assign layer1_outputs[554] = ~(layer0_outputs[2100]);
    assign layer1_outputs[555] = (layer0_outputs[1569]) & ~(layer0_outputs[6046]);
    assign layer1_outputs[556] = (layer0_outputs[5084]) ^ (layer0_outputs[5798]);
    assign layer1_outputs[557] = 1'b0;
    assign layer1_outputs[558] = ~(layer0_outputs[6333]) | (layer0_outputs[2985]);
    assign layer1_outputs[559] = ~(layer0_outputs[4998]);
    assign layer1_outputs[560] = (layer0_outputs[5725]) & (layer0_outputs[7874]);
    assign layer1_outputs[561] = layer0_outputs[7643];
    assign layer1_outputs[562] = ~(layer0_outputs[10621]) | (layer0_outputs[7867]);
    assign layer1_outputs[563] = (layer0_outputs[6628]) & (layer0_outputs[683]);
    assign layer1_outputs[564] = ~(layer0_outputs[9531]);
    assign layer1_outputs[565] = (layer0_outputs[1143]) & ~(layer0_outputs[6333]);
    assign layer1_outputs[566] = ~(layer0_outputs[11224]) | (layer0_outputs[4035]);
    assign layer1_outputs[567] = ~((layer0_outputs[4164]) ^ (layer0_outputs[5906]));
    assign layer1_outputs[568] = ~(layer0_outputs[1347]);
    assign layer1_outputs[569] = ~(layer0_outputs[10025]);
    assign layer1_outputs[570] = ~(layer0_outputs[10832]);
    assign layer1_outputs[571] = ~(layer0_outputs[9898]);
    assign layer1_outputs[572] = (layer0_outputs[3828]) ^ (layer0_outputs[12660]);
    assign layer1_outputs[573] = layer0_outputs[1278];
    assign layer1_outputs[574] = ~((layer0_outputs[6079]) ^ (layer0_outputs[10707]));
    assign layer1_outputs[575] = ~((layer0_outputs[12329]) ^ (layer0_outputs[7055]));
    assign layer1_outputs[576] = ~((layer0_outputs[7945]) | (layer0_outputs[10235]));
    assign layer1_outputs[577] = ~((layer0_outputs[11090]) | (layer0_outputs[11685]));
    assign layer1_outputs[578] = ~(layer0_outputs[682]) | (layer0_outputs[5144]);
    assign layer1_outputs[579] = (layer0_outputs[3099]) & ~(layer0_outputs[4330]);
    assign layer1_outputs[580] = ~((layer0_outputs[6560]) & (layer0_outputs[9228]));
    assign layer1_outputs[581] = (layer0_outputs[5891]) ^ (layer0_outputs[10144]);
    assign layer1_outputs[582] = ~(layer0_outputs[6349]);
    assign layer1_outputs[583] = (layer0_outputs[9916]) & ~(layer0_outputs[3602]);
    assign layer1_outputs[584] = (layer0_outputs[12687]) & ~(layer0_outputs[10246]);
    assign layer1_outputs[585] = ~((layer0_outputs[3616]) ^ (layer0_outputs[10806]));
    assign layer1_outputs[586] = ~(layer0_outputs[12418]) | (layer0_outputs[1211]);
    assign layer1_outputs[587] = layer0_outputs[7198];
    assign layer1_outputs[588] = ~(layer0_outputs[4505]);
    assign layer1_outputs[589] = (layer0_outputs[9054]) | (layer0_outputs[8699]);
    assign layer1_outputs[590] = layer0_outputs[6885];
    assign layer1_outputs[591] = ~(layer0_outputs[1139]);
    assign layer1_outputs[592] = (layer0_outputs[513]) & ~(layer0_outputs[9735]);
    assign layer1_outputs[593] = ~(layer0_outputs[10200]);
    assign layer1_outputs[594] = ~((layer0_outputs[9065]) ^ (layer0_outputs[2802]));
    assign layer1_outputs[595] = ~((layer0_outputs[1236]) ^ (layer0_outputs[11409]));
    assign layer1_outputs[596] = (layer0_outputs[7221]) & ~(layer0_outputs[2903]);
    assign layer1_outputs[597] = ~(layer0_outputs[3037]);
    assign layer1_outputs[598] = (layer0_outputs[5359]) & (layer0_outputs[3251]);
    assign layer1_outputs[599] = layer0_outputs[7928];
    assign layer1_outputs[600] = ~(layer0_outputs[599]);
    assign layer1_outputs[601] = (layer0_outputs[884]) & (layer0_outputs[6705]);
    assign layer1_outputs[602] = layer0_outputs[5715];
    assign layer1_outputs[603] = ~(layer0_outputs[2982]);
    assign layer1_outputs[604] = layer0_outputs[6049];
    assign layer1_outputs[605] = (layer0_outputs[8495]) & ~(layer0_outputs[3168]);
    assign layer1_outputs[606] = (layer0_outputs[10550]) & ~(layer0_outputs[3904]);
    assign layer1_outputs[607] = ~(layer0_outputs[424]);
    assign layer1_outputs[608] = ~(layer0_outputs[1242]) | (layer0_outputs[4951]);
    assign layer1_outputs[609] = ~((layer0_outputs[5409]) ^ (layer0_outputs[8821]));
    assign layer1_outputs[610] = ~((layer0_outputs[12464]) & (layer0_outputs[12144]));
    assign layer1_outputs[611] = ~(layer0_outputs[7570]);
    assign layer1_outputs[612] = ~(layer0_outputs[9593]) | (layer0_outputs[5097]);
    assign layer1_outputs[613] = ~(layer0_outputs[3207]);
    assign layer1_outputs[614] = ~(layer0_outputs[5911]);
    assign layer1_outputs[615] = layer0_outputs[9551];
    assign layer1_outputs[616] = 1'b0;
    assign layer1_outputs[617] = layer0_outputs[9518];
    assign layer1_outputs[618] = ~(layer0_outputs[1036]);
    assign layer1_outputs[619] = 1'b0;
    assign layer1_outputs[620] = layer0_outputs[6132];
    assign layer1_outputs[621] = (layer0_outputs[9922]) & (layer0_outputs[9737]);
    assign layer1_outputs[622] = layer0_outputs[10638];
    assign layer1_outputs[623] = ~((layer0_outputs[11398]) | (layer0_outputs[10424]));
    assign layer1_outputs[624] = layer0_outputs[12339];
    assign layer1_outputs[625] = ~(layer0_outputs[6109]) | (layer0_outputs[11898]);
    assign layer1_outputs[626] = layer0_outputs[6354];
    assign layer1_outputs[627] = ~(layer0_outputs[5503]);
    assign layer1_outputs[628] = ~((layer0_outputs[11731]) ^ (layer0_outputs[3154]));
    assign layer1_outputs[629] = ~(layer0_outputs[11673]) | (layer0_outputs[10511]);
    assign layer1_outputs[630] = ~(layer0_outputs[12529]);
    assign layer1_outputs[631] = (layer0_outputs[6483]) & (layer0_outputs[9712]);
    assign layer1_outputs[632] = layer0_outputs[9369];
    assign layer1_outputs[633] = (layer0_outputs[2613]) | (layer0_outputs[6871]);
    assign layer1_outputs[634] = (layer0_outputs[1752]) & (layer0_outputs[3958]);
    assign layer1_outputs[635] = ~(layer0_outputs[6345]);
    assign layer1_outputs[636] = (layer0_outputs[2140]) ^ (layer0_outputs[631]);
    assign layer1_outputs[637] = ~((layer0_outputs[6705]) & (layer0_outputs[1742]));
    assign layer1_outputs[638] = layer0_outputs[4182];
    assign layer1_outputs[639] = (layer0_outputs[8195]) & ~(layer0_outputs[4969]);
    assign layer1_outputs[640] = layer0_outputs[9871];
    assign layer1_outputs[641] = (layer0_outputs[4765]) & ~(layer0_outputs[5088]);
    assign layer1_outputs[642] = (layer0_outputs[6279]) ^ (layer0_outputs[12456]);
    assign layer1_outputs[643] = (layer0_outputs[2448]) | (layer0_outputs[1582]);
    assign layer1_outputs[644] = ~((layer0_outputs[6439]) & (layer0_outputs[9382]));
    assign layer1_outputs[645] = ~(layer0_outputs[11714]);
    assign layer1_outputs[646] = (layer0_outputs[12311]) & ~(layer0_outputs[4304]);
    assign layer1_outputs[647] = (layer0_outputs[11294]) ^ (layer0_outputs[11722]);
    assign layer1_outputs[648] = layer0_outputs[6189];
    assign layer1_outputs[649] = ~(layer0_outputs[5114]) | (layer0_outputs[11179]);
    assign layer1_outputs[650] = ~(layer0_outputs[10096]);
    assign layer1_outputs[651] = layer0_outputs[6488];
    assign layer1_outputs[652] = ~(layer0_outputs[5274]);
    assign layer1_outputs[653] = ~(layer0_outputs[3935]) | (layer0_outputs[11087]);
    assign layer1_outputs[654] = ~(layer0_outputs[8860]) | (layer0_outputs[9410]);
    assign layer1_outputs[655] = (layer0_outputs[2290]) & ~(layer0_outputs[7640]);
    assign layer1_outputs[656] = ~(layer0_outputs[10191]);
    assign layer1_outputs[657] = (layer0_outputs[3179]) ^ (layer0_outputs[6859]);
    assign layer1_outputs[658] = (layer0_outputs[7878]) ^ (layer0_outputs[9491]);
    assign layer1_outputs[659] = (layer0_outputs[1315]) & ~(layer0_outputs[9420]);
    assign layer1_outputs[660] = (layer0_outputs[3300]) ^ (layer0_outputs[758]);
    assign layer1_outputs[661] = (layer0_outputs[2523]) ^ (layer0_outputs[885]);
    assign layer1_outputs[662] = ~((layer0_outputs[12444]) | (layer0_outputs[5683]));
    assign layer1_outputs[663] = ~(layer0_outputs[9624]) | (layer0_outputs[3667]);
    assign layer1_outputs[664] = layer0_outputs[9765];
    assign layer1_outputs[665] = ~((layer0_outputs[8842]) | (layer0_outputs[6864]));
    assign layer1_outputs[666] = 1'b1;
    assign layer1_outputs[667] = ~(layer0_outputs[10349]);
    assign layer1_outputs[668] = (layer0_outputs[7671]) & (layer0_outputs[6252]);
    assign layer1_outputs[669] = ~((layer0_outputs[3868]) | (layer0_outputs[6789]));
    assign layer1_outputs[670] = (layer0_outputs[8020]) & ~(layer0_outputs[3853]);
    assign layer1_outputs[671] = ~((layer0_outputs[7504]) & (layer0_outputs[10588]));
    assign layer1_outputs[672] = layer0_outputs[416];
    assign layer1_outputs[673] = ~(layer0_outputs[5219]);
    assign layer1_outputs[674] = layer0_outputs[10760];
    assign layer1_outputs[675] = ~((layer0_outputs[9004]) | (layer0_outputs[7675]));
    assign layer1_outputs[676] = ~(layer0_outputs[1694]);
    assign layer1_outputs[677] = layer0_outputs[11053];
    assign layer1_outputs[678] = ~((layer0_outputs[7549]) ^ (layer0_outputs[7608]));
    assign layer1_outputs[679] = layer0_outputs[8302];
    assign layer1_outputs[680] = ~(layer0_outputs[12383]) | (layer0_outputs[4928]);
    assign layer1_outputs[681] = ~((layer0_outputs[9131]) & (layer0_outputs[9235]));
    assign layer1_outputs[682] = (layer0_outputs[7744]) & ~(layer0_outputs[10427]);
    assign layer1_outputs[683] = ~(layer0_outputs[9463]);
    assign layer1_outputs[684] = ~((layer0_outputs[12754]) | (layer0_outputs[2953]));
    assign layer1_outputs[685] = layer0_outputs[2145];
    assign layer1_outputs[686] = (layer0_outputs[813]) & (layer0_outputs[2231]);
    assign layer1_outputs[687] = 1'b1;
    assign layer1_outputs[688] = ~(layer0_outputs[6089]);
    assign layer1_outputs[689] = (layer0_outputs[10218]) & (layer0_outputs[3861]);
    assign layer1_outputs[690] = ~(layer0_outputs[9850]);
    assign layer1_outputs[691] = layer0_outputs[6771];
    assign layer1_outputs[692] = layer0_outputs[9949];
    assign layer1_outputs[693] = ~(layer0_outputs[12775]) | (layer0_outputs[6877]);
    assign layer1_outputs[694] = (layer0_outputs[12589]) ^ (layer0_outputs[513]);
    assign layer1_outputs[695] = ~(layer0_outputs[10933]);
    assign layer1_outputs[696] = (layer0_outputs[5137]) ^ (layer0_outputs[868]);
    assign layer1_outputs[697] = ~(layer0_outputs[12756]) | (layer0_outputs[8197]);
    assign layer1_outputs[698] = (layer0_outputs[3968]) ^ (layer0_outputs[8739]);
    assign layer1_outputs[699] = (layer0_outputs[11713]) & ~(layer0_outputs[8088]);
    assign layer1_outputs[700] = layer0_outputs[7566];
    assign layer1_outputs[701] = ~(layer0_outputs[2488]);
    assign layer1_outputs[702] = layer0_outputs[3054];
    assign layer1_outputs[703] = ~(layer0_outputs[6661]) | (layer0_outputs[7538]);
    assign layer1_outputs[704] = (layer0_outputs[322]) & ~(layer0_outputs[7135]);
    assign layer1_outputs[705] = ~(layer0_outputs[1986]);
    assign layer1_outputs[706] = ~(layer0_outputs[11318]);
    assign layer1_outputs[707] = layer0_outputs[3311];
    assign layer1_outputs[708] = (layer0_outputs[3614]) & ~(layer0_outputs[8616]);
    assign layer1_outputs[709] = ~(layer0_outputs[1913]) | (layer0_outputs[9590]);
    assign layer1_outputs[710] = ~(layer0_outputs[5628]);
    assign layer1_outputs[711] = layer0_outputs[6750];
    assign layer1_outputs[712] = ~(layer0_outputs[9523]);
    assign layer1_outputs[713] = ~(layer0_outputs[11131]);
    assign layer1_outputs[714] = ~(layer0_outputs[5053]);
    assign layer1_outputs[715] = (layer0_outputs[7203]) | (layer0_outputs[11905]);
    assign layer1_outputs[716] = ~((layer0_outputs[716]) & (layer0_outputs[7801]));
    assign layer1_outputs[717] = (layer0_outputs[3809]) & ~(layer0_outputs[12302]);
    assign layer1_outputs[718] = (layer0_outputs[10432]) & (layer0_outputs[925]);
    assign layer1_outputs[719] = (layer0_outputs[652]) & (layer0_outputs[5845]);
    assign layer1_outputs[720] = (layer0_outputs[7017]) & ~(layer0_outputs[6492]);
    assign layer1_outputs[721] = ~(layer0_outputs[2311]);
    assign layer1_outputs[722] = layer0_outputs[5557];
    assign layer1_outputs[723] = ~(layer0_outputs[4777]);
    assign layer1_outputs[724] = layer0_outputs[2856];
    assign layer1_outputs[725] = ~((layer0_outputs[5191]) & (layer0_outputs[2219]));
    assign layer1_outputs[726] = ~(layer0_outputs[12625]);
    assign layer1_outputs[727] = layer0_outputs[3176];
    assign layer1_outputs[728] = (layer0_outputs[2883]) & ~(layer0_outputs[9907]);
    assign layer1_outputs[729] = ~((layer0_outputs[998]) & (layer0_outputs[2986]));
    assign layer1_outputs[730] = ~((layer0_outputs[10028]) & (layer0_outputs[7798]));
    assign layer1_outputs[731] = layer0_outputs[4563];
    assign layer1_outputs[732] = ~((layer0_outputs[4651]) & (layer0_outputs[3935]));
    assign layer1_outputs[733] = ~(layer0_outputs[5501]);
    assign layer1_outputs[734] = 1'b0;
    assign layer1_outputs[735] = (layer0_outputs[5495]) & ~(layer0_outputs[5303]);
    assign layer1_outputs[736] = layer0_outputs[7386];
    assign layer1_outputs[737] = (layer0_outputs[5049]) | (layer0_outputs[6677]);
    assign layer1_outputs[738] = (layer0_outputs[4829]) & ~(layer0_outputs[12041]);
    assign layer1_outputs[739] = layer0_outputs[4824];
    assign layer1_outputs[740] = ~(layer0_outputs[7168]) | (layer0_outputs[698]);
    assign layer1_outputs[741] = 1'b1;
    assign layer1_outputs[742] = ~(layer0_outputs[2445]) | (layer0_outputs[74]);
    assign layer1_outputs[743] = (layer0_outputs[6334]) & ~(layer0_outputs[9533]);
    assign layer1_outputs[744] = ~(layer0_outputs[7292]) | (layer0_outputs[12619]);
    assign layer1_outputs[745] = layer0_outputs[287];
    assign layer1_outputs[746] = ~(layer0_outputs[2468]) | (layer0_outputs[9219]);
    assign layer1_outputs[747] = (layer0_outputs[3890]) ^ (layer0_outputs[8502]);
    assign layer1_outputs[748] = ~(layer0_outputs[6574]);
    assign layer1_outputs[749] = (layer0_outputs[1377]) ^ (layer0_outputs[2876]);
    assign layer1_outputs[750] = ~((layer0_outputs[8485]) | (layer0_outputs[8710]));
    assign layer1_outputs[751] = ~(layer0_outputs[635]);
    assign layer1_outputs[752] = ~(layer0_outputs[6881]) | (layer0_outputs[8812]);
    assign layer1_outputs[753] = (layer0_outputs[5060]) | (layer0_outputs[10485]);
    assign layer1_outputs[754] = ~(layer0_outputs[3660]) | (layer0_outputs[6129]);
    assign layer1_outputs[755] = ~(layer0_outputs[4888]);
    assign layer1_outputs[756] = ~(layer0_outputs[1702]);
    assign layer1_outputs[757] = ~(layer0_outputs[3318]);
    assign layer1_outputs[758] = ~((layer0_outputs[1713]) & (layer0_outputs[98]));
    assign layer1_outputs[759] = layer0_outputs[1971];
    assign layer1_outputs[760] = (layer0_outputs[12010]) & (layer0_outputs[10977]);
    assign layer1_outputs[761] = (layer0_outputs[8377]) & ~(layer0_outputs[8760]);
    assign layer1_outputs[762] = (layer0_outputs[4262]) & ~(layer0_outputs[5921]);
    assign layer1_outputs[763] = ~(layer0_outputs[10065]) | (layer0_outputs[3555]);
    assign layer1_outputs[764] = (layer0_outputs[6119]) ^ (layer0_outputs[8590]);
    assign layer1_outputs[765] = ~(layer0_outputs[2186]) | (layer0_outputs[10121]);
    assign layer1_outputs[766] = (layer0_outputs[10818]) ^ (layer0_outputs[4311]);
    assign layer1_outputs[767] = ~((layer0_outputs[10185]) | (layer0_outputs[11919]));
    assign layer1_outputs[768] = (layer0_outputs[360]) & ~(layer0_outputs[4533]);
    assign layer1_outputs[769] = layer0_outputs[6058];
    assign layer1_outputs[770] = ~((layer0_outputs[5629]) ^ (layer0_outputs[10617]));
    assign layer1_outputs[771] = ~(layer0_outputs[3385]);
    assign layer1_outputs[772] = ~(layer0_outputs[2629]) | (layer0_outputs[3257]);
    assign layer1_outputs[773] = ~(layer0_outputs[2726]);
    assign layer1_outputs[774] = layer0_outputs[1637];
    assign layer1_outputs[775] = (layer0_outputs[5515]) & (layer0_outputs[6245]);
    assign layer1_outputs[776] = ~((layer0_outputs[6527]) | (layer0_outputs[8334]));
    assign layer1_outputs[777] = layer0_outputs[7848];
    assign layer1_outputs[778] = layer0_outputs[12615];
    assign layer1_outputs[779] = (layer0_outputs[5664]) & ~(layer0_outputs[10523]);
    assign layer1_outputs[780] = (layer0_outputs[1045]) | (layer0_outputs[10277]);
    assign layer1_outputs[781] = ~((layer0_outputs[6228]) ^ (layer0_outputs[8597]));
    assign layer1_outputs[782] = layer0_outputs[2803];
    assign layer1_outputs[783] = ~(layer0_outputs[5366]) | (layer0_outputs[8985]);
    assign layer1_outputs[784] = layer0_outputs[2563];
    assign layer1_outputs[785] = layer0_outputs[3443];
    assign layer1_outputs[786] = (layer0_outputs[4971]) ^ (layer0_outputs[2651]);
    assign layer1_outputs[787] = ~(layer0_outputs[1153]);
    assign layer1_outputs[788] = layer0_outputs[12211];
    assign layer1_outputs[789] = ~(layer0_outputs[12008]);
    assign layer1_outputs[790] = (layer0_outputs[3293]) ^ (layer0_outputs[3631]);
    assign layer1_outputs[791] = ~(layer0_outputs[7266]);
    assign layer1_outputs[792] = (layer0_outputs[3165]) ^ (layer0_outputs[3047]);
    assign layer1_outputs[793] = (layer0_outputs[7740]) & ~(layer0_outputs[2172]);
    assign layer1_outputs[794] = ~((layer0_outputs[10182]) | (layer0_outputs[6793]));
    assign layer1_outputs[795] = ~((layer0_outputs[7682]) | (layer0_outputs[2497]));
    assign layer1_outputs[796] = layer0_outputs[10227];
    assign layer1_outputs[797] = layer0_outputs[11057];
    assign layer1_outputs[798] = layer0_outputs[5269];
    assign layer1_outputs[799] = ~(layer0_outputs[12656]) | (layer0_outputs[10315]);
    assign layer1_outputs[800] = (layer0_outputs[10119]) & ~(layer0_outputs[8384]);
    assign layer1_outputs[801] = layer0_outputs[6054];
    assign layer1_outputs[802] = layer0_outputs[12601];
    assign layer1_outputs[803] = ~(layer0_outputs[2369]) | (layer0_outputs[6160]);
    assign layer1_outputs[804] = ~((layer0_outputs[7529]) | (layer0_outputs[6964]));
    assign layer1_outputs[805] = (layer0_outputs[1030]) & ~(layer0_outputs[1628]);
    assign layer1_outputs[806] = (layer0_outputs[9175]) & (layer0_outputs[8220]);
    assign layer1_outputs[807] = ~(layer0_outputs[12637]);
    assign layer1_outputs[808] = layer0_outputs[9105];
    assign layer1_outputs[809] = ~((layer0_outputs[2848]) | (layer0_outputs[364]));
    assign layer1_outputs[810] = layer0_outputs[1761];
    assign layer1_outputs[811] = layer0_outputs[10958];
    assign layer1_outputs[812] = ~(layer0_outputs[6710]);
    assign layer1_outputs[813] = ~(layer0_outputs[5595]) | (layer0_outputs[3775]);
    assign layer1_outputs[814] = (layer0_outputs[6404]) & ~(layer0_outputs[1605]);
    assign layer1_outputs[815] = ~(layer0_outputs[390]);
    assign layer1_outputs[816] = layer0_outputs[9243];
    assign layer1_outputs[817] = (layer0_outputs[2096]) & (layer0_outputs[3513]);
    assign layer1_outputs[818] = 1'b0;
    assign layer1_outputs[819] = ~(layer0_outputs[1054]);
    assign layer1_outputs[820] = (layer0_outputs[1701]) ^ (layer0_outputs[8966]);
    assign layer1_outputs[821] = ~((layer0_outputs[218]) ^ (layer0_outputs[5607]));
    assign layer1_outputs[822] = ~((layer0_outputs[8825]) ^ (layer0_outputs[5272]));
    assign layer1_outputs[823] = layer0_outputs[7617];
    assign layer1_outputs[824] = ~(layer0_outputs[6580]);
    assign layer1_outputs[825] = ~((layer0_outputs[5199]) & (layer0_outputs[10555]));
    assign layer1_outputs[826] = layer0_outputs[8088];
    assign layer1_outputs[827] = ~(layer0_outputs[4994]);
    assign layer1_outputs[828] = ~((layer0_outputs[10559]) | (layer0_outputs[1856]));
    assign layer1_outputs[829] = (layer0_outputs[9114]) & (layer0_outputs[1454]);
    assign layer1_outputs[830] = (layer0_outputs[4176]) & ~(layer0_outputs[4328]);
    assign layer1_outputs[831] = layer0_outputs[123];
    assign layer1_outputs[832] = ~(layer0_outputs[7815]) | (layer0_outputs[2416]);
    assign layer1_outputs[833] = layer0_outputs[10377];
    assign layer1_outputs[834] = (layer0_outputs[1158]) ^ (layer0_outputs[10868]);
    assign layer1_outputs[835] = layer0_outputs[12410];
    assign layer1_outputs[836] = ~(layer0_outputs[7517]);
    assign layer1_outputs[837] = ~(layer0_outputs[2827]);
    assign layer1_outputs[838] = ~(layer0_outputs[10026]) | (layer0_outputs[5720]);
    assign layer1_outputs[839] = ~(layer0_outputs[6788]) | (layer0_outputs[9394]);
    assign layer1_outputs[840] = ~((layer0_outputs[6495]) | (layer0_outputs[5646]));
    assign layer1_outputs[841] = layer0_outputs[5904];
    assign layer1_outputs[842] = ~(layer0_outputs[12433]);
    assign layer1_outputs[843] = ~(layer0_outputs[7284]) | (layer0_outputs[1427]);
    assign layer1_outputs[844] = layer0_outputs[10173];
    assign layer1_outputs[845] = (layer0_outputs[11421]) & (layer0_outputs[10753]);
    assign layer1_outputs[846] = ~((layer0_outputs[2114]) ^ (layer0_outputs[5342]));
    assign layer1_outputs[847] = layer0_outputs[3489];
    assign layer1_outputs[848] = ~(layer0_outputs[3724]);
    assign layer1_outputs[849] = (layer0_outputs[3362]) & ~(layer0_outputs[5893]);
    assign layer1_outputs[850] = 1'b1;
    assign layer1_outputs[851] = ~(layer0_outputs[7900]);
    assign layer1_outputs[852] = ~(layer0_outputs[8957]);
    assign layer1_outputs[853] = ~(layer0_outputs[8520]) | (layer0_outputs[4894]);
    assign layer1_outputs[854] = (layer0_outputs[8304]) & ~(layer0_outputs[1890]);
    assign layer1_outputs[855] = ~(layer0_outputs[1800]);
    assign layer1_outputs[856] = ~(layer0_outputs[7092]);
    assign layer1_outputs[857] = (layer0_outputs[5863]) ^ (layer0_outputs[8516]);
    assign layer1_outputs[858] = layer0_outputs[11737];
    assign layer1_outputs[859] = ~(layer0_outputs[10653]);
    assign layer1_outputs[860] = ~((layer0_outputs[7213]) | (layer0_outputs[1068]));
    assign layer1_outputs[861] = ~(layer0_outputs[8344]);
    assign layer1_outputs[862] = (layer0_outputs[8647]) | (layer0_outputs[8493]);
    assign layer1_outputs[863] = ~(layer0_outputs[487]);
    assign layer1_outputs[864] = layer0_outputs[4685];
    assign layer1_outputs[865] = ~(layer0_outputs[12355]);
    assign layer1_outputs[866] = layer0_outputs[11495];
    assign layer1_outputs[867] = layer0_outputs[12218];
    assign layer1_outputs[868] = ~(layer0_outputs[185]) | (layer0_outputs[2025]);
    assign layer1_outputs[869] = ~(layer0_outputs[2066]);
    assign layer1_outputs[870] = layer0_outputs[3082];
    assign layer1_outputs[871] = ~((layer0_outputs[1009]) & (layer0_outputs[2608]));
    assign layer1_outputs[872] = ~(layer0_outputs[6680]) | (layer0_outputs[5981]);
    assign layer1_outputs[873] = layer0_outputs[10245];
    assign layer1_outputs[874] = layer0_outputs[11781];
    assign layer1_outputs[875] = ~((layer0_outputs[62]) | (layer0_outputs[6307]));
    assign layer1_outputs[876] = layer0_outputs[11587];
    assign layer1_outputs[877] = (layer0_outputs[4090]) | (layer0_outputs[3637]);
    assign layer1_outputs[878] = (layer0_outputs[5345]) ^ (layer0_outputs[2704]);
    assign layer1_outputs[879] = layer0_outputs[8649];
    assign layer1_outputs[880] = ~(layer0_outputs[1412]);
    assign layer1_outputs[881] = layer0_outputs[3105];
    assign layer1_outputs[882] = layer0_outputs[12727];
    assign layer1_outputs[883] = ~((layer0_outputs[8675]) & (layer0_outputs[5173]));
    assign layer1_outputs[884] = layer0_outputs[6791];
    assign layer1_outputs[885] = layer0_outputs[6225];
    assign layer1_outputs[886] = ~(layer0_outputs[6622]);
    assign layer1_outputs[887] = ~(layer0_outputs[11522]);
    assign layer1_outputs[888] = ~((layer0_outputs[993]) | (layer0_outputs[1361]));
    assign layer1_outputs[889] = ~((layer0_outputs[10207]) ^ (layer0_outputs[4688]));
    assign layer1_outputs[890] = (layer0_outputs[7105]) & (layer0_outputs[17]);
    assign layer1_outputs[891] = ~(layer0_outputs[3634]);
    assign layer1_outputs[892] = ~(layer0_outputs[7978]);
    assign layer1_outputs[893] = (layer0_outputs[10882]) & ~(layer0_outputs[6966]);
    assign layer1_outputs[894] = ~(layer0_outputs[11409]);
    assign layer1_outputs[895] = layer0_outputs[5025];
    assign layer1_outputs[896] = ~((layer0_outputs[10862]) ^ (layer0_outputs[12306]));
    assign layer1_outputs[897] = (layer0_outputs[7420]) | (layer0_outputs[2116]);
    assign layer1_outputs[898] = layer0_outputs[887];
    assign layer1_outputs[899] = ~((layer0_outputs[12254]) | (layer0_outputs[9291]));
    assign layer1_outputs[900] = ~((layer0_outputs[11471]) ^ (layer0_outputs[5836]));
    assign layer1_outputs[901] = (layer0_outputs[10901]) ^ (layer0_outputs[790]);
    assign layer1_outputs[902] = ~((layer0_outputs[12264]) | (layer0_outputs[1810]));
    assign layer1_outputs[903] = ~(layer0_outputs[4948]);
    assign layer1_outputs[904] = (layer0_outputs[7340]) | (layer0_outputs[5148]);
    assign layer1_outputs[905] = (layer0_outputs[1520]) & ~(layer0_outputs[4933]);
    assign layer1_outputs[906] = ~(layer0_outputs[5626]);
    assign layer1_outputs[907] = (layer0_outputs[612]) & (layer0_outputs[2291]);
    assign layer1_outputs[908] = (layer0_outputs[398]) ^ (layer0_outputs[7761]);
    assign layer1_outputs[909] = (layer0_outputs[1666]) | (layer0_outputs[5196]);
    assign layer1_outputs[910] = layer0_outputs[3316];
    assign layer1_outputs[911] = (layer0_outputs[4157]) | (layer0_outputs[9789]);
    assign layer1_outputs[912] = ~((layer0_outputs[3954]) ^ (layer0_outputs[9451]));
    assign layer1_outputs[913] = ~(layer0_outputs[8472]);
    assign layer1_outputs[914] = layer0_outputs[8831];
    assign layer1_outputs[915] = (layer0_outputs[12564]) & ~(layer0_outputs[8114]);
    assign layer1_outputs[916] = (layer0_outputs[8900]) & ~(layer0_outputs[12446]);
    assign layer1_outputs[917] = ~((layer0_outputs[9549]) & (layer0_outputs[5301]));
    assign layer1_outputs[918] = (layer0_outputs[4660]) & ~(layer0_outputs[6364]);
    assign layer1_outputs[919] = (layer0_outputs[5638]) & ~(layer0_outputs[12335]);
    assign layer1_outputs[920] = ~(layer0_outputs[10130]) | (layer0_outputs[9789]);
    assign layer1_outputs[921] = (layer0_outputs[5759]) | (layer0_outputs[9748]);
    assign layer1_outputs[922] = layer0_outputs[5333];
    assign layer1_outputs[923] = ~(layer0_outputs[8204]) | (layer0_outputs[9129]);
    assign layer1_outputs[924] = layer0_outputs[5814];
    assign layer1_outputs[925] = (layer0_outputs[8312]) & ~(layer0_outputs[3012]);
    assign layer1_outputs[926] = (layer0_outputs[6041]) & ~(layer0_outputs[7637]);
    assign layer1_outputs[927] = layer0_outputs[4900];
    assign layer1_outputs[928] = ~((layer0_outputs[6212]) & (layer0_outputs[6654]));
    assign layer1_outputs[929] = (layer0_outputs[8202]) & ~(layer0_outputs[5686]);
    assign layer1_outputs[930] = layer0_outputs[11229];
    assign layer1_outputs[931] = layer0_outputs[10613];
    assign layer1_outputs[932] = (layer0_outputs[6449]) & ~(layer0_outputs[1819]);
    assign layer1_outputs[933] = ~((layer0_outputs[11185]) | (layer0_outputs[11395]));
    assign layer1_outputs[934] = ~(layer0_outputs[12492]) | (layer0_outputs[6549]);
    assign layer1_outputs[935] = layer0_outputs[8667];
    assign layer1_outputs[936] = ~((layer0_outputs[2809]) & (layer0_outputs[4718]));
    assign layer1_outputs[937] = ~(layer0_outputs[4076]);
    assign layer1_outputs[938] = ~((layer0_outputs[11410]) ^ (layer0_outputs[11633]));
    assign layer1_outputs[939] = layer0_outputs[1583];
    assign layer1_outputs[940] = (layer0_outputs[882]) | (layer0_outputs[897]);
    assign layer1_outputs[941] = ~(layer0_outputs[7278]) | (layer0_outputs[8203]);
    assign layer1_outputs[942] = ~((layer0_outputs[6887]) ^ (layer0_outputs[11376]));
    assign layer1_outputs[943] = ~(layer0_outputs[2188]);
    assign layer1_outputs[944] = ~((layer0_outputs[5687]) | (layer0_outputs[7893]));
    assign layer1_outputs[945] = ~(layer0_outputs[9128]);
    assign layer1_outputs[946] = layer0_outputs[5804];
    assign layer1_outputs[947] = layer0_outputs[2365];
    assign layer1_outputs[948] = ~(layer0_outputs[9841]);
    assign layer1_outputs[949] = ~(layer0_outputs[12679]);
    assign layer1_outputs[950] = (layer0_outputs[4836]) | (layer0_outputs[7817]);
    assign layer1_outputs[951] = ~((layer0_outputs[8581]) & (layer0_outputs[1364]));
    assign layer1_outputs[952] = layer0_outputs[3254];
    assign layer1_outputs[953] = (layer0_outputs[8270]) | (layer0_outputs[12685]);
    assign layer1_outputs[954] = ~(layer0_outputs[929]);
    assign layer1_outputs[955] = layer0_outputs[5932];
    assign layer1_outputs[956] = (layer0_outputs[1172]) & ~(layer0_outputs[11912]);
    assign layer1_outputs[957] = (layer0_outputs[3792]) | (layer0_outputs[4861]);
    assign layer1_outputs[958] = (layer0_outputs[7419]) & ~(layer0_outputs[7776]);
    assign layer1_outputs[959] = 1'b0;
    assign layer1_outputs[960] = (layer0_outputs[7209]) & ~(layer0_outputs[11394]);
    assign layer1_outputs[961] = (layer0_outputs[5289]) & ~(layer0_outputs[12678]);
    assign layer1_outputs[962] = ~(layer0_outputs[5480]) | (layer0_outputs[11611]);
    assign layer1_outputs[963] = (layer0_outputs[7783]) | (layer0_outputs[7655]);
    assign layer1_outputs[964] = ~(layer0_outputs[9630]);
    assign layer1_outputs[965] = (layer0_outputs[6703]) | (layer0_outputs[7155]);
    assign layer1_outputs[966] = layer0_outputs[8163];
    assign layer1_outputs[967] = (layer0_outputs[9578]) | (layer0_outputs[879]);
    assign layer1_outputs[968] = (layer0_outputs[7417]) | (layer0_outputs[12598]);
    assign layer1_outputs[969] = ~(layer0_outputs[9870]);
    assign layer1_outputs[970] = (layer0_outputs[11256]) & ~(layer0_outputs[6899]);
    assign layer1_outputs[971] = 1'b1;
    assign layer1_outputs[972] = ~(layer0_outputs[12412]);
    assign layer1_outputs[973] = (layer0_outputs[8330]) & ~(layer0_outputs[11183]);
    assign layer1_outputs[974] = ~(layer0_outputs[1987]) | (layer0_outputs[8679]);
    assign layer1_outputs[975] = (layer0_outputs[1611]) | (layer0_outputs[11996]);
    assign layer1_outputs[976] = (layer0_outputs[1163]) & ~(layer0_outputs[9799]);
    assign layer1_outputs[977] = layer0_outputs[10701];
    assign layer1_outputs[978] = (layer0_outputs[3696]) & ~(layer0_outputs[9304]);
    assign layer1_outputs[979] = ~((layer0_outputs[11132]) ^ (layer0_outputs[2508]));
    assign layer1_outputs[980] = ~(layer0_outputs[11259]) | (layer0_outputs[3417]);
    assign layer1_outputs[981] = layer0_outputs[1902];
    assign layer1_outputs[982] = (layer0_outputs[2836]) & ~(layer0_outputs[4457]);
    assign layer1_outputs[983] = ~(layer0_outputs[6857]);
    assign layer1_outputs[984] = ~(layer0_outputs[6869]);
    assign layer1_outputs[985] = layer0_outputs[5011];
    assign layer1_outputs[986] = (layer0_outputs[6844]) ^ (layer0_outputs[12222]);
    assign layer1_outputs[987] = ~(layer0_outputs[2414]) | (layer0_outputs[5250]);
    assign layer1_outputs[988] = (layer0_outputs[8251]) & ~(layer0_outputs[1946]);
    assign layer1_outputs[989] = (layer0_outputs[2957]) & (layer0_outputs[12366]);
    assign layer1_outputs[990] = (layer0_outputs[4919]) & (layer0_outputs[3349]);
    assign layer1_outputs[991] = (layer0_outputs[8026]) ^ (layer0_outputs[4801]);
    assign layer1_outputs[992] = ~(layer0_outputs[5614]) | (layer0_outputs[6619]);
    assign layer1_outputs[993] = 1'b1;
    assign layer1_outputs[994] = (layer0_outputs[11743]) & ~(layer0_outputs[1582]);
    assign layer1_outputs[995] = ~(layer0_outputs[1499]) | (layer0_outputs[6182]);
    assign layer1_outputs[996] = ~((layer0_outputs[2514]) | (layer0_outputs[5110]));
    assign layer1_outputs[997] = ~(layer0_outputs[7811]);
    assign layer1_outputs[998] = layer0_outputs[2274];
    assign layer1_outputs[999] = layer0_outputs[1504];
    assign layer1_outputs[1000] = 1'b0;
    assign layer1_outputs[1001] = ~(layer0_outputs[793]) | (layer0_outputs[6888]);
    assign layer1_outputs[1002] = (layer0_outputs[11444]) ^ (layer0_outputs[3141]);
    assign layer1_outputs[1003] = (layer0_outputs[2352]) & ~(layer0_outputs[11148]);
    assign layer1_outputs[1004] = ~((layer0_outputs[2622]) ^ (layer0_outputs[4122]));
    assign layer1_outputs[1005] = (layer0_outputs[3942]) & (layer0_outputs[12252]);
    assign layer1_outputs[1006] = ~(layer0_outputs[8621]) | (layer0_outputs[4795]);
    assign layer1_outputs[1007] = (layer0_outputs[7647]) & (layer0_outputs[3999]);
    assign layer1_outputs[1008] = (layer0_outputs[7461]) & ~(layer0_outputs[4385]);
    assign layer1_outputs[1009] = layer0_outputs[6634];
    assign layer1_outputs[1010] = ~(layer0_outputs[11017]);
    assign layer1_outputs[1011] = layer0_outputs[2837];
    assign layer1_outputs[1012] = ~(layer0_outputs[7550]) | (layer0_outputs[9890]);
    assign layer1_outputs[1013] = layer0_outputs[12499];
    assign layer1_outputs[1014] = (layer0_outputs[5456]) & ~(layer0_outputs[7654]);
    assign layer1_outputs[1015] = ~(layer0_outputs[8744]) | (layer0_outputs[8623]);
    assign layer1_outputs[1016] = ~((layer0_outputs[10488]) | (layer0_outputs[6231]));
    assign layer1_outputs[1017] = (layer0_outputs[7991]) & (layer0_outputs[878]);
    assign layer1_outputs[1018] = ~(layer0_outputs[1320]);
    assign layer1_outputs[1019] = (layer0_outputs[9619]) | (layer0_outputs[5734]);
    assign layer1_outputs[1020] = (layer0_outputs[4371]) | (layer0_outputs[7512]);
    assign layer1_outputs[1021] = (layer0_outputs[5315]) & ~(layer0_outputs[2935]);
    assign layer1_outputs[1022] = ~(layer0_outputs[2452]);
    assign layer1_outputs[1023] = ~(layer0_outputs[11545]) | (layer0_outputs[6438]);
    assign layer1_outputs[1024] = ~((layer0_outputs[1362]) ^ (layer0_outputs[6027]));
    assign layer1_outputs[1025] = layer0_outputs[10810];
    assign layer1_outputs[1026] = layer0_outputs[1781];
    assign layer1_outputs[1027] = layer0_outputs[11974];
    assign layer1_outputs[1028] = ~(layer0_outputs[12375]);
    assign layer1_outputs[1029] = (layer0_outputs[3011]) & (layer0_outputs[12237]);
    assign layer1_outputs[1030] = ~(layer0_outputs[952]);
    assign layer1_outputs[1031] = ~(layer0_outputs[1363]) | (layer0_outputs[9067]);
    assign layer1_outputs[1032] = (layer0_outputs[1774]) ^ (layer0_outputs[2167]);
    assign layer1_outputs[1033] = ~((layer0_outputs[9161]) | (layer0_outputs[9123]));
    assign layer1_outputs[1034] = ~(layer0_outputs[12289]);
    assign layer1_outputs[1035] = (layer0_outputs[12532]) ^ (layer0_outputs[7660]);
    assign layer1_outputs[1036] = (layer0_outputs[1209]) & (layer0_outputs[445]);
    assign layer1_outputs[1037] = layer0_outputs[10948];
    assign layer1_outputs[1038] = ~(layer0_outputs[6696]);
    assign layer1_outputs[1039] = (layer0_outputs[4043]) | (layer0_outputs[2909]);
    assign layer1_outputs[1040] = layer0_outputs[2423];
    assign layer1_outputs[1041] = ~((layer0_outputs[4236]) ^ (layer0_outputs[6005]));
    assign layer1_outputs[1042] = ~(layer0_outputs[4830]) | (layer0_outputs[7660]);
    assign layer1_outputs[1043] = ~(layer0_outputs[11742]) | (layer0_outputs[1445]);
    assign layer1_outputs[1044] = ~(layer0_outputs[11029]);
    assign layer1_outputs[1045] = ~(layer0_outputs[5054]);
    assign layer1_outputs[1046] = layer0_outputs[226];
    assign layer1_outputs[1047] = ~((layer0_outputs[3230]) & (layer0_outputs[12141]));
    assign layer1_outputs[1048] = ~(layer0_outputs[11019]) | (layer0_outputs[9389]);
    assign layer1_outputs[1049] = layer0_outputs[11067];
    assign layer1_outputs[1050] = ~((layer0_outputs[2990]) & (layer0_outputs[4729]));
    assign layer1_outputs[1051] = (layer0_outputs[532]) ^ (layer0_outputs[7636]);
    assign layer1_outputs[1052] = layer0_outputs[3781];
    assign layer1_outputs[1053] = layer0_outputs[4994];
    assign layer1_outputs[1054] = ~((layer0_outputs[7682]) | (layer0_outputs[11381]));
    assign layer1_outputs[1055] = 1'b1;
    assign layer1_outputs[1056] = layer0_outputs[7326];
    assign layer1_outputs[1057] = (layer0_outputs[5708]) & ~(layer0_outputs[9320]);
    assign layer1_outputs[1058] = ~(layer0_outputs[10103]) | (layer0_outputs[853]);
    assign layer1_outputs[1059] = ~(layer0_outputs[11140]);
    assign layer1_outputs[1060] = (layer0_outputs[2577]) & ~(layer0_outputs[8019]);
    assign layer1_outputs[1061] = layer0_outputs[12070];
    assign layer1_outputs[1062] = (layer0_outputs[6400]) & ~(layer0_outputs[9556]);
    assign layer1_outputs[1063] = layer0_outputs[9919];
    assign layer1_outputs[1064] = layer0_outputs[1088];
    assign layer1_outputs[1065] = (layer0_outputs[3428]) & ~(layer0_outputs[4690]);
    assign layer1_outputs[1066] = ~(layer0_outputs[10382]) | (layer0_outputs[10881]);
    assign layer1_outputs[1067] = ~(layer0_outputs[5933]) | (layer0_outputs[4864]);
    assign layer1_outputs[1068] = layer0_outputs[2605];
    assign layer1_outputs[1069] = layer0_outputs[7255];
    assign layer1_outputs[1070] = (layer0_outputs[8684]) & ~(layer0_outputs[1610]);
    assign layer1_outputs[1071] = ~(layer0_outputs[8032]) | (layer0_outputs[1113]);
    assign layer1_outputs[1072] = ~(layer0_outputs[12616]) | (layer0_outputs[3238]);
    assign layer1_outputs[1073] = layer0_outputs[9489];
    assign layer1_outputs[1074] = layer0_outputs[9348];
    assign layer1_outputs[1075] = layer0_outputs[395];
    assign layer1_outputs[1076] = layer0_outputs[3383];
    assign layer1_outputs[1077] = layer0_outputs[11315];
    assign layer1_outputs[1078] = (layer0_outputs[505]) ^ (layer0_outputs[12691]);
    assign layer1_outputs[1079] = ~(layer0_outputs[4310]);
    assign layer1_outputs[1080] = ~((layer0_outputs[9109]) ^ (layer0_outputs[6461]));
    assign layer1_outputs[1081] = (layer0_outputs[5263]) & ~(layer0_outputs[9412]);
    assign layer1_outputs[1082] = ~((layer0_outputs[8111]) ^ (layer0_outputs[6666]));
    assign layer1_outputs[1083] = ~(layer0_outputs[4458]) | (layer0_outputs[8916]);
    assign layer1_outputs[1084] = ~((layer0_outputs[2330]) | (layer0_outputs[3679]));
    assign layer1_outputs[1085] = (layer0_outputs[4849]) & (layer0_outputs[12670]);
    assign layer1_outputs[1086] = (layer0_outputs[3231]) ^ (layer0_outputs[11768]);
    assign layer1_outputs[1087] = ~(layer0_outputs[5553]);
    assign layer1_outputs[1088] = ~((layer0_outputs[941]) | (layer0_outputs[6106]));
    assign layer1_outputs[1089] = (layer0_outputs[4001]) ^ (layer0_outputs[11512]);
    assign layer1_outputs[1090] = ~(layer0_outputs[1298]);
    assign layer1_outputs[1091] = ~((layer0_outputs[4667]) | (layer0_outputs[9221]));
    assign layer1_outputs[1092] = ~((layer0_outputs[10305]) & (layer0_outputs[2686]));
    assign layer1_outputs[1093] = ~(layer0_outputs[10767]);
    assign layer1_outputs[1094] = ~(layer0_outputs[3460]);
    assign layer1_outputs[1095] = (layer0_outputs[6142]) & ~(layer0_outputs[2194]);
    assign layer1_outputs[1096] = ~((layer0_outputs[6867]) ^ (layer0_outputs[10516]));
    assign layer1_outputs[1097] = ~(layer0_outputs[3142]);
    assign layer1_outputs[1098] = (layer0_outputs[948]) & ~(layer0_outputs[12159]);
    assign layer1_outputs[1099] = layer0_outputs[5236];
    assign layer1_outputs[1100] = ~(layer0_outputs[11480]);
    assign layer1_outputs[1101] = (layer0_outputs[6260]) | (layer0_outputs[8008]);
    assign layer1_outputs[1102] = (layer0_outputs[6428]) & ~(layer0_outputs[5804]);
    assign layer1_outputs[1103] = layer0_outputs[3113];
    assign layer1_outputs[1104] = (layer0_outputs[353]) & ~(layer0_outputs[6548]);
    assign layer1_outputs[1105] = ~(layer0_outputs[2382]);
    assign layer1_outputs[1106] = ~(layer0_outputs[10841]) | (layer0_outputs[4252]);
    assign layer1_outputs[1107] = (layer0_outputs[6826]) ^ (layer0_outputs[7083]);
    assign layer1_outputs[1108] = (layer0_outputs[6133]) & (layer0_outputs[7184]);
    assign layer1_outputs[1109] = ~(layer0_outputs[3496]);
    assign layer1_outputs[1110] = (layer0_outputs[7853]) & ~(layer0_outputs[10196]);
    assign layer1_outputs[1111] = ~((layer0_outputs[12330]) ^ (layer0_outputs[8046]));
    assign layer1_outputs[1112] = ~(layer0_outputs[5371]);
    assign layer1_outputs[1113] = layer0_outputs[7762];
    assign layer1_outputs[1114] = (layer0_outputs[2923]) | (layer0_outputs[12184]);
    assign layer1_outputs[1115] = (layer0_outputs[12376]) ^ (layer0_outputs[1752]);
    assign layer1_outputs[1116] = ~((layer0_outputs[8477]) & (layer0_outputs[1386]));
    assign layer1_outputs[1117] = (layer0_outputs[5527]) ^ (layer0_outputs[9866]);
    assign layer1_outputs[1118] = layer0_outputs[3339];
    assign layer1_outputs[1119] = (layer0_outputs[1240]) ^ (layer0_outputs[3031]);
    assign layer1_outputs[1120] = ~(layer0_outputs[11014]);
    assign layer1_outputs[1121] = ~((layer0_outputs[4136]) & (layer0_outputs[4791]));
    assign layer1_outputs[1122] = layer0_outputs[4356];
    assign layer1_outputs[1123] = (layer0_outputs[11568]) & ~(layer0_outputs[10962]);
    assign layer1_outputs[1124] = (layer0_outputs[11012]) ^ (layer0_outputs[11245]);
    assign layer1_outputs[1125] = ~((layer0_outputs[7866]) & (layer0_outputs[7230]));
    assign layer1_outputs[1126] = layer0_outputs[2605];
    assign layer1_outputs[1127] = layer0_outputs[5091];
    assign layer1_outputs[1128] = ~(layer0_outputs[2247]);
    assign layer1_outputs[1129] = ~(layer0_outputs[5990]);
    assign layer1_outputs[1130] = (layer0_outputs[666]) & ~(layer0_outputs[8338]);
    assign layer1_outputs[1131] = layer0_outputs[8984];
    assign layer1_outputs[1132] = ~(layer0_outputs[12739]) | (layer0_outputs[6570]);
    assign layer1_outputs[1133] = ~(layer0_outputs[12363]);
    assign layer1_outputs[1134] = layer0_outputs[4194];
    assign layer1_outputs[1135] = ~(layer0_outputs[9955]) | (layer0_outputs[9682]);
    assign layer1_outputs[1136] = (layer0_outputs[8018]) & ~(layer0_outputs[8053]);
    assign layer1_outputs[1137] = (layer0_outputs[11057]) & (layer0_outputs[9524]);
    assign layer1_outputs[1138] = ~((layer0_outputs[2979]) ^ (layer0_outputs[954]));
    assign layer1_outputs[1139] = ~(layer0_outputs[4703]);
    assign layer1_outputs[1140] = (layer0_outputs[7225]) & ~(layer0_outputs[7046]);
    assign layer1_outputs[1141] = ~(layer0_outputs[12394]);
    assign layer1_outputs[1142] = (layer0_outputs[92]) ^ (layer0_outputs[10482]);
    assign layer1_outputs[1143] = layer0_outputs[6710];
    assign layer1_outputs[1144] = (layer0_outputs[11178]) ^ (layer0_outputs[2587]);
    assign layer1_outputs[1145] = ~(layer0_outputs[650]);
    assign layer1_outputs[1146] = ~(layer0_outputs[8425]);
    assign layer1_outputs[1147] = ~(layer0_outputs[5340]) | (layer0_outputs[3379]);
    assign layer1_outputs[1148] = ~((layer0_outputs[8592]) | (layer0_outputs[1563]));
    assign layer1_outputs[1149] = ~(layer0_outputs[3888]) | (layer0_outputs[2353]);
    assign layer1_outputs[1150] = ~((layer0_outputs[5893]) & (layer0_outputs[5564]));
    assign layer1_outputs[1151] = ~(layer0_outputs[4908]) | (layer0_outputs[11044]);
    assign layer1_outputs[1152] = ~(layer0_outputs[11483]);
    assign layer1_outputs[1153] = ~(layer0_outputs[1632]);
    assign layer1_outputs[1154] = ~((layer0_outputs[8320]) | (layer0_outputs[12286]));
    assign layer1_outputs[1155] = ~((layer0_outputs[4770]) ^ (layer0_outputs[8434]));
    assign layer1_outputs[1156] = (layer0_outputs[7108]) & (layer0_outputs[3704]);
    assign layer1_outputs[1157] = ~(layer0_outputs[341]);
    assign layer1_outputs[1158] = ~(layer0_outputs[12758]);
    assign layer1_outputs[1159] = layer0_outputs[6753];
    assign layer1_outputs[1160] = (layer0_outputs[6594]) & ~(layer0_outputs[7437]);
    assign layer1_outputs[1161] = layer0_outputs[232];
    assign layer1_outputs[1162] = ~((layer0_outputs[2366]) | (layer0_outputs[1297]));
    assign layer1_outputs[1163] = ~(layer0_outputs[3826]);
    assign layer1_outputs[1164] = ~(layer0_outputs[1371]) | (layer0_outputs[3997]);
    assign layer1_outputs[1165] = ~(layer0_outputs[12504]) | (layer0_outputs[6528]);
    assign layer1_outputs[1166] = ~(layer0_outputs[11955]);
    assign layer1_outputs[1167] = ~((layer0_outputs[9020]) & (layer0_outputs[3591]));
    assign layer1_outputs[1168] = ~((layer0_outputs[1877]) ^ (layer0_outputs[10763]));
    assign layer1_outputs[1169] = ~(layer0_outputs[10892]) | (layer0_outputs[3607]);
    assign layer1_outputs[1170] = (layer0_outputs[11250]) | (layer0_outputs[1847]);
    assign layer1_outputs[1171] = ~(layer0_outputs[8864]);
    assign layer1_outputs[1172] = ~((layer0_outputs[10625]) | (layer0_outputs[1574]));
    assign layer1_outputs[1173] = ~(layer0_outputs[5647]) | (layer0_outputs[6778]);
    assign layer1_outputs[1174] = layer0_outputs[5694];
    assign layer1_outputs[1175] = ~(layer0_outputs[9801]);
    assign layer1_outputs[1176] = (layer0_outputs[10360]) & (layer0_outputs[5580]);
    assign layer1_outputs[1177] = 1'b1;
    assign layer1_outputs[1178] = layer0_outputs[669];
    assign layer1_outputs[1179] = (layer0_outputs[8093]) & ~(layer0_outputs[10090]);
    assign layer1_outputs[1180] = (layer0_outputs[11994]) & (layer0_outputs[584]);
    assign layer1_outputs[1181] = ~((layer0_outputs[6300]) & (layer0_outputs[1669]));
    assign layer1_outputs[1182] = (layer0_outputs[12382]) & ~(layer0_outputs[6581]);
    assign layer1_outputs[1183] = ~(layer0_outputs[9194]) | (layer0_outputs[9708]);
    assign layer1_outputs[1184] = ~(layer0_outputs[5491]) | (layer0_outputs[5901]);
    assign layer1_outputs[1185] = ~((layer0_outputs[1063]) & (layer0_outputs[3804]));
    assign layer1_outputs[1186] = (layer0_outputs[4652]) & ~(layer0_outputs[5142]);
    assign layer1_outputs[1187] = layer0_outputs[11068];
    assign layer1_outputs[1188] = (layer0_outputs[7843]) ^ (layer0_outputs[7243]);
    assign layer1_outputs[1189] = ~((layer0_outputs[12592]) | (layer0_outputs[3796]));
    assign layer1_outputs[1190] = (layer0_outputs[3113]) & ~(layer0_outputs[4246]);
    assign layer1_outputs[1191] = ~(layer0_outputs[3585]) | (layer0_outputs[5192]);
    assign layer1_outputs[1192] = layer0_outputs[6944];
    assign layer1_outputs[1193] = (layer0_outputs[8528]) | (layer0_outputs[7419]);
    assign layer1_outputs[1194] = ~(layer0_outputs[10411]);
    assign layer1_outputs[1195] = (layer0_outputs[1868]) & ~(layer0_outputs[5402]);
    assign layer1_outputs[1196] = layer0_outputs[7498];
    assign layer1_outputs[1197] = ~((layer0_outputs[8798]) ^ (layer0_outputs[10928]));
    assign layer1_outputs[1198] = (layer0_outputs[9821]) & ~(layer0_outputs[5539]);
    assign layer1_outputs[1199] = (layer0_outputs[69]) & ~(layer0_outputs[5610]);
    assign layer1_outputs[1200] = ~((layer0_outputs[4370]) & (layer0_outputs[8415]));
    assign layer1_outputs[1201] = layer0_outputs[11155];
    assign layer1_outputs[1202] = (layer0_outputs[1382]) & (layer0_outputs[11808]);
    assign layer1_outputs[1203] = layer0_outputs[1146];
    assign layer1_outputs[1204] = layer0_outputs[12238];
    assign layer1_outputs[1205] = layer0_outputs[6762];
    assign layer1_outputs[1206] = layer0_outputs[4817];
    assign layer1_outputs[1207] = ~((layer0_outputs[2300]) | (layer0_outputs[721]));
    assign layer1_outputs[1208] = (layer0_outputs[2920]) | (layer0_outputs[9460]);
    assign layer1_outputs[1209] = ~((layer0_outputs[3218]) & (layer0_outputs[5611]));
    assign layer1_outputs[1210] = ~(layer0_outputs[12538]);
    assign layer1_outputs[1211] = layer0_outputs[5294];
    assign layer1_outputs[1212] = ~((layer0_outputs[7104]) | (layer0_outputs[5936]));
    assign layer1_outputs[1213] = layer0_outputs[7124];
    assign layer1_outputs[1214] = layer0_outputs[2748];
    assign layer1_outputs[1215] = (layer0_outputs[10729]) & ~(layer0_outputs[5457]);
    assign layer1_outputs[1216] = layer0_outputs[8653];
    assign layer1_outputs[1217] = layer0_outputs[5419];
    assign layer1_outputs[1218] = (layer0_outputs[10300]) & ~(layer0_outputs[2921]);
    assign layer1_outputs[1219] = (layer0_outputs[2585]) | (layer0_outputs[6131]);
    assign layer1_outputs[1220] = layer0_outputs[7465];
    assign layer1_outputs[1221] = layer0_outputs[725];
    assign layer1_outputs[1222] = (layer0_outputs[6105]) ^ (layer0_outputs[9289]);
    assign layer1_outputs[1223] = ~(layer0_outputs[5737]);
    assign layer1_outputs[1224] = 1'b0;
    assign layer1_outputs[1225] = ~(layer0_outputs[3145]) | (layer0_outputs[8272]);
    assign layer1_outputs[1226] = ~(layer0_outputs[1477]);
    assign layer1_outputs[1227] = ~(layer0_outputs[2644]);
    assign layer1_outputs[1228] = layer0_outputs[1845];
    assign layer1_outputs[1229] = layer0_outputs[5293];
    assign layer1_outputs[1230] = ~((layer0_outputs[11439]) & (layer0_outputs[3343]));
    assign layer1_outputs[1231] = ~(layer0_outputs[1689]);
    assign layer1_outputs[1232] = (layer0_outputs[5493]) & ~(layer0_outputs[3967]);
    assign layer1_outputs[1233] = (layer0_outputs[1513]) & ~(layer0_outputs[1777]);
    assign layer1_outputs[1234] = ~((layer0_outputs[2991]) ^ (layer0_outputs[2894]));
    assign layer1_outputs[1235] = layer0_outputs[11839];
    assign layer1_outputs[1236] = ~(layer0_outputs[10123]) | (layer0_outputs[5740]);
    assign layer1_outputs[1237] = ~(layer0_outputs[1439]);
    assign layer1_outputs[1238] = layer0_outputs[9];
    assign layer1_outputs[1239] = (layer0_outputs[5274]) ^ (layer0_outputs[11488]);
    assign layer1_outputs[1240] = ~(layer0_outputs[1394]);
    assign layer1_outputs[1241] = ~((layer0_outputs[10451]) ^ (layer0_outputs[11374]));
    assign layer1_outputs[1242] = ~((layer0_outputs[6466]) | (layer0_outputs[4009]));
    assign layer1_outputs[1243] = ~((layer0_outputs[708]) & (layer0_outputs[12593]));
    assign layer1_outputs[1244] = ~(layer0_outputs[5490]) | (layer0_outputs[5802]);
    assign layer1_outputs[1245] = ~(layer0_outputs[2993]);
    assign layer1_outputs[1246] = ~((layer0_outputs[5586]) | (layer0_outputs[7363]));
    assign layer1_outputs[1247] = ~((layer0_outputs[6746]) & (layer0_outputs[6219]));
    assign layer1_outputs[1248] = ~((layer0_outputs[9578]) | (layer0_outputs[11991]));
    assign layer1_outputs[1249] = (layer0_outputs[1665]) & ~(layer0_outputs[1255]);
    assign layer1_outputs[1250] = (layer0_outputs[10372]) & ~(layer0_outputs[1973]);
    assign layer1_outputs[1251] = ~((layer0_outputs[505]) ^ (layer0_outputs[1077]));
    assign layer1_outputs[1252] = ~((layer0_outputs[7876]) | (layer0_outputs[8355]));
    assign layer1_outputs[1253] = ~(layer0_outputs[5930]) | (layer0_outputs[9791]);
    assign layer1_outputs[1254] = layer0_outputs[11133];
    assign layer1_outputs[1255] = ~(layer0_outputs[3111]);
    assign layer1_outputs[1256] = layer0_outputs[3848];
    assign layer1_outputs[1257] = ~((layer0_outputs[2378]) ^ (layer0_outputs[11998]));
    assign layer1_outputs[1258] = ~((layer0_outputs[4874]) & (layer0_outputs[2051]));
    assign layer1_outputs[1259] = ~(layer0_outputs[8322]);
    assign layer1_outputs[1260] = ~(layer0_outputs[4805]) | (layer0_outputs[2615]);
    assign layer1_outputs[1261] = ~((layer0_outputs[5361]) & (layer0_outputs[9341]));
    assign layer1_outputs[1262] = layer0_outputs[10275];
    assign layer1_outputs[1263] = ~((layer0_outputs[4206]) | (layer0_outputs[5697]));
    assign layer1_outputs[1264] = layer0_outputs[12738];
    assign layer1_outputs[1265] = (layer0_outputs[3990]) & (layer0_outputs[10720]);
    assign layer1_outputs[1266] = ~(layer0_outputs[5283]) | (layer0_outputs[5593]);
    assign layer1_outputs[1267] = (layer0_outputs[4118]) & (layer0_outputs[9412]);
    assign layer1_outputs[1268] = (layer0_outputs[4267]) | (layer0_outputs[12035]);
    assign layer1_outputs[1269] = ~(layer0_outputs[11646]) | (layer0_outputs[9205]);
    assign layer1_outputs[1270] = (layer0_outputs[3558]) | (layer0_outputs[10062]);
    assign layer1_outputs[1271] = ~((layer0_outputs[12441]) & (layer0_outputs[4187]));
    assign layer1_outputs[1272] = (layer0_outputs[6806]) & ~(layer0_outputs[7324]);
    assign layer1_outputs[1273] = ~((layer0_outputs[5742]) & (layer0_outputs[764]));
    assign layer1_outputs[1274] = ~((layer0_outputs[621]) | (layer0_outputs[3976]));
    assign layer1_outputs[1275] = (layer0_outputs[8002]) ^ (layer0_outputs[4617]);
    assign layer1_outputs[1276] = layer0_outputs[10149];
    assign layer1_outputs[1277] = ~(layer0_outputs[9965]);
    assign layer1_outputs[1278] = (layer0_outputs[5937]) | (layer0_outputs[9209]);
    assign layer1_outputs[1279] = layer0_outputs[12726];
    assign layer1_outputs[1280] = (layer0_outputs[8269]) | (layer0_outputs[8640]);
    assign layer1_outputs[1281] = layer0_outputs[699];
    assign layer1_outputs[1282] = ~((layer0_outputs[366]) | (layer0_outputs[1640]));
    assign layer1_outputs[1283] = ~(layer0_outputs[5542]);
    assign layer1_outputs[1284] = ~(layer0_outputs[251]) | (layer0_outputs[3712]);
    assign layer1_outputs[1285] = (layer0_outputs[12595]) & (layer0_outputs[11978]);
    assign layer1_outputs[1286] = layer0_outputs[4335];
    assign layer1_outputs[1287] = ~((layer0_outputs[12631]) | (layer0_outputs[5445]));
    assign layer1_outputs[1288] = (layer0_outputs[10877]) | (layer0_outputs[3920]);
    assign layer1_outputs[1289] = layer0_outputs[10862];
    assign layer1_outputs[1290] = (layer0_outputs[8805]) | (layer0_outputs[9295]);
    assign layer1_outputs[1291] = ~(layer0_outputs[996]);
    assign layer1_outputs[1292] = layer0_outputs[11322];
    assign layer1_outputs[1293] = ~(layer0_outputs[4308]);
    assign layer1_outputs[1294] = (layer0_outputs[4437]) & (layer0_outputs[7778]);
    assign layer1_outputs[1295] = (layer0_outputs[5838]) & ~(layer0_outputs[10022]);
    assign layer1_outputs[1296] = ~(layer0_outputs[5815]);
    assign layer1_outputs[1297] = (layer0_outputs[4599]) & ~(layer0_outputs[12295]);
    assign layer1_outputs[1298] = 1'b1;
    assign layer1_outputs[1299] = layer0_outputs[11564];
    assign layer1_outputs[1300] = layer0_outputs[9534];
    assign layer1_outputs[1301] = ~(layer0_outputs[7018]) | (layer0_outputs[3455]);
    assign layer1_outputs[1302] = ~(layer0_outputs[12158]) | (layer0_outputs[6749]);
    assign layer1_outputs[1303] = ~(layer0_outputs[2039]) | (layer0_outputs[2852]);
    assign layer1_outputs[1304] = ~((layer0_outputs[1259]) | (layer0_outputs[4751]));
    assign layer1_outputs[1305] = layer0_outputs[678];
    assign layer1_outputs[1306] = ~((layer0_outputs[5685]) & (layer0_outputs[4746]));
    assign layer1_outputs[1307] = (layer0_outputs[7953]) & ~(layer0_outputs[7676]);
    assign layer1_outputs[1308] = ~(layer0_outputs[6812]) | (layer0_outputs[1409]);
    assign layer1_outputs[1309] = layer0_outputs[2945];
    assign layer1_outputs[1310] = ~(layer0_outputs[5941]);
    assign layer1_outputs[1311] = (layer0_outputs[7927]) ^ (layer0_outputs[6462]);
    assign layer1_outputs[1312] = ~((layer0_outputs[1688]) | (layer0_outputs[470]));
    assign layer1_outputs[1313] = ~(layer0_outputs[6529]);
    assign layer1_outputs[1314] = (layer0_outputs[10014]) & ~(layer0_outputs[2777]);
    assign layer1_outputs[1315] = ~(layer0_outputs[1704]);
    assign layer1_outputs[1316] = layer0_outputs[4453];
    assign layer1_outputs[1317] = (layer0_outputs[263]) & (layer0_outputs[9447]);
    assign layer1_outputs[1318] = (layer0_outputs[12772]) & ~(layer0_outputs[665]);
    assign layer1_outputs[1319] = ~(layer0_outputs[5088]);
    assign layer1_outputs[1320] = (layer0_outputs[12297]) ^ (layer0_outputs[7621]);
    assign layer1_outputs[1321] = ~(layer0_outputs[11844]);
    assign layer1_outputs[1322] = ~(layer0_outputs[3391]) | (layer0_outputs[10713]);
    assign layer1_outputs[1323] = ~((layer0_outputs[2697]) & (layer0_outputs[3243]));
    assign layer1_outputs[1324] = ~(layer0_outputs[8320]) | (layer0_outputs[725]);
    assign layer1_outputs[1325] = layer0_outputs[11787];
    assign layer1_outputs[1326] = ~(layer0_outputs[1653]);
    assign layer1_outputs[1327] = ~((layer0_outputs[5725]) | (layer0_outputs[2805]));
    assign layer1_outputs[1328] = ~((layer0_outputs[1475]) ^ (layer0_outputs[4093]));
    assign layer1_outputs[1329] = ~((layer0_outputs[3528]) ^ (layer0_outputs[9515]));
    assign layer1_outputs[1330] = ~(layer0_outputs[2220]);
    assign layer1_outputs[1331] = ~((layer0_outputs[3003]) | (layer0_outputs[2340]));
    assign layer1_outputs[1332] = (layer0_outputs[4369]) & ~(layer0_outputs[12606]);
    assign layer1_outputs[1333] = ~((layer0_outputs[10260]) | (layer0_outputs[1539]));
    assign layer1_outputs[1334] = (layer0_outputs[6926]) | (layer0_outputs[11735]);
    assign layer1_outputs[1335] = layer0_outputs[664];
    assign layer1_outputs[1336] = ~(layer0_outputs[861]);
    assign layer1_outputs[1337] = (layer0_outputs[8559]) | (layer0_outputs[9833]);
    assign layer1_outputs[1338] = ~(layer0_outputs[3150]) | (layer0_outputs[5027]);
    assign layer1_outputs[1339] = ~(layer0_outputs[7654]) | (layer0_outputs[11114]);
    assign layer1_outputs[1340] = ~((layer0_outputs[7645]) & (layer0_outputs[890]));
    assign layer1_outputs[1341] = layer0_outputs[8563];
    assign layer1_outputs[1342] = ~((layer0_outputs[3989]) | (layer0_outputs[11418]));
    assign layer1_outputs[1343] = ~((layer0_outputs[8616]) | (layer0_outputs[7829]));
    assign layer1_outputs[1344] = (layer0_outputs[1969]) ^ (layer0_outputs[5474]);
    assign layer1_outputs[1345] = ~(layer0_outputs[11761]) | (layer0_outputs[2461]);
    assign layer1_outputs[1346] = ~((layer0_outputs[9777]) & (layer0_outputs[6088]));
    assign layer1_outputs[1347] = layer0_outputs[12461];
    assign layer1_outputs[1348] = ~(layer0_outputs[6433]);
    assign layer1_outputs[1349] = ~(layer0_outputs[1460]);
    assign layer1_outputs[1350] = ~(layer0_outputs[6882]);
    assign layer1_outputs[1351] = ~(layer0_outputs[3040]);
    assign layer1_outputs[1352] = 1'b0;
    assign layer1_outputs[1353] = (layer0_outputs[12276]) ^ (layer0_outputs[8166]);
    assign layer1_outputs[1354] = ~((layer0_outputs[10985]) & (layer0_outputs[2871]));
    assign layer1_outputs[1355] = ~(layer0_outputs[8217]);
    assign layer1_outputs[1356] = ~(layer0_outputs[265]);
    assign layer1_outputs[1357] = ~(layer0_outputs[2114]);
    assign layer1_outputs[1358] = ~((layer0_outputs[10189]) | (layer0_outputs[11692]));
    assign layer1_outputs[1359] = ~((layer0_outputs[11006]) & (layer0_outputs[7576]));
    assign layer1_outputs[1360] = ~(layer0_outputs[5928]);
    assign layer1_outputs[1361] = 1'b0;
    assign layer1_outputs[1362] = layer0_outputs[4662];
    assign layer1_outputs[1363] = layer0_outputs[347];
    assign layer1_outputs[1364] = (layer0_outputs[6195]) | (layer0_outputs[8949]);
    assign layer1_outputs[1365] = (layer0_outputs[1956]) & ~(layer0_outputs[4028]);
    assign layer1_outputs[1366] = ~((layer0_outputs[3017]) & (layer0_outputs[8668]));
    assign layer1_outputs[1367] = ~(layer0_outputs[8346]);
    assign layer1_outputs[1368] = (layer0_outputs[8907]) ^ (layer0_outputs[12040]);
    assign layer1_outputs[1369] = (layer0_outputs[191]) | (layer0_outputs[5003]);
    assign layer1_outputs[1370] = layer0_outputs[6693];
    assign layer1_outputs[1371] = layer0_outputs[8772];
    assign layer1_outputs[1372] = (layer0_outputs[11621]) | (layer0_outputs[10910]);
    assign layer1_outputs[1373] = layer0_outputs[6734];
    assign layer1_outputs[1374] = (layer0_outputs[7837]) & ~(layer0_outputs[9395]);
    assign layer1_outputs[1375] = 1'b0;
    assign layer1_outputs[1376] = (layer0_outputs[10818]) & (layer0_outputs[12337]);
    assign layer1_outputs[1377] = layer0_outputs[5217];
    assign layer1_outputs[1378] = ~(layer0_outputs[4821]);
    assign layer1_outputs[1379] = layer0_outputs[10171];
    assign layer1_outputs[1380] = ~(layer0_outputs[8725]);
    assign layer1_outputs[1381] = (layer0_outputs[8124]) ^ (layer0_outputs[8092]);
    assign layer1_outputs[1382] = (layer0_outputs[9557]) & ~(layer0_outputs[4098]);
    assign layer1_outputs[1383] = layer0_outputs[2967];
    assign layer1_outputs[1384] = layer0_outputs[8795];
    assign layer1_outputs[1385] = layer0_outputs[12733];
    assign layer1_outputs[1386] = (layer0_outputs[6479]) & (layer0_outputs[2400]);
    assign layer1_outputs[1387] = layer0_outputs[11556];
    assign layer1_outputs[1388] = layer0_outputs[7575];
    assign layer1_outputs[1389] = ~(layer0_outputs[6363]);
    assign layer1_outputs[1390] = (layer0_outputs[11578]) & ~(layer0_outputs[8874]);
    assign layer1_outputs[1391] = ~(layer0_outputs[1269]) | (layer0_outputs[11749]);
    assign layer1_outputs[1392] = ~(layer0_outputs[8413]) | (layer0_outputs[1527]);
    assign layer1_outputs[1393] = layer0_outputs[12556];
    assign layer1_outputs[1394] = ~(layer0_outputs[10034]);
    assign layer1_outputs[1395] = ~(layer0_outputs[4102]);
    assign layer1_outputs[1396] = ~((layer0_outputs[10501]) & (layer0_outputs[11917]));
    assign layer1_outputs[1397] = ~((layer0_outputs[1768]) & (layer0_outputs[8725]));
    assign layer1_outputs[1398] = layer0_outputs[12032];
    assign layer1_outputs[1399] = (layer0_outputs[4567]) ^ (layer0_outputs[7965]);
    assign layer1_outputs[1400] = (layer0_outputs[2094]) & ~(layer0_outputs[1404]);
    assign layer1_outputs[1401] = (layer0_outputs[2569]) & ~(layer0_outputs[5569]);
    assign layer1_outputs[1402] = ~(layer0_outputs[12671]);
    assign layer1_outputs[1403] = layer0_outputs[8993];
    assign layer1_outputs[1404] = ~(layer0_outputs[7877]);
    assign layer1_outputs[1405] = layer0_outputs[11776];
    assign layer1_outputs[1406] = ~(layer0_outputs[1732]) | (layer0_outputs[12735]);
    assign layer1_outputs[1407] = (layer0_outputs[2341]) & ~(layer0_outputs[2056]);
    assign layer1_outputs[1408] = ~((layer0_outputs[1359]) & (layer0_outputs[7361]));
    assign layer1_outputs[1409] = ~((layer0_outputs[6848]) & (layer0_outputs[6538]));
    assign layer1_outputs[1410] = 1'b1;
    assign layer1_outputs[1411] = (layer0_outputs[2285]) ^ (layer0_outputs[927]);
    assign layer1_outputs[1412] = ~(layer0_outputs[2576]) | (layer0_outputs[7209]);
    assign layer1_outputs[1413] = ~(layer0_outputs[7477]);
    assign layer1_outputs[1414] = (layer0_outputs[1700]) ^ (layer0_outputs[11396]);
    assign layer1_outputs[1415] = 1'b1;
    assign layer1_outputs[1416] = layer0_outputs[1944];
    assign layer1_outputs[1417] = ~(layer0_outputs[11025]) | (layer0_outputs[8090]);
    assign layer1_outputs[1418] = ~(layer0_outputs[12428]);
    assign layer1_outputs[1419] = ~(layer0_outputs[6000]) | (layer0_outputs[10134]);
    assign layer1_outputs[1420] = ~(layer0_outputs[9217]);
    assign layer1_outputs[1421] = ~((layer0_outputs[4464]) | (layer0_outputs[4944]));
    assign layer1_outputs[1422] = (layer0_outputs[11597]) & (layer0_outputs[10729]);
    assign layer1_outputs[1423] = ~(layer0_outputs[9003]);
    assign layer1_outputs[1424] = ~(layer0_outputs[6490]);
    assign layer1_outputs[1425] = (layer0_outputs[3162]) & ~(layer0_outputs[5187]);
    assign layer1_outputs[1426] = ~(layer0_outputs[10607]);
    assign layer1_outputs[1427] = (layer0_outputs[6807]) & ~(layer0_outputs[7392]);
    assign layer1_outputs[1428] = layer0_outputs[1646];
    assign layer1_outputs[1429] = layer0_outputs[4143];
    assign layer1_outputs[1430] = ~(layer0_outputs[1846]);
    assign layer1_outputs[1431] = ~(layer0_outputs[8727]);
    assign layer1_outputs[1432] = layer0_outputs[5069];
    assign layer1_outputs[1433] = layer0_outputs[338];
    assign layer1_outputs[1434] = ~(layer0_outputs[11264]);
    assign layer1_outputs[1435] = layer0_outputs[1984];
    assign layer1_outputs[1436] = ~(layer0_outputs[6606]);
    assign layer1_outputs[1437] = layer0_outputs[457];
    assign layer1_outputs[1438] = ~(layer0_outputs[5822]);
    assign layer1_outputs[1439] = (layer0_outputs[676]) ^ (layer0_outputs[4037]);
    assign layer1_outputs[1440] = (layer0_outputs[12320]) & (layer0_outputs[4501]);
    assign layer1_outputs[1441] = layer0_outputs[385];
    assign layer1_outputs[1442] = (layer0_outputs[2477]) & (layer0_outputs[10281]);
    assign layer1_outputs[1443] = ~((layer0_outputs[4458]) & (layer0_outputs[2714]));
    assign layer1_outputs[1444] = layer0_outputs[12424];
    assign layer1_outputs[1445] = ~(layer0_outputs[8138]);
    assign layer1_outputs[1446] = 1'b0;
    assign layer1_outputs[1447] = layer0_outputs[1832];
    assign layer1_outputs[1448] = ~(layer0_outputs[1056]);
    assign layer1_outputs[1449] = (layer0_outputs[11638]) & (layer0_outputs[10441]);
    assign layer1_outputs[1450] = ~(layer0_outputs[7666]);
    assign layer1_outputs[1451] = ~((layer0_outputs[6397]) ^ (layer0_outputs[1136]));
    assign layer1_outputs[1452] = ~(layer0_outputs[10979]) | (layer0_outputs[6315]);
    assign layer1_outputs[1453] = (layer0_outputs[8362]) & ~(layer0_outputs[2889]);
    assign layer1_outputs[1454] = ~(layer0_outputs[6063]);
    assign layer1_outputs[1455] = (layer0_outputs[12224]) ^ (layer0_outputs[9533]);
    assign layer1_outputs[1456] = (layer0_outputs[9037]) & ~(layer0_outputs[4025]);
    assign layer1_outputs[1457] = ~((layer0_outputs[8138]) & (layer0_outputs[2811]));
    assign layer1_outputs[1458] = ~((layer0_outputs[5448]) | (layer0_outputs[7727]));
    assign layer1_outputs[1459] = ~(layer0_outputs[2001]) | (layer0_outputs[5509]);
    assign layer1_outputs[1460] = ~((layer0_outputs[12699]) ^ (layer0_outputs[12750]));
    assign layer1_outputs[1461] = layer0_outputs[6732];
    assign layer1_outputs[1462] = layer0_outputs[7181];
    assign layer1_outputs[1463] = ~(layer0_outputs[1611]) | (layer0_outputs[2942]);
    assign layer1_outputs[1464] = ~(layer0_outputs[6110]);
    assign layer1_outputs[1465] = layer0_outputs[9181];
    assign layer1_outputs[1466] = (layer0_outputs[5609]) & (layer0_outputs[6892]);
    assign layer1_outputs[1467] = ~((layer0_outputs[4347]) ^ (layer0_outputs[4856]));
    assign layer1_outputs[1468] = (layer0_outputs[12692]) & (layer0_outputs[3973]);
    assign layer1_outputs[1469] = layer0_outputs[4042];
    assign layer1_outputs[1470] = ~((layer0_outputs[2835]) ^ (layer0_outputs[455]));
    assign layer1_outputs[1471] = ~(layer0_outputs[6017]) | (layer0_outputs[2062]);
    assign layer1_outputs[1472] = ~(layer0_outputs[5989]);
    assign layer1_outputs[1473] = ~(layer0_outputs[6490]);
    assign layer1_outputs[1474] = layer0_outputs[5749];
    assign layer1_outputs[1475] = ~(layer0_outputs[1197]) | (layer0_outputs[11230]);
    assign layer1_outputs[1476] = ~(layer0_outputs[11831]);
    assign layer1_outputs[1477] = ~(layer0_outputs[10117]);
    assign layer1_outputs[1478] = (layer0_outputs[7677]) & (layer0_outputs[4057]);
    assign layer1_outputs[1479] = ~(layer0_outputs[12276]);
    assign layer1_outputs[1480] = ~(layer0_outputs[3549]);
    assign layer1_outputs[1481] = (layer0_outputs[752]) & (layer0_outputs[2754]);
    assign layer1_outputs[1482] = layer0_outputs[692];
    assign layer1_outputs[1483] = 1'b0;
    assign layer1_outputs[1484] = ~((layer0_outputs[12097]) ^ (layer0_outputs[9706]));
    assign layer1_outputs[1485] = ~(layer0_outputs[6417]);
    assign layer1_outputs[1486] = ~(layer0_outputs[1251]);
    assign layer1_outputs[1487] = (layer0_outputs[3958]) ^ (layer0_outputs[5831]);
    assign layer1_outputs[1488] = (layer0_outputs[10804]) & (layer0_outputs[9819]);
    assign layer1_outputs[1489] = ~((layer0_outputs[1889]) | (layer0_outputs[5604]));
    assign layer1_outputs[1490] = layer0_outputs[995];
    assign layer1_outputs[1491] = ~(layer0_outputs[3163]) | (layer0_outputs[1950]);
    assign layer1_outputs[1492] = (layer0_outputs[11016]) ^ (layer0_outputs[8767]);
    assign layer1_outputs[1493] = (layer0_outputs[10810]) & ~(layer0_outputs[7425]);
    assign layer1_outputs[1494] = ~((layer0_outputs[10242]) | (layer0_outputs[2357]));
    assign layer1_outputs[1495] = ~(layer0_outputs[5057]);
    assign layer1_outputs[1496] = ~(layer0_outputs[6895]);
    assign layer1_outputs[1497] = ~((layer0_outputs[6158]) & (layer0_outputs[9173]));
    assign layer1_outputs[1498] = (layer0_outputs[7912]) & (layer0_outputs[3547]);
    assign layer1_outputs[1499] = layer0_outputs[4549];
    assign layer1_outputs[1500] = ~(layer0_outputs[12613]) | (layer0_outputs[10237]);
    assign layer1_outputs[1501] = (layer0_outputs[769]) | (layer0_outputs[3090]);
    assign layer1_outputs[1502] = (layer0_outputs[11478]) & ~(layer0_outputs[10132]);
    assign layer1_outputs[1503] = (layer0_outputs[11858]) & ~(layer0_outputs[1462]);
    assign layer1_outputs[1504] = ~((layer0_outputs[5055]) & (layer0_outputs[9107]));
    assign layer1_outputs[1505] = layer0_outputs[8552];
    assign layer1_outputs[1506] = (layer0_outputs[11474]) | (layer0_outputs[33]);
    assign layer1_outputs[1507] = ~(layer0_outputs[6920]);
    assign layer1_outputs[1508] = ~(layer0_outputs[7118]);
    assign layer1_outputs[1509] = ~(layer0_outputs[9513]);
    assign layer1_outputs[1510] = (layer0_outputs[5510]) & ~(layer0_outputs[3965]);
    assign layer1_outputs[1511] = (layer0_outputs[8761]) | (layer0_outputs[7423]);
    assign layer1_outputs[1512] = layer0_outputs[2345];
    assign layer1_outputs[1513] = ~((layer0_outputs[7584]) & (layer0_outputs[6305]));
    assign layer1_outputs[1514] = ~((layer0_outputs[6998]) & (layer0_outputs[6048]));
    assign layer1_outputs[1515] = ~(layer0_outputs[10212]);
    assign layer1_outputs[1516] = (layer0_outputs[9541]) & ~(layer0_outputs[4783]);
    assign layer1_outputs[1517] = ~((layer0_outputs[5180]) ^ (layer0_outputs[7110]));
    assign layer1_outputs[1518] = (layer0_outputs[9609]) & (layer0_outputs[5242]);
    assign layer1_outputs[1519] = (layer0_outputs[9180]) & ~(layer0_outputs[2061]);
    assign layer1_outputs[1520] = ~(layer0_outputs[1805]);
    assign layer1_outputs[1521] = (layer0_outputs[3884]) & (layer0_outputs[3903]);
    assign layer1_outputs[1522] = layer0_outputs[10358];
    assign layer1_outputs[1523] = (layer0_outputs[10294]) & (layer0_outputs[839]);
    assign layer1_outputs[1524] = ~(layer0_outputs[2690]);
    assign layer1_outputs[1525] = (layer0_outputs[4543]) ^ (layer0_outputs[6457]);
    assign layer1_outputs[1526] = (layer0_outputs[5412]) & ~(layer0_outputs[5762]);
    assign layer1_outputs[1527] = ~(layer0_outputs[9855]);
    assign layer1_outputs[1528] = (layer0_outputs[4985]) ^ (layer0_outputs[7748]);
    assign layer1_outputs[1529] = layer0_outputs[8371];
    assign layer1_outputs[1530] = layer0_outputs[10611];
    assign layer1_outputs[1531] = (layer0_outputs[1922]) | (layer0_outputs[10382]);
    assign layer1_outputs[1532] = (layer0_outputs[7102]) | (layer0_outputs[6711]);
    assign layer1_outputs[1533] = ~(layer0_outputs[9652]);
    assign layer1_outputs[1534] = ~(layer0_outputs[7838]);
    assign layer1_outputs[1535] = (layer0_outputs[10924]) | (layer0_outputs[1262]);
    assign layer1_outputs[1536] = ~(layer0_outputs[11513]);
    assign layer1_outputs[1537] = (layer0_outputs[2863]) ^ (layer0_outputs[1098]);
    assign layer1_outputs[1538] = (layer0_outputs[9408]) & ~(layer0_outputs[83]);
    assign layer1_outputs[1539] = layer0_outputs[11563];
    assign layer1_outputs[1540] = (layer0_outputs[201]) & ~(layer0_outputs[6697]);
    assign layer1_outputs[1541] = (layer0_outputs[10180]) | (layer0_outputs[10509]);
    assign layer1_outputs[1542] = (layer0_outputs[4709]) | (layer0_outputs[9118]);
    assign layer1_outputs[1543] = layer0_outputs[2532];
    assign layer1_outputs[1544] = ~((layer0_outputs[5760]) & (layer0_outputs[4798]));
    assign layer1_outputs[1545] = (layer0_outputs[489]) & ~(layer0_outputs[5069]);
    assign layer1_outputs[1546] = ~(layer0_outputs[3799]);
    assign layer1_outputs[1547] = (layer0_outputs[6733]) & ~(layer0_outputs[1734]);
    assign layer1_outputs[1548] = ~(layer0_outputs[6946]);
    assign layer1_outputs[1549] = ~(layer0_outputs[820]);
    assign layer1_outputs[1550] = (layer0_outputs[311]) & ~(layer0_outputs[2375]);
    assign layer1_outputs[1551] = (layer0_outputs[8263]) & (layer0_outputs[447]);
    assign layer1_outputs[1552] = ~(layer0_outputs[9986]) | (layer0_outputs[9645]);
    assign layer1_outputs[1553] = ~(layer0_outputs[9630]);
    assign layer1_outputs[1554] = ~(layer0_outputs[8288]);
    assign layer1_outputs[1555] = layer0_outputs[4881];
    assign layer1_outputs[1556] = ~(layer0_outputs[9828]);
    assign layer1_outputs[1557] = ~(layer0_outputs[8434]);
    assign layer1_outputs[1558] = ~((layer0_outputs[12632]) | (layer0_outputs[3987]));
    assign layer1_outputs[1559] = ~(layer0_outputs[3815]);
    assign layer1_outputs[1560] = layer0_outputs[8697];
    assign layer1_outputs[1561] = layer0_outputs[1033];
    assign layer1_outputs[1562] = layer0_outputs[10331];
    assign layer1_outputs[1563] = layer0_outputs[4830];
    assign layer1_outputs[1564] = (layer0_outputs[9658]) & (layer0_outputs[10922]);
    assign layer1_outputs[1565] = (layer0_outputs[404]) & ~(layer0_outputs[9028]);
    assign layer1_outputs[1566] = ~((layer0_outputs[11584]) & (layer0_outputs[8557]));
    assign layer1_outputs[1567] = layer0_outputs[12708];
    assign layer1_outputs[1568] = (layer0_outputs[8294]) & ~(layer0_outputs[8888]);
    assign layer1_outputs[1569] = ~(layer0_outputs[5794]) | (layer0_outputs[8838]);
    assign layer1_outputs[1570] = ~((layer0_outputs[9969]) & (layer0_outputs[4926]));
    assign layer1_outputs[1571] = ~(layer0_outputs[2698]);
    assign layer1_outputs[1572] = layer0_outputs[15];
    assign layer1_outputs[1573] = ~((layer0_outputs[4289]) | (layer0_outputs[2690]));
    assign layer1_outputs[1574] = layer0_outputs[4895];
    assign layer1_outputs[1575] = ~((layer0_outputs[4984]) ^ (layer0_outputs[3149]));
    assign layer1_outputs[1576] = ~(layer0_outputs[5667]);
    assign layer1_outputs[1577] = ~(layer0_outputs[6539]) | (layer0_outputs[7860]);
    assign layer1_outputs[1578] = ~(layer0_outputs[221]);
    assign layer1_outputs[1579] = layer0_outputs[10960];
    assign layer1_outputs[1580] = (layer0_outputs[4377]) ^ (layer0_outputs[10072]);
    assign layer1_outputs[1581] = ~((layer0_outputs[3031]) | (layer0_outputs[1856]));
    assign layer1_outputs[1582] = ~(layer0_outputs[8068]);
    assign layer1_outputs[1583] = ~((layer0_outputs[749]) | (layer0_outputs[7256]));
    assign layer1_outputs[1584] = ~(layer0_outputs[10834]);
    assign layer1_outputs[1585] = layer0_outputs[4862];
    assign layer1_outputs[1586] = layer0_outputs[6943];
    assign layer1_outputs[1587] = ~(layer0_outputs[2125]);
    assign layer1_outputs[1588] = (layer0_outputs[4399]) & (layer0_outputs[8923]);
    assign layer1_outputs[1589] = ~(layer0_outputs[4216]);
    assign layer1_outputs[1590] = ~((layer0_outputs[145]) & (layer0_outputs[11956]));
    assign layer1_outputs[1591] = ~(layer0_outputs[7470]);
    assign layer1_outputs[1592] = (layer0_outputs[5113]) ^ (layer0_outputs[1667]);
    assign layer1_outputs[1593] = layer0_outputs[4761];
    assign layer1_outputs[1594] = ~((layer0_outputs[9073]) ^ (layer0_outputs[5288]));
    assign layer1_outputs[1595] = ~(layer0_outputs[6127]) | (layer0_outputs[1528]);
    assign layer1_outputs[1596] = ~(layer0_outputs[229]);
    assign layer1_outputs[1597] = layer0_outputs[8051];
    assign layer1_outputs[1598] = (layer0_outputs[12371]) & ~(layer0_outputs[1332]);
    assign layer1_outputs[1599] = layer0_outputs[10586];
    assign layer1_outputs[1600] = ~((layer0_outputs[12077]) & (layer0_outputs[10303]));
    assign layer1_outputs[1601] = (layer0_outputs[10659]) & ~(layer0_outputs[10780]);
    assign layer1_outputs[1602] = ~(layer0_outputs[7428]) | (layer0_outputs[9036]);
    assign layer1_outputs[1603] = ~(layer0_outputs[8264]) | (layer0_outputs[7532]);
    assign layer1_outputs[1604] = ~(layer0_outputs[1807]);
    assign layer1_outputs[1605] = ~(layer0_outputs[4927]);
    assign layer1_outputs[1606] = ~((layer0_outputs[11710]) ^ (layer0_outputs[1756]));
    assign layer1_outputs[1607] = ~(layer0_outputs[6556]);
    assign layer1_outputs[1608] = (layer0_outputs[10452]) & ~(layer0_outputs[759]);
    assign layer1_outputs[1609] = (layer0_outputs[6907]) & ~(layer0_outputs[11374]);
    assign layer1_outputs[1610] = (layer0_outputs[8289]) | (layer0_outputs[6507]);
    assign layer1_outputs[1611] = layer0_outputs[12425];
    assign layer1_outputs[1612] = ~(layer0_outputs[12096]);
    assign layer1_outputs[1613] = ~((layer0_outputs[12762]) | (layer0_outputs[1586]));
    assign layer1_outputs[1614] = ~((layer0_outputs[10942]) ^ (layer0_outputs[12542]));
    assign layer1_outputs[1615] = layer0_outputs[9013];
    assign layer1_outputs[1616] = ~(layer0_outputs[9266]);
    assign layer1_outputs[1617] = ~(layer0_outputs[4398]);
    assign layer1_outputs[1618] = ~(layer0_outputs[12508]) | (layer0_outputs[6696]);
    assign layer1_outputs[1619] = (layer0_outputs[703]) | (layer0_outputs[8123]);
    assign layer1_outputs[1620] = layer0_outputs[1211];
    assign layer1_outputs[1621] = ~((layer0_outputs[5154]) & (layer0_outputs[401]));
    assign layer1_outputs[1622] = ~(layer0_outputs[579]);
    assign layer1_outputs[1623] = ~(layer0_outputs[9601]) | (layer0_outputs[5332]);
    assign layer1_outputs[1624] = (layer0_outputs[3704]) | (layer0_outputs[8125]);
    assign layer1_outputs[1625] = ~(layer0_outputs[11449]);
    assign layer1_outputs[1626] = (layer0_outputs[2010]) | (layer0_outputs[12739]);
    assign layer1_outputs[1627] = layer0_outputs[6151];
    assign layer1_outputs[1628] = ~(layer0_outputs[12328]);
    assign layer1_outputs[1629] = ~(layer0_outputs[11441]);
    assign layer1_outputs[1630] = ~(layer0_outputs[10183]);
    assign layer1_outputs[1631] = ~(layer0_outputs[584]) | (layer0_outputs[8618]);
    assign layer1_outputs[1632] = (layer0_outputs[947]) ^ (layer0_outputs[1030]);
    assign layer1_outputs[1633] = ~(layer0_outputs[10393]);
    assign layer1_outputs[1634] = ~(layer0_outputs[12746]);
    assign layer1_outputs[1635] = layer0_outputs[4837];
    assign layer1_outputs[1636] = layer0_outputs[8507];
    assign layer1_outputs[1637] = ~((layer0_outputs[11390]) ^ (layer0_outputs[11007]));
    assign layer1_outputs[1638] = ~(layer0_outputs[6451]) | (layer0_outputs[6157]);
    assign layer1_outputs[1639] = (layer0_outputs[10402]) ^ (layer0_outputs[11078]);
    assign layer1_outputs[1640] = ~((layer0_outputs[3072]) & (layer0_outputs[11882]));
    assign layer1_outputs[1641] = (layer0_outputs[4427]) ^ (layer0_outputs[10241]);
    assign layer1_outputs[1642] = (layer0_outputs[3673]) & ~(layer0_outputs[667]);
    assign layer1_outputs[1643] = ~(layer0_outputs[10657]) | (layer0_outputs[4108]);
    assign layer1_outputs[1644] = (layer0_outputs[11332]) & ~(layer0_outputs[6903]);
    assign layer1_outputs[1645] = layer0_outputs[1674];
    assign layer1_outputs[1646] = ~(layer0_outputs[4665]);
    assign layer1_outputs[1647] = ~((layer0_outputs[9008]) | (layer0_outputs[831]));
    assign layer1_outputs[1648] = ~(layer0_outputs[1324]);
    assign layer1_outputs[1649] = (layer0_outputs[648]) & (layer0_outputs[2513]);
    assign layer1_outputs[1650] = layer0_outputs[8155];
    assign layer1_outputs[1651] = ~(layer0_outputs[7730]);
    assign layer1_outputs[1652] = layer0_outputs[8302];
    assign layer1_outputs[1653] = layer0_outputs[9296];
    assign layer1_outputs[1654] = (layer0_outputs[3449]) & (layer0_outputs[1321]);
    assign layer1_outputs[1655] = layer0_outputs[10945];
    assign layer1_outputs[1656] = ~(layer0_outputs[5617]) | (layer0_outputs[10263]);
    assign layer1_outputs[1657] = ~((layer0_outputs[5782]) ^ (layer0_outputs[12312]));
    assign layer1_outputs[1658] = layer0_outputs[10598];
    assign layer1_outputs[1659] = ~(layer0_outputs[2007]);
    assign layer1_outputs[1660] = ~(layer0_outputs[3818]);
    assign layer1_outputs[1661] = layer0_outputs[2964];
    assign layer1_outputs[1662] = ~((layer0_outputs[2992]) & (layer0_outputs[7015]));
    assign layer1_outputs[1663] = ~(layer0_outputs[6413]);
    assign layer1_outputs[1664] = ~(layer0_outputs[11520]);
    assign layer1_outputs[1665] = ~((layer0_outputs[560]) ^ (layer0_outputs[12338]));
    assign layer1_outputs[1666] = (layer0_outputs[983]) & ~(layer0_outputs[6435]);
    assign layer1_outputs[1667] = ~(layer0_outputs[11674]);
    assign layer1_outputs[1668] = ~(layer0_outputs[3411]) | (layer0_outputs[12707]);
    assign layer1_outputs[1669] = (layer0_outputs[11872]) & ~(layer0_outputs[6946]);
    assign layer1_outputs[1670] = 1'b0;
    assign layer1_outputs[1671] = (layer0_outputs[1299]) & (layer0_outputs[1041]);
    assign layer1_outputs[1672] = layer0_outputs[2726];
    assign layer1_outputs[1673] = layer0_outputs[3257];
    assign layer1_outputs[1674] = ~(layer0_outputs[9163]) | (layer0_outputs[470]);
    assign layer1_outputs[1675] = ~((layer0_outputs[4197]) ^ (layer0_outputs[7127]));
    assign layer1_outputs[1676] = (layer0_outputs[9479]) & ~(layer0_outputs[9157]);
    assign layer1_outputs[1677] = layer0_outputs[4244];
    assign layer1_outputs[1678] = ~(layer0_outputs[235]);
    assign layer1_outputs[1679] = (layer0_outputs[2717]) & ~(layer0_outputs[8215]);
    assign layer1_outputs[1680] = layer0_outputs[9704];
    assign layer1_outputs[1681] = (layer0_outputs[5269]) & ~(layer0_outputs[2606]);
    assign layer1_outputs[1682] = (layer0_outputs[3203]) ^ (layer0_outputs[8041]);
    assign layer1_outputs[1683] = layer0_outputs[12225];
    assign layer1_outputs[1684] = ~(layer0_outputs[2342]) | (layer0_outputs[4285]);
    assign layer1_outputs[1685] = layer0_outputs[10334];
    assign layer1_outputs[1686] = ~((layer0_outputs[12364]) | (layer0_outputs[5806]));
    assign layer1_outputs[1687] = ~(layer0_outputs[1082]);
    assign layer1_outputs[1688] = ~(layer0_outputs[3390]);
    assign layer1_outputs[1689] = ~(layer0_outputs[2256]);
    assign layer1_outputs[1690] = (layer0_outputs[11205]) & ~(layer0_outputs[6994]);
    assign layer1_outputs[1691] = ~(layer0_outputs[2225]);
    assign layer1_outputs[1692] = (layer0_outputs[4353]) ^ (layer0_outputs[102]);
    assign layer1_outputs[1693] = (layer0_outputs[7986]) | (layer0_outputs[8885]);
    assign layer1_outputs[1694] = ~((layer0_outputs[6508]) ^ (layer0_outputs[8071]));
    assign layer1_outputs[1695] = layer0_outputs[6558];
    assign layer1_outputs[1696] = (layer0_outputs[6624]) & ~(layer0_outputs[2374]);
    assign layer1_outputs[1697] = ~(layer0_outputs[4463]) | (layer0_outputs[12272]);
    assign layer1_outputs[1698] = ~(layer0_outputs[2517]);
    assign layer1_outputs[1699] = (layer0_outputs[12052]) | (layer0_outputs[6257]);
    assign layer1_outputs[1700] = ~(layer0_outputs[8052]) | (layer0_outputs[11663]);
    assign layer1_outputs[1701] = (layer0_outputs[1279]) & ~(layer0_outputs[9204]);
    assign layer1_outputs[1702] = ~(layer0_outputs[11145]) | (layer0_outputs[2631]);
    assign layer1_outputs[1703] = ~((layer0_outputs[11940]) & (layer0_outputs[6827]));
    assign layer1_outputs[1704] = ~(layer0_outputs[3026]) | (layer0_outputs[3028]);
    assign layer1_outputs[1705] = ~(layer0_outputs[9953]);
    assign layer1_outputs[1706] = ~((layer0_outputs[5985]) | (layer0_outputs[12125]));
    assign layer1_outputs[1707] = 1'b1;
    assign layer1_outputs[1708] = ~(layer0_outputs[9849]) | (layer0_outputs[12064]);
    assign layer1_outputs[1709] = ~(layer0_outputs[12085]);
    assign layer1_outputs[1710] = layer0_outputs[1912];
    assign layer1_outputs[1711] = ~(layer0_outputs[4230]);
    assign layer1_outputs[1712] = ~(layer0_outputs[11447]);
    assign layer1_outputs[1713] = ~(layer0_outputs[11570]) | (layer0_outputs[12540]);
    assign layer1_outputs[1714] = ~(layer0_outputs[540]);
    assign layer1_outputs[1715] = (layer0_outputs[10967]) ^ (layer0_outputs[10310]);
    assign layer1_outputs[1716] = 1'b0;
    assign layer1_outputs[1717] = ~((layer0_outputs[1872]) | (layer0_outputs[436]));
    assign layer1_outputs[1718] = ~(layer0_outputs[1921]);
    assign layer1_outputs[1719] = ~(layer0_outputs[8609]);
    assign layer1_outputs[1720] = layer0_outputs[9868];
    assign layer1_outputs[1721] = ~(layer0_outputs[10542]);
    assign layer1_outputs[1722] = layer0_outputs[12677];
    assign layer1_outputs[1723] = (layer0_outputs[11175]) & ~(layer0_outputs[2741]);
    assign layer1_outputs[1724] = layer0_outputs[71];
    assign layer1_outputs[1725] = ~(layer0_outputs[3]) | (layer0_outputs[4512]);
    assign layer1_outputs[1726] = (layer0_outputs[5138]) & (layer0_outputs[6771]);
    assign layer1_outputs[1727] = layer0_outputs[9399];
    assign layer1_outputs[1728] = ~(layer0_outputs[11964]);
    assign layer1_outputs[1729] = ~((layer0_outputs[628]) ^ (layer0_outputs[11158]));
    assign layer1_outputs[1730] = (layer0_outputs[1202]) ^ (layer0_outputs[7331]);
    assign layer1_outputs[1731] = ~(layer0_outputs[4029]);
    assign layer1_outputs[1732] = (layer0_outputs[10937]) & (layer0_outputs[7354]);
    assign layer1_outputs[1733] = (layer0_outputs[12719]) & (layer0_outputs[7107]);
    assign layer1_outputs[1734] = ~(layer0_outputs[4496]);
    assign layer1_outputs[1735] = ~(layer0_outputs[10632]) | (layer0_outputs[2367]);
    assign layer1_outputs[1736] = ~(layer0_outputs[2152]);
    assign layer1_outputs[1737] = layer0_outputs[7923];
    assign layer1_outputs[1738] = ~(layer0_outputs[10796]);
    assign layer1_outputs[1739] = ~((layer0_outputs[7883]) | (layer0_outputs[972]));
    assign layer1_outputs[1740] = ~((layer0_outputs[11378]) | (layer0_outputs[9935]));
    assign layer1_outputs[1741] = ~((layer0_outputs[8523]) | (layer0_outputs[2200]));
    assign layer1_outputs[1742] = ~(layer0_outputs[3662]);
    assign layer1_outputs[1743] = ~(layer0_outputs[1026]);
    assign layer1_outputs[1744] = layer0_outputs[11927];
    assign layer1_outputs[1745] = ~(layer0_outputs[2778]) | (layer0_outputs[12470]);
    assign layer1_outputs[1746] = layer0_outputs[7499];
    assign layer1_outputs[1747] = ~(layer0_outputs[11709]);
    assign layer1_outputs[1748] = ~((layer0_outputs[9683]) ^ (layer0_outputs[2000]));
    assign layer1_outputs[1749] = ~((layer0_outputs[762]) ^ (layer0_outputs[5511]));
    assign layer1_outputs[1750] = (layer0_outputs[4674]) & (layer0_outputs[2795]);
    assign layer1_outputs[1751] = (layer0_outputs[9582]) & ~(layer0_outputs[6]);
    assign layer1_outputs[1752] = ~(layer0_outputs[5108]) | (layer0_outputs[9042]);
    assign layer1_outputs[1753] = ~(layer0_outputs[2499]) | (layer0_outputs[8897]);
    assign layer1_outputs[1754] = layer0_outputs[1302];
    assign layer1_outputs[1755] = ~(layer0_outputs[6203]);
    assign layer1_outputs[1756] = ~(layer0_outputs[1795]);
    assign layer1_outputs[1757] = ~((layer0_outputs[11584]) ^ (layer0_outputs[574]));
    assign layer1_outputs[1758] = (layer0_outputs[4412]) & ~(layer0_outputs[4714]);
    assign layer1_outputs[1759] = (layer0_outputs[3181]) & ~(layer0_outputs[10981]);
    assign layer1_outputs[1760] = ~((layer0_outputs[12634]) ^ (layer0_outputs[989]));
    assign layer1_outputs[1761] = ~((layer0_outputs[8950]) & (layer0_outputs[9832]));
    assign layer1_outputs[1762] = ~((layer0_outputs[7549]) ^ (layer0_outputs[9703]));
    assign layer1_outputs[1763] = (layer0_outputs[9535]) & ~(layer0_outputs[8213]);
    assign layer1_outputs[1764] = ~(layer0_outputs[6530]) | (layer0_outputs[7010]);
    assign layer1_outputs[1765] = layer0_outputs[599];
    assign layer1_outputs[1766] = ~(layer0_outputs[8967]) | (layer0_outputs[5044]);
    assign layer1_outputs[1767] = ~(layer0_outputs[3135]) | (layer0_outputs[8562]);
    assign layer1_outputs[1768] = layer0_outputs[9066];
    assign layer1_outputs[1769] = ~(layer0_outputs[5638]) | (layer0_outputs[107]);
    assign layer1_outputs[1770] = ~(layer0_outputs[4152]);
    assign layer1_outputs[1771] = ~(layer0_outputs[6030]) | (layer0_outputs[3741]);
    assign layer1_outputs[1772] = (layer0_outputs[4428]) & (layer0_outputs[11961]);
    assign layer1_outputs[1773] = ~((layer0_outputs[11710]) | (layer0_outputs[8883]));
    assign layer1_outputs[1774] = (layer0_outputs[2229]) | (layer0_outputs[3785]);
    assign layer1_outputs[1775] = ~(layer0_outputs[1060]);
    assign layer1_outputs[1776] = ~((layer0_outputs[12273]) ^ (layer0_outputs[1851]));
    assign layer1_outputs[1777] = layer0_outputs[8840];
    assign layer1_outputs[1778] = ~(layer0_outputs[5512]);
    assign layer1_outputs[1779] = ~((layer0_outputs[880]) | (layer0_outputs[7525]));
    assign layer1_outputs[1780] = 1'b1;
    assign layer1_outputs[1781] = layer0_outputs[4137];
    assign layer1_outputs[1782] = (layer0_outputs[1844]) & ~(layer0_outputs[11127]);
    assign layer1_outputs[1783] = (layer0_outputs[2672]) | (layer0_outputs[331]);
    assign layer1_outputs[1784] = (layer0_outputs[510]) | (layer0_outputs[1099]);
    assign layer1_outputs[1785] = (layer0_outputs[1755]) & ~(layer0_outputs[11774]);
    assign layer1_outputs[1786] = ~((layer0_outputs[8326]) ^ (layer0_outputs[10257]));
    assign layer1_outputs[1787] = (layer0_outputs[5270]) | (layer0_outputs[5095]);
    assign layer1_outputs[1788] = ~(layer0_outputs[3883]) | (layer0_outputs[8119]);
    assign layer1_outputs[1789] = ~(layer0_outputs[12118]);
    assign layer1_outputs[1790] = ~(layer0_outputs[173]);
    assign layer1_outputs[1791] = ~((layer0_outputs[2980]) ^ (layer0_outputs[12321]));
    assign layer1_outputs[1792] = layer0_outputs[7215];
    assign layer1_outputs[1793] = ~((layer0_outputs[9012]) | (layer0_outputs[5934]));
    assign layer1_outputs[1794] = layer0_outputs[981];
    assign layer1_outputs[1795] = (layer0_outputs[5689]) ^ (layer0_outputs[4878]);
    assign layer1_outputs[1796] = ~(layer0_outputs[10625]);
    assign layer1_outputs[1797] = ~((layer0_outputs[8394]) & (layer0_outputs[7114]));
    assign layer1_outputs[1798] = ~(layer0_outputs[6018]);
    assign layer1_outputs[1799] = ~(layer0_outputs[6013]);
    assign layer1_outputs[1800] = ~(layer0_outputs[6723]);
    assign layer1_outputs[1801] = ~((layer0_outputs[11834]) ^ (layer0_outputs[4137]));
    assign layer1_outputs[1802] = (layer0_outputs[5413]) & (layer0_outputs[11856]);
    assign layer1_outputs[1803] = ~((layer0_outputs[4692]) & (layer0_outputs[10077]));
    assign layer1_outputs[1804] = ~(layer0_outputs[3014]);
    assign layer1_outputs[1805] = (layer0_outputs[10073]) & ~(layer0_outputs[6655]);
    assign layer1_outputs[1806] = (layer0_outputs[10009]) & ~(layer0_outputs[8953]);
    assign layer1_outputs[1807] = ~(layer0_outputs[10921]);
    assign layer1_outputs[1808] = (layer0_outputs[11187]) & (layer0_outputs[10224]);
    assign layer1_outputs[1809] = (layer0_outputs[6877]) & ~(layer0_outputs[2017]);
    assign layer1_outputs[1810] = layer0_outputs[2271];
    assign layer1_outputs[1811] = ~(layer0_outputs[3726]);
    assign layer1_outputs[1812] = (layer0_outputs[6884]) ^ (layer0_outputs[951]);
    assign layer1_outputs[1813] = ~(layer0_outputs[2115]);
    assign layer1_outputs[1814] = (layer0_outputs[8752]) & (layer0_outputs[8505]);
    assign layer1_outputs[1815] = ~((layer0_outputs[9885]) & (layer0_outputs[11797]));
    assign layer1_outputs[1816] = ~(layer0_outputs[620]);
    assign layer1_outputs[1817] = ~((layer0_outputs[672]) ^ (layer0_outputs[198]));
    assign layer1_outputs[1818] = (layer0_outputs[7998]) & (layer0_outputs[9363]);
    assign layer1_outputs[1819] = layer0_outputs[2955];
    assign layer1_outputs[1820] = (layer0_outputs[2473]) | (layer0_outputs[6870]);
    assign layer1_outputs[1821] = (layer0_outputs[4775]) & (layer0_outputs[2213]);
    assign layer1_outputs[1822] = layer0_outputs[12303];
    assign layer1_outputs[1823] = ~((layer0_outputs[11899]) ^ (layer0_outputs[7355]));
    assign layer1_outputs[1824] = layer0_outputs[2176];
    assign layer1_outputs[1825] = ~((layer0_outputs[7486]) ^ (layer0_outputs[2117]));
    assign layer1_outputs[1826] = (layer0_outputs[5348]) | (layer0_outputs[8408]);
    assign layer1_outputs[1827] = ~(layer0_outputs[10544]);
    assign layer1_outputs[1828] = (layer0_outputs[2289]) | (layer0_outputs[8290]);
    assign layer1_outputs[1829] = (layer0_outputs[7534]) | (layer0_outputs[7414]);
    assign layer1_outputs[1830] = layer0_outputs[12372];
    assign layer1_outputs[1831] = layer0_outputs[1199];
    assign layer1_outputs[1832] = layer0_outputs[25];
    assign layer1_outputs[1833] = (layer0_outputs[2594]) & ~(layer0_outputs[506]);
    assign layer1_outputs[1834] = (layer0_outputs[5684]) & ~(layer0_outputs[707]);
    assign layer1_outputs[1835] = ~((layer0_outputs[11033]) ^ (layer0_outputs[2027]));
    assign layer1_outputs[1836] = ~(layer0_outputs[6085]) | (layer0_outputs[9422]);
    assign layer1_outputs[1837] = (layer0_outputs[4449]) & ~(layer0_outputs[5170]);
    assign layer1_outputs[1838] = ~(layer0_outputs[7610]);
    assign layer1_outputs[1839] = (layer0_outputs[9655]) & ~(layer0_outputs[3841]);
    assign layer1_outputs[1840] = layer0_outputs[1622];
    assign layer1_outputs[1841] = ~((layer0_outputs[11816]) ^ (layer0_outputs[10324]));
    assign layer1_outputs[1842] = layer0_outputs[3996];
    assign layer1_outputs[1843] = ~(layer0_outputs[2381]);
    assign layer1_outputs[1844] = ~(layer0_outputs[6708]);
    assign layer1_outputs[1845] = (layer0_outputs[12715]) ^ (layer0_outputs[6251]);
    assign layer1_outputs[1846] = layer0_outputs[2738];
    assign layer1_outputs[1847] = (layer0_outputs[6874]) ^ (layer0_outputs[10458]);
    assign layer1_outputs[1848] = layer0_outputs[5700];
    assign layer1_outputs[1849] = layer0_outputs[6596];
    assign layer1_outputs[1850] = (layer0_outputs[2521]) | (layer0_outputs[7372]);
    assign layer1_outputs[1851] = (layer0_outputs[2295]) & ~(layer0_outputs[12627]);
    assign layer1_outputs[1852] = (layer0_outputs[4623]) | (layer0_outputs[1651]);
    assign layer1_outputs[1853] = ~(layer0_outputs[3154]);
    assign layer1_outputs[1854] = (layer0_outputs[5862]) & ~(layer0_outputs[1131]);
    assign layer1_outputs[1855] = 1'b1;
    assign layer1_outputs[1856] = ~(layer0_outputs[2888]);
    assign layer1_outputs[1857] = ~(layer0_outputs[8932]) | (layer0_outputs[9077]);
    assign layer1_outputs[1858] = ~(layer0_outputs[1094]);
    assign layer1_outputs[1859] = layer0_outputs[540];
    assign layer1_outputs[1860] = ~(layer0_outputs[2268]) | (layer0_outputs[5840]);
    assign layer1_outputs[1861] = ~((layer0_outputs[7024]) & (layer0_outputs[10178]));
    assign layer1_outputs[1862] = ~(layer0_outputs[10187]) | (layer0_outputs[1101]);
    assign layer1_outputs[1863] = (layer0_outputs[11407]) & (layer0_outputs[11549]);
    assign layer1_outputs[1864] = 1'b0;
    assign layer1_outputs[1865] = (layer0_outputs[11339]) & (layer0_outputs[8536]);
    assign layer1_outputs[1866] = ~((layer0_outputs[11317]) | (layer0_outputs[6883]));
    assign layer1_outputs[1867] = layer0_outputs[3248];
    assign layer1_outputs[1868] = (layer0_outputs[11699]) & ~(layer0_outputs[2009]);
    assign layer1_outputs[1869] = ~((layer0_outputs[5012]) ^ (layer0_outputs[8551]));
    assign layer1_outputs[1870] = (layer0_outputs[2260]) | (layer0_outputs[11237]);
    assign layer1_outputs[1871] = ~(layer0_outputs[3094]);
    assign layer1_outputs[1872] = ~(layer0_outputs[3273]);
    assign layer1_outputs[1873] = (layer0_outputs[1081]) & ~(layer0_outputs[7779]);
    assign layer1_outputs[1874] = ~(layer0_outputs[12712]);
    assign layer1_outputs[1875] = ~((layer0_outputs[2306]) ^ (layer0_outputs[10859]));
    assign layer1_outputs[1876] = (layer0_outputs[9089]) | (layer0_outputs[5765]);
    assign layer1_outputs[1877] = ~(layer0_outputs[2224]);
    assign layer1_outputs[1878] = layer0_outputs[5587];
    assign layer1_outputs[1879] = ~(layer0_outputs[3965]) | (layer0_outputs[9997]);
    assign layer1_outputs[1880] = (layer0_outputs[5711]) & ~(layer0_outputs[356]);
    assign layer1_outputs[1881] = ~((layer0_outputs[9870]) & (layer0_outputs[6039]));
    assign layer1_outputs[1882] = (layer0_outputs[180]) & ~(layer0_outputs[8568]);
    assign layer1_outputs[1883] = layer0_outputs[6765];
    assign layer1_outputs[1884] = 1'b0;
    assign layer1_outputs[1885] = ~(layer0_outputs[1682]);
    assign layer1_outputs[1886] = ~(layer0_outputs[2944]) | (layer0_outputs[11648]);
    assign layer1_outputs[1887] = ~(layer0_outputs[2960]);
    assign layer1_outputs[1888] = ~((layer0_outputs[9951]) ^ (layer0_outputs[2780]));
    assign layer1_outputs[1889] = ~(layer0_outputs[11836]);
    assign layer1_outputs[1890] = ~(layer0_outputs[11384]);
    assign layer1_outputs[1891] = (layer0_outputs[1327]) ^ (layer0_outputs[4214]);
    assign layer1_outputs[1892] = ~((layer0_outputs[688]) ^ (layer0_outputs[5062]));
    assign layer1_outputs[1893] = layer0_outputs[9706];
    assign layer1_outputs[1894] = ~((layer0_outputs[9805]) | (layer0_outputs[3645]));
    assign layer1_outputs[1895] = ~(layer0_outputs[9166]);
    assign layer1_outputs[1896] = ~((layer0_outputs[11943]) ^ (layer0_outputs[7411]));
    assign layer1_outputs[1897] = ~(layer0_outputs[8325]);
    assign layer1_outputs[1898] = layer0_outputs[4952];
    assign layer1_outputs[1899] = ~(layer0_outputs[4619]);
    assign layer1_outputs[1900] = ~(layer0_outputs[6406]);
    assign layer1_outputs[1901] = (layer0_outputs[9114]) & ~(layer0_outputs[111]);
    assign layer1_outputs[1902] = layer0_outputs[11507];
    assign layer1_outputs[1903] = layer0_outputs[439];
    assign layer1_outputs[1904] = (layer0_outputs[3265]) & (layer0_outputs[6098]);
    assign layer1_outputs[1905] = layer0_outputs[110];
    assign layer1_outputs[1906] = ~((layer0_outputs[10604]) & (layer0_outputs[10940]));
    assign layer1_outputs[1907] = (layer0_outputs[1838]) & ~(layer0_outputs[7830]);
    assign layer1_outputs[1908] = ~(layer0_outputs[10328]);
    assign layer1_outputs[1909] = ~(layer0_outputs[2004]);
    assign layer1_outputs[1910] = (layer0_outputs[3603]) & (layer0_outputs[6140]);
    assign layer1_outputs[1911] = layer0_outputs[7235];
    assign layer1_outputs[1912] = ~(layer0_outputs[2041]);
    assign layer1_outputs[1913] = ~(layer0_outputs[9873]) | (layer0_outputs[4893]);
    assign layer1_outputs[1914] = layer0_outputs[10628];
    assign layer1_outputs[1915] = layer0_outputs[8142];
    assign layer1_outputs[1916] = ~(layer0_outputs[11578]);
    assign layer1_outputs[1917] = ~(layer0_outputs[10964]);
    assign layer1_outputs[1918] = (layer0_outputs[9560]) & ~(layer0_outputs[12569]);
    assign layer1_outputs[1919] = ~(layer0_outputs[9271]);
    assign layer1_outputs[1920] = ~((layer0_outputs[7907]) ^ (layer0_outputs[8494]));
    assign layer1_outputs[1921] = ~(layer0_outputs[11881]);
    assign layer1_outputs[1922] = ~(layer0_outputs[165]);
    assign layer1_outputs[1923] = ~((layer0_outputs[5421]) | (layer0_outputs[4212]));
    assign layer1_outputs[1924] = (layer0_outputs[6727]) ^ (layer0_outputs[12781]);
    assign layer1_outputs[1925] = layer0_outputs[4412];
    assign layer1_outputs[1926] = (layer0_outputs[7859]) | (layer0_outputs[11252]);
    assign layer1_outputs[1927] = (layer0_outputs[307]) & ~(layer0_outputs[4992]);
    assign layer1_outputs[1928] = ~(layer0_outputs[9950]);
    assign layer1_outputs[1929] = ~(layer0_outputs[10105]) | (layer0_outputs[2377]);
    assign layer1_outputs[1930] = ~(layer0_outputs[7561]);
    assign layer1_outputs[1931] = 1'b1;
    assign layer1_outputs[1932] = (layer0_outputs[7262]) & (layer0_outputs[6999]);
    assign layer1_outputs[1933] = ~(layer0_outputs[7376]);
    assign layer1_outputs[1934] = 1'b0;
    assign layer1_outputs[1935] = ~(layer0_outputs[10597]) | (layer0_outputs[6026]);
    assign layer1_outputs[1936] = layer0_outputs[7981];
    assign layer1_outputs[1937] = layer0_outputs[2595];
    assign layer1_outputs[1938] = layer0_outputs[8893];
    assign layer1_outputs[1939] = ~(layer0_outputs[9248]);
    assign layer1_outputs[1940] = ~(layer0_outputs[1601]) | (layer0_outputs[12247]);
    assign layer1_outputs[1941] = layer0_outputs[6878];
    assign layer1_outputs[1942] = ~(layer0_outputs[1422]);
    assign layer1_outputs[1943] = ~(layer0_outputs[3978]) | (layer0_outputs[7806]);
    assign layer1_outputs[1944] = ~(layer0_outputs[9778]);
    assign layer1_outputs[1945] = layer0_outputs[10695];
    assign layer1_outputs[1946] = layer0_outputs[3180];
    assign layer1_outputs[1947] = ~(layer0_outputs[1900]);
    assign layer1_outputs[1948] = (layer0_outputs[7351]) ^ (layer0_outputs[6820]);
    assign layer1_outputs[1949] = layer0_outputs[12285];
    assign layer1_outputs[1950] = (layer0_outputs[3852]) | (layer0_outputs[171]);
    assign layer1_outputs[1951] = (layer0_outputs[1899]) | (layer0_outputs[8085]);
    assign layer1_outputs[1952] = layer0_outputs[3511];
    assign layer1_outputs[1953] = ~(layer0_outputs[7593]) | (layer0_outputs[10607]);
    assign layer1_outputs[1954] = (layer0_outputs[2619]) & (layer0_outputs[10145]);
    assign layer1_outputs[1955] = (layer0_outputs[9828]) ^ (layer0_outputs[12615]);
    assign layer1_outputs[1956] = (layer0_outputs[12126]) & ~(layer0_outputs[6921]);
    assign layer1_outputs[1957] = ~(layer0_outputs[8694]);
    assign layer1_outputs[1958] = ~(layer0_outputs[4377]) | (layer0_outputs[2160]);
    assign layer1_outputs[1959] = (layer0_outputs[9879]) ^ (layer0_outputs[7056]);
    assign layer1_outputs[1960] = ~((layer0_outputs[11743]) | (layer0_outputs[7360]));
    assign layer1_outputs[1961] = ~(layer0_outputs[11603]);
    assign layer1_outputs[1962] = ~(layer0_outputs[5253]) | (layer0_outputs[8710]);
    assign layer1_outputs[1963] = ~(layer0_outputs[12689]);
    assign layer1_outputs[1964] = (layer0_outputs[7345]) & (layer0_outputs[209]);
    assign layer1_outputs[1965] = ~(layer0_outputs[1670]);
    assign layer1_outputs[1966] = ~(layer0_outputs[9978]) | (layer0_outputs[5741]);
    assign layer1_outputs[1967] = ~((layer0_outputs[2083]) & (layer0_outputs[3228]));
    assign layer1_outputs[1968] = ~(layer0_outputs[2102]);
    assign layer1_outputs[1969] = ~(layer0_outputs[1848]);
    assign layer1_outputs[1970] = ~(layer0_outputs[12248]);
    assign layer1_outputs[1971] = layer0_outputs[12651];
    assign layer1_outputs[1972] = ~(layer0_outputs[3398]);
    assign layer1_outputs[1973] = ~((layer0_outputs[3927]) ^ (layer0_outputs[6372]));
    assign layer1_outputs[1974] = layer0_outputs[6471];
    assign layer1_outputs[1975] = ~((layer0_outputs[1065]) & (layer0_outputs[3320]));
    assign layer1_outputs[1976] = ~(layer0_outputs[12467]);
    assign layer1_outputs[1977] = (layer0_outputs[1088]) & ~(layer0_outputs[116]);
    assign layer1_outputs[1978] = ~(layer0_outputs[413]);
    assign layer1_outputs[1979] = (layer0_outputs[6515]) & ~(layer0_outputs[11447]);
    assign layer1_outputs[1980] = ~(layer0_outputs[5811]) | (layer0_outputs[921]);
    assign layer1_outputs[1981] = layer0_outputs[4477];
    assign layer1_outputs[1982] = (layer0_outputs[3175]) | (layer0_outputs[10930]);
    assign layer1_outputs[1983] = layer0_outputs[4549];
    assign layer1_outputs[1984] = ~(layer0_outputs[9745]);
    assign layer1_outputs[1985] = ~(layer0_outputs[2720]) | (layer0_outputs[4743]);
    assign layer1_outputs[1986] = ~((layer0_outputs[10426]) | (layer0_outputs[10988]));
    assign layer1_outputs[1987] = layer0_outputs[5292];
    assign layer1_outputs[1988] = layer0_outputs[7988];
    assign layer1_outputs[1989] = ~((layer0_outputs[8346]) & (layer0_outputs[2448]));
    assign layer1_outputs[1990] = (layer0_outputs[277]) & ~(layer0_outputs[5781]);
    assign layer1_outputs[1991] = (layer0_outputs[458]) ^ (layer0_outputs[6081]);
    assign layer1_outputs[1992] = layer0_outputs[11080];
    assign layer1_outputs[1993] = ~((layer0_outputs[11318]) & (layer0_outputs[993]));
    assign layer1_outputs[1994] = ~((layer0_outputs[5182]) ^ (layer0_outputs[7618]));
    assign layer1_outputs[1995] = ~(layer0_outputs[10233]) | (layer0_outputs[12752]);
    assign layer1_outputs[1996] = (layer0_outputs[11193]) & ~(layer0_outputs[9306]);
    assign layer1_outputs[1997] = (layer0_outputs[7294]) ^ (layer0_outputs[7703]);
    assign layer1_outputs[1998] = ~(layer0_outputs[5319]);
    assign layer1_outputs[1999] = ~((layer0_outputs[6158]) | (layer0_outputs[9196]));
    assign layer1_outputs[2000] = ~(layer0_outputs[12431]);
    assign layer1_outputs[2001] = layer0_outputs[9130];
    assign layer1_outputs[2002] = ~(layer0_outputs[7160]);
    assign layer1_outputs[2003] = (layer0_outputs[3839]) & (layer0_outputs[6600]);
    assign layer1_outputs[2004] = (layer0_outputs[2271]) | (layer0_outputs[8028]);
    assign layer1_outputs[2005] = layer0_outputs[6858];
    assign layer1_outputs[2006] = ~((layer0_outputs[12539]) & (layer0_outputs[4724]));
    assign layer1_outputs[2007] = ~(layer0_outputs[7113]);
    assign layer1_outputs[2008] = (layer0_outputs[6663]) ^ (layer0_outputs[2441]);
    assign layer1_outputs[2009] = ~((layer0_outputs[12270]) & (layer0_outputs[4007]));
    assign layer1_outputs[2010] = ~(layer0_outputs[8128]) | (layer0_outputs[9525]);
    assign layer1_outputs[2011] = layer0_outputs[4100];
    assign layer1_outputs[2012] = (layer0_outputs[6537]) ^ (layer0_outputs[9305]);
    assign layer1_outputs[2013] = ~(layer0_outputs[3407]);
    assign layer1_outputs[2014] = (layer0_outputs[2368]) | (layer0_outputs[4813]);
    assign layer1_outputs[2015] = (layer0_outputs[6887]) | (layer0_outputs[1991]);
    assign layer1_outputs[2016] = ~((layer0_outputs[12138]) ^ (layer0_outputs[9550]));
    assign layer1_outputs[2017] = ~(layer0_outputs[5508]);
    assign layer1_outputs[2018] = ~(layer0_outputs[6648]) | (layer0_outputs[10350]);
    assign layer1_outputs[2019] = layer0_outputs[5056];
    assign layer1_outputs[2020] = ~(layer0_outputs[9933]);
    assign layer1_outputs[2021] = ~((layer0_outputs[3816]) ^ (layer0_outputs[2184]));
    assign layer1_outputs[2022] = ~((layer0_outputs[8993]) ^ (layer0_outputs[3291]));
    assign layer1_outputs[2023] = layer0_outputs[11958];
    assign layer1_outputs[2024] = layer0_outputs[12747];
    assign layer1_outputs[2025] = (layer0_outputs[11993]) | (layer0_outputs[7063]);
    assign layer1_outputs[2026] = ~(layer0_outputs[7094]);
    assign layer1_outputs[2027] = layer0_outputs[10093];
    assign layer1_outputs[2028] = ~((layer0_outputs[10196]) & (layer0_outputs[774]));
    assign layer1_outputs[2029] = (layer0_outputs[689]) | (layer0_outputs[11876]);
    assign layer1_outputs[2030] = (layer0_outputs[5828]) & (layer0_outputs[5631]);
    assign layer1_outputs[2031] = ~(layer0_outputs[188]);
    assign layer1_outputs[2032] = (layer0_outputs[9047]) | (layer0_outputs[3491]);
    assign layer1_outputs[2033] = ~(layer0_outputs[3399]);
    assign layer1_outputs[2034] = ~(layer0_outputs[11211]) | (layer0_outputs[2546]);
    assign layer1_outputs[2035] = ~(layer0_outputs[571]) | (layer0_outputs[3682]);
    assign layer1_outputs[2036] = (layer0_outputs[8866]) & ~(layer0_outputs[9406]);
    assign layer1_outputs[2037] = (layer0_outputs[3820]) & ~(layer0_outputs[1708]);
    assign layer1_outputs[2038] = 1'b0;
    assign layer1_outputs[2039] = layer0_outputs[4850];
    assign layer1_outputs[2040] = ~(layer0_outputs[5872]) | (layer0_outputs[12201]);
    assign layer1_outputs[2041] = (layer0_outputs[5966]) & ~(layer0_outputs[12094]);
    assign layer1_outputs[2042] = ~((layer0_outputs[6388]) | (layer0_outputs[7217]));
    assign layer1_outputs[2043] = (layer0_outputs[3380]) & (layer0_outputs[5368]);
    assign layer1_outputs[2044] = layer0_outputs[1776];
    assign layer1_outputs[2045] = ~(layer0_outputs[9709]);
    assign layer1_outputs[2046] = ~(layer0_outputs[12046]) | (layer0_outputs[5553]);
    assign layer1_outputs[2047] = ~(layer0_outputs[5703]);
    assign layer1_outputs[2048] = layer0_outputs[9456];
    assign layer1_outputs[2049] = layer0_outputs[5771];
    assign layer1_outputs[2050] = ~((layer0_outputs[6945]) | (layer0_outputs[11031]));
    assign layer1_outputs[2051] = ~(layer0_outputs[3900]) | (layer0_outputs[9854]);
    assign layer1_outputs[2052] = (layer0_outputs[4826]) & ~(layer0_outputs[506]);
    assign layer1_outputs[2053] = ~(layer0_outputs[28]);
    assign layer1_outputs[2054] = (layer0_outputs[535]) & (layer0_outputs[5907]);
    assign layer1_outputs[2055] = ~((layer0_outputs[2616]) | (layer0_outputs[8812]));
    assign layer1_outputs[2056] = ~(layer0_outputs[10034]);
    assign layer1_outputs[2057] = ~(layer0_outputs[10968]);
    assign layer1_outputs[2058] = 1'b1;
    assign layer1_outputs[2059] = layer0_outputs[6706];
    assign layer1_outputs[2060] = (layer0_outputs[2911]) & ~(layer0_outputs[9903]);
    assign layer1_outputs[2061] = ~(layer0_outputs[609]) | (layer0_outputs[4577]);
    assign layer1_outputs[2062] = (layer0_outputs[3443]) & ~(layer0_outputs[10997]);
    assign layer1_outputs[2063] = ~(layer0_outputs[11833]) | (layer0_outputs[1280]);
    assign layer1_outputs[2064] = (layer0_outputs[8965]) & (layer0_outputs[3275]);
    assign layer1_outputs[2065] = (layer0_outputs[5696]) | (layer0_outputs[8595]);
    assign layer1_outputs[2066] = (layer0_outputs[2891]) & ~(layer0_outputs[10579]);
    assign layer1_outputs[2067] = layer0_outputs[11110];
    assign layer1_outputs[2068] = (layer0_outputs[5303]) & ~(layer0_outputs[1036]);
    assign layer1_outputs[2069] = 1'b1;
    assign layer1_outputs[2070] = 1'b0;
    assign layer1_outputs[2071] = ~((layer0_outputs[5984]) ^ (layer0_outputs[12695]));
    assign layer1_outputs[2072] = ~(layer0_outputs[12086]);
    assign layer1_outputs[2073] = ~(layer0_outputs[11979]);
    assign layer1_outputs[2074] = (layer0_outputs[7148]) & ~(layer0_outputs[5700]);
    assign layer1_outputs[2075] = ~((layer0_outputs[10144]) | (layer0_outputs[5032]));
    assign layer1_outputs[2076] = 1'b0;
    assign layer1_outputs[2077] = ~((layer0_outputs[12733]) | (layer0_outputs[5885]));
    assign layer1_outputs[2078] = ~(layer0_outputs[573]) | (layer0_outputs[9691]);
    assign layer1_outputs[2079] = ~(layer0_outputs[12722]) | (layer0_outputs[5471]);
    assign layer1_outputs[2080] = ~(layer0_outputs[11561]) | (layer0_outputs[6729]);
    assign layer1_outputs[2081] = (layer0_outputs[8293]) ^ (layer0_outputs[8730]);
    assign layer1_outputs[2082] = ~(layer0_outputs[5772]) | (layer0_outputs[12473]);
    assign layer1_outputs[2083] = layer0_outputs[11323];
    assign layer1_outputs[2084] = layer0_outputs[11853];
    assign layer1_outputs[2085] = ~(layer0_outputs[447]);
    assign layer1_outputs[2086] = layer0_outputs[3847];
    assign layer1_outputs[2087] = ~((layer0_outputs[9170]) | (layer0_outputs[5427]));
    assign layer1_outputs[2088] = (layer0_outputs[9914]) & ~(layer0_outputs[1131]);
    assign layer1_outputs[2089] = (layer0_outputs[7707]) ^ (layer0_outputs[4450]);
    assign layer1_outputs[2090] = (layer0_outputs[553]) & (layer0_outputs[12310]);
    assign layer1_outputs[2091] = ~((layer0_outputs[4745]) | (layer0_outputs[8534]));
    assign layer1_outputs[2092] = ~(layer0_outputs[2421]) | (layer0_outputs[3574]);
    assign layer1_outputs[2093] = ~(layer0_outputs[5780]) | (layer0_outputs[378]);
    assign layer1_outputs[2094] = ~((layer0_outputs[12717]) & (layer0_outputs[1757]));
    assign layer1_outputs[2095] = ~(layer0_outputs[9235]) | (layer0_outputs[6943]);
    assign layer1_outputs[2096] = ~(layer0_outputs[8532]);
    assign layer1_outputs[2097] = (layer0_outputs[4661]) ^ (layer0_outputs[2896]);
    assign layer1_outputs[2098] = ~(layer0_outputs[12688]) | (layer0_outputs[1347]);
    assign layer1_outputs[2099] = ~(layer0_outputs[2456]) | (layer0_outputs[1444]);
    assign layer1_outputs[2100] = ~(layer0_outputs[3126]);
    assign layer1_outputs[2101] = layer0_outputs[1147];
    assign layer1_outputs[2102] = ~(layer0_outputs[2460]) | (layer0_outputs[8516]);
    assign layer1_outputs[2103] = layer0_outputs[5026];
    assign layer1_outputs[2104] = ~(layer0_outputs[5352]);
    assign layer1_outputs[2105] = ~(layer0_outputs[3418]);
    assign layer1_outputs[2106] = 1'b0;
    assign layer1_outputs[2107] = layer0_outputs[6919];
    assign layer1_outputs[2108] = ~(layer0_outputs[492]) | (layer0_outputs[5165]);
    assign layer1_outputs[2109] = layer0_outputs[7925];
    assign layer1_outputs[2110] = layer0_outputs[5637];
    assign layer1_outputs[2111] = (layer0_outputs[12436]) & ~(layer0_outputs[5455]);
    assign layer1_outputs[2112] = layer0_outputs[10133];
    assign layer1_outputs[2113] = ~(layer0_outputs[8482]);
    assign layer1_outputs[2114] = 1'b1;
    assign layer1_outputs[2115] = ~((layer0_outputs[1273]) | (layer0_outputs[1428]));
    assign layer1_outputs[2116] = ~(layer0_outputs[11673]);
    assign layer1_outputs[2117] = ~(layer0_outputs[9389]);
    assign layer1_outputs[2118] = layer0_outputs[4793];
    assign layer1_outputs[2119] = ~(layer0_outputs[10068]) | (layer0_outputs[3349]);
    assign layer1_outputs[2120] = (layer0_outputs[11569]) & ~(layer0_outputs[12268]);
    assign layer1_outputs[2121] = layer0_outputs[10285];
    assign layer1_outputs[2122] = (layer0_outputs[1596]) | (layer0_outputs[3936]);
    assign layer1_outputs[2123] = ~(layer0_outputs[8783]) | (layer0_outputs[6342]);
    assign layer1_outputs[2124] = (layer0_outputs[5263]) & ~(layer0_outputs[4743]);
    assign layer1_outputs[2125] = (layer0_outputs[6843]) & (layer0_outputs[3583]);
    assign layer1_outputs[2126] = ~(layer0_outputs[720]) | (layer0_outputs[10512]);
    assign layer1_outputs[2127] = layer0_outputs[9487];
    assign layer1_outputs[2128] = ~(layer0_outputs[2016]);
    assign layer1_outputs[2129] = ~((layer0_outputs[733]) ^ (layer0_outputs[746]));
    assign layer1_outputs[2130] = (layer0_outputs[12738]) & ~(layer0_outputs[8841]);
    assign layer1_outputs[2131] = layer0_outputs[250];
    assign layer1_outputs[2132] = (layer0_outputs[6265]) ^ (layer0_outputs[9597]);
    assign layer1_outputs[2133] = layer0_outputs[39];
    assign layer1_outputs[2134] = ~(layer0_outputs[6866]);
    assign layer1_outputs[2135] = ~(layer0_outputs[11516]);
    assign layer1_outputs[2136] = ~(layer0_outputs[10964]) | (layer0_outputs[4369]);
    assign layer1_outputs[2137] = (layer0_outputs[6576]) & ~(layer0_outputs[8557]);
    assign layer1_outputs[2138] = layer0_outputs[558];
    assign layer1_outputs[2139] = (layer0_outputs[289]) | (layer0_outputs[2204]);
    assign layer1_outputs[2140] = layer0_outputs[6118];
    assign layer1_outputs[2141] = layer0_outputs[1047];
    assign layer1_outputs[2142] = (layer0_outputs[2289]) & (layer0_outputs[45]);
    assign layer1_outputs[2143] = ~(layer0_outputs[454]);
    assign layer1_outputs[2144] = layer0_outputs[4915];
    assign layer1_outputs[2145] = layer0_outputs[2692];
    assign layer1_outputs[2146] = ~(layer0_outputs[2064]);
    assign layer1_outputs[2147] = ~(layer0_outputs[1212]) | (layer0_outputs[5423]);
    assign layer1_outputs[2148] = ~((layer0_outputs[6502]) ^ (layer0_outputs[5373]));
    assign layer1_outputs[2149] = (layer0_outputs[4758]) & ~(layer0_outputs[10008]);
    assign layer1_outputs[2150] = ~(layer0_outputs[9959]) | (layer0_outputs[1964]);
    assign layer1_outputs[2151] = ~(layer0_outputs[9544]);
    assign layer1_outputs[2152] = (layer0_outputs[1465]) | (layer0_outputs[10223]);
    assign layer1_outputs[2153] = (layer0_outputs[1572]) | (layer0_outputs[8790]);
    assign layer1_outputs[2154] = (layer0_outputs[5963]) & ~(layer0_outputs[2446]);
    assign layer1_outputs[2155] = (layer0_outputs[5449]) & ~(layer0_outputs[3723]);
    assign layer1_outputs[2156] = ~(layer0_outputs[6238]);
    assign layer1_outputs[2157] = ~((layer0_outputs[11348]) & (layer0_outputs[1193]));
    assign layer1_outputs[2158] = ~((layer0_outputs[6664]) | (layer0_outputs[3739]));
    assign layer1_outputs[2159] = ~((layer0_outputs[11530]) ^ (layer0_outputs[5306]));
    assign layer1_outputs[2160] = ~(layer0_outputs[9313]);
    assign layer1_outputs[2161] = (layer0_outputs[3352]) & ~(layer0_outputs[2230]);
    assign layer1_outputs[2162] = ~(layer0_outputs[5240]);
    assign layer1_outputs[2163] = ~(layer0_outputs[12241]);
    assign layer1_outputs[2164] = (layer0_outputs[2312]) & ~(layer0_outputs[11210]);
    assign layer1_outputs[2165] = layer0_outputs[10995];
    assign layer1_outputs[2166] = (layer0_outputs[7768]) & ~(layer0_outputs[1874]);
    assign layer1_outputs[2167] = ~(layer0_outputs[10401]);
    assign layer1_outputs[2168] = ~(layer0_outputs[1756]);
    assign layer1_outputs[2169] = ~(layer0_outputs[10386]);
    assign layer1_outputs[2170] = (layer0_outputs[3344]) & ~(layer0_outputs[7179]);
    assign layer1_outputs[2171] = ~(layer0_outputs[2190]) | (layer0_outputs[4717]);
    assign layer1_outputs[2172] = (layer0_outputs[6198]) ^ (layer0_outputs[7154]);
    assign layer1_outputs[2173] = layer0_outputs[12727];
    assign layer1_outputs[2174] = (layer0_outputs[12465]) | (layer0_outputs[10687]);
    assign layer1_outputs[2175] = layer0_outputs[1025];
    assign layer1_outputs[2176] = ~(layer0_outputs[1830]);
    assign layer1_outputs[2177] = ~(layer0_outputs[8121]);
    assign layer1_outputs[2178] = ~((layer0_outputs[3083]) ^ (layer0_outputs[1140]));
    assign layer1_outputs[2179] = ~(layer0_outputs[10285]);
    assign layer1_outputs[2180] = layer0_outputs[9579];
    assign layer1_outputs[2181] = layer0_outputs[43];
    assign layer1_outputs[2182] = (layer0_outputs[2838]) & ~(layer0_outputs[7679]);
    assign layer1_outputs[2183] = ~((layer0_outputs[2165]) | (layer0_outputs[3180]));
    assign layer1_outputs[2184] = layer0_outputs[10992];
    assign layer1_outputs[2185] = ~((layer0_outputs[1804]) ^ (layer0_outputs[663]));
    assign layer1_outputs[2186] = ~(layer0_outputs[7913]) | (layer0_outputs[3199]);
    assign layer1_outputs[2187] = ~((layer0_outputs[228]) | (layer0_outputs[1901]));
    assign layer1_outputs[2188] = ~(layer0_outputs[9426]);
    assign layer1_outputs[2189] = ~(layer0_outputs[3163]);
    assign layer1_outputs[2190] = layer0_outputs[1236];
    assign layer1_outputs[2191] = layer0_outputs[10487];
    assign layer1_outputs[2192] = layer0_outputs[12562];
    assign layer1_outputs[2193] = ~((layer0_outputs[9501]) & (layer0_outputs[41]));
    assign layer1_outputs[2194] = ~(layer0_outputs[7697]);
    assign layer1_outputs[2195] = (layer0_outputs[4397]) & ~(layer0_outputs[6493]);
    assign layer1_outputs[2196] = ~(layer0_outputs[12006]);
    assign layer1_outputs[2197] = ~(layer0_outputs[6268]);
    assign layer1_outputs[2198] = layer0_outputs[2655];
    assign layer1_outputs[2199] = ~(layer0_outputs[6523]);
    assign layer1_outputs[2200] = ~((layer0_outputs[4613]) ^ (layer0_outputs[7609]));
    assign layer1_outputs[2201] = ~(layer0_outputs[7917]);
    assign layer1_outputs[2202] = ~(layer0_outputs[8244]) | (layer0_outputs[9895]);
    assign layer1_outputs[2203] = (layer0_outputs[5466]) & ~(layer0_outputs[1869]);
    assign layer1_outputs[2204] = layer0_outputs[12110];
    assign layer1_outputs[2205] = (layer0_outputs[2823]) & ~(layer0_outputs[5810]);
    assign layer1_outputs[2206] = ~(layer0_outputs[11265]);
    assign layer1_outputs[2207] = ~((layer0_outputs[9448]) | (layer0_outputs[5152]));
    assign layer1_outputs[2208] = ~(layer0_outputs[12744]) | (layer0_outputs[4586]);
    assign layer1_outputs[2209] = layer0_outputs[11285];
    assign layer1_outputs[2210] = 1'b1;
    assign layer1_outputs[2211] = (layer0_outputs[2029]) & ~(layer0_outputs[6746]);
    assign layer1_outputs[2212] = layer0_outputs[1985];
    assign layer1_outputs[2213] = ~(layer0_outputs[5016]) | (layer0_outputs[4715]);
    assign layer1_outputs[2214] = (layer0_outputs[11413]) | (layer0_outputs[3008]);
    assign layer1_outputs[2215] = ~((layer0_outputs[7193]) ^ (layer0_outputs[4516]));
    assign layer1_outputs[2216] = layer0_outputs[11239];
    assign layer1_outputs[2217] = ~(layer0_outputs[5043]);
    assign layer1_outputs[2218] = ~(layer0_outputs[12205]);
    assign layer1_outputs[2219] = (layer0_outputs[5510]) & ~(layer0_outputs[2617]);
    assign layer1_outputs[2220] = layer0_outputs[3978];
    assign layer1_outputs[2221] = ~(layer0_outputs[8896]) | (layer0_outputs[3024]);
    assign layer1_outputs[2222] = (layer0_outputs[3261]) ^ (layer0_outputs[12690]);
    assign layer1_outputs[2223] = ~(layer0_outputs[11149]) | (layer0_outputs[9542]);
    assign layer1_outputs[2224] = ~((layer0_outputs[3540]) | (layer0_outputs[2240]));
    assign layer1_outputs[2225] = ~(layer0_outputs[8829]);
    assign layer1_outputs[2226] = ~(layer0_outputs[12725]);
    assign layer1_outputs[2227] = (layer0_outputs[10472]) & ~(layer0_outputs[996]);
    assign layer1_outputs[2228] = (layer0_outputs[5350]) & ~(layer0_outputs[11359]);
    assign layer1_outputs[2229] = layer0_outputs[9650];
    assign layer1_outputs[2230] = (layer0_outputs[12660]) & ~(layer0_outputs[3170]);
    assign layer1_outputs[2231] = (layer0_outputs[8917]) & (layer0_outputs[3301]);
    assign layer1_outputs[2232] = ~(layer0_outputs[9719]) | (layer0_outputs[3101]);
    assign layer1_outputs[2233] = ~(layer0_outputs[7711]) | (layer0_outputs[11970]);
    assign layer1_outputs[2234] = layer0_outputs[4491];
    assign layer1_outputs[2235] = ~(layer0_outputs[2668]) | (layer0_outputs[10238]);
    assign layer1_outputs[2236] = ~((layer0_outputs[12504]) & (layer0_outputs[3886]));
    assign layer1_outputs[2237] = ~((layer0_outputs[6601]) & (layer0_outputs[9934]));
    assign layer1_outputs[2238] = (layer0_outputs[10307]) & ~(layer0_outputs[3621]);
    assign layer1_outputs[2239] = (layer0_outputs[10526]) ^ (layer0_outputs[5719]);
    assign layer1_outputs[2240] = ~((layer0_outputs[10260]) ^ (layer0_outputs[9027]));
    assign layer1_outputs[2241] = layer0_outputs[6653];
    assign layer1_outputs[2242] = layer0_outputs[1336];
    assign layer1_outputs[2243] = (layer0_outputs[5543]) & ~(layer0_outputs[10735]);
    assign layer1_outputs[2244] = ~((layer0_outputs[5856]) & (layer0_outputs[8738]));
    assign layer1_outputs[2245] = ~((layer0_outputs[766]) | (layer0_outputs[1028]));
    assign layer1_outputs[2246] = ~(layer0_outputs[7725]);
    assign layer1_outputs[2247] = (layer0_outputs[9929]) & ~(layer0_outputs[7694]);
    assign layer1_outputs[2248] = layer0_outputs[991];
    assign layer1_outputs[2249] = (layer0_outputs[11060]) & (layer0_outputs[3585]);
    assign layer1_outputs[2250] = ~(layer0_outputs[10639]);
    assign layer1_outputs[2251] = (layer0_outputs[4972]) & ~(layer0_outputs[3517]);
    assign layer1_outputs[2252] = layer0_outputs[8030];
    assign layer1_outputs[2253] = (layer0_outputs[8784]) & (layer0_outputs[315]);
    assign layer1_outputs[2254] = layer0_outputs[8295];
    assign layer1_outputs[2255] = layer0_outputs[2589];
    assign layer1_outputs[2256] = ~(layer0_outputs[1203]);
    assign layer1_outputs[2257] = layer0_outputs[12767];
    assign layer1_outputs[2258] = ~(layer0_outputs[3434]);
    assign layer1_outputs[2259] = 1'b1;
    assign layer1_outputs[2260] = (layer0_outputs[10240]) & ~(layer0_outputs[164]);
    assign layer1_outputs[2261] = ~((layer0_outputs[4646]) & (layer0_outputs[11024]));
    assign layer1_outputs[2262] = ~(layer0_outputs[5469]);
    assign layer1_outputs[2263] = layer0_outputs[9846];
    assign layer1_outputs[2264] = ~(layer0_outputs[3151]) | (layer0_outputs[12402]);
    assign layer1_outputs[2265] = layer0_outputs[1867];
    assign layer1_outputs[2266] = layer0_outputs[12208];
    assign layer1_outputs[2267] = (layer0_outputs[854]) | (layer0_outputs[6190]);
    assign layer1_outputs[2268] = layer0_outputs[2950];
    assign layer1_outputs[2269] = (layer0_outputs[10431]) & ~(layer0_outputs[2724]);
    assign layer1_outputs[2270] = (layer0_outputs[8662]) & ~(layer0_outputs[1676]);
    assign layer1_outputs[2271] = (layer0_outputs[9659]) | (layer0_outputs[6575]);
    assign layer1_outputs[2272] = (layer0_outputs[1864]) & ~(layer0_outputs[12391]);
    assign layer1_outputs[2273] = (layer0_outputs[8981]) ^ (layer0_outputs[3972]);
    assign layer1_outputs[2274] = ~(layer0_outputs[5493]);
    assign layer1_outputs[2275] = (layer0_outputs[10755]) | (layer0_outputs[11537]);
    assign layer1_outputs[2276] = layer0_outputs[4482];
    assign layer1_outputs[2277] = layer0_outputs[815];
    assign layer1_outputs[2278] = ~(layer0_outputs[11197]);
    assign layer1_outputs[2279] = (layer0_outputs[10562]) & ~(layer0_outputs[5208]);
    assign layer1_outputs[2280] = (layer0_outputs[5705]) & ~(layer0_outputs[1833]);
    assign layer1_outputs[2281] = ~((layer0_outputs[12757]) & (layer0_outputs[9343]));
    assign layer1_outputs[2282] = layer0_outputs[9183];
    assign layer1_outputs[2283] = (layer0_outputs[2602]) & (layer0_outputs[7896]);
    assign layer1_outputs[2284] = ~(layer0_outputs[10658]) | (layer0_outputs[2265]);
    assign layer1_outputs[2285] = (layer0_outputs[5537]) | (layer0_outputs[10509]);
    assign layer1_outputs[2286] = (layer0_outputs[65]) & ~(layer0_outputs[9294]);
    assign layer1_outputs[2287] = (layer0_outputs[1730]) & ~(layer0_outputs[11934]);
    assign layer1_outputs[2288] = ~((layer0_outputs[11088]) | (layer0_outputs[7338]));
    assign layer1_outputs[2289] = layer0_outputs[6830];
    assign layer1_outputs[2290] = ~((layer0_outputs[12015]) ^ (layer0_outputs[5847]));
    assign layer1_outputs[2291] = ~((layer0_outputs[2607]) ^ (layer0_outputs[11792]));
    assign layer1_outputs[2292] = (layer0_outputs[4146]) ^ (layer0_outputs[9125]);
    assign layer1_outputs[2293] = ~(layer0_outputs[942]);
    assign layer1_outputs[2294] = ~(layer0_outputs[12251]);
    assign layer1_outputs[2295] = (layer0_outputs[354]) & (layer0_outputs[8089]);
    assign layer1_outputs[2296] = ~(layer0_outputs[11998]);
    assign layer1_outputs[2297] = (layer0_outputs[2756]) & ~(layer0_outputs[3611]);
    assign layer1_outputs[2298] = ~((layer0_outputs[11151]) ^ (layer0_outputs[9768]));
    assign layer1_outputs[2299] = (layer0_outputs[6558]) ^ (layer0_outputs[4274]);
    assign layer1_outputs[2300] = (layer0_outputs[10864]) | (layer0_outputs[8473]);
    assign layer1_outputs[2301] = (layer0_outputs[5809]) | (layer0_outputs[8736]);
    assign layer1_outputs[2302] = ~((layer0_outputs[3866]) & (layer0_outputs[3253]));
    assign layer1_outputs[2303] = ~(layer0_outputs[8294]) | (layer0_outputs[11890]);
    assign layer1_outputs[2304] = layer0_outputs[7631];
    assign layer1_outputs[2305] = (layer0_outputs[2562]) ^ (layer0_outputs[10029]);
    assign layer1_outputs[2306] = ~(layer0_outputs[12775]);
    assign layer1_outputs[2307] = (layer0_outputs[7176]) & (layer0_outputs[12371]);
    assign layer1_outputs[2308] = ~(layer0_outputs[5253]) | (layer0_outputs[7077]);
    assign layer1_outputs[2309] = ~(layer0_outputs[7844]);
    assign layer1_outputs[2310] = ~(layer0_outputs[11840]) | (layer0_outputs[695]);
    assign layer1_outputs[2311] = ~(layer0_outputs[6050]);
    assign layer1_outputs[2312] = ~((layer0_outputs[8921]) ^ (layer0_outputs[8361]));
    assign layer1_outputs[2313] = (layer0_outputs[9119]) & ~(layer0_outputs[1989]);
    assign layer1_outputs[2314] = layer0_outputs[713];
    assign layer1_outputs[2315] = layer0_outputs[2049];
    assign layer1_outputs[2316] = ~(layer0_outputs[5694]);
    assign layer1_outputs[2317] = (layer0_outputs[11581]) & ~(layer0_outputs[4205]);
    assign layer1_outputs[2318] = layer0_outputs[6075];
    assign layer1_outputs[2319] = (layer0_outputs[12396]) & ~(layer0_outputs[3196]);
    assign layer1_outputs[2320] = ~(layer0_outputs[8431]) | (layer0_outputs[9402]);
    assign layer1_outputs[2321] = ~(layer0_outputs[8162]);
    assign layer1_outputs[2322] = ~(layer0_outputs[6563]) | (layer0_outputs[1812]);
    assign layer1_outputs[2323] = (layer0_outputs[1064]) & ~(layer0_outputs[7467]);
    assign layer1_outputs[2324] = (layer0_outputs[11411]) | (layer0_outputs[8878]);
    assign layer1_outputs[2325] = (layer0_outputs[6269]) | (layer0_outputs[4850]);
    assign layer1_outputs[2326] = layer0_outputs[7746];
    assign layer1_outputs[2327] = ~((layer0_outputs[1652]) & (layer0_outputs[4746]));
    assign layer1_outputs[2328] = ~(layer0_outputs[12611]) | (layer0_outputs[10605]);
    assign layer1_outputs[2329] = ~((layer0_outputs[4829]) & (layer0_outputs[5417]));
    assign layer1_outputs[2330] = ~(layer0_outputs[1928]);
    assign layer1_outputs[2331] = layer0_outputs[3519];
    assign layer1_outputs[2332] = ~(layer0_outputs[9647]);
    assign layer1_outputs[2333] = ~(layer0_outputs[12753]) | (layer0_outputs[12040]);
    assign layer1_outputs[2334] = ~(layer0_outputs[11700]);
    assign layer1_outputs[2335] = layer0_outputs[11295];
    assign layer1_outputs[2336] = (layer0_outputs[6248]) ^ (layer0_outputs[3007]);
    assign layer1_outputs[2337] = (layer0_outputs[573]) | (layer0_outputs[5562]);
    assign layer1_outputs[2338] = ~(layer0_outputs[2766]);
    assign layer1_outputs[2339] = ~(layer0_outputs[10385]);
    assign layer1_outputs[2340] = ~((layer0_outputs[7142]) ^ (layer0_outputs[3079]));
    assign layer1_outputs[2341] = ~(layer0_outputs[7088]);
    assign layer1_outputs[2342] = ~(layer0_outputs[1226]);
    assign layer1_outputs[2343] = (layer0_outputs[5916]) & ~(layer0_outputs[1378]);
    assign layer1_outputs[2344] = ~((layer0_outputs[6855]) | (layer0_outputs[1647]));
    assign layer1_outputs[2345] = (layer0_outputs[6429]) & ~(layer0_outputs[2357]);
    assign layer1_outputs[2346] = (layer0_outputs[8081]) & ~(layer0_outputs[12409]);
    assign layer1_outputs[2347] = ~(layer0_outputs[2634]) | (layer0_outputs[8334]);
    assign layer1_outputs[2348] = ~((layer0_outputs[5184]) | (layer0_outputs[2394]));
    assign layer1_outputs[2349] = ~((layer0_outputs[4248]) | (layer0_outputs[11360]));
    assign layer1_outputs[2350] = ~(layer0_outputs[10662]);
    assign layer1_outputs[2351] = (layer0_outputs[550]) & ~(layer0_outputs[12346]);
    assign layer1_outputs[2352] = layer0_outputs[223];
    assign layer1_outputs[2353] = layer0_outputs[1599];
    assign layer1_outputs[2354] = ~(layer0_outputs[2110]);
    assign layer1_outputs[2355] = ~(layer0_outputs[6009]);
    assign layer1_outputs[2356] = ~(layer0_outputs[2405]);
    assign layer1_outputs[2357] = (layer0_outputs[7685]) ^ (layer0_outputs[11522]);
    assign layer1_outputs[2358] = ~((layer0_outputs[2460]) ^ (layer0_outputs[7542]));
    assign layer1_outputs[2359] = ~(layer0_outputs[9385]);
    assign layer1_outputs[2360] = (layer0_outputs[4668]) ^ (layer0_outputs[289]);
    assign layer1_outputs[2361] = ~(layer0_outputs[6699]);
    assign layer1_outputs[2362] = ~((layer0_outputs[8142]) ^ (layer0_outputs[4273]));
    assign layer1_outputs[2363] = ~((layer0_outputs[10079]) & (layer0_outputs[6757]));
    assign layer1_outputs[2364] = ~(layer0_outputs[4117]);
    assign layer1_outputs[2365] = (layer0_outputs[5952]) | (layer0_outputs[10622]);
    assign layer1_outputs[2366] = 1'b1;
    assign layer1_outputs[2367] = ~(layer0_outputs[5566]) | (layer0_outputs[678]);
    assign layer1_outputs[2368] = (layer0_outputs[3279]) | (layer0_outputs[12247]);
    assign layer1_outputs[2369] = layer0_outputs[9178];
    assign layer1_outputs[2370] = layer0_outputs[2675];
    assign layer1_outputs[2371] = ~(layer0_outputs[4044]);
    assign layer1_outputs[2372] = ~(layer0_outputs[1432]) | (layer0_outputs[1699]);
    assign layer1_outputs[2373] = ~(layer0_outputs[7600]);
    assign layer1_outputs[2374] = layer0_outputs[1404];
    assign layer1_outputs[2375] = ~((layer0_outputs[8420]) | (layer0_outputs[10366]));
    assign layer1_outputs[2376] = ~(layer0_outputs[7326]);
    assign layer1_outputs[2377] = (layer0_outputs[5119]) | (layer0_outputs[11236]);
    assign layer1_outputs[2378] = ~(layer0_outputs[3051]);
    assign layer1_outputs[2379] = (layer0_outputs[10825]) & (layer0_outputs[562]);
    assign layer1_outputs[2380] = ~(layer0_outputs[2336]);
    assign layer1_outputs[2381] = ~(layer0_outputs[7772]) | (layer0_outputs[9807]);
    assign layer1_outputs[2382] = 1'b0;
    assign layer1_outputs[2383] = layer0_outputs[4146];
    assign layer1_outputs[2384] = (layer0_outputs[7314]) ^ (layer0_outputs[10435]);
    assign layer1_outputs[2385] = (layer0_outputs[6912]) & ~(layer0_outputs[3229]);
    assign layer1_outputs[2386] = layer0_outputs[12018];
    assign layer1_outputs[2387] = (layer0_outputs[5717]) | (layer0_outputs[11064]);
    assign layer1_outputs[2388] = layer0_outputs[5605];
    assign layer1_outputs[2389] = layer0_outputs[11143];
    assign layer1_outputs[2390] = ~(layer0_outputs[8682]);
    assign layer1_outputs[2391] = layer0_outputs[5669];
    assign layer1_outputs[2392] = (layer0_outputs[9194]) | (layer0_outputs[4189]);
    assign layer1_outputs[2393] = layer0_outputs[5642];
    assign layer1_outputs[2394] = (layer0_outputs[7627]) & (layer0_outputs[3664]);
    assign layer1_outputs[2395] = ~(layer0_outputs[174]);
    assign layer1_outputs[2396] = (layer0_outputs[3226]) ^ (layer0_outputs[12755]);
    assign layer1_outputs[2397] = layer0_outputs[11069];
    assign layer1_outputs[2398] = (layer0_outputs[11826]) ^ (layer0_outputs[9112]);
    assign layer1_outputs[2399] = (layer0_outputs[12636]) & ~(layer0_outputs[8999]);
    assign layer1_outputs[2400] = (layer0_outputs[191]) & (layer0_outputs[9753]);
    assign layer1_outputs[2401] = ~(layer0_outputs[12488]) | (layer0_outputs[5484]);
    assign layer1_outputs[2402] = (layer0_outputs[8144]) & ~(layer0_outputs[280]);
    assign layer1_outputs[2403] = layer0_outputs[9390];
    assign layer1_outputs[2404] = (layer0_outputs[10156]) & (layer0_outputs[858]);
    assign layer1_outputs[2405] = ~((layer0_outputs[2380]) ^ (layer0_outputs[926]));
    assign layer1_outputs[2406] = ~(layer0_outputs[7061]);
    assign layer1_outputs[2407] = ~(layer0_outputs[3068]);
    assign layer1_outputs[2408] = (layer0_outputs[12474]) & ~(layer0_outputs[9082]);
    assign layer1_outputs[2409] = (layer0_outputs[4975]) & (layer0_outputs[10087]);
    assign layer1_outputs[2410] = (layer0_outputs[6932]) & (layer0_outputs[6838]);
    assign layer1_outputs[2411] = (layer0_outputs[10775]) & ~(layer0_outputs[352]);
    assign layer1_outputs[2412] = layer0_outputs[8773];
    assign layer1_outputs[2413] = ~(layer0_outputs[4119]);
    assign layer1_outputs[2414] = layer0_outputs[10696];
    assign layer1_outputs[2415] = layer0_outputs[12630];
    assign layer1_outputs[2416] = (layer0_outputs[12030]) & ~(layer0_outputs[8344]);
    assign layer1_outputs[2417] = ~(layer0_outputs[6172]);
    assign layer1_outputs[2418] = ~((layer0_outputs[3423]) & (layer0_outputs[9798]));
    assign layer1_outputs[2419] = 1'b0;
    assign layer1_outputs[2420] = ~(layer0_outputs[1754]) | (layer0_outputs[10666]);
    assign layer1_outputs[2421] = layer0_outputs[6448];
    assign layer1_outputs[2422] = ~(layer0_outputs[11330]) | (layer0_outputs[2866]);
    assign layer1_outputs[2423] = (layer0_outputs[10209]) ^ (layer0_outputs[6320]);
    assign layer1_outputs[2424] = ~(layer0_outputs[964]);
    assign layer1_outputs[2425] = ~(layer0_outputs[8332]);
    assign layer1_outputs[2426] = ~((layer0_outputs[10731]) | (layer0_outputs[9359]));
    assign layer1_outputs[2427] = layer0_outputs[431];
    assign layer1_outputs[2428] = ~(layer0_outputs[4420]);
    assign layer1_outputs[2429] = (layer0_outputs[8052]) & (layer0_outputs[6311]);
    assign layer1_outputs[2430] = layer0_outputs[6994];
    assign layer1_outputs[2431] = 1'b1;
    assign layer1_outputs[2432] = (layer0_outputs[7888]) & ~(layer0_outputs[5149]);
    assign layer1_outputs[2433] = ~(layer0_outputs[7416]);
    assign layer1_outputs[2434] = ~(layer0_outputs[4949]);
    assign layer1_outputs[2435] = ~((layer0_outputs[11301]) & (layer0_outputs[42]));
    assign layer1_outputs[2436] = layer0_outputs[8389];
    assign layer1_outputs[2437] = ~((layer0_outputs[1812]) ^ (layer0_outputs[6716]));
    assign layer1_outputs[2438] = ~((layer0_outputs[4586]) & (layer0_outputs[10213]));
    assign layer1_outputs[2439] = (layer0_outputs[12271]) ^ (layer0_outputs[4845]);
    assign layer1_outputs[2440] = layer0_outputs[288];
    assign layer1_outputs[2441] = layer0_outputs[4229];
    assign layer1_outputs[2442] = (layer0_outputs[7831]) | (layer0_outputs[328]);
    assign layer1_outputs[2443] = ~(layer0_outputs[3468]);
    assign layer1_outputs[2444] = (layer0_outputs[4667]) & ~(layer0_outputs[10140]);
    assign layer1_outputs[2445] = (layer0_outputs[7138]) & ~(layer0_outputs[8436]);
    assign layer1_outputs[2446] = ~((layer0_outputs[10980]) & (layer0_outputs[2810]));
    assign layer1_outputs[2447] = ~((layer0_outputs[12417]) ^ (layer0_outputs[6083]));
    assign layer1_outputs[2448] = layer0_outputs[6093];
    assign layer1_outputs[2449] = (layer0_outputs[701]) | (layer0_outputs[9277]);
    assign layer1_outputs[2450] = layer0_outputs[6533];
    assign layer1_outputs[2451] = ~(layer0_outputs[3052]) | (layer0_outputs[10448]);
    assign layer1_outputs[2452] = ~(layer0_outputs[11184]);
    assign layer1_outputs[2453] = (layer0_outputs[2692]) & ~(layer0_outputs[8697]);
    assign layer1_outputs[2454] = ~(layer0_outputs[4816]);
    assign layer1_outputs[2455] = (layer0_outputs[12156]) & (layer0_outputs[9564]);
    assign layer1_outputs[2456] = ~((layer0_outputs[12633]) ^ (layer0_outputs[11323]));
    assign layer1_outputs[2457] = ~(layer0_outputs[4831]) | (layer0_outputs[10314]);
    assign layer1_outputs[2458] = layer0_outputs[1920];
    assign layer1_outputs[2459] = layer0_outputs[3782];
    assign layer1_outputs[2460] = (layer0_outputs[9707]) ^ (layer0_outputs[6228]);
    assign layer1_outputs[2461] = layer0_outputs[10179];
    assign layer1_outputs[2462] = layer0_outputs[6126];
    assign layer1_outputs[2463] = ~(layer0_outputs[10137]);
    assign layer1_outputs[2464] = ~((layer0_outputs[4012]) ^ (layer0_outputs[1614]));
    assign layer1_outputs[2465] = ~(layer0_outputs[8758]);
    assign layer1_outputs[2466] = (layer0_outputs[12068]) ^ (layer0_outputs[3345]);
    assign layer1_outputs[2467] = 1'b1;
    assign layer1_outputs[2468] = (layer0_outputs[3432]) & (layer0_outputs[983]);
    assign layer1_outputs[2469] = (layer0_outputs[5797]) & ~(layer0_outputs[6330]);
    assign layer1_outputs[2470] = (layer0_outputs[5007]) | (layer0_outputs[8321]);
    assign layer1_outputs[2471] = ~(layer0_outputs[8154]) | (layer0_outputs[10887]);
    assign layer1_outputs[2472] = (layer0_outputs[988]) & ~(layer0_outputs[10421]);
    assign layer1_outputs[2473] = layer0_outputs[5050];
    assign layer1_outputs[2474] = (layer0_outputs[6554]) & (layer0_outputs[6210]);
    assign layer1_outputs[2475] = ~(layer0_outputs[4949]);
    assign layer1_outputs[2476] = ~(layer0_outputs[10900]);
    assign layer1_outputs[2477] = ~(layer0_outputs[9292]);
    assign layer1_outputs[2478] = ~(layer0_outputs[12291]) | (layer0_outputs[8071]);
    assign layer1_outputs[2479] = ~(layer0_outputs[4003]);
    assign layer1_outputs[2480] = layer0_outputs[3641];
    assign layer1_outputs[2481] = ~(layer0_outputs[7588]);
    assign layer1_outputs[2482] = ~(layer0_outputs[3743]);
    assign layer1_outputs[2483] = ~((layer0_outputs[8985]) & (layer0_outputs[9491]));
    assign layer1_outputs[2484] = layer0_outputs[11083];
    assign layer1_outputs[2485] = ~((layer0_outputs[11041]) & (layer0_outputs[2944]));
    assign layer1_outputs[2486] = layer0_outputs[7851];
    assign layer1_outputs[2487] = layer0_outputs[8521];
    assign layer1_outputs[2488] = ~((layer0_outputs[11843]) & (layer0_outputs[3887]));
    assign layer1_outputs[2489] = layer0_outputs[10153];
    assign layer1_outputs[2490] = layer0_outputs[11110];
    assign layer1_outputs[2491] = 1'b0;
    assign layer1_outputs[2492] = (layer0_outputs[10776]) & ~(layer0_outputs[888]);
    assign layer1_outputs[2493] = layer0_outputs[2375];
    assign layer1_outputs[2494] = ~((layer0_outputs[7724]) | (layer0_outputs[846]));
    assign layer1_outputs[2495] = ~(layer0_outputs[6172]) | (layer0_outputs[6933]);
    assign layer1_outputs[2496] = (layer0_outputs[379]) | (layer0_outputs[9540]);
    assign layer1_outputs[2497] = (layer0_outputs[1818]) & (layer0_outputs[6871]);
    assign layer1_outputs[2498] = (layer0_outputs[8349]) & ~(layer0_outputs[1831]);
    assign layer1_outputs[2499] = layer0_outputs[12638];
    assign layer1_outputs[2500] = ~((layer0_outputs[4529]) | (layer0_outputs[7113]));
    assign layer1_outputs[2501] = layer0_outputs[3525];
    assign layer1_outputs[2502] = ~((layer0_outputs[2373]) ^ (layer0_outputs[5449]));
    assign layer1_outputs[2503] = ~(layer0_outputs[9659]) | (layer0_outputs[5354]);
    assign layer1_outputs[2504] = ~(layer0_outputs[2505]) | (layer0_outputs[561]);
    assign layer1_outputs[2505] = ~(layer0_outputs[4409]) | (layer0_outputs[8470]);
    assign layer1_outputs[2506] = (layer0_outputs[6588]) & ~(layer0_outputs[9401]);
    assign layer1_outputs[2507] = (layer0_outputs[399]) & (layer0_outputs[4059]);
    assign layer1_outputs[2508] = (layer0_outputs[3358]) | (layer0_outputs[9086]);
    assign layer1_outputs[2509] = ~(layer0_outputs[3115]) | (layer0_outputs[7162]);
    assign layer1_outputs[2510] = ~(layer0_outputs[7088]);
    assign layer1_outputs[2511] = ~(layer0_outputs[9642]);
    assign layer1_outputs[2512] = ~((layer0_outputs[9092]) ^ (layer0_outputs[6577]));
    assign layer1_outputs[2513] = ~((layer0_outputs[11745]) | (layer0_outputs[4290]));
    assign layer1_outputs[2514] = ~(layer0_outputs[6688]);
    assign layer1_outputs[2515] = layer0_outputs[6911];
    assign layer1_outputs[2516] = layer0_outputs[6483];
    assign layer1_outputs[2517] = ~(layer0_outputs[1883]);
    assign layer1_outputs[2518] = layer0_outputs[11514];
    assign layer1_outputs[2519] = ~(layer0_outputs[1968]);
    assign layer1_outputs[2520] = 1'b0;
    assign layer1_outputs[2521] = ~(layer0_outputs[8178]);
    assign layer1_outputs[2522] = (layer0_outputs[5684]) & (layer0_outputs[10635]);
    assign layer1_outputs[2523] = ~((layer0_outputs[6196]) & (layer0_outputs[5307]));
    assign layer1_outputs[2524] = layer0_outputs[9991];
    assign layer1_outputs[2525] = ~(layer0_outputs[4135]);
    assign layer1_outputs[2526] = ~(layer0_outputs[4957]);
    assign layer1_outputs[2527] = (layer0_outputs[5892]) & ~(layer0_outputs[4844]);
    assign layer1_outputs[2528] = layer0_outputs[6961];
    assign layer1_outputs[2529] = (layer0_outputs[8184]) ^ (layer0_outputs[11043]);
    assign layer1_outputs[2530] = (layer0_outputs[8378]) | (layer0_outputs[5970]);
    assign layer1_outputs[2531] = layer0_outputs[7809];
    assign layer1_outputs[2532] = ~(layer0_outputs[12627]);
    assign layer1_outputs[2533] = ~(layer0_outputs[12435]);
    assign layer1_outputs[2534] = ~((layer0_outputs[1809]) ^ (layer0_outputs[6368]));
    assign layer1_outputs[2535] = ~(layer0_outputs[2284]);
    assign layer1_outputs[2536] = ~(layer0_outputs[6589]);
    assign layer1_outputs[2537] = ~(layer0_outputs[3720]);
    assign layer1_outputs[2538] = layer0_outputs[10010];
    assign layer1_outputs[2539] = (layer0_outputs[10346]) & ~(layer0_outputs[3745]);
    assign layer1_outputs[2540] = layer0_outputs[1753];
    assign layer1_outputs[2541] = ~((layer0_outputs[249]) & (layer0_outputs[3368]));
    assign layer1_outputs[2542] = ~((layer0_outputs[9823]) ^ (layer0_outputs[5328]));
    assign layer1_outputs[2543] = ~(layer0_outputs[8692]);
    assign layer1_outputs[2544] = ~((layer0_outputs[10145]) | (layer0_outputs[10825]));
    assign layer1_outputs[2545] = ~((layer0_outputs[2499]) & (layer0_outputs[11000]));
    assign layer1_outputs[2546] = (layer0_outputs[11262]) & (layer0_outputs[288]);
    assign layer1_outputs[2547] = ~((layer0_outputs[10115]) ^ (layer0_outputs[12111]));
    assign layer1_outputs[2548] = (layer0_outputs[11467]) & ~(layer0_outputs[3799]);
    assign layer1_outputs[2549] = layer0_outputs[11039];
    assign layer1_outputs[2550] = ~(layer0_outputs[7632]);
    assign layer1_outputs[2551] = ~(layer0_outputs[11290]) | (layer0_outputs[12306]);
    assign layer1_outputs[2552] = (layer0_outputs[278]) ^ (layer0_outputs[3055]);
    assign layer1_outputs[2553] = layer0_outputs[11335];
    assign layer1_outputs[2554] = ~(layer0_outputs[11388]) | (layer0_outputs[8439]);
    assign layer1_outputs[2555] = ~((layer0_outputs[11030]) | (layer0_outputs[1826]));
    assign layer1_outputs[2556] = (layer0_outputs[1311]) & ~(layer0_outputs[7095]);
    assign layer1_outputs[2557] = (layer0_outputs[842]) & ~(layer0_outputs[11548]);
    assign layer1_outputs[2558] = ~(layer0_outputs[11051]) | (layer0_outputs[11558]);
    assign layer1_outputs[2559] = (layer0_outputs[2913]) ^ (layer0_outputs[6332]);
    assign layer1_outputs[2560] = layer0_outputs[4906];
    assign layer1_outputs[2561] = layer0_outputs[10736];
    assign layer1_outputs[2562] = ~(layer0_outputs[12452]) | (layer0_outputs[5478]);
    assign layer1_outputs[2563] = ~(layer0_outputs[1496]) | (layer0_outputs[2702]);
    assign layer1_outputs[2564] = layer0_outputs[4181];
    assign layer1_outputs[2565] = ~(layer0_outputs[11840]);
    assign layer1_outputs[2566] = ~(layer0_outputs[11663]) | (layer0_outputs[12581]);
    assign layer1_outputs[2567] = ~(layer0_outputs[3281]);
    assign layer1_outputs[2568] = layer0_outputs[10102];
    assign layer1_outputs[2569] = ~((layer0_outputs[6774]) ^ (layer0_outputs[6393]));
    assign layer1_outputs[2570] = (layer0_outputs[2402]) & ~(layer0_outputs[1010]);
    assign layer1_outputs[2571] = ~((layer0_outputs[4929]) ^ (layer0_outputs[11042]));
    assign layer1_outputs[2572] = layer0_outputs[3307];
    assign layer1_outputs[2573] = layer0_outputs[5198];
    assign layer1_outputs[2574] = ~(layer0_outputs[10764]);
    assign layer1_outputs[2575] = ~(layer0_outputs[5305]) | (layer0_outputs[11889]);
    assign layer1_outputs[2576] = ~(layer0_outputs[8894]) | (layer0_outputs[620]);
    assign layer1_outputs[2577] = (layer0_outputs[9088]) | (layer0_outputs[6741]);
    assign layer1_outputs[2578] = ~((layer0_outputs[10934]) ^ (layer0_outputs[1534]));
    assign layer1_outputs[2579] = ~(layer0_outputs[198]) | (layer0_outputs[4636]);
    assign layer1_outputs[2580] = ~(layer0_outputs[5946]) | (layer0_outputs[12182]);
    assign layer1_outputs[2581] = ~(layer0_outputs[6060]);
    assign layer1_outputs[2582] = ~(layer0_outputs[3630]);
    assign layer1_outputs[2583] = ~((layer0_outputs[8962]) | (layer0_outputs[382]));
    assign layer1_outputs[2584] = layer0_outputs[11595];
    assign layer1_outputs[2585] = ~((layer0_outputs[6343]) & (layer0_outputs[7171]));
    assign layer1_outputs[2586] = (layer0_outputs[1580]) & (layer0_outputs[6230]);
    assign layer1_outputs[2587] = ~(layer0_outputs[11999]);
    assign layer1_outputs[2588] = ~(layer0_outputs[9509]) | (layer0_outputs[239]);
    assign layer1_outputs[2589] = layer0_outputs[434];
    assign layer1_outputs[2590] = ~(layer0_outputs[4266]);
    assign layer1_outputs[2591] = (layer0_outputs[7141]) & ~(layer0_outputs[4150]);
    assign layer1_outputs[2592] = 1'b0;
    assign layer1_outputs[2593] = ~(layer0_outputs[12702]);
    assign layer1_outputs[2594] = layer0_outputs[12556];
    assign layer1_outputs[2595] = (layer0_outputs[5259]) | (layer0_outputs[5061]);
    assign layer1_outputs[2596] = (layer0_outputs[12260]) ^ (layer0_outputs[9204]);
    assign layer1_outputs[2597] = ~((layer0_outputs[1276]) & (layer0_outputs[3543]));
    assign layer1_outputs[2598] = ~(layer0_outputs[9104]);
    assign layer1_outputs[2599] = (layer0_outputs[7818]) & (layer0_outputs[12137]);
    assign layer1_outputs[2600] = ~(layer0_outputs[200]) | (layer0_outputs[11560]);
    assign layer1_outputs[2601] = layer0_outputs[3758];
    assign layer1_outputs[2602] = ~(layer0_outputs[11347]);
    assign layer1_outputs[2603] = ~(layer0_outputs[1417]);
    assign layer1_outputs[2604] = ~(layer0_outputs[12544]);
    assign layer1_outputs[2605] = (layer0_outputs[4982]) & ~(layer0_outputs[1650]);
    assign layer1_outputs[2606] = (layer0_outputs[9694]) & ~(layer0_outputs[1798]);
    assign layer1_outputs[2607] = ~((layer0_outputs[6985]) ^ (layer0_outputs[7139]));
    assign layer1_outputs[2608] = (layer0_outputs[11097]) & (layer0_outputs[5461]);
    assign layer1_outputs[2609] = layer0_outputs[1831];
    assign layer1_outputs[2610] = (layer0_outputs[9681]) | (layer0_outputs[9982]);
    assign layer1_outputs[2611] = 1'b0;
    assign layer1_outputs[2612] = 1'b0;
    assign layer1_outputs[2613] = layer0_outputs[5131];
    assign layer1_outputs[2614] = ~(layer0_outputs[6347]);
    assign layer1_outputs[2615] = (layer0_outputs[12617]) ^ (layer0_outputs[2126]);
    assign layer1_outputs[2616] = 1'b0;
    assign layer1_outputs[2617] = ~((layer0_outputs[10951]) & (layer0_outputs[4339]));
    assign layer1_outputs[2618] = 1'b1;
    assign layer1_outputs[2619] = (layer0_outputs[11816]) & (layer0_outputs[8266]);
    assign layer1_outputs[2620] = ~(layer0_outputs[2267]);
    assign layer1_outputs[2621] = ~(layer0_outputs[9475]);
    assign layer1_outputs[2622] = ~((layer0_outputs[11911]) & (layer0_outputs[196]));
    assign layer1_outputs[2623] = (layer0_outputs[9948]) ^ (layer0_outputs[10621]);
    assign layer1_outputs[2624] = layer0_outputs[6355];
    assign layer1_outputs[2625] = (layer0_outputs[3995]) & ~(layer0_outputs[7643]);
    assign layer1_outputs[2626] = ~(layer0_outputs[3351]) | (layer0_outputs[2496]);
    assign layer1_outputs[2627] = ~((layer0_outputs[8632]) | (layer0_outputs[5850]));
    assign layer1_outputs[2628] = ~(layer0_outputs[5552]);
    assign layer1_outputs[2629] = (layer0_outputs[12267]) & (layer0_outputs[472]);
    assign layer1_outputs[2630] = ~(layer0_outputs[3330]) | (layer0_outputs[5115]);
    assign layer1_outputs[2631] = layer0_outputs[5656];
    assign layer1_outputs[2632] = 1'b1;
    assign layer1_outputs[2633] = layer0_outputs[12766];
    assign layer1_outputs[2634] = ~(layer0_outputs[2789]) | (layer0_outputs[9006]);
    assign layer1_outputs[2635] = ~((layer0_outputs[52]) & (layer0_outputs[5854]));
    assign layer1_outputs[2636] = (layer0_outputs[5817]) ^ (layer0_outputs[10601]);
    assign layer1_outputs[2637] = ~((layer0_outputs[6369]) & (layer0_outputs[907]));
    assign layer1_outputs[2638] = ~(layer0_outputs[4912]);
    assign layer1_outputs[2639] = layer0_outputs[6134];
    assign layer1_outputs[2640] = ~((layer0_outputs[1579]) & (layer0_outputs[7678]));
    assign layer1_outputs[2641] = (layer0_outputs[9933]) & ~(layer0_outputs[1840]);
    assign layer1_outputs[2642] = (layer0_outputs[821]) & ~(layer0_outputs[3302]);
    assign layer1_outputs[2643] = ~(layer0_outputs[7091]) | (layer0_outputs[9824]);
    assign layer1_outputs[2644] = layer0_outputs[6016];
    assign layer1_outputs[2645] = ~(layer0_outputs[2998]);
    assign layer1_outputs[2646] = ~(layer0_outputs[5001]);
    assign layer1_outputs[2647] = layer0_outputs[12210];
    assign layer1_outputs[2648] = layer0_outputs[4265];
    assign layer1_outputs[2649] = ~(layer0_outputs[1341]) | (layer0_outputs[9045]);
    assign layer1_outputs[2650] = ~((layer0_outputs[7082]) & (layer0_outputs[657]));
    assign layer1_outputs[2651] = ~(layer0_outputs[11429]);
    assign layer1_outputs[2652] = layer0_outputs[2516];
    assign layer1_outputs[2653] = layer0_outputs[6849];
    assign layer1_outputs[2654] = layer0_outputs[593];
    assign layer1_outputs[2655] = ~(layer0_outputs[1037]);
    assign layer1_outputs[2656] = ~(layer0_outputs[12196]);
    assign layer1_outputs[2657] = (layer0_outputs[10417]) ^ (layer0_outputs[3159]);
    assign layer1_outputs[2658] = (layer0_outputs[8380]) & ~(layer0_outputs[1937]);
    assign layer1_outputs[2659] = 1'b1;
    assign layer1_outputs[2660] = ~(layer0_outputs[12256]);
    assign layer1_outputs[2661] = ~(layer0_outputs[9798]) | (layer0_outputs[10569]);
    assign layer1_outputs[2662] = ~(layer0_outputs[504]);
    assign layer1_outputs[2663] = (layer0_outputs[4967]) & ~(layer0_outputs[5025]);
    assign layer1_outputs[2664] = layer0_outputs[3613];
    assign layer1_outputs[2665] = ~((layer0_outputs[6045]) ^ (layer0_outputs[7263]));
    assign layer1_outputs[2666] = ~(layer0_outputs[8383]) | (layer0_outputs[12272]);
    assign layer1_outputs[2667] = (layer0_outputs[8729]) & ~(layer0_outputs[11590]);
    assign layer1_outputs[2668] = ~(layer0_outputs[10291]);
    assign layer1_outputs[2669] = (layer0_outputs[9345]) & ~(layer0_outputs[2746]);
    assign layer1_outputs[2670] = ~(layer0_outputs[11959]);
    assign layer1_outputs[2671] = ~(layer0_outputs[7006]);
    assign layer1_outputs[2672] = ~(layer0_outputs[7283]);
    assign layer1_outputs[2673] = ~((layer0_outputs[7605]) | (layer0_outputs[8213]));
    assign layer1_outputs[2674] = ~(layer0_outputs[742]);
    assign layer1_outputs[2675] = (layer0_outputs[2318]) | (layer0_outputs[2793]);
    assign layer1_outputs[2676] = (layer0_outputs[10030]) | (layer0_outputs[5613]);
    assign layer1_outputs[2677] = ~(layer0_outputs[1457]) | (layer0_outputs[10207]);
    assign layer1_outputs[2678] = ~(layer0_outputs[471]);
    assign layer1_outputs[2679] = (layer0_outputs[10519]) | (layer0_outputs[1948]);
    assign layer1_outputs[2680] = ~((layer0_outputs[7702]) & (layer0_outputs[7177]));
    assign layer1_outputs[2681] = ~(layer0_outputs[3297]);
    assign layer1_outputs[2682] = (layer0_outputs[8250]) & ~(layer0_outputs[11218]);
    assign layer1_outputs[2683] = ~(layer0_outputs[9841]);
    assign layer1_outputs[2684] = layer0_outputs[9864];
    assign layer1_outputs[2685] = layer0_outputs[6440];
    assign layer1_outputs[2686] = ~(layer0_outputs[2069]) | (layer0_outputs[4336]);
    assign layer1_outputs[2687] = ~((layer0_outputs[22]) ^ (layer0_outputs[1970]));
    assign layer1_outputs[2688] = (layer0_outputs[3289]) ^ (layer0_outputs[36]);
    assign layer1_outputs[2689] = ~((layer0_outputs[12259]) ^ (layer0_outputs[6133]));
    assign layer1_outputs[2690] = ~(layer0_outputs[9608]);
    assign layer1_outputs[2691] = ~((layer0_outputs[511]) ^ (layer0_outputs[11371]));
    assign layer1_outputs[2692] = ~(layer0_outputs[6287]);
    assign layer1_outputs[2693] = ~((layer0_outputs[7301]) & (layer0_outputs[11809]));
    assign layer1_outputs[2694] = (layer0_outputs[10016]) | (layer0_outputs[7433]);
    assign layer1_outputs[2695] = (layer0_outputs[3000]) ^ (layer0_outputs[3979]);
    assign layer1_outputs[2696] = (layer0_outputs[7736]) & ~(layer0_outputs[4699]);
    assign layer1_outputs[2697] = ~(layer0_outputs[6000]);
    assign layer1_outputs[2698] = (layer0_outputs[6767]) & ~(layer0_outputs[6856]);
    assign layer1_outputs[2699] = ~(layer0_outputs[4107]);
    assign layer1_outputs[2700] = layer0_outputs[4182];
    assign layer1_outputs[2701] = (layer0_outputs[11267]) & ~(layer0_outputs[6007]);
    assign layer1_outputs[2702] = ~(layer0_outputs[4104]);
    assign layer1_outputs[2703] = (layer0_outputs[5791]) & (layer0_outputs[98]);
    assign layer1_outputs[2704] = ~(layer0_outputs[11926]);
    assign layer1_outputs[2705] = ~(layer0_outputs[7843]);
    assign layer1_outputs[2706] = ~((layer0_outputs[1382]) ^ (layer0_outputs[9324]));
    assign layer1_outputs[2707] = layer0_outputs[4866];
    assign layer1_outputs[2708] = (layer0_outputs[1933]) & ~(layer0_outputs[12697]);
    assign layer1_outputs[2709] = ~(layer0_outputs[10079]);
    assign layer1_outputs[2710] = (layer0_outputs[8274]) | (layer0_outputs[12214]);
    assign layer1_outputs[2711] = ~(layer0_outputs[9731]);
    assign layer1_outputs[2712] = (layer0_outputs[11999]) & (layer0_outputs[9620]);
    assign layer1_outputs[2713] = ~(layer0_outputs[9700]);
    assign layer1_outputs[2714] = layer0_outputs[6587];
    assign layer1_outputs[2715] = ~(layer0_outputs[6043]);
    assign layer1_outputs[2716] = ~(layer0_outputs[7321]) | (layer0_outputs[8867]);
    assign layer1_outputs[2717] = (layer0_outputs[5660]) | (layer0_outputs[5255]);
    assign layer1_outputs[2718] = layer0_outputs[6519];
    assign layer1_outputs[2719] = 1'b1;
    assign layer1_outputs[2720] = ~(layer0_outputs[9568]) | (layer0_outputs[7716]);
    assign layer1_outputs[2721] = (layer0_outputs[306]) ^ (layer0_outputs[9598]);
    assign layer1_outputs[2722] = ~((layer0_outputs[3238]) ^ (layer0_outputs[9793]));
    assign layer1_outputs[2723] = layer0_outputs[9390];
    assign layer1_outputs[2724] = (layer0_outputs[10739]) ^ (layer0_outputs[1596]);
    assign layer1_outputs[2725] = ~(layer0_outputs[276]);
    assign layer1_outputs[2726] = layer0_outputs[796];
    assign layer1_outputs[2727] = ~(layer0_outputs[8718]);
    assign layer1_outputs[2728] = ~((layer0_outputs[6652]) | (layer0_outputs[4]));
    assign layer1_outputs[2729] = ~(layer0_outputs[12279]);
    assign layer1_outputs[2730] = (layer0_outputs[10852]) ^ (layer0_outputs[7911]);
    assign layer1_outputs[2731] = ~(layer0_outputs[8927]);
    assign layer1_outputs[2732] = ~(layer0_outputs[2873]);
    assign layer1_outputs[2733] = (layer0_outputs[3123]) & ~(layer0_outputs[8587]);
    assign layer1_outputs[2734] = ~((layer0_outputs[12080]) ^ (layer0_outputs[4188]));
    assign layer1_outputs[2735] = ~(layer0_outputs[5633]) | (layer0_outputs[4395]);
    assign layer1_outputs[2736] = (layer0_outputs[10959]) ^ (layer0_outputs[2082]);
    assign layer1_outputs[2737] = ~(layer0_outputs[495]);
    assign layer1_outputs[2738] = ~(layer0_outputs[1871]);
    assign layer1_outputs[2739] = ~(layer0_outputs[10244]) | (layer0_outputs[9159]);
    assign layer1_outputs[2740] = (layer0_outputs[89]) & ~(layer0_outputs[11362]);
    assign layer1_outputs[2741] = (layer0_outputs[1553]) & (layer0_outputs[486]);
    assign layer1_outputs[2742] = layer0_outputs[11583];
    assign layer1_outputs[2743] = 1'b1;
    assign layer1_outputs[2744] = ~((layer0_outputs[6237]) ^ (layer0_outputs[12494]));
    assign layer1_outputs[2745] = ~(layer0_outputs[5161]);
    assign layer1_outputs[2746] = layer0_outputs[2338];
    assign layer1_outputs[2747] = 1'b0;
    assign layer1_outputs[2748] = (layer0_outputs[2287]) & ~(layer0_outputs[2701]);
    assign layer1_outputs[2749] = ~((layer0_outputs[2904]) ^ (layer0_outputs[9251]));
    assign layer1_outputs[2750] = ~(layer0_outputs[5746]);
    assign layer1_outputs[2751] = ~(layer0_outputs[4654]);
    assign layer1_outputs[2752] = ~((layer0_outputs[9914]) | (layer0_outputs[10053]));
    assign layer1_outputs[2753] = layer0_outputs[4096];
    assign layer1_outputs[2754] = layer0_outputs[3053];
    assign layer1_outputs[2755] = 1'b1;
    assign layer1_outputs[2756] = layer0_outputs[3395];
    assign layer1_outputs[2757] = (layer0_outputs[2939]) | (layer0_outputs[12438]);
    assign layer1_outputs[2758] = layer0_outputs[11810];
    assign layer1_outputs[2759] = (layer0_outputs[8247]) & ~(layer0_outputs[4635]);
    assign layer1_outputs[2760] = layer0_outputs[4856];
    assign layer1_outputs[2761] = layer0_outputs[3397];
    assign layer1_outputs[2762] = ~((layer0_outputs[10637]) | (layer0_outputs[9453]));
    assign layer1_outputs[2763] = layer0_outputs[4973];
    assign layer1_outputs[2764] = (layer0_outputs[9662]) ^ (layer0_outputs[11654]);
    assign layer1_outputs[2765] = ~(layer0_outputs[1546]);
    assign layer1_outputs[2766] = layer0_outputs[10634];
    assign layer1_outputs[2767] = ~(layer0_outputs[3554]);
    assign layer1_outputs[2768] = (layer0_outputs[5762]) | (layer0_outputs[10405]);
    assign layer1_outputs[2769] = (layer0_outputs[1921]) ^ (layer0_outputs[3549]);
    assign layer1_outputs[2770] = layer0_outputs[2090];
    assign layer1_outputs[2771] = ~((layer0_outputs[8529]) & (layer0_outputs[11692]));
    assign layer1_outputs[2772] = 1'b1;
    assign layer1_outputs[2773] = ~(layer0_outputs[3789]);
    assign layer1_outputs[2774] = layer0_outputs[11948];
    assign layer1_outputs[2775] = (layer0_outputs[8268]) | (layer0_outputs[5977]);
    assign layer1_outputs[2776] = ~(layer0_outputs[9650]);
    assign layer1_outputs[2777] = ~(layer0_outputs[4591]);
    assign layer1_outputs[2778] = ~(layer0_outputs[9660]);
    assign layer1_outputs[2779] = (layer0_outputs[7118]) ^ (layer0_outputs[3668]);
    assign layer1_outputs[2780] = ~(layer0_outputs[5534]);
    assign layer1_outputs[2781] = (layer0_outputs[4336]) ^ (layer0_outputs[11038]);
    assign layer1_outputs[2782] = ~((layer0_outputs[9620]) | (layer0_outputs[2298]));
    assign layer1_outputs[2783] = (layer0_outputs[10312]) | (layer0_outputs[7920]);
    assign layer1_outputs[2784] = 1'b0;
    assign layer1_outputs[2785] = (layer0_outputs[409]) & ~(layer0_outputs[7610]);
    assign layer1_outputs[2786] = layer0_outputs[5524];
    assign layer1_outputs[2787] = ~(layer0_outputs[11800]);
    assign layer1_outputs[2788] = (layer0_outputs[4034]) | (layer0_outputs[4343]);
    assign layer1_outputs[2789] = ~(layer0_outputs[687]) | (layer0_outputs[757]);
    assign layer1_outputs[2790] = layer0_outputs[4004];
    assign layer1_outputs[2791] = ~((layer0_outputs[5419]) ^ (layer0_outputs[4255]));
    assign layer1_outputs[2792] = layer0_outputs[2363];
    assign layer1_outputs[2793] = ~((layer0_outputs[10849]) & (layer0_outputs[3140]));
    assign layer1_outputs[2794] = layer0_outputs[12207];
    assign layer1_outputs[2795] = layer0_outputs[9679];
    assign layer1_outputs[2796] = ~(layer0_outputs[7001]);
    assign layer1_outputs[2797] = (layer0_outputs[12096]) | (layer0_outputs[9690]);
    assign layer1_outputs[2798] = (layer0_outputs[11592]) & (layer0_outputs[8526]);
    assign layer1_outputs[2799] = ~((layer0_outputs[1063]) | (layer0_outputs[6718]));
    assign layer1_outputs[2800] = ~(layer0_outputs[2234]);
    assign layer1_outputs[2801] = ~(layer0_outputs[9671]);
    assign layer1_outputs[2802] = ~(layer0_outputs[7045]);
    assign layer1_outputs[2803] = (layer0_outputs[1229]) & (layer0_outputs[2647]);
    assign layer1_outputs[2804] = ~((layer0_outputs[6203]) & (layer0_outputs[3139]));
    assign layer1_outputs[2805] = layer0_outputs[12598];
    assign layer1_outputs[2806] = ~(layer0_outputs[1528]) | (layer0_outputs[2817]);
    assign layer1_outputs[2807] = layer0_outputs[4261];
    assign layer1_outputs[2808] = (layer0_outputs[12110]) ^ (layer0_outputs[7606]);
    assign layer1_outputs[2809] = (layer0_outputs[789]) ^ (layer0_outputs[11487]);
    assign layer1_outputs[2810] = layer0_outputs[4737];
    assign layer1_outputs[2811] = (layer0_outputs[253]) ^ (layer0_outputs[6035]);
    assign layer1_outputs[2812] = (layer0_outputs[5818]) & ~(layer0_outputs[10432]);
    assign layer1_outputs[2813] = ~((layer0_outputs[9195]) ^ (layer0_outputs[7447]));
    assign layer1_outputs[2814] = layer0_outputs[10176];
    assign layer1_outputs[2815] = ~(layer0_outputs[2861]);
    assign layer1_outputs[2816] = layer0_outputs[2715];
    assign layer1_outputs[2817] = ~((layer0_outputs[8034]) & (layer0_outputs[5831]));
    assign layer1_outputs[2818] = ~(layer0_outputs[9576]);
    assign layer1_outputs[2819] = ~((layer0_outputs[12795]) ^ (layer0_outputs[9641]));
    assign layer1_outputs[2820] = ~((layer0_outputs[11683]) | (layer0_outputs[2910]));
    assign layer1_outputs[2821] = ~(layer0_outputs[7296]) | (layer0_outputs[6293]);
    assign layer1_outputs[2822] = (layer0_outputs[12320]) & (layer0_outputs[3479]);
    assign layer1_outputs[2823] = ~(layer0_outputs[2052]);
    assign layer1_outputs[2824] = layer0_outputs[3050];
    assign layer1_outputs[2825] = (layer0_outputs[10938]) & (layer0_outputs[8116]);
    assign layer1_outputs[2826] = ~(layer0_outputs[1717]);
    assign layer1_outputs[2827] = 1'b1;
    assign layer1_outputs[2828] = (layer0_outputs[12478]) & ~(layer0_outputs[6636]);
    assign layer1_outputs[2829] = layer0_outputs[2829];
    assign layer1_outputs[2830] = ~(layer0_outputs[9856]) | (layer0_outputs[3471]);
    assign layer1_outputs[2831] = ~(layer0_outputs[6108]);
    assign layer1_outputs[2832] = ~(layer0_outputs[4946]);
    assign layer1_outputs[2833] = ~(layer0_outputs[8735]);
    assign layer1_outputs[2834] = ~((layer0_outputs[8869]) ^ (layer0_outputs[2368]));
    assign layer1_outputs[2835] = layer0_outputs[8843];
    assign layer1_outputs[2836] = ~((layer0_outputs[8846]) & (layer0_outputs[7164]));
    assign layer1_outputs[2837] = ~(layer0_outputs[2625]);
    assign layer1_outputs[2838] = ~(layer0_outputs[12186]);
    assign layer1_outputs[2839] = ~(layer0_outputs[7093]) | (layer0_outputs[2730]);
    assign layer1_outputs[2840] = ~(layer0_outputs[12378]);
    assign layer1_outputs[2841] = (layer0_outputs[8234]) ^ (layer0_outputs[4237]);
    assign layer1_outputs[2842] = layer0_outputs[11634];
    assign layer1_outputs[2843] = ~((layer0_outputs[4338]) ^ (layer0_outputs[1253]));
    assign layer1_outputs[2844] = (layer0_outputs[12339]) & ~(layer0_outputs[3084]);
    assign layer1_outputs[2845] = ~(layer0_outputs[7260]);
    assign layer1_outputs[2846] = ~(layer0_outputs[2650]);
    assign layer1_outputs[2847] = (layer0_outputs[8908]) & (layer0_outputs[3989]);
    assign layer1_outputs[2848] = layer0_outputs[8683];
    assign layer1_outputs[2849] = (layer0_outputs[4061]) & ~(layer0_outputs[1910]);
    assign layer1_outputs[2850] = (layer0_outputs[5744]) | (layer0_outputs[7690]);
    assign layer1_outputs[2851] = ~((layer0_outputs[6780]) | (layer0_outputs[5773]));
    assign layer1_outputs[2852] = ~(layer0_outputs[6656]) | (layer0_outputs[326]);
    assign layer1_outputs[2853] = ~(layer0_outputs[12559]);
    assign layer1_outputs[2854] = (layer0_outputs[6317]) & ~(layer0_outputs[10788]);
    assign layer1_outputs[2855] = layer0_outputs[348];
    assign layer1_outputs[2856] = ~((layer0_outputs[11657]) & (layer0_outputs[530]));
    assign layer1_outputs[2857] = layer0_outputs[12571];
    assign layer1_outputs[2858] = ~(layer0_outputs[8944]);
    assign layer1_outputs[2859] = layer0_outputs[11870];
    assign layer1_outputs[2860] = (layer0_outputs[2073]) & ~(layer0_outputs[11905]);
    assign layer1_outputs[2861] = ~(layer0_outputs[1161]);
    assign layer1_outputs[2862] = ~(layer0_outputs[10100]);
    assign layer1_outputs[2863] = (layer0_outputs[87]) ^ (layer0_outputs[5433]);
    assign layer1_outputs[2864] = layer0_outputs[3633];
    assign layer1_outputs[2865] = ~(layer0_outputs[8666]) | (layer0_outputs[12134]);
    assign layer1_outputs[2866] = layer0_outputs[11038];
    assign layer1_outputs[2867] = ~(layer0_outputs[9811]);
    assign layer1_outputs[2868] = ~(layer0_outputs[9364]) | (layer0_outputs[1733]);
    assign layer1_outputs[2869] = ~(layer0_outputs[3039]);
    assign layer1_outputs[2870] = ~(layer0_outputs[10888]);
    assign layer1_outputs[2871] = layer0_outputs[2727];
    assign layer1_outputs[2872] = ~(layer0_outputs[4268]) | (layer0_outputs[1472]);
    assign layer1_outputs[2873] = ~(layer0_outputs[6695]) | (layer0_outputs[2550]);
    assign layer1_outputs[2874] = 1'b1;
    assign layer1_outputs[2875] = (layer0_outputs[4496]) ^ (layer0_outputs[5670]);
    assign layer1_outputs[2876] = (layer0_outputs[7410]) & ~(layer0_outputs[2963]);
    assign layer1_outputs[2877] = ~(layer0_outputs[9332]);
    assign layer1_outputs[2878] = ~((layer0_outputs[5133]) | (layer0_outputs[4430]));
    assign layer1_outputs[2879] = (layer0_outputs[7515]) & (layer0_outputs[7718]);
    assign layer1_outputs[2880] = layer0_outputs[9532];
    assign layer1_outputs[2881] = (layer0_outputs[529]) | (layer0_outputs[249]);
    assign layer1_outputs[2882] = ~(layer0_outputs[11654]);
    assign layer1_outputs[2883] = (layer0_outputs[1963]) & ~(layer0_outputs[235]);
    assign layer1_outputs[2884] = (layer0_outputs[11721]) | (layer0_outputs[9955]);
    assign layer1_outputs[2885] = (layer0_outputs[4583]) ^ (layer0_outputs[4070]);
    assign layer1_outputs[2886] = ~((layer0_outputs[4572]) & (layer0_outputs[7531]));
    assign layer1_outputs[2887] = layer0_outputs[323];
    assign layer1_outputs[2888] = ~((layer0_outputs[3242]) | (layer0_outputs[10912]));
    assign layer1_outputs[2889] = ~(layer0_outputs[4416]) | (layer0_outputs[1535]);
    assign layer1_outputs[2890] = 1'b1;
    assign layer1_outputs[2891] = ~((layer0_outputs[515]) | (layer0_outputs[9565]));
    assign layer1_outputs[2892] = layer0_outputs[3895];
    assign layer1_outputs[2893] = (layer0_outputs[12659]) & ~(layer0_outputs[651]);
    assign layer1_outputs[2894] = ~(layer0_outputs[6104]);
    assign layer1_outputs[2895] = layer0_outputs[5896];
    assign layer1_outputs[2896] = (layer0_outputs[415]) | (layer0_outputs[5656]);
    assign layer1_outputs[2897] = (layer0_outputs[11876]) & ~(layer0_outputs[11910]);
    assign layer1_outputs[2898] = ~(layer0_outputs[8450]);
    assign layer1_outputs[2899] = ~(layer0_outputs[4562]) | (layer0_outputs[5653]);
    assign layer1_outputs[2900] = (layer0_outputs[9723]) & ~(layer0_outputs[6614]);
    assign layer1_outputs[2901] = ~((layer0_outputs[6738]) ^ (layer0_outputs[8814]));
    assign layer1_outputs[2902] = layer0_outputs[9963];
    assign layer1_outputs[2903] = ~((layer0_outputs[2419]) & (layer0_outputs[4540]));
    assign layer1_outputs[2904] = (layer0_outputs[5117]) & ~(layer0_outputs[8618]);
    assign layer1_outputs[2905] = ~(layer0_outputs[3812]) | (layer0_outputs[7962]);
    assign layer1_outputs[2906] = layer0_outputs[11356];
    assign layer1_outputs[2907] = ~((layer0_outputs[3284]) | (layer0_outputs[12794]));
    assign layer1_outputs[2908] = ~(layer0_outputs[6645]) | (layer0_outputs[1061]);
    assign layer1_outputs[2909] = (layer0_outputs[152]) & (layer0_outputs[5998]);
    assign layer1_outputs[2910] = ~(layer0_outputs[8474]);
    assign layer1_outputs[2911] = (layer0_outputs[12290]) & (layer0_outputs[5766]);
    assign layer1_outputs[2912] = layer0_outputs[5731];
    assign layer1_outputs[2913] = (layer0_outputs[6950]) | (layer0_outputs[11525]);
    assign layer1_outputs[2914] = ~(layer0_outputs[859]) | (layer0_outputs[12718]);
    assign layer1_outputs[2915] = layer0_outputs[6544];
    assign layer1_outputs[2916] = ~(layer0_outputs[822]);
    assign layer1_outputs[2917] = ~(layer0_outputs[520]) | (layer0_outputs[2560]);
    assign layer1_outputs[2918] = ~(layer0_outputs[1]);
    assign layer1_outputs[2919] = ~((layer0_outputs[830]) & (layer0_outputs[1581]));
    assign layer1_outputs[2920] = (layer0_outputs[8977]) | (layer0_outputs[1232]);
    assign layer1_outputs[2921] = ~(layer0_outputs[7803]);
    assign layer1_outputs[2922] = (layer0_outputs[6098]) | (layer0_outputs[309]);
    assign layer1_outputs[2923] = ~(layer0_outputs[2395]) | (layer0_outputs[11414]);
    assign layer1_outputs[2924] = ~(layer0_outputs[9836]);
    assign layer1_outputs[2925] = ~((layer0_outputs[11465]) | (layer0_outputs[12650]));
    assign layer1_outputs[2926] = (layer0_outputs[4728]) | (layer0_outputs[5205]);
    assign layer1_outputs[2927] = ~(layer0_outputs[1011]);
    assign layer1_outputs[2928] = (layer0_outputs[10711]) & (layer0_outputs[3779]);
    assign layer1_outputs[2929] = ~(layer0_outputs[12149]);
    assign layer1_outputs[2930] = 1'b0;
    assign layer1_outputs[2931] = (layer0_outputs[3324]) & ~(layer0_outputs[1701]);
    assign layer1_outputs[2932] = (layer0_outputs[9047]) & ~(layer0_outputs[2250]);
    assign layer1_outputs[2933] = ~(layer0_outputs[9383]) | (layer0_outputs[8532]);
    assign layer1_outputs[2934] = ~((layer0_outputs[6270]) ^ (layer0_outputs[1938]));
    assign layer1_outputs[2935] = 1'b0;
    assign layer1_outputs[2936] = ~((layer0_outputs[7232]) ^ (layer0_outputs[11553]));
    assign layer1_outputs[2937] = layer0_outputs[9181];
    assign layer1_outputs[2938] = ~(layer0_outputs[11732]);
    assign layer1_outputs[2939] = ~(layer0_outputs[1770]);
    assign layer1_outputs[2940] = (layer0_outputs[11291]) & (layer0_outputs[9500]);
    assign layer1_outputs[2941] = ~(layer0_outputs[5008]);
    assign layer1_outputs[2942] = layer0_outputs[11805];
    assign layer1_outputs[2943] = ~((layer0_outputs[9116]) ^ (layer0_outputs[9780]));
    assign layer1_outputs[2944] = (layer0_outputs[2693]) & ~(layer0_outputs[11443]);
    assign layer1_outputs[2945] = ~(layer0_outputs[1517]) | (layer0_outputs[11624]);
    assign layer1_outputs[2946] = ~(layer0_outputs[508]) | (layer0_outputs[6197]);
    assign layer1_outputs[2947] = ~(layer0_outputs[1986]);
    assign layer1_outputs[2948] = layer0_outputs[12154];
    assign layer1_outputs[2949] = ~(layer0_outputs[12150]) | (layer0_outputs[1454]);
    assign layer1_outputs[2950] = layer0_outputs[12579];
    assign layer1_outputs[2951] = ~(layer0_outputs[5229]);
    assign layer1_outputs[2952] = ~(layer0_outputs[9305]) | (layer0_outputs[4955]);
    assign layer1_outputs[2953] = (layer0_outputs[4241]) & ~(layer0_outputs[5120]);
    assign layer1_outputs[2954] = (layer0_outputs[7790]) ^ (layer0_outputs[4702]);
    assign layer1_outputs[2955] = layer0_outputs[4537];
    assign layer1_outputs[2956] = layer0_outputs[9900];
    assign layer1_outputs[2957] = ~(layer0_outputs[5558]);
    assign layer1_outputs[2958] = (layer0_outputs[1413]) & (layer0_outputs[5964]);
    assign layer1_outputs[2959] = (layer0_outputs[10677]) & ~(layer0_outputs[3322]);
    assign layer1_outputs[2960] = ~(layer0_outputs[11217]);
    assign layer1_outputs[2961] = layer0_outputs[11295];
    assign layer1_outputs[2962] = ~((layer0_outputs[8510]) & (layer0_outputs[12529]));
    assign layer1_outputs[2963] = ~(layer0_outputs[2037]);
    assign layer1_outputs[2964] = ~(layer0_outputs[4472]);
    assign layer1_outputs[2965] = layer0_outputs[9864];
    assign layer1_outputs[2966] = ~((layer0_outputs[8909]) | (layer0_outputs[1898]));
    assign layer1_outputs[2967] = ~(layer0_outputs[7378]);
    assign layer1_outputs[2968] = ~((layer0_outputs[11046]) & (layer0_outputs[2303]));
    assign layer1_outputs[2969] = (layer0_outputs[12294]) & ~(layer0_outputs[1805]);
    assign layer1_outputs[2970] = (layer0_outputs[706]) | (layer0_outputs[66]);
    assign layer1_outputs[2971] = (layer0_outputs[1931]) & ~(layer0_outputs[880]);
    assign layer1_outputs[2972] = ~(layer0_outputs[3826]) | (layer0_outputs[7664]);
    assign layer1_outputs[2973] = (layer0_outputs[2412]) & (layer0_outputs[241]);
    assign layer1_outputs[2974] = layer0_outputs[3941];
    assign layer1_outputs[2975] = layer0_outputs[6202];
    assign layer1_outputs[2976] = ~(layer0_outputs[5872]) | (layer0_outputs[7407]);
    assign layer1_outputs[2977] = (layer0_outputs[6984]) & ~(layer0_outputs[5579]);
    assign layer1_outputs[2978] = 1'b0;
    assign layer1_outputs[2979] = ~(layer0_outputs[5327]);
    assign layer1_outputs[2980] = layer0_outputs[10130];
    assign layer1_outputs[2981] = layer0_outputs[1229];
    assign layer1_outputs[2982] = (layer0_outputs[35]) & (layer0_outputs[1892]);
    assign layer1_outputs[2983] = ~(layer0_outputs[2057]);
    assign layer1_outputs[2984] = (layer0_outputs[4864]) & ~(layer0_outputs[9380]);
    assign layer1_outputs[2985] = ~((layer0_outputs[2323]) | (layer0_outputs[1188]));
    assign layer1_outputs[2986] = ~(layer0_outputs[3153]) | (layer0_outputs[12359]);
    assign layer1_outputs[2987] = (layer0_outputs[7191]) ^ (layer0_outputs[7799]);
    assign layer1_outputs[2988] = (layer0_outputs[11801]) & ~(layer0_outputs[90]);
    assign layer1_outputs[2989] = layer0_outputs[456];
    assign layer1_outputs[2990] = ~(layer0_outputs[9103]) | (layer0_outputs[6678]);
    assign layer1_outputs[2991] = ~(layer0_outputs[2042]) | (layer0_outputs[488]);
    assign layer1_outputs[2992] = layer0_outputs[1104];
    assign layer1_outputs[2993] = (layer0_outputs[9148]) & (layer0_outputs[9515]);
    assign layer1_outputs[2994] = ~((layer0_outputs[8343]) ^ (layer0_outputs[419]));
    assign layer1_outputs[2995] = ~((layer0_outputs[8925]) | (layer0_outputs[11502]));
    assign layer1_outputs[2996] = ~((layer0_outputs[4217]) & (layer0_outputs[7421]));
    assign layer1_outputs[2997] = layer0_outputs[9229];
    assign layer1_outputs[2998] = ~(layer0_outputs[12400]);
    assign layer1_outputs[2999] = ~((layer0_outputs[11570]) ^ (layer0_outputs[6744]));
    assign layer1_outputs[3000] = ~(layer0_outputs[2884]);
    assign layer1_outputs[3001] = layer0_outputs[2792];
    assign layer1_outputs[3002] = layer0_outputs[6709];
    assign layer1_outputs[3003] = ~((layer0_outputs[5933]) ^ (layer0_outputs[11850]));
    assign layer1_outputs[3004] = ~(layer0_outputs[5564]);
    assign layer1_outputs[3005] = (layer0_outputs[7217]) & ~(layer0_outputs[10927]);
    assign layer1_outputs[3006] = ~(layer0_outputs[11159]);
    assign layer1_outputs[3007] = ~(layer0_outputs[12324]) | (layer0_outputs[3576]);
    assign layer1_outputs[3008] = (layer0_outputs[3597]) & ~(layer0_outputs[11498]);
    assign layer1_outputs[3009] = layer0_outputs[11250];
    assign layer1_outputs[3010] = ~((layer0_outputs[3010]) | (layer0_outputs[7211]));
    assign layer1_outputs[3011] = 1'b0;
    assign layer1_outputs[3012] = (layer0_outputs[12169]) & (layer0_outputs[3656]);
    assign layer1_outputs[3013] = (layer0_outputs[6156]) & ~(layer0_outputs[6463]);
    assign layer1_outputs[3014] = ~(layer0_outputs[3017]) | (layer0_outputs[10013]);
    assign layer1_outputs[3015] = (layer0_outputs[11094]) & ~(layer0_outputs[3784]);
    assign layer1_outputs[3016] = (layer0_outputs[8844]) & ~(layer0_outputs[12479]);
    assign layer1_outputs[3017] = ~((layer0_outputs[935]) | (layer0_outputs[7785]));
    assign layer1_outputs[3018] = layer0_outputs[11372];
    assign layer1_outputs[3019] = ~(layer0_outputs[9050]) | (layer0_outputs[8385]);
    assign layer1_outputs[3020] = (layer0_outputs[1209]) & ~(layer0_outputs[1511]);
    assign layer1_outputs[3021] = ~(layer0_outputs[3379]);
    assign layer1_outputs[3022] = ~(layer0_outputs[10576]);
    assign layer1_outputs[3023] = ~(layer0_outputs[325]);
    assign layer1_outputs[3024] = ~(layer0_outputs[7086]) | (layer0_outputs[11463]);
    assign layer1_outputs[3025] = (layer0_outputs[10294]) & ~(layer0_outputs[2484]);
    assign layer1_outputs[3026] = (layer0_outputs[8865]) | (layer0_outputs[8421]);
    assign layer1_outputs[3027] = (layer0_outputs[4692]) & (layer0_outputs[7300]);
    assign layer1_outputs[3028] = (layer0_outputs[5572]) & (layer0_outputs[2427]);
    assign layer1_outputs[3029] = (layer0_outputs[5963]) & ~(layer0_outputs[12754]);
    assign layer1_outputs[3030] = (layer0_outputs[12132]) ^ (layer0_outputs[2713]);
    assign layer1_outputs[3031] = ~((layer0_outputs[6725]) & (layer0_outputs[6740]));
    assign layer1_outputs[3032] = ~(layer0_outputs[3494]) | (layer0_outputs[5568]);
    assign layer1_outputs[3033] = ~((layer0_outputs[1961]) | (layer0_outputs[9566]));
    assign layer1_outputs[3034] = layer0_outputs[5161];
    assign layer1_outputs[3035] = ~((layer0_outputs[2720]) ^ (layer0_outputs[316]));
    assign layer1_outputs[3036] = layer0_outputs[8397];
    assign layer1_outputs[3037] = ~((layer0_outputs[7183]) ^ (layer0_outputs[11519]));
    assign layer1_outputs[3038] = ~(layer0_outputs[9788]);
    assign layer1_outputs[3039] = (layer0_outputs[4535]) | (layer0_outputs[3956]);
    assign layer1_outputs[3040] = ~(layer0_outputs[4352]);
    assign layer1_outputs[3041] = ~((layer0_outputs[2164]) | (layer0_outputs[1947]));
    assign layer1_outputs[3042] = (layer0_outputs[6403]) & ~(layer0_outputs[10577]);
    assign layer1_outputs[3043] = ~((layer0_outputs[4673]) ^ (layer0_outputs[530]));
    assign layer1_outputs[3044] = ~(layer0_outputs[10434]);
    assign layer1_outputs[3045] = (layer0_outputs[4718]) & (layer0_outputs[8904]);
    assign layer1_outputs[3046] = ~((layer0_outputs[2915]) | (layer0_outputs[8149]));
    assign layer1_outputs[3047] = (layer0_outputs[10085]) & ~(layer0_outputs[613]);
    assign layer1_outputs[3048] = ~(layer0_outputs[7261]);
    assign layer1_outputs[3049] = layer0_outputs[9146];
    assign layer1_outputs[3050] = layer0_outputs[7034];
    assign layer1_outputs[3051] = 1'b0;
    assign layer1_outputs[3052] = (layer0_outputs[5094]) & ~(layer0_outputs[1307]);
    assign layer1_outputs[3053] = layer0_outputs[2283];
    assign layer1_outputs[3054] = ~((layer0_outputs[11599]) | (layer0_outputs[5776]));
    assign layer1_outputs[3055] = ~(layer0_outputs[5902]);
    assign layer1_outputs[3056] = ~(layer0_outputs[5036]);
    assign layer1_outputs[3057] = layer0_outputs[403];
    assign layer1_outputs[3058] = (layer0_outputs[10909]) ^ (layer0_outputs[11961]);
    assign layer1_outputs[3059] = ~((layer0_outputs[6249]) ^ (layer0_outputs[5596]));
    assign layer1_outputs[3060] = ~(layer0_outputs[1434]) | (layer0_outputs[5067]);
    assign layer1_outputs[3061] = ~((layer0_outputs[8445]) | (layer0_outputs[4341]));
    assign layer1_outputs[3062] = layer0_outputs[4605];
    assign layer1_outputs[3063] = 1'b1;
    assign layer1_outputs[3064] = ~((layer0_outputs[9316]) & (layer0_outputs[6559]));
    assign layer1_outputs[3065] = layer0_outputs[8889];
    assign layer1_outputs[3066] = ~(layer0_outputs[1275]);
    assign layer1_outputs[3067] = layer0_outputs[722];
    assign layer1_outputs[3068] = 1'b1;
    assign layer1_outputs[3069] = (layer0_outputs[6305]) ^ (layer0_outputs[4283]);
    assign layer1_outputs[3070] = ~(layer0_outputs[10016]);
    assign layer1_outputs[3071] = (layer0_outputs[1903]) & (layer0_outputs[3772]);
    assign layer1_outputs[3072] = ~((layer0_outputs[12268]) | (layer0_outputs[11632]));
    assign layer1_outputs[3073] = ~(layer0_outputs[6958]);
    assign layer1_outputs[3074] = (layer0_outputs[11442]) ^ (layer0_outputs[572]);
    assign layer1_outputs[3075] = 1'b1;
    assign layer1_outputs[3076] = ~((layer0_outputs[8076]) | (layer0_outputs[2306]));
    assign layer1_outputs[3077] = layer0_outputs[12295];
    assign layer1_outputs[3078] = ~((layer0_outputs[8847]) & (layer0_outputs[11969]));
    assign layer1_outputs[3079] = ~((layer0_outputs[3015]) ^ (layer0_outputs[10446]));
    assign layer1_outputs[3080] = ~(layer0_outputs[4651]) | (layer0_outputs[7384]);
    assign layer1_outputs[3081] = ~((layer0_outputs[1919]) & (layer0_outputs[8177]));
    assign layer1_outputs[3082] = ~(layer0_outputs[4337]);
    assign layer1_outputs[3083] = ~(layer0_outputs[5193]);
    assign layer1_outputs[3084] = ~(layer0_outputs[5772]);
    assign layer1_outputs[3085] = (layer0_outputs[397]) & ~(layer0_outputs[10972]);
    assign layer1_outputs[3086] = ~(layer0_outputs[7503]) | (layer0_outputs[12748]);
    assign layer1_outputs[3087] = ~(layer0_outputs[11942]);
    assign layer1_outputs[3088] = (layer0_outputs[6893]) & ~(layer0_outputs[6878]);
    assign layer1_outputs[3089] = (layer0_outputs[10955]) & ~(layer0_outputs[6185]);
    assign layer1_outputs[3090] = layer0_outputs[11100];
    assign layer1_outputs[3091] = (layer0_outputs[10069]) | (layer0_outputs[9587]);
    assign layer1_outputs[3092] = ~(layer0_outputs[9560]) | (layer0_outputs[6615]);
    assign layer1_outputs[3093] = layer0_outputs[1152];
    assign layer1_outputs[3094] = ~(layer0_outputs[12215]);
    assign layer1_outputs[3095] = (layer0_outputs[8523]) & (layer0_outputs[10474]);
    assign layer1_outputs[3096] = ~(layer0_outputs[9212]);
    assign layer1_outputs[3097] = (layer0_outputs[592]) & ~(layer0_outputs[7710]);
    assign layer1_outputs[3098] = (layer0_outputs[444]) & (layer0_outputs[2434]);
    assign layer1_outputs[3099] = ~(layer0_outputs[11308]) | (layer0_outputs[10919]);
    assign layer1_outputs[3100] = ~(layer0_outputs[6934]) | (layer0_outputs[373]);
    assign layer1_outputs[3101] = ~(layer0_outputs[8381]) | (layer0_outputs[6659]);
    assign layer1_outputs[3102] = ~((layer0_outputs[12604]) & (layer0_outputs[8080]));
    assign layer1_outputs[3103] = ~((layer0_outputs[6772]) ^ (layer0_outputs[5077]));
    assign layer1_outputs[3104] = 1'b1;
    assign layer1_outputs[3105] = ~(layer0_outputs[11794]) | (layer0_outputs[3911]);
    assign layer1_outputs[3106] = ~((layer0_outputs[4472]) ^ (layer0_outputs[4618]));
    assign layer1_outputs[3107] = (layer0_outputs[12181]) & (layer0_outputs[4547]);
    assign layer1_outputs[3108] = ~(layer0_outputs[6273]);
    assign layer1_outputs[3109] = 1'b0;
    assign layer1_outputs[3110] = ~(layer0_outputs[6578]);
    assign layer1_outputs[3111] = ~((layer0_outputs[7653]) | (layer0_outputs[1643]));
    assign layer1_outputs[3112] = ~(layer0_outputs[7223]);
    assign layer1_outputs[3113] = (layer0_outputs[2197]) | (layer0_outputs[7722]);
    assign layer1_outputs[3114] = (layer0_outputs[6480]) & (layer0_outputs[2538]);
    assign layer1_outputs[3115] = layer0_outputs[7136];
    assign layer1_outputs[3116] = ~((layer0_outputs[4669]) | (layer0_outputs[5051]));
    assign layer1_outputs[3117] = ~(layer0_outputs[9300]);
    assign layer1_outputs[3118] = (layer0_outputs[6578]) ^ (layer0_outputs[2785]);
    assign layer1_outputs[3119] = ~(layer0_outputs[11893]);
    assign layer1_outputs[3120] = ~(layer0_outputs[11056]) | (layer0_outputs[3438]);
    assign layer1_outputs[3121] = 1'b0;
    assign layer1_outputs[3122] = layer0_outputs[5891];
    assign layer1_outputs[3123] = layer0_outputs[3532];
    assign layer1_outputs[3124] = ~(layer0_outputs[4868]) | (layer0_outputs[10134]);
    assign layer1_outputs[3125] = layer0_outputs[12059];
    assign layer1_outputs[3126] = (layer0_outputs[1975]) & (layer0_outputs[8637]);
    assign layer1_outputs[3127] = (layer0_outputs[3185]) ^ (layer0_outputs[1470]);
    assign layer1_outputs[3128] = (layer0_outputs[10812]) & (layer0_outputs[6612]);
    assign layer1_outputs[3129] = layer0_outputs[8613];
    assign layer1_outputs[3130] = ~((layer0_outputs[7136]) | (layer0_outputs[5377]));
    assign layer1_outputs[3131] = ~(layer0_outputs[2841]);
    assign layer1_outputs[3132] = 1'b1;
    assign layer1_outputs[3133] = ~((layer0_outputs[12140]) | (layer0_outputs[1484]));
    assign layer1_outputs[3134] = ~((layer0_outputs[5953]) & (layer0_outputs[67]));
    assign layer1_outputs[3135] = layer0_outputs[10971];
    assign layer1_outputs[3136] = ~(layer0_outputs[11785]);
    assign layer1_outputs[3137] = (layer0_outputs[7106]) | (layer0_outputs[7960]);
    assign layer1_outputs[3138] = ~(layer0_outputs[4232]) | (layer0_outputs[12549]);
    assign layer1_outputs[3139] = ~((layer0_outputs[6293]) | (layer0_outputs[7882]));
    assign layer1_outputs[3140] = ~((layer0_outputs[2293]) | (layer0_outputs[1154]));
    assign layer1_outputs[3141] = layer0_outputs[1299];
    assign layer1_outputs[3142] = (layer0_outputs[10998]) & ~(layer0_outputs[12076]);
    assign layer1_outputs[3143] = ~((layer0_outputs[2795]) | (layer0_outputs[4814]));
    assign layer1_outputs[3144] = (layer0_outputs[2850]) & ~(layer0_outputs[7636]);
    assign layer1_outputs[3145] = (layer0_outputs[478]) ^ (layer0_outputs[12348]);
    assign layer1_outputs[3146] = ~((layer0_outputs[11741]) ^ (layer0_outputs[7269]));
    assign layer1_outputs[3147] = 1'b1;
    assign layer1_outputs[3148] = (layer0_outputs[10362]) & ~(layer0_outputs[5748]);
    assign layer1_outputs[3149] = ~(layer0_outputs[222]);
    assign layer1_outputs[3150] = ~(layer0_outputs[325]);
    assign layer1_outputs[3151] = (layer0_outputs[2990]) & ~(layer0_outputs[9480]);
    assign layer1_outputs[3152] = ~(layer0_outputs[1384]);
    assign layer1_outputs[3153] = ~(layer0_outputs[3874]);
    assign layer1_outputs[3154] = ~(layer0_outputs[9979]);
    assign layer1_outputs[3155] = layer0_outputs[10217];
    assign layer1_outputs[3156] = layer0_outputs[12100];
    assign layer1_outputs[3157] = (layer0_outputs[12061]) | (layer0_outputs[2119]);
    assign layer1_outputs[3158] = ~(layer0_outputs[9030]);
    assign layer1_outputs[3159] = (layer0_outputs[12038]) ^ (layer0_outputs[10853]);
    assign layer1_outputs[3160] = (layer0_outputs[5673]) & (layer0_outputs[8141]);
    assign layer1_outputs[3161] = ~(layer0_outputs[8495]) | (layer0_outputs[4744]);
    assign layer1_outputs[3162] = layer0_outputs[10731];
    assign layer1_outputs[3163] = 1'b0;
    assign layer1_outputs[3164] = (layer0_outputs[4588]) ^ (layer0_outputs[1854]);
    assign layer1_outputs[3165] = (layer0_outputs[9530]) & (layer0_outputs[9124]);
    assign layer1_outputs[3166] = ~(layer0_outputs[3869]);
    assign layer1_outputs[3167] = layer0_outputs[5761];
    assign layer1_outputs[3168] = ~((layer0_outputs[2740]) ^ (layer0_outputs[7028]));
    assign layer1_outputs[3169] = (layer0_outputs[5813]) & ~(layer0_outputs[194]);
    assign layer1_outputs[3170] = layer0_outputs[7344];
    assign layer1_outputs[3171] = (layer0_outputs[1507]) ^ (layer0_outputs[9238]);
    assign layer1_outputs[3172] = ~((layer0_outputs[7376]) ^ (layer0_outputs[5636]));
    assign layer1_outputs[3173] = (layer0_outputs[10596]) & ~(layer0_outputs[6148]);
    assign layer1_outputs[3174] = ~(layer0_outputs[3333]);
    assign layer1_outputs[3175] = (layer0_outputs[4507]) & (layer0_outputs[443]);
    assign layer1_outputs[3176] = ~(layer0_outputs[11185]) | (layer0_outputs[7060]);
    assign layer1_outputs[3177] = ~((layer0_outputs[12476]) ^ (layer0_outputs[3298]));
    assign layer1_outputs[3178] = ~(layer0_outputs[4456]);
    assign layer1_outputs[3179] = layer0_outputs[1649];
    assign layer1_outputs[3180] = ~((layer0_outputs[9948]) | (layer0_outputs[4440]));
    assign layer1_outputs[3181] = (layer0_outputs[2078]) & (layer0_outputs[8133]);
    assign layer1_outputs[3182] = ~(layer0_outputs[1685]) | (layer0_outputs[2513]);
    assign layer1_outputs[3183] = 1'b0;
    assign layer1_outputs[3184] = ~((layer0_outputs[6200]) & (layer0_outputs[10091]));
    assign layer1_outputs[3185] = (layer0_outputs[8986]) | (layer0_outputs[5593]);
    assign layer1_outputs[3186] = layer0_outputs[7201];
    assign layer1_outputs[3187] = ~(layer0_outputs[12162]);
    assign layer1_outputs[3188] = 1'b0;
    assign layer1_outputs[3189] = ~((layer0_outputs[9485]) ^ (layer0_outputs[796]));
    assign layer1_outputs[3190] = ~((layer0_outputs[11757]) & (layer0_outputs[8757]));
    assign layer1_outputs[3191] = layer0_outputs[2694];
    assign layer1_outputs[3192] = ~((layer0_outputs[2919]) | (layer0_outputs[3170]));
    assign layer1_outputs[3193] = (layer0_outputs[2652]) | (layer0_outputs[6104]);
    assign layer1_outputs[3194] = (layer0_outputs[6915]) & (layer0_outputs[6822]);
    assign layer1_outputs[3195] = ~(layer0_outputs[4810]) | (layer0_outputs[6835]);
    assign layer1_outputs[3196] = (layer0_outputs[3684]) ^ (layer0_outputs[8121]);
    assign layer1_outputs[3197] = layer0_outputs[9571];
    assign layer1_outputs[3198] = ~(layer0_outputs[2591]);
    assign layer1_outputs[3199] = layer0_outputs[4681];
    assign layer1_outputs[3200] = ~((layer0_outputs[7210]) | (layer0_outputs[11305]));
    assign layer1_outputs[3201] = ~(layer0_outputs[11280]) | (layer0_outputs[10040]);
    assign layer1_outputs[3202] = layer0_outputs[10529];
    assign layer1_outputs[3203] = ~((layer0_outputs[2979]) & (layer0_outputs[53]));
    assign layer1_outputs[3204] = (layer0_outputs[2220]) & ~(layer0_outputs[259]);
    assign layer1_outputs[3205] = ~((layer0_outputs[11321]) | (layer0_outputs[10038]));
    assign layer1_outputs[3206] = layer0_outputs[2399];
    assign layer1_outputs[3207] = ~(layer0_outputs[12282]);
    assign layer1_outputs[3208] = layer0_outputs[7911];
    assign layer1_outputs[3209] = ~(layer0_outputs[1877]);
    assign layer1_outputs[3210] = ~((layer0_outputs[6181]) ^ (layer0_outputs[709]));
    assign layer1_outputs[3211] = ~(layer0_outputs[6164]) | (layer0_outputs[12256]);
    assign layer1_outputs[3212] = ~(layer0_outputs[2084]) | (layer0_outputs[4980]);
    assign layer1_outputs[3213] = ~(layer0_outputs[9097]);
    assign layer1_outputs[3214] = (layer0_outputs[913]) & ~(layer0_outputs[7791]);
    assign layer1_outputs[3215] = layer0_outputs[1119];
    assign layer1_outputs[3216] = ~((layer0_outputs[4340]) & (layer0_outputs[7323]));
    assign layer1_outputs[3217] = layer0_outputs[2546];
    assign layer1_outputs[3218] = ~(layer0_outputs[8246]) | (layer0_outputs[10339]);
    assign layer1_outputs[3219] = ~((layer0_outputs[489]) & (layer0_outputs[10084]));
    assign layer1_outputs[3220] = layer0_outputs[10782];
    assign layer1_outputs[3221] = layer0_outputs[8047];
    assign layer1_outputs[3222] = (layer0_outputs[8507]) ^ (layer0_outputs[8254]);
    assign layer1_outputs[3223] = ~(layer0_outputs[4602]);
    assign layer1_outputs[3224] = (layer0_outputs[8336]) ^ (layer0_outputs[1171]);
    assign layer1_outputs[3225] = ~(layer0_outputs[6819]);
    assign layer1_outputs[3226] = (layer0_outputs[2366]) | (layer0_outputs[11094]);
    assign layer1_outputs[3227] = ~(layer0_outputs[7017]);
    assign layer1_outputs[3228] = ~((layer0_outputs[9529]) | (layer0_outputs[677]));
    assign layer1_outputs[3229] = (layer0_outputs[6123]) | (layer0_outputs[4560]);
    assign layer1_outputs[3230] = (layer0_outputs[1263]) ^ (layer0_outputs[2669]);
    assign layer1_outputs[3231] = (layer0_outputs[593]) | (layer0_outputs[805]);
    assign layer1_outputs[3232] = ~(layer0_outputs[8147]);
    assign layer1_outputs[3233] = ~(layer0_outputs[2639]) | (layer0_outputs[2356]);
    assign layer1_outputs[3234] = ~((layer0_outputs[876]) ^ (layer0_outputs[5775]));
    assign layer1_outputs[3235] = (layer0_outputs[10063]) & ~(layer0_outputs[6476]);
    assign layer1_outputs[3236] = ~(layer0_outputs[5286]);
    assign layer1_outputs[3237] = layer0_outputs[824];
    assign layer1_outputs[3238] = ~(layer0_outputs[5867]);
    assign layer1_outputs[3239] = ~(layer0_outputs[12496]) | (layer0_outputs[11386]);
    assign layer1_outputs[3240] = (layer0_outputs[9219]) & ~(layer0_outputs[10257]);
    assign layer1_outputs[3241] = ~((layer0_outputs[11877]) & (layer0_outputs[10949]));
    assign layer1_outputs[3242] = ~((layer0_outputs[6275]) | (layer0_outputs[11445]));
    assign layer1_outputs[3243] = ~(layer0_outputs[4469]);
    assign layer1_outputs[3244] = (layer0_outputs[12326]) ^ (layer0_outputs[4645]);
    assign layer1_outputs[3245] = ~(layer0_outputs[9108]);
    assign layer1_outputs[3246] = layer0_outputs[1218];
    assign layer1_outputs[3247] = ~(layer0_outputs[6540]);
    assign layer1_outputs[3248] = (layer0_outputs[9508]) & ~(layer0_outputs[11406]);
    assign layer1_outputs[3249] = layer0_outputs[948];
    assign layer1_outputs[3250] = ~(layer0_outputs[290]);
    assign layer1_outputs[3251] = (layer0_outputs[3277]) & ~(layer0_outputs[8900]);
    assign layer1_outputs[3252] = ~((layer0_outputs[9191]) & (layer0_outputs[7097]));
    assign layer1_outputs[3253] = layer0_outputs[647];
    assign layer1_outputs[3254] = (layer0_outputs[10268]) & ~(layer0_outputs[8648]);
    assign layer1_outputs[3255] = (layer0_outputs[6990]) & ~(layer0_outputs[5533]);
    assign layer1_outputs[3256] = layer0_outputs[6637];
    assign layer1_outputs[3257] = ~(layer0_outputs[7574]);
    assign layer1_outputs[3258] = ~(layer0_outputs[11177]);
    assign layer1_outputs[3259] = ~((layer0_outputs[9280]) ^ (layer0_outputs[3467]));
    assign layer1_outputs[3260] = layer0_outputs[4349];
    assign layer1_outputs[3261] = ~((layer0_outputs[3842]) | (layer0_outputs[481]));
    assign layer1_outputs[3262] = (layer0_outputs[801]) & ~(layer0_outputs[1232]);
    assign layer1_outputs[3263] = ~((layer0_outputs[4105]) | (layer0_outputs[9136]));
    assign layer1_outputs[3264] = 1'b0;
    assign layer1_outputs[3265] = layer0_outputs[3153];
    assign layer1_outputs[3266] = (layer0_outputs[4821]) & ~(layer0_outputs[10357]);
    assign layer1_outputs[3267] = ~((layer0_outputs[11651]) & (layer0_outputs[12703]));
    assign layer1_outputs[3268] = ~(layer0_outputs[6016]);
    assign layer1_outputs[3269] = ~(layer0_outputs[11598]) | (layer0_outputs[10641]);
    assign layer1_outputs[3270] = (layer0_outputs[10937]) & ~(layer0_outputs[10147]);
    assign layer1_outputs[3271] = (layer0_outputs[102]) & ~(layer0_outputs[4681]);
    assign layer1_outputs[3272] = (layer0_outputs[9325]) & ~(layer0_outputs[9838]);
    assign layer1_outputs[3273] = ~(layer0_outputs[2348]) | (layer0_outputs[1160]);
    assign layer1_outputs[3274] = ~((layer0_outputs[8628]) | (layer0_outputs[9177]));
    assign layer1_outputs[3275] = layer0_outputs[934];
    assign layer1_outputs[3276] = 1'b1;
    assign layer1_outputs[3277] = ~(layer0_outputs[54]) | (layer0_outputs[7709]);
    assign layer1_outputs[3278] = layer0_outputs[1602];
    assign layer1_outputs[3279] = (layer0_outputs[6580]) & ~(layer0_outputs[3315]);
    assign layer1_outputs[3280] = ~(layer0_outputs[10083]) | (layer0_outputs[10618]);
    assign layer1_outputs[3281] = layer0_outputs[12444];
    assign layer1_outputs[3282] = (layer0_outputs[7556]) ^ (layer0_outputs[2143]);
    assign layer1_outputs[3283] = layer0_outputs[11766];
    assign layer1_outputs[3284] = layer0_outputs[1402];
    assign layer1_outputs[3285] = layer0_outputs[12239];
    assign layer1_outputs[3286] = ~((layer0_outputs[10051]) | (layer0_outputs[1123]));
    assign layer1_outputs[3287] = layer0_outputs[4577];
    assign layer1_outputs[3288] = layer0_outputs[9355];
    assign layer1_outputs[3289] = ~((layer0_outputs[3329]) & (layer0_outputs[7764]));
    assign layer1_outputs[3290] = ~(layer0_outputs[7277]);
    assign layer1_outputs[3291] = layer0_outputs[5815];
    assign layer1_outputs[3292] = (layer0_outputs[7079]) ^ (layer0_outputs[705]);
    assign layer1_outputs[3293] = ~(layer0_outputs[1834]) | (layer0_outputs[6115]);
    assign layer1_outputs[3294] = ~((layer0_outputs[9700]) & (layer0_outputs[2445]));
    assign layer1_outputs[3295] = ~((layer0_outputs[6416]) | (layer0_outputs[11200]));
    assign layer1_outputs[3296] = (layer0_outputs[1420]) ^ (layer0_outputs[11198]);
    assign layer1_outputs[3297] = layer0_outputs[770];
    assign layer1_outputs[3298] = (layer0_outputs[3917]) | (layer0_outputs[9921]);
    assign layer1_outputs[3299] = ~(layer0_outputs[12102]);
    assign layer1_outputs[3300] = layer0_outputs[4141];
    assign layer1_outputs[3301] = ~((layer0_outputs[3672]) & (layer0_outputs[847]));
    assign layer1_outputs[3302] = ~((layer0_outputs[8430]) | (layer0_outputs[4457]));
    assign layer1_outputs[3303] = ~((layer0_outputs[8469]) ^ (layer0_outputs[10381]));
    assign layer1_outputs[3304] = layer0_outputs[10287];
    assign layer1_outputs[3305] = (layer0_outputs[4953]) | (layer0_outputs[12180]);
    assign layer1_outputs[3306] = layer0_outputs[6322];
    assign layer1_outputs[3307] = (layer0_outputs[11226]) | (layer0_outputs[8758]);
    assign layer1_outputs[3308] = (layer0_outputs[4825]) ^ (layer0_outputs[8443]);
    assign layer1_outputs[3309] = ~(layer0_outputs[8949]);
    assign layer1_outputs[3310] = ~(layer0_outputs[7268]) | (layer0_outputs[8033]);
    assign layer1_outputs[3311] = layer0_outputs[2530];
    assign layer1_outputs[3312] = 1'b1;
    assign layer1_outputs[3313] = (layer0_outputs[8049]) | (layer0_outputs[10573]);
    assign layer1_outputs[3314] = ~((layer0_outputs[2390]) ^ (layer0_outputs[3236]));
    assign layer1_outputs[3315] = ~((layer0_outputs[2950]) ^ (layer0_outputs[4699]));
    assign layer1_outputs[3316] = layer0_outputs[5204];
    assign layer1_outputs[3317] = (layer0_outputs[5128]) & ~(layer0_outputs[424]);
    assign layer1_outputs[3318] = (layer0_outputs[11348]) | (layer0_outputs[9111]);
    assign layer1_outputs[3319] = ~(layer0_outputs[2766]);
    assign layer1_outputs[3320] = (layer0_outputs[4682]) & ~(layer0_outputs[4358]);
    assign layer1_outputs[3321] = ~((layer0_outputs[4789]) & (layer0_outputs[9360]));
    assign layer1_outputs[3322] = ~(layer0_outputs[2783]);
    assign layer1_outputs[3323] = layer0_outputs[11849];
    assign layer1_outputs[3324] = ~(layer0_outputs[7115]) | (layer0_outputs[7454]);
    assign layer1_outputs[3325] = ~(layer0_outputs[8466]);
    assign layer1_outputs[3326] = ~((layer0_outputs[6752]) | (layer0_outputs[5905]));
    assign layer1_outputs[3327] = layer0_outputs[3495];
    assign layer1_outputs[3328] = ~(layer0_outputs[9411]) | (layer0_outputs[62]);
    assign layer1_outputs[3329] = layer0_outputs[3051];
    assign layer1_outputs[3330] = ~(layer0_outputs[11062]) | (layer0_outputs[8265]);
    assign layer1_outputs[3331] = ~(layer0_outputs[11479]) | (layer0_outputs[3427]);
    assign layer1_outputs[3332] = (layer0_outputs[6103]) ^ (layer0_outputs[9451]);
    assign layer1_outputs[3333] = ~(layer0_outputs[2940]) | (layer0_outputs[1801]);
    assign layer1_outputs[3334] = ~(layer0_outputs[1248]);
    assign layer1_outputs[3335] = ~(layer0_outputs[6560]);
    assign layer1_outputs[3336] = 1'b1;
    assign layer1_outputs[3337] = ~((layer0_outputs[461]) & (layer0_outputs[4951]));
    assign layer1_outputs[3338] = (layer0_outputs[12522]) | (layer0_outputs[2240]);
    assign layer1_outputs[3339] = ~(layer0_outputs[2695]);
    assign layer1_outputs[3340] = layer0_outputs[8701];
    assign layer1_outputs[3341] = layer0_outputs[9673];
    assign layer1_outputs[3342] = ~(layer0_outputs[12635]) | (layer0_outputs[3144]);
    assign layer1_outputs[3343] = (layer0_outputs[11436]) & (layer0_outputs[10563]);
    assign layer1_outputs[3344] = ~(layer0_outputs[12361]) | (layer0_outputs[2765]);
    assign layer1_outputs[3345] = ~((layer0_outputs[6185]) | (layer0_outputs[11236]));
    assign layer1_outputs[3346] = layer0_outputs[3502];
    assign layer1_outputs[3347] = ~(layer0_outputs[9159]);
    assign layer1_outputs[3348] = layer0_outputs[1609];
    assign layer1_outputs[3349] = (layer0_outputs[5291]) | (layer0_outputs[901]);
    assign layer1_outputs[3350] = ~((layer0_outputs[12091]) ^ (layer0_outputs[1301]));
    assign layer1_outputs[3351] = layer0_outputs[8022];
    assign layer1_outputs[3352] = ~(layer0_outputs[4374]) | (layer0_outputs[875]);
    assign layer1_outputs[3353] = ~(layer0_outputs[11309]);
    assign layer1_outputs[3354] = ~((layer0_outputs[6826]) | (layer0_outputs[9709]));
    assign layer1_outputs[3355] = ~((layer0_outputs[2308]) | (layer0_outputs[2019]));
    assign layer1_outputs[3356] = ~(layer0_outputs[1361]);
    assign layer1_outputs[3357] = (layer0_outputs[2864]) & (layer0_outputs[3623]);
    assign layer1_outputs[3358] = (layer0_outputs[12195]) & ~(layer0_outputs[11771]);
    assign layer1_outputs[3359] = ~((layer0_outputs[3187]) | (layer0_outputs[8707]));
    assign layer1_outputs[3360] = layer0_outputs[11368];
    assign layer1_outputs[3361] = (layer0_outputs[6121]) ^ (layer0_outputs[8464]);
    assign layer1_outputs[3362] = ~(layer0_outputs[4075]);
    assign layer1_outputs[3363] = (layer0_outputs[1266]) & ~(layer0_outputs[4658]);
    assign layer1_outputs[3364] = ~((layer0_outputs[251]) ^ (layer0_outputs[2101]));
    assign layer1_outputs[3365] = ~((layer0_outputs[5437]) | (layer0_outputs[9216]));
    assign layer1_outputs[3366] = layer0_outputs[4180];
    assign layer1_outputs[3367] = ~((layer0_outputs[1271]) | (layer0_outputs[9210]));
    assign layer1_outputs[3368] = ~(layer0_outputs[2628]);
    assign layer1_outputs[3369] = (layer0_outputs[933]) & ~(layer0_outputs[12763]);
    assign layer1_outputs[3370] = ~(layer0_outputs[6088]);
    assign layer1_outputs[3371] = layer0_outputs[10889];
    assign layer1_outputs[3372] = (layer0_outputs[7076]) & ~(layer0_outputs[4812]);
    assign layer1_outputs[3373] = (layer0_outputs[9260]) & (layer0_outputs[4763]);
    assign layer1_outputs[3374] = layer0_outputs[9858];
    assign layer1_outputs[3375] = (layer0_outputs[3961]) ^ (layer0_outputs[9427]);
    assign layer1_outputs[3376] = ~((layer0_outputs[4545]) & (layer0_outputs[9031]));
    assign layer1_outputs[3377] = layer0_outputs[4151];
    assign layer1_outputs[3378] = ~(layer0_outputs[5136]);
    assign layer1_outputs[3379] = (layer0_outputs[6575]) | (layer0_outputs[183]);
    assign layer1_outputs[3380] = ~(layer0_outputs[5749]);
    assign layer1_outputs[3381] = ~((layer0_outputs[3402]) | (layer0_outputs[12005]));
    assign layer1_outputs[3382] = ~((layer0_outputs[11135]) ^ (layer0_outputs[7650]));
    assign layer1_outputs[3383] = (layer0_outputs[883]) ^ (layer0_outputs[392]);
    assign layer1_outputs[3384] = ~(layer0_outputs[11683]) | (layer0_outputs[10994]);
    assign layer1_outputs[3385] = ~(layer0_outputs[2252]);
    assign layer1_outputs[3386] = ~(layer0_outputs[9975]);
    assign layer1_outputs[3387] = layer0_outputs[9003];
    assign layer1_outputs[3388] = 1'b0;
    assign layer1_outputs[3389] = ~(layer0_outputs[9497]);
    assign layer1_outputs[3390] = (layer0_outputs[9568]) & (layer0_outputs[3741]);
    assign layer1_outputs[3391] = layer0_outputs[6111];
    assign layer1_outputs[3392] = ~(layer0_outputs[7429]);
    assign layer1_outputs[3393] = (layer0_outputs[11283]) & ~(layer0_outputs[6956]);
    assign layer1_outputs[3394] = ~((layer0_outputs[528]) ^ (layer0_outputs[1241]));
    assign layer1_outputs[3395] = ~(layer0_outputs[10282]);
    assign layer1_outputs[3396] = (layer0_outputs[7241]) & ~(layer0_outputs[9883]);
    assign layer1_outputs[3397] = ~(layer0_outputs[12497]);
    assign layer1_outputs[3398] = (layer0_outputs[3686]) & ~(layer0_outputs[5846]);
    assign layer1_outputs[3399] = ~((layer0_outputs[3580]) & (layer0_outputs[5066]));
    assign layer1_outputs[3400] = (layer0_outputs[1842]) & (layer0_outputs[11314]);
    assign layer1_outputs[3401] = layer0_outputs[4341];
    assign layer1_outputs[3402] = (layer0_outputs[5766]) | (layer0_outputs[9759]);
    assign layer1_outputs[3403] = (layer0_outputs[8267]) & ~(layer0_outputs[9959]);
    assign layer1_outputs[3404] = ~(layer0_outputs[10897]) | (layer0_outputs[10728]);
    assign layer1_outputs[3405] = layer0_outputs[12703];
    assign layer1_outputs[3406] = ~(layer0_outputs[7370]) | (layer0_outputs[8086]);
    assign layer1_outputs[3407] = (layer0_outputs[9849]) | (layer0_outputs[2942]);
    assign layer1_outputs[3408] = (layer0_outputs[10754]) & ~(layer0_outputs[4616]);
    assign layer1_outputs[3409] = ~((layer0_outputs[8731]) ^ (layer0_outputs[832]));
    assign layer1_outputs[3410] = (layer0_outputs[5834]) & (layer0_outputs[10165]);
    assign layer1_outputs[3411] = layer0_outputs[12011];
    assign layer1_outputs[3412] = 1'b0;
    assign layer1_outputs[3413] = ~(layer0_outputs[7075]);
    assign layer1_outputs[3414] = ~(layer0_outputs[7144]) | (layer0_outputs[10784]);
    assign layer1_outputs[3415] = ~((layer0_outputs[1568]) & (layer0_outputs[3562]));
    assign layer1_outputs[3416] = (layer0_outputs[6155]) & ~(layer0_outputs[12784]);
    assign layer1_outputs[3417] = ~(layer0_outputs[4352]);
    assign layer1_outputs[3418] = ~(layer0_outputs[7288]) | (layer0_outputs[10004]);
    assign layer1_outputs[3419] = ~(layer0_outputs[7337]) | (layer0_outputs[6118]);
    assign layer1_outputs[3420] = ~(layer0_outputs[4193]) | (layer0_outputs[12588]);
    assign layer1_outputs[3421] = layer0_outputs[604];
    assign layer1_outputs[3422] = ~(layer0_outputs[4245]);
    assign layer1_outputs[3423] = ~((layer0_outputs[12527]) & (layer0_outputs[1571]));
    assign layer1_outputs[3424] = ~(layer0_outputs[8137]) | (layer0_outputs[11909]);
    assign layer1_outputs[3425] = ~(layer0_outputs[2532]);
    assign layer1_outputs[3426] = ~((layer0_outputs[9255]) ^ (layer0_outputs[9762]));
    assign layer1_outputs[3427] = (layer0_outputs[130]) ^ (layer0_outputs[6419]);
    assign layer1_outputs[3428] = ~(layer0_outputs[11150]) | (layer0_outputs[8547]);
    assign layer1_outputs[3429] = layer0_outputs[11574];
    assign layer1_outputs[3430] = layer0_outputs[1258];
    assign layer1_outputs[3431] = ~(layer0_outputs[656]) | (layer0_outputs[11199]);
    assign layer1_outputs[3432] = layer0_outputs[1531];
    assign layer1_outputs[3433] = ~((layer0_outputs[833]) & (layer0_outputs[5028]));
    assign layer1_outputs[3434] = (layer0_outputs[6593]) & (layer0_outputs[5796]);
    assign layer1_outputs[3435] = ~((layer0_outputs[10006]) & (layer0_outputs[2168]));
    assign layer1_outputs[3436] = ~(layer0_outputs[7929]);
    assign layer1_outputs[3437] = ~((layer0_outputs[11975]) ^ (layer0_outputs[6437]));
    assign layer1_outputs[3438] = (layer0_outputs[2010]) & (layer0_outputs[5633]);
    assign layer1_outputs[3439] = layer0_outputs[8458];
    assign layer1_outputs[3440] = (layer0_outputs[6128]) & (layer0_outputs[2832]);
    assign layer1_outputs[3441] = 1'b1;
    assign layer1_outputs[3442] = ~(layer0_outputs[12053]);
    assign layer1_outputs[3443] = ~(layer0_outputs[6652]) | (layer0_outputs[7306]);
    assign layer1_outputs[3444] = ~(layer0_outputs[1679]);
    assign layer1_outputs[3445] = ~(layer0_outputs[7626]);
    assign layer1_outputs[3446] = (layer0_outputs[4020]) | (layer0_outputs[285]);
    assign layer1_outputs[3447] = (layer0_outputs[11609]) & (layer0_outputs[10722]);
    assign layer1_outputs[3448] = ~(layer0_outputs[8854]);
    assign layer1_outputs[3449] = (layer0_outputs[2308]) & ~(layer0_outputs[6539]);
    assign layer1_outputs[3450] = layer0_outputs[3765];
    assign layer1_outputs[3451] = (layer0_outputs[1290]) & ~(layer0_outputs[1618]);
    assign layer1_outputs[3452] = ~(layer0_outputs[984]) | (layer0_outputs[8073]);
    assign layer1_outputs[3453] = layer0_outputs[918];
    assign layer1_outputs[3454] = ~((layer0_outputs[275]) | (layer0_outputs[6290]));
    assign layer1_outputs[3455] = ~(layer0_outputs[9153]);
    assign layer1_outputs[3456] = layer0_outputs[9740];
    assign layer1_outputs[3457] = 1'b0;
    assign layer1_outputs[3458] = ~(layer0_outputs[6803]);
    assign layer1_outputs[3459] = (layer0_outputs[9827]) & (layer0_outputs[4242]);
    assign layer1_outputs[3460] = ~(layer0_outputs[1679]);
    assign layer1_outputs[3461] = ~((layer0_outputs[9154]) | (layer0_outputs[5627]));
    assign layer1_outputs[3462] = ~((layer0_outputs[1483]) ^ (layer0_outputs[2799]));
    assign layer1_outputs[3463] = ~(layer0_outputs[5950]);
    assign layer1_outputs[3464] = ~((layer0_outputs[4969]) & (layer0_outputs[8380]));
    assign layer1_outputs[3465] = layer0_outputs[6673];
    assign layer1_outputs[3466] = layer0_outputs[9654];
    assign layer1_outputs[3467] = (layer0_outputs[7462]) & ~(layer0_outputs[6282]);
    assign layer1_outputs[3468] = ~(layer0_outputs[4539]);
    assign layer1_outputs[3469] = (layer0_outputs[8392]) | (layer0_outputs[3915]);
    assign layer1_outputs[3470] = ~(layer0_outputs[9749]);
    assign layer1_outputs[3471] = ~((layer0_outputs[2922]) ^ (layer0_outputs[1562]));
    assign layer1_outputs[3472] = layer0_outputs[12122];
    assign layer1_outputs[3473] = (layer0_outputs[2023]) & ~(layer0_outputs[5147]);
    assign layer1_outputs[3474] = layer0_outputs[2319];
    assign layer1_outputs[3475] = (layer0_outputs[2661]) | (layer0_outputs[8745]);
    assign layer1_outputs[3476] = (layer0_outputs[480]) & ~(layer0_outputs[3246]);
    assign layer1_outputs[3477] = (layer0_outputs[10089]) & ~(layer0_outputs[3767]);
    assign layer1_outputs[3478] = ~(layer0_outputs[2074]) | (layer0_outputs[10969]);
    assign layer1_outputs[3479] = ~(layer0_outputs[2404]);
    assign layer1_outputs[3480] = ~((layer0_outputs[10580]) | (layer0_outputs[12709]));
    assign layer1_outputs[3481] = (layer0_outputs[9586]) & ~(layer0_outputs[6037]);
    assign layer1_outputs[3482] = ~((layer0_outputs[3372]) | (layer0_outputs[4607]));
    assign layer1_outputs[3483] = layer0_outputs[8742];
    assign layer1_outputs[3484] = ~(layer0_outputs[1218]);
    assign layer1_outputs[3485] = (layer0_outputs[9270]) & ~(layer0_outputs[2839]);
    assign layer1_outputs[3486] = (layer0_outputs[3670]) & ~(layer0_outputs[2818]);
    assign layer1_outputs[3487] = layer0_outputs[4848];
    assign layer1_outputs[3488] = (layer0_outputs[10754]) & ~(layer0_outputs[9256]);
    assign layer1_outputs[3489] = ~((layer0_outputs[3069]) & (layer0_outputs[6478]));
    assign layer1_outputs[3490] = 1'b1;
    assign layer1_outputs[3491] = ~(layer0_outputs[9250]) | (layer0_outputs[6761]);
    assign layer1_outputs[3492] = ~(layer0_outputs[2919]);
    assign layer1_outputs[3493] = ~(layer0_outputs[6314]) | (layer0_outputs[463]);
    assign layer1_outputs[3494] = (layer0_outputs[12776]) ^ (layer0_outputs[1004]);
    assign layer1_outputs[3495] = layer0_outputs[4277];
    assign layer1_outputs[3496] = (layer0_outputs[8518]) ^ (layer0_outputs[9221]);
    assign layer1_outputs[3497] = (layer0_outputs[3026]) & ~(layer0_outputs[4803]);
    assign layer1_outputs[3498] = ~((layer0_outputs[11802]) ^ (layer0_outputs[11861]));
    assign layer1_outputs[3499] = (layer0_outputs[5947]) & ~(layer0_outputs[8384]);
    assign layer1_outputs[3500] = ~((layer0_outputs[8376]) & (layer0_outputs[8004]));
    assign layer1_outputs[3501] = ~((layer0_outputs[4511]) | (layer0_outputs[1184]));
    assign layer1_outputs[3502] = layer0_outputs[10252];
    assign layer1_outputs[3503] = (layer0_outputs[12277]) | (layer0_outputs[3146]);
    assign layer1_outputs[3504] = (layer0_outputs[4615]) & ~(layer0_outputs[10921]);
    assign layer1_outputs[3505] = layer0_outputs[2251];
    assign layer1_outputs[3506] = 1'b1;
    assign layer1_outputs[3507] = (layer0_outputs[4986]) & (layer0_outputs[763]);
    assign layer1_outputs[3508] = (layer0_outputs[3114]) & (layer0_outputs[1546]);
    assign layer1_outputs[3509] = (layer0_outputs[12711]) ^ (layer0_outputs[11532]);
    assign layer1_outputs[3510] = ~(layer0_outputs[7489]) | (layer0_outputs[10433]);
    assign layer1_outputs[3511] = (layer0_outputs[6187]) & ~(layer0_outputs[76]);
    assign layer1_outputs[3512] = (layer0_outputs[4027]) | (layer0_outputs[10195]);
    assign layer1_outputs[3513] = (layer0_outputs[3860]) & (layer0_outputs[8629]);
    assign layer1_outputs[3514] = layer0_outputs[1661];
    assign layer1_outputs[3515] = (layer0_outputs[3601]) & ~(layer0_outputs[867]);
    assign layer1_outputs[3516] = (layer0_outputs[9954]) | (layer0_outputs[5842]);
    assign layer1_outputs[3517] = 1'b0;
    assign layer1_outputs[3518] = 1'b0;
    assign layer1_outputs[3519] = ~((layer0_outputs[2371]) | (layer0_outputs[1439]));
    assign layer1_outputs[3520] = (layer0_outputs[2242]) ^ (layer0_outputs[4508]);
    assign layer1_outputs[3521] = ~((layer0_outputs[5293]) | (layer0_outputs[4238]));
    assign layer1_outputs[3522] = (layer0_outputs[10015]) ^ (layer0_outputs[8587]);
    assign layer1_outputs[3523] = ~(layer0_outputs[4364]) | (layer0_outputs[2130]);
    assign layer1_outputs[3524] = layer0_outputs[7139];
    assign layer1_outputs[3525] = (layer0_outputs[5406]) & (layer0_outputs[1268]);
    assign layer1_outputs[3526] = ~(layer0_outputs[810]);
    assign layer1_outputs[3527] = layer0_outputs[12711];
    assign layer1_outputs[3528] = (layer0_outputs[3683]) & ~(layer0_outputs[7808]);
    assign layer1_outputs[3529] = layer0_outputs[6959];
    assign layer1_outputs[3530] = ~(layer0_outputs[11027]) | (layer0_outputs[10177]);
    assign layer1_outputs[3531] = ~(layer0_outputs[10362]);
    assign layer1_outputs[3532] = ~(layer0_outputs[5121]) | (layer0_outputs[9994]);
    assign layer1_outputs[3533] = 1'b1;
    assign layer1_outputs[3534] = ~(layer0_outputs[4993]);
    assign layer1_outputs[3535] = 1'b0;
    assign layer1_outputs[3536] = 1'b1;
    assign layer1_outputs[3537] = ~((layer0_outputs[2268]) & (layer0_outputs[10681]));
    assign layer1_outputs[3538] = layer0_outputs[10404];
    assign layer1_outputs[3539] = (layer0_outputs[12019]) ^ (layer0_outputs[766]);
    assign layer1_outputs[3540] = ~((layer0_outputs[1222]) ^ (layer0_outputs[7493]));
    assign layer1_outputs[3541] = (layer0_outputs[11393]) & (layer0_outputs[4505]);
    assign layer1_outputs[3542] = ~((layer0_outputs[1797]) ^ (layer0_outputs[12318]));
    assign layer1_outputs[3543] = layer0_outputs[3245];
    assign layer1_outputs[3544] = ~(layer0_outputs[12648]) | (layer0_outputs[5646]);
    assign layer1_outputs[3545] = layer0_outputs[3659];
    assign layer1_outputs[3546] = ~((layer0_outputs[1193]) ^ (layer0_outputs[316]));
    assign layer1_outputs[3547] = (layer0_outputs[11322]) & (layer0_outputs[516]);
    assign layer1_outputs[3548] = ~((layer0_outputs[7936]) ^ (layer0_outputs[2845]));
    assign layer1_outputs[3549] = ~((layer0_outputs[11088]) & (layer0_outputs[10395]));
    assign layer1_outputs[3550] = ~(layer0_outputs[3825]);
    assign layer1_outputs[3551] = ~(layer0_outputs[6730]);
    assign layer1_outputs[3552] = ~(layer0_outputs[7231]);
    assign layer1_outputs[3553] = layer0_outputs[3674];
    assign layer1_outputs[3554] = (layer0_outputs[9583]) | (layer0_outputs[10598]);
    assign layer1_outputs[3555] = 1'b0;
    assign layer1_outputs[3556] = layer0_outputs[11593];
    assign layer1_outputs[3557] = (layer0_outputs[4240]) | (layer0_outputs[1109]);
    assign layer1_outputs[3558] = (layer0_outputs[3442]) & (layer0_outputs[4513]);
    assign layer1_outputs[3559] = ~(layer0_outputs[5260]) | (layer0_outputs[2305]);
    assign layer1_outputs[3560] = ~((layer0_outputs[6367]) ^ (layer0_outputs[3041]));
    assign layer1_outputs[3561] = (layer0_outputs[3577]) | (layer0_outputs[1518]);
    assign layer1_outputs[3562] = (layer0_outputs[5771]) & (layer0_outputs[8580]);
    assign layer1_outputs[3563] = layer0_outputs[1808];
    assign layer1_outputs[3564] = ~(layer0_outputs[18]);
    assign layer1_outputs[3565] = ~(layer0_outputs[11605]);
    assign layer1_outputs[3566] = 1'b1;
    assign layer1_outputs[3567] = ~(layer0_outputs[2152]);
    assign layer1_outputs[3568] = ~((layer0_outputs[1844]) | (layer0_outputs[6747]));
    assign layer1_outputs[3569] = (layer0_outputs[566]) ^ (layer0_outputs[8024]);
    assign layer1_outputs[3570] = layer0_outputs[6782];
    assign layer1_outputs[3571] = layer0_outputs[2500];
    assign layer1_outputs[3572] = layer0_outputs[1530];
    assign layer1_outputs[3573] = ~(layer0_outputs[7683]);
    assign layer1_outputs[3574] = (layer0_outputs[1115]) ^ (layer0_outputs[2599]);
    assign layer1_outputs[3575] = (layer0_outputs[7897]) & ~(layer0_outputs[11195]);
    assign layer1_outputs[3576] = ~(layer0_outputs[8375]) | (layer0_outputs[11676]);
    assign layer1_outputs[3577] = (layer0_outputs[7993]) | (layer0_outputs[99]);
    assign layer1_outputs[3578] = layer0_outputs[5911];
    assign layer1_outputs[3579] = layer0_outputs[9618];
    assign layer1_outputs[3580] = (layer0_outputs[7123]) & ~(layer0_outputs[1100]);
    assign layer1_outputs[3581] = (layer0_outputs[10356]) | (layer0_outputs[8467]);
    assign layer1_outputs[3582] = (layer0_outputs[2050]) & (layer0_outputs[2218]);
    assign layer1_outputs[3583] = 1'b0;
    assign layer1_outputs[3584] = layer0_outputs[9455];
    assign layer1_outputs[3585] = (layer0_outputs[8308]) ^ (layer0_outputs[2773]);
    assign layer1_outputs[3586] = ~((layer0_outputs[11277]) ^ (layer0_outputs[894]));
    assign layer1_outputs[3587] = ~(layer0_outputs[12429]);
    assign layer1_outputs[3588] = ~(layer0_outputs[6709]) | (layer0_outputs[8585]);
    assign layer1_outputs[3589] = ~(layer0_outputs[10527]);
    assign layer1_outputs[3590] = layer0_outputs[9595];
    assign layer1_outputs[3591] = ~(layer0_outputs[8888]) | (layer0_outputs[4706]);
    assign layer1_outputs[3592] = (layer0_outputs[2112]) & (layer0_outputs[8537]);
    assign layer1_outputs[3593] = layer0_outputs[10104];
    assign layer1_outputs[3594] = (layer0_outputs[4322]) & (layer0_outputs[7440]);
    assign layer1_outputs[3595] = (layer0_outputs[3000]) ^ (layer0_outputs[11937]);
    assign layer1_outputs[3596] = ~(layer0_outputs[1775]) | (layer0_outputs[11750]);
    assign layer1_outputs[3597] = ~((layer0_outputs[12794]) ^ (layer0_outputs[7630]));
    assign layer1_outputs[3598] = (layer0_outputs[6288]) | (layer0_outputs[11848]);
    assign layer1_outputs[3599] = (layer0_outputs[7105]) & (layer0_outputs[945]);
    assign layer1_outputs[3600] = (layer0_outputs[12468]) & (layer0_outputs[6303]);
    assign layer1_outputs[3601] = ~(layer0_outputs[830]);
    assign layer1_outputs[3602] = ~((layer0_outputs[12054]) & (layer0_outputs[8468]));
    assign layer1_outputs[3603] = (layer0_outputs[4067]) | (layer0_outputs[11237]);
    assign layer1_outputs[3604] = ~(layer0_outputs[4560]) | (layer0_outputs[9553]);
    assign layer1_outputs[3605] = 1'b0;
    assign layer1_outputs[3606] = layer0_outputs[8215];
    assign layer1_outputs[3607] = layer0_outputs[11637];
    assign layer1_outputs[3608] = (layer0_outputs[2891]) ^ (layer0_outputs[10396]);
    assign layer1_outputs[3609] = ~((layer0_outputs[6239]) ^ (layer0_outputs[6053]));
    assign layer1_outputs[3610] = ~(layer0_outputs[5382]) | (layer0_outputs[3811]);
    assign layer1_outputs[3611] = ~(layer0_outputs[1078]) | (layer0_outputs[7970]);
    assign layer1_outputs[3612] = layer0_outputs[10788];
    assign layer1_outputs[3613] = ~((layer0_outputs[6337]) & (layer0_outputs[7917]));
    assign layer1_outputs[3614] = layer0_outputs[8550];
    assign layer1_outputs[3615] = ~((layer0_outputs[10956]) ^ (layer0_outputs[9570]));
    assign layer1_outputs[3616] = layer0_outputs[10890];
    assign layer1_outputs[3617] = layer0_outputs[8144];
    assign layer1_outputs[3618] = (layer0_outputs[3230]) | (layer0_outputs[9756]);
    assign layer1_outputs[3619] = ~(layer0_outputs[9495]) | (layer0_outputs[7188]);
    assign layer1_outputs[3620] = 1'b1;
    assign layer1_outputs[3621] = layer0_outputs[4425];
    assign layer1_outputs[3622] = (layer0_outputs[1145]) | (layer0_outputs[1111]);
    assign layer1_outputs[3623] = ~((layer0_outputs[5924]) & (layer0_outputs[2707]));
    assign layer1_outputs[3624] = layer0_outputs[5923];
    assign layer1_outputs[3625] = (layer0_outputs[4904]) & ~(layer0_outputs[337]);
    assign layer1_outputs[3626] = (layer0_outputs[4695]) & ~(layer0_outputs[10990]);
    assign layer1_outputs[3627] = ~(layer0_outputs[2651]);
    assign layer1_outputs[3628] = layer0_outputs[7073];
    assign layer1_outputs[3629] = ~(layer0_outputs[10747]);
    assign layer1_outputs[3630] = layer0_outputs[4121];
    assign layer1_outputs[3631] = (layer0_outputs[2344]) | (layer0_outputs[3085]);
    assign layer1_outputs[3632] = ~(layer0_outputs[9278]);
    assign layer1_outputs[3633] = (layer0_outputs[6676]) ^ (layer0_outputs[5498]);
    assign layer1_outputs[3634] = layer0_outputs[8638];
    assign layer1_outputs[3635] = ~((layer0_outputs[4393]) & (layer0_outputs[10035]));
    assign layer1_outputs[3636] = ~(layer0_outputs[10323]);
    assign layer1_outputs[3637] = 1'b1;
    assign layer1_outputs[3638] = layer0_outputs[10901];
    assign layer1_outputs[3639] = 1'b0;
    assign layer1_outputs[3640] = ~(layer0_outputs[551]) | (layer0_outputs[5132]);
    assign layer1_outputs[3641] = ~(layer0_outputs[6343]);
    assign layer1_outputs[3642] = (layer0_outputs[7134]) & (layer0_outputs[1698]);
    assign layer1_outputs[3643] = ~((layer0_outputs[3802]) & (layer0_outputs[10531]));
    assign layer1_outputs[3644] = ~(layer0_outputs[7941]) | (layer0_outputs[9937]);
    assign layer1_outputs[3645] = (layer0_outputs[6496]) | (layer0_outputs[2598]);
    assign layer1_outputs[3646] = ~((layer0_outputs[7668]) ^ (layer0_outputs[4434]));
    assign layer1_outputs[3647] = ~(layer0_outputs[11701]);
    assign layer1_outputs[3648] = ~((layer0_outputs[12658]) ^ (layer0_outputs[10039]));
    assign layer1_outputs[3649] = ~((layer0_outputs[2665]) | (layer0_outputs[5865]));
    assign layer1_outputs[3650] = layer0_outputs[4934];
    assign layer1_outputs[3651] = ~((layer0_outputs[4465]) & (layer0_outputs[10309]));
    assign layer1_outputs[3652] = ~(layer0_outputs[10710]);
    assign layer1_outputs[3653] = ~((layer0_outputs[12790]) ^ (layer0_outputs[11858]));
    assign layer1_outputs[3654] = (layer0_outputs[12570]) | (layer0_outputs[4132]);
    assign layer1_outputs[3655] = (layer0_outputs[2657]) ^ (layer0_outputs[6050]);
    assign layer1_outputs[3656] = ~(layer0_outputs[6845]);
    assign layer1_outputs[3657] = (layer0_outputs[5369]) ^ (layer0_outputs[831]);
    assign layer1_outputs[3658] = (layer0_outputs[9835]) ^ (layer0_outputs[4938]);
    assign layer1_outputs[3659] = layer0_outputs[63];
    assign layer1_outputs[3660] = 1'b0;
    assign layer1_outputs[3661] = (layer0_outputs[2067]) & ~(layer0_outputs[10605]);
    assign layer1_outputs[3662] = ~(layer0_outputs[6040]) | (layer0_outputs[12515]);
    assign layer1_outputs[3663] = ~(layer0_outputs[7558]) | (layer0_outputs[6142]);
    assign layer1_outputs[3664] = layer0_outputs[5658];
    assign layer1_outputs[3665] = ~(layer0_outputs[3748]) | (layer0_outputs[12503]);
    assign layer1_outputs[3666] = ~((layer0_outputs[393]) & (layer0_outputs[9199]));
    assign layer1_outputs[3667] = layer0_outputs[2503];
    assign layer1_outputs[3668] = ~((layer0_outputs[9110]) & (layer0_outputs[8452]));
    assign layer1_outputs[3669] = layer0_outputs[868];
    assign layer1_outputs[3670] = layer0_outputs[11687];
    assign layer1_outputs[3671] = ~(layer0_outputs[4664]) | (layer0_outputs[5023]);
    assign layer1_outputs[3672] = ~(layer0_outputs[6500]) | (layer0_outputs[12017]);
    assign layer1_outputs[3673] = layer0_outputs[2362];
    assign layer1_outputs[3674] = ~(layer0_outputs[9855]) | (layer0_outputs[7805]);
    assign layer1_outputs[3675] = ~((layer0_outputs[5096]) | (layer0_outputs[1161]));
    assign layer1_outputs[3676] = layer0_outputs[822];
    assign layer1_outputs[3677] = ~(layer0_outputs[11649]);
    assign layer1_outputs[3678] = ~(layer0_outputs[5950]);
    assign layer1_outputs[3679] = ~((layer0_outputs[11600]) | (layer0_outputs[10844]));
    assign layer1_outputs[3680] = ~((layer0_outputs[5989]) & (layer0_outputs[12624]));
    assign layer1_outputs[3681] = layer0_outputs[7145];
    assign layer1_outputs[3682] = ~((layer0_outputs[6940]) & (layer0_outputs[547]));
    assign layer1_outputs[3683] = ~(layer0_outputs[2297]) | (layer0_outputs[11435]);
    assign layer1_outputs[3684] = (layer0_outputs[3087]) | (layer0_outputs[3342]);
    assign layer1_outputs[3685] = ~(layer0_outputs[11829]);
    assign layer1_outputs[3686] = ~(layer0_outputs[8379]);
    assign layer1_outputs[3687] = ~(layer0_outputs[1424]) | (layer0_outputs[4631]);
    assign layer1_outputs[3688] = (layer0_outputs[7132]) ^ (layer0_outputs[5033]);
    assign layer1_outputs[3689] = ~(layer0_outputs[4231]) | (layer0_outputs[5188]);
    assign layer1_outputs[3690] = (layer0_outputs[1915]) | (layer0_outputs[10770]);
    assign layer1_outputs[3691] = (layer0_outputs[3750]) & (layer0_outputs[5505]);
    assign layer1_outputs[3692] = ~(layer0_outputs[10740]) | (layer0_outputs[8853]);
    assign layer1_outputs[3693] = layer0_outputs[11959];
    assign layer1_outputs[3694] = ~((layer0_outputs[7976]) ^ (layer0_outputs[3165]));
    assign layer1_outputs[3695] = layer0_outputs[8010];
    assign layer1_outputs[3696] = ~(layer0_outputs[213]);
    assign layer1_outputs[3697] = ~(layer0_outputs[12005]);
    assign layer1_outputs[3698] = layer0_outputs[2433];
    assign layer1_outputs[3699] = ~(layer0_outputs[1713]);
    assign layer1_outputs[3700] = ~(layer0_outputs[7980]) | (layer0_outputs[3862]);
    assign layer1_outputs[3701] = layer0_outputs[926];
    assign layer1_outputs[3702] = 1'b0;
    assign layer1_outputs[3703] = ~((layer0_outputs[5079]) ^ (layer0_outputs[1223]));
    assign layer1_outputs[3704] = (layer0_outputs[2638]) & (layer0_outputs[8227]);
    assign layer1_outputs[3705] = layer0_outputs[1255];
    assign layer1_outputs[3706] = layer0_outputs[8601];
    assign layer1_outputs[3707] = (layer0_outputs[7086]) & ~(layer0_outputs[792]);
    assign layer1_outputs[3708] = layer0_outputs[10706];
    assign layer1_outputs[3709] = ~(layer0_outputs[908]);
    assign layer1_outputs[3710] = layer0_outputs[7886];
    assign layer1_outputs[3711] = ~(layer0_outputs[11895]);
    assign layer1_outputs[3712] = layer0_outputs[12545];
    assign layer1_outputs[3713] = (layer0_outputs[384]) | (layer0_outputs[8340]);
    assign layer1_outputs[3714] = ~(layer0_outputs[7727]);
    assign layer1_outputs[3715] = (layer0_outputs[3234]) | (layer0_outputs[10755]);
    assign layer1_outputs[3716] = layer0_outputs[6286];
    assign layer1_outputs[3717] = ~(layer0_outputs[3559]);
    assign layer1_outputs[3718] = ~((layer0_outputs[6986]) & (layer0_outputs[5949]));
    assign layer1_outputs[3719] = (layer0_outputs[1452]) ^ (layer0_outputs[11792]);
    assign layer1_outputs[3720] = ~(layer0_outputs[4031]) | (layer0_outputs[11001]);
    assign layer1_outputs[3721] = (layer0_outputs[8003]) ^ (layer0_outputs[3157]);
    assign layer1_outputs[3722] = (layer0_outputs[12771]) & (layer0_outputs[10293]);
    assign layer1_outputs[3723] = ~((layer0_outputs[4160]) ^ (layer0_outputs[8462]));
    assign layer1_outputs[3724] = (layer0_outputs[754]) ^ (layer0_outputs[8326]);
    assign layer1_outputs[3725] = ~((layer0_outputs[11571]) | (layer0_outputs[10746]));
    assign layer1_outputs[3726] = ~(layer0_outputs[11580]);
    assign layer1_outputs[3727] = (layer0_outputs[7830]) ^ (layer0_outputs[1456]);
    assign layer1_outputs[3728] = (layer0_outputs[7591]) & ~(layer0_outputs[5447]);
    assign layer1_outputs[3729] = layer0_outputs[10299];
    assign layer1_outputs[3730] = layer0_outputs[7403];
    assign layer1_outputs[3731] = 1'b0;
    assign layer1_outputs[3732] = ~(layer0_outputs[3685]);
    assign layer1_outputs[3733] = 1'b0;
    assign layer1_outputs[3734] = ~(layer0_outputs[47]);
    assign layer1_outputs[3735] = ~((layer0_outputs[4358]) ^ (layer0_outputs[11404]));
    assign layer1_outputs[3736] = (layer0_outputs[1773]) | (layer0_outputs[2813]);
    assign layer1_outputs[3737] = ~(layer0_outputs[6789]);
    assign layer1_outputs[3738] = ~(layer0_outputs[1247]);
    assign layer1_outputs[3739] = (layer0_outputs[11029]) & ~(layer0_outputs[12381]);
    assign layer1_outputs[3740] = ~((layer0_outputs[2325]) & (layer0_outputs[8486]));
    assign layer1_outputs[3741] = (layer0_outputs[10717]) ^ (layer0_outputs[8794]);
    assign layer1_outputs[3742] = (layer0_outputs[12362]) & (layer0_outputs[1909]);
    assign layer1_outputs[3743] = ~(layer0_outputs[1726]) | (layer0_outputs[2133]);
    assign layer1_outputs[3744] = 1'b0;
    assign layer1_outputs[3745] = layer0_outputs[6757];
    assign layer1_outputs[3746] = layer0_outputs[2211];
    assign layer1_outputs[3747] = (layer0_outputs[11649]) ^ (layer0_outputs[3454]);
    assign layer1_outputs[3748] = ~((layer0_outputs[10654]) | (layer0_outputs[6137]));
    assign layer1_outputs[3749] = ~((layer0_outputs[253]) ^ (layer0_outputs[2798]));
    assign layer1_outputs[3750] = (layer0_outputs[6256]) ^ (layer0_outputs[11863]);
    assign layer1_outputs[3751] = (layer0_outputs[7718]) | (layer0_outputs[1021]);
    assign layer1_outputs[3752] = ~(layer0_outputs[7526]);
    assign layer1_outputs[3753] = ~((layer0_outputs[4753]) ^ (layer0_outputs[3210]));
    assign layer1_outputs[3754] = ~((layer0_outputs[2273]) ^ (layer0_outputs[6632]));
    assign layer1_outputs[3755] = (layer0_outputs[8510]) & ~(layer0_outputs[2688]);
    assign layer1_outputs[3756] = layer0_outputs[6304];
    assign layer1_outputs[3757] = ~(layer0_outputs[7598]);
    assign layer1_outputs[3758] = ~((layer0_outputs[4624]) | (layer0_outputs[7708]));
    assign layer1_outputs[3759] = ~(layer0_outputs[3214]);
    assign layer1_outputs[3760] = 1'b0;
    assign layer1_outputs[3761] = ~((layer0_outputs[1981]) ^ (layer0_outputs[10973]));
    assign layer1_outputs[3762] = layer0_outputs[11539];
    assign layer1_outputs[3763] = layer0_outputs[10112];
    assign layer1_outputs[3764] = (layer0_outputs[6391]) & ~(layer0_outputs[11451]);
    assign layer1_outputs[3765] = ~(layer0_outputs[6357]);
    assign layer1_outputs[3766] = ~(layer0_outputs[11845]);
    assign layer1_outputs[3767] = ~((layer0_outputs[2543]) | (layer0_outputs[11870]));
    assign layer1_outputs[3768] = (layer0_outputs[3887]) & ~(layer0_outputs[4835]);
    assign layer1_outputs[3769] = ~(layer0_outputs[2008]) | (layer0_outputs[11904]);
    assign layer1_outputs[3770] = (layer0_outputs[10442]) & ~(layer0_outputs[3760]);
    assign layer1_outputs[3771] = (layer0_outputs[2506]) & (layer0_outputs[8004]);
    assign layer1_outputs[3772] = (layer0_outputs[11962]) & ~(layer0_outputs[5829]);
    assign layer1_outputs[3773] = (layer0_outputs[6958]) | (layer0_outputs[11459]);
    assign layer1_outputs[3774] = (layer0_outputs[94]) ^ (layer0_outputs[992]);
    assign layer1_outputs[3775] = (layer0_outputs[3979]) ^ (layer0_outputs[1980]);
    assign layer1_outputs[3776] = ~(layer0_outputs[11141]) | (layer0_outputs[601]);
    assign layer1_outputs[3777] = layer0_outputs[7844];
    assign layer1_outputs[3778] = (layer0_outputs[2]) & ~(layer0_outputs[5379]);
    assign layer1_outputs[3779] = ~((layer0_outputs[9643]) ^ (layer0_outputs[6027]));
    assign layer1_outputs[3780] = ~(layer0_outputs[11111]);
    assign layer1_outputs[3781] = ~(layer0_outputs[10656]);
    assign layer1_outputs[3782] = ~(layer0_outputs[3173]);
    assign layer1_outputs[3783] = ~(layer0_outputs[2856]);
    assign layer1_outputs[3784] = ~(layer0_outputs[5605]);
    assign layer1_outputs[3785] = ~(layer0_outputs[4535]);
    assign layer1_outputs[3786] = ~((layer0_outputs[9253]) ^ (layer0_outputs[387]));
    assign layer1_outputs[3787] = ~(layer0_outputs[10674]) | (layer0_outputs[1891]);
    assign layer1_outputs[3788] = layer0_outputs[5257];
    assign layer1_outputs[3789] = ~(layer0_outputs[6740]);
    assign layer1_outputs[3790] = layer0_outputs[6399];
    assign layer1_outputs[3791] = (layer0_outputs[6188]) | (layer0_outputs[2918]);
    assign layer1_outputs[3792] = ~(layer0_outputs[1038]);
    assign layer1_outputs[3793] = layer0_outputs[10791];
    assign layer1_outputs[3794] = ~(layer0_outputs[749]) | (layer0_outputs[7916]);
    assign layer1_outputs[3795] = layer0_outputs[8584];
    assign layer1_outputs[3796] = (layer0_outputs[9744]) | (layer0_outputs[7409]);
    assign layer1_outputs[3797] = ~((layer0_outputs[1080]) & (layer0_outputs[3463]));
    assign layer1_outputs[3798] = 1'b0;
    assign layer1_outputs[3799] = (layer0_outputs[4800]) & (layer0_outputs[11963]);
    assign layer1_outputs[3800] = layer0_outputs[11737];
    assign layer1_outputs[3801] = ~(layer0_outputs[6444]);
    assign layer1_outputs[3802] = (layer0_outputs[519]) & ~(layer0_outputs[1418]);
    assign layer1_outputs[3803] = layer0_outputs[4322];
    assign layer1_outputs[3804] = 1'b0;
    assign layer1_outputs[3805] = (layer0_outputs[3155]) & ~(layer0_outputs[4049]);
    assign layer1_outputs[3806] = layer0_outputs[4918];
    assign layer1_outputs[3807] = ~((layer0_outputs[1001]) ^ (layer0_outputs[2384]));
    assign layer1_outputs[3808] = layer0_outputs[1815];
    assign layer1_outputs[3809] = ~(layer0_outputs[3723]);
    assign layer1_outputs[3810] = ~((layer0_outputs[9546]) & (layer0_outputs[1774]));
    assign layer1_outputs[3811] = layer0_outputs[6638];
    assign layer1_outputs[3812] = (layer0_outputs[7828]) | (layer0_outputs[10463]);
    assign layer1_outputs[3813] = (layer0_outputs[4640]) & ~(layer0_outputs[5404]);
    assign layer1_outputs[3814] = layer0_outputs[9703];
    assign layer1_outputs[3815] = ~((layer0_outputs[2948]) & (layer0_outputs[1682]));
    assign layer1_outputs[3816] = (layer0_outputs[7532]) & (layer0_outputs[5520]);
    assign layer1_outputs[3817] = layer0_outputs[9545];
    assign layer1_outputs[3818] = ~(layer0_outputs[12316]);
    assign layer1_outputs[3819] = ~(layer0_outputs[12012]);
    assign layer1_outputs[3820] = ~((layer0_outputs[3347]) | (layer0_outputs[11028]));
    assign layer1_outputs[3821] = layer0_outputs[10045];
    assign layer1_outputs[3822] = ~(layer0_outputs[7809]) | (layer0_outputs[7344]);
    assign layer1_outputs[3823] = layer0_outputs[9302];
    assign layer1_outputs[3824] = layer0_outputs[362];
    assign layer1_outputs[3825] = ~((layer0_outputs[7281]) | (layer0_outputs[9719]));
    assign layer1_outputs[3826] = (layer0_outputs[300]) ^ (layer0_outputs[9707]);
    assign layer1_outputs[3827] = ~((layer0_outputs[2089]) ^ (layer0_outputs[11912]));
    assign layer1_outputs[3828] = ~((layer0_outputs[7049]) & (layer0_outputs[860]));
    assign layer1_outputs[3829] = (layer0_outputs[11334]) ^ (layer0_outputs[3478]);
    assign layer1_outputs[3830] = ~(layer0_outputs[7149]);
    assign layer1_outputs[3831] = ~((layer0_outputs[10545]) ^ (layer0_outputs[9033]));
    assign layer1_outputs[3832] = ~(layer0_outputs[4747]) | (layer0_outputs[7540]);
    assign layer1_outputs[3833] = ~(layer0_outputs[1529]);
    assign layer1_outputs[3834] = ~((layer0_outputs[8157]) & (layer0_outputs[10120]));
    assign layer1_outputs[3835] = layer0_outputs[10246];
    assign layer1_outputs[3836] = (layer0_outputs[12693]) & ~(layer0_outputs[1525]);
    assign layer1_outputs[3837] = layer0_outputs[9730];
    assign layer1_outputs[3838] = ~((layer0_outputs[266]) & (layer0_outputs[8746]));
    assign layer1_outputs[3839] = ~(layer0_outputs[1318]);
    assign layer1_outputs[3840] = (layer0_outputs[11101]) | (layer0_outputs[12226]);
    assign layer1_outputs[3841] = ~(layer0_outputs[12265]) | (layer0_outputs[9859]);
    assign layer1_outputs[3842] = (layer0_outputs[3044]) & ~(layer0_outputs[2870]);
    assign layer1_outputs[3843] = layer0_outputs[826];
    assign layer1_outputs[3844] = (layer0_outputs[10960]) & ~(layer0_outputs[2171]);
    assign layer1_outputs[3845] = ~(layer0_outputs[5712]);
    assign layer1_outputs[3846] = ~((layer0_outputs[6420]) & (layer0_outputs[10021]));
    assign layer1_outputs[3847] = layer0_outputs[6982];
    assign layer1_outputs[3848] = (layer0_outputs[6971]) & (layer0_outputs[12431]);
    assign layer1_outputs[3849] = layer0_outputs[6607];
    assign layer1_outputs[3850] = (layer0_outputs[4653]) & ~(layer0_outputs[11146]);
    assign layer1_outputs[3851] = (layer0_outputs[2494]) & (layer0_outputs[4040]);
    assign layer1_outputs[3852] = (layer0_outputs[11506]) & (layer0_outputs[4942]);
    assign layer1_outputs[3853] = ~(layer0_outputs[5445]) | (layer0_outputs[12663]);
    assign layer1_outputs[3854] = (layer0_outputs[642]) & ~(layer0_outputs[10875]);
    assign layer1_outputs[3855] = (layer0_outputs[9049]) | (layer0_outputs[6702]);
    assign layer1_outputs[3856] = layer0_outputs[3481];
    assign layer1_outputs[3857] = (layer0_outputs[449]) ^ (layer0_outputs[4767]);
    assign layer1_outputs[3858] = ~(layer0_outputs[10765]);
    assign layer1_outputs[3859] = (layer0_outputs[8212]) ^ (layer0_outputs[1262]);
    assign layer1_outputs[3860] = layer0_outputs[12414];
    assign layer1_outputs[3861] = ~(layer0_outputs[3319]) | (layer0_outputs[3108]);
    assign layer1_outputs[3862] = ~(layer0_outputs[4776]) | (layer0_outputs[8328]);
    assign layer1_outputs[3863] = ~(layer0_outputs[3057]);
    assign layer1_outputs[3864] = layer0_outputs[8546];
    assign layer1_outputs[3865] = ~(layer0_outputs[3204]) | (layer0_outputs[11719]);
    assign layer1_outputs[3866] = ~(layer0_outputs[1755]);
    assign layer1_outputs[3867] = (layer0_outputs[8609]) & ~(layer0_outputs[4591]);
    assign layer1_outputs[3868] = (layer0_outputs[4456]) & (layer0_outputs[5895]);
    assign layer1_outputs[3869] = (layer0_outputs[11971]) & ~(layer0_outputs[9868]);
    assign layer1_outputs[3870] = layer0_outputs[7098];
    assign layer1_outputs[3871] = (layer0_outputs[12148]) ^ (layer0_outputs[12719]);
    assign layer1_outputs[3872] = (layer0_outputs[12632]) & ~(layer0_outputs[12420]);
    assign layer1_outputs[3873] = (layer0_outputs[582]) & (layer0_outputs[7884]);
    assign layer1_outputs[3874] = layer0_outputs[4108];
    assign layer1_outputs[3875] = ~((layer0_outputs[6624]) & (layer0_outputs[9506]));
    assign layer1_outputs[3876] = ~(layer0_outputs[8463]);
    assign layer1_outputs[3877] = layer0_outputs[12071];
    assign layer1_outputs[3878] = ~((layer0_outputs[1558]) ^ (layer0_outputs[6969]));
    assign layer1_outputs[3879] = (layer0_outputs[1742]) & ~(layer0_outputs[8920]);
    assign layer1_outputs[3880] = 1'b0;
    assign layer1_outputs[3881] = ~(layer0_outputs[7052]);
    assign layer1_outputs[3882] = ~(layer0_outputs[10714]);
    assign layer1_outputs[3883] = ~(layer0_outputs[11760]);
    assign layer1_outputs[3884] = ~((layer0_outputs[5462]) & (layer0_outputs[10163]));
    assign layer1_outputs[3885] = ~(layer0_outputs[5287]);
    assign layer1_outputs[3886] = (layer0_outputs[4270]) & (layer0_outputs[4345]);
    assign layer1_outputs[3887] = ~((layer0_outputs[2612]) & (layer0_outputs[11592]));
    assign layer1_outputs[3888] = (layer0_outputs[2055]) & ~(layer0_outputs[10649]);
    assign layer1_outputs[3889] = (layer0_outputs[9405]) | (layer0_outputs[5506]);
    assign layer1_outputs[3890] = ~((layer0_outputs[5384]) ^ (layer0_outputs[889]));
    assign layer1_outputs[3891] = ~((layer0_outputs[11035]) ^ (layer0_outputs[780]));
    assign layer1_outputs[3892] = ~(layer0_outputs[964]) | (layer0_outputs[3134]);
    assign layer1_outputs[3893] = layer0_outputs[9595];
    assign layer1_outputs[3894] = ~(layer0_outputs[4704]);
    assign layer1_outputs[3895] = ~(layer0_outputs[3535]) | (layer0_outputs[494]);
    assign layer1_outputs[3896] = ~((layer0_outputs[8940]) ^ (layer0_outputs[9115]));
    assign layer1_outputs[3897] = ~(layer0_outputs[1806]);
    assign layer1_outputs[3898] = (layer0_outputs[5268]) ^ (layer0_outputs[1962]);
    assign layer1_outputs[3899] = ~(layer0_outputs[1167]);
    assign layer1_outputs[3900] = (layer0_outputs[12117]) & ~(layer0_outputs[12104]);
    assign layer1_outputs[3901] = layer0_outputs[814];
    assign layer1_outputs[3902] = (layer0_outputs[3553]) & (layer0_outputs[2590]);
    assign layer1_outputs[3903] = ~(layer0_outputs[8374]);
    assign layer1_outputs[3904] = (layer0_outputs[3839]) & ~(layer0_outputs[2409]);
    assign layer1_outputs[3905] = ~(layer0_outputs[10724]) | (layer0_outputs[9701]);
    assign layer1_outputs[3906] = ~(layer0_outputs[5394]) | (layer0_outputs[6987]);
    assign layer1_outputs[3907] = (layer0_outputs[4103]) ^ (layer0_outputs[11113]);
    assign layer1_outputs[3908] = layer0_outputs[3216];
    assign layer1_outputs[3909] = ~(layer0_outputs[4760]);
    assign layer1_outputs[3910] = ~((layer0_outputs[12332]) | (layer0_outputs[2555]));
    assign layer1_outputs[3911] = (layer0_outputs[2831]) | (layer0_outputs[5805]);
    assign layer1_outputs[3912] = ~(layer0_outputs[9873]) | (layer0_outputs[9530]);
    assign layer1_outputs[3913] = (layer0_outputs[7121]) & (layer0_outputs[1958]);
    assign layer1_outputs[3914] = ~(layer0_outputs[12612]);
    assign layer1_outputs[3915] = layer0_outputs[646];
    assign layer1_outputs[3916] = (layer0_outputs[6299]) & ~(layer0_outputs[7548]);
    assign layer1_outputs[3917] = (layer0_outputs[2148]) ^ (layer0_outputs[804]);
    assign layer1_outputs[3918] = ~((layer0_outputs[1736]) ^ (layer0_outputs[10565]));
    assign layer1_outputs[3919] = (layer0_outputs[12349]) ^ (layer0_outputs[1627]);
    assign layer1_outputs[3920] = ~(layer0_outputs[6100]);
    assign layer1_outputs[3921] = (layer0_outputs[2551]) | (layer0_outputs[7426]);
    assign layer1_outputs[3922] = ~(layer0_outputs[4973]);
    assign layer1_outputs[3923] = ~((layer0_outputs[545]) & (layer0_outputs[7274]));
    assign layer1_outputs[3924] = ~(layer0_outputs[160]);
    assign layer1_outputs[3925] = ~((layer0_outputs[5984]) & (layer0_outputs[4430]));
    assign layer1_outputs[3926] = ~((layer0_outputs[10041]) ^ (layer0_outputs[12586]));
    assign layer1_outputs[3927] = (layer0_outputs[481]) & (layer0_outputs[10673]);
    assign layer1_outputs[3928] = ~(layer0_outputs[7692]);
    assign layer1_outputs[3929] = ~(layer0_outputs[1185]);
    assign layer1_outputs[3930] = ~((layer0_outputs[5423]) & (layer0_outputs[8974]));
    assign layer1_outputs[3931] = ~((layer0_outputs[8760]) ^ (layer0_outputs[8423]));
    assign layer1_outputs[3932] = ~(layer0_outputs[1658]);
    assign layer1_outputs[3933] = (layer0_outputs[3347]) & ~(layer0_outputs[12183]);
    assign layer1_outputs[3934] = ~((layer0_outputs[4937]) | (layer0_outputs[1836]));
    assign layer1_outputs[3935] = ~(layer0_outputs[12404]);
    assign layer1_outputs[3936] = (layer0_outputs[7394]) & ~(layer0_outputs[7800]);
    assign layer1_outputs[3937] = layer0_outputs[9954];
    assign layer1_outputs[3938] = 1'b0;
    assign layer1_outputs[3939] = (layer0_outputs[11296]) & (layer0_outputs[12035]);
    assign layer1_outputs[3940] = (layer0_outputs[2543]) | (layer0_outputs[9957]);
    assign layer1_outputs[3941] = ~(layer0_outputs[484]) | (layer0_outputs[11041]);
    assign layer1_outputs[3942] = (layer0_outputs[4404]) & (layer0_outputs[3529]);
    assign layer1_outputs[3943] = ~(layer0_outputs[3949]);
    assign layer1_outputs[3944] = ~(layer0_outputs[283]);
    assign layer1_outputs[3945] = layer0_outputs[3035];
    assign layer1_outputs[3946] = (layer0_outputs[1190]) & ~(layer0_outputs[3840]);
    assign layer1_outputs[3947] = ~((layer0_outputs[2333]) ^ (layer0_outputs[6842]));
    assign layer1_outputs[3948] = (layer0_outputs[324]) & ~(layer0_outputs[5176]);
    assign layer1_outputs[3949] = ~(layer0_outputs[6275]) | (layer0_outputs[9227]);
    assign layer1_outputs[3950] = (layer0_outputs[8569]) & ~(layer0_outputs[3884]);
    assign layer1_outputs[3951] = (layer0_outputs[12789]) & ~(layer0_outputs[6408]);
    assign layer1_outputs[3952] = (layer0_outputs[8203]) ^ (layer0_outputs[3070]);
    assign layer1_outputs[3953] = ~(layer0_outputs[7977]);
    assign layer1_outputs[3954] = (layer0_outputs[4902]) ^ (layer0_outputs[6467]);
    assign layer1_outputs[3955] = (layer0_outputs[7039]) ^ (layer0_outputs[1473]);
    assign layer1_outputs[3956] = ~((layer0_outputs[914]) | (layer0_outputs[12283]));
    assign layer1_outputs[3957] = (layer0_outputs[12245]) & ~(layer0_outputs[5640]);
    assign layer1_outputs[3958] = layer0_outputs[1851];
    assign layer1_outputs[3959] = ~(layer0_outputs[7688]);
    assign layer1_outputs[3960] = (layer0_outputs[6360]) & ~(layer0_outputs[7120]);
    assign layer1_outputs[3961] = (layer0_outputs[12535]) ^ (layer0_outputs[12509]);
    assign layer1_outputs[3962] = ~(layer0_outputs[6673]);
    assign layer1_outputs[3963] = ~((layer0_outputs[1170]) | (layer0_outputs[12362]));
    assign layer1_outputs[3964] = ~(layer0_outputs[8478]);
    assign layer1_outputs[3965] = (layer0_outputs[6070]) & ~(layer0_outputs[11344]);
    assign layer1_outputs[3966] = ~((layer0_outputs[9323]) | (layer0_outputs[11244]));
    assign layer1_outputs[3967] = ~(layer0_outputs[6102]) | (layer0_outputs[5753]);
    assign layer1_outputs[3968] = ~(layer0_outputs[7202]);
    assign layer1_outputs[3969] = layer0_outputs[4477];
    assign layer1_outputs[3970] = ~(layer0_outputs[9989]) | (layer0_outputs[11829]);
    assign layer1_outputs[3971] = layer0_outputs[10238];
    assign layer1_outputs[3972] = (layer0_outputs[3621]) | (layer0_outputs[4417]);
    assign layer1_outputs[3973] = layer0_outputs[3763];
    assign layer1_outputs[3974] = layer0_outputs[4025];
    assign layer1_outputs[3975] = ~(layer0_outputs[75]);
    assign layer1_outputs[3976] = (layer0_outputs[11910]) & ~(layer0_outputs[1186]);
    assign layer1_outputs[3977] = ~(layer0_outputs[3382]) | (layer0_outputs[7053]);
    assign layer1_outputs[3978] = 1'b1;
    assign layer1_outputs[3979] = ~(layer0_outputs[10688]);
    assign layer1_outputs[3980] = (layer0_outputs[7012]) & ~(layer0_outputs[3787]);
    assign layer1_outputs[3981] = ~((layer0_outputs[1626]) | (layer0_outputs[5236]));
    assign layer1_outputs[3982] = ~((layer0_outputs[2158]) | (layer0_outputs[2572]));
    assign layer1_outputs[3983] = 1'b1;
    assign layer1_outputs[3984] = ~(layer0_outputs[2770]) | (layer0_outputs[12152]);
    assign layer1_outputs[3985] = ~(layer0_outputs[2992]);
    assign layer1_outputs[3986] = layer0_outputs[6942];
    assign layer1_outputs[3987] = 1'b1;
    assign layer1_outputs[3988] = layer0_outputs[6402];
    assign layer1_outputs[3989] = ~((layer0_outputs[3373]) & (layer0_outputs[7197]));
    assign layer1_outputs[3990] = (layer0_outputs[10188]) | (layer0_outputs[7831]);
    assign layer1_outputs[3991] = ~(layer0_outputs[11058]) | (layer0_outputs[4670]);
    assign layer1_outputs[3992] = ~(layer0_outputs[3266]) | (layer0_outputs[753]);
    assign layer1_outputs[3993] = 1'b0;
    assign layer1_outputs[3994] = ~(layer0_outputs[10596]) | (layer0_outputs[6724]);
    assign layer1_outputs[3995] = ~(layer0_outputs[8603]) | (layer0_outputs[3335]);
    assign layer1_outputs[3996] = 1'b0;
    assign layer1_outputs[3997] = (layer0_outputs[7740]) & ~(layer0_outputs[11751]);
    assign layer1_outputs[3998] = ~((layer0_outputs[8579]) | (layer0_outputs[9672]));
    assign layer1_outputs[3999] = layer0_outputs[4971];
    assign layer1_outputs[4000] = layer0_outputs[6190];
    assign layer1_outputs[4001] = ~(layer0_outputs[12516]);
    assign layer1_outputs[4002] = (layer0_outputs[11559]) | (layer0_outputs[10576]);
    assign layer1_outputs[4003] = layer0_outputs[10097];
    assign layer1_outputs[4004] = layer0_outputs[2053];
    assign layer1_outputs[4005] = (layer0_outputs[12766]) | (layer0_outputs[208]);
    assign layer1_outputs[4006] = ~((layer0_outputs[8886]) & (layer0_outputs[6287]));
    assign layer1_outputs[4007] = ~((layer0_outputs[681]) ^ (layer0_outputs[2654]));
    assign layer1_outputs[4008] = layer0_outputs[3137];
    assign layer1_outputs[4009] = ~(layer0_outputs[12164]);
    assign layer1_outputs[4010] = layer0_outputs[8651];
    assign layer1_outputs[4011] = (layer0_outputs[627]) & ~(layer0_outputs[8719]);
    assign layer1_outputs[4012] = ~(layer0_outputs[1323]);
    assign layer1_outputs[4013] = ~(layer0_outputs[769]);
    assign layer1_outputs[4014] = layer0_outputs[5925];
    assign layer1_outputs[4015] = (layer0_outputs[12241]) & (layer0_outputs[12099]);
    assign layer1_outputs[4016] = (layer0_outputs[8364]) & (layer0_outputs[6410]);
    assign layer1_outputs[4017] = (layer0_outputs[7130]) & ~(layer0_outputs[2235]);
    assign layer1_outputs[4018] = (layer0_outputs[9749]) & ~(layer0_outputs[8453]);
    assign layer1_outputs[4019] = (layer0_outputs[9999]) | (layer0_outputs[10022]);
    assign layer1_outputs[4020] = ~(layer0_outputs[8630]);
    assign layer1_outputs[4021] = layer0_outputs[5874];
    assign layer1_outputs[4022] = (layer0_outputs[4893]) ^ (layer0_outputs[12078]);
    assign layer1_outputs[4023] = ~((layer0_outputs[970]) ^ (layer0_outputs[3327]));
    assign layer1_outputs[4024] = layer0_outputs[233];
    assign layer1_outputs[4025] = ~(layer0_outputs[3622]);
    assign layer1_outputs[4026] = (layer0_outputs[5828]) | (layer0_outputs[3588]);
    assign layer1_outputs[4027] = ~((layer0_outputs[6779]) | (layer0_outputs[5044]));
    assign layer1_outputs[4028] = ~((layer0_outputs[3226]) & (layer0_outputs[818]));
    assign layer1_outputs[4029] = ~(layer0_outputs[11641]) | (layer0_outputs[8193]);
    assign layer1_outputs[4030] = layer0_outputs[5084];
    assign layer1_outputs[4031] = ~(layer0_outputs[5992]) | (layer0_outputs[2946]);
    assign layer1_outputs[4032] = ~(layer0_outputs[2097]);
    assign layer1_outputs[4033] = ~((layer0_outputs[4628]) & (layer0_outputs[5930]));
    assign layer1_outputs[4034] = ~(layer0_outputs[7955]);
    assign layer1_outputs[4035] = ~(layer0_outputs[8652]);
    assign layer1_outputs[4036] = ~(layer0_outputs[3025]);
    assign layer1_outputs[4037] = ~((layer0_outputs[7608]) & (layer0_outputs[1287]));
    assign layer1_outputs[4038] = layer0_outputs[5488];
    assign layer1_outputs[4039] = (layer0_outputs[7822]) | (layer0_outputs[6940]);
    assign layer1_outputs[4040] = layer0_outputs[7445];
    assign layer1_outputs[4041] = layer0_outputs[12603];
    assign layer1_outputs[4042] = ~(layer0_outputs[12451]);
    assign layer1_outputs[4043] = layer0_outputs[6418];
    assign layer1_outputs[4044] = ~(layer0_outputs[6220]) | (layer0_outputs[7863]);
    assign layer1_outputs[4045] = (layer0_outputs[8851]) ^ (layer0_outputs[9014]);
    assign layer1_outputs[4046] = ~(layer0_outputs[4065]);
    assign layer1_outputs[4047] = ~(layer0_outputs[7311]);
    assign layer1_outputs[4048] = (layer0_outputs[9699]) ^ (layer0_outputs[10519]);
    assign layer1_outputs[4049] = (layer0_outputs[9026]) & ~(layer0_outputs[290]);
    assign layer1_outputs[4050] = ~((layer0_outputs[7052]) & (layer0_outputs[7856]));
    assign layer1_outputs[4051] = ~(layer0_outputs[1625]) | (layer0_outputs[2421]);
    assign layer1_outputs[4052] = (layer0_outputs[3595]) & ~(layer0_outputs[6765]);
    assign layer1_outputs[4053] = layer0_outputs[3643];
    assign layer1_outputs[4054] = ~((layer0_outputs[2807]) & (layer0_outputs[1764]));
    assign layer1_outputs[4055] = (layer0_outputs[97]) & (layer0_outputs[4752]);
    assign layer1_outputs[4056] = ~(layer0_outputs[3367]);
    assign layer1_outputs[4057] = layer0_outputs[16];
    assign layer1_outputs[4058] = ~(layer0_outputs[9026]);
    assign layer1_outputs[4059] = ~((layer0_outputs[5844]) | (layer0_outputs[12163]));
    assign layer1_outputs[4060] = ~(layer0_outputs[896]);
    assign layer1_outputs[4061] = layer0_outputs[7877];
    assign layer1_outputs[4062] = layer0_outputs[10666];
    assign layer1_outputs[4063] = ~(layer0_outputs[8990]);
    assign layer1_outputs[4064] = ~((layer0_outputs[6952]) & (layer0_outputs[5598]));
    assign layer1_outputs[4065] = (layer0_outputs[5839]) ^ (layer0_outputs[2527]);
    assign layer1_outputs[4066] = (layer0_outputs[8733]) | (layer0_outputs[967]);
    assign layer1_outputs[4067] = ~(layer0_outputs[10471]);
    assign layer1_outputs[4068] = ~(layer0_outputs[1494]);
    assign layer1_outputs[4069] = ~(layer0_outputs[6450]);
    assign layer1_outputs[4070] = (layer0_outputs[4606]) & (layer0_outputs[11524]);
    assign layer1_outputs[4071] = ~(layer0_outputs[11354]);
    assign layer1_outputs[4072] = 1'b0;
    assign layer1_outputs[4073] = ~(layer0_outputs[4419]);
    assign layer1_outputs[4074] = (layer0_outputs[10560]) & ~(layer0_outputs[6634]);
    assign layer1_outputs[4075] = ~(layer0_outputs[355]);
    assign layer1_outputs[4076] = ~((layer0_outputs[6823]) | (layer0_outputs[9415]));
    assign layer1_outputs[4077] = layer0_outputs[8643];
    assign layer1_outputs[4078] = ~(layer0_outputs[521]) | (layer0_outputs[3514]);
    assign layer1_outputs[4079] = 1'b0;
    assign layer1_outputs[4080] = layer0_outputs[5175];
    assign layer1_outputs[4081] = (layer0_outputs[10833]) & ~(layer0_outputs[5776]);
    assign layer1_outputs[4082] = ~((layer0_outputs[8187]) ^ (layer0_outputs[1524]));
    assign layer1_outputs[4083] = layer0_outputs[1801];
    assign layer1_outputs[4084] = layer0_outputs[503];
    assign layer1_outputs[4085] = (layer0_outputs[1615]) | (layer0_outputs[8090]);
    assign layer1_outputs[4086] = 1'b1;
    assign layer1_outputs[4087] = layer0_outputs[10866];
    assign layer1_outputs[4088] = ~(layer0_outputs[710]);
    assign layer1_outputs[4089] = (layer0_outputs[12459]) & (layer0_outputs[8757]);
    assign layer1_outputs[4090] = layer0_outputs[5443];
    assign layer1_outputs[4091] = (layer0_outputs[11612]) | (layer0_outputs[4657]);
    assign layer1_outputs[4092] = layer0_outputs[82];
    assign layer1_outputs[4093] = ~(layer0_outputs[8291]) | (layer0_outputs[5991]);
    assign layer1_outputs[4094] = (layer0_outputs[1737]) & ~(layer0_outputs[4165]);
    assign layer1_outputs[4095] = ~((layer0_outputs[3524]) | (layer0_outputs[5410]));
    assign layer1_outputs[4096] = (layer0_outputs[11971]) ^ (layer0_outputs[6737]);
    assign layer1_outputs[4097] = ~(layer0_outputs[4536]);
    assign layer1_outputs[4098] = (layer0_outputs[365]) & ~(layer0_outputs[12165]);
    assign layer1_outputs[4099] = ~(layer0_outputs[9439]);
    assign layer1_outputs[4100] = (layer0_outputs[2511]) & (layer0_outputs[6308]);
    assign layer1_outputs[4101] = (layer0_outputs[2751]) & ~(layer0_outputs[5031]);
    assign layer1_outputs[4102] = ~(layer0_outputs[4030]);
    assign layer1_outputs[4103] = layer0_outputs[2138];
    assign layer1_outputs[4104] = layer0_outputs[10965];
    assign layer1_outputs[4105] = ~(layer0_outputs[4036]) | (layer0_outputs[2596]);
    assign layer1_outputs[4106] = ~(layer0_outputs[4222]) | (layer0_outputs[6832]);
    assign layer1_outputs[4107] = ~(layer0_outputs[7860]) | (layer0_outputs[2312]);
    assign layer1_outputs[4108] = ~(layer0_outputs[11260]);
    assign layer1_outputs[4109] = (layer0_outputs[5679]) & (layer0_outputs[11821]);
    assign layer1_outputs[4110] = ~((layer0_outputs[5483]) & (layer0_outputs[9267]));
    assign layer1_outputs[4111] = layer0_outputs[8877];
    assign layer1_outputs[4112] = ~((layer0_outputs[10309]) | (layer0_outputs[8503]));
    assign layer1_outputs[4113] = (layer0_outputs[8422]) & (layer0_outputs[8651]);
    assign layer1_outputs[4114] = ~((layer0_outputs[12469]) | (layer0_outputs[11773]));
    assign layer1_outputs[4115] = 1'b1;
    assign layer1_outputs[4116] = (layer0_outputs[907]) & ~(layer0_outputs[4254]);
    assign layer1_outputs[4117] = layer0_outputs[679];
    assign layer1_outputs[4118] = ~(layer0_outputs[2003]);
    assign layer1_outputs[4119] = layer0_outputs[1671];
    assign layer1_outputs[4120] = layer0_outputs[408];
    assign layer1_outputs[4121] = ~((layer0_outputs[4602]) & (layer0_outputs[4967]));
    assign layer1_outputs[4122] = 1'b0;
    assign layer1_outputs[4123] = (layer0_outputs[11886]) & ~(layer0_outputs[9886]);
    assign layer1_outputs[4124] = ~(layer0_outputs[5612]) | (layer0_outputs[10002]);
    assign layer1_outputs[4125] = (layer0_outputs[51]) & ~(layer0_outputs[10365]);
    assign layer1_outputs[4126] = layer0_outputs[617];
    assign layer1_outputs[4127] = ~(layer0_outputs[3011]) | (layer0_outputs[2945]);
    assign layer1_outputs[4128] = layer0_outputs[9396];
    assign layer1_outputs[4129] = (layer0_outputs[11165]) & ~(layer0_outputs[12088]);
    assign layer1_outputs[4130] = ~(layer0_outputs[4730]);
    assign layer1_outputs[4131] = ~(layer0_outputs[12217]) | (layer0_outputs[5037]);
    assign layer1_outputs[4132] = (layer0_outputs[6006]) & (layer0_outputs[12379]);
    assign layer1_outputs[4133] = ~((layer0_outputs[11434]) ^ (layer0_outputs[8769]));
    assign layer1_outputs[4134] = (layer0_outputs[11415]) & ~(layer0_outputs[2338]);
    assign layer1_outputs[4135] = (layer0_outputs[4312]) & (layer0_outputs[5011]);
    assign layer1_outputs[4136] = ~(layer0_outputs[10225]) | (layer0_outputs[2973]);
    assign layer1_outputs[4137] = (layer0_outputs[227]) & (layer0_outputs[4779]);
    assign layer1_outputs[4138] = layer0_outputs[106];
    assign layer1_outputs[4139] = (layer0_outputs[193]) ^ (layer0_outputs[5154]);
    assign layer1_outputs[4140] = layer0_outputs[5302];
    assign layer1_outputs[4141] = ~((layer0_outputs[10081]) ^ (layer0_outputs[5832]));
    assign layer1_outputs[4142] = ~(layer0_outputs[942]);
    assign layer1_outputs[4143] = (layer0_outputs[8518]) & ~(layer0_outputs[8764]);
    assign layer1_outputs[4144] = 1'b0;
    assign layer1_outputs[4145] = layer0_outputs[9368];
    assign layer1_outputs[4146] = ~(layer0_outputs[11172]) | (layer0_outputs[6517]);
    assign layer1_outputs[4147] = ~(layer0_outputs[1687]);
    assign layer1_outputs[4148] = layer0_outputs[12075];
    assign layer1_outputs[4149] = layer0_outputs[2166];
    assign layer1_outputs[4150] = 1'b1;
    assign layer1_outputs[4151] = (layer0_outputs[5029]) ^ (layer0_outputs[10686]);
    assign layer1_outputs[4152] = layer0_outputs[11945];
    assign layer1_outputs[4153] = ~(layer0_outputs[1292]);
    assign layer1_outputs[4154] = ~((layer0_outputs[644]) ^ (layer0_outputs[10915]));
    assign layer1_outputs[4155] = ~((layer0_outputs[12242]) | (layer0_outputs[5774]));
    assign layer1_outputs[4156] = ~(layer0_outputs[10247]) | (layer0_outputs[4988]);
    assign layer1_outputs[4157] = ~(layer0_outputs[6238]);
    assign layer1_outputs[4158] = ~((layer0_outputs[2390]) & (layer0_outputs[4106]));
    assign layer1_outputs[4159] = ~((layer0_outputs[8979]) & (layer0_outputs[812]));
    assign layer1_outputs[4160] = ~((layer0_outputs[2802]) | (layer0_outputs[4234]));
    assign layer1_outputs[4161] = (layer0_outputs[12569]) | (layer0_outputs[11390]);
    assign layer1_outputs[4162] = ~((layer0_outputs[276]) ^ (layer0_outputs[5677]));
    assign layer1_outputs[4163] = ~(layer0_outputs[10124]);
    assign layer1_outputs[4164] = ~((layer0_outputs[5690]) & (layer0_outputs[3346]));
    assign layer1_outputs[4165] = ~(layer0_outputs[5853]) | (layer0_outputs[9428]);
    assign layer1_outputs[4166] = ~(layer0_outputs[7699]);
    assign layer1_outputs[4167] = (layer0_outputs[8785]) & (layer0_outputs[10354]);
    assign layer1_outputs[4168] = (layer0_outputs[12579]) & ~(layer0_outputs[7412]);
    assign layer1_outputs[4169] = layer0_outputs[6595];
    assign layer1_outputs[4170] = (layer0_outputs[11153]) | (layer0_outputs[6609]);
    assign layer1_outputs[4171] = ~(layer0_outputs[974]);
    assign layer1_outputs[4172] = ~(layer0_outputs[6526]);
    assign layer1_outputs[4173] = (layer0_outputs[5956]) | (layer0_outputs[11247]);
    assign layer1_outputs[4174] = layer0_outputs[7524];
    assign layer1_outputs[4175] = ~(layer0_outputs[3663]);
    assign layer1_outputs[4176] = ~(layer0_outputs[4918]);
    assign layer1_outputs[4177] = (layer0_outputs[646]) & (layer0_outputs[4232]);
    assign layer1_outputs[4178] = ~(layer0_outputs[4225]);
    assign layer1_outputs[4179] = ~(layer0_outputs[12728]);
    assign layer1_outputs[4180] = (layer0_outputs[1629]) & ~(layer0_outputs[4348]);
    assign layer1_outputs[4181] = ~(layer0_outputs[9467]) | (layer0_outputs[4067]);
    assign layer1_outputs[4182] = layer0_outputs[7576];
    assign layer1_outputs[4183] = layer0_outputs[7975];
    assign layer1_outputs[4184] = ~((layer0_outputs[5873]) & (layer0_outputs[0]));
    assign layer1_outputs[4185] = ~(layer0_outputs[865]);
    assign layer1_outputs[4186] = ~(layer0_outputs[159]);
    assign layer1_outputs[4187] = (layer0_outputs[12232]) & ~(layer0_outputs[5496]);
    assign layer1_outputs[4188] = (layer0_outputs[11089]) & ~(layer0_outputs[12013]);
    assign layer1_outputs[4189] = ~((layer0_outputs[9739]) & (layer0_outputs[6836]));
    assign layer1_outputs[4190] = (layer0_outputs[7774]) | (layer0_outputs[7759]);
    assign layer1_outputs[4191] = (layer0_outputs[7613]) ^ (layer0_outputs[517]);
    assign layer1_outputs[4192] = ~(layer0_outputs[10252]) | (layer0_outputs[2104]);
    assign layer1_outputs[4193] = (layer0_outputs[1656]) | (layer0_outputs[8154]);
    assign layer1_outputs[4194] = ~(layer0_outputs[3247]);
    assign layer1_outputs[4195] = layer0_outputs[12032];
    assign layer1_outputs[4196] = 1'b0;
    assign layer1_outputs[4197] = layer0_outputs[2336];
    assign layer1_outputs[4198] = (layer0_outputs[8457]) & (layer0_outputs[5658]);
    assign layer1_outputs[4199] = ~(layer0_outputs[12748]);
    assign layer1_outputs[4200] = layer0_outputs[6092];
    assign layer1_outputs[4201] = (layer0_outputs[11600]) | (layer0_outputs[9113]);
    assign layer1_outputs[4202] = ~(layer0_outputs[3338]) | (layer0_outputs[2764]);
    assign layer1_outputs[4203] = layer0_outputs[3717];
    assign layer1_outputs[4204] = (layer0_outputs[10631]) | (layer0_outputs[4738]);
    assign layer1_outputs[4205] = (layer0_outputs[5024]) & ~(layer0_outputs[9967]);
    assign layer1_outputs[4206] = (layer0_outputs[2038]) & (layer0_outputs[792]);
    assign layer1_outputs[4207] = 1'b0;
    assign layer1_outputs[4208] = (layer0_outputs[6141]) & ~(layer0_outputs[11960]);
    assign layer1_outputs[4209] = (layer0_outputs[1239]) ^ (layer0_outputs[12137]);
    assign layer1_outputs[4210] = ~((layer0_outputs[2416]) & (layer0_outputs[8584]));
    assign layer1_outputs[4211] = ~(layer0_outputs[2284]) | (layer0_outputs[11892]);
    assign layer1_outputs[4212] = (layer0_outputs[6239]) | (layer0_outputs[3053]);
    assign layer1_outputs[4213] = ~((layer0_outputs[9085]) ^ (layer0_outputs[6453]));
    assign layer1_outputs[4214] = layer0_outputs[1069];
    assign layer1_outputs[4215] = (layer0_outputs[6795]) & ~(layer0_outputs[7641]);
    assign layer1_outputs[4216] = layer0_outputs[8072];
    assign layer1_outputs[4217] = ~((layer0_outputs[5846]) ^ (layer0_outputs[11951]));
    assign layer1_outputs[4218] = layer0_outputs[11171];
    assign layer1_outputs[4219] = (layer0_outputs[12554]) & ~(layer0_outputs[6949]);
    assign layer1_outputs[4220] = ~(layer0_outputs[5735]);
    assign layer1_outputs[4221] = layer0_outputs[11597];
    assign layer1_outputs[4222] = ~(layer0_outputs[11747]);
    assign layer1_outputs[4223] = ~(layer0_outputs[757]);
    assign layer1_outputs[4224] = ~(layer0_outputs[11500]);
    assign layer1_outputs[4225] = (layer0_outputs[8671]) & ~(layer0_outputs[12021]);
    assign layer1_outputs[4226] = ~((layer0_outputs[4815]) | (layer0_outputs[9164]));
    assign layer1_outputs[4227] = (layer0_outputs[2678]) & ~(layer0_outputs[1850]);
    assign layer1_outputs[4228] = ~(layer0_outputs[11604]);
    assign layer1_outputs[4229] = layer0_outputs[3060];
    assign layer1_outputs[4230] = (layer0_outputs[5648]) | (layer0_outputs[6121]);
    assign layer1_outputs[4231] = ~(layer0_outputs[10539]);
    assign layer1_outputs[4232] = ~((layer0_outputs[3982]) | (layer0_outputs[357]));
    assign layer1_outputs[4233] = (layer0_outputs[3495]) & (layer0_outputs[3794]);
    assign layer1_outputs[4234] = ~(layer0_outputs[7071]);
    assign layer1_outputs[4235] = layer0_outputs[3459];
    assign layer1_outputs[4236] = ~(layer0_outputs[8661]);
    assign layer1_outputs[4237] = ~(layer0_outputs[2070]) | (layer0_outputs[1186]);
    assign layer1_outputs[4238] = layer0_outputs[1029];
    assign layer1_outputs[4239] = ~(layer0_outputs[2695]) | (layer0_outputs[8714]);
    assign layer1_outputs[4240] = (layer0_outputs[9556]) ^ (layer0_outputs[12540]);
    assign layer1_outputs[4241] = ~((layer0_outputs[4224]) ^ (layer0_outputs[12597]));
    assign layer1_outputs[4242] = ~((layer0_outputs[3721]) & (layer0_outputs[7864]));
    assign layer1_outputs[4243] = ~(layer0_outputs[11757]);
    assign layer1_outputs[4244] = (layer0_outputs[12437]) & ~(layer0_outputs[6824]);
    assign layer1_outputs[4245] = (layer0_outputs[6572]) & ~(layer0_outputs[2488]);
    assign layer1_outputs[4246] = 1'b0;
    assign layer1_outputs[4247] = ~((layer0_outputs[11121]) ^ (layer0_outputs[5845]));
    assign layer1_outputs[4248] = ~(layer0_outputs[1819]) | (layer0_outputs[1924]);
    assign layer1_outputs[4249] = ~((layer0_outputs[9684]) & (layer0_outputs[1376]));
    assign layer1_outputs[4250] = layer0_outputs[2881];
    assign layer1_outputs[4251] = ~(layer0_outputs[7902]);
    assign layer1_outputs[4252] = (layer0_outputs[5201]) & (layer0_outputs[2699]);
    assign layer1_outputs[4253] = ~(layer0_outputs[3708]);
    assign layer1_outputs[4254] = ~(layer0_outputs[2625]);
    assign layer1_outputs[4255] = ~(layer0_outputs[9635]);
    assign layer1_outputs[4256] = (layer0_outputs[12778]) | (layer0_outputs[8539]);
    assign layer1_outputs[4257] = ~((layer0_outputs[2001]) & (layer0_outputs[317]));
    assign layer1_outputs[4258] = layer0_outputs[3687];
    assign layer1_outputs[4259] = ~((layer0_outputs[2840]) & (layer0_outputs[2977]));
    assign layer1_outputs[4260] = layer0_outputs[1897];
    assign layer1_outputs[4261] = ~(layer0_outputs[4883]);
    assign layer1_outputs[4262] = ~((layer0_outputs[11555]) & (layer0_outputs[5210]));
    assign layer1_outputs[4263] = (layer0_outputs[9057]) & ~(layer0_outputs[9202]);
    assign layer1_outputs[4264] = ~(layer0_outputs[4782]);
    assign layer1_outputs[4265] = ~((layer0_outputs[5306]) | (layer0_outputs[11308]));
    assign layer1_outputs[4266] = ~(layer0_outputs[11769]);
    assign layer1_outputs[4267] = ~((layer0_outputs[10211]) ^ (layer0_outputs[10003]));
    assign layer1_outputs[4268] = (layer0_outputs[6817]) & ~(layer0_outputs[7234]);
    assign layer1_outputs[4269] = (layer0_outputs[11033]) | (layer0_outputs[8222]);
    assign layer1_outputs[4270] = ~(layer0_outputs[155]) | (layer0_outputs[607]);
    assign layer1_outputs[4271] = ~(layer0_outputs[7625]);
    assign layer1_outputs[4272] = ~(layer0_outputs[10280]);
    assign layer1_outputs[4273] = ~(layer0_outputs[4343]);
    assign layer1_outputs[4274] = ~((layer0_outputs[6069]) & (layer0_outputs[7446]));
    assign layer1_outputs[4275] = (layer0_outputs[9915]) & ~(layer0_outputs[8890]);
    assign layer1_outputs[4276] = ~((layer0_outputs[2376]) ^ (layer0_outputs[4541]));
    assign layer1_outputs[4277] = (layer0_outputs[10265]) & ~(layer0_outputs[9053]);
    assign layer1_outputs[4278] = layer0_outputs[7812];
    assign layer1_outputs[4279] = layer0_outputs[2786];
    assign layer1_outputs[4280] = ~(layer0_outputs[7355]);
    assign layer1_outputs[4281] = layer0_outputs[1716];
    assign layer1_outputs[4282] = layer0_outputs[11109];
    assign layer1_outputs[4283] = layer0_outputs[6655];
    assign layer1_outputs[4284] = (layer0_outputs[3493]) | (layer0_outputs[5668]);
    assign layer1_outputs[4285] = layer0_outputs[2939];
    assign layer1_outputs[4286] = ~(layer0_outputs[6161]);
    assign layer1_outputs[4287] = (layer0_outputs[5405]) ^ (layer0_outputs[1459]);
    assign layer1_outputs[4288] = ~(layer0_outputs[6393]);
    assign layer1_outputs[4289] = ~(layer0_outputs[10391]);
    assign layer1_outputs[4290] = ~((layer0_outputs[6384]) ^ (layer0_outputs[708]));
    assign layer1_outputs[4291] = ~(layer0_outputs[7717]);
    assign layer1_outputs[4292] = ~((layer0_outputs[5988]) & (layer0_outputs[8029]));
    assign layer1_outputs[4293] = ~(layer0_outputs[8265]);
    assign layer1_outputs[4294] = layer0_outputs[6362];
    assign layer1_outputs[4295] = ~(layer0_outputs[2175]);
    assign layer1_outputs[4296] = ~(layer0_outputs[11228]);
    assign layer1_outputs[4297] = ~((layer0_outputs[10838]) ^ (layer0_outputs[5135]));
    assign layer1_outputs[4298] = (layer0_outputs[5245]) ^ (layer0_outputs[5663]);
    assign layer1_outputs[4299] = (layer0_outputs[6082]) & ~(layer0_outputs[1046]);
    assign layer1_outputs[4300] = ~((layer0_outputs[5712]) | (layer0_outputs[10179]));
    assign layer1_outputs[4301] = layer0_outputs[7485];
    assign layer1_outputs[4302] = (layer0_outputs[2972]) | (layer0_outputs[7516]);
    assign layer1_outputs[4303] = ~(layer0_outputs[6676]);
    assign layer1_outputs[4304] = (layer0_outputs[10684]) | (layer0_outputs[11634]);
    assign layer1_outputs[4305] = (layer0_outputs[11426]) & ~(layer0_outputs[4081]);
    assign layer1_outputs[4306] = ~((layer0_outputs[11711]) | (layer0_outputs[11763]));
    assign layer1_outputs[4307] = (layer0_outputs[12420]) ^ (layer0_outputs[10420]);
    assign layer1_outputs[4308] = layer0_outputs[4447];
    assign layer1_outputs[4309] = ~(layer0_outputs[5232]) | (layer0_outputs[10037]);
    assign layer1_outputs[4310] = ~(layer0_outputs[10936]);
    assign layer1_outputs[4311] = (layer0_outputs[11664]) ^ (layer0_outputs[7250]);
    assign layer1_outputs[4312] = ~(layer0_outputs[12593]) | (layer0_outputs[4554]);
    assign layer1_outputs[4313] = (layer0_outputs[9897]) ^ (layer0_outputs[9286]);
    assign layer1_outputs[4314] = ~((layer0_outputs[2493]) ^ (layer0_outputs[6837]));
    assign layer1_outputs[4315] = ~(layer0_outputs[5149]);
    assign layer1_outputs[4316] = ~((layer0_outputs[9247]) ^ (layer0_outputs[8391]));
    assign layer1_outputs[4317] = layer0_outputs[8301];
    assign layer1_outputs[4318] = ~(layer0_outputs[12657]) | (layer0_outputs[4391]);
    assign layer1_outputs[4319] = layer0_outputs[3462];
    assign layer1_outputs[4320] = ~((layer0_outputs[11425]) ^ (layer0_outputs[4172]));
    assign layer1_outputs[4321] = ~((layer0_outputs[900]) | (layer0_outputs[10423]));
    assign layer1_outputs[4322] = 1'b1;
    assign layer1_outputs[4323] = ~(layer0_outputs[6220]) | (layer0_outputs[8738]);
    assign layer1_outputs[4324] = ~(layer0_outputs[10793]);
    assign layer1_outputs[4325] = ~((layer0_outputs[6135]) | (layer0_outputs[9652]));
    assign layer1_outputs[4326] = layer0_outputs[4936];
    assign layer1_outputs[4327] = ~(layer0_outputs[10490]) | (layer0_outputs[11835]);
    assign layer1_outputs[4328] = (layer0_outputs[3931]) & (layer0_outputs[3100]);
    assign layer1_outputs[4329] = layer0_outputs[12430];
    assign layer1_outputs[4330] = (layer0_outputs[10993]) & (layer0_outputs[9877]);
    assign layer1_outputs[4331] = layer0_outputs[5121];
    assign layer1_outputs[4332] = ~((layer0_outputs[6193]) & (layer0_outputs[7390]));
    assign layer1_outputs[4333] = layer0_outputs[3606];
    assign layer1_outputs[4334] = ~((layer0_outputs[4736]) & (layer0_outputs[1219]));
    assign layer1_outputs[4335] = ~((layer0_outputs[3610]) ^ (layer0_outputs[4943]));
    assign layer1_outputs[4336] = ~(layer0_outputs[5759]);
    assign layer1_outputs[4337] = ~(layer0_outputs[5866]);
    assign layer1_outputs[4338] = (layer0_outputs[7379]) & (layer0_outputs[5005]);
    assign layer1_outputs[4339] = (layer0_outputs[6173]) ^ (layer0_outputs[5969]);
    assign layer1_outputs[4340] = ~(layer0_outputs[3675]) | (layer0_outputs[1771]);
    assign layer1_outputs[4341] = layer0_outputs[11814];
    assign layer1_outputs[4342] = (layer0_outputs[60]) | (layer0_outputs[6552]);
    assign layer1_outputs[4343] = (layer0_outputs[12525]) & ~(layer0_outputs[4198]);
    assign layer1_outputs[4344] = ~(layer0_outputs[238]) | (layer0_outputs[1181]);
    assign layer1_outputs[4345] = ~((layer0_outputs[2470]) | (layer0_outputs[3251]));
    assign layer1_outputs[4346] = ~(layer0_outputs[12779]);
    assign layer1_outputs[4347] = ~(layer0_outputs[917]);
    assign layer1_outputs[4348] = ~((layer0_outputs[12031]) | (layer0_outputs[11283]));
    assign layer1_outputs[4349] = 1'b0;
    assign layer1_outputs[4350] = (layer0_outputs[2170]) & (layer0_outputs[8525]);
    assign layer1_outputs[4351] = layer0_outputs[9792];
    assign layer1_outputs[4352] = ~((layer0_outputs[5470]) ^ (layer0_outputs[3019]));
    assign layer1_outputs[4353] = ~(layer0_outputs[8175]) | (layer0_outputs[6521]);
    assign layer1_outputs[4354] = ~(layer0_outputs[9862]);
    assign layer1_outputs[4355] = (layer0_outputs[5687]) & ~(layer0_outputs[1886]);
    assign layer1_outputs[4356] = ~(layer0_outputs[4689]) | (layer0_outputs[5474]);
    assign layer1_outputs[4357] = 1'b1;
    assign layer1_outputs[4358] = ~(layer0_outputs[960]);
    assign layer1_outputs[4359] = layer0_outputs[3878];
    assign layer1_outputs[4360] = (layer0_outputs[12625]) & ~(layer0_outputs[7324]);
    assign layer1_outputs[4361] = layer0_outputs[10584];
    assign layer1_outputs[4362] = ~((layer0_outputs[11775]) & (layer0_outputs[10581]));
    assign layer1_outputs[4363] = (layer0_outputs[7998]) | (layer0_outputs[10932]);
    assign layer1_outputs[4364] = layer0_outputs[5630];
    assign layer1_outputs[4365] = 1'b0;
    assign layer1_outputs[4366] = ~((layer0_outputs[7568]) & (layer0_outputs[12751]));
    assign layer1_outputs[4367] = ~((layer0_outputs[5456]) | (layer0_outputs[5103]));
    assign layer1_outputs[4368] = (layer0_outputs[11301]) & (layer0_outputs[5980]);
    assign layer1_outputs[4369] = (layer0_outputs[9504]) & ~(layer0_outputs[12626]);
    assign layer1_outputs[4370] = layer0_outputs[3739];
    assign layer1_outputs[4371] = ~((layer0_outputs[4150]) ^ (layer0_outputs[12084]));
    assign layer1_outputs[4372] = ~(layer0_outputs[6235]);
    assign layer1_outputs[4373] = layer0_outputs[2202];
    assign layer1_outputs[4374] = ~((layer0_outputs[10629]) | (layer0_outputs[9311]));
    assign layer1_outputs[4375] = ~(layer0_outputs[11466]);
    assign layer1_outputs[4376] = ~(layer0_outputs[11342]);
    assign layer1_outputs[4377] = ~(layer0_outputs[9298]);
    assign layer1_outputs[4378] = ~((layer0_outputs[10996]) & (layer0_outputs[11640]));
    assign layer1_outputs[4379] = ~(layer0_outputs[11556]);
    assign layer1_outputs[4380] = ~(layer0_outputs[5086]);
    assign layer1_outputs[4381] = ~((layer0_outputs[1275]) & (layer0_outputs[10920]));
    assign layer1_outputs[4382] = ~(layer0_outputs[12089]) | (layer0_outputs[5052]);
    assign layer1_outputs[4383] = ~((layer0_outputs[1760]) ^ (layer0_outputs[12675]));
    assign layer1_outputs[4384] = (layer0_outputs[597]) & ~(layer0_outputs[6335]);
    assign layer1_outputs[4385] = layer0_outputs[9391];
    assign layer1_outputs[4386] = ~(layer0_outputs[7070]) | (layer0_outputs[7089]);
    assign layer1_outputs[4387] = layer0_outputs[894];
    assign layer1_outputs[4388] = ~((layer0_outputs[5908]) & (layer0_outputs[1743]));
    assign layer1_outputs[4389] = ~(layer0_outputs[5105]);
    assign layer1_outputs[4390] = ~(layer0_outputs[9353]);
    assign layer1_outputs[4391] = ~((layer0_outputs[7767]) | (layer0_outputs[9094]));
    assign layer1_outputs[4392] = ~(layer0_outputs[10056]);
    assign layer1_outputs[4393] = ~(layer0_outputs[77]) | (layer0_outputs[5714]);
    assign layer1_outputs[4394] = 1'b1;
    assign layer1_outputs[4395] = layer0_outputs[2628];
    assign layer1_outputs[4396] = (layer0_outputs[1121]) ^ (layer0_outputs[12330]);
    assign layer1_outputs[4397] = layer0_outputs[2554];
    assign layer1_outputs[4398] = layer0_outputs[5922];
    assign layer1_outputs[4399] = ~(layer0_outputs[11739]);
    assign layer1_outputs[4400] = layer0_outputs[3749];
    assign layer1_outputs[4401] = layer0_outputs[12570];
    assign layer1_outputs[4402] = (layer0_outputs[10675]) & ~(layer0_outputs[1384]);
    assign layer1_outputs[4403] = ~((layer0_outputs[9400]) | (layer0_outputs[9957]));
    assign layer1_outputs[4404] = (layer0_outputs[6213]) ^ (layer0_outputs[9042]);
    assign layer1_outputs[4405] = ~((layer0_outputs[5202]) & (layer0_outputs[5594]));
    assign layer1_outputs[4406] = layer0_outputs[9631];
    assign layer1_outputs[4407] = layer0_outputs[10114];
    assign layer1_outputs[4408] = ~(layer0_outputs[2473]);
    assign layer1_outputs[4409] = layer0_outputs[11317];
    assign layer1_outputs[4410] = layer0_outputs[3936];
    assign layer1_outputs[4411] = ~((layer0_outputs[9044]) | (layer0_outputs[7747]));
    assign layer1_outputs[4412] = layer0_outputs[3976];
    assign layer1_outputs[4413] = layer0_outputs[8399];
    assign layer1_outputs[4414] = (layer0_outputs[4050]) & ~(layer0_outputs[748]);
    assign layer1_outputs[4415] = ~((layer0_outputs[8373]) ^ (layer0_outputs[11167]));
    assign layer1_outputs[4416] = ~(layer0_outputs[10330]);
    assign layer1_outputs[4417] = ~(layer0_outputs[4532]);
    assign layer1_outputs[4418] = ~(layer0_outputs[11048]);
    assign layer1_outputs[4419] = layer0_outputs[5726];
    assign layer1_outputs[4420] = layer0_outputs[8177];
    assign layer1_outputs[4421] = (layer0_outputs[10860]) & ~(layer0_outputs[8902]);
    assign layer1_outputs[4422] = ~(layer0_outputs[6051]) | (layer0_outputs[10053]);
    assign layer1_outputs[4423] = ~(layer0_outputs[7016]) | (layer0_outputs[12530]);
    assign layer1_outputs[4424] = layer0_outputs[4584];
    assign layer1_outputs[4425] = ~(layer0_outputs[9090]) | (layer0_outputs[1429]);
    assign layer1_outputs[4426] = (layer0_outputs[7444]) & ~(layer0_outputs[4103]);
    assign layer1_outputs[4427] = ~(layer0_outputs[4892]) | (layer0_outputs[7865]);
    assign layer1_outputs[4428] = ~((layer0_outputs[10717]) | (layer0_outputs[9081]));
    assign layer1_outputs[4429] = layer0_outputs[2693];
    assign layer1_outputs[4430] = ~((layer0_outputs[6041]) & (layer0_outputs[11100]));
    assign layer1_outputs[4431] = (layer0_outputs[10346]) ^ (layer0_outputs[6854]);
    assign layer1_outputs[4432] = (layer0_outputs[8694]) ^ (layer0_outputs[6715]);
    assign layer1_outputs[4433] = layer0_outputs[3914];
    assign layer1_outputs[4434] = layer0_outputs[2253];
    assign layer1_outputs[4435] = (layer0_outputs[4280]) & ~(layer0_outputs[5997]);
    assign layer1_outputs[4436] = (layer0_outputs[2880]) & (layer0_outputs[8001]);
    assign layer1_outputs[4437] = (layer0_outputs[4636]) & (layer0_outputs[11706]);
    assign layer1_outputs[4438] = layer0_outputs[2318];
    assign layer1_outputs[4439] = layer0_outputs[10352];
    assign layer1_outputs[4440] = ~(layer0_outputs[1201]);
    assign layer1_outputs[4441] = (layer0_outputs[10157]) & (layer0_outputs[10601]);
    assign layer1_outputs[4442] = ~(layer0_outputs[2440]) | (layer0_outputs[3428]);
    assign layer1_outputs[4443] = ~(layer0_outputs[8394]) | (layer0_outputs[402]);
    assign layer1_outputs[4444] = ~(layer0_outputs[699]);
    assign layer1_outputs[4445] = ~(layer0_outputs[5453]);
    assign layer1_outputs[4446] = (layer0_outputs[7868]) | (layer0_outputs[4497]);
    assign layer1_outputs[4447] = layer0_outputs[9310];
    assign layer1_outputs[4448] = (layer0_outputs[8763]) & ~(layer0_outputs[1375]);
    assign layer1_outputs[4449] = (layer0_outputs[6011]) ^ (layer0_outputs[6214]);
    assign layer1_outputs[4450] = ~((layer0_outputs[2092]) | (layer0_outputs[3608]));
    assign layer1_outputs[4451] = ~(layer0_outputs[2266]);
    assign layer1_outputs[4452] = layer0_outputs[496];
    assign layer1_outputs[4453] = ~((layer0_outputs[11319]) | (layer0_outputs[4462]));
    assign layer1_outputs[4454] = ~((layer0_outputs[4988]) ^ (layer0_outputs[8802]));
    assign layer1_outputs[4455] = ~((layer0_outputs[1821]) | (layer0_outputs[5729]));
    assign layer1_outputs[4456] = ~(layer0_outputs[3687]);
    assign layer1_outputs[4457] = layer0_outputs[10292];
    assign layer1_outputs[4458] = ~(layer0_outputs[12012]) | (layer0_outputs[9905]);
    assign layer1_outputs[4459] = 1'b1;
    assign layer1_outputs[4460] = (layer0_outputs[4201]) | (layer0_outputs[3224]);
    assign layer1_outputs[4461] = ~(layer0_outputs[4419]) | (layer0_outputs[4985]);
    assign layer1_outputs[4462] = ~(layer0_outputs[3878]) | (layer0_outputs[11343]);
    assign layer1_outputs[4463] = layer0_outputs[6375];
    assign layer1_outputs[4464] = (layer0_outputs[2933]) & ~(layer0_outputs[11343]);
    assign layer1_outputs[4465] = ~((layer0_outputs[10741]) | (layer0_outputs[10515]));
    assign layer1_outputs[4466] = ~(layer0_outputs[2987]) | (layer0_outputs[7825]);
    assign layer1_outputs[4467] = ~(layer0_outputs[7380]);
    assign layer1_outputs[4468] = 1'b1;
    assign layer1_outputs[4469] = (layer0_outputs[1995]) & ~(layer0_outputs[4715]);
    assign layer1_outputs[4470] = ~(layer0_outputs[4422]) | (layer0_outputs[9748]);
    assign layer1_outputs[4471] = (layer0_outputs[438]) & (layer0_outputs[1284]);
    assign layer1_outputs[4472] = layer0_outputs[4196];
    assign layer1_outputs[4473] = (layer0_outputs[7037]) ^ (layer0_outputs[11534]);
    assign layer1_outputs[4474] = ~((layer0_outputs[4226]) ^ (layer0_outputs[131]));
    assign layer1_outputs[4475] = (layer0_outputs[7798]) | (layer0_outputs[6350]);
    assign layer1_outputs[4476] = ~(layer0_outputs[6751]) | (layer0_outputs[6424]);
    assign layer1_outputs[4477] = ~(layer0_outputs[11786]) | (layer0_outputs[9184]);
    assign layer1_outputs[4478] = (layer0_outputs[12654]) ^ (layer0_outputs[10171]);
    assign layer1_outputs[4479] = layer0_outputs[359];
    assign layer1_outputs[4480] = ~(layer0_outputs[12442]) | (layer0_outputs[6685]);
    assign layer1_outputs[4481] = (layer0_outputs[12231]) | (layer0_outputs[2013]);
    assign layer1_outputs[4482] = ~(layer0_outputs[12495]) | (layer0_outputs[12293]);
    assign layer1_outputs[4483] = ~(layer0_outputs[2932]) | (layer0_outputs[6204]);
    assign layer1_outputs[4484] = (layer0_outputs[2658]) & ~(layer0_outputs[9189]);
    assign layer1_outputs[4485] = layer0_outputs[11773];
    assign layer1_outputs[4486] = layer0_outputs[1694];
    assign layer1_outputs[4487] = (layer0_outputs[3196]) | (layer0_outputs[3515]);
    assign layer1_outputs[4488] = (layer0_outputs[9646]) & ~(layer0_outputs[10152]);
    assign layer1_outputs[4489] = layer0_outputs[6682];
    assign layer1_outputs[4490] = ~((layer0_outputs[3324]) ^ (layer0_outputs[3882]));
    assign layer1_outputs[4491] = layer0_outputs[3229];
    assign layer1_outputs[4492] = ~((layer0_outputs[9106]) ^ (layer0_outputs[7545]));
    assign layer1_outputs[4493] = (layer0_outputs[12462]) | (layer0_outputs[3578]);
    assign layer1_outputs[4494] = layer0_outputs[12171];
    assign layer1_outputs[4495] = (layer0_outputs[7642]) & (layer0_outputs[11789]);
    assign layer1_outputs[4496] = (layer0_outputs[9306]) & (layer0_outputs[1685]);
    assign layer1_outputs[4497] = ~((layer0_outputs[7644]) & (layer0_outputs[12039]));
    assign layer1_outputs[4498] = layer0_outputs[7657];
    assign layer1_outputs[4499] = ~((layer0_outputs[1712]) & (layer0_outputs[7353]));
    assign layer1_outputs[4500] = (layer0_outputs[1007]) | (layer0_outputs[3097]);
    assign layer1_outputs[4501] = ~((layer0_outputs[12142]) | (layer0_outputs[11968]));
    assign layer1_outputs[4502] = ~((layer0_outputs[8509]) & (layer0_outputs[557]));
    assign layer1_outputs[4503] = ~(layer0_outputs[3211]) | (layer0_outputs[7264]);
    assign layer1_outputs[4504] = (layer0_outputs[7296]) | (layer0_outputs[11279]);
    assign layer1_outputs[4505] = (layer0_outputs[12691]) & (layer0_outputs[6908]);
    assign layer1_outputs[4506] = ~(layer0_outputs[4159]);
    assign layer1_outputs[4507] = (layer0_outputs[10679]) & ~(layer0_outputs[686]);
    assign layer1_outputs[4508] = (layer0_outputs[8647]) & (layer0_outputs[9599]);
    assign layer1_outputs[4509] = (layer0_outputs[6280]) & (layer0_outputs[4498]);
    assign layer1_outputs[4510] = ~(layer0_outputs[6708]) | (layer0_outputs[5138]);
    assign layer1_outputs[4511] = ~((layer0_outputs[8598]) & (layer0_outputs[1952]));
    assign layer1_outputs[4512] = ~(layer0_outputs[8718]);
    assign layer1_outputs[4513] = (layer0_outputs[10807]) | (layer0_outputs[7242]);
    assign layer1_outputs[4514] = (layer0_outputs[7629]) | (layer0_outputs[2401]);
    assign layer1_outputs[4515] = (layer0_outputs[12622]) | (layer0_outputs[12108]);
    assign layer1_outputs[4516] = ~(layer0_outputs[5702]) | (layer0_outputs[12176]);
    assign layer1_outputs[4517] = (layer0_outputs[128]) ^ (layer0_outputs[6782]);
    assign layer1_outputs[4518] = (layer0_outputs[6136]) & (layer0_outputs[8772]);
    assign layer1_outputs[4519] = layer0_outputs[1057];
    assign layer1_outputs[4520] = ~((layer0_outputs[11800]) | (layer0_outputs[7925]));
    assign layer1_outputs[4521] = (layer0_outputs[841]) ^ (layer0_outputs[6439]);
    assign layer1_outputs[4522] = ~(layer0_outputs[3107]);
    assign layer1_outputs[4523] = (layer0_outputs[6096]) & (layer0_outputs[9322]);
    assign layer1_outputs[4524] = ~(layer0_outputs[1983]) | (layer0_outputs[11823]);
    assign layer1_outputs[4525] = ~((layer0_outputs[6355]) & (layer0_outputs[2288]));
    assign layer1_outputs[4526] = ~(layer0_outputs[8227]) | (layer0_outputs[8643]);
    assign layer1_outputs[4527] = layer0_outputs[2972];
    assign layer1_outputs[4528] = (layer0_outputs[6534]) & ~(layer0_outputs[5151]);
    assign layer1_outputs[4529] = ~(layer0_outputs[12296]);
    assign layer1_outputs[4530] = ~((layer0_outputs[9839]) & (layer0_outputs[7339]));
    assign layer1_outputs[4531] = (layer0_outputs[12353]) & ~(layer0_outputs[3959]);
    assign layer1_outputs[4532] = ~((layer0_outputs[8053]) & (layer0_outputs[1855]));
    assign layer1_outputs[4533] = layer0_outputs[5285];
    assign layer1_outputs[4534] = layer0_outputs[7886];
    assign layer1_outputs[4535] = ~(layer0_outputs[8631]) | (layer0_outputs[5369]);
    assign layer1_outputs[4536] = layer0_outputs[12449];
    assign layer1_outputs[4537] = layer0_outputs[9860];
    assign layer1_outputs[4538] = ~((layer0_outputs[145]) | (layer0_outputs[1865]));
    assign layer1_outputs[4539] = ~(layer0_outputs[761]) | (layer0_outputs[9736]);
    assign layer1_outputs[4540] = ~(layer0_outputs[9431]);
    assign layer1_outputs[4541] = ~(layer0_outputs[3336]);
    assign layer1_outputs[4542] = (layer0_outputs[10381]) ^ (layer0_outputs[3755]);
    assign layer1_outputs[4543] = layer0_outputs[5223];
    assign layer1_outputs[4544] = layer0_outputs[4264];
    assign layer1_outputs[4545] = ~(layer0_outputs[9928]);
    assign layer1_outputs[4546] = (layer0_outputs[3263]) & ~(layer0_outputs[2744]);
    assign layer1_outputs[4547] = ~((layer0_outputs[275]) & (layer0_outputs[12563]));
    assign layer1_outputs[4548] = ~(layer0_outputs[5674]);
    assign layer1_outputs[4549] = (layer0_outputs[5644]) & ~(layer0_outputs[1478]);
    assign layer1_outputs[4550] = (layer0_outputs[9586]) & (layer0_outputs[5563]);
    assign layer1_outputs[4551] = ~(layer0_outputs[10395]);
    assign layer1_outputs[4552] = 1'b1;
    assign layer1_outputs[4553] = ~((layer0_outputs[5295]) | (layer0_outputs[5900]));
    assign layer1_outputs[4554] = layer0_outputs[7322];
    assign layer1_outputs[4555] = ~((layer0_outputs[1517]) | (layer0_outputs[8836]));
    assign layer1_outputs[4556] = ~((layer0_outputs[9368]) | (layer0_outputs[5944]));
    assign layer1_outputs[4557] = (layer0_outputs[3678]) & (layer0_outputs[5752]);
    assign layer1_outputs[4558] = ~(layer0_outputs[4495]) | (layer0_outputs[3334]);
    assign layer1_outputs[4559] = (layer0_outputs[1791]) & ~(layer0_outputs[11855]);
    assign layer1_outputs[4560] = ~((layer0_outputs[2282]) | (layer0_outputs[12667]));
    assign layer1_outputs[4561] = ~((layer0_outputs[893]) & (layer0_outputs[7667]));
    assign layer1_outputs[4562] = ~(layer0_outputs[11730]) | (layer0_outputs[11915]);
    assign layer1_outputs[4563] = ~(layer0_outputs[8186]);
    assign layer1_outputs[4564] = layer0_outputs[1419];
    assign layer1_outputs[4565] = ~(layer0_outputs[12401]);
    assign layer1_outputs[4566] = ~(layer0_outputs[1488]) | (layer0_outputs[2451]);
    assign layer1_outputs[4567] = (layer0_outputs[244]) & ~(layer0_outputs[3873]);
    assign layer1_outputs[4568] = layer0_outputs[1741];
    assign layer1_outputs[4569] = layer0_outputs[291];
    assign layer1_outputs[4570] = ~((layer0_outputs[9051]) & (layer0_outputs[5534]));
    assign layer1_outputs[4571] = ~((layer0_outputs[1002]) & (layer0_outputs[3483]));
    assign layer1_outputs[4572] = layer0_outputs[5203];
    assign layer1_outputs[4573] = layer0_outputs[2848];
    assign layer1_outputs[4574] = (layer0_outputs[8365]) ^ (layer0_outputs[1624]);
    assign layer1_outputs[4575] = ~(layer0_outputs[6244]);
    assign layer1_outputs[4576] = (layer0_outputs[12516]) & ~(layer0_outputs[9168]);
    assign layer1_outputs[4577] = ~((layer0_outputs[10694]) | (layer0_outputs[2486]));
    assign layer1_outputs[4578] = ~(layer0_outputs[12043]) | (layer0_outputs[3183]);
    assign layer1_outputs[4579] = ~(layer0_outputs[6640]);
    assign layer1_outputs[4580] = ~((layer0_outputs[6837]) & (layer0_outputs[1778]));
    assign layer1_outputs[4581] = layer0_outputs[12187];
    assign layer1_outputs[4582] = ~(layer0_outputs[5496]) | (layer0_outputs[11304]);
    assign layer1_outputs[4583] = ~((layer0_outputs[694]) | (layer0_outputs[10535]));
    assign layer1_outputs[4584] = (layer0_outputs[1501]) ^ (layer0_outputs[117]);
    assign layer1_outputs[4585] = ~(layer0_outputs[9211]) | (layer0_outputs[324]);
    assign layer1_outputs[4586] = layer0_outputs[12642];
    assign layer1_outputs[4587] = layer0_outputs[7348];
    assign layer1_outputs[4588] = ~(layer0_outputs[4455]);
    assign layer1_outputs[4589] = layer0_outputs[1830];
    assign layer1_outputs[4590] = (layer0_outputs[9307]) & ~(layer0_outputs[9601]);
    assign layer1_outputs[4591] = ~(layer0_outputs[10534]) | (layer0_outputs[8724]);
    assign layer1_outputs[4592] = ~(layer0_outputs[459]);
    assign layer1_outputs[4593] = layer0_outputs[3604];
    assign layer1_outputs[4594] = ~(layer0_outputs[7288]) | (layer0_outputs[834]);
    assign layer1_outputs[4595] = ~(layer0_outputs[3287]);
    assign layer1_outputs[4596] = layer0_outputs[10315];
    assign layer1_outputs[4597] = (layer0_outputs[4486]) & ~(layer0_outputs[4020]);
    assign layer1_outputs[4598] = ~(layer0_outputs[5133]);
    assign layer1_outputs[4599] = ~(layer0_outputs[2006]) | (layer0_outputs[10555]);
    assign layer1_outputs[4600] = ~(layer0_outputs[3641]);
    assign layer1_outputs[4601] = ~(layer0_outputs[8120]);
    assign layer1_outputs[4602] = ~(layer0_outputs[5315]) | (layer0_outputs[2973]);
    assign layer1_outputs[4603] = layer0_outputs[8483];
    assign layer1_outputs[4604] = ~(layer0_outputs[2834]) | (layer0_outputs[2420]);
    assign layer1_outputs[4605] = ~(layer0_outputs[6208]);
    assign layer1_outputs[4606] = (layer0_outputs[5118]) & (layer0_outputs[10971]);
    assign layer1_outputs[4607] = layer0_outputs[12415];
    assign layer1_outputs[4608] = (layer0_outputs[7929]) | (layer0_outputs[11244]);
    assign layer1_outputs[4609] = layer0_outputs[4433];
    assign layer1_outputs[4610] = (layer0_outputs[2022]) & (layer0_outputs[6541]);
    assign layer1_outputs[4611] = (layer0_outputs[7475]) & ~(layer0_outputs[5926]);
    assign layer1_outputs[4612] = (layer0_outputs[6458]) ^ (layer0_outputs[6672]);
    assign layer1_outputs[4613] = (layer0_outputs[1560]) & ~(layer0_outputs[1796]);
    assign layer1_outputs[4614] = ~(layer0_outputs[5213]) | (layer0_outputs[423]);
    assign layer1_outputs[4615] = (layer0_outputs[5688]) & (layer0_outputs[9448]);
    assign layer1_outputs[4616] = layer0_outputs[12580];
    assign layer1_outputs[4617] = ~(layer0_outputs[591]) | (layer0_outputs[6251]);
    assign layer1_outputs[4618] = layer0_outputs[10345];
    assign layer1_outputs[4619] = (layer0_outputs[1132]) & ~(layer0_outputs[3888]);
    assign layer1_outputs[4620] = ~(layer0_outputs[9912]);
    assign layer1_outputs[4621] = ~(layer0_outputs[4524]) | (layer0_outputs[11054]);
    assign layer1_outputs[4622] = ~(layer0_outputs[9070]) | (layer0_outputs[5074]);
    assign layer1_outputs[4623] = ~(layer0_outputs[7187]);
    assign layer1_outputs[4624] = ~((layer0_outputs[3450]) | (layer0_outputs[2653]));
    assign layer1_outputs[4625] = ~(layer0_outputs[7294]) | (layer0_outputs[9253]);
    assign layer1_outputs[4626] = 1'b1;
    assign layer1_outputs[4627] = ~(layer0_outputs[730]);
    assign layer1_outputs[4628] = (layer0_outputs[6886]) & ~(layer0_outputs[9321]);
    assign layer1_outputs[4629] = layer0_outputs[1825];
    assign layer1_outputs[4630] = ~(layer0_outputs[2650]);
    assign layer1_outputs[4631] = ~((layer0_outputs[3584]) & (layer0_outputs[912]));
    assign layer1_outputs[4632] = ~(layer0_outputs[8743]);
    assign layer1_outputs[4633] = (layer0_outputs[1293]) & (layer0_outputs[4373]);
    assign layer1_outputs[4634] = ~((layer0_outputs[209]) | (layer0_outputs[8988]));
    assign layer1_outputs[4635] = ~(layer0_outputs[12060]) | (layer0_outputs[2255]);
    assign layer1_outputs[4636] = ~((layer0_outputs[654]) ^ (layer0_outputs[8583]));
    assign layer1_outputs[4637] = (layer0_outputs[10643]) | (layer0_outputs[715]);
    assign layer1_outputs[4638] = ~(layer0_outputs[630]) | (layer0_outputs[4995]);
    assign layer1_outputs[4639] = ~((layer0_outputs[10704]) & (layer0_outputs[3488]));
    assign layer1_outputs[4640] = ~(layer0_outputs[9344]);
    assign layer1_outputs[4641] = (layer0_outputs[2491]) & ~(layer0_outputs[9059]);
    assign layer1_outputs[4642] = ~((layer0_outputs[2970]) ^ (layer0_outputs[7999]));
    assign layer1_outputs[4643] = 1'b1;
    assign layer1_outputs[4644] = layer0_outputs[294];
    assign layer1_outputs[4645] = ~((layer0_outputs[3819]) & (layer0_outputs[11550]));
    assign layer1_outputs[4646] = ~(layer0_outputs[5033]) | (layer0_outputs[222]);
    assign layer1_outputs[4647] = layer0_outputs[10745];
    assign layer1_outputs[4648] = ~(layer0_outputs[5784]);
    assign layer1_outputs[4649] = (layer0_outputs[6189]) & (layer0_outputs[6338]);
    assign layer1_outputs[4650] = ~(layer0_outputs[4855]);
    assign layer1_outputs[4651] = (layer0_outputs[9765]) & ~(layer0_outputs[3946]);
    assign layer1_outputs[4652] = 1'b0;
    assign layer1_outputs[4653] = layer0_outputs[16];
    assign layer1_outputs[4654] = ~(layer0_outputs[4175]);
    assign layer1_outputs[4655] = layer0_outputs[5202];
    assign layer1_outputs[4656] = layer0_outputs[7003];
    assign layer1_outputs[4657] = ~(layer0_outputs[8176]);
    assign layer1_outputs[4658] = ~((layer0_outputs[3222]) & (layer0_outputs[5318]));
    assign layer1_outputs[4659] = layer0_outputs[3363];
    assign layer1_outputs[4660] = 1'b0;
    assign layer1_outputs[4661] = (layer0_outputs[6371]) & ~(layer0_outputs[11281]);
    assign layer1_outputs[4662] = (layer0_outputs[772]) | (layer0_outputs[5820]);
    assign layer1_outputs[4663] = ~(layer0_outputs[6010]);
    assign layer1_outputs[4664] = ~(layer0_outputs[11103]);
    assign layer1_outputs[4665] = ~(layer0_outputs[6928]);
    assign layer1_outputs[4666] = (layer0_outputs[3168]) ^ (layer0_outputs[8362]);
    assign layer1_outputs[4667] = layer0_outputs[170];
    assign layer1_outputs[4668] = ~(layer0_outputs[10700]);
    assign layer1_outputs[4669] = (layer0_outputs[11049]) & ~(layer0_outputs[2565]);
    assign layer1_outputs[4670] = ~(layer0_outputs[4882]);
    assign layer1_outputs[4671] = (layer0_outputs[5162]) & ~(layer0_outputs[723]);
    assign layer1_outputs[4672] = ~(layer0_outputs[9540]) | (layer0_outputs[7383]);
    assign layer1_outputs[4673] = (layer0_outputs[427]) & ~(layer0_outputs[6618]);
    assign layer1_outputs[4674] = ~(layer0_outputs[2045]);
    assign layer1_outputs[4675] = (layer0_outputs[2059]) ^ (layer0_outputs[12363]);
    assign layer1_outputs[4676] = (layer0_outputs[7316]) ^ (layer0_outputs[9051]);
    assign layer1_outputs[4677] = ~((layer0_outputs[7827]) | (layer0_outputs[2700]));
    assign layer1_outputs[4678] = ~(layer0_outputs[6681]) | (layer0_outputs[1279]);
    assign layer1_outputs[4679] = ~(layer0_outputs[11214]);
    assign layer1_outputs[4680] = ~((layer0_outputs[4086]) & (layer0_outputs[8512]));
    assign layer1_outputs[4681] = (layer0_outputs[8081]) & ~(layer0_outputs[1706]);
    assign layer1_outputs[4682] = (layer0_outputs[8315]) & (layer0_outputs[3464]);
    assign layer1_outputs[4683] = ~(layer0_outputs[11693]) | (layer0_outputs[2233]);
    assign layer1_outputs[4684] = layer0_outputs[8060];
    assign layer1_outputs[4685] = layer0_outputs[2535];
    assign layer1_outputs[4686] = layer0_outputs[5940];
    assign layer1_outputs[4687] = ~(layer0_outputs[8276]);
    assign layer1_outputs[4688] = ~(layer0_outputs[7399]);
    assign layer1_outputs[4689] = ~(layer0_outputs[6874]);
    assign layer1_outputs[4690] = 1'b0;
    assign layer1_outputs[4691] = ~(layer0_outputs[693]);
    assign layer1_outputs[4692] = (layer0_outputs[10518]) & ~(layer0_outputs[5281]);
    assign layer1_outputs[4693] = layer0_outputs[6168];
    assign layer1_outputs[4694] = (layer0_outputs[2351]) & (layer0_outputs[4979]);
    assign layer1_outputs[4695] = (layer0_outputs[9040]) ^ (layer0_outputs[12798]);
    assign layer1_outputs[4696] = (layer0_outputs[6077]) & ~(layer0_outputs[12300]);
    assign layer1_outputs[4697] = (layer0_outputs[24]) & ~(layer0_outputs[1260]);
    assign layer1_outputs[4698] = layer0_outputs[12419];
    assign layer1_outputs[4699] = 1'b1;
    assign layer1_outputs[4700] = ~(layer0_outputs[10916]);
    assign layer1_outputs[4701] = layer0_outputs[8080];
    assign layer1_outputs[4702] = layer0_outputs[971];
    assign layer1_outputs[4703] = ~(layer0_outputs[3842]) | (layer0_outputs[8698]);
    assign layer1_outputs[4704] = ~((layer0_outputs[9964]) ^ (layer0_outputs[10172]));
    assign layer1_outputs[4705] = (layer0_outputs[1996]) ^ (layer0_outputs[4958]);
    assign layer1_outputs[4706] = ~(layer0_outputs[11652]);
    assign layer1_outputs[4707] = ~((layer0_outputs[4165]) | (layer0_outputs[9791]));
    assign layer1_outputs[4708] = layer0_outputs[6485];
    assign layer1_outputs[4709] = ~((layer0_outputs[2905]) ^ (layer0_outputs[2505]));
    assign layer1_outputs[4710] = ~(layer0_outputs[6551]);
    assign layer1_outputs[4711] = layer0_outputs[6114];
    assign layer1_outputs[4712] = ~(layer0_outputs[8123]);
    assign layer1_outputs[4713] = ~((layer0_outputs[3964]) | (layer0_outputs[11990]));
    assign layer1_outputs[4714] = ~(layer0_outputs[4576]);
    assign layer1_outputs[4715] = ~(layer0_outputs[7646]);
    assign layer1_outputs[4716] = ~((layer0_outputs[8837]) ^ (layer0_outputs[2514]));
    assign layer1_outputs[4717] = (layer0_outputs[11053]) & (layer0_outputs[9445]);
    assign layer1_outputs[4718] = ~((layer0_outputs[1191]) ^ (layer0_outputs[65]));
    assign layer1_outputs[4719] = (layer0_outputs[3038]) & ~(layer0_outputs[10027]);
    assign layer1_outputs[4720] = layer0_outputs[5123];
    assign layer1_outputs[4721] = ~((layer0_outputs[8970]) | (layer0_outputs[6273]));
    assign layer1_outputs[4722] = ~((layer0_outputs[11955]) & (layer0_outputs[12128]));
    assign layer1_outputs[4723] = 1'b0;
    assign layer1_outputs[4724] = (layer0_outputs[6731]) & ~(layer0_outputs[124]);
    assign layer1_outputs[4725] = layer0_outputs[10721];
    assign layer1_outputs[4726] = ~((layer0_outputs[11086]) & (layer0_outputs[3253]));
    assign layer1_outputs[4727] = (layer0_outputs[6307]) | (layer0_outputs[8808]);
    assign layer1_outputs[4728] = ~(layer0_outputs[7219]) | (layer0_outputs[8747]);
    assign layer1_outputs[4729] = layer0_outputs[9455];
    assign layer1_outputs[4730] = layer0_outputs[2800];
    assign layer1_outputs[4731] = layer0_outputs[5870];
    assign layer1_outputs[4732] = (layer0_outputs[11440]) & ~(layer0_outputs[11974]);
    assign layer1_outputs[4733] = (layer0_outputs[12736]) & ~(layer0_outputs[4520]);
    assign layer1_outputs[4734] = ~((layer0_outputs[5488]) ^ (layer0_outputs[4992]));
    assign layer1_outputs[4735] = ~((layer0_outputs[5386]) & (layer0_outputs[7497]));
    assign layer1_outputs[4736] = ~(layer0_outputs[2511]) | (layer0_outputs[1585]);
    assign layer1_outputs[4737] = ~((layer0_outputs[1953]) ^ (layer0_outputs[4739]));
    assign layer1_outputs[4738] = (layer0_outputs[7723]) & ~(layer0_outputs[11357]);
    assign layer1_outputs[4739] = layer0_outputs[1908];
    assign layer1_outputs[4740] = ~(layer0_outputs[11933]);
    assign layer1_outputs[4741] = ~(layer0_outputs[10263]) | (layer0_outputs[11093]);
    assign layer1_outputs[4742] = ~(layer0_outputs[3855]) | (layer0_outputs[5479]);
    assign layer1_outputs[4743] = layer0_outputs[6988];
    assign layer1_outputs[4744] = ~(layer0_outputs[3787]) | (layer0_outputs[1515]);
    assign layer1_outputs[4745] = ~(layer0_outputs[9837]);
    assign layer1_outputs[4746] = (layer0_outputs[5282]) & (layer0_outputs[8025]);
    assign layer1_outputs[4747] = layer0_outputs[11383];
    assign layer1_outputs[4748] = layer0_outputs[11194];
    assign layer1_outputs[4749] = layer0_outputs[10887];
    assign layer1_outputs[4750] = ~(layer0_outputs[4909]);
    assign layer1_outputs[4751] = ~(layer0_outputs[2358]);
    assign layer1_outputs[4752] = (layer0_outputs[6069]) & (layer0_outputs[5851]);
    assign layer1_outputs[4753] = ~((layer0_outputs[5415]) & (layer0_outputs[2801]));
    assign layer1_outputs[4754] = (layer0_outputs[3962]) & ~(layer0_outputs[2814]);
    assign layer1_outputs[4755] = (layer0_outputs[100]) | (layer0_outputs[8572]);
    assign layer1_outputs[4756] = (layer0_outputs[8031]) & ~(layer0_outputs[9216]);
    assign layer1_outputs[4757] = (layer0_outputs[34]) ^ (layer0_outputs[6353]);
    assign layer1_outputs[4758] = ~((layer0_outputs[4205]) ^ (layer0_outputs[1373]));
    assign layer1_outputs[4759] = layer0_outputs[7];
    assign layer1_outputs[4760] = layer0_outputs[6212];
    assign layer1_outputs[4761] = (layer0_outputs[4359]) & ~(layer0_outputs[1450]);
    assign layer1_outputs[4762] = layer0_outputs[11382];
    assign layer1_outputs[4763] = ~(layer0_outputs[7474]);
    assign layer1_outputs[4764] = ~(layer0_outputs[2442]);
    assign layer1_outputs[4765] = (layer0_outputs[5158]) | (layer0_outputs[3042]);
    assign layer1_outputs[4766] = ~(layer0_outputs[2476]) | (layer0_outputs[11572]);
    assign layer1_outputs[4767] = (layer0_outputs[873]) | (layer0_outputs[10506]);
    assign layer1_outputs[4768] = ~(layer0_outputs[8906]);
    assign layer1_outputs[4769] = (layer0_outputs[1185]) ^ (layer0_outputs[4585]);
    assign layer1_outputs[4770] = layer0_outputs[12281];
    assign layer1_outputs[4771] = (layer0_outputs[1871]) | (layer0_outputs[7073]);
    assign layer1_outputs[4772] = ~(layer0_outputs[5409]) | (layer0_outputs[7009]);
    assign layer1_outputs[4773] = (layer0_outputs[7342]) & (layer0_outputs[12464]);
    assign layer1_outputs[4774] = (layer0_outputs[4362]) | (layer0_outputs[4582]);
    assign layer1_outputs[4775] = ~(layer0_outputs[5329]) | (layer0_outputs[6341]);
    assign layer1_outputs[4776] = layer0_outputs[271];
    assign layer1_outputs[4777] = (layer0_outputs[3281]) ^ (layer0_outputs[11389]);
    assign layer1_outputs[4778] = layer0_outputs[8486];
    assign layer1_outputs[4779] = ~(layer0_outputs[11313]);
    assign layer1_outputs[4780] = ~(layer0_outputs[5287]);
    assign layer1_outputs[4781] = (layer0_outputs[8594]) & ~(layer0_outputs[3542]);
    assign layer1_outputs[4782] = layer0_outputs[852];
    assign layer1_outputs[4783] = layer0_outputs[12547];
    assign layer1_outputs[4784] = layer0_outputs[10585];
    assign layer1_outputs[4785] = ~(layer0_outputs[8969]);
    assign layer1_outputs[4786] = ~((layer0_outputs[11016]) | (layer0_outputs[2581]));
    assign layer1_outputs[4787] = (layer0_outputs[169]) ^ (layer0_outputs[11478]);
    assign layer1_outputs[4788] = ~(layer0_outputs[10933]);
    assign layer1_outputs[4789] = (layer0_outputs[3917]) & (layer0_outputs[4125]);
    assign layer1_outputs[4790] = layer0_outputs[11776];
    assign layer1_outputs[4791] = ~(layer0_outputs[11970]) | (layer0_outputs[3593]);
    assign layer1_outputs[4792] = (layer0_outputs[6620]) & ~(layer0_outputs[12774]);
    assign layer1_outputs[4793] = ~(layer0_outputs[361]);
    assign layer1_outputs[4794] = layer0_outputs[11449];
    assign layer1_outputs[4795] = 1'b1;
    assign layer1_outputs[4796] = ~(layer0_outputs[236]) | (layer0_outputs[4616]);
    assign layer1_outputs[4797] = layer0_outputs[9623];
    assign layer1_outputs[4798] = (layer0_outputs[7485]) & ~(layer0_outputs[4515]);
    assign layer1_outputs[4799] = ~(layer0_outputs[11756]);
    assign layer1_outputs[4800] = (layer0_outputs[3407]) & ~(layer0_outputs[2038]);
    assign layer1_outputs[4801] = ~((layer0_outputs[9418]) | (layer0_outputs[1015]));
    assign layer1_outputs[4802] = layer0_outputs[2150];
    assign layer1_outputs[4803] = layer0_outputs[9880];
    assign layer1_outputs[4804] = ~((layer0_outputs[576]) & (layer0_outputs[9548]));
    assign layer1_outputs[4805] = layer0_outputs[7208];
    assign layer1_outputs[4806] = (layer0_outputs[5002]) & (layer0_outputs[5652]);
    assign layer1_outputs[4807] = ~(layer0_outputs[4778]);
    assign layer1_outputs[4808] = ~((layer0_outputs[6491]) ^ (layer0_outputs[10939]));
    assign layer1_outputs[4809] = (layer0_outputs[2419]) & ~(layer0_outputs[587]);
    assign layer1_outputs[4810] = (layer0_outputs[12661]) | (layer0_outputs[2121]);
    assign layer1_outputs[4811] = (layer0_outputs[1647]) & ~(layer0_outputs[11161]);
    assign layer1_outputs[4812] = (layer0_outputs[12057]) ^ (layer0_outputs[9970]);
    assign layer1_outputs[4813] = ~(layer0_outputs[6254]);
    assign layer1_outputs[4814] = (layer0_outputs[8902]) ^ (layer0_outputs[1727]);
    assign layer1_outputs[4815] = (layer0_outputs[6402]) & (layer0_outputs[90]);
    assign layer1_outputs[4816] = ~((layer0_outputs[7771]) & (layer0_outputs[3559]));
    assign layer1_outputs[4817] = ~(layer0_outputs[9688]);
    assign layer1_outputs[4818] = (layer0_outputs[6610]) & ~(layer0_outputs[9439]);
    assign layer1_outputs[4819] = layer0_outputs[8005];
    assign layer1_outputs[4820] = (layer0_outputs[1707]) & ~(layer0_outputs[12298]);
    assign layer1_outputs[4821] = layer0_outputs[166];
    assign layer1_outputs[4822] = (layer0_outputs[1458]) & ~(layer0_outputs[279]);
    assign layer1_outputs[4823] = (layer0_outputs[10193]) & ~(layer0_outputs[1669]);
    assign layer1_outputs[4824] = (layer0_outputs[4706]) & ~(layer0_outputs[2135]);
    assign layer1_outputs[4825] = ~((layer0_outputs[9462]) | (layer0_outputs[72]));
    assign layer1_outputs[4826] = ~(layer0_outputs[4452]);
    assign layer1_outputs[4827] = (layer0_outputs[10732]) | (layer0_outputs[4275]);
    assign layer1_outputs[4828] = ~((layer0_outputs[1177]) | (layer0_outputs[814]));
    assign layer1_outputs[4829] = layer0_outputs[1124];
    assign layer1_outputs[4830] = ~((layer0_outputs[2962]) | (layer0_outputs[9069]));
    assign layer1_outputs[4831] = layer0_outputs[6122];
    assign layer1_outputs[4832] = ~(layer0_outputs[7390]);
    assign layer1_outputs[4833] = (layer0_outputs[3002]) | (layer0_outputs[12549]);
    assign layer1_outputs[4834] = (layer0_outputs[12596]) & (layer0_outputs[12184]);
    assign layer1_outputs[4835] = (layer0_outputs[2402]) & ~(layer0_outputs[8759]);
    assign layer1_outputs[4836] = (layer0_outputs[8078]) & ~(layer0_outputs[9775]);
    assign layer1_outputs[4837] = ~(layer0_outputs[614]) | (layer0_outputs[7986]);
    assign layer1_outputs[4838] = ~((layer0_outputs[11059]) | (layer0_outputs[6914]));
    assign layer1_outputs[4839] = (layer0_outputs[12166]) & ~(layer0_outputs[718]);
    assign layer1_outputs[4840] = (layer0_outputs[3159]) & ~(layer0_outputs[6223]);
    assign layer1_outputs[4841] = ~(layer0_outputs[491]);
    assign layer1_outputs[4842] = layer0_outputs[9648];
    assign layer1_outputs[4843] = (layer0_outputs[9664]) | (layer0_outputs[8423]);
    assign layer1_outputs[4844] = ~(layer0_outputs[6311]);
    assign layer1_outputs[4845] = (layer0_outputs[5190]) ^ (layer0_outputs[768]);
    assign layer1_outputs[4846] = ~((layer0_outputs[10336]) & (layer0_outputs[9539]));
    assign layer1_outputs[4847] = layer0_outputs[639];
    assign layer1_outputs[4848] = (layer0_outputs[5577]) | (layer0_outputs[6899]);
    assign layer1_outputs[4849] = ~((layer0_outputs[2503]) & (layer0_outputs[9772]));
    assign layer1_outputs[4850] = (layer0_outputs[10185]) & ~(layer0_outputs[10903]);
    assign layer1_outputs[4851] = (layer0_outputs[471]) & ~(layer0_outputs[11819]);
    assign layer1_outputs[4852] = ~((layer0_outputs[6870]) ^ (layer0_outputs[9257]));
    assign layer1_outputs[4853] = 1'b0;
    assign layer1_outputs[4854] = layer0_outputs[11727];
    assign layer1_outputs[4855] = 1'b0;
    assign layer1_outputs[4856] = ~(layer0_outputs[9852]);
    assign layer1_outputs[4857] = (layer0_outputs[6598]) & (layer0_outputs[11401]);
    assign layer1_outputs[4858] = ~(layer0_outputs[10356]) | (layer0_outputs[4107]);
    assign layer1_outputs[4859] = ~(layer0_outputs[9281]) | (layer0_outputs[10410]);
    assign layer1_outputs[4860] = ~((layer0_outputs[12635]) | (layer0_outputs[6250]));
    assign layer1_outputs[4861] = ~((layer0_outputs[3468]) | (layer0_outputs[11135]));
    assign layer1_outputs[4862] = ~(layer0_outputs[10075]) | (layer0_outputs[7845]);
    assign layer1_outputs[4863] = ~(layer0_outputs[4631]) | (layer0_outputs[9012]);
    assign layer1_outputs[4864] = (layer0_outputs[1101]) & (layer0_outputs[12668]);
    assign layer1_outputs[4865] = layer0_outputs[9653];
    assign layer1_outputs[4866] = ~(layer0_outputs[5907]);
    assign layer1_outputs[4867] = layer0_outputs[6762];
    assign layer1_outputs[4868] = ~(layer0_outputs[11923]);
    assign layer1_outputs[4869] = ~(layer0_outputs[1052]);
    assign layer1_outputs[4870] = ~(layer0_outputs[261]) | (layer0_outputs[29]);
    assign layer1_outputs[4871] = 1'b0;
    assign layer1_outputs[4872] = ~((layer0_outputs[6030]) ^ (layer0_outputs[1441]));
    assign layer1_outputs[4873] = ~((layer0_outputs[2031]) & (layer0_outputs[9179]));
    assign layer1_outputs[4874] = (layer0_outputs[9519]) ^ (layer0_outputs[5376]);
    assign layer1_outputs[4875] = ~(layer0_outputs[11136]);
    assign layer1_outputs[4876] = layer0_outputs[9804];
    assign layer1_outputs[4877] = layer0_outputs[8555];
    assign layer1_outputs[4878] = ~((layer0_outputs[5276]) | (layer0_outputs[11646]));
    assign layer1_outputs[4879] = (layer0_outputs[3812]) & (layer0_outputs[12522]);
    assign layer1_outputs[4880] = (layer0_outputs[5078]) & ~(layer0_outputs[3480]);
    assign layer1_outputs[4881] = layer0_outputs[12132];
    assign layer1_outputs[4882] = (layer0_outputs[3311]) | (layer0_outputs[4531]);
    assign layer1_outputs[4883] = ~((layer0_outputs[3221]) | (layer0_outputs[11338]));
    assign layer1_outputs[4884] = ~(layer0_outputs[9188]) | (layer0_outputs[9117]);
    assign layer1_outputs[4885] = (layer0_outputs[11081]) & ~(layer0_outputs[7174]);
    assign layer1_outputs[4886] = ~(layer0_outputs[259]);
    assign layer1_outputs[4887] = ~((layer0_outputs[7603]) | (layer0_outputs[1142]));
    assign layer1_outputs[4888] = (layer0_outputs[916]) ^ (layer0_outputs[8915]);
    assign layer1_outputs[4889] = ~(layer0_outputs[10189]);
    assign layer1_outputs[4890] = ~(layer0_outputs[7156]);
    assign layer1_outputs[4891] = (layer0_outputs[11070]) & ~(layer0_outputs[10116]);
    assign layer1_outputs[4892] = ~(layer0_outputs[1908]) | (layer0_outputs[3474]);
    assign layer1_outputs[4893] = ~((layer0_outputs[2192]) & (layer0_outputs[10682]));
    assign layer1_outputs[4894] = layer0_outputs[11758];
    assign layer1_outputs[4895] = (layer0_outputs[12358]) & (layer0_outputs[3209]);
    assign layer1_outputs[4896] = ~(layer0_outputs[5085]);
    assign layer1_outputs[4897] = (layer0_outputs[9024]) & ~(layer0_outputs[1896]);
    assign layer1_outputs[4898] = ~((layer0_outputs[9199]) | (layer0_outputs[1955]));
    assign layer1_outputs[4899] = (layer0_outputs[3525]) | (layer0_outputs[4781]);
    assign layer1_outputs[4900] = (layer0_outputs[6178]) & ~(layer0_outputs[7667]);
    assign layer1_outputs[4901] = ~(layer0_outputs[108]);
    assign layer1_outputs[4902] = ~((layer0_outputs[5696]) | (layer0_outputs[12465]));
    assign layer1_outputs[4903] = ~(layer0_outputs[9826]);
    assign layer1_outputs[4904] = ~(layer0_outputs[9741]);
    assign layer1_outputs[4905] = ~((layer0_outputs[7185]) | (layer0_outputs[5529]));
    assign layer1_outputs[4906] = ~(layer0_outputs[7087]);
    assign layer1_outputs[4907] = layer0_outputs[6021];
    assign layer1_outputs[4908] = (layer0_outputs[1447]) & ~(layer0_outputs[2966]);
    assign layer1_outputs[4909] = ~((layer0_outputs[6474]) | (layer0_outputs[3344]));
    assign layer1_outputs[4910] = ~(layer0_outputs[8387]);
    assign layer1_outputs[4911] = ~((layer0_outputs[11866]) ^ (layer0_outputs[11160]));
    assign layer1_outputs[4912] = ~(layer0_outputs[7123]);
    assign layer1_outputs[4913] = (layer0_outputs[1690]) & (layer0_outputs[7476]);
    assign layer1_outputs[4914] = ~(layer0_outputs[4167]) | (layer0_outputs[8483]);
    assign layer1_outputs[4915] = ~(layer0_outputs[10070]) | (layer0_outputs[10692]);
    assign layer1_outputs[4916] = ~(layer0_outputs[4840]);
    assign layer1_outputs[4917] = ~((layer0_outputs[6446]) ^ (layer0_outputs[2249]));
    assign layer1_outputs[4918] = layer0_outputs[1205];
    assign layer1_outputs[4919] = 1'b0;
    assign layer1_outputs[4920] = (layer0_outputs[5308]) | (layer0_outputs[3094]);
    assign layer1_outputs[4921] = layer0_outputs[711];
    assign layer1_outputs[4922] = (layer0_outputs[12472]) | (layer0_outputs[9757]);
    assign layer1_outputs[4923] = ~(layer0_outputs[2212]);
    assign layer1_outputs[4924] = ~((layer0_outputs[1762]) | (layer0_outputs[7406]));
    assign layer1_outputs[4925] = (layer0_outputs[532]) & ~(layer0_outputs[1237]);
    assign layer1_outputs[4926] = (layer0_outputs[6473]) & ~(layer0_outputs[5868]);
    assign layer1_outputs[4927] = ~(layer0_outputs[1664]) | (layer0_outputs[10047]);
    assign layer1_outputs[4928] = ~(layer0_outputs[10989]);
    assign layer1_outputs[4929] = layer0_outputs[7586];
    assign layer1_outputs[4930] = ~((layer0_outputs[2946]) & (layer0_outputs[2859]));
    assign layer1_outputs[4931] = (layer0_outputs[3952]) | (layer0_outputs[11360]);
    assign layer1_outputs[4932] = ~(layer0_outputs[4313]);
    assign layer1_outputs[4933] = ~(layer0_outputs[11149]) | (layer0_outputs[8676]);
    assign layer1_outputs[4934] = (layer0_outputs[3984]) & (layer0_outputs[12652]);
    assign layer1_outputs[4935] = (layer0_outputs[6794]) ^ (layer0_outputs[5205]);
    assign layer1_outputs[4936] = ~(layer0_outputs[5057]);
    assign layer1_outputs[4937] = ~(layer0_outputs[3215]) | (layer0_outputs[7249]);
    assign layer1_outputs[4938] = (layer0_outputs[5049]) & ~(layer0_outputs[11925]);
    assign layer1_outputs[4939] = layer0_outputs[1400];
    assign layer1_outputs[4940] = (layer0_outputs[10271]) ^ (layer0_outputs[11616]);
    assign layer1_outputs[4941] = (layer0_outputs[5823]) ^ (layer0_outputs[8005]);
    assign layer1_outputs[4942] = (layer0_outputs[11984]) & ~(layer0_outputs[1407]);
    assign layer1_outputs[4943] = ~(layer0_outputs[1609]);
    assign layer1_outputs[4944] = ~(layer0_outputs[4011]) | (layer0_outputs[6700]);
    assign layer1_outputs[4945] = ~(layer0_outputs[5311]);
    assign layer1_outputs[4946] = (layer0_outputs[3466]) & (layer0_outputs[4145]);
    assign layer1_outputs[4947] = (layer0_outputs[10841]) & ~(layer0_outputs[8269]);
    assign layer1_outputs[4948] = (layer0_outputs[1633]) & ~(layer0_outputs[9801]);
    assign layer1_outputs[4949] = (layer0_outputs[2983]) & (layer0_outputs[121]);
    assign layer1_outputs[4950] = (layer0_outputs[7358]) & ~(layer0_outputs[9055]);
    assign layer1_outputs[4951] = (layer0_outputs[9498]) & ~(layer0_outputs[7804]);
    assign layer1_outputs[4952] = (layer0_outputs[3201]) & ~(layer0_outputs[3001]);
    assign layer1_outputs[4953] = ~(layer0_outputs[826]);
    assign layer1_outputs[4954] = layer0_outputs[10582];
    assign layer1_outputs[4955] = layer0_outputs[5251];
    assign layer1_outputs[4956] = layer0_outputs[11384];
    assign layer1_outputs[4957] = (layer0_outputs[3983]) | (layer0_outputs[7967]);
    assign layer1_outputs[4958] = (layer0_outputs[10949]) & (layer0_outputs[10547]);
    assign layer1_outputs[4959] = (layer0_outputs[1103]) & ~(layer0_outputs[5692]);
    assign layer1_outputs[4960] = layer0_outputs[1127];
    assign layer1_outputs[4961] = ~(layer0_outputs[10500]);
    assign layer1_outputs[4962] = ~((layer0_outputs[2892]) | (layer0_outputs[8430]));
    assign layer1_outputs[4963] = layer0_outputs[2404];
    assign layer1_outputs[4964] = ~((layer0_outputs[11266]) & (layer0_outputs[927]));
    assign layer1_outputs[4965] = ~(layer0_outputs[3272]);
    assign layer1_outputs[4966] = ~(layer0_outputs[7134]) | (layer0_outputs[3372]);
    assign layer1_outputs[4967] = (layer0_outputs[11636]) ^ (layer0_outputs[4301]);
    assign layer1_outputs[4968] = layer0_outputs[11267];
    assign layer1_outputs[4969] = ~(layer0_outputs[5999]) | (layer0_outputs[11924]);
    assign layer1_outputs[4970] = ~(layer0_outputs[11837]);
    assign layer1_outputs[4971] = (layer0_outputs[6482]) & ~(layer0_outputs[12270]);
    assign layer1_outputs[4972] = (layer0_outputs[3496]) & ~(layer0_outputs[12212]);
    assign layer1_outputs[4973] = ~(layer0_outputs[10478]);
    assign layer1_outputs[4974] = ~((layer0_outputs[1783]) | (layer0_outputs[11450]));
    assign layer1_outputs[4975] = (layer0_outputs[2682]) & ~(layer0_outputs[3765]);
    assign layer1_outputs[4976] = ~(layer0_outputs[5158]) | (layer0_outputs[2583]);
    assign layer1_outputs[4977] = layer0_outputs[10214];
    assign layer1_outputs[4978] = (layer0_outputs[12240]) | (layer0_outputs[6535]);
    assign layer1_outputs[4979] = layer0_outputs[11667];
    assign layer1_outputs[4980] = (layer0_outputs[9024]) & ~(layer0_outputs[4749]);
    assign layer1_outputs[4981] = ~((layer0_outputs[3788]) ^ (layer0_outputs[690]));
    assign layer1_outputs[4982] = (layer0_outputs[11180]) & (layer0_outputs[5483]);
    assign layer1_outputs[4983] = (layer0_outputs[9129]) & ~(layer0_outputs[1296]);
    assign layer1_outputs[4984] = ~((layer0_outputs[3822]) ^ (layer0_outputs[1494]));
    assign layer1_outputs[4985] = ~((layer0_outputs[12195]) & (layer0_outputs[10855]));
    assign layer1_outputs[4986] = (layer0_outputs[968]) & (layer0_outputs[10747]);
    assign layer1_outputs[4987] = layer0_outputs[12679];
    assign layer1_outputs[4988] = ~(layer0_outputs[10300]) | (layer0_outputs[1022]);
    assign layer1_outputs[4989] = ~(layer0_outputs[2927]);
    assign layer1_outputs[4990] = (layer0_outputs[7808]) | (layer0_outputs[11073]);
    assign layer1_outputs[4991] = layer0_outputs[7431];
    assign layer1_outputs[4992] = ~(layer0_outputs[6044]);
    assign layer1_outputs[4993] = (layer0_outputs[5548]) | (layer0_outputs[6779]);
    assign layer1_outputs[4994] = ~(layer0_outputs[5721]);
    assign layer1_outputs[4995] = ~(layer0_outputs[10570]);
    assign layer1_outputs[4996] = ~(layer0_outputs[7004]);
    assign layer1_outputs[4997] = layer0_outputs[6972];
    assign layer1_outputs[4998] = ~(layer0_outputs[5619]);
    assign layer1_outputs[4999] = (layer0_outputs[3237]) | (layer0_outputs[2888]);
    assign layer1_outputs[5000] = ~((layer0_outputs[1864]) | (layer0_outputs[1175]));
    assign layer1_outputs[5001] = ~(layer0_outputs[4081]) | (layer0_outputs[1085]);
    assign layer1_outputs[5002] = ~(layer0_outputs[12489]) | (layer0_outputs[10498]);
    assign layer1_outputs[5003] = ~(layer0_outputs[8493]);
    assign layer1_outputs[5004] = ~(layer0_outputs[267]);
    assign layer1_outputs[5005] = ~(layer0_outputs[1464]);
    assign layer1_outputs[5006] = layer0_outputs[9034];
    assign layer1_outputs[5007] = ~((layer0_outputs[5176]) & (layer0_outputs[11151]));
    assign layer1_outputs[5008] = ~(layer0_outputs[10778]);
    assign layer1_outputs[5009] = ~(layer0_outputs[4296]);
    assign layer1_outputs[5010] = ~(layer0_outputs[10768]);
    assign layer1_outputs[5011] = ~((layer0_outputs[5748]) & (layer0_outputs[10040]));
    assign layer1_outputs[5012] = layer0_outputs[11387];
    assign layer1_outputs[5013] = ~(layer0_outputs[7339]);
    assign layer1_outputs[5014] = ~(layer0_outputs[9264]) | (layer0_outputs[400]);
    assign layer1_outputs[5015] = ~(layer0_outputs[2197]);
    assign layer1_outputs[5016] = (layer0_outputs[8823]) & (layer0_outputs[2301]);
    assign layer1_outputs[5017] = (layer0_outputs[11345]) & ~(layer0_outputs[7318]);
    assign layer1_outputs[5018] = ~((layer0_outputs[12399]) & (layer0_outputs[5763]));
    assign layer1_outputs[5019] = layer0_outputs[12168];
    assign layer1_outputs[5020] = ~(layer0_outputs[6564]) | (layer0_outputs[391]);
    assign layer1_outputs[5021] = layer0_outputs[10287];
    assign layer1_outputs[5022] = (layer0_outputs[11804]) & (layer0_outputs[6470]);
    assign layer1_outputs[5023] = layer0_outputs[10201];
    assign layer1_outputs[5024] = layer0_outputs[1575];
    assign layer1_outputs[5025] = ~(layer0_outputs[7029]) | (layer0_outputs[7878]);
    assign layer1_outputs[5026] = ~(layer0_outputs[8037]) | (layer0_outputs[6942]);
    assign layer1_outputs[5027] = (layer0_outputs[2277]) | (layer0_outputs[8262]);
    assign layer1_outputs[5028] = ~((layer0_outputs[4325]) | (layer0_outputs[8132]));
    assign layer1_outputs[5029] = 1'b0;
    assign layer1_outputs[5030] = ~(layer0_outputs[6766]) | (layer0_outputs[12172]);
    assign layer1_outputs[5031] = ~(layer0_outputs[9689]);
    assign layer1_outputs[5032] = (layer0_outputs[6167]) | (layer0_outputs[4269]);
    assign layer1_outputs[5033] = layer0_outputs[4945];
    assign layer1_outputs[5034] = ~((layer0_outputs[11464]) | (layer0_outputs[2646]));
    assign layer1_outputs[5035] = layer0_outputs[2212];
    assign layer1_outputs[5036] = (layer0_outputs[7275]) & (layer0_outputs[5378]);
    assign layer1_outputs[5037] = (layer0_outputs[12366]) & ~(layer0_outputs[1171]);
    assign layer1_outputs[5038] = (layer0_outputs[11288]) ^ (layer0_outputs[565]);
    assign layer1_outputs[5039] = ~((layer0_outputs[2294]) ^ (layer0_outputs[5204]));
    assign layer1_outputs[5040] = (layer0_outputs[4116]) & ~(layer0_outputs[8886]);
    assign layer1_outputs[5041] = ~(layer0_outputs[10192]) | (layer0_outputs[7466]);
    assign layer1_outputs[5042] = layer0_outputs[6127];
    assign layer1_outputs[5043] = (layer0_outputs[982]) & ~(layer0_outputs[6470]);
    assign layer1_outputs[5044] = layer0_outputs[3821];
    assign layer1_outputs[5045] = ~((layer0_outputs[10352]) | (layer0_outputs[1278]));
    assign layer1_outputs[5046] = 1'b0;
    assign layer1_outputs[5047] = ~((layer0_outputs[12573]) ^ (layer0_outputs[3491]));
    assign layer1_outputs[5048] = ~((layer0_outputs[3689]) | (layer0_outputs[3416]));
    assign layer1_outputs[5049] = ~((layer0_outputs[8644]) | (layer0_outputs[11538]));
    assign layer1_outputs[5050] = (layer0_outputs[3569]) & (layer0_outputs[7117]);
    assign layer1_outputs[5051] = layer0_outputs[5464];
    assign layer1_outputs[5052] = (layer0_outputs[230]) & ~(layer0_outputs[11931]);
    assign layer1_outputs[5053] = ~((layer0_outputs[8118]) | (layer0_outputs[8]));
    assign layer1_outputs[5054] = (layer0_outputs[3800]) | (layer0_outputs[6011]);
    assign layer1_outputs[5055] = (layer0_outputs[10902]) & (layer0_outputs[7732]);
    assign layer1_outputs[5056] = (layer0_outputs[3619]) & (layer0_outputs[5358]);
    assign layer1_outputs[5057] = ~(layer0_outputs[4265]) | (layer0_outputs[2211]);
    assign layer1_outputs[5058] = ~(layer0_outputs[11428]);
    assign layer1_outputs[5059] = (layer0_outputs[8416]) & (layer0_outputs[152]);
    assign layer1_outputs[5060] = ~(layer0_outputs[5335]) | (layer0_outputs[1390]);
    assign layer1_outputs[5061] = ~(layer0_outputs[10095]) | (layer0_outputs[6885]);
    assign layer1_outputs[5062] = layer0_outputs[9372];
    assign layer1_outputs[5063] = (layer0_outputs[7714]) & ~(layer0_outputs[689]);
    assign layer1_outputs[5064] = 1'b1;
    assign layer1_outputs[5065] = layer0_outputs[3804];
    assign layer1_outputs[5066] = ~(layer0_outputs[10153]) | (layer0_outputs[252]);
    assign layer1_outputs[5067] = (layer0_outputs[10273]) & ~(layer0_outputs[5284]);
    assign layer1_outputs[5068] = (layer0_outputs[2957]) & (layer0_outputs[8933]);
    assign layer1_outputs[5069] = ~(layer0_outputs[12167]);
    assign layer1_outputs[5070] = ~(layer0_outputs[5458]) | (layer0_outputs[5980]);
    assign layer1_outputs[5071] = (layer0_outputs[7238]) & ~(layer0_outputs[4373]);
    assign layer1_outputs[5072] = (layer0_outputs[835]) & ~(layer0_outputs[9579]);
    assign layer1_outputs[5073] = layer0_outputs[6854];
    assign layer1_outputs[5074] = ~(layer0_outputs[11377]) | (layer0_outputs[1863]);
    assign layer1_outputs[5075] = (layer0_outputs[7932]) & ~(layer0_outputs[5200]);
    assign layer1_outputs[5076] = layer0_outputs[2346];
    assign layer1_outputs[5077] = (layer0_outputs[9956]) | (layer0_outputs[1308]);
    assign layer1_outputs[5078] = (layer0_outputs[4247]) & ~(layer0_outputs[103]);
    assign layer1_outputs[5079] = ~(layer0_outputs[11003]) | (layer0_outputs[6796]);
    assign layer1_outputs[5080] = (layer0_outputs[3295]) & ~(layer0_outputs[3877]);
    assign layer1_outputs[5081] = ~(layer0_outputs[8112]) | (layer0_outputs[6065]);
    assign layer1_outputs[5082] = layer0_outputs[4275];
    assign layer1_outputs[5083] = ~((layer0_outputs[1165]) & (layer0_outputs[4454]));
    assign layer1_outputs[5084] = ~(layer0_outputs[6377]);
    assign layer1_outputs[5085] = (layer0_outputs[4161]) & ~(layer0_outputs[9708]);
    assign layer1_outputs[5086] = ~((layer0_outputs[10060]) ^ (layer0_outputs[784]));
    assign layer1_outputs[5087] = ~((layer0_outputs[9143]) & (layer0_outputs[3513]));
    assign layer1_outputs[5088] = layer0_outputs[3103];
    assign layer1_outputs[5089] = (layer0_outputs[550]) & ~(layer0_outputs[11435]);
    assign layer1_outputs[5090] = 1'b0;
    assign layer1_outputs[5091] = layer0_outputs[6643];
    assign layer1_outputs[5092] = (layer0_outputs[7968]) | (layer0_outputs[422]);
    assign layer1_outputs[5093] = (layer0_outputs[4815]) | (layer0_outputs[9161]);
    assign layer1_outputs[5094] = (layer0_outputs[6263]) & ~(layer0_outputs[3172]);
    assign layer1_outputs[5095] = ~(layer0_outputs[4527]);
    assign layer1_outputs[5096] = ~(layer0_outputs[5799]);
    assign layer1_outputs[5097] = (layer0_outputs[3264]) & (layer0_outputs[6701]);
    assign layer1_outputs[5098] = ~(layer0_outputs[8263]);
    assign layer1_outputs[5099] = ~(layer0_outputs[4251]) | (layer0_outputs[1476]);
    assign layer1_outputs[5100] = ~((layer0_outputs[425]) | (layer0_outputs[7524]));
    assign layer1_outputs[5101] = ~(layer0_outputs[3614]) | (layer0_outputs[2755]);
    assign layer1_outputs[5102] = 1'b1;
    assign layer1_outputs[5103] = ~(layer0_outputs[8834]);
    assign layer1_outputs[5104] = ~(layer0_outputs[7195]);
    assign layer1_outputs[5105] = (layer0_outputs[4751]) & ~(layer0_outputs[2844]);
    assign layer1_outputs[5106] = (layer0_outputs[2395]) & (layer0_outputs[5601]);
    assign layer1_outputs[5107] = layer0_outputs[293];
    assign layer1_outputs[5108] = layer0_outputs[4094];
    assign layer1_outputs[5109] = (layer0_outputs[1550]) | (layer0_outputs[2557]);
    assign layer1_outputs[5110] = (layer0_outputs[11171]) & (layer0_outputs[6350]);
    assign layer1_outputs[5111] = (layer0_outputs[5961]) | (layer0_outputs[10102]);
    assign layer1_outputs[5112] = (layer0_outputs[4820]) & (layer0_outputs[520]);
    assign layer1_outputs[5113] = 1'b0;
    assign layer1_outputs[5114] = ~(layer0_outputs[4512]) | (layer0_outputs[5869]);
    assign layer1_outputs[5115] = ~((layer0_outputs[2272]) ^ (layer0_outputs[1451]));
    assign layer1_outputs[5116] = ~((layer0_outputs[1469]) | (layer0_outputs[7019]));
    assign layer1_outputs[5117] = ~(layer0_outputs[6608]) | (layer0_outputs[12622]);
    assign layer1_outputs[5118] = ~(layer0_outputs[1941]);
    assign layer1_outputs[5119] = (layer0_outputs[5692]) | (layer0_outputs[11188]);
    assign layer1_outputs[5120] = (layer0_outputs[6024]) & (layer0_outputs[9898]);
    assign layer1_outputs[5121] = ~(layer0_outputs[4521]);
    assign layer1_outputs[5122] = ~(layer0_outputs[2415]);
    assign layer1_outputs[5123] = (layer0_outputs[7970]) & (layer0_outputs[4207]);
    assign layer1_outputs[5124] = ~(layer0_outputs[670]);
    assign layer1_outputs[5125] = ~((layer0_outputs[3462]) & (layer0_outputs[11454]));
    assign layer1_outputs[5126] = ~((layer0_outputs[7719]) & (layer0_outputs[1443]));
    assign layer1_outputs[5127] = layer0_outputs[4382];
    assign layer1_outputs[5128] = ~(layer0_outputs[7841]) | (layer0_outputs[3775]);
    assign layer1_outputs[5129] = ~(layer0_outputs[12481]);
    assign layer1_outputs[5130] = (layer0_outputs[2932]) & (layer0_outputs[11455]);
    assign layer1_outputs[5131] = (layer0_outputs[4112]) ^ (layer0_outputs[2073]);
    assign layer1_outputs[5132] = layer0_outputs[5650];
    assign layer1_outputs[5133] = (layer0_outputs[4268]) & ~(layer0_outputs[4556]);
    assign layer1_outputs[5134] = ~(layer0_outputs[12713]);
    assign layer1_outputs[5135] = (layer0_outputs[3806]) & ~(layer0_outputs[2352]);
    assign layer1_outputs[5136] = ~((layer0_outputs[3222]) & (layer0_outputs[2673]));
    assign layer1_outputs[5137] = (layer0_outputs[1053]) | (layer0_outputs[12623]);
    assign layer1_outputs[5138] = (layer0_outputs[8641]) & ~(layer0_outputs[11722]);
    assign layer1_outputs[5139] = (layer0_outputs[1793]) | (layer0_outputs[12050]);
    assign layer1_outputs[5140] = ~((layer0_outputs[9497]) | (layer0_outputs[4234]));
    assign layer1_outputs[5141] = ~(layer0_outputs[9819]);
    assign layer1_outputs[5142] = (layer0_outputs[4748]) & (layer0_outputs[1416]);
    assign layer1_outputs[5143] = (layer0_outputs[6269]) & (layer0_outputs[387]);
    assign layer1_outputs[5144] = (layer0_outputs[1198]) | (layer0_outputs[4201]);
    assign layer1_outputs[5145] = ~(layer0_outputs[6385]) | (layer0_outputs[2241]);
    assign layer1_outputs[5146] = ~(layer0_outputs[7922]);
    assign layer1_outputs[5147] = layer0_outputs[161];
    assign layer1_outputs[5148] = layer0_outputs[8544];
    assign layer1_outputs[5149] = layer0_outputs[4923];
    assign layer1_outputs[5150] = (layer0_outputs[12548]) & ~(layer0_outputs[4384]);
    assign layer1_outputs[5151] = 1'b0;
    assign layer1_outputs[5152] = layer0_outputs[10473];
    assign layer1_outputs[5153] = (layer0_outputs[10320]) & ~(layer0_outputs[10184]);
    assign layer1_outputs[5154] = (layer0_outputs[4642]) & ~(layer0_outputs[1137]);
    assign layer1_outputs[5155] = layer0_outputs[6237];
    assign layer1_outputs[5156] = ~(layer0_outputs[10436]);
    assign layer1_outputs[5157] = layer0_outputs[11357];
    assign layer1_outputs[5158] = (layer0_outputs[11795]) ^ (layer0_outputs[8298]);
    assign layer1_outputs[5159] = (layer0_outputs[8057]) | (layer0_outputs[7954]);
    assign layer1_outputs[5160] = ~((layer0_outputs[11684]) & (layer0_outputs[1448]));
    assign layer1_outputs[5161] = ~((layer0_outputs[10409]) | (layer0_outputs[4140]));
    assign layer1_outputs[5162] = (layer0_outputs[5974]) & (layer0_outputs[11417]);
    assign layer1_outputs[5163] = ~(layer0_outputs[3138]);
    assign layer1_outputs[5164] = ~((layer0_outputs[10523]) | (layer0_outputs[10894]));
    assign layer1_outputs[5165] = layer0_outputs[9974];
    assign layer1_outputs[5166] = (layer0_outputs[4409]) & (layer0_outputs[10192]);
    assign layer1_outputs[5167] = (layer0_outputs[4529]) | (layer0_outputs[4879]);
    assign layer1_outputs[5168] = (layer0_outputs[8658]) & ~(layer0_outputs[8337]);
    assign layer1_outputs[5169] = ~(layer0_outputs[5968]);
    assign layer1_outputs[5170] = ~(layer0_outputs[7905]);
    assign layer1_outputs[5171] = ~((layer0_outputs[3921]) & (layer0_outputs[11901]));
    assign layer1_outputs[5172] = ~(layer0_outputs[10648]) | (layer0_outputs[2830]);
    assign layer1_outputs[5173] = (layer0_outputs[8174]) ^ (layer0_outputs[5958]);
    assign layer1_outputs[5174] = layer0_outputs[6798];
    assign layer1_outputs[5175] = ~(layer0_outputs[1648]);
    assign layer1_outputs[5176] = (layer0_outputs[4883]) | (layer0_outputs[6830]);
    assign layer1_outputs[5177] = ~(layer0_outputs[8789]) | (layer0_outputs[1272]);
    assign layer1_outputs[5178] = ~((layer0_outputs[2623]) | (layer0_outputs[274]));
    assign layer1_outputs[5179] = ~((layer0_outputs[8429]) | (layer0_outputs[1271]));
    assign layer1_outputs[5180] = ~((layer0_outputs[2624]) & (layer0_outputs[5540]));
    assign layer1_outputs[5181] = layer0_outputs[9016];
    assign layer1_outputs[5182] = (layer0_outputs[8941]) & ~(layer0_outputs[6906]);
    assign layer1_outputs[5183] = ~(layer0_outputs[765]) | (layer0_outputs[10809]);
    assign layer1_outputs[5184] = ~(layer0_outputs[6383]);
    assign layer1_outputs[5185] = layer0_outputs[1512];
    assign layer1_outputs[5186] = ~((layer0_outputs[2870]) ^ (layer0_outputs[7521]));
    assign layer1_outputs[5187] = ~(layer0_outputs[7497]);
    assign layer1_outputs[5188] = ~(layer0_outputs[5816]) | (layer0_outputs[8771]);
    assign layer1_outputs[5189] = ~(layer0_outputs[8884]);
    assign layer1_outputs[5190] = (layer0_outputs[492]) | (layer0_outputs[12486]);
    assign layer1_outputs[5191] = ~(layer0_outputs[7869]) | (layer0_outputs[11977]);
    assign layer1_outputs[5192] = 1'b0;
    assign layer1_outputs[5193] = 1'b1;
    assign layer1_outputs[5194] = ~(layer0_outputs[3087]) | (layer0_outputs[10440]);
    assign layer1_outputs[5195] = ~(layer0_outputs[1035]);
    assign layer1_outputs[5196] = (layer0_outputs[6514]) ^ (layer0_outputs[8393]);
    assign layer1_outputs[5197] = ~(layer0_outputs[4080]);
    assign layer1_outputs[5198] = (layer0_outputs[11550]) & (layer0_outputs[9396]);
    assign layer1_outputs[5199] = layer0_outputs[5504];
    assign layer1_outputs[5200] = layer0_outputs[6863];
    assign layer1_outputs[5201] = ~(layer0_outputs[8278]);
    assign layer1_outputs[5202] = (layer0_outputs[498]) & (layer0_outputs[5169]);
    assign layer1_outputs[5203] = (layer0_outputs[683]) & ~(layer0_outputs[5858]);
    assign layer1_outputs[5204] = ~((layer0_outputs[7478]) & (layer0_outputs[2969]));
    assign layer1_outputs[5205] = (layer0_outputs[4158]) & ~(layer0_outputs[2173]);
    assign layer1_outputs[5206] = layer0_outputs[7001];
    assign layer1_outputs[5207] = (layer0_outputs[199]) & ~(layer0_outputs[5151]);
    assign layer1_outputs[5208] = ~((layer0_outputs[12267]) ^ (layer0_outputs[3642]));
    assign layer1_outputs[5209] = ~(layer0_outputs[1244]);
    assign layer1_outputs[5210] = ~((layer0_outputs[9817]) | (layer0_outputs[5058]));
    assign layer1_outputs[5211] = ~((layer0_outputs[7701]) | (layer0_outputs[11625]));
    assign layer1_outputs[5212] = ~((layer0_outputs[9884]) | (layer0_outputs[10508]));
    assign layer1_outputs[5213] = ~(layer0_outputs[11827]);
    assign layer1_outputs[5214] = layer0_outputs[286];
    assign layer1_outputs[5215] = layer0_outputs[11159];
    assign layer1_outputs[5216] = (layer0_outputs[12389]) | (layer0_outputs[12300]);
    assign layer1_outputs[5217] = ~(layer0_outputs[2520]) | (layer0_outputs[2864]);
    assign layer1_outputs[5218] = (layer0_outputs[12304]) ^ (layer0_outputs[10389]);
    assign layer1_outputs[5219] = ~(layer0_outputs[7454]);
    assign layer1_outputs[5220] = ~(layer0_outputs[12346]);
    assign layer1_outputs[5221] = ~(layer0_outputs[5385]) | (layer0_outputs[467]);
    assign layer1_outputs[5222] = ~(layer0_outputs[10122]) | (layer0_outputs[5460]);
    assign layer1_outputs[5223] = (layer0_outputs[9500]) | (layer0_outputs[7557]);
    assign layer1_outputs[5224] = ~(layer0_outputs[9817]);
    assign layer1_outputs[5225] = 1'b1;
    assign layer1_outputs[5226] = ~(layer0_outputs[1206]);
    assign layer1_outputs[5227] = ~((layer0_outputs[9068]) | (layer0_outputs[9125]));
    assign layer1_outputs[5228] = (layer0_outputs[6335]) & ~(layer0_outputs[12206]);
    assign layer1_outputs[5229] = ~(layer0_outputs[10471]) | (layer0_outputs[8252]);
    assign layer1_outputs[5230] = ~(layer0_outputs[2480]);
    assign layer1_outputs[5231] = ~(layer0_outputs[2593]);
    assign layer1_outputs[5232] = layer0_outputs[1879];
    assign layer1_outputs[5233] = layer0_outputs[4191];
    assign layer1_outputs[5234] = (layer0_outputs[7006]) ^ (layer0_outputs[11143]);
    assign layer1_outputs[5235] = layer0_outputs[12079];
    assign layer1_outputs[5236] = layer0_outputs[12273];
    assign layer1_outputs[5237] = ~(layer0_outputs[9943]) | (layer0_outputs[375]);
    assign layer1_outputs[5238] = ~(layer0_outputs[7987]);
    assign layer1_outputs[5239] = ~(layer0_outputs[9070]);
    assign layer1_outputs[5240] = (layer0_outputs[1556]) & ~(layer0_outputs[2975]);
    assign layer1_outputs[5241] = layer0_outputs[262];
    assign layer1_outputs[5242] = (layer0_outputs[4242]) & ~(layer0_outputs[9767]);
    assign layer1_outputs[5243] = layer0_outputs[3780];
    assign layer1_outputs[5244] = ~((layer0_outputs[9674]) & (layer0_outputs[7187]));
    assign layer1_outputs[5245] = ~(layer0_outputs[10987]);
    assign layer1_outputs[5246] = ~((layer0_outputs[10064]) ^ (layer0_outputs[2796]));
    assign layer1_outputs[5247] = ~(layer0_outputs[3204]) | (layer0_outputs[3212]);
    assign layer1_outputs[5248] = ~(layer0_outputs[9498]);
    assign layer1_outputs[5249] = ~(layer0_outputs[11658]) | (layer0_outputs[10620]);
    assign layer1_outputs[5250] = ~(layer0_outputs[9812]) | (layer0_outputs[9325]);
    assign layer1_outputs[5251] = ~(layer0_outputs[9019]) | (layer0_outputs[1455]);
    assign layer1_outputs[5252] = ~((layer0_outputs[6876]) | (layer0_outputs[12445]));
    assign layer1_outputs[5253] = ~(layer0_outputs[10854]);
    assign layer1_outputs[5254] = ~(layer0_outputs[1633]) | (layer0_outputs[1399]);
    assign layer1_outputs[5255] = ~(layer0_outputs[11366]);
    assign layer1_outputs[5256] = (layer0_outputs[5363]) | (layer0_outputs[9830]);
    assign layer1_outputs[5257] = ~(layer0_outputs[11681]) | (layer0_outputs[10377]);
    assign layer1_outputs[5258] = 1'b1;
    assign layer1_outputs[5259] = ~(layer0_outputs[7375]) | (layer0_outputs[7211]);
    assign layer1_outputs[5260] = (layer0_outputs[254]) & ~(layer0_outputs[382]);
    assign layer1_outputs[5261] = ~(layer0_outputs[86]);
    assign layer1_outputs[5262] = ~((layer0_outputs[2195]) | (layer0_outputs[5942]));
    assign layer1_outputs[5263] = ~((layer0_outputs[2453]) & (layer0_outputs[2301]));
    assign layer1_outputs[5264] = (layer0_outputs[1841]) ^ (layer0_outputs[11585]);
    assign layer1_outputs[5265] = (layer0_outputs[11872]) ^ (layer0_outputs[2787]);
    assign layer1_outputs[5266] = (layer0_outputs[11156]) ^ (layer0_outputs[9504]);
    assign layer1_outputs[5267] = ~(layer0_outputs[665]);
    assign layer1_outputs[5268] = (layer0_outputs[10556]) & ~(layer0_outputs[7989]);
    assign layer1_outputs[5269] = ~(layer0_outputs[9624]);
    assign layer1_outputs[5270] = (layer0_outputs[2464]) & ~(layer0_outputs[3366]);
    assign layer1_outputs[5271] = layer0_outputs[585];
    assign layer1_outputs[5272] = ~(layer0_outputs[360]) | (layer0_outputs[567]);
    assign layer1_outputs[5273] = (layer0_outputs[5745]) & ~(layer0_outputs[12206]);
    assign layer1_outputs[5274] = ~(layer0_outputs[7705]);
    assign layer1_outputs[5275] = ~(layer0_outputs[10276]) | (layer0_outputs[5657]);
    assign layer1_outputs[5276] = layer0_outputs[6851];
    assign layer1_outputs[5277] = ~(layer0_outputs[4557]);
    assign layer1_outputs[5278] = layer0_outputs[4672];
    assign layer1_outputs[5279] = layer0_outputs[3064];
    assign layer1_outputs[5280] = ~(layer0_outputs[12210]);
    assign layer1_outputs[5281] = layer0_outputs[7395];
    assign layer1_outputs[5282] = ~(layer0_outputs[7368]) | (layer0_outputs[4082]);
    assign layer1_outputs[5283] = 1'b0;
    assign layer1_outputs[5284] = ~(layer0_outputs[2067]) | (layer0_outputs[2464]);
    assign layer1_outputs[5285] = ~(layer0_outputs[5796]);
    assign layer1_outputs[5286] = ~(layer0_outputs[12023]) | (layer0_outputs[8935]);
    assign layer1_outputs[5287] = layer0_outputs[6486];
    assign layer1_outputs[5288] = layer0_outputs[8212];
    assign layer1_outputs[5289] = layer0_outputs[7240];
    assign layer1_outputs[5290] = 1'b1;
    assign layer1_outputs[5291] = layer0_outputs[11544];
    assign layer1_outputs[5292] = ~(layer0_outputs[1606]) | (layer0_outputs[10142]);
    assign layer1_outputs[5293] = ~(layer0_outputs[2910]);
    assign layer1_outputs[5294] = ~((layer0_outputs[7002]) | (layer0_outputs[5507]));
    assign layer1_outputs[5295] = ~((layer0_outputs[10883]) ^ (layer0_outputs[10895]));
    assign layer1_outputs[5296] = (layer0_outputs[7589]) ^ (layer0_outputs[8337]);
    assign layer1_outputs[5297] = ~((layer0_outputs[3074]) | (layer0_outputs[6934]));
    assign layer1_outputs[5298] = ~(layer0_outputs[1733]);
    assign layer1_outputs[5299] = ~(layer0_outputs[9921]) | (layer0_outputs[11916]);
    assign layer1_outputs[5300] = ~(layer0_outputs[304]);
    assign layer1_outputs[5301] = (layer0_outputs[5225]) & ~(layer0_outputs[9482]);
    assign layer1_outputs[5302] = ~((layer0_outputs[7543]) ^ (layer0_outputs[12242]));
    assign layer1_outputs[5303] = ~(layer0_outputs[5020]) | (layer0_outputs[5109]);
    assign layer1_outputs[5304] = (layer0_outputs[2378]) & ~(layer0_outputs[2542]);
    assign layer1_outputs[5305] = layer0_outputs[12497];
    assign layer1_outputs[5306] = ~(layer0_outputs[10131]);
    assign layer1_outputs[5307] = (layer0_outputs[8909]) & ~(layer0_outputs[5860]);
    assign layer1_outputs[5308] = layer0_outputs[8245];
    assign layer1_outputs[5309] = layer0_outputs[6543];
    assign layer1_outputs[5310] = (layer0_outputs[299]) & ~(layer0_outputs[1238]);
    assign layer1_outputs[5311] = layer0_outputs[1448];
    assign layer1_outputs[5312] = ~(layer0_outputs[5999]);
    assign layer1_outputs[5313] = (layer0_outputs[9569]) ^ (layer0_outputs[8797]);
    assign layer1_outputs[5314] = ~(layer0_outputs[7481]) | (layer0_outputs[12762]);
    assign layer1_outputs[5315] = ~(layer0_outputs[3283]) | (layer0_outputs[8038]);
    assign layer1_outputs[5316] = (layer0_outputs[3174]) ^ (layer0_outputs[8708]);
    assign layer1_outputs[5317] = ~(layer0_outputs[8822]);
    assign layer1_outputs[5318] = ~(layer0_outputs[6414]);
    assign layer1_outputs[5319] = layer0_outputs[1426];
    assign layer1_outputs[5320] = ~(layer0_outputs[6152]);
    assign layer1_outputs[5321] = (layer0_outputs[7601]) | (layer0_outputs[7963]);
    assign layer1_outputs[5322] = (layer0_outputs[5763]) & ~(layer0_outputs[9982]);
    assign layer1_outputs[5323] = 1'b0;
    assign layer1_outputs[5324] = layer0_outputs[4802];
    assign layer1_outputs[5325] = ~((layer0_outputs[773]) & (layer0_outputs[11509]));
    assign layer1_outputs[5326] = ~(layer0_outputs[11666]);
    assign layer1_outputs[5327] = (layer0_outputs[2206]) | (layer0_outputs[11712]);
    assign layer1_outputs[5328] = ~(layer0_outputs[182]);
    assign layer1_outputs[5329] = (layer0_outputs[10261]) & (layer0_outputs[10995]);
    assign layer1_outputs[5330] = (layer0_outputs[3208]) | (layer0_outputs[5921]);
    assign layer1_outputs[5331] = (layer0_outputs[5958]) & ~(layer0_outputs[7373]);
    assign layer1_outputs[5332] = ~(layer0_outputs[2182]) | (layer0_outputs[1587]);
    assign layer1_outputs[5333] = ~((layer0_outputs[4475]) | (layer0_outputs[5799]));
    assign layer1_outputs[5334] = layer0_outputs[1585];
    assign layer1_outputs[5335] = layer0_outputs[10633];
    assign layer1_outputs[5336] = ~(layer0_outputs[7309]);
    assign layer1_outputs[5337] = (layer0_outputs[8649]) & ~(layer0_outputs[12724]);
    assign layer1_outputs[5338] = layer0_outputs[7350];
    assign layer1_outputs[5339] = 1'b1;
    assign layer1_outputs[5340] = ~((layer0_outputs[6649]) | (layer0_outputs[6547]));
    assign layer1_outputs[5341] = layer0_outputs[4984];
    assign layer1_outputs[5342] = (layer0_outputs[11575]) ^ (layer0_outputs[6859]);
    assign layer1_outputs[5343] = layer0_outputs[939];
    assign layer1_outputs[5344] = ~((layer0_outputs[1033]) & (layer0_outputs[8610]));
    assign layer1_outputs[5345] = layer0_outputs[6435];
    assign layer1_outputs[5346] = layer0_outputs[5330];
    assign layer1_outputs[5347] = ~(layer0_outputs[3439]);
    assign layer1_outputs[5348] = ~(layer0_outputs[6611]);
    assign layer1_outputs[5349] = layer0_outputs[4333];
    assign layer1_outputs[5350] = (layer0_outputs[10009]) & (layer0_outputs[7842]);
    assign layer1_outputs[5351] = layer0_outputs[7008];
    assign layer1_outputs[5352] = layer0_outputs[8182];
    assign layer1_outputs[5353] = layer0_outputs[10822];
    assign layer1_outputs[5354] = 1'b0;
    assign layer1_outputs[5355] = ~(layer0_outputs[5081]);
    assign layer1_outputs[5356] = ~(layer0_outputs[10275]);
    assign layer1_outputs[5357] = layer0_outputs[781];
    assign layer1_outputs[5358] = (layer0_outputs[8074]) & ~(layer0_outputs[2667]);
    assign layer1_outputs[5359] = (layer0_outputs[12061]) & ~(layer0_outputs[7131]);
    assign layer1_outputs[5360] = (layer0_outputs[8788]) | (layer0_outputs[3639]);
    assign layer1_outputs[5361] = layer0_outputs[7939];
    assign layer1_outputs[5362] = ~((layer0_outputs[6240]) | (layer0_outputs[9089]));
    assign layer1_outputs[5363] = ~(layer0_outputs[8223]);
    assign layer1_outputs[5364] = layer0_outputs[5309];
    assign layer1_outputs[5365] = layer0_outputs[7133];
    assign layer1_outputs[5366] = ~(layer0_outputs[6527]);
    assign layer1_outputs[5367] = ~(layer0_outputs[11297]) | (layer0_outputs[8806]);
    assign layer1_outputs[5368] = (layer0_outputs[1099]) & (layer0_outputs[6684]);
    assign layer1_outputs[5369] = ~(layer0_outputs[3963]);
    assign layer1_outputs[5370] = layer0_outputs[1977];
    assign layer1_outputs[5371] = ~(layer0_outputs[1743]);
    assign layer1_outputs[5372] = ~((layer0_outputs[3328]) | (layer0_outputs[7649]));
    assign layer1_outputs[5373] = ~((layer0_outputs[11284]) | (layer0_outputs[6792]));
    assign layer1_outputs[5374] = ~(layer0_outputs[1192]);
    assign layer1_outputs[5375] = (layer0_outputs[7368]) ^ (layer0_outputs[9298]);
    assign layer1_outputs[5376] = ~(layer0_outputs[6760]);
    assign layer1_outputs[5377] = ~(layer0_outputs[1827]) | (layer0_outputs[5235]);
    assign layer1_outputs[5378] = ~((layer0_outputs[4396]) | (layer0_outputs[1040]));
    assign layer1_outputs[5379] = layer0_outputs[10004];
    assign layer1_outputs[5380] = (layer0_outputs[9160]) ^ (layer0_outputs[7161]);
    assign layer1_outputs[5381] = layer0_outputs[1924];
    assign layer1_outputs[5382] = layer0_outputs[2777];
    assign layer1_outputs[5383] = ~(layer0_outputs[4355]);
    assign layer1_outputs[5384] = ~(layer0_outputs[10886]) | (layer0_outputs[6147]);
    assign layer1_outputs[5385] = ~((layer0_outputs[2275]) | (layer0_outputs[10850]));
    assign layer1_outputs[5386] = ~(layer0_outputs[8181]) | (layer0_outputs[10829]);
    assign layer1_outputs[5387] = ~(layer0_outputs[11350]) | (layer0_outputs[6292]);
    assign layer1_outputs[5388] = layer0_outputs[11186];
    assign layer1_outputs[5389] = layer0_outputs[12690];
    assign layer1_outputs[5390] = (layer0_outputs[10454]) & (layer0_outputs[11699]);
    assign layer1_outputs[5391] = ~((layer0_outputs[10228]) & (layer0_outputs[512]));
    assign layer1_outputs[5392] = layer0_outputs[4441];
    assign layer1_outputs[5393] = ~(layer0_outputs[6408]) | (layer0_outputs[5859]);
    assign layer1_outputs[5394] = ~((layer0_outputs[4193]) & (layer0_outputs[3414]));
    assign layer1_outputs[5395] = (layer0_outputs[8026]) & ~(layer0_outputs[10364]);
    assign layer1_outputs[5396] = ~((layer0_outputs[5279]) & (layer0_outputs[4091]));
    assign layer1_outputs[5397] = ~(layer0_outputs[5101]);
    assign layer1_outputs[5398] = (layer0_outputs[888]) ^ (layer0_outputs[388]);
    assign layer1_outputs[5399] = layer0_outputs[11957];
    assign layer1_outputs[5400] = ~(layer0_outputs[10558]);
    assign layer1_outputs[5401] = layer0_outputs[2379];
    assign layer1_outputs[5402] = layer0_outputs[9465];
    assign layer1_outputs[5403] = ~((layer0_outputs[4292]) | (layer0_outputs[12672]));
    assign layer1_outputs[5404] = layer0_outputs[5639];
    assign layer1_outputs[5405] = layer0_outputs[6219];
    assign layer1_outputs[5406] = (layer0_outputs[9983]) | (layer0_outputs[5106]);
    assign layer1_outputs[5407] = ~(layer0_outputs[10687]) | (layer0_outputs[4517]);
    assign layer1_outputs[5408] = ~(layer0_outputs[5197]);
    assign layer1_outputs[5409] = layer0_outputs[6981];
    assign layer1_outputs[5410] = ~(layer0_outputs[828]) | (layer0_outputs[4079]);
    assign layer1_outputs[5411] = layer0_outputs[5091];
    assign layer1_outputs[5412] = ~(layer0_outputs[9773]);
    assign layer1_outputs[5413] = 1'b0;
    assign layer1_outputs[5414] = ~((layer0_outputs[510]) | (layer0_outputs[4296]));
    assign layer1_outputs[5415] = (layer0_outputs[10848]) & (layer0_outputs[7700]);
    assign layer1_outputs[5416] = 1'b1;
    assign layer1_outputs[5417] = ~(layer0_outputs[7075]);
    assign layer1_outputs[5418] = ~(layer0_outputs[4684]);
    assign layer1_outputs[5419] = 1'b1;
    assign layer1_outputs[5420] = ~(layer0_outputs[8313]);
    assign layer1_outputs[5421] = (layer0_outputs[12194]) & (layer0_outputs[1587]);
    assign layer1_outputs[5422] = ~(layer0_outputs[6728]) | (layer0_outputs[5841]);
    assign layer1_outputs[5423] = ~((layer0_outputs[9142]) & (layer0_outputs[5401]));
    assign layer1_outputs[5424] = layer0_outputs[6049];
    assign layer1_outputs[5425] = ~(layer0_outputs[7020]);
    assign layer1_outputs[5426] = layer0_outputs[10867];
    assign layer1_outputs[5427] = ~(layer0_outputs[843]) | (layer0_outputs[4069]);
    assign layer1_outputs[5428] = layer0_outputs[9392];
    assign layer1_outputs[5429] = layer0_outputs[4134];
    assign layer1_outputs[5430] = (layer0_outputs[7267]) & ~(layer0_outputs[10575]);
    assign layer1_outputs[5431] = ~(layer0_outputs[10567]);
    assign layer1_outputs[5432] = 1'b1;
    assign layer1_outputs[5433] = layer0_outputs[6019];
    assign layer1_outputs[5434] = ~(layer0_outputs[1216]);
    assign layer1_outputs[5435] = ~((layer0_outputs[4677]) & (layer0_outputs[7140]));
    assign layer1_outputs[5436] = layer0_outputs[1928];
    assign layer1_outputs[5437] = ~((layer0_outputs[6767]) & (layer0_outputs[1048]));
    assign layer1_outputs[5438] = ~(layer0_outputs[11783]) | (layer0_outputs[5000]);
    assign layer1_outputs[5439] = ~((layer0_outputs[5899]) ^ (layer0_outputs[3757]));
    assign layer1_outputs[5440] = (layer0_outputs[9913]) & ~(layer0_outputs[6592]);
    assign layer1_outputs[5441] = ~(layer0_outputs[1474]) | (layer0_outputs[321]);
    assign layer1_outputs[5442] = ~(layer0_outputs[4074]);
    assign layer1_outputs[5443] = ~((layer0_outputs[2140]) ^ (layer0_outputs[3102]));
    assign layer1_outputs[5444] = (layer0_outputs[3126]) ^ (layer0_outputs[1156]);
    assign layer1_outputs[5445] = ~(layer0_outputs[10746]) | (layer0_outputs[6391]);
    assign layer1_outputs[5446] = ~(layer0_outputs[5745]) | (layer0_outputs[4959]);
    assign layer1_outputs[5447] = layer0_outputs[10181];
    assign layer1_outputs[5448] = (layer0_outputs[2200]) & ~(layer0_outputs[490]);
    assign layer1_outputs[5449] = ~(layer0_outputs[4999]) | (layer0_outputs[2131]);
    assign layer1_outputs[5450] = ~(layer0_outputs[5374]) | (layer0_outputs[11708]);
    assign layer1_outputs[5451] = (layer0_outputs[2291]) & ~(layer0_outputs[9201]);
    assign layer1_outputs[5452] = (layer0_outputs[758]) | (layer0_outputs[3152]);
    assign layer1_outputs[5453] = layer0_outputs[8039];
    assign layer1_outputs[5454] = ~(layer0_outputs[1560]);
    assign layer1_outputs[5455] = ~(layer0_outputs[8409]);
    assign layer1_outputs[5456] = ~(layer0_outputs[7891]);
    assign layer1_outputs[5457] = (layer0_outputs[3005]) ^ (layer0_outputs[7459]);
    assign layer1_outputs[5458] = ~(layer0_outputs[4280]);
    assign layer1_outputs[5459] = layer0_outputs[1073];
    assign layer1_outputs[5460] = (layer0_outputs[11160]) & ~(layer0_outputs[2788]);
    assign layer1_outputs[5461] = (layer0_outputs[9573]) ^ (layer0_outputs[8575]);
    assign layer1_outputs[5462] = ~((layer0_outputs[2674]) ^ (layer0_outputs[3194]));
    assign layer1_outputs[5463] = ~(layer0_outputs[745]);
    assign layer1_outputs[5464] = layer0_outputs[6688];
    assign layer1_outputs[5465] = ~(layer0_outputs[12513]);
    assign layer1_outputs[5466] = (layer0_outputs[443]) & ~(layer0_outputs[4899]);
    assign layer1_outputs[5467] = (layer0_outputs[8189]) & ~(layer0_outputs[2434]);
    assign layer1_outputs[5468] = layer0_outputs[10270];
    assign layer1_outputs[5469] = ~(layer0_outputs[7192]) | (layer0_outputs[8127]);
    assign layer1_outputs[5470] = (layer0_outputs[6451]) & (layer0_outputs[2847]);
    assign layer1_outputs[5471] = layer0_outputs[3239];
    assign layer1_outputs[5472] = layer0_outputs[4231];
    assign layer1_outputs[5473] = (layer0_outputs[7995]) & ~(layer0_outputs[8531]);
    assign layer1_outputs[5474] = ~(layer0_outputs[3191]) | (layer0_outputs[2641]);
    assign layer1_outputs[5475] = layer0_outputs[1676];
    assign layer1_outputs[5476] = ~(layer0_outputs[1882]);
    assign layer1_outputs[5477] = ~(layer0_outputs[7494]);
    assign layer1_outputs[5478] = (layer0_outputs[6785]) & ~(layer0_outputs[7796]);
    assign layer1_outputs[5479] = 1'b1;
    assign layer1_outputs[5480] = ~(layer0_outputs[1786]) | (layer0_outputs[8634]);
    assign layer1_outputs[5481] = ~(layer0_outputs[12162]) | (layer0_outputs[11223]);
    assign layer1_outputs[5482] = (layer0_outputs[1695]) & ~(layer0_outputs[1440]);
    assign layer1_outputs[5483] = (layer0_outputs[3880]) & ~(layer0_outputs[1027]);
    assign layer1_outputs[5484] = ~(layer0_outputs[1338]) | (layer0_outputs[3564]);
    assign layer1_outputs[5485] = layer0_outputs[5418];
    assign layer1_outputs[5486] = (layer0_outputs[10306]) & ~(layer0_outputs[2015]);
    assign layer1_outputs[5487] = ~(layer0_outputs[864]);
    assign layer1_outputs[5488] = layer0_outputs[1965];
    assign layer1_outputs[5489] = ~((layer0_outputs[902]) | (layer0_outputs[11393]));
    assign layer1_outputs[5490] = ~(layer0_outputs[8377]) | (layer0_outputs[9993]);
    assign layer1_outputs[5491] = layer0_outputs[5155];
    assign layer1_outputs[5492] = ~(layer0_outputs[6407]) | (layer0_outputs[2442]);
    assign layer1_outputs[5493] = (layer0_outputs[1552]) & ~(layer0_outputs[2899]);
    assign layer1_outputs[5494] = (layer0_outputs[8190]) & ~(layer0_outputs[6939]);
    assign layer1_outputs[5495] = ~(layer0_outputs[2400]);
    assign layer1_outputs[5496] = (layer0_outputs[11619]) & ~(layer0_outputs[10977]);
    assign layer1_outputs[5497] = layer0_outputs[5444];
    assign layer1_outputs[5498] = (layer0_outputs[2640]) & ~(layer0_outputs[3050]);
    assign layer1_outputs[5499] = (layer0_outputs[11755]) & ~(layer0_outputs[1369]);
    assign layer1_outputs[5500] = ~(layer0_outputs[6951]);
    assign layer1_outputs[5501] = ~(layer0_outputs[11530]) | (layer0_outputs[6623]);
    assign layer1_outputs[5502] = (layer0_outputs[915]) & ~(layer0_outputs[3071]);
    assign layer1_outputs[5503] = ~((layer0_outputs[2254]) & (layer0_outputs[5434]));
    assign layer1_outputs[5504] = ~((layer0_outputs[5586]) | (layer0_outputs[3669]));
    assign layer1_outputs[5505] = ~(layer0_outputs[12447]);
    assign layer1_outputs[5506] = ~(layer0_outputs[2332]) | (layer0_outputs[3607]);
    assign layer1_outputs[5507] = (layer0_outputs[8034]) & ~(layer0_outputs[10931]);
    assign layer1_outputs[5508] = layer0_outputs[3596];
    assign layer1_outputs[5509] = (layer0_outputs[4657]) & ~(layer0_outputs[4084]);
    assign layer1_outputs[5510] = (layer0_outputs[953]) | (layer0_outputs[6546]);
    assign layer1_outputs[5511] = (layer0_outputs[2550]) ^ (layer0_outputs[1351]);
    assign layer1_outputs[5512] = layer0_outputs[12255];
    assign layer1_outputs[5513] = ~(layer0_outputs[2731]);
    assign layer1_outputs[5514] = ~(layer0_outputs[11811]) | (layer0_outputs[3588]);
    assign layer1_outputs[5515] = layer0_outputs[12354];
    assign layer1_outputs[5516] = layer0_outputs[7420];
    assign layer1_outputs[5517] = layer0_outputs[10047];
    assign layer1_outputs[5518] = ~(layer0_outputs[5858]) | (layer0_outputs[4609]);
    assign layer1_outputs[5519] = (layer0_outputs[12457]) & (layer0_outputs[10236]);
    assign layer1_outputs[5520] = (layer0_outputs[3086]) | (layer0_outputs[911]);
    assign layer1_outputs[5521] = (layer0_outputs[9546]) & ~(layer0_outputs[6116]);
    assign layer1_outputs[5522] = ~((layer0_outputs[4839]) | (layer0_outputs[746]));
    assign layer1_outputs[5523] = (layer0_outputs[1226]) | (layer0_outputs[6292]);
    assign layer1_outputs[5524] = ~((layer0_outputs[8248]) ^ (layer0_outputs[7958]));
    assign layer1_outputs[5525] = ~(layer0_outputs[6822]);
    assign layer1_outputs[5526] = layer0_outputs[8488];
    assign layer1_outputs[5527] = ~((layer0_outputs[6513]) & (layer0_outputs[5672]));
    assign layer1_outputs[5528] = layer0_outputs[12322];
    assign layer1_outputs[5529] = layer0_outputs[4566];
    assign layer1_outputs[5530] = (layer0_outputs[4206]) | (layer0_outputs[5526]);
    assign layer1_outputs[5531] = layer0_outputs[5556];
    assign layer1_outputs[5532] = ~(layer0_outputs[11741]);
    assign layer1_outputs[5533] = (layer0_outputs[12410]) | (layer0_outputs[8045]);
    assign layer1_outputs[5534] = ~(layer0_outputs[10699]);
    assign layer1_outputs[5535] = ~(layer0_outputs[9509]);
    assign layer1_outputs[5536] = (layer0_outputs[8136]) ^ (layer0_outputs[1603]);
    assign layer1_outputs[5537] = layer0_outputs[3438];
    assign layer1_outputs[5538] = (layer0_outputs[8356]) & ~(layer0_outputs[3148]);
    assign layer1_outputs[5539] = ~(layer0_outputs[7408]);
    assign layer1_outputs[5540] = (layer0_outputs[12412]) & ~(layer0_outputs[1245]);
    assign layer1_outputs[5541] = layer0_outputs[7400];
    assign layer1_outputs[5542] = ~(layer0_outputs[3314]);
    assign layer1_outputs[5543] = 1'b1;
    assign layer1_outputs[5544] = (layer0_outputs[1581]) ^ (layer0_outputs[6591]);
    assign layer1_outputs[5545] = ~(layer0_outputs[7090]);
    assign layer1_outputs[5546] = layer0_outputs[3341];
    assign layer1_outputs[5547] = (layer0_outputs[8438]) | (layer0_outputs[5527]);
    assign layer1_outputs[5548] = layer0_outputs[1327];
    assign layer1_outputs[5549] = (layer0_outputs[5348]) ^ (layer0_outputs[1881]);
    assign layer1_outputs[5550] = ~(layer0_outputs[5186]);
    assign layer1_outputs[5551] = ~((layer0_outputs[2478]) | (layer0_outputs[11479]));
    assign layer1_outputs[5552] = ~((layer0_outputs[2498]) & (layer0_outputs[1163]));
    assign layer1_outputs[5553] = 1'b0;
    assign layer1_outputs[5554] = (layer0_outputs[8508]) | (layer0_outputs[1150]);
    assign layer1_outputs[5555] = ~((layer0_outputs[12090]) & (layer0_outputs[764]));
    assign layer1_outputs[5556] = ~((layer0_outputs[10916]) & (layer0_outputs[5323]));
    assign layer1_outputs[5557] = 1'b1;
    assign layer1_outputs[5558] = ~(layer0_outputs[10229]);
    assign layer1_outputs[5559] = ~(layer0_outputs[1062]) | (layer0_outputs[11363]);
    assign layer1_outputs[5560] = layer0_outputs[6146];
    assign layer1_outputs[5561] = ~(layer0_outputs[11620]) | (layer0_outputs[3167]);
    assign layer1_outputs[5562] = ~(layer0_outputs[2866]) | (layer0_outputs[12233]);
    assign layer1_outputs[5563] = layer0_outputs[7500];
    assign layer1_outputs[5564] = (layer0_outputs[11848]) & ~(layer0_outputs[8381]);
    assign layer1_outputs[5565] = ~((layer0_outputs[383]) | (layer0_outputs[10698]));
    assign layer1_outputs[5566] = (layer0_outputs[6321]) & (layer0_outputs[12190]);
    assign layer1_outputs[5567] = ~((layer0_outputs[8014]) ^ (layer0_outputs[8347]));
    assign layer1_outputs[5568] = (layer0_outputs[6744]) & ~(layer0_outputs[11076]);
    assign layer1_outputs[5569] = ~(layer0_outputs[8408]) | (layer0_outputs[8129]);
    assign layer1_outputs[5570] = ~(layer0_outputs[768]);
    assign layer1_outputs[5571] = ~((layer0_outputs[11269]) & (layer0_outputs[12546]));
    assign layer1_outputs[5572] = ~((layer0_outputs[12689]) & (layer0_outputs[3702]));
    assign layer1_outputs[5573] = ~(layer0_outputs[12131]);
    assign layer1_outputs[5574] = (layer0_outputs[5266]) & (layer0_outputs[10407]);
    assign layer1_outputs[5575] = (layer0_outputs[10428]) | (layer0_outputs[2949]);
    assign layer1_outputs[5576] = layer0_outputs[7565];
    assign layer1_outputs[5577] = ~((layer0_outputs[6499]) ^ (layer0_outputs[784]));
    assign layer1_outputs[5578] = layer0_outputs[11477];
    assign layer1_outputs[5579] = ~((layer0_outputs[8822]) | (layer0_outputs[4252]));
    assign layer1_outputs[5580] = ~(layer0_outputs[10368]) | (layer0_outputs[12325]);
    assign layer1_outputs[5581] = layer0_outputs[5676];
    assign layer1_outputs[5582] = ~(layer0_outputs[6752]) | (layer0_outputs[7035]);
    assign layer1_outputs[5583] = layer0_outputs[12237];
    assign layer1_outputs[5584] = ~(layer0_outputs[11603]);
    assign layer1_outputs[5585] = 1'b1;
    assign layer1_outputs[5586] = (layer0_outputs[12381]) & ~(layer0_outputs[11843]);
    assign layer1_outputs[5587] = ~((layer0_outputs[11450]) & (layer0_outputs[1380]));
    assign layer1_outputs[5588] = layer0_outputs[5060];
    assign layer1_outputs[5589] = ~(layer0_outputs[105]);
    assign layer1_outputs[5590] = layer0_outputs[12777];
    assign layer1_outputs[5591] = layer0_outputs[8746];
    assign layer1_outputs[5592] = 1'b1;
    assign layer1_outputs[5593] = (layer0_outputs[4939]) ^ (layer0_outputs[8020]);
    assign layer1_outputs[5594] = ~(layer0_outputs[11602]);
    assign layer1_outputs[5595] = (layer0_outputs[11099]) | (layer0_outputs[9193]);
    assign layer1_outputs[5596] = ~(layer0_outputs[12783]) | (layer0_outputs[8628]);
    assign layer1_outputs[5597] = layer0_outputs[3377];
    assign layer1_outputs[5598] = layer0_outputs[7488];
    assign layer1_outputs[5599] = (layer0_outputs[104]) ^ (layer0_outputs[8003]);
    assign layer1_outputs[5600] = ~(layer0_outputs[4650]);
    assign layer1_outputs[5601] = ~((layer0_outputs[6504]) & (layer0_outputs[5588]));
    assign layer1_outputs[5602] = layer0_outputs[2775];
    assign layer1_outputs[5603] = ~(layer0_outputs[12368]);
    assign layer1_outputs[5604] = (layer0_outputs[5030]) & (layer0_outputs[3546]);
    assign layer1_outputs[5605] = ~(layer0_outputs[1577]);
    assign layer1_outputs[5606] = layer0_outputs[10012];
    assign layer1_outputs[5607] = layer0_outputs[1204];
    assign layer1_outputs[5608] = ~((layer0_outputs[8446]) ^ (layer0_outputs[6441]));
    assign layer1_outputs[5609] = layer0_outputs[6227];
    assign layer1_outputs[5610] = ~(layer0_outputs[11179]);
    assign layer1_outputs[5611] = 1'b1;
    assign layer1_outputs[5612] = (layer0_outputs[6977]) & ~(layer0_outputs[1929]);
    assign layer1_outputs[5613] = ~(layer0_outputs[9866]) | (layer0_outputs[1199]);
    assign layer1_outputs[5614] = (layer0_outputs[6083]) & (layer0_outputs[7071]);
    assign layer1_outputs[5615] = 1'b1;
    assign layer1_outputs[5616] = ~(layer0_outputs[3666]) | (layer0_outputs[4707]);
    assign layer1_outputs[5617] = layer0_outputs[3415];
    assign layer1_outputs[5618] = ~((layer0_outputs[3]) ^ (layer0_outputs[1104]));
    assign layer1_outputs[5619] = layer0_outputs[7099];
    assign layer1_outputs[5620] = layer0_outputs[11168];
    assign layer1_outputs[5621] = (layer0_outputs[3575]) | (layer0_outputs[2912]);
    assign layer1_outputs[5622] = layer0_outputs[10630];
    assign layer1_outputs[5623] = 1'b0;
    assign layer1_outputs[5624] = (layer0_outputs[1266]) & ~(layer0_outputs[1916]);
    assign layer1_outputs[5625] = ~((layer0_outputs[4346]) | (layer0_outputs[8958]));
    assign layer1_outputs[5626] = ~(layer0_outputs[10839]) | (layer0_outputs[9116]);
    assign layer1_outputs[5627] = ~(layer0_outputs[7205]);
    assign layer1_outputs[5628] = ~((layer0_outputs[5304]) ^ (layer0_outputs[7874]));
    assign layer1_outputs[5629] = layer0_outputs[9060];
    assign layer1_outputs[5630] = ~((layer0_outputs[4123]) | (layer0_outputs[12729]));
    assign layer1_outputs[5631] = layer0_outputs[3579];
    assign layer1_outputs[5632] = (layer0_outputs[9189]) ^ (layer0_outputs[219]);
    assign layer1_outputs[5633] = ~(layer0_outputs[5463]);
    assign layer1_outputs[5634] = layer0_outputs[9430];
    assign layer1_outputs[5635] = ~((layer0_outputs[9071]) | (layer0_outputs[11714]));
    assign layer1_outputs[5636] = layer0_outputs[2024];
    assign layer1_outputs[5637] = ~(layer0_outputs[10175]);
    assign layer1_outputs[5638] = ~(layer0_outputs[3849]);
    assign layer1_outputs[5639] = ~(layer0_outputs[6773]) | (layer0_outputs[6191]);
    assign layer1_outputs[5640] = layer0_outputs[11718];
    assign layer1_outputs[5641] = ~((layer0_outputs[312]) ^ (layer0_outputs[2978]));
    assign layer1_outputs[5642] = ~(layer0_outputs[7704]) | (layer0_outputs[4847]);
    assign layer1_outputs[5643] = ~(layer0_outputs[2920]) | (layer0_outputs[617]);
    assign layer1_outputs[5644] = ~(layer0_outputs[3551]) | (layer0_outputs[11465]);
    assign layer1_outputs[5645] = (layer0_outputs[1518]) & ~(layer0_outputs[3107]);
    assign layer1_outputs[5646] = ~(layer0_outputs[12115]);
    assign layer1_outputs[5647] = ~(layer0_outputs[9095]);
    assign layer1_outputs[5648] = (layer0_outputs[7196]) & ~(layer0_outputs[5647]);
    assign layer1_outputs[5649] = layer0_outputs[5473];
    assign layer1_outputs[5650] = ~(layer0_outputs[1370]);
    assign layer1_outputs[5651] = (layer0_outputs[3853]) | (layer0_outputs[4522]);
    assign layer1_outputs[5652] = (layer0_outputs[10031]) ^ (layer0_outputs[2827]);
    assign layer1_outputs[5653] = ~(layer0_outputs[1261]);
    assign layer1_outputs[5654] = ~((layer0_outputs[11669]) ^ (layer0_outputs[11894]));
    assign layer1_outputs[5655] = ~((layer0_outputs[1882]) & (layer0_outputs[2663]));
    assign layer1_outputs[5656] = ~(layer0_outputs[9387]);
    assign layer1_outputs[5657] = ~((layer0_outputs[2859]) ^ (layer0_outputs[8027]));
    assign layer1_outputs[5658] = 1'b0;
    assign layer1_outputs[5659] = 1'b1;
    assign layer1_outputs[5660] = ~(layer0_outputs[12716]) | (layer0_outputs[2164]);
    assign layer1_outputs[5661] = ~((layer0_outputs[2080]) | (layer0_outputs[3725]));
    assign layer1_outputs[5662] = ~(layer0_outputs[6398]);
    assign layer1_outputs[5663] = ~(layer0_outputs[3791]) | (layer0_outputs[2893]);
    assign layer1_outputs[5664] = (layer0_outputs[7680]) & ~(layer0_outputs[9623]);
    assign layer1_outputs[5665] = layer0_outputs[11921];
    assign layer1_outputs[5666] = (layer0_outputs[9733]) & (layer0_outputs[4173]);
    assign layer1_outputs[5667] = ~(layer0_outputs[5324]);
    assign layer1_outputs[5668] = layer0_outputs[129];
    assign layer1_outputs[5669] = layer0_outputs[4042];
    assign layer1_outputs[5670] = ~(layer0_outputs[8157]) | (layer0_outputs[6694]);
    assign layer1_outputs[5671] = layer0_outputs[4945];
    assign layer1_outputs[5672] = layer0_outputs[4474];
    assign layer1_outputs[5673] = layer0_outputs[2371];
    assign layer1_outputs[5674] = (layer0_outputs[4391]) & ~(layer0_outputs[6823]);
    assign layer1_outputs[5675] = (layer0_outputs[10813]) & (layer0_outputs[9134]);
    assign layer1_outputs[5676] = ~((layer0_outputs[8062]) ^ (layer0_outputs[6468]));
    assign layer1_outputs[5677] = ~((layer0_outputs[4780]) & (layer0_outputs[5148]));
    assign layer1_outputs[5678] = layer0_outputs[1839];
    assign layer1_outputs[5679] = (layer0_outputs[5685]) ^ (layer0_outputs[9394]);
    assign layer1_outputs[5680] = ~((layer0_outputs[4705]) ^ (layer0_outputs[12655]));
    assign layer1_outputs[5681] = (layer0_outputs[9823]) | (layer0_outputs[2819]);
    assign layer1_outputs[5682] = ~(layer0_outputs[364]);
    assign layer1_outputs[5683] = ~(layer0_outputs[7333]);
    assign layer1_outputs[5684] = ~(layer0_outputs[9584]);
    assign layer1_outputs[5685] = ~((layer0_outputs[4168]) | (layer0_outputs[4392]));
    assign layer1_outputs[5686] = layer0_outputs[8491];
    assign layer1_outputs[5687] = ~(layer0_outputs[3343]);
    assign layer1_outputs[5688] = layer0_outputs[479];
    assign layer1_outputs[5689] = layer0_outputs[11593];
    assign layer1_outputs[5690] = layer0_outputs[3504];
    assign layer1_outputs[5691] = (layer0_outputs[9656]) & ~(layer0_outputs[3040]);
    assign layer1_outputs[5692] = layer0_outputs[10787];
    assign layer1_outputs[5693] = 1'b0;
    assign layer1_outputs[5694] = ~(layer0_outputs[6876]) | (layer0_outputs[7516]);
    assign layer1_outputs[5695] = (layer0_outputs[9174]) & ~(layer0_outputs[6585]);
    assign layer1_outputs[5696] = layer0_outputs[9691];
    assign layer1_outputs[5697] = ~(layer0_outputs[3670]);
    assign layer1_outputs[5698] = ~((layer0_outputs[6669]) ^ (layer0_outputs[5279]));
    assign layer1_outputs[5699] = ~((layer0_outputs[1664]) | (layer0_outputs[5603]));
    assign layer1_outputs[5700] = layer0_outputs[9445];
    assign layer1_outputs[5701] = ~(layer0_outputs[5982]) | (layer0_outputs[10460]);
    assign layer1_outputs[5702] = layer0_outputs[4121];
    assign layer1_outputs[5703] = ~((layer0_outputs[4559]) & (layer0_outputs[8517]));
    assign layer1_outputs[5704] = ~((layer0_outputs[2705]) ^ (layer0_outputs[8086]));
    assign layer1_outputs[5705] = ~(layer0_outputs[1740]);
    assign layer1_outputs[5706] = layer0_outputs[1353];
    assign layer1_outputs[5707] = layer0_outputs[4544];
    assign layer1_outputs[5708] = ~((layer0_outputs[10779]) ^ (layer0_outputs[5522]));
    assign layer1_outputs[5709] = layer0_outputs[3911];
    assign layer1_outputs[5710] = (layer0_outputs[3097]) & ~(layer0_outputs[11711]);
    assign layer1_outputs[5711] = ~(layer0_outputs[2512]);
    assign layer1_outputs[5712] = ~((layer0_outputs[7603]) & (layer0_outputs[11417]));
    assign layer1_outputs[5713] = ~((layer0_outputs[7229]) ^ (layer0_outputs[8016]));
    assign layer1_outputs[5714] = ~(layer0_outputs[1345]);
    assign layer1_outputs[5715] = (layer0_outputs[4596]) & ~(layer0_outputs[10306]);
    assign layer1_outputs[5716] = ~((layer0_outputs[12796]) ^ (layer0_outputs[7445]));
    assign layer1_outputs[5717] = layer0_outputs[9554];
    assign layer1_outputs[5718] = layer0_outputs[9329];
    assign layer1_outputs[5719] = (layer0_outputs[4807]) | (layer0_outputs[5726]);
    assign layer1_outputs[5720] = ~(layer0_outputs[3067]);
    assign layer1_outputs[5721] = ~(layer0_outputs[8300]);
    assign layer1_outputs[5722] = ~(layer0_outputs[2076]);
    assign layer1_outputs[5723] = ~(layer0_outputs[3069]);
    assign layer1_outputs[5724] = ~((layer0_outputs[2047]) ^ (layer0_outputs[10759]));
    assign layer1_outputs[5725] = ~((layer0_outputs[7442]) ^ (layer0_outputs[1591]));
    assign layer1_outputs[5726] = 1'b1;
    assign layer1_outputs[5727] = layer0_outputs[5339];
    assign layer1_outputs[5728] = ~((layer0_outputs[6689]) ^ (layer0_outputs[3061]));
    assign layer1_outputs[5729] = (layer0_outputs[7387]) | (layer0_outputs[3776]);
    assign layer1_outputs[5730] = ~(layer0_outputs[4135]);
    assign layer1_outputs[5731] = ~(layer0_outputs[12072]) | (layer0_outputs[3543]);
    assign layer1_outputs[5732] = ~((layer0_outputs[12668]) | (layer0_outputs[12553]));
    assign layer1_outputs[5733] = layer0_outputs[11918];
    assign layer1_outputs[5734] = ~((layer0_outputs[6736]) & (layer0_outputs[6135]));
    assign layer1_outputs[5735] = ~(layer0_outputs[5550]);
    assign layer1_outputs[5736] = (layer0_outputs[9600]) & ~(layer0_outputs[7513]);
    assign layer1_outputs[5737] = (layer0_outputs[10104]) & ~(layer0_outputs[7763]);
    assign layer1_outputs[5738] = ~(layer0_outputs[8911]) | (layer0_outputs[1540]);
    assign layer1_outputs[5739] = layer0_outputs[10696];
    assign layer1_outputs[5740] = ~(layer0_outputs[3590]);
    assign layer1_outputs[5741] = ~(layer0_outputs[3348]);
    assign layer1_outputs[5742] = ~(layer0_outputs[2443]);
    assign layer1_outputs[5743] = (layer0_outputs[7307]) | (layer0_outputs[11978]);
    assign layer1_outputs[5744] = (layer0_outputs[3424]) ^ (layer0_outputs[9589]);
    assign layer1_outputs[5745] = ~(layer0_outputs[7304]);
    assign layer1_outputs[5746] = (layer0_outputs[3655]) & ~(layer0_outputs[12793]);
    assign layer1_outputs[5747] = layer0_outputs[11013];
    assign layer1_outputs[5748] = 1'b0;
    assign layer1_outputs[5749] = ~(layer0_outputs[2223]);
    assign layer1_outputs[5750] = (layer0_outputs[767]) ^ (layer0_outputs[8691]);
    assign layer1_outputs[5751] = (layer0_outputs[2879]) ^ (layer0_outputs[2017]);
    assign layer1_outputs[5752] = ~(layer0_outputs[5322]) | (layer0_outputs[9525]);
    assign layer1_outputs[5753] = layer0_outputs[1644];
    assign layer1_outputs[5754] = layer0_outputs[9183];
    assign layer1_outputs[5755] = ~((layer0_outputs[1637]) | (layer0_outputs[7846]));
    assign layer1_outputs[5756] = ~(layer0_outputs[4923]) | (layer0_outputs[8980]);
    assign layer1_outputs[5757] = ~((layer0_outputs[1189]) ^ (layer0_outputs[6223]));
    assign layer1_outputs[5758] = (layer0_outputs[9254]) | (layer0_outputs[1888]);
    assign layer1_outputs[5759] = ~((layer0_outputs[2875]) & (layer0_outputs[6640]));
    assign layer1_outputs[5760] = ~((layer0_outputs[5913]) & (layer0_outputs[3100]));
    assign layer1_outputs[5761] = (layer0_outputs[460]) & (layer0_outputs[10492]);
    assign layer1_outputs[5762] = ~((layer0_outputs[690]) | (layer0_outputs[7924]));
    assign layer1_outputs[5763] = (layer0_outputs[10647]) & (layer0_outputs[10427]);
    assign layer1_outputs[5764] = (layer0_outputs[744]) | (layer0_outputs[468]);
    assign layer1_outputs[5765] = (layer0_outputs[6786]) ^ (layer0_outputs[8792]);
    assign layer1_outputs[5766] = layer0_outputs[2865];
    assign layer1_outputs[5767] = (layer0_outputs[10211]) ^ (layer0_outputs[5339]);
    assign layer1_outputs[5768] = ~((layer0_outputs[8393]) ^ (layer0_outputs[5821]));
    assign layer1_outputs[5769] = 1'b0;
    assign layer1_outputs[5770] = (layer0_outputs[12069]) | (layer0_outputs[12442]);
    assign layer1_outputs[5771] = layer0_outputs[5000];
    assign layer1_outputs[5772] = layer0_outputs[5239];
    assign layer1_outputs[5773] = ~(layer0_outputs[8187]);
    assign layer1_outputs[5774] = 1'b0;
    assign layer1_outputs[5775] = ~((layer0_outputs[10181]) ^ (layer0_outputs[3260]));
    assign layer1_outputs[5776] = layer0_outputs[4383];
    assign layer1_outputs[5777] = ~(layer0_outputs[2447]) | (layer0_outputs[9282]);
    assign layer1_outputs[5778] = (layer0_outputs[991]) | (layer0_outputs[1201]);
    assign layer1_outputs[5779] = ~(layer0_outputs[8422]);
    assign layer1_outputs[5780] = ~(layer0_outputs[6606]) | (layer0_outputs[12193]);
    assign layer1_outputs[5781] = 1'b1;
    assign layer1_outputs[5782] = (layer0_outputs[11221]) & ~(layer0_outputs[7567]);
    assign layer1_outputs[5783] = ~(layer0_outputs[3548]);
    assign layer1_outputs[5784] = 1'b0;
    assign layer1_outputs[5785] = (layer0_outputs[4803]) & ~(layer0_outputs[8565]);
    assign layer1_outputs[5786] = layer0_outputs[6035];
    assign layer1_outputs[5787] = ~(layer0_outputs[650]);
    assign layer1_outputs[5788] = (layer0_outputs[12594]) | (layer0_outputs[5174]);
    assign layer1_outputs[5789] = (layer0_outputs[4467]) & (layer0_outputs[7337]);
    assign layer1_outputs[5790] = layer0_outputs[6365];
    assign layer1_outputs[5791] = ~((layer0_outputs[1554]) & (layer0_outputs[4501]));
    assign layer1_outputs[5792] = ~(layer0_outputs[1588]);
    assign layer1_outputs[5793] = (layer0_outputs[12610]) & (layer0_outputs[3681]);
    assign layer1_outputs[5794] = layer0_outputs[9127];
    assign layer1_outputs[5795] = ~(layer0_outputs[2544]);
    assign layer1_outputs[5796] = (layer0_outputs[11286]) & ~(layer0_outputs[1855]);
    assign layer1_outputs[5797] = layer0_outputs[417];
    assign layer1_outputs[5798] = ~(layer0_outputs[8720]);
    assign layer1_outputs[5799] = (layer0_outputs[12608]) & ~(layer0_outputs[245]);
    assign layer1_outputs[5800] = (layer0_outputs[12460]) ^ (layer0_outputs[575]);
    assign layer1_outputs[5801] = ~(layer0_outputs[2548]) | (layer0_outputs[8632]);
    assign layer1_outputs[5802] = ~(layer0_outputs[242]);
    assign layer1_outputs[5803] = ~(layer0_outputs[2781]);
    assign layer1_outputs[5804] = (layer0_outputs[12416]) & ~(layer0_outputs[9794]);
    assign layer1_outputs[5805] = (layer0_outputs[9149]) & (layer0_outputs[597]);
    assign layer1_outputs[5806] = (layer0_outputs[8489]) & ~(layer0_outputs[1085]);
    assign layer1_outputs[5807] = ~(layer0_outputs[7805]) | (layer0_outputs[2937]);
    assign layer1_outputs[5808] = (layer0_outputs[11868]) ^ (layer0_outputs[601]);
    assign layer1_outputs[5809] = ~((layer0_outputs[7613]) ^ (layer0_outputs[10694]));
    assign layer1_outputs[5810] = ~(layer0_outputs[2549]) | (layer0_outputs[2194]);
    assign layer1_outputs[5811] = ~(layer0_outputs[9764]) | (layer0_outputs[1412]);
    assign layer1_outputs[5812] = ~((layer0_outputs[12131]) | (layer0_outputs[9409]));
    assign layer1_outputs[5813] = (layer0_outputs[8614]) & (layer0_outputs[11729]);
    assign layer1_outputs[5814] = ~(layer0_outputs[2604]);
    assign layer1_outputs[5815] = (layer0_outputs[4570]) & ~(layer0_outputs[9315]);
    assign layer1_outputs[5816] = ~(layer0_outputs[4315]) | (layer0_outputs[8645]);
    assign layer1_outputs[5817] = ~(layer0_outputs[5058]);
    assign layer1_outputs[5818] = ~(layer0_outputs[3120]) | (layer0_outputs[8627]);
    assign layer1_outputs[5819] = ~(layer0_outputs[8102]);
    assign layer1_outputs[5820] = layer0_outputs[2544];
    assign layer1_outputs[5821] = ~(layer0_outputs[12261]);
    assign layer1_outputs[5822] = (layer0_outputs[4809]) & (layer0_outputs[3336]);
    assign layer1_outputs[5823] = ~(layer0_outputs[6735]);
    assign layer1_outputs[5824] = ~(layer0_outputs[12433]);
    assign layer1_outputs[5825] = (layer0_outputs[11533]) ^ (layer0_outputs[9239]);
    assign layer1_outputs[5826] = 1'b0;
    assign layer1_outputs[5827] = ~((layer0_outputs[1502]) ^ (layer0_outputs[5331]));
    assign layer1_outputs[5828] = (layer0_outputs[95]) & (layer0_outputs[5190]);
    assign layer1_outputs[5829] = layer0_outputs[432];
    assign layer1_outputs[5830] = 1'b0;
    assign layer1_outputs[5831] = ~(layer0_outputs[10642]) | (layer0_outputs[12029]);
    assign layer1_outputs[5832] = ~(layer0_outputs[7409]) | (layer0_outputs[4770]);
    assign layer1_outputs[5833] = layer0_outputs[9427];
    assign layer1_outputs[5834] = layer0_outputs[1480];
    assign layer1_outputs[5835] = (layer0_outputs[11777]) & ~(layer0_outputs[1531]);
    assign layer1_outputs[5836] = ~(layer0_outputs[2051]);
    assign layer1_outputs[5837] = (layer0_outputs[9400]) ^ (layer0_outputs[2401]);
    assign layer1_outputs[5838] = ~(layer0_outputs[1912]);
    assign layer1_outputs[5839] = ~(layer0_outputs[9800]) | (layer0_outputs[4475]);
    assign layer1_outputs[5840] = ~(layer0_outputs[12077]);
    assign layer1_outputs[5841] = layer0_outputs[5465];
    assign layer1_outputs[5842] = ~((layer0_outputs[8712]) | (layer0_outputs[7230]));
    assign layer1_outputs[5843] = (layer0_outputs[10554]) & ~(layer0_outputs[2232]);
    assign layer1_outputs[5844] = layer0_outputs[4518];
    assign layer1_outputs[5845] = ~((layer0_outputs[11933]) & (layer0_outputs[2826]));
    assign layer1_outputs[5846] = (layer0_outputs[6434]) & ~(layer0_outputs[5320]);
    assign layer1_outputs[5847] = ~((layer0_outputs[11957]) ^ (layer0_outputs[11542]));
    assign layer1_outputs[5848] = ~((layer0_outputs[11624]) | (layer0_outputs[8596]));
    assign layer1_outputs[5849] = 1'b1;
    assign layer1_outputs[5850] = ~(layer0_outputs[12317]) | (layer0_outputs[12424]);
    assign layer1_outputs[5851] = ~(layer0_outputs[3382]);
    assign layer1_outputs[5852] = (layer0_outputs[4643]) & ~(layer0_outputs[10978]);
    assign layer1_outputs[5853] = (layer0_outputs[3034]) & ~(layer0_outputs[5615]);
    assign layer1_outputs[5854] = (layer0_outputs[3647]) & ~(layer0_outputs[9474]);
    assign layer1_outputs[5855] = layer0_outputs[4532];
    assign layer1_outputs[5856] = layer0_outputs[11894];
    assign layer1_outputs[5857] = ~((layer0_outputs[6242]) ^ (layer0_outputs[6721]));
    assign layer1_outputs[5858] = ~((layer0_outputs[6339]) ^ (layer0_outputs[5422]));
    assign layer1_outputs[5859] = (layer0_outputs[192]) | (layer0_outputs[9033]);
    assign layer1_outputs[5860] = ~(layer0_outputs[11212]);
    assign layer1_outputs[5861] = ~(layer0_outputs[9188]);
    assign layer1_outputs[5862] = (layer0_outputs[5928]) & ~(layer0_outputs[1746]);
    assign layer1_outputs[5863] = (layer0_outputs[8808]) & ~(layer0_outputs[6267]);
    assign layer1_outputs[5864] = ~(layer0_outputs[2310]);
    assign layer1_outputs[5865] = (layer0_outputs[8232]) & (layer0_outputs[7943]);
    assign layer1_outputs[5866] = (layer0_outputs[7058]) & (layer0_outputs[1113]);
    assign layer1_outputs[5867] = ~(layer0_outputs[6494]);
    assign layer1_outputs[5868] = layer0_outputs[6283];
    assign layer1_outputs[5869] = ~(layer0_outputs[3307]);
    assign layer1_outputs[5870] = (layer0_outputs[595]) | (layer0_outputs[7624]);
    assign layer1_outputs[5871] = layer0_outputs[8514];
    assign layer1_outputs[5872] = layer0_outputs[5509];
    assign layer1_outputs[5873] = ~(layer0_outputs[2657]);
    assign layer1_outputs[5874] = ~(layer0_outputs[6409]);
    assign layer1_outputs[5875] = (layer0_outputs[12259]) & ~(layer0_outputs[9883]);
    assign layer1_outputs[5876] = layer0_outputs[3754];
    assign layer1_outputs[5877] = ~((layer0_outputs[7343]) | (layer0_outputs[11835]));
    assign layer1_outputs[5878] = ~(layer0_outputs[12398]);
    assign layer1_outputs[5879] = (layer0_outputs[11032]) ^ (layer0_outputs[8410]);
    assign layer1_outputs[5880] = ~(layer0_outputs[10936]);
    assign layer1_outputs[5881] = layer0_outputs[7269];
    assign layer1_outputs[5882] = ~(layer0_outputs[1618]);
    assign layer1_outputs[5883] = (layer0_outputs[544]) | (layer0_outputs[9755]);
    assign layer1_outputs[5884] = ~(layer0_outputs[6570]);
    assign layer1_outputs[5885] = ~(layer0_outputs[10763]);
    assign layer1_outputs[5886] = layer0_outputs[8211];
    assign layer1_outputs[5887] = ~((layer0_outputs[3925]) | (layer0_outputs[2536]));
    assign layer1_outputs[5888] = (layer0_outputs[8402]) & ~(layer0_outputs[1988]);
    assign layer1_outputs[5889] = 1'b0;
    assign layer1_outputs[5890] = ~((layer0_outputs[147]) & (layer0_outputs[11632]));
    assign layer1_outputs[5891] = (layer0_outputs[12157]) & ~(layer0_outputs[12068]);
    assign layer1_outputs[5892] = (layer0_outputs[9115]) ^ (layer0_outputs[5362]);
    assign layer1_outputs[5893] = layer0_outputs[11086];
    assign layer1_outputs[5894] = (layer0_outputs[12169]) | (layer0_outputs[1941]);
    assign layer1_outputs[5895] = ~(layer0_outputs[3903]) | (layer0_outputs[5132]);
    assign layer1_outputs[5896] = layer0_outputs[10659];
    assign layer1_outputs[5897] = (layer0_outputs[75]) & (layer0_outputs[8792]);
    assign layer1_outputs[5898] = layer0_outputs[3632];
    assign layer1_outputs[5899] = ~(layer0_outputs[7129]) | (layer0_outputs[8695]);
    assign layer1_outputs[5900] = ~(layer0_outputs[9618]);
    assign layer1_outputs[5901] = ~((layer0_outputs[5475]) ^ (layer0_outputs[4479]));
    assign layer1_outputs[5902] = ~((layer0_outputs[4990]) | (layer0_outputs[11645]));
    assign layer1_outputs[5903] = ~(layer0_outputs[10098]);
    assign layer1_outputs[5904] = (layer0_outputs[67]) & ~(layer0_outputs[2951]);
    assign layer1_outputs[5905] = ~(layer0_outputs[12177]);
    assign layer1_outputs[5906] = ~(layer0_outputs[130]);
    assign layer1_outputs[5907] = ~(layer0_outputs[2698]);
    assign layer1_outputs[5908] = ~(layer0_outputs[1635]) | (layer0_outputs[2119]);
    assign layer1_outputs[5909] = layer0_outputs[4346];
    assign layer1_outputs[5910] = ~(layer0_outputs[4095]);
    assign layer1_outputs[5911] = (layer0_outputs[5234]) & ~(layer0_outputs[12369]);
    assign layer1_outputs[5912] = ~(layer0_outputs[8924]) | (layer0_outputs[9334]);
    assign layer1_outputs[5913] = (layer0_outputs[957]) & (layer0_outputs[12014]);
    assign layer1_outputs[5914] = ~(layer0_outputs[5334]);
    assign layer1_outputs[5915] = (layer0_outputs[5782]) | (layer0_outputs[5707]);
    assign layer1_outputs[5916] = ~(layer0_outputs[1358]);
    assign layer1_outputs[5917] = (layer0_outputs[10363]) & ~(layer0_outputs[7254]);
    assign layer1_outputs[5918] = ~(layer0_outputs[1724]);
    assign layer1_outputs[5919] = (layer0_outputs[1573]) ^ (layer0_outputs[4691]);
    assign layer1_outputs[5920] = (layer0_outputs[5473]) & (layer0_outputs[7972]);
    assign layer1_outputs[5921] = ~(layer0_outputs[4937]);
    assign layer1_outputs[5922] = ~(layer0_outputs[7341]) | (layer0_outputs[4729]);
    assign layer1_outputs[5923] = (layer0_outputs[10571]) | (layer0_outputs[9607]);
    assign layer1_outputs[5924] = layer0_outputs[565];
    assign layer1_outputs[5925] = ~((layer0_outputs[12065]) ^ (layer0_outputs[9207]));
    assign layer1_outputs[5926] = ~(layer0_outputs[4287]);
    assign layer1_outputs[5927] = ~(layer0_outputs[5539]);
    assign layer1_outputs[5928] = (layer0_outputs[10623]) & ~(layer0_outputs[7988]);
    assign layer1_outputs[5929] = ~(layer0_outputs[2467]) | (layer0_outputs[7815]);
    assign layer1_outputs[5930] = layer0_outputs[6965];
    assign layer1_outputs[5931] = ~((layer0_outputs[9869]) | (layer0_outputs[5934]));
    assign layer1_outputs[5932] = layer0_outputs[19];
    assign layer1_outputs[5933] = ~((layer0_outputs[3767]) & (layer0_outputs[1567]));
    assign layer1_outputs[5934] = ~((layer0_outputs[10317]) & (layer0_outputs[10615]));
    assign layer1_outputs[5935] = ~((layer0_outputs[4590]) & (layer0_outputs[6829]));
    assign layer1_outputs[5936] = ~(layer0_outputs[12045]);
    assign layer1_outputs[5937] = ~(layer0_outputs[9044]);
    assign layer1_outputs[5938] = ~(layer0_outputs[8013]) | (layer0_outputs[8547]);
    assign layer1_outputs[5939] = (layer0_outputs[9289]) & ~(layer0_outputs[5817]);
    assign layer1_outputs[5940] = ~((layer0_outputs[2307]) ^ (layer0_outputs[12617]));
    assign layer1_outputs[5941] = layer0_outputs[5829];
    assign layer1_outputs[5942] = (layer0_outputs[7096]) ^ (layer0_outputs[10547]);
    assign layer1_outputs[5943] = ~((layer0_outputs[8748]) ^ (layer0_outputs[5051]));
    assign layer1_outputs[5944] = ~(layer0_outputs[4575]);
    assign layer1_outputs[5945] = ~(layer0_outputs[8854]) | (layer0_outputs[4759]);
    assign layer1_outputs[5946] = layer0_outputs[5179];
    assign layer1_outputs[5947] = layer0_outputs[5708];
    assign layer1_outputs[5948] = (layer0_outputs[6643]) | (layer0_outputs[5981]);
    assign layer1_outputs[5949] = (layer0_outputs[5384]) & (layer0_outputs[297]);
    assign layer1_outputs[5950] = (layer0_outputs[8527]) & (layer0_outputs[10769]);
    assign layer1_outputs[5951] = ~(layer0_outputs[4668]);
    assign layer1_outputs[5952] = layer0_outputs[3118];
    assign layer1_outputs[5953] = ~(layer0_outputs[4306]);
    assign layer1_outputs[5954] = layer0_outputs[11482];
    assign layer1_outputs[5955] = ~(layer0_outputs[4202]);
    assign layer1_outputs[5956] = ~(layer0_outputs[6977]);
    assign layer1_outputs[5957] = (layer0_outputs[8318]) ^ (layer0_outputs[380]);
    assign layer1_outputs[5958] = (layer0_outputs[8293]) & ~(layer0_outputs[1095]);
    assign layer1_outputs[5959] = (layer0_outputs[7575]) & ~(layer0_outputs[7214]);
    assign layer1_outputs[5960] = layer0_outputs[3848];
    assign layer1_outputs[5961] = ~(layer0_outputs[5278]);
    assign layer1_outputs[5962] = ~((layer0_outputs[11540]) ^ (layer0_outputs[12554]));
    assign layer1_outputs[5963] = ~(layer0_outputs[10858]) | (layer0_outputs[5264]);
    assign layer1_outputs[5964] = (layer0_outputs[11098]) ^ (layer0_outputs[1174]);
    assign layer1_outputs[5965] = layer0_outputs[12356];
    assign layer1_outputs[5966] = (layer0_outputs[2244]) ^ (layer0_outputs[9627]);
    assign layer1_outputs[5967] = (layer0_outputs[7836]) & ~(layer0_outputs[12425]);
    assign layer1_outputs[5968] = (layer0_outputs[352]) & ~(layer0_outputs[8225]);
    assign layer1_outputs[5969] = ~(layer0_outputs[2718]) | (layer0_outputs[6145]);
    assign layer1_outputs[5970] = ~((layer0_outputs[2818]) & (layer0_outputs[7990]));
    assign layer1_outputs[5971] = ~(layer0_outputs[6585]);
    assign layer1_outputs[5972] = (layer0_outputs[805]) ^ (layer0_outputs[9825]);
    assign layer1_outputs[5973] = (layer0_outputs[6234]) ^ (layer0_outputs[7686]);
    assign layer1_outputs[5974] = layer0_outputs[6592];
    assign layer1_outputs[5975] = layer0_outputs[10168];
    assign layer1_outputs[5976] = (layer0_outputs[4407]) & (layer0_outputs[8980]);
    assign layer1_outputs[5977] = (layer0_outputs[8398]) & ~(layer0_outputs[9979]);
    assign layer1_outputs[5978] = (layer0_outputs[9470]) & ~(layer0_outputs[9365]);
    assign layer1_outputs[5979] = ~(layer0_outputs[80]) | (layer0_outputs[9269]);
    assign layer1_outputs[5980] = ~(layer0_outputs[8894]) | (layer0_outputs[5596]);
    assign layer1_outputs[5981] = layer0_outputs[8501];
    assign layer1_outputs[5982] = (layer0_outputs[1152]) | (layer0_outputs[635]);
    assign layer1_outputs[5983] = layer0_outputs[8625];
    assign layer1_outputs[5984] = layer0_outputs[5570];
    assign layer1_outputs[5985] = ~(layer0_outputs[10220]) | (layer0_outputs[1542]);
    assign layer1_outputs[5986] = (layer0_outputs[9834]) & (layer0_outputs[12331]);
    assign layer1_outputs[5987] = (layer0_outputs[1604]) & ~(layer0_outputs[11138]);
    assign layer1_outputs[5988] = (layer0_outputs[11311]) & ~(layer0_outputs[4772]);
    assign layer1_outputs[5989] = (layer0_outputs[10994]) ^ (layer0_outputs[6967]);
    assign layer1_outputs[5990] = ~((layer0_outputs[3006]) & (layer0_outputs[4445]));
    assign layer1_outputs[5991] = (layer0_outputs[3327]) ^ (layer0_outputs[5843]);
    assign layer1_outputs[5992] = (layer0_outputs[5104]) & ~(layer0_outputs[435]);
    assign layer1_outputs[5993] = (layer0_outputs[5046]) & ~(layer0_outputs[10489]);
    assign layer1_outputs[5994] = ~(layer0_outputs[1606]) | (layer0_outputs[1522]);
    assign layer1_outputs[5995] = ~(layer0_outputs[4019]);
    assign layer1_outputs[5996] = layer0_outputs[171];
    assign layer1_outputs[5997] = ~(layer0_outputs[5231]) | (layer0_outputs[8153]);
    assign layer1_outputs[5998] = (layer0_outputs[12207]) & ~(layer0_outputs[10802]);
    assign layer1_outputs[5999] = ~(layer0_outputs[144]) | (layer0_outputs[5375]);
    assign layer1_outputs[6000] = layer0_outputs[8528];
    assign layer1_outputs[6001] = ~((layer0_outputs[12358]) & (layer0_outputs[9507]));
    assign layer1_outputs[6002] = layer0_outputs[8720];
    assign layer1_outputs[6003] = (layer0_outputs[366]) ^ (layer0_outputs[12396]);
    assign layer1_outputs[6004] = ~((layer0_outputs[11473]) | (layer0_outputs[6304]));
    assign layer1_outputs[6005] = layer0_outputs[6551];
    assign layer1_outputs[6006] = (layer0_outputs[2839]) & ~(layer0_outputs[5296]);
    assign layer1_outputs[6007] = (layer0_outputs[4070]) & (layer0_outputs[12486]);
    assign layer1_outputs[6008] = layer0_outputs[3342];
    assign layer1_outputs[6009] = ~((layer0_outputs[4402]) & (layer0_outputs[9146]));
    assign layer1_outputs[6010] = (layer0_outputs[1373]) & ~(layer0_outputs[4436]);
    assign layer1_outputs[6011] = layer0_outputs[7304];
    assign layer1_outputs[6012] = ~(layer0_outputs[7302]);
    assign layer1_outputs[6013] = layer0_outputs[4448];
    assign layer1_outputs[6014] = (layer0_outputs[10199]) ^ (layer0_outputs[8559]);
    assign layer1_outputs[6015] = ~((layer0_outputs[7357]) ^ (layer0_outputs[4443]));
    assign layer1_outputs[6016] = (layer0_outputs[9536]) & ~(layer0_outputs[5542]);
    assign layer1_outputs[6017] = (layer0_outputs[2732]) | (layer0_outputs[8152]);
    assign layer1_outputs[6018] = (layer0_outputs[2337]) & ~(layer0_outputs[1909]);
    assign layer1_outputs[6019] = (layer0_outputs[10065]) ^ (layer0_outputs[4062]);
    assign layer1_outputs[6020] = ~((layer0_outputs[74]) ^ (layer0_outputs[12115]));
    assign layer1_outputs[6021] = ~(layer0_outputs[1719]);
    assign layer1_outputs[6022] = ~((layer0_outputs[11080]) | (layer0_outputs[5518]));
    assign layer1_outputs[6023] = (layer0_outputs[11213]) & (layer0_outputs[1195]);
    assign layer1_outputs[6024] = ~((layer0_outputs[4749]) & (layer0_outputs[7028]));
    assign layer1_outputs[6025] = ~(layer0_outputs[7300]);
    assign layer1_outputs[6026] = (layer0_outputs[4617]) & (layer0_outputs[11847]);
    assign layer1_outputs[6027] = ~(layer0_outputs[12675]);
    assign layer1_outputs[6028] = layer0_outputs[3584];
    assign layer1_outputs[6029] = ~((layer0_outputs[11658]) ^ (layer0_outputs[1959]));
    assign layer1_outputs[6030] = ~((layer0_outputs[1748]) & (layer0_outputs[4317]));
    assign layer1_outputs[6031] = ~(layer0_outputs[5861]) | (layer0_outputs[9460]);
    assign layer1_outputs[6032] = (layer0_outputs[10778]) ^ (layer0_outputs[8863]);
    assign layer1_outputs[6033] = (layer0_outputs[2851]) | (layer0_outputs[7410]);
    assign layer1_outputs[6034] = (layer0_outputs[10890]) & ~(layer0_outputs[10061]);
    assign layer1_outputs[6035] = layer0_outputs[9725];
    assign layer1_outputs[6036] = ~(layer0_outputs[4414]) | (layer0_outputs[5002]);
    assign layer1_outputs[6037] = ~(layer0_outputs[11432]);
    assign layer1_outputs[6038] = layer0_outputs[9550];
    assign layer1_outputs[6039] = (layer0_outputs[10816]) & (layer0_outputs[10194]);
    assign layer1_outputs[6040] = ~(layer0_outputs[7334]);
    assign layer1_outputs[6041] = (layer0_outputs[6421]) & ~(layer0_outputs[3843]);
    assign layer1_outputs[6042] = 1'b1;
    assign layer1_outputs[6043] = ~((layer0_outputs[4898]) | (layer0_outputs[1346]));
    assign layer1_outputs[6044] = ~((layer0_outputs[4494]) & (layer0_outputs[9594]));
    assign layer1_outputs[6045] = ~(layer0_outputs[3764]) | (layer0_outputs[8721]);
    assign layer1_outputs[6046] = ~((layer0_outputs[3686]) | (layer0_outputs[9486]));
    assign layer1_outputs[6047] = ~((layer0_outputs[3521]) | (layer0_outputs[12151]));
    assign layer1_outputs[6048] = ~(layer0_outputs[4921]);
    assign layer1_outputs[6049] = layer0_outputs[3164];
    assign layer1_outputs[6050] = (layer0_outputs[6460]) | (layer0_outputs[7207]);
    assign layer1_outputs[6051] = ~(layer0_outputs[96]);
    assign layer1_outputs[6052] = (layer0_outputs[1589]) & ~(layer0_outputs[1070]);
    assign layer1_outputs[6053] = (layer0_outputs[3712]) ^ (layer0_outputs[807]);
    assign layer1_outputs[6054] = ~(layer0_outputs[8159]);
    assign layer1_outputs[6055] = layer0_outputs[9984];
    assign layer1_outputs[6056] = 1'b0;
    assign layer1_outputs[6057] = layer0_outputs[9995];
    assign layer1_outputs[6058] = (layer0_outputs[11296]) & ~(layer0_outputs[12634]);
    assign layer1_outputs[6059] = (layer0_outputs[2071]) ^ (layer0_outputs[562]);
    assign layer1_outputs[6060] = ~(layer0_outputs[11809]) | (layer0_outputs[11791]);
    assign layer1_outputs[6061] = ~(layer0_outputs[3340]);
    assign layer1_outputs[6062] = ~(layer0_outputs[9260]) | (layer0_outputs[6418]);
    assign layer1_outputs[6063] = ~(layer0_outputs[871]);
    assign layer1_outputs[6064] = ~(layer0_outputs[3941]);
    assign layer1_outputs[6065] = layer0_outputs[8924];
    assign layer1_outputs[6066] = (layer0_outputs[10531]) & ~(layer0_outputs[2997]);
    assign layer1_outputs[6067] = 1'b0;
    assign layer1_outputs[6068] = (layer0_outputs[10408]) & ~(layer0_outputs[5751]);
    assign layer1_outputs[6069] = (layer0_outputs[7143]) | (layer0_outputs[5]);
    assign layer1_outputs[6070] = layer0_outputs[12353];
    assign layer1_outputs[6071] = layer0_outputs[7675];
    assign layer1_outputs[6072] = layer0_outputs[7821];
    assign layer1_outputs[6073] = (layer0_outputs[10842]) | (layer0_outputs[11484]);
    assign layer1_outputs[6074] = ~(layer0_outputs[5146]);
    assign layer1_outputs[6075] = ~(layer0_outputs[8871]) | (layer0_outputs[10636]);
    assign layer1_outputs[6076] = layer0_outputs[12629];
    assign layer1_outputs[6077] = (layer0_outputs[7813]) ^ (layer0_outputs[3598]);
    assign layer1_outputs[6078] = layer0_outputs[2081];
    assign layer1_outputs[6079] = (layer0_outputs[7424]) & ~(layer0_outputs[4436]);
    assign layer1_outputs[6080] = ~(layer0_outputs[7612]);
    assign layer1_outputs[6081] = (layer0_outputs[12223]) | (layer0_outputs[12361]);
    assign layer1_outputs[6082] = (layer0_outputs[10215]) ^ (layer0_outputs[3430]);
    assign layer1_outputs[6083] = (layer0_outputs[5630]) | (layer0_outputs[3740]);
    assign layer1_outputs[6084] = (layer0_outputs[1039]) ^ (layer0_outputs[6441]);
    assign layer1_outputs[6085] = ~(layer0_outputs[8556]) | (layer0_outputs[12723]);
    assign layer1_outputs[6086] = (layer0_outputs[7128]) | (layer0_outputs[3657]);
    assign layer1_outputs[6087] = (layer0_outputs[10878]) & ~(layer0_outputs[5046]);
    assign layer1_outputs[6088] = ~(layer0_outputs[8620]);
    assign layer1_outputs[6089] = (layer0_outputs[12049]) ^ (layer0_outputs[5364]);
    assign layer1_outputs[6090] = ~((layer0_outputs[3866]) & (layer0_outputs[2276]));
    assign layer1_outputs[6091] = layer0_outputs[9337];
    assign layer1_outputs[6092] = (layer0_outputs[516]) | (layer0_outputs[5392]);
    assign layer1_outputs[6093] = ~(layer0_outputs[5492]);
    assign layer1_outputs[6094] = layer0_outputs[4797];
    assign layer1_outputs[6095] = ~(layer0_outputs[10575]) | (layer0_outputs[8193]);
    assign layer1_outputs[6096] = 1'b1;
    assign layer1_outputs[6097] = ~(layer0_outputs[2136]) | (layer0_outputs[4317]);
    assign layer1_outputs[6098] = layer0_outputs[12133];
    assign layer1_outputs[6099] = ~(layer0_outputs[6727]);
    assign layer1_outputs[6100] = (layer0_outputs[6091]) & (layer0_outputs[6386]);
    assign layer1_outputs[6101] = ~(layer0_outputs[2124]);
    assign layer1_outputs[6102] = (layer0_outputs[11746]) ^ (layer0_outputs[6182]);
    assign layer1_outputs[6103] = layer0_outputs[2639];
    assign layer1_outputs[6104] = (layer0_outputs[6671]) & (layer0_outputs[2769]);
    assign layer1_outputs[6105] = (layer0_outputs[2814]) | (layer0_outputs[4488]);
    assign layer1_outputs[6106] = (layer0_outputs[10861]) | (layer0_outputs[4877]);
    assign layer1_outputs[6107] = 1'b1;
    assign layer1_outputs[6108] = ~(layer0_outputs[6236]);
    assign layer1_outputs[6109] = ~(layer0_outputs[9477]);
    assign layer1_outputs[6110] = ~(layer0_outputs[6452]);
    assign layer1_outputs[6111] = (layer0_outputs[11734]) & (layer0_outputs[2682]);
    assign layer1_outputs[6112] = ~((layer0_outputs[3556]) ^ (layer0_outputs[3451]));
    assign layer1_outputs[6113] = ~(layer0_outputs[9770]);
    assign layer1_outputs[6114] = (layer0_outputs[3910]) | (layer0_outputs[4897]);
    assign layer1_outputs[6115] = (layer0_outputs[9505]) & ~(layer0_outputs[2479]);
    assign layer1_outputs[6116] = ~(layer0_outputs[9990]);
    assign layer1_outputs[6117] = layer0_outputs[12105];
    assign layer1_outputs[6118] = layer0_outputs[8357];
    assign layer1_outputs[6119] = layer0_outputs[12049];
    assign layer1_outputs[6120] = (layer0_outputs[736]) & (layer0_outputs[1223]);
    assign layer1_outputs[6121] = layer0_outputs[7163];
    assign layer1_outputs[6122] = ~((layer0_outputs[4379]) | (layer0_outputs[11192]));
    assign layer1_outputs[6123] = ~(layer0_outputs[2329]) | (layer0_outputs[12523]);
    assign layer1_outputs[6124] = (layer0_outputs[12515]) & ~(layer0_outputs[2187]);
    assign layer1_outputs[6125] = (layer0_outputs[11852]) & (layer0_outputs[32]);
    assign layer1_outputs[6126] = (layer0_outputs[1943]) | (layer0_outputs[3572]);
    assign layer1_outputs[6127] = layer0_outputs[11778];
    assign layer1_outputs[6128] = (layer0_outputs[9319]) | (layer0_outputs[4905]);
    assign layer1_outputs[6129] = (layer0_outputs[11557]) & ~(layer0_outputs[9584]);
    assign layer1_outputs[6130] = ~((layer0_outputs[7031]) & (layer0_outputs[12198]));
    assign layer1_outputs[6131] = ~((layer0_outputs[11020]) & (layer0_outputs[12557]));
    assign layer1_outputs[6132] = (layer0_outputs[142]) | (layer0_outputs[2646]);
    assign layer1_outputs[6133] = 1'b1;
    assign layer1_outputs[6134] = ~(layer0_outputs[2846]);
    assign layer1_outputs[6135] = ~(layer0_outputs[4899]);
    assign layer1_outputs[6136] = layer0_outputs[554];
    assign layer1_outputs[6137] = layer0_outputs[4857];
    assign layer1_outputs[6138] = ~(layer0_outputs[10273]) | (layer0_outputs[5905]);
    assign layer1_outputs[6139] = (layer0_outputs[10190]) | (layer0_outputs[1511]);
    assign layer1_outputs[6140] = (layer0_outputs[5594]) | (layer0_outputs[8160]);
    assign layer1_outputs[6141] = layer0_outputs[5159];
    assign layer1_outputs[6142] = ~((layer0_outputs[4010]) | (layer0_outputs[6536]));
    assign layer1_outputs[6143] = (layer0_outputs[12620]) & (layer0_outputs[6472]);
    assign layer1_outputs[6144] = ~((layer0_outputs[7855]) & (layer0_outputs[6834]));
    assign layer1_outputs[6145] = layer0_outputs[7857];
    assign layer1_outputs[6146] = ~((layer0_outputs[12342]) ^ (layer0_outputs[1978]));
    assign layer1_outputs[6147] = layer0_outputs[10340];
    assign layer1_outputs[6148] = ~(layer0_outputs[6130]);
    assign layer1_outputs[6149] = ~(layer0_outputs[2586]);
    assign layer1_outputs[6150] = (layer0_outputs[1090]) & ~(layer0_outputs[9152]);
    assign layer1_outputs[6151] = 1'b0;
    assign layer1_outputs[6152] = (layer0_outputs[10373]) & ~(layer0_outputs[10453]);
    assign layer1_outputs[6153] = (layer0_outputs[10870]) & (layer0_outputs[4058]);
    assign layer1_outputs[6154] = (layer0_outputs[7893]) & ~(layer0_outputs[9613]);
    assign layer1_outputs[6155] = ~((layer0_outputs[11248]) ^ (layer0_outputs[6297]));
    assign layer1_outputs[6156] = ~(layer0_outputs[5512]);
    assign layer1_outputs[6157] = 1'b0;
    assign layer1_outputs[6158] = ~((layer0_outputs[9459]) | (layer0_outputs[10787]));
    assign layer1_outputs[6159] = ~(layer0_outputs[3391]) | (layer0_outputs[2343]);
    assign layer1_outputs[6160] = layer0_outputs[986];
    assign layer1_outputs[6161] = 1'b0;
    assign layer1_outputs[6162] = ~(layer0_outputs[6412]) | (layer0_outputs[12699]);
    assign layer1_outputs[6163] = ~((layer0_outputs[4309]) ^ (layer0_outputs[9512]));
    assign layer1_outputs[6164] = (layer0_outputs[9978]) ^ (layer0_outputs[6276]);
    assign layer1_outputs[6165] = ~((layer0_outputs[1002]) & (layer0_outputs[8506]));
    assign layer1_outputs[6166] = ~(layer0_outputs[4660]) | (layer0_outputs[5824]);
    assign layer1_outputs[6167] = (layer0_outputs[11471]) | (layer0_outputs[6815]);
    assign layer1_outputs[6168] = (layer0_outputs[2226]) & ~(layer0_outputs[2518]);
    assign layer1_outputs[6169] = layer0_outputs[1878];
    assign layer1_outputs[6170] = ~(layer0_outputs[2246]) | (layer0_outputs[6622]);
    assign layer1_outputs[6171] = ~(layer0_outputs[5026]);
    assign layer1_outputs[6172] = ~((layer0_outputs[9130]) ^ (layer0_outputs[11486]));
    assign layer1_outputs[6173] = layer0_outputs[7248];
    assign layer1_outputs[6174] = ~((layer0_outputs[128]) | (layer0_outputs[1207]));
    assign layer1_outputs[6175] = ~(layer0_outputs[12423]);
    assign layer1_outputs[6176] = (layer0_outputs[2791]) & ~(layer0_outputs[11729]);
    assign layer1_outputs[6177] = ~(layer0_outputs[6459]) | (layer0_outputs[8462]);
    assign layer1_outputs[6178] = layer0_outputs[8926];
    assign layer1_outputs[6179] = layer0_outputs[2855];
    assign layer1_outputs[6180] = (layer0_outputs[4047]) & ~(layer0_outputs[5218]);
    assign layer1_outputs[6181] = ~(layer0_outputs[3151]);
    assign layer1_outputs[6182] = (layer0_outputs[1697]) | (layer0_outputs[1617]);
    assign layer1_outputs[6183] = ~((layer0_outputs[7108]) & (layer0_outputs[4514]));
    assign layer1_outputs[6184] = layer0_outputs[8110];
    assign layer1_outputs[6185] = ~((layer0_outputs[2712]) ^ (layer0_outputs[1957]));
    assign layer1_outputs[6186] = layer0_outputs[11637];
    assign layer1_outputs[6187] = (layer0_outputs[1902]) & ~(layer0_outputs[2437]);
    assign layer1_outputs[6188] = ~((layer0_outputs[8372]) ^ (layer0_outputs[4728]));
    assign layer1_outputs[6189] = ~(layer0_outputs[8781]);
    assign layer1_outputs[6190] = (layer0_outputs[4017]) & ~(layer0_outputs[12373]);
    assign layer1_outputs[6191] = layer0_outputs[6572];
    assign layer1_outputs[6192] = layer0_outputs[12704];
    assign layer1_outputs[6193] = layer0_outputs[10805];
    assign layer1_outputs[6194] = ~((layer0_outputs[11528]) | (layer0_outputs[1749]));
    assign layer1_outputs[6195] = layer0_outputs[1319];
    assign layer1_outputs[6196] = (layer0_outputs[7810]) | (layer0_outputs[394]);
    assign layer1_outputs[6197] = ~(layer0_outputs[12246]);
    assign layer1_outputs[6198] = ~(layer0_outputs[7330]);
    assign layer1_outputs[6199] = (layer0_outputs[9853]) ^ (layer0_outputs[2036]);
    assign layer1_outputs[6200] = (layer0_outputs[1738]) & ~(layer0_outputs[497]);
    assign layer1_outputs[6201] = layer0_outputs[2091];
    assign layer1_outputs[6202] = layer0_outputs[9494];
    assign layer1_outputs[6203] = ~((layer0_outputs[12676]) | (layer0_outputs[656]));
    assign layer1_outputs[6204] = ~(layer0_outputs[4492]);
    assign layer1_outputs[6205] = ~((layer0_outputs[6210]) & (layer0_outputs[7826]));
    assign layer1_outputs[6206] = layer0_outputs[2418];
    assign layer1_outputs[6207] = ~((layer0_outputs[9238]) & (layer0_outputs[2664]));
    assign layer1_outputs[6208] = ~(layer0_outputs[7953]);
    assign layer1_outputs[6209] = ~(layer0_outputs[4269]);
    assign layer1_outputs[6210] = layer0_outputs[12297];
    assign layer1_outputs[6211] = (layer0_outputs[6221]) & ~(layer0_outputs[4245]);
    assign layer1_outputs[6212] = ~(layer0_outputs[4399]);
    assign layer1_outputs[6213] = (layer0_outputs[7492]) & ~(layer0_outputs[1822]);
    assign layer1_outputs[6214] = ~(layer0_outputs[7579]);
    assign layer1_outputs[6215] = (layer0_outputs[569]) ^ (layer0_outputs[2006]);
    assign layer1_outputs[6216] = ~((layer0_outputs[11253]) | (layer0_outputs[4845]));
    assign layer1_outputs[6217] = ~((layer0_outputs[4438]) ^ (layer0_outputs[6023]));
    assign layer1_outputs[6218] = ~((layer0_outputs[12792]) | (layer0_outputs[9015]));
    assign layer1_outputs[6219] = layer0_outputs[4495];
    assign layer1_outputs[6220] = (layer0_outputs[5101]) ^ (layer0_outputs[9326]);
    assign layer1_outputs[6221] = (layer0_outputs[12543]) & ~(layer0_outputs[7538]);
    assign layer1_outputs[6222] = (layer0_outputs[466]) ^ (layer0_outputs[110]);
    assign layer1_outputs[6223] = layer0_outputs[8038];
    assign layer1_outputs[6224] = ~((layer0_outputs[8104]) ^ (layer0_outputs[9091]));
    assign layer1_outputs[6225] = ~(layer0_outputs[11182]);
    assign layer1_outputs[6226] = (layer0_outputs[5589]) & ~(layer0_outputs[6143]);
    assign layer1_outputs[6227] = (layer0_outputs[2417]) & (layer0_outputs[6679]);
    assign layer1_outputs[6228] = (layer0_outputs[3370]) & ~(layer0_outputs[9692]);
    assign layer1_outputs[6229] = 1'b0;
    assign layer1_outputs[6230] = ~(layer0_outputs[11351]) | (layer0_outputs[10200]);
    assign layer1_outputs[6231] = ~(layer0_outputs[97]);
    assign layer1_outputs[6232] = layer0_outputs[9912];
    assign layer1_outputs[6233] = layer0_outputs[7683];
    assign layer1_outputs[6234] = 1'b0;
    assign layer1_outputs[6235] = (layer0_outputs[10952]) & ~(layer0_outputs[5102]);
    assign layer1_outputs[6236] = layer0_outputs[10751];
    assign layer1_outputs[6237] = layer0_outputs[1200];
    assign layer1_outputs[6238] = layer0_outputs[12604];
    assign layer1_outputs[6239] = (layer0_outputs[10979]) & (layer0_outputs[8921]);
    assign layer1_outputs[6240] = ~((layer0_outputs[6843]) ^ (layer0_outputs[8297]));
    assign layer1_outputs[6241] = (layer0_outputs[6433]) & ~(layer0_outputs[5392]);
    assign layer1_outputs[6242] = ~((layer0_outputs[12263]) | (layer0_outputs[1815]));
    assign layer1_outputs[6243] = (layer0_outputs[3795]) & ~(layer0_outputs[8128]);
    assign layer1_outputs[6244] = (layer0_outputs[2394]) ^ (layer0_outputs[9133]);
    assign layer1_outputs[6245] = ~(layer0_outputs[193]);
    assign layer1_outputs[6246] = (layer0_outputs[1813]) ^ (layer0_outputs[10982]);
    assign layer1_outputs[6247] = layer0_outputs[1243];
    assign layer1_outputs[6248] = ~(layer0_outputs[3675]);
    assign layer1_outputs[6249] = ~((layer0_outputs[2556]) & (layer0_outputs[5198]));
    assign layer1_outputs[6250] = ~((layer0_outputs[287]) | (layer0_outputs[11299]));
    assign layer1_outputs[6251] = (layer0_outputs[2912]) & (layer0_outputs[1012]);
    assign layer1_outputs[6252] = 1'b1;
    assign layer1_outputs[6253] = ~(layer0_outputs[2731]);
    assign layer1_outputs[6254] = layer0_outputs[4287];
    assign layer1_outputs[6255] = ~((layer0_outputs[7268]) ^ (layer0_outputs[12591]));
    assign layer1_outputs[6256] = ~(layer0_outputs[10505]);
    assign layer1_outputs[6257] = (layer0_outputs[11630]) & ~(layer0_outputs[9769]);
    assign layer1_outputs[6258] = layer0_outputs[10107];
    assign layer1_outputs[6259] = ~(layer0_outputs[12112]);
    assign layer1_outputs[6260] = layer0_outputs[10768];
    assign layer1_outputs[6261] = (layer0_outputs[2237]) & (layer0_outputs[6103]);
    assign layer1_outputs[6262] = ~((layer0_outputs[5951]) & (layer0_outputs[973]));
    assign layer1_outputs[6263] = layer0_outputs[9936];
    assign layer1_outputs[6264] = ~((layer0_outputs[4571]) & (layer0_outputs[380]));
    assign layer1_outputs[6265] = layer0_outputs[12734];
    assign layer1_outputs[6266] = layer0_outputs[6953];
    assign layer1_outputs[6267] = ~((layer0_outputs[9513]) & (layer0_outputs[5601]));
    assign layer1_outputs[6268] = layer0_outputs[8576];
    assign layer1_outputs[6269] = 1'b1;
    assign layer1_outputs[6270] = (layer0_outputs[8704]) & ~(layer0_outputs[4007]);
    assign layer1_outputs[6271] = layer0_outputs[9693];
    assign layer1_outputs[6272] = ~(layer0_outputs[5664]);
    assign layer1_outputs[6273] = ~((layer0_outputs[8228]) & (layer0_outputs[7543]));
    assign layer1_outputs[6274] = (layer0_outputs[4288]) ^ (layer0_outputs[9523]);
    assign layer1_outputs[6275] = layer0_outputs[12296];
    assign layer1_outputs[6276] = layer0_outputs[1449];
    assign layer1_outputs[6277] = 1'b1;
    assign layer1_outputs[6278] = layer0_outputs[7819];
    assign layer1_outputs[6279] = ~(layer0_outputs[7544]) | (layer0_outputs[7691]);
    assign layer1_outputs[6280] = (layer0_outputs[10795]) & ~(layer0_outputs[7596]);
    assign layer1_outputs[6281] = (layer0_outputs[9711]) & ~(layer0_outputs[10871]);
    assign layer1_outputs[6282] = (layer0_outputs[120]) & ~(layer0_outputs[7606]);
    assign layer1_outputs[6283] = ~(layer0_outputs[2991]);
    assign layer1_outputs[6284] = (layer0_outputs[3243]) ^ (layer0_outputs[4164]);
    assign layer1_outputs[6285] = (layer0_outputs[7716]) | (layer0_outputs[6199]);
    assign layer1_outputs[6286] = layer0_outputs[12028];
    assign layer1_outputs[6287] = ~(layer0_outputs[4960]);
    assign layer1_outputs[6288] = layer0_outputs[9962];
    assign layer1_outputs[6289] = ~(layer0_outputs[10595]) | (layer0_outputs[9809]);
    assign layer1_outputs[6290] = (layer0_outputs[4987]) & (layer0_outputs[6862]);
    assign layer1_outputs[6291] = (layer0_outputs[9435]) ^ (layer0_outputs[4051]);
    assign layer1_outputs[6292] = ~(layer0_outputs[12774]);
    assign layer1_outputs[6293] = ~(layer0_outputs[11162]);
    assign layer1_outputs[6294] = layer0_outputs[7427];
    assign layer1_outputs[6295] = ~((layer0_outputs[7918]) | (layer0_outputs[7616]));
    assign layer1_outputs[6296] = (layer0_outputs[10684]) & ~(layer0_outputs[6618]);
    assign layer1_outputs[6297] = ~((layer0_outputs[8497]) | (layer0_outputs[6801]));
    assign layer1_outputs[6298] = (layer0_outputs[11420]) & ~(layer0_outputs[9259]);
    assign layer1_outputs[6299] = ~(layer0_outputs[753]);
    assign layer1_outputs[6300] = layer0_outputs[3467];
    assign layer1_outputs[6301] = layer0_outputs[7803];
    assign layer1_outputs[6302] = ~(layer0_outputs[12202]) | (layer0_outputs[10129]);
    assign layer1_outputs[6303] = ~(layer0_outputs[8243]) | (layer0_outputs[6241]);
    assign layer1_outputs[6304] = (layer0_outputs[5944]) & (layer0_outputs[8570]);
    assign layer1_outputs[6305] = ~(layer0_outputs[7714]);
    assign layer1_outputs[6306] = (layer0_outputs[9913]) | (layer0_outputs[4711]);
    assign layer1_outputs[6307] = (layer0_outputs[5753]) | (layer0_outputs[9443]);
    assign layer1_outputs[6308] = ~(layer0_outputs[6896]);
    assign layer1_outputs[6309] = (layer0_outputs[11908]) & (layer0_outputs[8847]);
    assign layer1_outputs[6310] = layer0_outputs[3942];
    assign layer1_outputs[6311] = (layer0_outputs[651]) | (layer0_outputs[9710]);
    assign layer1_outputs[6312] = (layer0_outputs[6062]) | (layer0_outputs[5969]);
    assign layer1_outputs[6313] = ~((layer0_outputs[12471]) & (layer0_outputs[4611]));
    assign layer1_outputs[6314] = layer0_outputs[7510];
    assign layer1_outputs[6315] = ~(layer0_outputs[9122]);
    assign layer1_outputs[6316] = layer0_outputs[2853];
    assign layer1_outputs[6317] = ~(layer0_outputs[4919]) | (layer0_outputs[3582]);
    assign layer1_outputs[6318] = (layer0_outputs[2315]) | (layer0_outputs[10689]);
    assign layer1_outputs[6319] = ~(layer0_outputs[7522]);
    assign layer1_outputs[6320] = ~(layer0_outputs[1642]) | (layer0_outputs[99]);
    assign layer1_outputs[6321] = ~(layer0_outputs[1149]) | (layer0_outputs[11547]);
    assign layer1_outputs[6322] = ~(layer0_outputs[7948]);
    assign layer1_outputs[6323] = ~((layer0_outputs[2292]) & (layer0_outputs[1491]));
    assign layer1_outputs[6324] = ~(layer0_outputs[9213]) | (layer0_outputs[8832]);
    assign layer1_outputs[6325] = ~(layer0_outputs[10232]);
    assign layer1_outputs[6326] = ~(layer0_outputs[20]);
    assign layer1_outputs[6327] = ~((layer0_outputs[7825]) & (layer0_outputs[6657]));
    assign layer1_outputs[6328] = layer0_outputs[6320];
    assign layer1_outputs[6329] = ~(layer0_outputs[136]) | (layer0_outputs[5777]);
    assign layer1_outputs[6330] = ~(layer0_outputs[8149]) | (layer0_outputs[8713]);
    assign layer1_outputs[6331] = ~(layer0_outputs[3772]);
    assign layer1_outputs[6332] = (layer0_outputs[8680]) | (layer0_outputs[3707]);
    assign layer1_outputs[6333] = ~((layer0_outputs[9782]) | (layer0_outputs[4422]));
    assign layer1_outputs[6334] = ~((layer0_outputs[12539]) & (layer0_outputs[3536]));
    assign layer1_outputs[6335] = (layer0_outputs[11326]) | (layer0_outputs[11446]);
    assign layer1_outputs[6336] = (layer0_outputs[1381]) & ~(layer0_outputs[10534]);
    assign layer1_outputs[6337] = (layer0_outputs[10665]) & (layer0_outputs[11452]);
    assign layer1_outputs[6338] = layer0_outputs[12186];
    assign layer1_outputs[6339] = (layer0_outputs[6602]) & ~(layer0_outputs[12299]);
    assign layer1_outputs[6340] = (layer0_outputs[12199]) ^ (layer0_outputs[418]);
    assign layer1_outputs[6341] = layer0_outputs[7694];
    assign layer1_outputs[6342] = ~(layer0_outputs[10556]) | (layer0_outputs[6149]);
    assign layer1_outputs[6343] = ~((layer0_outputs[5194]) ^ (layer0_outputs[4451]));
    assign layer1_outputs[6344] = (layer0_outputs[10554]) | (layer0_outputs[1675]);
    assign layer1_outputs[6345] = ~(layer0_outputs[6046]) | (layer0_outputs[2387]);
    assign layer1_outputs[6346] = (layer0_outputs[4972]) & ~(layer0_outputs[38]);
    assign layer1_outputs[6347] = ~(layer0_outputs[2003]) | (layer0_outputs[1991]);
    assign layer1_outputs[6348] = (layer0_outputs[5920]) & ~(layer0_outputs[1172]);
    assign layer1_outputs[6349] = ~(layer0_outputs[449]) | (layer0_outputs[825]);
    assign layer1_outputs[6350] = ~((layer0_outputs[228]) | (layer0_outputs[12543]));
    assign layer1_outputs[6351] = ~(layer0_outputs[858]) | (layer0_outputs[12407]);
    assign layer1_outputs[6352] = ~(layer0_outputs[11771]) | (layer0_outputs[8065]);
    assign layer1_outputs[6353] = ~((layer0_outputs[10600]) ^ (layer0_outputs[5425]));
    assign layer1_outputs[6354] = layer0_outputs[1720];
    assign layer1_outputs[6355] = ~(layer0_outputs[11462]) | (layer0_outputs[5812]);
    assign layer1_outputs[6356] = ~(layer0_outputs[2654]) | (layer0_outputs[8082]);
    assign layer1_outputs[6357] = ~(layer0_outputs[3010]);
    assign layer1_outputs[6358] = ~(layer0_outputs[3700]);
    assign layer1_outputs[6359] = layer0_outputs[11698];
    assign layer1_outputs[6360] = layer0_outputs[570];
    assign layer1_outputs[6361] = ~(layer0_outputs[6129]);
    assign layer1_outputs[6362] = ~(layer0_outputs[4450]);
    assign layer1_outputs[6363] = (layer0_outputs[5248]) & ~(layer0_outputs[9786]);
    assign layer1_outputs[6364] = ~((layer0_outputs[4321]) & (layer0_outputs[3242]));
    assign layer1_outputs[6365] = ~((layer0_outputs[4974]) | (layer0_outputs[7897]));
    assign layer1_outputs[6366] = (layer0_outputs[12121]) & (layer0_outputs[1824]);
    assign layer1_outputs[6367] = ~(layer0_outputs[5235]);
    assign layer1_outputs[6368] = layer0_outputs[3331];
    assign layer1_outputs[6369] = ~(layer0_outputs[7863]) | (layer0_outputs[5768]);
    assign layer1_outputs[6370] = ~((layer0_outputs[11622]) & (layer0_outputs[6506]));
    assign layer1_outputs[6371] = ~(layer0_outputs[4637]);
    assign layer1_outputs[6372] = (layer0_outputs[11612]) & ~(layer0_outputs[7563]);
    assign layer1_outputs[6373] = ~(layer0_outputs[9932]);
    assign layer1_outputs[6374] = (layer0_outputs[1203]) ^ (layer0_outputs[1105]);
    assign layer1_outputs[6375] = (layer0_outputs[8331]) | (layer0_outputs[11825]);
    assign layer1_outputs[6376] = layer0_outputs[5003];
    assign layer1_outputs[6377] = (layer0_outputs[8620]) & (layer0_outputs[11395]);
    assign layer1_outputs[6378] = 1'b1;
    assign layer1_outputs[6379] = (layer0_outputs[10867]) & (layer0_outputs[8892]);
    assign layer1_outputs[6380] = ~(layer0_outputs[1317]) | (layer0_outputs[8665]);
    assign layer1_outputs[6381] = layer0_outputs[7690];
    assign layer1_outputs[6382] = ~((layer0_outputs[273]) & (layer0_outputs[5832]));
    assign layer1_outputs[6383] = layer0_outputs[3611];
    assign layer1_outputs[6384] = ~(layer0_outputs[11304]);
    assign layer1_outputs[6385] = ~((layer0_outputs[7931]) & (layer0_outputs[10559]));
    assign layer1_outputs[6386] = ~(layer0_outputs[2064]) | (layer0_outputs[8539]);
    assign layer1_outputs[6387] = layer0_outputs[11907];
    assign layer1_outputs[6388] = (layer0_outputs[1289]) & ~(layer0_outputs[10668]);
    assign layer1_outputs[6389] = ~((layer0_outputs[5096]) ^ (layer0_outputs[8729]));
    assign layer1_outputs[6390] = ~(layer0_outputs[8918]) | (layer0_outputs[4920]);
    assign layer1_outputs[6391] = ~(layer0_outputs[10050]);
    assign layer1_outputs[6392] = (layer0_outputs[6437]) & ~(layer0_outputs[1960]);
    assign layer1_outputs[6393] = ~(layer0_outputs[10943]) | (layer0_outputs[1670]);
    assign layer1_outputs[6394] = ~(layer0_outputs[5451]) | (layer0_outputs[11628]);
    assign layer1_outputs[6395] = layer0_outputs[5808];
    assign layer1_outputs[6396] = (layer0_outputs[8130]) & ~(layer0_outputs[9324]);
    assign layer1_outputs[6397] = ~(layer0_outputs[9032]);
    assign layer1_outputs[6398] = (layer0_outputs[10425]) | (layer0_outputs[3249]);
    assign layer1_outputs[6399] = ~(layer0_outputs[7842]);
    assign layer1_outputs[6400] = (layer0_outputs[1709]) ^ (layer0_outputs[9307]);
    assign layer1_outputs[6401] = layer0_outputs[1438];
    assign layer1_outputs[6402] = (layer0_outputs[9563]) & ~(layer0_outputs[4534]);
    assign layer1_outputs[6403] = layer0_outputs[6209];
    assign layer1_outputs[6404] = ~(layer0_outputs[2011]);
    assign layer1_outputs[6405] = ~((layer0_outputs[9805]) & (layer0_outputs[4062]));
    assign layer1_outputs[6406] = (layer0_outputs[7276]) ^ (layer0_outputs[8241]);
    assign layer1_outputs[6407] = layer0_outputs[6010];
    assign layer1_outputs[6408] = layer0_outputs[10750];
    assign layer1_outputs[6409] = (layer0_outputs[2510]) | (layer0_outputs[4362]);
    assign layer1_outputs[6410] = ~(layer0_outputs[296]) | (layer0_outputs[10270]);
    assign layer1_outputs[6411] = layer0_outputs[9241];
    assign layer1_outputs[6412] = ~(layer0_outputs[12463]) | (layer0_outputs[1026]);
    assign layer1_outputs[6413] = (layer0_outputs[9248]) | (layer0_outputs[26]);
    assign layer1_outputs[6414] = layer0_outputs[134];
    assign layer1_outputs[6415] = ~((layer0_outputs[6139]) & (layer0_outputs[5326]));
    assign layer1_outputs[6416] = layer0_outputs[3060];
    assign layer1_outputs[6417] = ~((layer0_outputs[8351]) | (layer0_outputs[5115]));
    assign layer1_outputs[6418] = ~(layer0_outputs[9657]);
    assign layer1_outputs[6419] = (layer0_outputs[4041]) & ~(layer0_outputs[11985]);
    assign layer1_outputs[6420] = ~(layer0_outputs[7750]);
    assign layer1_outputs[6421] = (layer0_outputs[8297]) ^ (layer0_outputs[2115]);
    assign layer1_outputs[6422] = 1'b0;
    assign layer1_outputs[6423] = ~((layer0_outputs[5431]) | (layer0_outputs[2149]));
    assign layer1_outputs[6424] = ~(layer0_outputs[797]);
    assign layer1_outputs[6425] = (layer0_outputs[8831]) & ~(layer0_outputs[5615]);
    assign layer1_outputs[6426] = ~(layer0_outputs[12437]) | (layer0_outputs[2541]);
    assign layer1_outputs[6427] = ~(layer0_outputs[3536]);
    assign layer1_outputs[6428] = layer0_outputs[486];
    assign layer1_outputs[6429] = layer0_outputs[11836];
    assign layer1_outputs[6430] = (layer0_outputs[10353]) & ~(layer0_outputs[8799]);
    assign layer1_outputs[6431] = layer0_outputs[895];
    assign layer1_outputs[6432] = ~(layer0_outputs[4659]) | (layer0_outputs[2278]);
    assign layer1_outputs[6433] = ~((layer0_outputs[11008]) ^ (layer0_outputs[11532]));
    assign layer1_outputs[6434] = layer0_outputs[2609];
    assign layer1_outputs[6435] = ~(layer0_outputs[3743]);
    assign layer1_outputs[6436] = layer0_outputs[10158];
    assign layer1_outputs[6437] = (layer0_outputs[9850]) | (layer0_outputs[368]);
    assign layer1_outputs[6438] = ~(layer0_outputs[1949]);
    assign layer1_outputs[6439] = ~((layer0_outputs[3912]) & (layer0_outputs[9198]));
    assign layer1_outputs[6440] = ~(layer0_outputs[7433]) | (layer0_outputs[5061]);
    assign layer1_outputs[6441] = ~((layer0_outputs[4486]) | (layer0_outputs[1285]));
    assign layer1_outputs[6442] = ~(layer0_outputs[2408]) | (layer0_outputs[9658]);
    assign layer1_outputs[6443] = ~(layer0_outputs[6738]) | (layer0_outputs[10720]);
    assign layer1_outputs[6444] = layer0_outputs[7465];
    assign layer1_outputs[6445] = (layer0_outputs[8091]) & (layer0_outputs[9701]);
    assign layer1_outputs[6446] = layer0_outputs[1787];
    assign layer1_outputs[6447] = ~(layer0_outputs[12620]);
    assign layer1_outputs[6448] = ~(layer0_outputs[10203]);
    assign layer1_outputs[6449] = (layer0_outputs[4588]) & ~(layer0_outputs[12752]);
    assign layer1_outputs[6450] = (layer0_outputs[10514]) & ~(layer0_outputs[6445]);
    assign layer1_outputs[6451] = (layer0_outputs[295]) | (layer0_outputs[6824]);
    assign layer1_outputs[6452] = (layer0_outputs[9413]) & (layer0_outputs[9284]);
    assign layer1_outputs[6453] = ~((layer0_outputs[8771]) & (layer0_outputs[7076]));
    assign layer1_outputs[6454] = (layer0_outputs[8348]) & ~(layer0_outputs[9815]);
    assign layer1_outputs[6455] = layer0_outputs[5209];
    assign layer1_outputs[6456] = ~((layer0_outputs[11081]) ^ (layer0_outputs[2993]));
    assign layer1_outputs[6457] = (layer0_outputs[12768]) & ~(layer0_outputs[136]);
    assign layer1_outputs[6458] = (layer0_outputs[8774]) & ~(layer0_outputs[987]);
    assign layer1_outputs[6459] = layer0_outputs[1020];
    assign layer1_outputs[6460] = ~(layer0_outputs[12023]) | (layer0_outputs[561]);
    assign layer1_outputs[6461] = ~(layer0_outputs[1031]);
    assign layer1_outputs[6462] = (layer0_outputs[1114]) & ~(layer0_outputs[2533]);
    assign layer1_outputs[6463] = layer0_outputs[5559];
    assign layer1_outputs[6464] = layer0_outputs[7822];
    assign layer1_outputs[6465] = layer0_outputs[1699];
    assign layer1_outputs[6466] = ~(layer0_outputs[9713]);
    assign layer1_outputs[6467] = (layer0_outputs[6973]) | (layer0_outputs[9340]);
    assign layer1_outputs[6468] = (layer0_outputs[9014]) ^ (layer0_outputs[10137]);
    assign layer1_outputs[6469] = ~(layer0_outputs[12026]);
    assign layer1_outputs[6470] = ~(layer0_outputs[5861]) | (layer0_outputs[6363]);
    assign layer1_outputs[6471] = ~((layer0_outputs[7406]) & (layer0_outputs[3706]));
    assign layer1_outputs[6472] = ~(layer0_outputs[1205]);
    assign layer1_outputs[6473] = ~(layer0_outputs[8065]);
    assign layer1_outputs[6474] = ~((layer0_outputs[7170]) | (layer0_outputs[5224]));
    assign layer1_outputs[6475] = ~((layer0_outputs[7133]) & (layer0_outputs[3666]));
    assign layer1_outputs[6476] = (layer0_outputs[3485]) & ~(layer0_outputs[11061]);
    assign layer1_outputs[6477] = (layer0_outputs[7114]) | (layer0_outputs[8087]);
    assign layer1_outputs[6478] = (layer0_outputs[3392]) | (layer0_outputs[8887]);
    assign layer1_outputs[6479] = (layer0_outputs[3872]) ^ (layer0_outputs[11662]);
    assign layer1_outputs[6480] = ~(layer0_outputs[1016]) | (layer0_outputs[11137]);
    assign layer1_outputs[6481] = 1'b1;
    assign layer1_outputs[6482] = ~(layer0_outputs[6012]) | (layer0_outputs[4691]);
    assign layer1_outputs[6483] = ~((layer0_outputs[5640]) ^ (layer0_outputs[3747]));
    assign layer1_outputs[6484] = 1'b1;
    assign layer1_outputs[6485] = ~(layer0_outputs[1049]);
    assign layer1_outputs[6486] = layer0_outputs[1544];
    assign layer1_outputs[6487] = (layer0_outputs[2030]) & (layer0_outputs[2545]);
    assign layer1_outputs[6488] = ~((layer0_outputs[6505]) ^ (layer0_outputs[1076]));
    assign layer1_outputs[6489] = ~(layer0_outputs[5555]);
    assign layer1_outputs[6490] = ~(layer0_outputs[4073]);
    assign layer1_outputs[6491] = ~(layer0_outputs[11889]);
    assign layer1_outputs[6492] = (layer0_outputs[1243]) & ~(layer0_outputs[9958]);
    assign layer1_outputs[6493] = ~(layer0_outputs[347]) | (layer0_outputs[8285]);
    assign layer1_outputs[6494] = ~(layer0_outputs[8610]);
    assign layer1_outputs[6495] = (layer0_outputs[8740]) & ~(layer0_outputs[8857]);
    assign layer1_outputs[6496] = ~(layer0_outputs[9756]);
    assign layer1_outputs[6497] = ~(layer0_outputs[6455]) | (layer0_outputs[2637]);
    assign layer1_outputs[6498] = (layer0_outputs[12214]) ^ (layer0_outputs[3205]);
    assign layer1_outputs[6499] = ~(layer0_outputs[6512]);
    assign layer1_outputs[6500] = ~(layer0_outputs[3612]);
    assign layer1_outputs[6501] = (layer0_outputs[1188]) & ~(layer0_outputs[3143]);
    assign layer1_outputs[6502] = layer0_outputs[11134];
    assign layer1_outputs[6503] = layer0_outputs[1230];
    assign layer1_outputs[6504] = (layer0_outputs[5886]) & ~(layer0_outputs[8405]);
    assign layer1_outputs[6505] = ~(layer0_outputs[3498]);
    assign layer1_outputs[6506] = ~(layer0_outputs[9]);
    assign layer1_outputs[6507] = layer0_outputs[5871];
    assign layer1_outputs[6508] = (layer0_outputs[8606]) | (layer0_outputs[1901]);
    assign layer1_outputs[6509] = (layer0_outputs[8774]) & ~(layer0_outputs[9888]);
    assign layer1_outputs[6510] = ~(layer0_outputs[7758]);
    assign layer1_outputs[6511] = ~((layer0_outputs[8487]) ^ (layer0_outputs[1603]));
    assign layer1_outputs[6512] = ~(layer0_outputs[5479]);
    assign layer1_outputs[6513] = layer0_outputs[10836];
    assign layer1_outputs[6514] = (layer0_outputs[9663]) & ~(layer0_outputs[10475]);
    assign layer1_outputs[6515] = (layer0_outputs[7223]) & ~(layer0_outputs[5673]);
    assign layer1_outputs[6516] = ~(layer0_outputs[11642]) | (layer0_outputs[6613]);
    assign layer1_outputs[6517] = (layer0_outputs[9113]) & ~(layer0_outputs[7959]);
    assign layer1_outputs[6518] = ~(layer0_outputs[4066]);
    assign layer1_outputs[6519] = (layer0_outputs[11412]) ^ (layer0_outputs[3235]);
    assign layer1_outputs[6520] = layer0_outputs[5583];
    assign layer1_outputs[6521] = ~((layer0_outputs[2811]) ^ (layer0_outputs[269]));
    assign layer1_outputs[6522] = (layer0_outputs[4514]) | (layer0_outputs[9963]);
    assign layer1_outputs[6523] = layer0_outputs[5451];
    assign layer1_outputs[6524] = layer0_outputs[12704];
    assign layer1_outputs[6525] = ~(layer0_outputs[9156]);
    assign layer1_outputs[6526] = layer0_outputs[4694];
    assign layer1_outputs[6527] = (layer0_outputs[12765]) & (layer0_outputs[807]);
    assign layer1_outputs[6528] = ~((layer0_outputs[1231]) | (layer0_outputs[2328]));
    assign layer1_outputs[6529] = (layer0_outputs[11469]) & ~(layer0_outputs[8479]);
    assign layer1_outputs[6530] = 1'b0;
    assign layer1_outputs[6531] = (layer0_outputs[878]) & (layer0_outputs[8287]);
    assign layer1_outputs[6532] = ~((layer0_outputs[4609]) & (layer0_outputs[1521]));
    assign layer1_outputs[6533] = ~(layer0_outputs[12591]);
    assign layer1_outputs[6534] = (layer0_outputs[4100]) & ~(layer0_outputs[2575]);
    assign layer1_outputs[6535] = (layer0_outputs[12245]) & (layer0_outputs[6463]);
    assign layer1_outputs[6536] = ~((layer0_outputs[6124]) | (layer0_outputs[9240]));
    assign layer1_outputs[6537] = (layer0_outputs[6373]) & ~(layer0_outputs[184]);
    assign layer1_outputs[6538] = ~((layer0_outputs[869]) & (layer0_outputs[11924]));
    assign layer1_outputs[6539] = layer0_outputs[10479];
    assign layer1_outputs[6540] = ~((layer0_outputs[10691]) & (layer0_outputs[8070]));
    assign layer1_outputs[6541] = ~((layer0_outputs[5244]) ^ (layer0_outputs[6107]));
    assign layer1_outputs[6542] = ~(layer0_outputs[12791]) | (layer0_outputs[4220]);
    assign layer1_outputs[6543] = layer0_outputs[1215];
    assign layer1_outputs[6544] = layer0_outputs[3075];
    assign layer1_outputs[6545] = layer0_outputs[6042];
    assign layer1_outputs[6546] = ~((layer0_outputs[1023]) | (layer0_outputs[6628]));
    assign layer1_outputs[6547] = ~((layer0_outputs[342]) | (layer0_outputs[11527]));
    assign layer1_outputs[6548] = layer0_outputs[11626];
    assign layer1_outputs[6549] = 1'b0;
    assign layer1_outputs[6550] = layer0_outputs[4673];
    assign layer1_outputs[6551] = (layer0_outputs[3699]) ^ (layer0_outputs[10785]);
    assign layer1_outputs[6552] = ~((layer0_outputs[12025]) & (layer0_outputs[2518]));
    assign layer1_outputs[6553] = 1'b1;
    assign layer1_outputs[6554] = layer0_outputs[300];
    assign layer1_outputs[6555] = (layer0_outputs[1213]) | (layer0_outputs[9479]);
    assign layer1_outputs[6556] = (layer0_outputs[8850]) & ~(layer0_outputs[751]);
    assign layer1_outputs[6557] = ~((layer0_outputs[6976]) & (layer0_outputs[9637]));
    assign layer1_outputs[6558] = (layer0_outputs[11403]) & ~(layer0_outputs[9162]);
    assign layer1_outputs[6559] = (layer0_outputs[10218]) ^ (layer0_outputs[8099]);
    assign layer1_outputs[6560] = (layer0_outputs[938]) & ~(layer0_outputs[8067]);
    assign layer1_outputs[6561] = (layer0_outputs[5760]) & ~(layer0_outputs[94]);
    assign layer1_outputs[6562] = ~(layer0_outputs[9353]);
    assign layer1_outputs[6563] = ~(layer0_outputs[460]) | (layer0_outputs[10897]);
    assign layer1_outputs[6564] = layer0_outputs[8436];
    assign layer1_outputs[6565] = (layer0_outputs[2209]) & ~(layer0_outputs[4900]);
    assign layer1_outputs[6566] = layer0_outputs[3964];
    assign layer1_outputs[6567] = ~(layer0_outputs[9016]);
    assign layer1_outputs[6568] = (layer0_outputs[12008]) | (layer0_outputs[985]);
    assign layer1_outputs[6569] = layer0_outputs[9716];
    assign layer1_outputs[6570] = ~((layer0_outputs[7297]) | (layer0_outputs[7824]));
    assign layer1_outputs[6571] = ~(layer0_outputs[12347]);
    assign layer1_outputs[6572] = layer0_outputs[9666];
    assign layer1_outputs[6573] = ~(layer0_outputs[8967]);
    assign layer1_outputs[6574] = (layer0_outputs[1692]) & ~(layer0_outputs[3828]);
    assign layer1_outputs[6575] = ~((layer0_outputs[5887]) | (layer0_outputs[8815]));
    assign layer1_outputs[6576] = (layer0_outputs[6872]) & ~(layer0_outputs[7541]);
    assign layer1_outputs[6577] = (layer0_outputs[2049]) & ~(layer0_outputs[336]);
    assign layer1_outputs[6578] = ~((layer0_outputs[5856]) & (layer0_outputs[1744]));
    assign layer1_outputs[6579] = layer0_outputs[10307];
    assign layer1_outputs[6580] = layer0_outputs[12150];
    assign layer1_outputs[6581] = ~((layer0_outputs[7638]) & (layer0_outputs[6703]));
    assign layer1_outputs[6582] = ~(layer0_outputs[5724]);
    assign layer1_outputs[6583] = ~(layer0_outputs[4954]) | (layer0_outputs[9098]);
    assign layer1_outputs[6584] = (layer0_outputs[8342]) ^ (layer0_outputs[10409]);
    assign layer1_outputs[6585] = layer0_outputs[10404];
    assign layer1_outputs[6586] = ~(layer0_outputs[512]) | (layer0_outputs[1809]);
    assign layer1_outputs[6587] = (layer0_outputs[5971]) | (layer0_outputs[4574]);
    assign layer1_outputs[6588] = layer0_outputs[6390];
    assign layer1_outputs[6589] = ~((layer0_outputs[10619]) | (layer0_outputs[12326]));
    assign layer1_outputs[6590] = ~(layer0_outputs[3927]) | (layer0_outputs[11697]);
    assign layer1_outputs[6591] = ~(layer0_outputs[6447]) | (layer0_outputs[2383]);
    assign layer1_outputs[6592] = (layer0_outputs[9149]) | (layer0_outputs[9392]);
    assign layer1_outputs[6593] = ~(layer0_outputs[1224]);
    assign layer1_outputs[6594] = (layer0_outputs[4015]) ^ (layer0_outputs[11785]);
    assign layer1_outputs[6595] = 1'b1;
    assign layer1_outputs[6596] = (layer0_outputs[11126]) & ~(layer0_outputs[2615]);
    assign layer1_outputs[6597] = layer0_outputs[10259];
    assign layer1_outputs[6598] = ~((layer0_outputs[8685]) | (layer0_outputs[2090]));
    assign layer1_outputs[6599] = layer0_outputs[10085];
    assign layer1_outputs[6600] = (layer0_outputs[10383]) & ~(layer0_outputs[11940]);
    assign layer1_outputs[6601] = layer0_outputs[751];
    assign layer1_outputs[6602] = ~(layer0_outputs[1655]);
    assign layer1_outputs[6603] = (layer0_outputs[4101]) ^ (layer0_outputs[7659]);
    assign layer1_outputs[6604] = layer0_outputs[3244];
    assign layer1_outputs[6605] = (layer0_outputs[6818]) | (layer0_outputs[410]);
    assign layer1_outputs[6606] = ~(layer0_outputs[12405]) | (layer0_outputs[2345]);
    assign layer1_outputs[6607] = (layer0_outputs[3868]) ^ (layer0_outputs[2110]);
    assign layer1_outputs[6608] = (layer0_outputs[10631]) ^ (layer0_outputs[3282]);
    assign layer1_outputs[6609] = 1'b1;
    assign layer1_outputs[6610] = layer0_outputs[3900];
    assign layer1_outputs[6611] = layer0_outputs[2752];
    assign layer1_outputs[6612] = layer0_outputs[3963];
    assign layer1_outputs[6613] = ~(layer0_outputs[6966]) | (layer0_outputs[10351]);
    assign layer1_outputs[6614] = ~(layer0_outputs[989]);
    assign layer1_outputs[6615] = layer0_outputs[11402];
    assign layer1_outputs[6616] = ~(layer0_outputs[1051]) | (layer0_outputs[626]);
    assign layer1_outputs[6617] = layer0_outputs[8613];
    assign layer1_outputs[6618] = (layer0_outputs[10726]) & (layer0_outputs[3119]);
    assign layer1_outputs[6619] = (layer0_outputs[9195]) & (layer0_outputs[7713]);
    assign layer1_outputs[6620] = ~((layer0_outputs[3797]) | (layer0_outputs[1453]));
    assign layer1_outputs[6621] = ~(layer0_outputs[1708]);
    assign layer1_outputs[6622] = ~(layer0_outputs[2837]);
    assign layer1_outputs[6623] = ~(layer0_outputs[7289]);
    assign layer1_outputs[6624] = layer0_outputs[6908];
    assign layer1_outputs[6625] = 1'b1;
    assign layer1_outputs[6626] = ~((layer0_outputs[2710]) ^ (layer0_outputs[9596]));
    assign layer1_outputs[6627] = (layer0_outputs[11587]) | (layer0_outputs[4365]);
    assign layer1_outputs[6628] = ~(layer0_outputs[36]) | (layer0_outputs[9097]);
    assign layer1_outputs[6629] = ~(layer0_outputs[4316]) | (layer0_outputs[2219]);
    assign layer1_outputs[6630] = ~((layer0_outputs[4948]) | (layer0_outputs[6267]));
    assign layer1_outputs[6631] = ~(layer0_outputs[7119]) | (layer0_outputs[1616]);
    assign layer1_outputs[6632] = layer0_outputs[10680];
    assign layer1_outputs[6633] = ~(layer0_outputs[9476]);
    assign layer1_outputs[6634] = ~(layer0_outputs[1040]);
    assign layer1_outputs[6635] = ~(layer0_outputs[2575]) | (layer0_outputs[4858]);
    assign layer1_outputs[6636] = ~(layer0_outputs[10325]);
    assign layer1_outputs[6637] = ~(layer0_outputs[7398]) | (layer0_outputs[9603]);
    assign layer1_outputs[6638] = ~((layer0_outputs[6552]) & (layer0_outputs[1939]));
    assign layer1_outputs[6639] = (layer0_outputs[9893]) & (layer0_outputs[10052]);
    assign layer1_outputs[6640] = (layer0_outputs[3023]) | (layer0_outputs[3509]);
    assign layer1_outputs[6641] = layer0_outputs[6753];
    assign layer1_outputs[6642] = ~(layer0_outputs[8734]) | (layer0_outputs[355]);
    assign layer1_outputs[6643] = ~(layer0_outputs[10565]);
    assign layer1_outputs[6644] = layer0_outputs[3206];
    assign layer1_outputs[6645] = layer0_outputs[4033];
    assign layer1_outputs[6646] = layer0_outputs[8992];
    assign layer1_outputs[6647] = (layer0_outputs[7405]) | (layer0_outputs[8329]);
    assign layer1_outputs[6648] = ~((layer0_outputs[3186]) & (layer0_outputs[11218]));
    assign layer1_outputs[6649] = layer0_outputs[12386];
    assign layer1_outputs[6650] = ~((layer0_outputs[160]) & (layer0_outputs[6787]));
    assign layer1_outputs[6651] = ~(layer0_outputs[8437]) | (layer0_outputs[654]);
    assign layer1_outputs[6652] = 1'b1;
    assign layer1_outputs[6653] = layer0_outputs[6113];
    assign layer1_outputs[6654] = ~((layer0_outputs[7345]) & (layer0_outputs[5801]));
    assign layer1_outputs[6655] = layer0_outputs[4421];
    assign layer1_outputs[6656] = (layer0_outputs[9591]) ^ (layer0_outputs[3727]);
    assign layer1_outputs[6657] = ~((layer0_outputs[790]) & (layer0_outputs[6412]));
    assign layer1_outputs[6658] = ~((layer0_outputs[6026]) | (layer0_outputs[5343]));
    assign layer1_outputs[6659] = ~(layer0_outputs[8752]);
    assign layer1_outputs[6660] = ~((layer0_outputs[5994]) & (layer0_outputs[3901]));
    assign layer1_outputs[6661] = ~((layer0_outputs[2582]) | (layer0_outputs[10634]));
    assign layer1_outputs[6662] = ~(layer0_outputs[4930]);
    assign layer1_outputs[6663] = ~((layer0_outputs[5323]) ^ (layer0_outputs[2088]));
    assign layer1_outputs[6664] = ~(layer0_outputs[11344]);
    assign layer1_outputs[6665] = (layer0_outputs[988]) & ~(layer0_outputs[1853]);
    assign layer1_outputs[6666] = layer0_outputs[372];
    assign layer1_outputs[6667] = (layer0_outputs[8133]) ^ (layer0_outputs[4530]);
    assign layer1_outputs[6668] = (layer0_outputs[1861]) & ~(layer0_outputs[2507]);
    assign layer1_outputs[6669] = 1'b0;
    assign layer1_outputs[6670] = layer0_outputs[12572];
    assign layer1_outputs[6671] = layer0_outputs[6075];
    assign layer1_outputs[6672] = layer0_outputs[11352];
    assign layer1_outputs[6673] = ~((layer0_outputs[2670]) & (layer0_outputs[12027]));
    assign layer1_outputs[6674] = ~((layer0_outputs[9358]) & (layer0_outputs[938]));
    assign layer1_outputs[6675] = ~(layer0_outputs[722]);
    assign layer1_outputs[6676] = layer0_outputs[4014];
    assign layer1_outputs[6677] = layer0_outputs[5183];
    assign layer1_outputs[6678] = layer0_outputs[638];
    assign layer1_outputs[6679] = ~(layer0_outputs[328]) | (layer0_outputs[1559]);
    assign layer1_outputs[6680] = ~(layer0_outputs[12505]) | (layer0_outputs[6255]);
    assign layer1_outputs[6681] = (layer0_outputs[12414]) ^ (layer0_outputs[1175]);
    assign layer1_outputs[6682] = (layer0_outputs[8109]) & (layer0_outputs[10699]);
    assign layer1_outputs[6683] = (layer0_outputs[256]) & (layer0_outputs[3037]);
    assign layer1_outputs[6684] = ~((layer0_outputs[11538]) ^ (layer0_outputs[5223]));
    assign layer1_outputs[6685] = ~(layer0_outputs[9179]);
    assign layer1_outputs[6686] = (layer0_outputs[10526]) & ~(layer0_outputs[11965]);
    assign layer1_outputs[6687] = layer0_outputs[2824];
    assign layer1_outputs[6688] = (layer0_outputs[10072]) & ~(layer0_outputs[11042]);
    assign layer1_outputs[6689] = (layer0_outputs[5635]) & ~(layer0_outputs[12678]);
    assign layer1_outputs[6690] = (layer0_outputs[5261]) & (layer0_outputs[8696]);
    assign layer1_outputs[6691] = ~((layer0_outputs[7736]) & (layer0_outputs[6694]));
    assign layer1_outputs[6692] = ~(layer0_outputs[21]) | (layer0_outputs[3908]);
    assign layer1_outputs[6693] = ~(layer0_outputs[1730]);
    assign layer1_outputs[6694] = (layer0_outputs[1393]) | (layer0_outputs[12441]);
    assign layer1_outputs[6695] = layer0_outputs[6800];
    assign layer1_outputs[6696] = ~((layer0_outputs[4396]) | (layer0_outputs[2854]));
    assign layer1_outputs[6697] = layer0_outputs[2427];
    assign layer1_outputs[6698] = ~(layer0_outputs[4196]);
    assign layer1_outputs[6699] = 1'b0;
    assign layer1_outputs[6700] = ~((layer0_outputs[10748]) | (layer0_outputs[2901]));
    assign layer1_outputs[6701] = ~(layer0_outputs[7152]);
    assign layer1_outputs[6702] = (layer0_outputs[8432]) | (layer0_outputs[9304]);
    assign layer1_outputs[6703] = layer0_outputs[11144];
    assign layer1_outputs[6704] = (layer0_outputs[9347]) & (layer0_outputs[146]);
    assign layer1_outputs[6705] = ~((layer0_outputs[3144]) ^ (layer0_outputs[850]));
    assign layer1_outputs[6706] = (layer0_outputs[1716]) | (layer0_outputs[8959]);
    assign layer1_outputs[6707] = ~(layer0_outputs[5250]) | (layer0_outputs[10267]);
    assign layer1_outputs[6708] = ~(layer0_outputs[9141]);
    assign layer1_outputs[6709] = (layer0_outputs[8565]) & (layer0_outputs[3381]);
    assign layer1_outputs[6710] = ~((layer0_outputs[12098]) | (layer0_outputs[6406]));
    assign layer1_outputs[6711] = (layer0_outputs[2035]) & (layer0_outputs[619]);
    assign layer1_outputs[6712] = ~(layer0_outputs[9420]);
    assign layer1_outputs[6713] = (layer0_outputs[7169]) & (layer0_outputs[9626]);
    assign layer1_outputs[6714] = layer0_outputs[6786];
    assign layer1_outputs[6715] = layer0_outputs[11095];
    assign layer1_outputs[6716] = (layer0_outputs[12445]) ^ (layer0_outputs[4382]);
    assign layer1_outputs[6717] = layer0_outputs[8253];
    assign layer1_outputs[6718] = layer0_outputs[10086];
    assign layer1_outputs[6719] = layer0_outputs[2833];
    assign layer1_outputs[6720] = (layer0_outputs[1770]) ^ (layer0_outputs[6644]);
    assign layer1_outputs[6721] = ~(layer0_outputs[8210]);
    assign layer1_outputs[6722] = ~((layer0_outputs[666]) & (layer0_outputs[9769]));
    assign layer1_outputs[6723] = (layer0_outputs[10918]) & ~(layer0_outputs[8333]);
    assign layer1_outputs[6724] = ~((layer0_outputs[9697]) ^ (layer0_outputs[6933]));
    assign layer1_outputs[6725] = (layer0_outputs[12298]) | (layer0_outputs[8505]);
    assign layer1_outputs[6726] = ~((layer0_outputs[11232]) & (layer0_outputs[3444]));
    assign layer1_outputs[6727] = layer0_outputs[527];
    assign layer1_outputs[6728] = (layer0_outputs[11277]) & ~(layer0_outputs[3574]);
    assign layer1_outputs[6729] = (layer0_outputs[2299]) & (layer0_outputs[11221]);
    assign layer1_outputs[6730] = layer0_outputs[10002];
    assign layer1_outputs[6731] = ~(layer0_outputs[413]);
    assign layer1_outputs[6732] = (layer0_outputs[10258]) & ~(layer0_outputs[7274]);
    assign layer1_outputs[6733] = layer0_outputs[26];
    assign layer1_outputs[6734] = ~(layer0_outputs[3009]);
    assign layer1_outputs[6735] = ~(layer0_outputs[11680]) | (layer0_outputs[3627]);
    assign layer1_outputs[6736] = (layer0_outputs[11483]) | (layer0_outputs[9166]);
    assign layer1_outputs[6737] = ~(layer0_outputs[1586]);
    assign layer1_outputs[6738] = ~(layer0_outputs[3624]) | (layer0_outputs[8002]);
    assign layer1_outputs[6739] = (layer0_outputs[1121]) & (layer0_outputs[1206]);
    assign layer1_outputs[6740] = (layer0_outputs[7849]) & ~(layer0_outputs[12409]);
    assign layer1_outputs[6741] = layer0_outputs[3313];
    assign layer1_outputs[6742] = layer0_outputs[1816];
    assign layer1_outputs[6743] = ~(layer0_outputs[11219]) | (layer0_outputs[9436]);
    assign layer1_outputs[6744] = ~((layer0_outputs[451]) | (layer0_outputs[2282]));
    assign layer1_outputs[6745] = (layer0_outputs[794]) | (layer0_outputs[3909]);
    assign layer1_outputs[6746] = 1'b1;
    assign layer1_outputs[6747] = ~(layer0_outputs[9758]) | (layer0_outputs[12548]);
    assign layer1_outputs[6748] = ~((layer0_outputs[5116]) ^ (layer0_outputs[10998]));
    assign layer1_outputs[6749] = ~(layer0_outputs[477]);
    assign layer1_outputs[6750] = (layer0_outputs[2897]) & ~(layer0_outputs[680]);
    assign layer1_outputs[6751] = layer0_outputs[2828];
    assign layer1_outputs[6752] = (layer0_outputs[3534]) | (layer0_outputs[1612]);
    assign layer1_outputs[6753] = ~(layer0_outputs[4174]);
    assign layer1_outputs[6754] = ~(layer0_outputs[4832]);
    assign layer1_outputs[6755] = (layer0_outputs[9224]) | (layer0_outputs[1210]);
    assign layer1_outputs[6756] = (layer0_outputs[3137]) ^ (layer0_outputs[7212]);
    assign layer1_outputs[6757] = ~(layer0_outputs[5227]) | (layer0_outputs[5739]);
    assign layer1_outputs[6758] = (layer0_outputs[10856]) & (layer0_outputs[10415]);
    assign layer1_outputs[6759] = layer0_outputs[8848];
    assign layer1_outputs[6760] = (layer0_outputs[11941]) & ~(layer0_outputs[5561]);
    assign layer1_outputs[6761] = (layer0_outputs[10254]) | (layer0_outputs[10442]);
    assign layer1_outputs[6762] = ~(layer0_outputs[8530]) | (layer0_outputs[12717]);
    assign layer1_outputs[6763] = (layer0_outputs[3854]) | (layer0_outputs[11834]);
    assign layer1_outputs[6764] = layer0_outputs[3114];
    assign layer1_outputs[6765] = layer0_outputs[5422];
    assign layer1_outputs[6766] = (layer0_outputs[8288]) & ~(layer0_outputs[7231]);
    assign layer1_outputs[6767] = (layer0_outputs[9215]) & (layer0_outputs[2722]);
    assign layer1_outputs[6768] = (layer0_outputs[6667]) ^ (layer0_outputs[7866]);
    assign layer1_outputs[6769] = ~(layer0_outputs[11130]) | (layer0_outputs[3644]);
    assign layer1_outputs[6770] = 1'b0;
    assign layer1_outputs[6771] = ~(layer0_outputs[10443]) | (layer0_outputs[9688]);
    assign layer1_outputs[6772] = ~((layer0_outputs[6795]) & (layer0_outputs[3421]));
    assign layer1_outputs[6773] = (layer0_outputs[313]) & (layer0_outputs[5171]);
    assign layer1_outputs[6774] = ~(layer0_outputs[10603]);
    assign layer1_outputs[6775] = layer0_outputs[3032];
    assign layer1_outputs[6776] = layer0_outputs[4117];
    assign layer1_outputs[6777] = layer0_outputs[12471];
    assign layer1_outputs[6778] = ~(layer0_outputs[545]);
    assign layer1_outputs[6779] = layer0_outputs[1926];
    assign layer1_outputs[6780] = ~((layer0_outputs[924]) & (layer0_outputs[1037]));
    assign layer1_outputs[6781] = ~(layer0_outputs[3179]) | (layer0_outputs[2311]);
    assign layer1_outputs[6782] = ~(layer0_outputs[5637]);
    assign layer1_outputs[6783] = layer0_outputs[6683];
    assign layer1_outputs[6784] = ~(layer0_outputs[7885]);
    assign layer1_outputs[6785] = layer0_outputs[10069];
    assign layer1_outputs[6786] = ~((layer0_outputs[5935]) | (layer0_outputs[2040]));
    assign layer1_outputs[6787] = (layer0_outputs[12528]) & ~(layer0_outputs[5863]);
    assign layer1_outputs[6788] = layer0_outputs[5431];
    assign layer1_outputs[6789] = (layer0_outputs[5783]) & (layer0_outputs[2131]);
    assign layer1_outputs[6790] = ~(layer0_outputs[1264]) | (layer0_outputs[5356]);
    assign layer1_outputs[6791] = (layer0_outputs[9617]) ^ (layer0_outputs[5455]);
    assign layer1_outputs[6792] = ~((layer0_outputs[11891]) & (layer0_outputs[8814]));
    assign layer1_outputs[6793] = (layer0_outputs[837]) ^ (layer0_outputs[10698]);
    assign layer1_outputs[6794] = layer0_outputs[3089];
    assign layer1_outputs[6795] = ~(layer0_outputs[425]);
    assign layer1_outputs[6796] = ~(layer0_outputs[1058]);
    assign layer1_outputs[6797] = ~(layer0_outputs[4444]);
    assign layer1_outputs[6798] = layer0_outputs[3394];
    assign layer1_outputs[6799] = ~(layer0_outputs[11123]);
    assign layer1_outputs[6800] = ~(layer0_outputs[6357]);
    assign layer1_outputs[6801] = ~(layer0_outputs[767]);
    assign layer1_outputs[6802] = (layer0_outputs[653]) & ~(layer0_outputs[899]);
    assign layer1_outputs[6803] = (layer0_outputs[12572]) & ~(layer0_outputs[6784]);
    assign layer1_outputs[6804] = ~(layer0_outputs[3098]);
    assign layer1_outputs[6805] = (layer0_outputs[53]) & ~(layer0_outputs[9872]);
    assign layer1_outputs[6806] = (layer0_outputs[4274]) | (layer0_outputs[8135]);
    assign layer1_outputs[6807] = layer0_outputs[1221];
    assign layer1_outputs[6808] = layer0_outputs[10950];
    assign layer1_outputs[6809] = ~(layer0_outputs[2934]);
    assign layer1_outputs[6810] = layer0_outputs[8563];
    assign layer1_outputs[6811] = ~(layer0_outputs[9641]);
    assign layer1_outputs[6812] = (layer0_outputs[7051]) & (layer0_outputs[7742]);
    assign layer1_outputs[6813] = ~((layer0_outputs[9005]) | (layer0_outputs[9205]));
    assign layer1_outputs[6814] = (layer0_outputs[4224]) ^ (layer0_outputs[772]);
    assign layer1_outputs[6815] = ~(layer0_outputs[7901]);
    assign layer1_outputs[6816] = layer0_outputs[8667];
    assign layer1_outputs[6817] = (layer0_outputs[7477]) & ~(layer0_outputs[2072]);
    assign layer1_outputs[6818] = (layer0_outputs[8103]) & ~(layer0_outputs[5885]);
    assign layer1_outputs[6819] = layer0_outputs[2679];
    assign layer1_outputs[6820] = ~(layer0_outputs[2354]);
    assign layer1_outputs[6821] = ~(layer0_outputs[6537]);
    assign layer1_outputs[6822] = (layer0_outputs[3672]) & ~(layer0_outputs[6369]);
    assign layer1_outputs[6823] = ~(layer0_outputs[3642]);
    assign layer1_outputs[6824] = (layer0_outputs[6481]) & (layer0_outputs[7486]);
    assign layer1_outputs[6825] = ~((layer0_outputs[9932]) & (layer0_outputs[839]));
    assign layer1_outputs[6826] = ~(layer0_outputs[7589]);
    assign layer1_outputs[6827] = layer0_outputs[9165];
    assign layer1_outputs[6828] = ~(layer0_outputs[9488]) | (layer0_outputs[5641]);
    assign layer1_outputs[6829] = (layer0_outputs[6177]) | (layer0_outputs[4186]);
    assign layer1_outputs[6830] = ~(layer0_outputs[2742]);
    assign layer1_outputs[6831] = ~(layer0_outputs[10948]) | (layer0_outputs[2020]);
    assign layer1_outputs[6832] = (layer0_outputs[750]) ^ (layer0_outputs[10718]);
    assign layer1_outputs[6833] = ~((layer0_outputs[6668]) & (layer0_outputs[2396]));
    assign layer1_outputs[6834] = ~(layer0_outputs[9615]);
    assign layer1_outputs[6835] = ~((layer0_outputs[8870]) | (layer0_outputs[652]));
    assign layer1_outputs[6836] = ~(layer0_outputs[603]) | (layer0_outputs[5508]);
    assign layer1_outputs[6837] = ~(layer0_outputs[11419]) | (layer0_outputs[7044]);
    assign layer1_outputs[6838] = ~(layer0_outputs[3339]);
    assign layer1_outputs[6839] = ~(layer0_outputs[2116]) | (layer0_outputs[11364]);
    assign layer1_outputs[6840] = ~(layer0_outputs[7912]) | (layer0_outputs[7879]);
    assign layer1_outputs[6841] = ~(layer0_outputs[9696]) | (layer0_outputs[5894]);
    assign layer1_outputs[6842] = ~(layer0_outputs[2524]) | (layer0_outputs[7579]);
    assign layer1_outputs[6843] = layer0_outputs[8041];
    assign layer1_outputs[6844] = (layer0_outputs[5721]) & (layer0_outputs[1796]);
    assign layer1_outputs[6845] = (layer0_outputs[3870]) ^ (layer0_outputs[8542]);
    assign layer1_outputs[6846] = ~(layer0_outputs[539]) | (layer0_outputs[9038]);
    assign layer1_outputs[6847] = (layer0_outputs[12352]) | (layer0_outputs[2480]);
    assign layer1_outputs[6848] = ~((layer0_outputs[850]) | (layer0_outputs[1050]));
    assign layer1_outputs[6849] = ~(layer0_outputs[3300]);
    assign layer1_outputs[6850] = ~(layer0_outputs[6565]);
    assign layer1_outputs[6851] = (layer0_outputs[6868]) | (layer0_outputs[6805]);
    assign layer1_outputs[6852] = (layer0_outputs[11421]) & ~(layer0_outputs[5439]);
    assign layer1_outputs[6853] = ~(layer0_outputs[1572]) | (layer0_outputs[9395]);
    assign layer1_outputs[6854] = ~((layer0_outputs[10880]) & (layer0_outputs[12575]));
    assign layer1_outputs[6855] = layer0_outputs[10682];
    assign layer1_outputs[6856] = (layer0_outputs[3637]) & ~(layer0_outputs[12009]);
    assign layer1_outputs[6857] = layer0_outputs[7000];
    assign layer1_outputs[6858] = ~(layer0_outputs[11724]);
    assign layer1_outputs[6859] = ~((layer0_outputs[11896]) & (layer0_outputs[9531]));
    assign layer1_outputs[6860] = 1'b0;
    assign layer1_outputs[6861] = layer0_outputs[6828];
    assign layer1_outputs[6862] = (layer0_outputs[11758]) & ~(layer0_outputs[9714]);
    assign layer1_outputs[6863] = ~((layer0_outputs[8451]) & (layer0_outputs[9002]));
    assign layer1_outputs[6864] = ~(layer0_outputs[8343]);
    assign layer1_outputs[6865] = layer0_outputs[2159];
    assign layer1_outputs[6866] = ~(layer0_outputs[8855]) | (layer0_outputs[1516]);
    assign layer1_outputs[6867] = ~(layer0_outputs[10311]);
    assign layer1_outputs[6868] = layer0_outputs[9640];
    assign layer1_outputs[6869] = layer0_outputs[8754];
    assign layer1_outputs[6870] = (layer0_outputs[1192]) & (layer0_outputs[8460]);
    assign layer1_outputs[6871] = layer0_outputs[875];
    assign layer1_outputs[6872] = ~(layer0_outputs[1125]);
    assign layer1_outputs[6873] = (layer0_outputs[6968]) | (layer0_outputs[10344]);
    assign layer1_outputs[6874] = ~(layer0_outputs[8353]) | (layer0_outputs[11480]);
    assign layer1_outputs[6875] = ~(layer0_outputs[7652]) | (layer0_outputs[9766]);
    assign layer1_outputs[6876] = (layer0_outputs[3893]) & ~(layer0_outputs[6207]);
    assign layer1_outputs[6877] = ~(layer0_outputs[12294]);
    assign layer1_outputs[6878] = ~((layer0_outputs[7639]) & (layer0_outputs[1674]));
    assign layer1_outputs[6879] = (layer0_outputs[8765]) | (layer0_outputs[5257]);
    assign layer1_outputs[6880] = layer0_outputs[6426];
    assign layer1_outputs[6881] = (layer0_outputs[4493]) & ~(layer0_outputs[9296]);
    assign layer1_outputs[6882] = ~(layer0_outputs[1253]) | (layer0_outputs[7041]);
    assign layer1_outputs[6883] = ~(layer0_outputs[4149]) | (layer0_outputs[9415]);
    assign layer1_outputs[6884] = (layer0_outputs[9064]) & ~(layer0_outputs[6783]);
    assign layer1_outputs[6885] = ~((layer0_outputs[5578]) ^ (layer0_outputs[2643]));
    assign layer1_outputs[6886] = (layer0_outputs[9378]) | (layer0_outputs[10836]);
    assign layer1_outputs[6887] = ~((layer0_outputs[12713]) ^ (layer0_outputs[3571]));
    assign layer1_outputs[6888] = ~((layer0_outputs[5843]) & (layer0_outputs[7634]));
    assign layer1_outputs[6889] = (layer0_outputs[10140]) & ~(layer0_outputs[7158]);
    assign layer1_outputs[6890] = ~((layer0_outputs[2685]) | (layer0_outputs[1032]));
    assign layer1_outputs[6891] = ~(layer0_outputs[4095]);
    assign layer1_outputs[6892] = ~(layer0_outputs[10437]);
    assign layer1_outputs[6893] = ~(layer0_outputs[5975]);
    assign layer1_outputs[6894] = ~(layer0_outputs[11877]);
    assign layer1_outputs[6895] = layer0_outputs[1110];
    assign layer1_outputs[6896] = layer0_outputs[8501];
    assign layer1_outputs[6897] = (layer0_outputs[4768]) | (layer0_outputs[1108]);
    assign layer1_outputs[6898] = (layer0_outputs[4851]) ^ (layer0_outputs[9336]);
    assign layer1_outputs[6899] = layer0_outputs[10048];
    assign layer1_outputs[6900] = ~(layer0_outputs[2745]);
    assign layer1_outputs[6901] = ~((layer0_outputs[4392]) & (layer0_outputs[4921]));
    assign layer1_outputs[6902] = layer0_outputs[5350];
    assign layer1_outputs[6903] = ~((layer0_outputs[3757]) | (layer0_outputs[52]));
    assign layer1_outputs[6904] = ~(layer0_outputs[9727]) | (layer0_outputs[442]);
    assign layer1_outputs[6905] = 1'b0;
    assign layer1_outputs[6906] = (layer0_outputs[7035]) & ~(layer0_outputs[3749]);
    assign layer1_outputs[6907] = layer0_outputs[11768];
    assign layer1_outputs[6908] = ~((layer0_outputs[8880]) | (layer0_outputs[12280]));
    assign layer1_outputs[6909] = (layer0_outputs[12323]) ^ (layer0_outputs[5962]);
    assign layer1_outputs[6910] = layer0_outputs[229];
    assign layer1_outputs[6911] = (layer0_outputs[7994]) & (layer0_outputs[12357]);
    assign layer1_outputs[6912] = ~((layer0_outputs[6992]) | (layer0_outputs[1110]));
    assign layer1_outputs[6913] = ~(layer0_outputs[7005]) | (layer0_outputs[12448]);
    assign layer1_outputs[6914] = (layer0_outputs[6891]) & (layer0_outputs[12639]);
    assign layer1_outputs[6915] = ~((layer0_outputs[9326]) & (layer0_outputs[11936]));
    assign layer1_outputs[6916] = (layer0_outputs[5977]) | (layer0_outputs[1395]);
    assign layer1_outputs[6917] = ~((layer0_outputs[7332]) ^ (layer0_outputs[8732]));
    assign layer1_outputs[6918] = layer0_outputs[4686];
    assign layer1_outputs[6919] = (layer0_outputs[10278]) & ~(layer0_outputs[10950]);
    assign layer1_outputs[6920] = (layer0_outputs[1071]) & ~(layer0_outputs[6980]);
    assign layer1_outputs[6921] = ~(layer0_outputs[3990]);
    assign layer1_outputs[6922] = ~((layer0_outputs[3177]) | (layer0_outputs[6787]));
    assign layer1_outputs[6923] = layer0_outputs[8796];
    assign layer1_outputs[6924] = layer0_outputs[10445];
    assign layer1_outputs[6925] = ~((layer0_outputs[8124]) & (layer0_outputs[7042]));
    assign layer1_outputs[6926] = ~(layer0_outputs[10248]);
    assign layer1_outputs[6927] = ~(layer0_outputs[2671]);
    assign layer1_outputs[6928] = layer0_outputs[7770];
    assign layer1_outputs[6929] = (layer0_outputs[1309]) ^ (layer0_outputs[3086]);
    assign layer1_outputs[6930] = ~((layer0_outputs[10056]) & (layer0_outputs[8151]));
    assign layer1_outputs[6931] = ~((layer0_outputs[11206]) ^ (layer0_outputs[7505]));
    assign layer1_outputs[6932] = ~((layer0_outputs[12761]) & (layer0_outputs[8296]));
    assign layer1_outputs[6933] = ~((layer0_outputs[3940]) ^ (layer0_outputs[1314]));
    assign layer1_outputs[6934] = ~(layer0_outputs[6897]) | (layer0_outputs[11227]);
    assign layer1_outputs[6935] = layer0_outputs[8951];
    assign layer1_outputs[6936] = ~(layer0_outputs[4775]);
    assign layer1_outputs[6937] = ~(layer0_outputs[502]);
    assign layer1_outputs[6938] = 1'b1;
    assign layer1_outputs[6939] = layer0_outputs[1481];
    assign layer1_outputs[6940] = ~(layer0_outputs[1923]) | (layer0_outputs[8015]);
    assign layer1_outputs[6941] = (layer0_outputs[2132]) | (layer0_outputs[11414]);
    assign layer1_outputs[6942] = (layer0_outputs[2309]) ^ (layer0_outputs[11307]);
    assign layer1_outputs[6943] = (layer0_outputs[8374]) & ~(layer0_outputs[12178]);
    assign layer1_outputs[6944] = 1'b1;
    assign layer1_outputs[6945] = ~(layer0_outputs[10978]) | (layer0_outputs[1138]);
    assign layer1_outputs[6946] = ~(layer0_outputs[10467]) | (layer0_outputs[10272]);
    assign layer1_outputs[6947] = ~(layer0_outputs[3766]);
    assign layer1_outputs[6948] = ~((layer0_outputs[9782]) & (layer0_outputs[1151]));
    assign layer1_outputs[6949] = ~((layer0_outputs[7680]) & (layer0_outputs[7701]));
    assign layer1_outputs[6950] = ~(layer0_outputs[7633]);
    assign layer1_outputs[6951] = ~((layer0_outputs[11303]) | (layer0_outputs[9190]));
    assign layer1_outputs[6952] = (layer0_outputs[1643]) & ~(layer0_outputs[1870]);
    assign layer1_outputs[6953] = ~(layer0_outputs[12787]);
    assign layer1_outputs[6954] = (layer0_outputs[2620]) & ~(layer0_outputs[5671]);
    assign layer1_outputs[6955] = layer0_outputs[4528];
    assign layer1_outputs[6956] = ~((layer0_outputs[4243]) & (layer0_outputs[2520]));
    assign layer1_outputs[6957] = ~(layer0_outputs[11302]);
    assign layer1_outputs[6958] = (layer0_outputs[3497]) & (layer0_outputs[11579]);
    assign layer1_outputs[6959] = (layer0_outputs[9218]) ^ (layer0_outputs[2180]);
    assign layer1_outputs[6960] = (layer0_outputs[8102]) & ~(layer0_outputs[11437]);
    assign layer1_outputs[6961] = (layer0_outputs[10057]) & (layer0_outputs[10265]);
    assign layer1_outputs[6962] = ~((layer0_outputs[11832]) & (layer0_outputs[4013]));
    assign layer1_outputs[6963] = 1'b0;
    assign layer1_outputs[6964] = 1'b1;
    assign layer1_outputs[6965] = (layer0_outputs[4858]) & (layer0_outputs[2002]);
    assign layer1_outputs[6966] = ~(layer0_outputs[8883]);
    assign layer1_outputs[6967] = layer0_outputs[11644];
    assign layer1_outputs[6968] = ~(layer0_outputs[4834]) | (layer0_outputs[12770]);
    assign layer1_outputs[6969] = layer0_outputs[10071];
    assign layer1_outputs[6970] = (layer0_outputs[12183]) & ~(layer0_outputs[10274]);
    assign layer1_outputs[6971] = (layer0_outputs[6965]) ^ (layer0_outputs[7099]);
    assign layer1_outputs[6972] = (layer0_outputs[4628]) ^ (layer0_outputs[2426]);
    assign layer1_outputs[6973] = layer0_outputs[5631];
    assign layer1_outputs[6974] = (layer0_outputs[4246]) | (layer0_outputs[396]);
    assign layer1_outputs[6975] = (layer0_outputs[7582]) & ~(layer0_outputs[11995]);
    assign layer1_outputs[6976] = (layer0_outputs[12127]) ^ (layer0_outputs[8657]);
    assign layer1_outputs[6977] = ~((layer0_outputs[4875]) ^ (layer0_outputs[9975]));
    assign layer1_outputs[6978] = (layer0_outputs[10543]) & ~(layer0_outputs[4045]);
    assign layer1_outputs[6979] = ~(layer0_outputs[12578]) | (layer0_outputs[8686]);
    assign layer1_outputs[6980] = ~(layer0_outputs[2248]) | (layer0_outputs[6014]);
    assign layer1_outputs[6981] = ~(layer0_outputs[10363]);
    assign layer1_outputs[6982] = (layer0_outputs[11405]) & ~(layer0_outputs[6586]);
    assign layer1_outputs[6983] = 1'b0;
    assign layer1_outputs[6984] = (layer0_outputs[1530]) ^ (layer0_outputs[5577]);
    assign layer1_outputs[6985] = ~((layer0_outputs[4835]) | (layer0_outputs[614]));
    assign layer1_outputs[6986] = ~(layer0_outputs[4157]);
    assign layer1_outputs[6987] = (layer0_outputs[10430]) & ~(layer0_outputs[2179]);
    assign layer1_outputs[6988] = ~((layer0_outputs[10113]) & (layer0_outputs[1892]));
    assign layer1_outputs[6989] = ~((layer0_outputs[9128]) | (layer0_outputs[3718]));
    assign layer1_outputs[6990] = (layer0_outputs[11779]) & (layer0_outputs[5282]);
    assign layer1_outputs[6991] = (layer0_outputs[10317]) & ~(layer0_outputs[3184]);
    assign layer1_outputs[6992] = (layer0_outputs[5420]) & ~(layer0_outputs[11821]);
    assign layer1_outputs[6993] = (layer0_outputs[2201]) & ~(layer0_outputs[10824]);
    assign layer1_outputs[6994] = (layer0_outputs[7439]) & ~(layer0_outputs[9847]);
    assign layer1_outputs[6995] = ~(layer0_outputs[10563]);
    assign layer1_outputs[6996] = (layer0_outputs[6593]) & ~(layer0_outputs[10043]);
    assign layer1_outputs[6997] = (layer0_outputs[8112]) & (layer0_outputs[9018]);
    assign layer1_outputs[6998] = (layer0_outputs[12421]) ^ (layer0_outputs[7151]);
    assign layer1_outputs[6999] = ~(layer0_outputs[4566]);
    assign layer1_outputs[7000] = (layer0_outputs[5252]) & ~(layer0_outputs[6884]);
    assign layer1_outputs[7001] = ~((layer0_outputs[9643]) | (layer0_outputs[6925]));
    assign layer1_outputs[7002] = ~(layer0_outputs[7491]);
    assign layer1_outputs[7003] = ~(layer0_outputs[11784]);
    assign layer1_outputs[7004] = ~((layer0_outputs[8562]) & (layer0_outputs[10714]));
    assign layer1_outputs[7005] = layer0_outputs[3619];
    assign layer1_outputs[7006] = layer0_outputs[1897];
    assign layer1_outputs[7007] = 1'b0;
    assign layer1_outputs[7008] = ~(layer0_outputs[2815]);
    assign layer1_outputs[7009] = ~(layer0_outputs[3969]);
    assign layer1_outputs[7010] = ~((layer0_outputs[12586]) & (layer0_outputs[2150]));
    assign layer1_outputs[7011] = ~(layer0_outputs[2855]);
    assign layer1_outputs[7012] = (layer0_outputs[5743]) & ~(layer0_outputs[11704]);
    assign layer1_outputs[7013] = (layer0_outputs[8807]) & (layer0_outputs[519]);
    assign layer1_outputs[7014] = (layer0_outputs[9076]) | (layer0_outputs[9143]);
    assign layer1_outputs[7015] = ~(layer0_outputs[4133]) | (layer0_outputs[6976]);
    assign layer1_outputs[7016] = ~(layer0_outputs[5166]) | (layer0_outputs[1288]);
    assign layer1_outputs[7017] = (layer0_outputs[3119]) | (layer0_outputs[3652]);
    assign layer1_outputs[7018] = ~((layer0_outputs[6889]) ^ (layer0_outputs[10709]));
    assign layer1_outputs[7019] = layer0_outputs[6006];
    assign layer1_outputs[7020] = layer0_outputs[6760];
    assign layer1_outputs[7021] = ~((layer0_outputs[5993]) | (layer0_outputs[11071]));
    assign layer1_outputs[7022] = (layer0_outputs[11631]) & (layer0_outputs[9774]);
    assign layer1_outputs[7023] = (layer0_outputs[1240]) & ~(layer0_outputs[5486]);
    assign layer1_outputs[7024] = ~(layer0_outputs[2205]);
    assign layer1_outputs[7025] = ~(layer0_outputs[7343]);
    assign layer1_outputs[7026] = ~((layer0_outputs[11169]) & (layer0_outputs[11594]));
    assign layer1_outputs[7027] = (layer0_outputs[4213]) & ~(layer0_outputs[2689]);
    assign layer1_outputs[7028] = (layer0_outputs[498]) | (layer0_outputs[9257]);
    assign layer1_outputs[7029] = (layer0_outputs[10588]) & ~(layer0_outputs[4603]);
    assign layer1_outputs[7030] = (layer0_outputs[11425]) & (layer0_outputs[1256]);
    assign layer1_outputs[7031] = ~(layer0_outputs[12274]);
    assign layer1_outputs[7032] = ~(layer0_outputs[2635]);
    assign layer1_outputs[7033] = layer0_outputs[5587];
    assign layer1_outputs[7034] = ~(layer0_outputs[6641]);
    assign layer1_outputs[7035] = 1'b0;
    assign layer1_outputs[7036] = ~(layer0_outputs[2261]) | (layer0_outputs[1286]);
    assign layer1_outputs[7037] = layer0_outputs[12480];
    assign layer1_outputs[7038] = (layer0_outputs[7924]) & ~(layer0_outputs[1645]);
    assign layer1_outputs[7039] = ~(layer0_outputs[2749]) | (layer0_outputs[10644]);
    assign layer1_outputs[7040] = (layer0_outputs[7252]) & ~(layer0_outputs[10125]);
    assign layer1_outputs[7041] = ~(layer0_outputs[11077]);
    assign layer1_outputs[7042] = (layer0_outputs[9355]) & ~(layer0_outputs[787]);
    assign layer1_outputs[7043] = (layer0_outputs[12289]) & ~(layer0_outputs[3788]);
    assign layer1_outputs[7044] = layer0_outputs[3117];
    assign layer1_outputs[7045] = layer0_outputs[4064];
    assign layer1_outputs[7046] = layer0_outputs[11845];
    assign layer1_outputs[7047] = layer0_outputs[3074];
    assign layer1_outputs[7048] = layer0_outputs[1790];
    assign layer1_outputs[7049] = (layer0_outputs[6379]) & ~(layer0_outputs[3849]);
    assign layer1_outputs[7050] = ~(layer0_outputs[6798]) | (layer0_outputs[911]);
    assign layer1_outputs[7051] = ~((layer0_outputs[7537]) | (layer0_outputs[8458]));
    assign layer1_outputs[7052] = ~(layer0_outputs[2235]) | (layer0_outputs[10987]);
    assign layer1_outputs[7053] = ~(layer0_outputs[3055]) | (layer0_outputs[8075]);
    assign layer1_outputs[7054] = (layer0_outputs[1003]) & (layer0_outputs[3817]);
    assign layer1_outputs[7055] = ~(layer0_outputs[2675]) | (layer0_outputs[10375]);
    assign layer1_outputs[7056] = 1'b1;
    assign layer1_outputs[7057] = (layer0_outputs[6112]) | (layer0_outputs[978]);
    assign layer1_outputs[7058] = ~(layer0_outputs[4485]);
    assign layer1_outputs[7059] = layer0_outputs[8983];
    assign layer1_outputs[7060] = (layer0_outputs[7949]) | (layer0_outputs[10564]);
    assign layer1_outputs[7061] = ~(layer0_outputs[1803]);
    assign layer1_outputs[7062] = ~(layer0_outputs[8329]) | (layer0_outputs[10852]);
    assign layer1_outputs[7063] = layer0_outputs[11026];
    assign layer1_outputs[7064] = ~((layer0_outputs[3321]) ^ (layer0_outputs[1372]));
    assign layer1_outputs[7065] = ~(layer0_outputs[1631]);
    assign layer1_outputs[7066] = ~(layer0_outputs[6553]);
    assign layer1_outputs[7067] = (layer0_outputs[3233]) & (layer0_outputs[1935]);
    assign layer1_outputs[7068] = ~(layer0_outputs[7089]);
    assign layer1_outputs[7069] = ~(layer0_outputs[4753]);
    assign layer1_outputs[7070] = (layer0_outputs[11235]) & (layer0_outputs[5385]);
    assign layer1_outputs[7071] = (layer0_outputs[10578]) & ~(layer0_outputs[3296]);
    assign layer1_outputs[7072] = ~(layer0_outputs[748]);
    assign layer1_outputs[7073] = ~((layer0_outputs[8072]) ^ (layer0_outputs[4607]));
    assign layer1_outputs[7074] = ~(layer0_outputs[7867]) | (layer0_outputs[4833]);
    assign layer1_outputs[7075] = layer0_outputs[4504];
    assign layer1_outputs[7076] = (layer0_outputs[1158]) & ~(layer0_outputs[2145]);
    assign layer1_outputs[7077] = layer0_outputs[6582];
    assign layer1_outputs[7078] = ~((layer0_outputs[6375]) ^ (layer0_outputs[930]));
    assign layer1_outputs[7079] = ~((layer0_outputs[4959]) ^ (layer0_outputs[6836]));
    assign layer1_outputs[7080] = layer0_outputs[2193];
    assign layer1_outputs[7081] = ~(layer0_outputs[8936]) | (layer0_outputs[12697]);
    assign layer1_outputs[7082] = (layer0_outputs[6948]) & (layer0_outputs[8654]);
    assign layer1_outputs[7083] = ~(layer0_outputs[5528]) | (layer0_outputs[9120]);
    assign layer1_outputs[7084] = layer0_outputs[8472];
    assign layer1_outputs[7085] = (layer0_outputs[6873]) & ~(layer0_outputs[11954]);
    assign layer1_outputs[7086] = layer0_outputs[6061];
    assign layer1_outputs[7087] = ~(layer0_outputs[7887]);
    assign layer1_outputs[7088] = 1'b0;
    assign layer1_outputs[7089] = ~(layer0_outputs[3109]);
    assign layer1_outputs[7090] = (layer0_outputs[8579]) & ~(layer0_outputs[8864]);
    assign layer1_outputs[7091] = ~((layer0_outputs[5801]) & (layer0_outputs[7735]));
    assign layer1_outputs[7092] = (layer0_outputs[2270]) & ~(layer0_outputs[9085]);
    assign layer1_outputs[7093] = ~(layer0_outputs[9175]);
    assign layer1_outputs[7094] = ~((layer0_outputs[1874]) ^ (layer0_outputs[107]));
    assign layer1_outputs[7095] = ~(layer0_outputs[5125]) | (layer0_outputs[7115]);
    assign layer1_outputs[7096] = layer0_outputs[9538];
    assign layer1_outputs[7097] = ~((layer0_outputs[1043]) & (layer0_outputs[10880]));
    assign layer1_outputs[7098] = ~((layer0_outputs[10727]) ^ (layer0_outputs[1729]));
    assign layer1_outputs[7099] = ~(layer0_outputs[10842]);
    assign layer1_outputs[7100] = ~(layer0_outputs[9751]);
    assign layer1_outputs[7101] = (layer0_outputs[5375]) & ~(layer0_outputs[3406]);
    assign layer1_outputs[7102] = ~((layer0_outputs[7434]) ^ (layer0_outputs[507]));
    assign layer1_outputs[7103] = ~((layer0_outputs[12651]) ^ (layer0_outputs[7239]));
    assign layer1_outputs[7104] = 1'b0;
    assign layer1_outputs[7105] = (layer0_outputs[3486]) ^ (layer0_outputs[10863]);
    assign layer1_outputs[7106] = (layer0_outputs[8830]) | (layer0_outputs[3401]);
    assign layer1_outputs[7107] = layer0_outputs[12357];
    assign layer1_outputs[7108] = 1'b1;
    assign layer1_outputs[7109] = layer0_outputs[8068];
    assign layer1_outputs[7110] = ~(layer0_outputs[224]);
    assign layer1_outputs[7111] = ~(layer0_outputs[1500]) | (layer0_outputs[8455]);
    assign layer1_outputs[7112] = (layer0_outputs[5222]) & ~(layer0_outputs[10087]);
    assign layer1_outputs[7113] = layer0_outputs[6258];
    assign layer1_outputs[7114] = ~(layer0_outputs[5360]);
    assign layer1_outputs[7115] = ~((layer0_outputs[8960]) | (layer0_outputs[11679]));
    assign layer1_outputs[7116] = (layer0_outputs[5180]) & ~(layer0_outputs[4769]);
    assign layer1_outputs[7117] = ~(layer0_outputs[5111]);
    assign layer1_outputs[7118] = (layer0_outputs[5666]) & (layer0_outputs[12209]);
    assign layer1_outputs[7119] = layer0_outputs[10302];
    assign layer1_outputs[7120] = (layer0_outputs[3030]) ^ (layer0_outputs[3326]);
    assign layer1_outputs[7121] = ~(layer0_outputs[12208]);
    assign layer1_outputs[7122] = ~(layer0_outputs[6719]);
    assign layer1_outputs[7123] = ~(layer0_outputs[1402]);
    assign layer1_outputs[7124] = layer0_outputs[5281];
    assign layer1_outputs[7125] = ~(layer0_outputs[4147]);
    assign layer1_outputs[7126] = ~(layer0_outputs[11272]) | (layer0_outputs[4010]);
    assign layer1_outputs[7127] = layer0_outputs[1839];
    assign layer1_outputs[7128] = ~(layer0_outputs[1899]);
    assign layer1_outputs[7129] = layer0_outputs[27];
    assign layer1_outputs[7130] = layer0_outputs[2431];
    assign layer1_outputs[7131] = ~(layer0_outputs[11381]);
    assign layer1_outputs[7132] = ~(layer0_outputs[7984]) | (layer0_outputs[1654]);
    assign layer1_outputs[7133] = (layer0_outputs[812]) & (layer0_outputs[9030]);
    assign layer1_outputs[7134] = (layer0_outputs[11536]) & ~(layer0_outputs[6987]);
    assign layer1_outputs[7135] = ~(layer0_outputs[5090]) | (layer0_outputs[8242]);
    assign layer1_outputs[7136] = (layer0_outputs[6138]) ^ (layer0_outputs[6236]);
    assign layer1_outputs[7137] = ~(layer0_outputs[2685]) | (layer0_outputs[4089]);
    assign layer1_outputs[7138] = (layer0_outputs[9676]) & ~(layer0_outputs[1660]);
    assign layer1_outputs[7139] = layer0_outputs[12573];
    assign layer1_outputs[7140] = ~((layer0_outputs[3158]) ^ (layer0_outputs[12246]));
    assign layer1_outputs[7141] = ~(layer0_outputs[6999]);
    assign layer1_outputs[7142] = (layer0_outputs[11707]) & ~(layer0_outputs[3957]);
    assign layer1_outputs[7143] = layer0_outputs[5955];
    assign layer1_outputs[7144] = layer0_outputs[2162];
    assign layer1_outputs[7145] = layer0_outputs[4793];
    assign layer1_outputs[7146] = ~((layer0_outputs[9112]) & (layer0_outputs[12613]));
    assign layer1_outputs[7147] = ~(layer0_outputs[8629]);
    assign layer1_outputs[7148] = (layer0_outputs[11415]) ^ (layer0_outputs[9261]);
    assign layer1_outputs[7149] = (layer0_outputs[10088]) ^ (layer0_outputs[12374]);
    assign layer1_outputs[7150] = ~((layer0_outputs[7919]) | (layer0_outputs[6758]));
    assign layer1_outputs[7151] = ~(layer0_outputs[1396]) | (layer0_outputs[3844]);
    assign layer1_outputs[7152] = layer0_outputs[3374];
    assign layer1_outputs[7153] = ~((layer0_outputs[282]) & (layer0_outputs[12630]));
    assign layer1_outputs[7154] = ~(layer0_outputs[1083]) | (layer0_outputs[1994]);
    assign layer1_outputs[7155] = layer0_outputs[10183];
    assign layer1_outputs[7156] = ~(layer0_outputs[2987]) | (layer0_outputs[10644]);
    assign layer1_outputs[7157] = (layer0_outputs[1722]) & (layer0_outputs[7054]);
    assign layer1_outputs[7158] = ~((layer0_outputs[1641]) | (layer0_outputs[4523]));
    assign layer1_outputs[7159] = ~(layer0_outputs[2708]);
    assign layer1_outputs[7160] = ~(layer0_outputs[833]);
    assign layer1_outputs[7161] = layer0_outputs[6597];
    assign layer1_outputs[7162] = ~(layer0_outputs[12527]) | (layer0_outputs[12166]);
    assign layer1_outputs[7163] = (layer0_outputs[8705]) & ~(layer0_outputs[8541]);
    assign layer1_outputs[7164] = (layer0_outputs[9364]) & ~(layer0_outputs[5127]);
    assign layer1_outputs[7165] = ~(layer0_outputs[7623]) | (layer0_outputs[8164]);
    assign layer1_outputs[7166] = layer0_outputs[9357];
    assign layer1_outputs[7167] = ~(layer0_outputs[12680]);
    assign layer1_outputs[7168] = ~(layer0_outputs[3781]);
    assign layer1_outputs[7169] = (layer0_outputs[11496]) | (layer0_outputs[9622]);
    assign layer1_outputs[7170] = (layer0_outputs[7732]) & ~(layer0_outputs[6875]);
    assign layer1_outputs[7171] = ~(layer0_outputs[11752]);
    assign layer1_outputs[7172] = ~(layer0_outputs[1405]);
    assign layer1_outputs[7173] = (layer0_outputs[9636]) ^ (layer0_outputs[9096]);
    assign layer1_outputs[7174] = layer0_outputs[7622];
    assign layer1_outputs[7175] = (layer0_outputs[7519]) ^ (layer0_outputs[5009]);
    assign layer1_outputs[7176] = ~((layer0_outputs[10740]) | (layer0_outputs[1736]));
    assign layer1_outputs[7177] = (layer0_outputs[1745]) & ~(layer0_outputs[6401]);
    assign layer1_outputs[7178] = 1'b0;
    assign layer1_outputs[7179] = ~((layer0_outputs[8608]) ^ (layer0_outputs[11936]));
    assign layer1_outputs[7180] = (layer0_outputs[2324]) & (layer0_outputs[2547]);
    assign layer1_outputs[7181] = ~(layer0_outputs[6079]);
    assign layer1_outputs[7182] = ~(layer0_outputs[9872]) | (layer0_outputs[4110]);
    assign layer1_outputs[7183] = layer0_outputs[7730];
    assign layer1_outputs[7184] = ~(layer0_outputs[7509]);
    assign layer1_outputs[7185] = 1'b0;
    assign layer1_outputs[7186] = ~(layer0_outputs[11826]);
    assign layer1_outputs[7187] = (layer0_outputs[3305]) ^ (layer0_outputs[8756]);
    assign layer1_outputs[7188] = ~(layer0_outputs[4478]);
    assign layer1_outputs[7189] = (layer0_outputs[7743]) | (layer0_outputs[3346]);
    assign layer1_outputs[7190] = (layer0_outputs[11817]) | (layer0_outputs[7529]);
    assign layer1_outputs[7191] = layer0_outputs[11115];
    assign layer1_outputs[7192] = (layer0_outputs[2808]) & ~(layer0_outputs[12605]);
    assign layer1_outputs[7193] = ~((layer0_outputs[9944]) | (layer0_outputs[11935]));
    assign layer1_outputs[7194] = ~(layer0_outputs[10286]) | (layer0_outputs[163]);
    assign layer1_outputs[7195] = ~((layer0_outputs[11400]) | (layer0_outputs[12266]));
    assign layer1_outputs[7196] = ~(layer0_outputs[10486]) | (layer0_outputs[5634]);
    assign layer1_outputs[7197] = ~(layer0_outputs[1111]);
    assign layer1_outputs[7198] = layer0_outputs[1542];
    assign layer1_outputs[7199] = layer0_outputs[3577];
    assign layer1_outputs[7200] = (layer0_outputs[2909]) | (layer0_outputs[4087]);
    assign layer1_outputs[7201] = layer0_outputs[11832];
    assign layer1_outputs[7202] = (layer0_outputs[12799]) & ~(layer0_outputs[7299]);
    assign layer1_outputs[7203] = layer0_outputs[4204];
    assign layer1_outputs[7204] = (layer0_outputs[3833]) & ~(layer0_outputs[3919]);
    assign layer1_outputs[7205] = layer0_outputs[8222];
    assign layer1_outputs[7206] = (layer0_outputs[3865]) & ~(layer0_outputs[1144]);
    assign layer1_outputs[7207] = ~((layer0_outputs[8228]) & (layer0_outputs[11455]));
    assign layer1_outputs[7208] = layer0_outputs[1166];
    assign layer1_outputs[7209] = (layer0_outputs[12112]) | (layer0_outputs[12221]);
    assign layer1_outputs[7210] = ~((layer0_outputs[4902]) | (layer0_outputs[7094]));
    assign layer1_outputs[7211] = (layer0_outputs[9567]) & ~(layer0_outputs[10394]);
    assign layer1_outputs[7212] = ~((layer0_outputs[8583]) | (layer0_outputs[10674]));
    assign layer1_outputs[7213] = (layer0_outputs[3442]) | (layer0_outputs[11118]);
    assign layer1_outputs[7214] = ~((layer0_outputs[10681]) & (layer0_outputs[4859]));
    assign layer1_outputs[7215] = 1'b1;
    assign layer1_outputs[7216] = ~((layer0_outputs[12643]) & (layer0_outputs[7771]));
    assign layer1_outputs[7217] = ~(layer0_outputs[11886]);
    assign layer1_outputs[7218] = (layer0_outputs[203]) & ~(layer0_outputs[12438]);
    assign layer1_outputs[7219] = layer0_outputs[6152];
    assign layer1_outputs[7220] = ~((layer0_outputs[1401]) | (layer0_outputs[2761]));
    assign layer1_outputs[7221] = (layer0_outputs[2832]) | (layer0_outputs[4592]);
    assign layer1_outputs[7222] = layer0_outputs[12102];
    assign layer1_outputs[7223] = layer0_outputs[587];
    assign layer1_outputs[7224] = ~(layer0_outputs[5273]);
    assign layer1_outputs[7225] = layer0_outputs[4573];
    assign layer1_outputs[7226] = layer0_outputs[5308];
    assign layer1_outputs[7227] = ~(layer0_outputs[8278]) | (layer0_outputs[5045]);
    assign layer1_outputs[7228] = (layer0_outputs[8703]) & ~(layer0_outputs[4853]);
    assign layer1_outputs[7229] = ~((layer0_outputs[3910]) | (layer0_outputs[3502]));
    assign layer1_outputs[7230] = ~(layer0_outputs[1100]);
    assign layer1_outputs[7231] = ~(layer0_outputs[1777]);
    assign layer1_outputs[7232] = (layer0_outputs[5214]) & (layer0_outputs[3938]);
    assign layer1_outputs[7233] = (layer0_outputs[10929]) | (layer0_outputs[10449]);
    assign layer1_outputs[7234] = ~(layer0_outputs[12683]);
    assign layer1_outputs[7235] = layer0_outputs[4431];
    assign layer1_outputs[7236] = ~(layer0_outputs[3400]) | (layer0_outputs[8319]);
    assign layer1_outputs[7237] = layer0_outputs[12742];
    assign layer1_outputs[7238] = ~((layer0_outputs[5833]) ^ (layer0_outputs[12094]));
    assign layer1_outputs[7239] = (layer0_outputs[9327]) | (layer0_outputs[4481]);
    assign layer1_outputs[7240] = ~(layer0_outputs[2162]) | (layer0_outputs[8572]);
    assign layer1_outputs[7241] = (layer0_outputs[7956]) & ~(layer0_outputs[5562]);
    assign layer1_outputs[7242] = (layer0_outputs[2512]) ^ (layer0_outputs[4489]);
    assign layer1_outputs[7243] = layer0_outputs[4952];
    assign layer1_outputs[7244] = layer0_outputs[11077];
    assign layer1_outputs[7245] = ~((layer0_outputs[9607]) | (layer0_outputs[8989]));
    assign layer1_outputs[7246] = ~(layer0_outputs[887]);
    assign layer1_outputs[7247] = layer0_outputs[5528];
    assign layer1_outputs[7248] = 1'b0;
    assign layer1_outputs[7249] = ~(layer0_outputs[11201]) | (layer0_outputs[4818]);
    assign layer1_outputs[7250] = (layer0_outputs[11864]) & (layer0_outputs[10135]);
    assign layer1_outputs[7251] = layer0_outputs[6301];
    assign layer1_outputs[7252] = ~(layer0_outputs[9614]);
    assign layer1_outputs[7253] = (layer0_outputs[10438]) ^ (layer0_outputs[7404]);
    assign layer1_outputs[7254] = ~((layer0_outputs[9291]) ^ (layer0_outputs[5518]));
    assign layer1_outputs[7255] = layer0_outputs[3822];
    assign layer1_outputs[7256] = layer0_outputs[8856];
    assign layer1_outputs[7257] = layer0_outputs[9802];
    assign layer1_outputs[7258] = (layer0_outputs[10985]) & ~(layer0_outputs[476]);
    assign layer1_outputs[7259] = (layer0_outputs[9100]) & ~(layer0_outputs[9220]);
    assign layer1_outputs[7260] = ~((layer0_outputs[1811]) & (layer0_outputs[12204]));
    assign layer1_outputs[7261] = layer0_outputs[2586];
    assign layer1_outputs[7262] = ~(layer0_outputs[8820]) | (layer0_outputs[2154]);
    assign layer1_outputs[7263] = ~(layer0_outputs[206]);
    assign layer1_outputs[7264] = (layer0_outputs[5211]) ^ (layer0_outputs[433]);
    assign layer1_outputs[7265] = ~(layer0_outputs[4527]);
    assign layer1_outputs[7266] = ~((layer0_outputs[6800]) & (layer0_outputs[849]));
    assign layer1_outputs[7267] = ~(layer0_outputs[5215]);
    assign layer1_outputs[7268] = ~((layer0_outputs[1274]) ^ (layer0_outputs[3353]));
    assign layer1_outputs[7269] = ~((layer0_outputs[5378]) ^ (layer0_outputs[7226]));
    assign layer1_outputs[7270] = layer0_outputs[10701];
    assign layer1_outputs[7271] = layer0_outputs[8404];
    assign layer1_outputs[7272] = (layer0_outputs[9924]) | (layer0_outputs[11588]);
    assign layer1_outputs[7273] = ~(layer0_outputs[965]) | (layer0_outputs[3455]);
    assign layer1_outputs[7274] = (layer0_outputs[11197]) & ~(layer0_outputs[11037]);
    assign layer1_outputs[7275] = 1'b1;
    assign layer1_outputs[7276] = ~(layer0_outputs[1514]);
    assign layer1_outputs[7277] = layer0_outputs[1526];
    assign layer1_outputs[7278] = (layer0_outputs[7349]) ^ (layer0_outputs[799]);
    assign layer1_outputs[7279] = (layer0_outputs[4569]) & ~(layer0_outputs[4796]);
    assign layer1_outputs[7280] = ~((layer0_outputs[1244]) ^ (layer0_outputs[10782]));
    assign layer1_outputs[7281] = (layer0_outputs[7008]) & ~(layer0_outputs[5864]);
    assign layer1_outputs[7282] = ~(layer0_outputs[11311]);
    assign layer1_outputs[7283] = ~(layer0_outputs[891]) | (layer0_outputs[5735]);
    assign layer1_outputs[7284] = (layer0_outputs[9675]) & ~(layer0_outputs[12455]);
    assign layer1_outputs[7285] = (layer0_outputs[6896]) & ~(layer0_outputs[6775]);
    assign layer1_outputs[7286] = ~((layer0_outputs[2952]) | (layer0_outputs[1576]));
    assign layer1_outputs[7287] = 1'b0;
    assign layer1_outputs[7288] = (layer0_outputs[2208]) & (layer0_outputs[7973]);
    assign layer1_outputs[7289] = ~((layer0_outputs[8094]) ^ (layer0_outputs[11245]));
    assign layer1_outputs[7290] = ~(layer0_outputs[8342]) | (layer0_outputs[7697]);
    assign layer1_outputs[7291] = layer0_outputs[332];
    assign layer1_outputs[7292] = layer0_outputs[9185];
    assign layer1_outputs[7293] = ~((layer0_outputs[3422]) | (layer0_outputs[6351]));
    assign layer1_outputs[7294] = (layer0_outputs[7819]) ^ (layer0_outputs[4410]);
    assign layer1_outputs[7295] = ~((layer0_outputs[2603]) | (layer0_outputs[4060]));
    assign layer1_outputs[7296] = layer0_outputs[12056];
    assign layer1_outputs[7297] = ~(layer0_outputs[10330]);
    assign layer1_outputs[7298] = ~(layer0_outputs[10873]) | (layer0_outputs[11329]);
    assign layer1_outputs[7299] = ~(layer0_outputs[4056]);
    assign layer1_outputs[7300] = layer0_outputs[11887];
    assign layer1_outputs[7301] = (layer0_outputs[4886]) & (layer0_outputs[8007]);
    assign layer1_outputs[7302] = ~(layer0_outputs[4526]);
    assign layer1_outputs[7303] = layer0_outputs[2659];
    assign layer1_outputs[7304] = ~(layer0_outputs[10894]);
    assign layer1_outputs[7305] = ~(layer0_outputs[10590]) | (layer0_outputs[11249]);
    assign layer1_outputs[7306] = ~((layer0_outputs[5909]) | (layer0_outputs[3078]));
    assign layer1_outputs[7307] = (layer0_outputs[2349]) | (layer0_outputs[9373]);
    assign layer1_outputs[7308] = (layer0_outputs[8879]) & ~(layer0_outputs[7899]);
    assign layer1_outputs[7309] = (layer0_outputs[5546]) | (layer0_outputs[7082]);
    assign layer1_outputs[7310] = ~(layer0_outputs[4411]);
    assign layer1_outputs[7311] = (layer0_outputs[11398]) & ~(layer0_outputs[3648]);
    assign layer1_outputs[7312] = (layer0_outputs[6382]) & ~(layer0_outputs[6646]);
    assign layer1_outputs[7313] = ~(layer0_outputs[11972]);
    assign layer1_outputs[7314] = 1'b1;
    assign layer1_outputs[7315] = (layer0_outputs[6087]) | (layer0_outputs[6171]);
    assign layer1_outputs[7316] = (layer0_outputs[12055]) | (layer0_outputs[12599]);
    assign layer1_outputs[7317] = layer0_outputs[7852];
    assign layer1_outputs[7318] = ~(layer0_outputs[7528]);
    assign layer1_outputs[7319] = layer0_outputs[864];
    assign layer1_outputs[7320] = ~((layer0_outputs[10194]) | (layer0_outputs[11700]));
    assign layer1_outputs[7321] = ~(layer0_outputs[12637]);
    assign layer1_outputs[7322] = ~((layer0_outputs[11207]) & (layer0_outputs[7614]));
    assign layer1_outputs[7323] = ~(layer0_outputs[5563]);
    assign layer1_outputs[7324] = (layer0_outputs[3759]) & (layer0_outputs[6651]);
    assign layer1_outputs[7325] = ~(layer0_outputs[6498]) | (layer0_outputs[8948]);
    assign layer1_outputs[7326] = layer0_outputs[7502];
    assign layer1_outputs[7327] = ~(layer0_outputs[10635]);
    assign layer1_outputs[7328] = (layer0_outputs[12550]) & ~(layer0_outputs[12629]);
    assign layer1_outputs[7329] = ~(layer0_outputs[9891]) | (layer0_outputs[10383]);
    assign layer1_outputs[7330] = (layer0_outputs[6224]) & ~(layer0_outputs[5241]);
    assign layer1_outputs[7331] = ~(layer0_outputs[1499]);
    assign layer1_outputs[7332] = (layer0_outputs[10221]) ^ (layer0_outputs[1710]);
    assign layer1_outputs[7333] = ~(layer0_outputs[1553]) | (layer0_outputs[2379]);
    assign layer1_outputs[7334] = (layer0_outputs[3225]) & ~(layer0_outputs[5211]);
    assign layer1_outputs[7335] = layer0_outputs[2191];
    assign layer1_outputs[7336] = ~(layer0_outputs[8355]) | (layer0_outputs[5164]);
    assign layer1_outputs[7337] = (layer0_outputs[12741]) & ~(layer0_outputs[9352]);
    assign layer1_outputs[7338] = ~((layer0_outputs[7726]) ^ (layer0_outputs[11113]));
    assign layer1_outputs[7339] = (layer0_outputs[12287]) & ~(layer0_outputs[7508]);
    assign layer1_outputs[7340] = ~((layer0_outputs[3266]) | (layer0_outputs[252]));
    assign layer1_outputs[7341] = (layer0_outputs[9303]) ^ (layer0_outputs[7904]);
    assign layer1_outputs[7342] = ~(layer0_outputs[2744]) | (layer0_outputs[4276]);
    assign layer1_outputs[7343] = ~(layer0_outputs[776]) | (layer0_outputs[12653]);
    assign layer1_outputs[7344] = layer0_outputs[4417];
    assign layer1_outputs[7345] = ~(layer0_outputs[284]) | (layer0_outputs[2606]);
    assign layer1_outputs[7346] = ~((layer0_outputs[8606]) | (layer0_outputs[334]));
    assign layer1_outputs[7347] = layer0_outputs[11863];
    assign layer1_outputs[7348] = (layer0_outputs[8634]) | (layer0_outputs[5]);
    assign layer1_outputs[7349] = (layer0_outputs[12536]) | (layer0_outputs[3583]);
    assign layer1_outputs[7350] = ~(layer0_outputs[8084]) | (layer0_outputs[8387]);
    assign layer1_outputs[7351] = ~(layer0_outputs[11290]);
    assign layer1_outputs[7352] = (layer0_outputs[5146]) & (layer0_outputs[12498]);
    assign layer1_outputs[7353] = ~(layer0_outputs[2094]) | (layer0_outputs[7696]);
    assign layer1_outputs[7354] = (layer0_outputs[11856]) & ~(layer0_outputs[6781]);
    assign layer1_outputs[7355] = ~(layer0_outputs[12707]);
    assign layer1_outputs[7356] = ~((layer0_outputs[4389]) ^ (layer0_outputs[1292]));
    assign layer1_outputs[7357] = ~(layer0_outputs[633]);
    assign layer1_outputs[7358] = layer0_outputs[2293];
    assign layer1_outputs[7359] = ~(layer0_outputs[3405]);
    assign layer1_outputs[7360] = ~(layer0_outputs[2118]);
    assign layer1_outputs[7361] = (layer0_outputs[1084]) & ~(layer0_outputs[2044]);
    assign layer1_outputs[7362] = (layer0_outputs[2627]) & (layer0_outputs[2100]);
    assign layer1_outputs[7363] = (layer0_outputs[9526]) & (layer0_outputs[11915]);
    assign layer1_outputs[7364] = layer0_outputs[5171];
    assign layer1_outputs[7365] = ~(layer0_outputs[10913]);
    assign layer1_outputs[7366] = ~((layer0_outputs[10243]) | (layer0_outputs[4082]));
    assign layer1_outputs[7367] = (layer0_outputs[2492]) & (layer0_outputs[2627]);
    assign layer1_outputs[7368] = ~((layer0_outputs[11433]) ^ (layer0_outputs[3021]));
    assign layer1_outputs[7369] = layer0_outputs[6422];
    assign layer1_outputs[7370] = ~((layer0_outputs[11688]) ^ (layer0_outputs[7327]));
    assign layer1_outputs[7371] = ~(layer0_outputs[10503]);
    assign layer1_outputs[7372] = ~((layer0_outputs[12597]) & (layer0_outputs[9435]));
    assign layer1_outputs[7373] = ~(layer0_outputs[10154]) | (layer0_outputs[4288]);
    assign layer1_outputs[7374] = (layer0_outputs[119]) & (layer0_outputs[3075]);
    assign layer1_outputs[7375] = layer0_outputs[3122];
    assign layer1_outputs[7376] = ~(layer0_outputs[1873]) | (layer0_outputs[3897]);
    assign layer1_outputs[7377] = ~((layer0_outputs[10702]) ^ (layer0_outputs[7492]));
    assign layer1_outputs[7378] = ~((layer0_outputs[3501]) | (layer0_outputs[2725]));
    assign layer1_outputs[7379] = ~((layer0_outputs[1858]) & (layer0_outputs[9331]));
    assign layer1_outputs[7380] = layer0_outputs[3108];
    assign layer1_outputs[7381] = (layer0_outputs[8650]) & (layer0_outputs[6460]);
    assign layer1_outputs[7382] = layer0_outputs[9424];
    assign layer1_outputs[7383] = ~((layer0_outputs[4828]) | (layer0_outputs[8508]));
    assign layer1_outputs[7384] = layer0_outputs[12463];
    assign layer1_outputs[7385] = ~(layer0_outputs[9226]) | (layer0_outputs[7908]);
    assign layer1_outputs[7386] = layer0_outputs[6647];
    assign layer1_outputs[7387] = layer0_outputs[5742];
    assign layer1_outputs[7388] = ~((layer0_outputs[10761]) & (layer0_outputs[7665]));
    assign layer1_outputs[7389] = ~(layer0_outputs[11636]);
    assign layer1_outputs[7390] = ~((layer0_outputs[4980]) | (layer0_outputs[1952]));
    assign layer1_outputs[7391] = ~((layer0_outputs[5098]) | (layer0_outputs[2267]));
    assign layer1_outputs[7392] = ~(layer0_outputs[51]);
    assign layer1_outputs[7393] = layer0_outputs[1160];
    assign layer1_outputs[7394] = ~(layer0_outputs[1690]) | (layer0_outputs[3647]);
    assign layer1_outputs[7395] = (layer0_outputs[9144]) | (layer0_outputs[10360]);
    assign layer1_outputs[7396] = 1'b0;
    assign layer1_outputs[7397] = ~((layer0_outputs[11932]) | (layer0_outputs[3970]));
    assign layer1_outputs[7398] = layer0_outputs[1894];
    assign layer1_outputs[7399] = (layer0_outputs[7612]) & (layer0_outputs[6468]);
    assign layer1_outputs[7400] = ~(layer0_outputs[7728]);
    assign layer1_outputs[7401] = layer0_outputs[12304];
    assign layer1_outputs[7402] = ~(layer0_outputs[4156]);
    assign layer1_outputs[7403] = ~((layer0_outputs[3618]) & (layer0_outputs[9526]));
    assign layer1_outputs[7404] = (layer0_outputs[6722]) & ~(layer0_outputs[2185]);
    assign layer1_outputs[7405] = ~((layer0_outputs[5249]) & (layer0_outputs[5094]));
    assign layer1_outputs[7406] = layer0_outputs[6957];
    assign layer1_outputs[7407] = (layer0_outputs[12447]) & ~(layer0_outputs[8012]);
    assign layer1_outputs[7408] = (layer0_outputs[7995]) ^ (layer0_outputs[2104]);
    assign layer1_outputs[7409] = layer0_outputs[3875];
    assign layer1_outputs[7410] = ~(layer0_outputs[6675]);
    assign layer1_outputs[7411] = ~(layer0_outputs[10484]) | (layer0_outputs[919]);
    assign layer1_outputs[7412] = ~(layer0_outputs[5714]);
    assign layer1_outputs[7413] = ~(layer0_outputs[12232]);
    assign layer1_outputs[7414] = (layer0_outputs[8385]) ^ (layer0_outputs[5226]);
    assign layer1_outputs[7415] = ~(layer0_outputs[11121]);
    assign layer1_outputs[7416] = layer0_outputs[12672];
    assign layer1_outputs[7417] = ~(layer0_outputs[1673]) | (layer0_outputs[10551]);
    assign layer1_outputs[7418] = ~((layer0_outputs[3713]) & (layer0_outputs[10847]));
    assign layer1_outputs[7419] = ~(layer0_outputs[12200]);
    assign layer1_outputs[7420] = layer0_outputs[4710];
    assign layer1_outputs[7421] = ~((layer0_outputs[9972]) | (layer0_outputs[11183]));
    assign layer1_outputs[7422] = layer0_outputs[464];
    assign layer1_outputs[7423] = layer0_outputs[11740];
    assign layer1_outputs[7424] = (layer0_outputs[1599]) & ~(layer0_outputs[10419]);
    assign layer1_outputs[7425] = (layer0_outputs[1998]) | (layer0_outputs[6201]);
    assign layer1_outputs[7426] = ~(layer0_outputs[846]);
    assign layer1_outputs[7427] = (layer0_outputs[11457]) & ~(layer0_outputs[7188]);
    assign layer1_outputs[7428] = ~(layer0_outputs[736]) | (layer0_outputs[9996]);
    assign layer1_outputs[7429] = ~((layer0_outputs[2504]) & (layer0_outputs[8927]));
    assign layer1_outputs[7430] = (layer0_outputs[10815]) & ~(layer0_outputs[7388]);
    assign layer1_outputs[7431] = ~(layer0_outputs[12177]) | (layer0_outputs[5357]);
    assign layer1_outputs[7432] = (layer0_outputs[1250]) & ~(layer0_outputs[2280]);
    assign layer1_outputs[7433] = ~((layer0_outputs[6494]) ^ (layer0_outputs[1251]));
    assign layer1_outputs[7434] = ~(layer0_outputs[3306]) | (layer0_outputs[8677]);
    assign layer1_outputs[7435] = ~(layer0_outputs[3433]) | (layer0_outputs[1339]);
    assign layer1_outputs[7436] = (layer0_outputs[12406]) ^ (layer0_outputs[11216]);
    assign layer1_outputs[7437] = layer0_outputs[2086];
    assign layer1_outputs[7438] = layer0_outputs[7523];
    assign layer1_outputs[7439] = ~(layer0_outputs[7964]) | (layer0_outputs[12235]);
    assign layer1_outputs[7440] = (layer0_outputs[3399]) & (layer0_outputs[11703]);
    assign layer1_outputs[7441] = (layer0_outputs[8192]) | (layer0_outputs[6697]);
    assign layer1_outputs[7442] = layer0_outputs[3322];
    assign layer1_outputs[7443] = layer0_outputs[881];
    assign layer1_outputs[7444] = (layer0_outputs[1442]) & ~(layer0_outputs[4989]);
    assign layer1_outputs[7445] = ~(layer0_outputs[12666]) | (layer0_outputs[12016]);
    assign layer1_outputs[7446] = (layer0_outputs[1527]) & (layer0_outputs[9692]);
    assign layer1_outputs[7447] = ~((layer0_outputs[10803]) ^ (layer0_outputs[3435]));
    assign layer1_outputs[7448] = layer0_outputs[2487];
    assign layer1_outputs[7449] = layer0_outputs[154];
    assign layer1_outputs[7450] = layer0_outputs[2754];
    assign layer1_outputs[7451] = ~(layer0_outputs[452]);
    assign layer1_outputs[7452] = ~((layer0_outputs[6187]) ^ (layer0_outputs[2930]));
    assign layer1_outputs[7453] = ~(layer0_outputs[3477]);
    assign layer1_outputs[7454] = ~(layer0_outputs[2534]) | (layer0_outputs[9339]);
    assign layer1_outputs[7455] = 1'b1;
    assign layer1_outputs[7456] = ~(layer0_outputs[10266]) | (layer0_outputs[12028]);
    assign layer1_outputs[7457] = (layer0_outputs[1865]) ^ (layer0_outputs[12308]);
    assign layer1_outputs[7458] = (layer0_outputs[3337]) & ~(layer0_outputs[2334]);
    assign layer1_outputs[7459] = ~((layer0_outputs[6124]) & (layer0_outputs[4152]));
    assign layer1_outputs[7460] = ~(layer0_outputs[1916]) | (layer0_outputs[5877]);
    assign layer1_outputs[7461] = ~(layer0_outputs[2399]) | (layer0_outputs[2236]);
    assign layer1_outputs[7462] = (layer0_outputs[11568]) & (layer0_outputs[12397]);
    assign layer1_outputs[7463] = (layer0_outputs[9083]) ^ (layer0_outputs[5167]);
    assign layer1_outputs[7464] = layer0_outputs[9388];
    assign layer1_outputs[7465] = ~(layer0_outputs[2822]);
    assign layer1_outputs[7466] = ~(layer0_outputs[10773]) | (layer0_outputs[9906]);
    assign layer1_outputs[7467] = ~(layer0_outputs[1880]);
    assign layer1_outputs[7468] = ~(layer0_outputs[1147]);
    assign layer1_outputs[7469] = layer0_outputs[11861];
    assign layer1_outputs[7470] = ~(layer0_outputs[12544]) | (layer0_outputs[6557]);
    assign layer1_outputs[7471] = (layer0_outputs[10795]) & ~(layer0_outputs[6373]);
    assign layer1_outputs[7472] = ~((layer0_outputs[8898]) & (layer0_outputs[9140]));
    assign layer1_outputs[7473] = (layer0_outputs[4109]) & ~(layer0_outputs[1829]);
    assign layer1_outputs[7474] = ~(layer0_outputs[2649]) | (layer0_outputs[11191]);
    assign layer1_outputs[7475] = ~((layer0_outputs[10413]) ^ (layer0_outputs[2174]));
    assign layer1_outputs[7476] = (layer0_outputs[7034]) | (layer0_outputs[899]);
    assign layer1_outputs[7477] = ~(layer0_outputs[3403]);
    assign layer1_outputs[7478] = (layer0_outputs[11855]) & ~(layer0_outputs[2391]);
    assign layer1_outputs[7479] = (layer0_outputs[11927]) & (layer0_outputs[480]);
    assign layer1_outputs[7480] = 1'b0;
    assign layer1_outputs[7481] = (layer0_outputs[3550]) & (layer0_outputs[1613]);
    assign layer1_outputs[7482] = ~((layer0_outputs[7184]) & (layer0_outputs[6170]));
    assign layer1_outputs[7483] = 1'b1;
    assign layer1_outputs[7484] = (layer0_outputs[6991]) | (layer0_outputs[8324]);
    assign layer1_outputs[7485] = ~((layer0_outputs[8503]) ^ (layer0_outputs[2767]));
    assign layer1_outputs[7486] = (layer0_outputs[10546]) & (layer0_outputs[12731]);
    assign layer1_outputs[7487] = layer0_outputs[5099];
    assign layer1_outputs[7488] = (layer0_outputs[1322]) & (layer0_outputs[3398]);
    assign layer1_outputs[7489] = ~((layer0_outputs[10044]) | (layer0_outputs[108]));
    assign layer1_outputs[7490] = ~(layer0_outputs[11085]);
    assign layer1_outputs[7491] = ~(layer0_outputs[5276]) | (layer0_outputs[931]);
    assign layer1_outputs[7492] = (layer0_outputs[10318]) & ~(layer0_outputs[6031]);
    assign layer1_outputs[7493] = ~((layer0_outputs[315]) | (layer0_outputs[10735]));
    assign layer1_outputs[7494] = ~(layer0_outputs[5347]) | (layer0_outputs[3737]);
    assign layer1_outputs[7495] = ~(layer0_outputs[5013]);
    assign layer1_outputs[7496] = layer0_outputs[406];
    assign layer1_outputs[7497] = layer0_outputs[4732];
    assign layer1_outputs[7498] = ~((layer0_outputs[11790]) ^ (layer0_outputs[5113]));
    assign layer1_outputs[7499] = ~(layer0_outputs[3578]);
    assign layer1_outputs[7500] = (layer0_outputs[5010]) | (layer0_outputs[3332]);
    assign layer1_outputs[7501] = layer0_outputs[9456];
    assign layer1_outputs[7502] = ~(layer0_outputs[4114]);
    assign layer1_outputs[7503] = (layer0_outputs[6737]) | (layer0_outputs[9230]);
    assign layer1_outputs[7504] = ~(layer0_outputs[11950]);
    assign layer1_outputs[7505] = ~(layer0_outputs[6588]);
    assign layer1_outputs[7506] = ~((layer0_outputs[5517]) & (layer0_outputs[6758]));
    assign layer1_outputs[7507] = (layer0_outputs[4766]) | (layer0_outputs[5575]);
    assign layer1_outputs[7508] = (layer0_outputs[9681]) | (layer0_outputs[10451]);
    assign layer1_outputs[7509] = ~(layer0_outputs[12308]) | (layer0_outputs[4515]);
    assign layer1_outputs[7510] = (layer0_outputs[5009]) ^ (layer0_outputs[1911]);
    assign layer1_outputs[7511] = (layer0_outputs[8064]) | (layer0_outputs[11108]);
    assign layer1_outputs[7512] = 1'b1;
    assign layer1_outputs[7513] = layer0_outputs[9800];
    assign layer1_outputs[7514] = ~(layer0_outputs[12197]) | (layer0_outputs[8500]);
    assign layer1_outputs[7515] = ~(layer0_outputs[7737]);
    assign layer1_outputs[7516] = ~(layer0_outputs[776]);
    assign layer1_outputs[7517] = 1'b0;
    assign layer1_outputs[7518] = layer0_outputs[7372];
    assign layer1_outputs[7519] = ~((layer0_outputs[12683]) & (layer0_outputs[11918]));
    assign layer1_outputs[7520] = (layer0_outputs[3801]) | (layer0_outputs[11328]);
    assign layer1_outputs[7521] = ~(layer0_outputs[12303]);
    assign layer1_outputs[7522] = ~((layer0_outputs[4735]) ^ (layer0_outputs[3879]));
    assign layer1_outputs[7523] = ~(layer0_outputs[4272]);
    assign layer1_outputs[7524] = 1'b0;
    assign layer1_outputs[7525] = ~((layer0_outputs[3413]) ^ (layer0_outputs[5871]));
    assign layer1_outputs[7526] = (layer0_outputs[9554]) | (layer0_outputs[197]);
    assign layer1_outputs[7527] = layer0_outputs[12271];
    assign layer1_outputs[7528] = (layer0_outputs[12260]) & ~(layer0_outputs[11744]);
    assign layer1_outputs[7529] = ~((layer0_outputs[4138]) ^ (layer0_outputs[10833]));
    assign layer1_outputs[7530] = ~(layer0_outputs[9585]) | (layer0_outputs[192]);
    assign layer1_outputs[7531] = ~((layer0_outputs[9693]) ^ (layer0_outputs[7546]));
    assign layer1_outputs[7532] = ~(layer0_outputs[139]);
    assign layer1_outputs[7533] = (layer0_outputs[429]) & (layer0_outputs[6180]);
    assign layer1_outputs[7534] = layer0_outputs[5676];
    assign layer1_outputs[7535] = (layer0_outputs[1481]) & (layer0_outputs[2447]);
    assign layer1_outputs[7536] = layer0_outputs[662];
    assign layer1_outputs[7537] = ~((layer0_outputs[7826]) & (layer0_outputs[7991]));
    assign layer1_outputs[7538] = (layer0_outputs[5125]) | (layer0_outputs[7495]);
    assign layer1_outputs[7539] = (layer0_outputs[3579]) ^ (layer0_outputs[7594]);
    assign layer1_outputs[7540] = (layer0_outputs[9186]) ^ (layer0_outputs[3104]);
    assign layer1_outputs[7541] = (layer0_outputs[7312]) ^ (layer0_outputs[12236]);
    assign layer1_outputs[7542] = layer0_outputs[7621];
    assign layer1_outputs[7543] = ~((layer0_outputs[12499]) ^ (layer0_outputs[11728]));
    assign layer1_outputs[7544] = ~((layer0_outputs[2608]) | (layer0_outputs[3404]));
    assign layer1_outputs[7545] = (layer0_outputs[2004]) & ~(layer0_outputs[8073]);
    assign layer1_outputs[7546] = ~((layer0_outputs[8678]) ^ (layer0_outputs[8210]));
    assign layer1_outputs[7547] = layer0_outputs[2549];
    assign layer1_outputs[7548] = (layer0_outputs[5316]) | (layer0_outputs[12523]);
    assign layer1_outputs[7549] = ~(layer0_outputs[8295]);
    assign layer1_outputs[7550] = ~(layer0_outputs[7870]);
    assign layer1_outputs[7551] = ~(layer0_outputs[9910]);
    assign layer1_outputs[7552] = layer0_outputs[2885];
    assign layer1_outputs[7553] = (layer0_outputs[9302]) | (layer0_outputs[1478]);
    assign layer1_outputs[7554] = (layer0_outputs[7569]) & ~(layer0_outputs[11993]);
    assign layer1_outputs[7555] = (layer0_outputs[6759]) & ~(layer0_outputs[10373]);
    assign layer1_outputs[7556] = (layer0_outputs[4134]) & ~(layer0_outputs[6743]);
    assign layer1_outputs[7557] = ~((layer0_outputs[7414]) ^ (layer0_outputs[11091]));
    assign layer1_outputs[7558] = ~(layer0_outputs[9976]);
    assign layer1_outputs[7559] = ~(layer0_outputs[8846]);
    assign layer1_outputs[7560] = ~(layer0_outputs[655]);
    assign layer1_outputs[7561] = (layer0_outputs[11286]) | (layer0_outputs[10267]);
    assign layer1_outputs[7562] = layer0_outputs[3223];
    assign layer1_outputs[7563] = layer0_outputs[2462];
    assign layer1_outputs[7564] = ~(layer0_outputs[3264]);
    assign layer1_outputs[7565] = layer0_outputs[9909];
    assign layer1_outputs[7566] = layer0_outputs[4238];
    assign layer1_outputs[7567] = ~(layer0_outputs[8100]);
    assign layer1_outputs[7568] = ~(layer0_outputs[1368]) | (layer0_outputs[1500]);
    assign layer1_outputs[7569] = ~(layer0_outputs[8699]) | (layer0_outputs[4655]);
    assign layer1_outputs[7570] = ~(layer0_outputs[1807]);
    assign layer1_outputs[7571] = ~(layer0_outputs[6295]) | (layer0_outputs[11124]);
    assign layer1_outputs[7572] = ~(layer0_outputs[5230]);
    assign layer1_outputs[7573] = (layer0_outputs[1789]) & ~(layer0_outputs[8567]);
    assign layer1_outputs[7574] = layer0_outputs[4634];
    assign layer1_outputs[7575] = layer0_outputs[10760];
    assign layer1_outputs[7576] = layer0_outputs[6802];
    assign layer1_outputs[7577] = (layer0_outputs[2980]) ^ (layer0_outputs[9718]);
    assign layer1_outputs[7578] = (layer0_outputs[11473]) ^ (layer0_outputs[11034]);
    assign layer1_outputs[7579] = 1'b1;
    assign layer1_outputs[7580] = (layer0_outputs[11043]) ^ (layer0_outputs[6038]);
    assign layer1_outputs[7581] = ~(layer0_outputs[10361]);
    assign layer1_outputs[7582] = layer0_outputs[6073];
    assign layer1_outputs[7583] = (layer0_outputs[12151]) & ~(layer0_outputs[11331]);
    assign layer1_outputs[7584] = ~(layer0_outputs[6092]);
    assign layer1_outputs[7585] = ~(layer0_outputs[4836]);
    assign layer1_outputs[7586] = layer0_outputs[4991];
    assign layer1_outputs[7587] = ~(layer0_outputs[9989]) | (layer0_outputs[7693]);
    assign layer1_outputs[7588] = (layer0_outputs[3488]) ^ (layer0_outputs[5597]);
    assign layer1_outputs[7589] = layer0_outputs[3724];
    assign layer1_outputs[7590] = ~(layer0_outputs[913]);
    assign layer1_outputs[7591] = ~(layer0_outputs[552]);
    assign layer1_outputs[7592] = ~(layer0_outputs[12123]);
    assign layer1_outputs[7593] = (layer0_outputs[10177]) & (layer0_outputs[8515]);
    assign layer1_outputs[7594] = ~((layer0_outputs[3132]) & (layer0_outputs[1343]));
    assign layer1_outputs[7595] = layer0_outputs[8995];
    assign layer1_outputs[7596] = ~((layer0_outputs[3517]) ^ (layer0_outputs[6317]));
    assign layer1_outputs[7597] = (layer0_outputs[2885]) & ~(layer0_outputs[11526]);
    assign layer1_outputs[7598] = ~(layer0_outputs[8469]) | (layer0_outputs[11102]);
    assign layer1_outputs[7599] = (layer0_outputs[7719]) ^ (layer0_outputs[8310]);
    assign layer1_outputs[7600] = layer0_outputs[4574];
    assign layer1_outputs[7601] = layer0_outputs[2806];
    assign layer1_outputs[7602] = ~(layer0_outputs[2664]) | (layer0_outputs[5480]);
    assign layer1_outputs[7603] = layer0_outputs[317];
    assign layer1_outputs[7604] = layer0_outputs[6323];
    assign layer1_outputs[7605] = ~(layer0_outputs[11938]);
    assign layer1_outputs[7606] = layer0_outputs[6955];
    assign layer1_outputs[7607] = (layer0_outputs[8335]) & (layer0_outputs[3057]);
    assign layer1_outputs[7608] = ~(layer0_outputs[10713]) | (layer0_outputs[11341]);
    assign layer1_outputs[7609] = ~((layer0_outputs[7054]) & (layer0_outputs[3843]));
    assign layer1_outputs[7610] = ~(layer0_outputs[6743]);
    assign layer1_outputs[7611] = (layer0_outputs[3084]) | (layer0_outputs[2678]);
    assign layer1_outputs[7612] = ~((layer0_outputs[11898]) | (layer0_outputs[9940]));
    assign layer1_outputs[7613] = layer0_outputs[4085];
    assign layer1_outputs[7614] = (layer0_outputs[836]) & ~(layer0_outputs[8180]);
    assign layer1_outputs[7615] = (layer0_outputs[7130]) & (layer0_outputs[5970]);
    assign layer1_outputs[7616] = (layer0_outputs[9210]) | (layer0_outputs[10445]);
    assign layer1_outputs[7617] = ~(layer0_outputs[7594]);
    assign layer1_outputs[7618] = ~((layer0_outputs[6067]) & (layer0_outputs[673]));
    assign layer1_outputs[7619] = layer0_outputs[2825];
    assign layer1_outputs[7620] = ~(layer0_outputs[4633]);
    assign layer1_outputs[7621] = (layer0_outputs[12107]) & (layer0_outputs[7763]);
    assign layer1_outputs[7622] = ~((layer0_outputs[4363]) ^ (layer0_outputs[6108]));
    assign layer1_outputs[7623] = layer0_outputs[9471];
    assign layer1_outputs[7624] = (layer0_outputs[4038]) ^ (layer0_outputs[10838]);
    assign layer1_outputs[7625] = (layer0_outputs[10622]) & (layer0_outputs[10781]);
    assign layer1_outputs[7626] = ~((layer0_outputs[8947]) | (layer0_outputs[7479]));
    assign layer1_outputs[7627] = (layer0_outputs[1828]) & ~(layer0_outputs[7393]);
    assign layer1_outputs[7628] = layer0_outputs[11177];
    assign layer1_outputs[7629] = ~((layer0_outputs[3419]) & (layer0_outputs[4630]));
    assign layer1_outputs[7630] = ~(layer0_outputs[3070]);
    assign layer1_outputs[7631] = ~(layer0_outputs[3654]) | (layer0_outputs[3071]);
    assign layer1_outputs[7632] = (layer0_outputs[4187]) & ~(layer0_outputs[4004]);
    assign layer1_outputs[7633] = ~((layer0_outputs[11671]) & (layer0_outputs[4562]));
    assign layer1_outputs[7634] = ~(layer0_outputs[10048]);
    assign layer1_outputs[7635] = ~((layer0_outputs[2806]) ^ (layer0_outputs[2328]));
    assign layer1_outputs[7636] = (layer0_outputs[8205]) & ~(layer0_outputs[3277]);
    assign layer1_outputs[7637] = (layer0_outputs[188]) | (layer0_outputs[4551]);
    assign layer1_outputs[7638] = ~(layer0_outputs[307]) | (layer0_outputs[1763]);
    assign layer1_outputs[7639] = ~(layer0_outputs[5620]);
    assign layer1_outputs[7640] = ~((layer0_outputs[11775]) & (layer0_outputs[12146]));
    assign layer1_outputs[7641] = ~(layer0_outputs[7780]) | (layer0_outputs[7422]);
    assign layer1_outputs[7642] = ~((layer0_outputs[5476]) | (layer0_outputs[8884]));
    assign layer1_outputs[7643] = ~(layer0_outputs[7724]);
    assign layer1_outputs[7644] = (layer0_outputs[3685]) | (layer0_outputs[12688]);
    assign layer1_outputs[7645] = (layer0_outputs[8194]) ^ (layer0_outputs[1267]);
    assign layer1_outputs[7646] = layer0_outputs[6639];
    assign layer1_outputs[7647] = (layer0_outputs[459]) ^ (layer0_outputs[1227]);
    assign layer1_outputs[7648] = (layer0_outputs[9346]) & ~(layer0_outputs[711]);
    assign layer1_outputs[7649] = (layer0_outputs[7607]) & ~(layer0_outputs[10332]);
    assign layer1_outputs[7650] = layer0_outputs[7820];
    assign layer1_outputs[7651] = ~(layer0_outputs[914]);
    assign layer1_outputs[7652] = ~((layer0_outputs[10962]) ^ (layer0_outputs[11101]));
    assign layer1_outputs[7653] = ~(layer0_outputs[7397]);
    assign layer1_outputs[7654] = ~((layer0_outputs[12129]) ^ (layer0_outputs[7103]));
    assign layer1_outputs[7655] = (layer0_outputs[9846]) ^ (layer0_outputs[4831]);
    assign layer1_outputs[7656] = ~((layer0_outputs[4072]) & (layer0_outputs[2960]));
    assign layer1_outputs[7657] = ~(layer0_outputs[11982]);
    assign layer1_outputs[7658] = 1'b1;
    assign layer1_outputs[7659] = layer0_outputs[10297];
    assign layer1_outputs[7660] = ~(layer0_outputs[4910]);
    assign layer1_outputs[7661] = (layer0_outputs[118]) ^ (layer0_outputs[604]);
    assign layer1_outputs[7662] = ~(layer0_outputs[310]) | (layer0_outputs[8743]);
    assign layer1_outputs[7663] = ~(layer0_outputs[5275]);
    assign layer1_outputs[7664] = layer0_outputs[9185];
    assign layer1_outputs[7665] = 1'b0;
    assign layer1_outputs[7666] = (layer0_outputs[9169]) & ~(layer0_outputs[3291]);
    assign layer1_outputs[7667] = layer0_outputs[7599];
    assign layer1_outputs[7668] = ~(layer0_outputs[785]);
    assign layer1_outputs[7669] = (layer0_outputs[8332]) & ~(layer0_outputs[9308]);
    assign layer1_outputs[7670] = (layer0_outputs[4716]) & (layer0_outputs[9785]);
    assign layer1_outputs[7671] = (layer0_outputs[10151]) & ~(layer0_outputs[1168]);
    assign layer1_outputs[7672] = (layer0_outputs[12392]) ^ (layer0_outputs[6012]);
    assign layer1_outputs[7673] = ~((layer0_outputs[11647]) ^ (layer0_outputs[1423]));
    assign layer1_outputs[7674] = ~(layer0_outputs[5818]) | (layer0_outputs[9442]);
    assign layer1_outputs[7675] = ~(layer0_outputs[2925]) | (layer0_outputs[5758]);
    assign layer1_outputs[7676] = layer0_outputs[2102];
    assign layer1_outputs[7677] = (layer0_outputs[9398]) & ~(layer0_outputs[4415]);
    assign layer1_outputs[7678] = ~(layer0_outputs[27]);
    assign layer1_outputs[7679] = layer0_outputs[3831];
    assign layer1_outputs[7680] = (layer0_outputs[9011]) & ~(layer0_outputs[2734]);
    assign layer1_outputs[7681] = ~(layer0_outputs[9694]) | (layer0_outputs[5912]);
    assign layer1_outputs[7682] = ~(layer0_outputs[7782]) | (layer0_outputs[7128]);
    assign layer1_outputs[7683] = ~((layer0_outputs[12133]) | (layer0_outputs[739]));
    assign layer1_outputs[7684] = (layer0_outputs[6120]) & ~(layer0_outputs[9418]);
    assign layer1_outputs[7685] = ~(layer0_outputs[803]) | (layer0_outputs[5600]);
    assign layer1_outputs[7686] = ~((layer0_outputs[9182]) & (layer0_outputs[11695]));
    assign layer1_outputs[7687] = (layer0_outputs[618]) & ~(layer0_outputs[9297]);
    assign layer1_outputs[7688] = (layer0_outputs[11468]) & ~(layer0_outputs[4247]);
    assign layer1_outputs[7689] = ~(layer0_outputs[8600]);
    assign layer1_outputs[7690] = ~((layer0_outputs[917]) & (layer0_outputs[7644]));
    assign layer1_outputs[7691] = ~(layer0_outputs[6735]) | (layer0_outputs[1650]);
    assign layer1_outputs[7692] = (layer0_outputs[5059]) | (layer0_outputs[10799]);
    assign layer1_outputs[7693] = (layer0_outputs[11934]) | (layer0_outputs[6568]);
    assign layer1_outputs[7694] = ~(layer0_outputs[9818]);
    assign layer1_outputs[7695] = ~(layer0_outputs[11630]);
    assign layer1_outputs[7696] = ~(layer0_outputs[8593]);
    assign layer1_outputs[7697] = ~(layer0_outputs[420]);
    assign layer1_outputs[7698] = ~((layer0_outputs[4597]) | (layer0_outputs[5408]));
    assign layer1_outputs[7699] = (layer0_outputs[5554]) | (layer0_outputs[762]);
    assign layer1_outputs[7700] = ~(layer0_outputs[5571]);
    assign layer1_outputs[7701] = ~((layer0_outputs[369]) ^ (layer0_outputs[4880]));
    assign layer1_outputs[7702] = ~(layer0_outputs[10327]);
    assign layer1_outputs[7703] = (layer0_outputs[1930]) & ~(layer0_outputs[5015]);
    assign layer1_outputs[7704] = ~((layer0_outputs[5960]) | (layer0_outputs[3626]));
    assign layer1_outputs[7705] = ~((layer0_outputs[2887]) & (layer0_outputs[6039]));
    assign layer1_outputs[7706] = (layer0_outputs[9466]) & ~(layer0_outputs[3385]);
    assign layer1_outputs[7707] = ~(layer0_outputs[11888]) | (layer0_outputs[10347]);
    assign layer1_outputs[7708] = 1'b1;
    assign layer1_outputs[7709] = (layer0_outputs[2708]) & (layer0_outputs[2078]);
    assign layer1_outputs[7710] = layer0_outputs[2418];
    assign layer1_outputs[7711] = layer0_outputs[437];
    assign layer1_outputs[7712] = ~(layer0_outputs[2921]);
    assign layer1_outputs[7713] = ~(layer0_outputs[2706]);
    assign layer1_outputs[7714] = (layer0_outputs[2388]) | (layer0_outputs[10984]);
    assign layer1_outputs[7715] = ~(layer0_outputs[10166]) | (layer0_outputs[6186]);
    assign layer1_outputs[7716] = (layer0_outputs[11116]) & ~(layer0_outputs[5010]);
    assign layer1_outputs[7717] = layer0_outputs[10240];
    assign layer1_outputs[7718] = layer0_outputs[8687];
    assign layer1_outputs[7719] = ~(layer0_outputs[1883]);
    assign layer1_outputs[7720] = ~((layer0_outputs[12789]) ^ (layer0_outputs[10311]));
    assign layer1_outputs[7721] = ~((layer0_outputs[8633]) | (layer0_outputs[8703]));
    assign layer1_outputs[7722] = ~(layer0_outputs[3865]) | (layer0_outputs[9642]);
    assign layer1_outputs[7723] = ~(layer0_outputs[9470]) | (layer0_outputs[8593]);
    assign layer1_outputs[7724] = 1'b0;
    assign layer1_outputs[7725] = ~(layer0_outputs[7741]) | (layer0_outputs[6131]);
    assign layer1_outputs[7726] = (layer0_outputs[950]) & (layer0_outputs[12092]);
    assign layer1_outputs[7727] = ~((layer0_outputs[1031]) | (layer0_outputs[3250]));
    assign layer1_outputs[7728] = ~(layer0_outputs[4092]);
    assign layer1_outputs[7729] = (layer0_outputs[5117]) & ~(layer0_outputs[5529]);
    assign layer1_outputs[7730] = ~(layer0_outputs[5689]) | (layer0_outputs[8194]);
    assign layer1_outputs[7731] = ~((layer0_outputs[3354]) ^ (layer0_outputs[2875]));
    assign layer1_outputs[7732] = ~(layer0_outputs[9537]) | (layer0_outputs[5080]);
    assign layer1_outputs[7733] = layer0_outputs[10430];
    assign layer1_outputs[7734] = ~(layer0_outputs[11231]);
    assign layer1_outputs[7735] = layer0_outputs[4122];
    assign layer1_outputs[7736] = ~(layer0_outputs[4488]);
    assign layer1_outputs[7737] = (layer0_outputs[3210]) & ~(layer0_outputs[4688]);
    assign layer1_outputs[7738] = ~(layer0_outputs[8801]) | (layer0_outputs[350]);
    assign layer1_outputs[7739] = ~(layer0_outputs[6395]) | (layer0_outputs[6916]);
    assign layer1_outputs[7740] = layer0_outputs[4656];
    assign layer1_outputs[7741] = ~(layer0_outputs[10325]) | (layer0_outputs[546]);
    assign layer1_outputs[7742] = ~(layer0_outputs[8286]) | (layer0_outputs[3729]);
    assign layer1_outputs[7743] = ~((layer0_outputs[6995]) | (layer0_outputs[11379]));
    assign layer1_outputs[7744] = (layer0_outputs[10628]) & (layer0_outputs[2485]);
    assign layer1_outputs[7745] = ~((layer0_outputs[6167]) | (layer0_outputs[340]));
    assign layer1_outputs[7746] = (layer0_outputs[488]) & ~(layer0_outputs[6968]);
    assign layer1_outputs[7747] = 1'b1;
    assign layer1_outputs[7748] = ~(layer0_outputs[7554]);
    assign layer1_outputs[7749] = layer0_outputs[8938];
    assign layer1_outputs[7750] = ~(layer0_outputs[10114]);
    assign layer1_outputs[7751] = (layer0_outputs[8664]) & (layer0_outputs[657]);
    assign layer1_outputs[7752] = ~(layer0_outputs[2683]);
    assign layer1_outputs[7753] = ~(layer0_outputs[2545]);
    assign layer1_outputs[7754] = ~(layer0_outputs[782]);
    assign layer1_outputs[7755] = ~(layer0_outputs[4711]);
    assign layer1_outputs[7756] = ~((layer0_outputs[3864]) | (layer0_outputs[7365]));
    assign layer1_outputs[7757] = (layer0_outputs[38]) & ~(layer0_outputs[1814]);
    assign layer1_outputs[7758] = layer0_outputs[2584];
    assign layer1_outputs[7759] = ~((layer0_outputs[3540]) & (layer0_outputs[836]));
    assign layer1_outputs[7760] = layer0_outputs[840];
    assign layer1_outputs[7761] = 1'b1;
    assign layer1_outputs[7762] = (layer0_outputs[886]) & ~(layer0_outputs[12382]);
    assign layer1_outputs[7763] = (layer0_outputs[7395]) & (layer0_outputs[12705]);
    assign layer1_outputs[7764] = ~((layer0_outputs[7247]) & (layer0_outputs[2663]));
    assign layer1_outputs[7765] = ~((layer0_outputs[7539]) | (layer0_outputs[6432]));
    assign layer1_outputs[7766] = (layer0_outputs[12467]) ^ (layer0_outputs[2091]);
    assign layer1_outputs[7767] = ~(layer0_outputs[8401]) | (layer0_outputs[1533]);
    assign layer1_outputs[7768] = ~(layer0_outputs[11191]);
    assign layer1_outputs[7769] = (layer0_outputs[3131]) | (layer0_outputs[7639]);
    assign layer1_outputs[7770] = 1'b1;
    assign layer1_outputs[7771] = ~(layer0_outputs[1136]);
    assign layer1_outputs[7772] = (layer0_outputs[1145]) & ~(layer0_outputs[3133]);
    assign layer1_outputs[7773] = ~((layer0_outputs[10938]) | (layer0_outputs[499]));
    assign layer1_outputs[7774] = (layer0_outputs[7881]) | (layer0_outputs[12365]);
    assign layer1_outputs[7775] = layer0_outputs[1543];
    assign layer1_outputs[7776] = ~((layer0_outputs[358]) | (layer0_outputs[9750]));
    assign layer1_outputs[7777] = (layer0_outputs[8659]) ^ (layer0_outputs[7832]);
    assign layer1_outputs[7778] = ~(layer0_outputs[7890]);
    assign layer1_outputs[7779] = layer0_outputs[12145];
    assign layer1_outputs[7780] = ~(layer0_outputs[6611]);
    assign layer1_outputs[7781] = (layer0_outputs[5395]) & (layer0_outputs[583]);
    assign layer1_outputs[7782] = (layer0_outputs[10375]) & ~(layer0_outputs[6902]);
    assign layer1_outputs[7783] = ~(layer0_outputs[3413]) | (layer0_outputs[6204]);
    assign layer1_outputs[7784] = ~(layer0_outputs[7794]);
    assign layer1_outputs[7785] = layer0_outputs[6719];
    assign layer1_outputs[7786] = ~(layer0_outputs[10163]) | (layer0_outputs[9052]);
    assign layer1_outputs[7787] = (layer0_outputs[2933]) & (layer0_outputs[8358]);
    assign layer1_outputs[7788] = layer0_outputs[9778];
    assign layer1_outputs[7789] = (layer0_outputs[4962]) ^ (layer0_outputs[8277]);
    assign layer1_outputs[7790] = (layer0_outputs[5313]) & (layer0_outputs[5900]);
    assign layer1_outputs[7791] = ~(layer0_outputs[7835]) | (layer0_outputs[1258]);
    assign layer1_outputs[7792] = ~((layer0_outputs[9135]) ^ (layer0_outputs[11012]));
    assign layer1_outputs[7793] = (layer0_outputs[691]) & (layer0_outputs[6784]);
    assign layer1_outputs[7794] = ~(layer0_outputs[3200]);
    assign layer1_outputs[7795] = ~(layer0_outputs[6015]) | (layer0_outputs[3615]);
    assign layer1_outputs[7796] = ~(layer0_outputs[3899]);
    assign layer1_outputs[7797] = ~(layer0_outputs[9147]);
    assign layer1_outputs[7798] = layer0_outputs[12154];
    assign layer1_outputs[7799] = ~(layer0_outputs[10500]);
    assign layer1_outputs[7800] = ~(layer0_outputs[6409]);
    assign layer1_outputs[7801] = (layer0_outputs[2568]) & ~(layer0_outputs[5041]);
    assign layer1_outputs[7802] = layer0_outputs[11140];
    assign layer1_outputs[7803] = (layer0_outputs[195]) & ~(layer0_outputs[5481]);
    assign layer1_outputs[7804] = layer0_outputs[6848];
    assign layer1_outputs[7805] = (layer0_outputs[6444]) & ~(layer0_outputs[7235]);
    assign layer1_outputs[7806] = ~(layer0_outputs[9367]) | (layer0_outputs[5571]);
    assign layer1_outputs[7807] = ~(layer0_outputs[2537]);
    assign layer1_outputs[7808] = ~(layer0_outputs[10673]);
    assign layer1_outputs[7809] = ~(layer0_outputs[1568]);
    assign layer1_outputs[7810] = (layer0_outputs[84]) | (layer0_outputs[11867]);
    assign layer1_outputs[7811] = layer0_outputs[960];
    assign layer1_outputs[7812] = ~(layer0_outputs[3846]) | (layer0_outputs[10629]);
    assign layer1_outputs[7813] = layer0_outputs[8070];
    assign layer1_outputs[7814] = layer0_outputs[11040];
    assign layer1_outputs[7815] = ~(layer0_outputs[9625]);
    assign layer1_outputs[7816] = layer0_outputs[12718];
    assign layer1_outputs[7817] = ~(layer0_outputs[7630]);
    assign layer1_outputs[7818] = (layer0_outputs[12351]) & ~(layer0_outputs[1436]);
    assign layer1_outputs[7819] = ~((layer0_outputs[12735]) & (layer0_outputs[5405]));
    assign layer1_outputs[7820] = ~(layer0_outputs[5238]) | (layer0_outputs[4492]);
    assign layer1_outputs[7821] = ~(layer0_outputs[4327]) | (layer0_outputs[5400]);
    assign layer1_outputs[7822] = layer0_outputs[12118];
    assign layer1_outputs[7823] = layer0_outputs[256];
    assign layer1_outputs[7824] = layer0_outputs[11668];
    assign layer1_outputs[7825] = (layer0_outputs[7653]) & ~(layer0_outputs[8566]);
    assign layer1_outputs[7826] = (layer0_outputs[11015]) & ~(layer0_outputs[1753]);
    assign layer1_outputs[7827] = ~(layer0_outputs[6064]);
    assign layer1_outputs[7828] = ~((layer0_outputs[6693]) & (layer0_outputs[10049]));
    assign layer1_outputs[7829] = ~(layer0_outputs[7244]);
    assign layer1_outputs[7830] = (layer0_outputs[6138]) & ~(layer0_outputs[11258]);
    assign layer1_outputs[7831] = ~(layer0_outputs[3509]) | (layer0_outputs[72]);
    assign layer1_outputs[7832] = layer0_outputs[10808];
    assign layer1_outputs[7833] = ~(layer0_outputs[10449]);
    assign layer1_outputs[7834] = ~(layer0_outputs[10390]);
    assign layer1_outputs[7835] = ~(layer0_outputs[7499]);
    assign layer1_outputs[7836] = layer0_outputs[10415];
    assign layer1_outputs[7837] = (layer0_outputs[448]) ^ (layer0_outputs[8602]);
    assign layer1_outputs[7838] = ~(layer0_outputs[9170]) | (layer0_outputs[5248]);
    assign layer1_outputs[7839] = ~(layer0_outputs[6382]) | (layer0_outputs[2552]);
    assign layer1_outputs[7840] = (layer0_outputs[3147]) & (layer0_outputs[2262]);
    assign layer1_outputs[7841] = layer0_outputs[8109];
    assign layer1_outputs[7842] = ~(layer0_outputs[9613]) | (layer0_outputs[2128]);
    assign layer1_outputs[7843] = ~((layer0_outputs[7657]) ^ (layer0_outputs[11055]));
    assign layer1_outputs[7844] = ~(layer0_outputs[2439]);
    assign layer1_outputs[7845] = ~(layer0_outputs[5628]);
    assign layer1_outputs[7846] = ~((layer0_outputs[8083]) | (layer0_outputs[7758]));
    assign layer1_outputs[7847] = layer0_outputs[4754];
    assign layer1_outputs[7848] = ~(layer0_outputs[824]);
    assign layer1_outputs[7849] = layer0_outputs[7966];
    assign layer1_outputs[7850] = 1'b0;
    assign layer1_outputs[7851] = ~(layer0_outputs[2765]);
    assign layer1_outputs[7852] = ~(layer0_outputs[5102]);
    assign layer1_outputs[7853] = (layer0_outputs[3644]) & ~(layer0_outputs[1241]);
    assign layer1_outputs[7854] = ~(layer0_outputs[12108]) | (layer0_outputs[4867]);
    assign layer1_outputs[7855] = ~(layer0_outputs[12139]);
    assign layer1_outputs[7856] = ~(layer0_outputs[1157]);
    assign layer1_outputs[7857] = ~(layer0_outputs[1979]);
    assign layer1_outputs[7858] = ~(layer0_outputs[6415]);
    assign layer1_outputs[7859] = layer0_outputs[11960];
    assign layer1_outputs[7860] = ~(layer0_outputs[2670]);
    assign layer1_outputs[7861] = 1'b0;
    assign layer1_outputs[7862] = ~(layer0_outputs[2463]);
    assign layer1_outputs[7863] = layer0_outputs[11709];
    assign layer1_outputs[7864] = ~((layer0_outputs[8]) & (layer0_outputs[11953]));
    assign layer1_outputs[7865] = ~(layer0_outputs[11413]);
    assign layer1_outputs[7866] = (layer0_outputs[8568]) ^ (layer0_outputs[6996]);
    assign layer1_outputs[7867] = ~(layer0_outputs[150]) | (layer0_outputs[3863]);
    assign layer1_outputs[7868] = (layer0_outputs[5538]) & ~(layer0_outputs[12734]);
    assign layer1_outputs[7869] = ~(layer0_outputs[2570]);
    assign layer1_outputs[7870] = ~(layer0_outputs[5608]);
    assign layer1_outputs[7871] = ~((layer0_outputs[4158]) & (layer0_outputs[12454]));
    assign layer1_outputs[7872] = ~(layer0_outputs[811]);
    assign layer1_outputs[7873] = (layer0_outputs[2396]) | (layer0_outputs[8594]);
    assign layer1_outputs[7874] = ~(layer0_outputs[944]);
    assign layer1_outputs[7875] = ~(layer0_outputs[2413]) | (layer0_outputs[11554]);
    assign layer1_outputs[7876] = ~(layer0_outputs[11852]);
    assign layer1_outputs[7877] = (layer0_outputs[4161]) ^ (layer0_outputs[3284]);
    assign layer1_outputs[7878] = ~((layer0_outputs[4308]) & (layer0_outputs[4145]));
    assign layer1_outputs[7879] = layer0_outputs[3485];
    assign layer1_outputs[7880] = ~((layer0_outputs[227]) & (layer0_outputs[5242]));
    assign layer1_outputs[7881] = ~(layer0_outputs[10057]) | (layer0_outputs[1793]);
    assign layer1_outputs[7882] = (layer0_outputs[1833]) & (layer0_outputs[5565]);
    assign layer1_outputs[7883] = ~((layer0_outputs[10014]) | (layer0_outputs[11919]));
    assign layer1_outputs[7884] = (layer0_outputs[11611]) ^ (layer0_outputs[11881]);
    assign layer1_outputs[7885] = layer0_outputs[10716];
    assign layer1_outputs[7886] = layer0_outputs[549];
    assign layer1_outputs[7887] = layer0_outputs[9351];
    assign layer1_outputs[7888] = 1'b0;
    assign layer1_outputs[7889] = ~((layer0_outputs[3156]) & (layer0_outputs[11551]));
    assign layer1_outputs[7890] = (layer0_outputs[9463]) & (layer0_outputs[2022]);
    assign layer1_outputs[7891] = ~(layer0_outputs[3059]);
    assign layer1_outputs[7892] = ~((layer0_outputs[6922]) ^ (layer0_outputs[12384]));
    assign layer1_outputs[7893] = (layer0_outputs[10210]) & (layer0_outputs[11625]);
    assign layer1_outputs[7894] = ~(layer0_outputs[1102]) | (layer0_outputs[671]);
    assign layer1_outputs[7895] = (layer0_outputs[172]) & ~(layer0_outputs[6091]);
    assign layer1_outputs[7896] = ~((layer0_outputs[5365]) & (layer0_outputs[7580]));
    assign layer1_outputs[7897] = ~((layer0_outputs[1506]) & (layer0_outputs[11136]));
    assign layer1_outputs[7898] = (layer0_outputs[8261]) & ~(layer0_outputs[2903]);
    assign layer1_outputs[7899] = 1'b0;
    assign layer1_outputs[7900] = (layer0_outputs[168]) | (layer0_outputs[10324]);
    assign layer1_outputs[7901] = 1'b1;
    assign layer1_outputs[7902] = (layer0_outputs[2728]) & (layer0_outputs[5300]);
    assign layer1_outputs[7903] = (layer0_outputs[5833]) & ~(layer0_outputs[2780]);
    assign layer1_outputs[7904] = ~(layer0_outputs[11608]) | (layer0_outputs[12314]);
    assign layer1_outputs[7905] = layer0_outputs[3239];
    assign layer1_outputs[7906] = layer0_outputs[2472];
    assign layer1_outputs[7907] = (layer0_outputs[1489]) | (layer0_outputs[12340]);
    assign layer1_outputs[7908] = (layer0_outputs[5949]) & ~(layer0_outputs[2737]);
    assign layer1_outputs[7909] = ~(layer0_outputs[10440]);
    assign layer1_outputs[7910] = ~((layer0_outputs[10961]) & (layer0_outputs[4344]));
    assign layer1_outputs[7911] = layer0_outputs[729];
    assign layer1_outputs[7912] = ~((layer0_outputs[6523]) | (layer0_outputs[8397]));
    assign layer1_outputs[7913] = ~((layer0_outputs[1955]) | (layer0_outputs[10917]));
    assign layer1_outputs[7914] = (layer0_outputs[11981]) ^ (layer0_outputs[2176]);
    assign layer1_outputs[7915] = ~(layer0_outputs[9290]);
    assign layer1_outputs[7916] = (layer0_outputs[12347]) & ~(layer0_outputs[1248]);
    assign layer1_outputs[7917] = layer0_outputs[10406];
    assign layer1_outputs[7918] = layer0_outputs[11698];
    assign layer1_outputs[7919] = 1'b1;
    assign layer1_outputs[7920] = layer0_outputs[7369];
    assign layer1_outputs[7921] = (layer0_outputs[3189]) | (layer0_outputs[10322]);
    assign layer1_outputs[7922] = (layer0_outputs[3851]) & (layer0_outputs[1634]);
    assign layer1_outputs[7923] = (layer0_outputs[6347]) | (layer0_outputs[8671]);
    assign layer1_outputs[7924] = ~(layer0_outputs[9385]);
    assign layer1_outputs[7925] = layer0_outputs[8876];
    assign layer1_outputs[7926] = ~(layer0_outputs[3599]) | (layer0_outputs[5770]);
    assign layer1_outputs[7927] = layer0_outputs[10703];
    assign layer1_outputs[7928] = (layer0_outputs[5857]) ^ (layer0_outputs[8195]);
    assign layer1_outputs[7929] = ~((layer0_outputs[8912]) & (layer0_outputs[2984]));
    assign layer1_outputs[7930] = layer0_outputs[9920];
    assign layer1_outputs[7931] = ~((layer0_outputs[9824]) ^ (layer0_outputs[10092]));
    assign layer1_outputs[7932] = ~((layer0_outputs[10910]) | (layer0_outputs[1640]));
    assign layer1_outputs[7933] = ~(layer0_outputs[606]);
    assign layer1_outputs[7934] = ~(layer0_outputs[2443]) | (layer0_outputs[1337]);
    assign layer1_outputs[7935] = ~((layer0_outputs[4202]) | (layer0_outputs[11434]));
    assign layer1_outputs[7936] = ~(layer0_outputs[10384]) | (layer0_outputs[3951]);
    assign layer1_outputs[7937] = layer0_outputs[6489];
    assign layer1_outputs[7938] = ~(layer0_outputs[6821]);
    assign layer1_outputs[7939] = (layer0_outputs[11204]) ^ (layer0_outputs[6626]);
    assign layer1_outputs[7940] = (layer0_outputs[11476]) | (layer0_outputs[816]);
    assign layer1_outputs[7941] = layer0_outputs[3353];
    assign layer1_outputs[7942] = (layer0_outputs[10237]) | (layer0_outputs[11989]);
    assign layer1_outputs[7943] = layer0_outputs[9288];
    assign layer1_outputs[7944] = ~(layer0_outputs[11917]) | (layer0_outputs[4938]);
    assign layer1_outputs[7945] = ~((layer0_outputs[5324]) | (layer0_outputs[12058]));
    assign layer1_outputs[7946] = ~(layer0_outputs[3895]);
    assign layer1_outputs[7947] = ~(layer0_outputs[9285]) | (layer0_outputs[7766]);
    assign layer1_outputs[7948] = layer0_outputs[11679];
    assign layer1_outputs[7949] = ~((layer0_outputs[11992]) ^ (layer0_outputs[3774]));
    assign layer1_outputs[7950] = ~(layer0_outputs[7681]) | (layer0_outputs[11904]);
    assign layer1_outputs[7951] = ~(layer0_outputs[6930]);
    assign layer1_outputs[7952] = layer0_outputs[6106];
    assign layer1_outputs[7953] = ~((layer0_outputs[10100]) & (layer0_outputs[8383]));
    assign layer1_outputs[7954] = ~(layer0_outputs[5221]) | (layer0_outputs[1857]);
    assign layer1_outputs[7955] = (layer0_outputs[3047]) ^ (layer0_outputs[12401]);
    assign layer1_outputs[7956] = layer0_outputs[12601];
    assign layer1_outputs[7957] = layer0_outputs[6613];
    assign layer1_outputs[7958] = ~(layer0_outputs[5076]);
    assign layer1_outputs[7959] = layer0_outputs[5398];
    assign layer1_outputs[7960] = ~((layer0_outputs[5653]) ^ (layer0_outputs[11050]));
    assign layer1_outputs[7961] = layer0_outputs[863];
    assign layer1_outputs[7962] = (layer0_outputs[8723]) ^ (layer0_outputs[2127]);
    assign layer1_outputs[7963] = layer0_outputs[12656];
    assign layer1_outputs[7964] = ~(layer0_outputs[7065]) | (layer0_outputs[12025]);
    assign layer1_outputs[7965] = ~((layer0_outputs[2564]) | (layer0_outputs[8424]));
    assign layer1_outputs[7966] = layer0_outputs[5156];
    assign layer1_outputs[7967] = ~(layer0_outputs[8067]);
    assign layer1_outputs[7968] = (layer0_outputs[2533]) ^ (layer0_outputs[11762]);
    assign layer1_outputs[7969] = (layer0_outputs[1747]) & (layer0_outputs[8877]);
    assign layer1_outputs[7970] = ~((layer0_outputs[5902]) ^ (layer0_outputs[7025]));
    assign layer1_outputs[7971] = ~((layer0_outputs[3562]) & (layer0_outputs[5383]));
    assign layer1_outputs[7972] = (layer0_outputs[8950]) | (layer0_outputs[3716]);
    assign layer1_outputs[7973] = (layer0_outputs[7692]) & (layer0_outputs[12780]);
    assign layer1_outputs[7974] = ~(layer0_outputs[2640]) | (layer0_outputs[7298]);
    assign layer1_outputs[7975] = ~(layer0_outputs[7382]);
    assign layer1_outputs[7976] = ~(layer0_outputs[10777]);
    assign layer1_outputs[7977] = layer0_outputs[9075];
    assign layer1_outputs[7978] = ~(layer0_outputs[1316]);
    assign layer1_outputs[7979] = ~(layer0_outputs[9417]) | (layer0_outputs[7275]);
    assign layer1_outputs[7980] = (layer0_outputs[12084]) & (layer0_outputs[4294]);
    assign layer1_outputs[7981] = (layer0_outputs[6461]) ^ (layer0_outputs[3290]);
    assign layer1_outputs[7982] = (layer0_outputs[1394]) ^ (layer0_outputs[2790]);
    assign layer1_outputs[7983] = ~(layer0_outputs[7892]);
    assign layer1_outputs[7984] = ~(layer0_outputs[7117]);
    assign layer1_outputs[7985] = ~(layer0_outputs[7791]);
    assign layer1_outputs[7986] = (layer0_outputs[9458]) & (layer0_outputs[2428]);
    assign layer1_outputs[7987] = ~(layer0_outputs[8601]) | (layer0_outputs[9639]);
    assign layer1_outputs[7988] = layer0_outputs[10198];
    assign layer1_outputs[7989] = 1'b0;
    assign layer1_outputs[7990] = (layer0_outputs[8180]) & ~(layer0_outputs[12085]);
    assign layer1_outputs[7991] = layer0_outputs[3048];
    assign layer1_outputs[7992] = ~((layer0_outputs[1666]) | (layer0_outputs[2658]));
    assign layer1_outputs[7993] = ~(layer0_outputs[8762]);
    assign layer1_outputs[7994] = (layer0_outputs[250]) & (layer0_outputs[3998]);
    assign layer1_outputs[7995] = layer0_outputs[7480];
    assign layer1_outputs[7996] = ~(layer0_outputs[10139]);
    assign layer1_outputs[7997] = ~(layer0_outputs[12600]) | (layer0_outputs[7165]);
    assign layer1_outputs[7998] = ~(layer0_outputs[8689]);
    assign layer1_outputs[7999] = (layer0_outputs[7750]) ^ (layer0_outputs[916]);
    assign layer1_outputs[8000] = ~((layer0_outputs[478]) | (layer0_outputs[7637]));
    assign layer1_outputs[8001] = layer0_outputs[2373];
    assign layer1_outputs[8002] = (layer0_outputs[2215]) ^ (layer0_outputs[2804]);
    assign layer1_outputs[8003] = (layer0_outputs[10633]) & ~(layer0_outputs[11372]);
    assign layer1_outputs[8004] = layer0_outputs[6935];
    assign layer1_outputs[8005] = layer0_outputs[10374];
    assign layer1_outputs[8006] = layer0_outputs[11158];
    assign layer1_outputs[8007] = (layer0_outputs[2032]) ^ (layer0_outputs[7487]);
    assign layer1_outputs[8008] = layer0_outputs[9335];
    assign layer1_outputs[8009] = (layer0_outputs[537]) & ~(layer0_outputs[10703]);
    assign layer1_outputs[8010] = ~(layer0_outputs[7746]);
    assign layer1_outputs[8011] = ~(layer0_outputs[3448]) | (layer0_outputs[9815]);
    assign layer1_outputs[8012] = ~((layer0_outputs[5723]) & (layer0_outputs[4695]));
    assign layer1_outputs[8013] = (layer0_outputs[10041]) & ~(layer0_outputs[1885]);
    assign layer1_outputs[8014] = ~(layer0_outputs[7552]);
    assign layer1_outputs[8015] = ~(layer0_outputs[10752]) | (layer0_outputs[6254]);
    assign layer1_outputs[8016] = ~(layer0_outputs[3396]);
    assign layer1_outputs[8017] = layer0_outputs[7302];
    assign layer1_outputs[8018] = ~(layer0_outputs[9583]);
    assign layer1_outputs[8019] = ~(layer0_outputs[2214]);
    assign layer1_outputs[8020] = layer0_outputs[7194];
    assign layer1_outputs[8021] = (layer0_outputs[8538]) & ~(layer0_outputs[7032]);
    assign layer1_outputs[8022] = ~((layer0_outputs[12101]) ^ (layer0_outputs[5386]));
    assign layer1_outputs[8023] = (layer0_outputs[856]) & ~(layer0_outputs[6313]);
    assign layer1_outputs[8024] = ~(layer0_outputs[2515]);
    assign layer1_outputs[8025] = (layer0_outputs[7559]) & ~(layer0_outputs[10434]);
    assign layer1_outputs[8026] = layer0_outputs[5812];
    assign layer1_outputs[8027] = layer0_outputs[7625];
    assign layer1_outputs[8028] = layer0_outputs[2405];
    assign layer1_outputs[8029] = 1'b1;
    assign layer1_outputs[8030] = (layer0_outputs[4131]) & ~(layer0_outputs[5754]);
    assign layer1_outputs[8031] = (layer0_outputs[1127]) & ~(layer0_outputs[2632]);
    assign layer1_outputs[8032] = layer0_outputs[4248];
    assign layer1_outputs[8033] = ~(layer0_outputs[6289]);
    assign layer1_outputs[8034] = (layer0_outputs[568]) & (layer0_outputs[1065]);
    assign layer1_outputs[8035] = ~((layer0_outputs[11332]) & (layer0_outputs[6387]));
    assign layer1_outputs[8036] = ~((layer0_outputs[11930]) & (layer0_outputs[1115]));
    assign layer1_outputs[8037] = layer0_outputs[6506];
    assign layer1_outputs[8038] = ~((layer0_outputs[7587]) ^ (layer0_outputs[1619]));
    assign layer1_outputs[8039] = ~(layer0_outputs[5478]);
    assign layer1_outputs[8040] = ~(layer0_outputs[738]) | (layer0_outputs[1503]);
    assign layer1_outputs[8041] = layer0_outputs[2239];
    assign layer1_outputs[8042] = (layer0_outputs[308]) & (layer0_outputs[11299]);
    assign layer1_outputs[8043] = ~(layer0_outputs[9905]);
    assign layer1_outputs[8044] = (layer0_outputs[5284]) & ~(layer0_outputs[1315]);
    assign layer1_outputs[8045] = layer0_outputs[4623];
    assign layer1_outputs[8046] = ~(layer0_outputs[1781]) | (layer0_outputs[2350]);
    assign layer1_outputs[8047] = ~((layer0_outputs[6675]) | (layer0_outputs[12518]));
    assign layer1_outputs[8048] = ~(layer0_outputs[3649]);
    assign layer1_outputs[8049] = ~((layer0_outputs[2500]) ^ (layer0_outputs[10331]));
    assign layer1_outputs[8050] = ~((layer0_outputs[1907]) | (layer0_outputs[1905]));
    assign layer1_outputs[8051] = (layer0_outputs[8571]) ^ (layer0_outputs[1543]);
    assign layer1_outputs[8052] = 1'b1;
    assign layer1_outputs[8053] = ~(layer0_outputs[12000]);
    assign layer1_outputs[8054] = layer0_outputs[7571];
    assign layer1_outputs[8055] = ~((layer0_outputs[6603]) & (layer0_outputs[7859]));
    assign layer1_outputs[8056] = ~((layer0_outputs[9639]) | (layer0_outputs[7490]));
    assign layer1_outputs[8057] = ~((layer0_outputs[8117]) & (layer0_outputs[8938]));
    assign layer1_outputs[8058] = ~((layer0_outputs[7655]) ^ (layer0_outputs[3867]));
    assign layer1_outputs[8059] = layer0_outputs[4840];
    assign layer1_outputs[8060] = ~((layer0_outputs[6842]) & (layer0_outputs[5882]));
    assign layer1_outputs[8061] = (layer0_outputs[11897]) & (layer0_outputs[176]);
    assign layer1_outputs[8062] = ~(layer0_outputs[3894]);
    assign layer1_outputs[8063] = (layer0_outputs[6687]) & (layer0_outputs[5260]);
    assign layer1_outputs[8064] = (layer0_outputs[10847]) & (layer0_outputs[4393]);
    assign layer1_outputs[8065] = layer0_outputs[624];
    assign layer1_outputs[8066] = ~(layer0_outputs[9571]);
    assign layer1_outputs[8067] = (layer0_outputs[11752]) | (layer0_outputs[10541]);
    assign layer1_outputs[8068] = ~((layer0_outputs[1441]) ^ (layer0_outputs[9505]));
    assign layer1_outputs[8069] = ~(layer0_outputs[10835]) | (layer0_outputs[11759]);
    assign layer1_outputs[8070] = layer0_outputs[8270];
    assign layer1_outputs[8071] = (layer0_outputs[9009]) ^ (layer0_outputs[538]);
    assign layer1_outputs[8072] = layer0_outputs[9807];
    assign layer1_outputs[8073] = (layer0_outputs[123]) ^ (layer0_outputs[4545]);
    assign layer1_outputs[8074] = (layer0_outputs[7354]) & (layer0_outputs[8753]);
    assign layer1_outputs[8075] = ~(layer0_outputs[2618]) | (layer0_outputs[5788]);
    assign layer1_outputs[8076] = layer0_outputs[4595];
    assign layer1_outputs[8077] = layer0_outputs[9419];
    assign layer1_outputs[8078] = (layer0_outputs[6309]) & (layer0_outputs[10609]);
    assign layer1_outputs[8079] = ~(layer0_outputs[10272]);
    assign layer1_outputs[8080] = ~(layer0_outputs[1788]) | (layer0_outputs[3435]);
    assign layer1_outputs[8081] = ~(layer0_outputs[9334]) | (layer0_outputs[5717]);
    assign layer1_outputs[8082] = ~((layer0_outputs[440]) & (layer0_outputs[8991]));
    assign layer1_outputs[8083] = (layer0_outputs[1154]) ^ (layer0_outputs[2415]);
    assign layer1_outputs[8084] = layer0_outputs[5952];
    assign layer1_outputs[8085] = ~(layer0_outputs[956]) | (layer0_outputs[2702]);
    assign layer1_outputs[8086] = ~((layer0_outputs[9600]) & (layer0_outputs[9945]));
    assign layer1_outputs[8087] = ~(layer0_outputs[1750]) | (layer0_outputs[6557]);
    assign layer1_outputs[8088] = ~(layer0_outputs[7014]) | (layer0_outputs[10665]);
    assign layer1_outputs[8089] = layer0_outputs[3905];
    assign layer1_outputs[8090] = ~(layer0_outputs[11907]);
    assign layer1_outputs[8091] = layer0_outputs[10174];
    assign layer1_outputs[8092] = (layer0_outputs[12682]) & (layer0_outputs[976]);
    assign layer1_outputs[8093] = (layer0_outputs[8867]) ^ (layer0_outputs[844]);
    assign layer1_outputs[8094] = ~((layer0_outputs[7352]) & (layer0_outputs[1887]));
    assign layer1_outputs[8095] = ~(layer0_outputs[6978]);
    assign layer1_outputs[8096] = layer0_outputs[8931];
    assign layer1_outputs[8097] = ~((layer0_outputs[10824]) | (layer0_outputs[11010]));
    assign layer1_outputs[8098] = layer0_outputs[9318];
    assign layer1_outputs[8099] = layer0_outputs[10139];
    assign layer1_outputs[8100] = (layer0_outputs[8826]) & ~(layer0_outputs[6145]);
    assign layer1_outputs[8101] = ~((layer0_outputs[1112]) & (layer0_outputs[1984]));
    assign layer1_outputs[8102] = ~(layer0_outputs[5157]) | (layer0_outputs[700]);
    assign layer1_outputs[8103] = (layer0_outputs[1937]) & (layer0_outputs[5607]);
    assign layer1_outputs[8104] = layer0_outputs[5853];
    assign layer1_outputs[8105] = (layer0_outputs[12440]) & (layer0_outputs[6004]);
    assign layer1_outputs[8106] = (layer0_outputs[3683]) & ~(layer0_outputs[8357]);
    assign layer1_outputs[8107] = ~(layer0_outputs[44]);
    assign layer1_outputs[8108] = ~(layer0_outputs[9616]);
    assign layer1_outputs[8109] = (layer0_outputs[3694]) | (layer0_outputs[6869]);
    assign layer1_outputs[8110] = layer0_outputs[7583];
    assign layer1_outputs[8111] = ~((layer0_outputs[5195]) ^ (layer0_outputs[4112]));
    assign layer1_outputs[8112] = layer0_outputs[8990];
    assign layer1_outputs[8113] = 1'b1;
    assign layer1_outputs[8114] = ~(layer0_outputs[3067]);
    assign layer1_outputs[8115] = (layer0_outputs[9558]) & (layer0_outputs[1426]);
    assign layer1_outputs[8116] = ~(layer0_outputs[12258]) | (layer0_outputs[8908]);
    assign layer1_outputs[8117] = ~((layer0_outputs[1686]) | (layer0_outputs[10774]));
    assign layer1_outputs[8118] = ~((layer0_outputs[6160]) & (layer0_outputs[1840]));
    assign layer1_outputs[8119] = ~(layer0_outputs[4029]);
    assign layer1_outputs[8120] = (layer0_outputs[3573]) & (layer0_outputs[7935]);
    assign layer1_outputs[8121] = ~(layer0_outputs[8433]);
    assign layer1_outputs[8122] = layer0_outputs[420];
    assign layer1_outputs[8123] = ~(layer0_outputs[9277]);
    assign layer1_outputs[8124] = layer0_outputs[5840];
    assign layer1_outputs[8125] = (layer0_outputs[7958]) & ~(layer0_outputs[3188]);
    assign layer1_outputs[8126] = layer0_outputs[4381];
    assign layer1_outputs[8127] = ~(layer0_outputs[3921]);
    assign layer1_outputs[8128] = ~((layer0_outputs[6051]) ^ (layer0_outputs[5499]));
    assign layer1_outputs[8129] = ~((layer0_outputs[2260]) & (layer0_outputs[241]));
    assign layer1_outputs[8130] = ~(layer0_outputs[4819]) | (layer0_outputs[10017]);
    assign layer1_outputs[8131] = ~(layer0_outputs[5967]);
    assign layer1_outputs[8132] = layer0_outputs[6322];
    assign layer1_outputs[8133] = ~(layer0_outputs[4191]);
    assign layer1_outputs[8134] = (layer0_outputs[10193]) ^ (layer0_outputs[3975]);
    assign layer1_outputs[8135] = layer0_outputs[1259];
    assign layer1_outputs[8136] = ~(layer0_outputs[7437]);
    assign layer1_outputs[8137] = (layer0_outputs[4790]) & ~(layer0_outputs[3874]);
    assign layer1_outputs[8138] = ~(layer0_outputs[5787]);
    assign layer1_outputs[8139] = layer0_outputs[920];
    assign layer1_outputs[8140] = (layer0_outputs[10591]) | (layer0_outputs[8875]);
    assign layer1_outputs[8141] = layer0_outputs[11196];
    assign layer1_outputs[8142] = ~(layer0_outputs[11298]);
    assign layer1_outputs[8143] = layer0_outputs[1385];
    assign layer1_outputs[8144] = ~((layer0_outputs[5237]) & (layer0_outputs[11788]));
    assign layer1_outputs[8145] = ~(layer0_outputs[6576]);
    assign layer1_outputs[8146] = ~(layer0_outputs[528]);
    assign layer1_outputs[8147] = ~(layer0_outputs[7738]);
    assign layer1_outputs[8148] = layer0_outputs[12099];
    assign layer1_outputs[8149] = ~(layer0_outputs[3289]);
    assign layer1_outputs[8150] = layer0_outputs[9902];
    assign layer1_outputs[8151] = ~((layer0_outputs[31]) | (layer0_outputs[4077]));
    assign layer1_outputs[8152] = layer0_outputs[9956];
    assign layer1_outputs[8153] = ~((layer0_outputs[3840]) ^ (layer0_outputs[6745]));
    assign layer1_outputs[8154] = (layer0_outputs[5320]) & ~(layer0_outputs[10353]);
    assign layer1_outputs[8155] = layer0_outputs[127];
    assign layer1_outputs[8156] = ~((layer0_outputs[10305]) & (layer0_outputs[1818]));
    assign layer1_outputs[8157] = ~(layer0_outputs[1772]) | (layer0_outputs[4413]);
    assign layer1_outputs[8158] = layer0_outputs[9423];
    assign layer1_outputs[8159] = ~(layer0_outputs[12712]);
    assign layer1_outputs[8160] = ~(layer0_outputs[697]);
    assign layer1_outputs[8161] = layer0_outputs[2340];
    assign layer1_outputs[8162] = (layer0_outputs[1683]) & ~(layer0_outputs[2762]);
    assign layer1_outputs[8163] = ~(layer0_outputs[8717]);
    assign layer1_outputs[8164] = ~(layer0_outputs[1008]);
    assign layer1_outputs[8165] = (layer0_outputs[6754]) | (layer0_outputs[4621]);
    assign layer1_outputs[8166] = 1'b0;
    assign layer1_outputs[8167] = (layer0_outputs[11922]) ^ (layer0_outputs[4401]);
    assign layer1_outputs[8168] = (layer0_outputs[5674]) & (layer0_outputs[4805]);
    assign layer1_outputs[8169] = layer0_outputs[11990];
    assign layer1_outputs[8170] = ~(layer0_outputs[9163]);
    assign layer1_outputs[8171] = (layer0_outputs[3220]) & ~(layer0_outputs[10403]);
    assign layer1_outputs[8172] = ~(layer0_outputs[740]);
    assign layer1_outputs[8173] = (layer0_outputs[11956]) & (layer0_outputs[2704]);
    assign layer1_outputs[8174] = ~((layer0_outputs[11326]) | (layer0_outputs[6799]));
    assign layer1_outputs[8175] = layer0_outputs[4990];
    assign layer1_outputs[8176] = ~(layer0_outputs[167]);
    assign layer1_outputs[8177] = (layer0_outputs[2417]) & (layer0_outputs[6970]);
    assign layer1_outputs[8178] = (layer0_outputs[9249]) | (layer0_outputs[9029]);
    assign layer1_outputs[8179] = ~((layer0_outputs[2322]) | (layer0_outputs[2553]));
    assign layer1_outputs[8180] = ~(layer0_outputs[1884]) | (layer0_outputs[5018]);
    assign layer1_outputs[8181] = (layer0_outputs[5632]) ^ (layer0_outputs[2587]);
    assign layer1_outputs[8182] = 1'b1;
    assign layer1_outputs[8183] = (layer0_outputs[3396]) & ~(layer0_outputs[7160]);
    assign layer1_outputs[8184] = ~(layer0_outputs[2858]);
    assign layer1_outputs[8185] = ~((layer0_outputs[7272]) | (layer0_outputs[12793]));
    assign layer1_outputs[8186] = layer0_outputs[7698];
    assign layer1_outputs[8187] = layer0_outputs[5185];
    assign layer1_outputs[8188] = (layer0_outputs[326]) & ~(layer0_outputs[9829]);
    assign layer1_outputs[8189] = ~(layer0_outputs[3512]);
    assign layer1_outputs[8190] = layer0_outputs[8106];
    assign layer1_outputs[8191] = ~(layer0_outputs[21]) | (layer0_outputs[8839]);
    assign layer1_outputs[8192] = layer0_outputs[4349];
    assign layer1_outputs[8193] = (layer0_outputs[7316]) ^ (layer0_outputs[3021]);
    assign layer1_outputs[8194] = layer0_outputs[10785];
    assign layer1_outputs[8195] = ~(layer0_outputs[9453]);
    assign layer1_outputs[8196] = ~(layer0_outputs[3320]);
    assign layer1_outputs[8197] = (layer0_outputs[6918]) & (layer0_outputs[4853]);
    assign layer1_outputs[8198] = ~((layer0_outputs[6501]) ^ (layer0_outputs[5208]));
    assign layer1_outputs[8199] = ~(layer0_outputs[2770]);
    assign layer1_outputs[8200] = (layer0_outputs[4410]) & ~(layer0_outputs[7544]);
    assign layer1_outputs[8201] = 1'b0;
    assign layer1_outputs[8202] = (layer0_outputs[1273]) ^ (layer0_outputs[1055]);
    assign layer1_outputs[8203] = layer0_outputs[3980];
    assign layer1_outputs[8204] = layer0_outputs[906];
    assign layer1_outputs[8205] = 1'b0;
    assign layer1_outputs[8206] = ~(layer0_outputs[12130]) | (layer0_outputs[9281]);
    assign layer1_outputs[8207] = ~(layer0_outputs[10321]);
    assign layer1_outputs[8208] = ~(layer0_outputs[3847]);
    assign layer1_outputs[8209] = ~((layer0_outputs[5304]) | (layer0_outputs[8676]));
    assign layer1_outputs[8210] = ~(layer0_outputs[405]);
    assign layer1_outputs[8211] = ~(layer0_outputs[9464]) | (layer0_outputs[9947]);
    assign layer1_outputs[8212] = (layer0_outputs[3904]) & ~(layer0_outputs[8705]);
    assign layer1_outputs[8213] = (layer0_outputs[11857]) & ~(layer0_outputs[718]);
    assign layer1_outputs[8214] = ~((layer0_outputs[2869]) & (layer0_outputs[7468]));
    assign layer1_outputs[8215] = (layer0_outputs[1367]) | (layer0_outputs[2065]);
    assign layer1_outputs[8216] = ~(layer0_outputs[10870]);
    assign layer1_outputs[8217] = ~((layer0_outputs[11717]) | (layer0_outputs[6096]));
    assign layer1_outputs[8218] = 1'b0;
    assign layer1_outputs[8219] = (layer0_outputs[10186]) & (layer0_outputs[6633]);
    assign layer1_outputs[8220] = ~(layer0_outputs[9169]);
    assign layer1_outputs[8221] = layer0_outputs[2333];
    assign layer1_outputs[8222] = ~(layer0_outputs[1894]);
    assign layer1_outputs[8223] = ~((layer0_outputs[2982]) ^ (layer0_outputs[84]));
    assign layer1_outputs[8224] = 1'b0;
    assign layer1_outputs[8225] = layer0_outputs[12611];
    assign layer1_outputs[8226] = (layer0_outputs[10809]) | (layer0_outputs[4804]);
    assign layer1_outputs[8227] = ~(layer0_outputs[4946]) | (layer0_outputs[12135]);
    assign layer1_outputs[8228] = ~(layer0_outputs[10705]);
    assign layer1_outputs[8229] = ~(layer0_outputs[6905]);
    assign layer1_outputs[8230] = ~(layer0_outputs[12018]);
    assign layer1_outputs[8231] = (layer0_outputs[3490]) | (layer0_outputs[7249]);
    assign layer1_outputs[8232] = layer0_outputs[6359];
    assign layer1_outputs[8233] = (layer0_outputs[8407]) & ~(layer0_outputs[1677]);
    assign layer1_outputs[8234] = ~(layer0_outputs[5270]) | (layer0_outputs[12048]);
    assign layer1_outputs[8235] = layer0_outputs[5070];
    assign layer1_outputs[8236] = ~(layer0_outputs[8544]);
    assign layer1_outputs[8237] = ~((layer0_outputs[8110]) ^ (layer0_outputs[10707]));
    assign layer1_outputs[8238] = (layer0_outputs[4767]) & ~(layer0_outputs[6284]);
    assign layer1_outputs[8239] = ~((layer0_outputs[6018]) | (layer0_outputs[8440]));
    assign layer1_outputs[8240] = ~((layer0_outputs[3891]) ^ (layer0_outputs[12109]));
    assign layer1_outputs[8241] = layer0_outputs[1913];
    assign layer1_outputs[8242] = layer0_outputs[9629];
    assign layer1_outputs[8243] = 1'b1;
    assign layer1_outputs[8244] = ~(layer0_outputs[7030]) | (layer0_outputs[3751]);
    assign layer1_outputs[8245] = ~(layer0_outputs[10113]);
    assign layer1_outputs[8246] = layer0_outputs[6845];
    assign layer1_outputs[8247] = layer0_outputs[11942];
    assign layer1_outputs[8248] = ~((layer0_outputs[5122]) ^ (layer0_outputs[8794]));
    assign layer1_outputs[8249] = layer0_outputs[9739];
    assign layer1_outputs[8250] = layer0_outputs[8398];
    assign layer1_outputs[8251] = (layer0_outputs[10730]) & (layer0_outputs[6808]);
    assign layer1_outputs[8252] = ~(layer0_outputs[3681]);
    assign layer1_outputs[8253] = ~(layer0_outputs[4526]) | (layer0_outputs[11333]);
    assign layer1_outputs[8254] = (layer0_outputs[5785]) & ~(layer0_outputs[5327]);
    assign layer1_outputs[8255] = ~((layer0_outputs[4647]) ^ (layer0_outputs[5590]));
    assign layer1_outputs[8256] = 1'b1;
    assign layer1_outputs[8257] = (layer0_outputs[7165]) & (layer0_outputs[11922]);
    assign layer1_outputs[8258] = ~(layer0_outputs[9069]);
    assign layer1_outputs[8259] = ~((layer0_outputs[11208]) | (layer0_outputs[11134]));
    assign layer1_outputs[8260] = ~((layer0_outputs[3004]) & (layer0_outputs[2996]));
    assign layer1_outputs[8261] = ~(layer0_outputs[8249]) | (layer0_outputs[3321]);
    assign layer1_outputs[8262] = layer0_outputs[11039];
    assign layer1_outputs[8263] = ~(layer0_outputs[3360]) | (layer0_outputs[3420]);
    assign layer1_outputs[8264] = ~((layer0_outputs[8043]) & (layer0_outputs[755]));
    assign layer1_outputs[8265] = ~((layer0_outputs[4924]) | (layer0_outputs[6939]));
    assign layer1_outputs[8266] = ~((layer0_outputs[215]) ^ (layer0_outputs[5083]));
    assign layer1_outputs[8267] = ~((layer0_outputs[113]) & (layer0_outputs[2482]));
    assign layer1_outputs[8268] = (layer0_outputs[466]) ^ (layer0_outputs[6993]);
    assign layer1_outputs[8269] = ~((layer0_outputs[1313]) ^ (layer0_outputs[6438]));
    assign layer1_outputs[8270] = ~(layer0_outputs[4359]) | (layer0_outputs[12293]);
    assign layer1_outputs[8271] = (layer0_outputs[8089]) & (layer0_outputs[7837]);
    assign layer1_outputs[8272] = ~((layer0_outputs[12492]) ^ (layer0_outputs[2279]));
    assign layer1_outputs[8273] = ~(layer0_outputs[7446]) | (layer0_outputs[1329]);
    assign layer1_outputs[8274] = ~(layer0_outputs[9964]) | (layer0_outputs[10402]);
    assign layer1_outputs[8275] = ~(layer0_outputs[7738]);
    assign layer1_outputs[8276] = ~((layer0_outputs[4115]) | (layer0_outputs[11571]));
    assign layer1_outputs[8277] = (layer0_outputs[9908]) & (layer0_outputs[4027]);
    assign layer1_outputs[8278] = 1'b0;
    assign layer1_outputs[8279] = layer0_outputs[6810];
    assign layer1_outputs[8280] = (layer0_outputs[248]) & ~(layer0_outputs[6360]);
    assign layer1_outputs[8281] = layer0_outputs[9197];
    assign layer1_outputs[8282] = layer0_outputs[1385];
    assign layer1_outputs[8283] = (layer0_outputs[7408]) & ~(layer0_outputs[6892]);
    assign layer1_outputs[8284] = (layer0_outputs[2370]) ^ (layer0_outputs[11482]);
    assign layer1_outputs[8285] = ~(layer0_outputs[8895]);
    assign layer1_outputs[8286] = ~(layer0_outputs[12334]) | (layer0_outputs[9438]);
    assign layer1_outputs[8287] = (layer0_outputs[11085]) & (layer0_outputs[7580]);
    assign layer1_outputs[8288] = (layer0_outputs[3594]) & (layer0_outputs[6264]);
    assign layer1_outputs[8289] = ~(layer0_outputs[1792]);
    assign layer1_outputs[8290] = layer0_outputs[4754];
    assign layer1_outputs[8291] = layer0_outputs[2604];
    assign layer1_outputs[8292] = (layer0_outputs[2759]) & ~(layer0_outputs[11215]);
    assign layer1_outputs[8293] = ~((layer0_outputs[7974]) | (layer0_outputs[12]));
    assign layer1_outputs[8294] = ~(layer0_outputs[11747]);
    assign layer1_outputs[8295] = (layer0_outputs[8825]) ^ (layer0_outputs[6255]);
    assign layer1_outputs[8296] = ~(layer0_outputs[6057]);
    assign layer1_outputs[8297] = (layer0_outputs[7007]) & ~(layer0_outputs[10508]);
    assign layer1_outputs[8298] = ~(layer0_outputs[6029]);
    assign layer1_outputs[8299] = ~(layer0_outputs[10256]);
    assign layer1_outputs[8300] = ~(layer0_outputs[9492]);
    assign layer1_outputs[8301] = 1'b1;
    assign layer1_outputs[8302] = ~((layer0_outputs[11305]) ^ (layer0_outputs[7087]));
    assign layer1_outputs[8303] = ~(layer0_outputs[2600]);
    assign layer1_outputs[8304] = layer0_outputs[3661];
    assign layer1_outputs[8305] = ~((layer0_outputs[5372]) | (layer0_outputs[957]));
    assign layer1_outputs[8306] = layer0_outputs[7879];
    assign layer1_outputs[8307] = layer0_outputs[11370];
    assign layer1_outputs[8308] = (layer0_outputs[7429]) & ~(layer0_outputs[10422]);
    assign layer1_outputs[8309] = ~(layer0_outputs[10993]);
    assign layer1_outputs[8310] = layer0_outputs[9792];
    assign layer1_outputs[8311] = ~(layer0_outputs[564]);
    assign layer1_outputs[8312] = ~(layer0_outputs[64]);
    assign layer1_outputs[8313] = layer0_outputs[5458];
    assign layer1_outputs[8314] = layer0_outputs[11359];
    assign layer1_outputs[8315] = layer0_outputs[92];
    assign layer1_outputs[8316] = (layer0_outputs[3993]) | (layer0_outputs[2186]);
    assign layer1_outputs[8317] = ~(layer0_outputs[11194]);
    assign layer1_outputs[8318] = layer0_outputs[4839];
    assign layer1_outputs[8319] = layer0_outputs[10466];
    assign layer1_outputs[8320] = ~(layer0_outputs[9035]);
    assign layer1_outputs[8321] = (layer0_outputs[8082]) ^ (layer0_outputs[11157]);
    assign layer1_outputs[8322] = (layer0_outputs[5987]) | (layer0_outputs[740]);
    assign layer1_outputs[8323] = ~(layer0_outputs[7649]);
    assign layer1_outputs[8324] = ~(layer0_outputs[7930]);
    assign layer1_outputs[8325] = ~(layer0_outputs[268]);
    assign layer1_outputs[8326] = ~(layer0_outputs[2493]);
    assign layer1_outputs[8327] = ~((layer0_outputs[1794]) ^ (layer0_outputs[12261]));
    assign layer1_outputs[8328] = (layer0_outputs[5182]) & ~(layer0_outputs[9875]);
    assign layer1_outputs[8329] = ~(layer0_outputs[10689]) | (layer0_outputs[11929]);
    assign layer1_outputs[8330] = ~((layer0_outputs[1390]) | (layer0_outputs[4538]));
    assign layer1_outputs[8331] = (layer0_outputs[7698]) & ~(layer0_outputs[12037]);
    assign layer1_outputs[8332] = (layer0_outputs[6963]) & ~(layer0_outputs[12074]);
    assign layer1_outputs[8333] = ~(layer0_outputs[11988]);
    assign layer1_outputs[8334] = ~(layer0_outputs[5068]);
    assign layer1_outputs[8335] = ~(layer0_outputs[3437]) | (layer0_outputs[7443]);
    assign layer1_outputs[8336] = ~(layer0_outputs[7027]);
    assign layer1_outputs[8337] = layer0_outputs[10221];
    assign layer1_outputs[8338] = (layer0_outputs[5996]) & ~(layer0_outputs[3668]);
    assign layer1_outputs[8339] = (layer0_outputs[7679]) | (layer0_outputs[11656]);
    assign layer1_outputs[8340] = (layer0_outputs[5716]) | (layer0_outputs[12777]);
    assign layer1_outputs[8341] = ~(layer0_outputs[6761]) | (layer0_outputs[12377]);
    assign layer1_outputs[8342] = ~((layer0_outputs[6095]) | (layer0_outputs[11219]));
    assign layer1_outputs[8343] = (layer0_outputs[4843]) & ~(layer0_outputs[494]);
    assign layer1_outputs[8344] = ~(layer0_outputs[12644]) | (layer0_outputs[8403]);
    assign layer1_outputs[8345] = (layer0_outputs[11731]) & ~(layer0_outputs[11623]);
    assign layer1_outputs[8346] = layer0_outputs[2666];
    assign layer1_outputs[8347] = ~((layer0_outputs[3890]) & (layer0_outputs[5212]));
    assign layer1_outputs[8348] = ~(layer0_outputs[1648]) | (layer0_outputs[9087]);
    assign layer1_outputs[8349] = ~((layer0_outputs[5039]) ^ (layer0_outputs[10884]));
    assign layer1_outputs[8350] = ~(layer0_outputs[427]);
    assign layer1_outputs[8351] = ~(layer0_outputs[12168]) | (layer0_outputs[6895]);
    assign layer1_outputs[8352] = ~(layer0_outputs[10380]);
    assign layer1_outputs[8353] = (layer0_outputs[9502]) & ~(layer0_outputs[9724]);
    assign layer1_outputs[8354] = layer0_outputs[7226];
    assign layer1_outputs[8355] = layer0_outputs[7491];
    assign layer1_outputs[8356] = layer0_outputs[8851];
    assign layer1_outputs[8357] = ~(layer0_outputs[10683]);
    assign layer1_outputs[8358] = ~((layer0_outputs[11214]) & (layer0_outputs[7167]));
    assign layer1_outputs[8359] = (layer0_outputs[2147]) & ~(layer0_outputs[12590]);
    assign layer1_outputs[8360] = (layer0_outputs[10403]) & (layer0_outputs[10514]);
    assign layer1_outputs[8361] = layer0_outputs[7691];
    assign layer1_outputs[8362] = ~(layer0_outputs[7709]);
    assign layer1_outputs[8363] = ~(layer0_outputs[10773]);
    assign layer1_outputs[8364] = ~(layer0_outputs[6519]);
    assign layer1_outputs[8365] = layer0_outputs[11190];
    assign layer1_outputs[8366] = (layer0_outputs[10561]) & (layer0_outputs[452]);
    assign layer1_outputs[8367] = layer0_outputs[4332];
    assign layer1_outputs[8368] = ~(layer0_outputs[6176]);
    assign layer1_outputs[8369] = layer0_outputs[2257];
    assign layer1_outputs[8370] = ~(layer0_outputs[2238]);
    assign layer1_outputs[8371] = (layer0_outputs[10453]) & (layer0_outputs[1605]);
    assign layer1_outputs[8372] = ~(layer0_outputs[6499]);
    assign layer1_outputs[8373] = ~(layer0_outputs[6773]) | (layer0_outputs[7839]);
    assign layer1_outputs[8374] = ~(layer0_outputs[7253]);
    assign layer1_outputs[8375] = ~((layer0_outputs[4033]) & (layer0_outputs[6625]));
    assign layer1_outputs[8376] = ~(layer0_outputs[12129]) | (layer0_outputs[11525]);
    assign layer1_outputs[8377] = (layer0_outputs[8199]) & ~(layer0_outputs[11678]);
    assign layer1_outputs[8378] = layer0_outputs[11167];
    assign layer1_outputs[8379] = ~((layer0_outputs[11765]) | (layer0_outputs[10959]));
    assign layer1_outputs[8380] = ~(layer0_outputs[4499]);
    assign layer1_outputs[8381] = ~(layer0_outputs[3121]) | (layer0_outputs[5859]);
    assign layer1_outputs[8382] = (layer0_outputs[9021]) & ~(layer0_outputs[2729]);
    assign layer1_outputs[8383] = ~(layer0_outputs[7802]) | (layer0_outputs[6619]);
    assign layer1_outputs[8384] = ~((layer0_outputs[10958]) ^ (layer0_outputs[6032]));
    assign layer1_outputs[8385] = layer0_outputs[12558];
    assign layer1_outputs[8386] = layer0_outputs[7935];
    assign layer1_outputs[8387] = (layer0_outputs[11031]) | (layer0_outputs[10074]);
    assign layer1_outputs[8388] = layer0_outputs[11022];
    assign layer1_outputs[8389] = ~(layer0_outputs[2599]);
    assign layer1_outputs[8390] = (layer0_outputs[6410]) & ~(layer0_outputs[7832]);
    assign layer1_outputs[8391] = (layer0_outputs[9939]) & ~(layer0_outputs[1859]);
    assign layer1_outputs[8392] = 1'b0;
    assign layer1_outputs[8393] = ~((layer0_outputs[2509]) ^ (layer0_outputs[8591]));
    assign layer1_outputs[8394] = 1'b1;
    assign layer1_outputs[8395] = 1'b0;
    assign layer1_outputs[8396] = ~((layer0_outputs[9567]) ^ (layer0_outputs[10913]));
    assign layer1_outputs[8397] = (layer0_outputs[963]) & ~(layer0_outputs[1023]);
    assign layer1_outputs[8398] = ~(layer0_outputs[8641]);
    assign layer1_outputs[8399] = layer0_outputs[7453];
    assign layer1_outputs[8400] = ~(layer0_outputs[1779]);
    assign layer1_outputs[8401] = ~(layer0_outputs[10023]) | (layer0_outputs[1683]);
    assign layer1_outputs[8402] = ~((layer0_outputs[10452]) & (layer0_outputs[5351]));
    assign layer1_outputs[8403] = layer0_outputs[5460];
    assign layer1_outputs[8404] = ~(layer0_outputs[4388]) | (layer0_outputs[8612]);
    assign layer1_outputs[8405] = (layer0_outputs[3262]) & (layer0_outputs[2411]);
    assign layer1_outputs[8406] = (layer0_outputs[12317]) & ~(layer0_outputs[2502]);
    assign layer1_outputs[8407] = layer0_outputs[12589];
    assign layer1_outputs[8408] = layer0_outputs[9718];
    assign layer1_outputs[8409] = (layer0_outputs[4896]) | (layer0_outputs[5038]);
    assign layer1_outputs[8410] = ~((layer0_outputs[45]) & (layer0_outputs[8828]));
    assign layer1_outputs[8411] = (layer0_outputs[9918]) & ~(layer0_outputs[8642]);
    assign layer1_outputs[8412] = ~((layer0_outputs[5380]) ^ (layer0_outputs[1180]));
    assign layer1_outputs[8413] = layer0_outputs[349];
    assign layer1_outputs[8414] = layer0_outputs[12229];
    assign layer1_outputs[8415] = (layer0_outputs[9667]) ^ (layer0_outputs[9783]);
    assign layer1_outputs[8416] = ~((layer0_outputs[6071]) & (layer0_outputs[1852]));
    assign layer1_outputs[8417] = ~(layer0_outputs[1130]);
    assign layer1_outputs[8418] = layer0_outputs[6840];
    assign layer1_outputs[8419] = (layer0_outputs[3673]) & (layer0_outputs[7963]);
    assign layer1_outputs[8420] = (layer0_outputs[7356]) & (layer0_outputs[7940]);
    assign layer1_outputs[8421] = ~(layer0_outputs[747]) | (layer0_outputs[5197]);
    assign layer1_outputs[8422] = (layer0_outputs[181]) & ~(layer0_outputs[4429]);
    assign layer1_outputs[8423] = (layer0_outputs[1943]) ^ (layer0_outputs[5655]);
    assign layer1_outputs[8424] = layer0_outputs[9147];
    assign layer1_outputs[8425] = layer0_outputs[2753];
    assign layer1_outputs[8426] = (layer0_outputs[602]) & ~(layer0_outputs[5550]);
    assign layer1_outputs[8427] = ~((layer0_outputs[6864]) ^ (layer0_outputs[157]));
    assign layer1_outputs[8428] = ~((layer0_outputs[10174]) & (layer0_outputs[168]));
    assign layer1_outputs[8429] = ~((layer0_outputs[9312]) ^ (layer0_outputs[11129]));
    assign layer1_outputs[8430] = (layer0_outputs[3827]) | (layer0_outputs[8010]);
    assign layer1_outputs[8431] = (layer0_outputs[1146]) & ~(layer0_outputs[10234]);
    assign layer1_outputs[8432] = ~(layer0_outputs[9429]);
    assign layer1_outputs[8433] = (layer0_outputs[8582]) & (layer0_outputs[7039]);
    assign layer1_outputs[8434] = layer0_outputs[11790];
    assign layer1_outputs[8435] = (layer0_outputs[1019]) & (layer0_outputs[12456]);
    assign layer1_outputs[8436] = ~(layer0_outputs[7907]);
    assign layer1_outputs[8437] = layer0_outputs[6149];
    assign layer1_outputs[8438] = (layer0_outputs[2938]) & (layer0_outputs[1359]);
    assign layer1_outputs[8439] = (layer0_outputs[10573]) | (layer0_outputs[10202]);
    assign layer1_outputs[8440] = ~(layer0_outputs[645]) | (layer0_outputs[1010]);
    assign layer1_outputs[8441] = (layer0_outputs[3371]) & ~(layer0_outputs[2603]);
    assign layer1_outputs[8442] = ~(layer0_outputs[8366]);
    assign layer1_outputs[8443] = layer0_outputs[322];
    assign layer1_outputs[8444] = layer0_outputs[10672];
    assign layer1_outputs[8445] = ~(layer0_outputs[12517]);
    assign layer1_outputs[8446] = ~((layer0_outputs[7881]) | (layer0_outputs[8595]));
    assign layer1_outputs[8447] = ~(layer0_outputs[6868]);
    assign layer1_outputs[8448] = (layer0_outputs[591]) & (layer0_outputs[2028]);
    assign layer1_outputs[8449] = layer0_outputs[9231];
    assign layer1_outputs[8450] = ~(layer0_outputs[1488]);
    assign layer1_outputs[8451] = ~((layer0_outputs[8432]) & (layer0_outputs[6059]));
    assign layer1_outputs[8452] = (layer0_outputs[9674]) & ~(layer0_outputs[9763]);
    assign layer1_outputs[8453] = (layer0_outputs[4931]) & (layer0_outputs[112]);
    assign layer1_outputs[8454] = layer0_outputs[4459];
    assign layer1_outputs[8455] = (layer0_outputs[1415]) & (layer0_outputs[5906]);
    assign layer1_outputs[8456] = ~(layer0_outputs[3955]);
    assign layer1_outputs[8457] = layer0_outputs[2042];
    assign layer1_outputs[8458] = layer0_outputs[5361];
    assign layer1_outputs[8459] = layer0_outputs[11200];
    assign layer1_outputs[8460] = layer0_outputs[4625];
    assign layer1_outputs[8461] = ~((layer0_outputs[1365]) | (layer0_outputs[7310]));
    assign layer1_outputs[8462] = (layer0_outputs[6656]) & ~(layer0_outputs[11458]);
    assign layer1_outputs[8463] = (layer0_outputs[2380]) & (layer0_outputs[10290]);
    assign layer1_outputs[8464] = ~((layer0_outputs[10156]) & (layer0_outputs[12457]));
    assign layer1_outputs[8465] = layer0_outputs[10966];
    assign layer1_outputs[8466] = layer0_outputs[5232];
    assign layer1_outputs[8467] = ~((layer0_outputs[9998]) ^ (layer0_outputs[12662]));
    assign layer1_outputs[8468] = (layer0_outputs[8457]) & (layer0_outputs[2907]);
    assign layer1_outputs[8469] = ~(layer0_outputs[12388]);
    assign layer1_outputs[8470] = ~((layer0_outputs[3433]) & (layer0_outputs[10992]));
    assign layer1_outputs[8471] = ~((layer0_outputs[11092]) & (layer0_outputs[7717]));
    assign layer1_outputs[8472] = layer0_outputs[3814];
    assign layer1_outputs[8473] = layer0_outputs[1574];
    assign layer1_outputs[8474] = layer0_outputs[5848];
    assign layer1_outputs[8475] = layer0_outputs[12531];
    assign layer1_outputs[8476] = ~(layer0_outputs[6362]) | (layer0_outputs[3461]);
    assign layer1_outputs[8477] = ~((layer0_outputs[6986]) | (layer0_outputs[3671]));
    assign layer1_outputs[8478] = (layer0_outputs[450]) & ~(layer0_outputs[7507]);
    assign layer1_outputs[8479] = layer0_outputs[11361];
    assign layer1_outputs[8480] = ~(layer0_outputs[2287]) | (layer0_outputs[12017]);
    assign layer1_outputs[8481] = (layer0_outputs[2483]) | (layer0_outputs[2437]);
    assign layer1_outputs[8482] = ~(layer0_outputs[11280]) | (layer0_outputs[5538]);
    assign layer1_outputs[8483] = ~(layer0_outputs[7695]);
    assign layer1_outputs[8484] = ~(layer0_outputs[2713]) | (layer0_outputs[8895]);
    assign layer1_outputs[8485] = ~(layer0_outputs[990]);
    assign layer1_outputs[8486] = ~(layer0_outputs[5153]) | (layer0_outputs[8241]);
    assign layer1_outputs[8487] = (layer0_outputs[12654]) ^ (layer0_outputs[3805]);
    assign layer1_outputs[8488] = ~((layer0_outputs[3861]) | (layer0_outputs[1294]));
    assign layer1_outputs[8489] = (layer0_outputs[9104]) | (layer0_outputs[7197]);
    assign layer1_outputs[8490] = ~((layer0_outputs[5704]) | (layer0_outputs[5077]));
    assign layer1_outputs[8491] = layer0_outputs[4166];
    assign layer1_outputs[8492] = ~(layer0_outputs[7045]);
    assign layer1_outputs[8493] = (layer0_outputs[4324]) & ~(layer0_outputs[2108]);
    assign layer1_outputs[8494] = layer0_outputs[5396];
    assign layer1_outputs[8495] = layer0_outputs[8543];
    assign layer1_outputs[8496] = ~(layer0_outputs[2681]);
    assign layer1_outputs[8497] = ~(layer0_outputs[7564]);
    assign layer1_outputs[8498] = ~((layer0_outputs[1059]) & (layer0_outputs[4032]));
    assign layer1_outputs[8499] = ~(layer0_outputs[3139]) | (layer0_outputs[9610]);
    assign layer1_outputs[8500] = ~((layer0_outputs[10313]) ^ (layer0_outputs[11315]));
    assign layer1_outputs[8501] = layer0_outputs[5441];
    assign layer1_outputs[8502] = ~(layer0_outputs[2087]);
    assign layer1_outputs[8503] = (layer0_outputs[8937]) ^ (layer0_outputs[12485]);
    assign layer1_outputs[8504] = ~(layer0_outputs[9667]);
    assign layer1_outputs[8505] = ~(layer0_outputs[3625]);
    assign layer1_outputs[8506] = ~(layer0_outputs[9726]);
    assign layer1_outputs[8507] = ~(layer0_outputs[6326]);
    assign layer1_outputs[8508] = ~(layer0_outputs[10545]);
    assign layer1_outputs[8509] = ~(layer0_outputs[11648]);
    assign layer1_outputs[8510] = ~((layer0_outputs[7729]) & (layer0_outputs[11045]));
    assign layer1_outputs[8511] = layer0_outputs[3225];
    assign layer1_outputs[8512] = ~((layer0_outputs[1132]) & (layer0_outputs[2085]));
    assign layer1_outputs[8513] = ~(layer0_outputs[3854]) | (layer0_outputs[2384]);
    assign layer1_outputs[8514] = ~((layer0_outputs[1074]) & (layer0_outputs[4213]));
    assign layer1_outputs[8515] = ~(layer0_outputs[5844]);
    assign layer1_outputs[8516] = ~(layer0_outputs[8619]);
    assign layer1_outputs[8517] = ~(layer0_outputs[11580]);
    assign layer1_outputs[8518] = (layer0_outputs[12426]) & ~(layer0_outputs[8953]);
    assign layer1_outputs[8519] = ~((layer0_outputs[10281]) & (layer0_outputs[6434]));
    assign layer1_outputs[8520] = ~((layer0_outputs[4914]) | (layer0_outputs[1680]));
    assign layer1_outputs[8521] = ~(layer0_outputs[6556]);
    assign layer1_outputs[8522] = (layer0_outputs[10026]) | (layer0_outputs[1133]);
    assign layer1_outputs[8523] = (layer0_outputs[2687]) & ~(layer0_outputs[7785]);
    assign layer1_outputs[8524] = ~((layer0_outputs[2129]) | (layer0_outputs[7591]));
    assign layer1_outputs[8525] = (layer0_outputs[12521]) | (layer0_outputs[6376]);
    assign layer1_outputs[8526] = layer0_outputs[7426];
    assign layer1_outputs[8527] = (layer0_outputs[7531]) ^ (layer0_outputs[11313]);
    assign layer1_outputs[8528] = (layer0_outputs[8431]) & ~(layer0_outputs[10024]);
    assign layer1_outputs[8529] = (layer0_outputs[319]) & ~(layer0_outputs[351]);
    assign layer1_outputs[8530] = (layer0_outputs[9328]) & ~(layer0_outputs[2561]);
    assign layer1_outputs[8531] = ~((layer0_outputs[6061]) & (layer0_outputs[6853]));
    assign layer1_outputs[8532] = layer0_outputs[8185];
    assign layer1_outputs[8533] = (layer0_outputs[11373]) & ~(layer0_outputs[1723]);
    assign layer1_outputs[8534] = ~(layer0_outputs[12665]);
    assign layer1_outputs[8535] = layer0_outputs[12026];
    assign layer1_outputs[8536] = ~(layer0_outputs[7369]);
    assign layer1_outputs[8537] = ~(layer0_outputs[6413]) | (layer0_outputs[9300]);
    assign layer1_outputs[8538] = ~((layer0_outputs[9386]) ^ (layer0_outputs[8932]));
    assign layer1_outputs[8539] = layer0_outputs[4968];
    assign layer1_outputs[8540] = ~(layer0_outputs[9111]);
    assign layer1_outputs[8541] = ~((layer0_outputs[4538]) ^ (layer0_outputs[750]));
    assign layer1_outputs[8542] = layer0_outputs[9524];
    assign layer1_outputs[8543] = layer0_outputs[7876];
    assign layer1_outputs[8544] = ~(layer0_outputs[2189]);
    assign layer1_outputs[8545] = layer0_outputs[2084];
    assign layer1_outputs[8546] = layer0_outputs[3358];
    assign layer1_outputs[8547] = ~(layer0_outputs[2984]);
    assign layer1_outputs[8548] = (layer0_outputs[3750]) & ~(layer0_outputs[12359]);
    assign layer1_outputs[8549] = ~(layer0_outputs[1536]);
    assign layer1_outputs[8550] = (layer0_outputs[7870]) & ~(layer0_outputs[129]);
    assign layer1_outputs[8551] = ~((layer0_outputs[11620]) | (layer0_outputs[8273]));
    assign layer1_outputs[8552] = ~(layer0_outputs[1148]);
    assign layer1_outputs[8553] = ~(layer0_outputs[4085]) | (layer0_outputs[7787]);
    assign layer1_outputs[8554] = ~((layer0_outputs[8126]) & (layer0_outputs[10302]));
    assign layer1_outputs[8555] = layer0_outputs[7634];
    assign layer1_outputs[8556] = ~((layer0_outputs[5894]) ^ (layer0_outputs[10549]));
    assign layer1_outputs[8557] = (layer0_outputs[6068]) & ~(layer0_outputs[4433]);
    assign layer1_outputs[8558] = ~(layer0_outputs[1167]);
    assign layer1_outputs[8559] = (layer0_outputs[6632]) ^ (layer0_outputs[10488]);
    assign layer1_outputs[8560] = (layer0_outputs[6485]) & (layer0_outputs[463]);
    assign layer1_outputs[8561] = ~(layer0_outputs[8345]);
    assign layer1_outputs[8562] = (layer0_outputs[12248]) & ~(layer0_outputs[4696]);
    assign layer1_outputs[8563] = ~(layer0_outputs[10504]);
    assign layer1_outputs[8564] = ~((layer0_outputs[4794]) & (layer0_outputs[9008]));
    assign layer1_outputs[8565] = layer0_outputs[2347];
    assign layer1_outputs[8566] = layer0_outputs[10520];
    assign layer1_outputs[8567] = ~(layer0_outputs[6166]) | (layer0_outputs[1357]);
    assign layer1_outputs[8568] = ~(layer0_outputs[8229]);
    assign layer1_outputs[8569] = ~(layer0_outputs[9213]) | (layer0_outputs[2889]);
    assign layer1_outputs[8570] = ~(layer0_outputs[2199]);
    assign layer1_outputs[8571] = ~((layer0_outputs[9994]) & (layer0_outputs[8291]));
    assign layer1_outputs[8572] = ~(layer0_outputs[2452]);
    assign layer1_outputs[8573] = ~(layer0_outputs[11156]);
    assign layer1_outputs[8574] = ~(layer0_outputs[11365]) | (layer0_outputs[175]);
    assign layer1_outputs[8575] = layer0_outputs[11817];
    assign layer1_outputs[8576] = layer0_outputs[9926];
    assign layer1_outputs[8577] = ~(layer0_outputs[7503]);
    assign layer1_outputs[8578] = ~((layer0_outputs[1601]) | (layer0_outputs[286]));
    assign layer1_outputs[8579] = (layer0_outputs[2259]) | (layer0_outputs[12010]);
    assign layer1_outputs[8580] = layer0_outputs[1252];
    assign layer1_outputs[8581] = layer0_outputs[6838];
    assign layer1_outputs[8582] = (layer0_outputs[12323]) ^ (layer0_outputs[339]);
    assign layer1_outputs[8583] = ~(layer0_outputs[638]);
    assign layer1_outputs[8584] = (layer0_outputs[8218]) & (layer0_outputs[1598]);
    assign layer1_outputs[8585] = ~((layer0_outputs[7262]) & (layer0_outputs[7164]));
    assign layer1_outputs[8586] = layer0_outputs[1816];
    assign layer1_outputs[8587] = ~(layer0_outputs[2943]) | (layer0_outputs[4001]);
    assign layer1_outputs[8588] = (layer0_outputs[7002]) & (layer0_outputs[4432]);
    assign layer1_outputs[8589] = ~(layer0_outputs[7583]);
    assign layer1_outputs[8590] = ~((layer0_outputs[5800]) ^ (layer0_outputs[240]));
    assign layer1_outputs[8591] = ~(layer0_outputs[8627]);
    assign layer1_outputs[8592] = ~(layer0_outputs[8542]);
    assign layer1_outputs[8593] = ~(layer0_outputs[10227]) | (layer0_outputs[11373]);
    assign layer1_outputs[8594] = ~(layer0_outputs[9100]) | (layer0_outputs[6763]);
    assign layer1_outputs[8595] = ~(layer0_outputs[10357]);
    assign layer1_outputs[8596] = layer0_outputs[4068];
    assign layer1_outputs[8597] = 1'b1;
    assign layer1_outputs[8598] = (layer0_outputs[3575]) & ~(layer0_outputs[6024]);
    assign layer1_outputs[8599] = layer0_outputs[10290];
    assign layer1_outputs[8600] = ~(layer0_outputs[4665]) | (layer0_outputs[5544]);
    assign layer1_outputs[8601] = ~((layer0_outputs[7792]) & (layer0_outputs[7411]));
    assign layer1_outputs[8602] = ~(layer0_outputs[5193]) | (layer0_outputs[11537]);
    assign layer1_outputs[8603] = (layer0_outputs[4006]) ^ (layer0_outputs[3431]);
    assign layer1_outputs[8604] = layer0_outputs[9393];
    assign layer1_outputs[8605] = ~(layer0_outputs[8789]);
    assign layer1_outputs[8606] = layer0_outputs[4162];
    assign layer1_outputs[8607] = (layer0_outputs[4823]) & (layer0_outputs[234]);
    assign layer1_outputs[8608] = (layer0_outputs[8221]) & ~(layer0_outputs[3593]);
    assign layer1_outputs[8609] = (layer0_outputs[6607]) | (layer0_outputs[7609]);
    assign layer1_outputs[8610] = layer0_outputs[6310];
    assign layer1_outputs[8611] = ~(layer0_outputs[8781]);
    assign layer1_outputs[8612] = ~(layer0_outputs[1300]) | (layer0_outputs[7620]);
    assign layer1_outputs[8613] = ~(layer0_outputs[6474]);
    assign layer1_outputs[8614] = (layer0_outputs[11623]) ^ (layer0_outputs[11098]);
    assign layer1_outputs[8615] = (layer0_outputs[147]) ^ (layer0_outputs[1514]);
    assign layer1_outputs[8616] = (layer0_outputs[4297]) & (layer0_outputs[6186]);
    assign layer1_outputs[8617] = ~((layer0_outputs[731]) ^ (layer0_outputs[8048]));
    assign layer1_outputs[8618] = ~(layer0_outputs[9483]);
    assign layer1_outputs[8619] = layer0_outputs[10039];
    assign layer1_outputs[8620] = (layer0_outputs[12576]) & (layer0_outputs[8235]);
    assign layer1_outputs[8621] = layer0_outputs[2322];
    assign layer1_outputs[8622] = layer0_outputs[6366];
    assign layer1_outputs[8623] = ~(layer0_outputs[9484]) | (layer0_outputs[12257]);
    assign layer1_outputs[8624] = (layer0_outputs[12322]) & ~(layer0_outputs[3530]);
    assign layer1_outputs[8625] = (layer0_outputs[9839]) & ~(layer0_outputs[1249]);
    assign layer1_outputs[8626] = ~(layer0_outputs[558]) | (layer0_outputs[6911]);
    assign layer1_outputs[8627] = 1'b0;
    assign layer1_outputs[8628] = ~(layer0_outputs[12274]) | (layer0_outputs[5680]);
    assign layer1_outputs[8629] = (layer0_outputs[3062]) | (layer0_outputs[4302]);
    assign layer1_outputs[8630] = layer0_outputs[9117];
    assign layer1_outputs[8631] = ~((layer0_outputs[4713]) | (layer0_outputs[9101]));
    assign layer1_outputs[8632] = ~((layer0_outputs[7513]) & (layer0_outputs[2653]));
    assign layer1_outputs[8633] = ~(layer0_outputs[11601]) | (layer0_outputs[10618]);
    assign layer1_outputs[8634] = layer0_outputs[1204];
    assign layer1_outputs[8635] = ~((layer0_outputs[1228]) & (layer0_outputs[7107]));
    assign layer1_outputs[8636] = ~(layer0_outputs[5342]);
    assign layer1_outputs[8637] = ~(layer0_outputs[3881]);
    assign layer1_outputs[8638] = (layer0_outputs[8675]) ^ (layer0_outputs[920]);
    assign layer1_outputs[8639] = layer0_outputs[9606];
    assign layer1_outputs[8640] = (layer0_outputs[5669]) & ~(layer0_outputs[8309]);
    assign layer1_outputs[8641] = (layer0_outputs[10239]) & ~(layer0_outputs[12568]);
    assign layer1_outputs[8642] = ~(layer0_outputs[7937]);
    assign layer1_outputs[8643] = ~(layer0_outputs[5680]);
    assign layer1_outputs[8644] = ~(layer0_outputs[9293]) | (layer0_outputs[4267]);
    assign layer1_outputs[8645] = (layer0_outputs[4485]) & (layer0_outputs[1592]);
    assign layer1_outputs[8646] = ~(layer0_outputs[9825]);
    assign layer1_outputs[8647] = ~((layer0_outputs[10400]) ^ (layer0_outputs[4026]));
    assign layer1_outputs[8648] = ~(layer0_outputs[12340]) | (layer0_outputs[2123]);
    assign layer1_outputs[8649] = layer0_outputs[4697];
    assign layer1_outputs[8650] = layer0_outputs[11075];
    assign layer1_outputs[8651] = layer0_outputs[1739];
    assign layer1_outputs[8652] = layer0_outputs[7794];
    assign layer1_outputs[8653] = layer0_outputs[12533];
    assign layer1_outputs[8654] = ~((layer0_outputs[6780]) ^ (layer0_outputs[11096]));
    assign layer1_outputs[8655] = layer0_outputs[9804];
    assign layer1_outputs[8656] = ~(layer0_outputs[2799]) | (layer0_outputs[3746]);
    assign layer1_outputs[8657] = (layer0_outputs[4644]) & ~(layer0_outputs[4021]);
    assign layer1_outputs[8658] = layer0_outputs[5290];
    assign layer1_outputs[8659] = (layer0_outputs[3232]) & (layer0_outputs[4940]);
    assign layer1_outputs[8660] = (layer0_outputs[10401]) & (layer0_outputs[1005]);
    assign layer1_outputs[8661] = layer0_outputs[9538];
    assign layer1_outputs[8662] = layer0_outputs[243];
    assign layer1_outputs[8663] = layer0_outputs[2943];
    assign layer1_outputs[8664] = ~(layer0_outputs[12482]);
    assign layer1_outputs[8665] = layer0_outputs[6491];
    assign layer1_outputs[8666] = ~(layer0_outputs[6014]);
    assign layer1_outputs[8667] = (layer0_outputs[5842]) & ~(layer0_outputs[9000]);
    assign layer1_outputs[8668] = 1'b1;
    assign layer1_outputs[8669] = ~(layer0_outputs[2529]);
    assign layer1_outputs[8670] = (layer0_outputs[9848]) ^ (layer0_outputs[4168]);
    assign layer1_outputs[8671] = layer0_outputs[820];
    assign layer1_outputs[8672] = ~((layer0_outputs[2531]) & (layer0_outputs[3974]));
    assign layer1_outputs[8673] = (layer0_outputs[1825]) & (layer0_outputs[2393]);
    assign layer1_outputs[8674] = 1'b0;
    assign layer1_outputs[8675] = layer0_outputs[5663];
    assign layer1_outputs[8676] = (layer0_outputs[12067]) & ~(layer0_outputs[3658]);
    assign layer1_outputs[8677] = (layer0_outputs[5662]) & ~(layer0_outputs[179]);
    assign layer1_outputs[8678] = 1'b0;
    assign layer1_outputs[8679] = ~(layer0_outputs[10467]);
    assign layer1_outputs[8680] = ~(layer0_outputs[367]);
    assign layer1_outputs[8681] = ~(layer0_outputs[1007]) | (layer0_outputs[12192]);
    assign layer1_outputs[8682] = layer0_outputs[9854];
    assign layer1_outputs[8683] = ~(layer0_outputs[1893]) | (layer0_outputs[9678]);
    assign layer1_outputs[8684] = ~(layer0_outputs[928]) | (layer0_outputs[11497]);
    assign layer1_outputs[8685] = ~((layer0_outputs[6909]) | (layer0_outputs[4842]));
    assign layer1_outputs[8686] = ~(layer0_outputs[370]);
    assign layer1_outputs[8687] = (layer0_outputs[15]) ^ (layer0_outputs[6601]);
    assign layer1_outputs[8688] = ~(layer0_outputs[345]);
    assign layer1_outputs[8689] = ~((layer0_outputs[5095]) ^ (layer0_outputs[9218]));
    assign layer1_outputs[8690] = ~(layer0_outputs[6630]) | (layer0_outputs[10431]);
    assign layer1_outputs[8691] = layer0_outputs[11281];
    assign layer1_outputs[8692] = layer0_outputs[3380];
    assign layer1_outputs[8693] = ~(layer0_outputs[10337]) | (layer0_outputs[4363]);
    assign layer1_outputs[8694] = ~(layer0_outputs[9031]) | (layer0_outputs[3312]);
    assign layer1_outputs[8695] = layer0_outputs[12072];
    assign layer1_outputs[8696] = ~(layer0_outputs[6256]);
    assign layer1_outputs[8697] = (layer0_outputs[1811]) ^ (layer0_outputs[426]);
    assign layer1_outputs[8698] = (layer0_outputs[10389]) ^ (layer0_outputs[6573]);
    assign layer1_outputs[8699] = layer0_outputs[6120];
    assign layer1_outputs[8700] = (layer0_outputs[8818]) | (layer0_outputs[3508]);
    assign layer1_outputs[8701] = ~((layer0_outputs[6432]) | (layer0_outputs[1972]));
    assign layer1_outputs[8702] = layer0_outputs[2242];
    assign layer1_outputs[8703] = layer0_outputs[3476];
    assign layer1_outputs[8704] = ~(layer0_outputs[3044]);
    assign layer1_outputs[8705] = ~(layer0_outputs[3479]);
    assign layer1_outputs[8706] = (layer0_outputs[5140]) & (layer0_outputs[474]);
    assign layer1_outputs[8707] = layer0_outputs[1177];
    assign layer1_outputs[8708] = ~(layer0_outputs[5004]);
    assign layer1_outputs[8709] = ~(layer0_outputs[4926]) | (layer0_outputs[7861]);
    assign layer1_outputs[8710] = (layer0_outputs[7510]) | (layer0_outputs[7960]);
    assign layer1_outputs[8711] = (layer0_outputs[6286]) & (layer0_outputs[2893]);
    assign layer1_outputs[8712] = ~((layer0_outputs[9080]) & (layer0_outputs[8474]));
    assign layer1_outputs[8713] = ~(layer0_outputs[9985]);
    assign layer1_outputs[8714] = ~((layer0_outputs[10372]) ^ (layer0_outputs[2923]));
    assign layer1_outputs[8715] = ~(layer0_outputs[4209]);
    assign layer1_outputs[8716] = (layer0_outputs[11489]) & ~(layer0_outputs[3477]);
    assign layer1_outputs[8717] = layer0_outputs[3232];
    assign layer1_outputs[8718] = ~(layer0_outputs[2574]) | (layer0_outputs[4339]);
    assign layer1_outputs[8719] = ~(layer0_outputs[1638]);
    assign layer1_outputs[8720] = ~((layer0_outputs[5280]) | (layer0_outputs[8582]));
    assign layer1_outputs[8721] = ~(layer0_outputs[11006]);
    assign layer1_outputs[8722] = layer0_outputs[6996];
    assign layer1_outputs[8723] = (layer0_outputs[4088]) | (layer0_outputs[8025]);
    assign layer1_outputs[8724] = ~(layer0_outputs[8391]);
    assign layer1_outputs[8725] = (layer0_outputs[262]) & ~(layer0_outputs[5296]);
    assign layer1_outputs[8726] = layer0_outputs[8406];
    assign layer1_outputs[8727] = (layer0_outputs[10343]) & ~(layer0_outputs[3875]);
    assign layer1_outputs[8728] = layer0_outputs[11430];
    assign layer1_outputs[8729] = ~(layer0_outputs[7940]);
    assign layer1_outputs[8730] = ~((layer0_outputs[7373]) ^ (layer0_outputs[12045]));
    assign layer1_outputs[8731] = ~(layer0_outputs[8009]) | (layer0_outputs[10840]);
    assign layer1_outputs[8732] = ~(layer0_outputs[2005]);
    assign layer1_outputs[8733] = ~(layer0_outputs[3019]);
    assign layer1_outputs[8734] = (layer0_outputs[627]) & ~(layer0_outputs[4500]);
    assign layer1_outputs[8735] = ~(layer0_outputs[4911]);
    assign layer1_outputs[8736] = layer0_outputs[5610];
    assign layer1_outputs[8737] = (layer0_outputs[3295]) | (layer0_outputs[8202]);
    assign layer1_outputs[8738] = ~((layer0_outputs[583]) ^ (layer0_outputs[9960]));
    assign layer1_outputs[8739] = layer0_outputs[6211];
    assign layer1_outputs[8740] = 1'b1;
    assign layer1_outputs[8741] = layer0_outputs[11647];
    assign layer1_outputs[8742] = ~(layer0_outputs[7036]) | (layer0_outputs[11947]);
    assign layer1_outputs[8743] = ~((layer0_outputs[9676]) & (layer0_outputs[1126]));
    assign layer1_outputs[8744] = ~(layer0_outputs[6036]);
    assign layer1_outputs[8745] = ~(layer0_outputs[9421]);
    assign layer1_outputs[8746] = ~((layer0_outputs[11452]) & (layer0_outputs[10803]));
    assign layer1_outputs[8747] = layer0_outputs[9256];
    assign layer1_outputs[8748] = (layer0_outputs[11958]) & (layer0_outputs[6057]);
    assign layer1_outputs[8749] = ~((layer0_outputs[8427]) | (layer0_outputs[9137]));
    assign layer1_outputs[8750] = ~(layer0_outputs[6086]);
    assign layer1_outputs[8751] = (layer0_outputs[11534]) & (layer0_outputs[696]);
    assign layer1_outputs[8752] = 1'b0;
    assign layer1_outputs[8753] = ~(layer0_outputs[6584]);
    assign layer1_outputs[8754] = ~(layer0_outputs[226]);
    assign layer1_outputs[8755] = ~((layer0_outputs[1555]) | (layer0_outputs[1490]));
    assign layer1_outputs[8756] = ~((layer0_outputs[12380]) & (layer0_outputs[5442]));
    assign layer1_outputs[8757] = layer0_outputs[959];
    assign layer1_outputs[8758] = (layer0_outputs[3482]) | (layer0_outputs[5100]);
    assign layer1_outputs[8759] = (layer0_outputs[5497]) | (layer0_outputs[4932]);
    assign layer1_outputs[8760] = layer0_outputs[7868];
    assign layer1_outputs[8761] = ~(layer0_outputs[1975]);
    assign layer1_outputs[8762] = ~(layer0_outputs[5145]) | (layer0_outputs[6961]);
    assign layer1_outputs[8763] = (layer0_outputs[10335]) & (layer0_outputs[508]);
    assign layer1_outputs[8764] = layer0_outputs[12191];
    assign layer1_outputs[8765] = ~(layer0_outputs[8707]);
    assign layer1_outputs[8766] = ~(layer0_outputs[11092]);
    assign layer1_outputs[8767] = 1'b0;
    assign layer1_outputs[8768] = (layer0_outputs[12218]) & ~(layer0_outputs[1055]);
    assign layer1_outputs[8769] = ~((layer0_outputs[2819]) | (layer0_outputs[6354]));
    assign layer1_outputs[8770] = layer0_outputs[5376];
    assign layer1_outputs[8771] = ~(layer0_outputs[7483]);
    assign layer1_outputs[8772] = (layer0_outputs[8496]) & ~(layer0_outputs[3268]);
    assign layer1_outputs[8773] = layer0_outputs[1659];
    assign layer1_outputs[8774] = ~(layer0_outputs[1417]) | (layer0_outputs[12002]);
    assign layer1_outputs[8775] = (layer0_outputs[2868]) ^ (layer0_outputs[9371]);
    assign layer1_outputs[8776] = ~((layer0_outputs[7665]) | (layer0_outputs[10323]));
    assign layer1_outputs[8777] = (layer0_outputs[10586]) | (layer0_outputs[3250]);
    assign layer1_outputs[8778] = ~((layer0_outputs[7687]) & (layer0_outputs[356]));
    assign layer1_outputs[8779] = (layer0_outputs[1732]) & ~(layer0_outputs[8958]);
    assign layer1_outputs[8780] = (layer0_outputs[6126]) & (layer0_outputs[8292]);
    assign layer1_outputs[8781] = (layer0_outputs[2897]) & (layer0_outputs[10438]);
    assign layer1_outputs[8782] = (layer0_outputs[10595]) | (layer0_outputs[2954]);
    assign layer1_outputs[8783] = ~((layer0_outputs[283]) | (layer0_outputs[4503]));
    assign layer1_outputs[8784] = (layer0_outputs[2077]) & ~(layer0_outputs[5024]);
    assign layer1_outputs[8785] = ~((layer0_outputs[11103]) ^ (layer0_outputs[11599]));
    assign layer1_outputs[8786] = ~(layer0_outputs[4811]) | (layer0_outputs[2966]);
    assign layer1_outputs[8787] = (layer0_outputs[8925]) & (layer0_outputs[4542]);
    assign layer1_outputs[8788] = 1'b1;
    assign layer1_outputs[8789] = (layer0_outputs[3554]) ^ (layer0_outputs[4580]);
    assign layer1_outputs[8790] = ~(layer0_outputs[2785]);
    assign layer1_outputs[8791] = ~(layer0_outputs[1486]) | (layer0_outputs[8243]);
    assign layer1_outputs[8792] = ~((layer0_outputs[4093]) ^ (layer0_outputs[1687]));
    assign layer1_outputs[8793] = ~((layer0_outputs[5186]) & (layer0_outputs[10654]));
    assign layer1_outputs[8794] = ~(layer0_outputs[4022]);
    assign layer1_outputs[8795] = 1'b0;
    assign layer1_outputs[8796] = ~(layer0_outputs[6532]) | (layer0_outputs[3530]);
    assign layer1_outputs[8797] = ~((layer0_outputs[374]) ^ (layer0_outputs[10015]));
    assign layer1_outputs[8798] = ~(layer0_outputs[3500]) | (layer0_outputs[6306]);
    assign layer1_outputs[8799] = ~(layer0_outputs[3650]) | (layer0_outputs[4578]);
    assign layer1_outputs[8800] = ~((layer0_outputs[5018]) & (layer0_outputs[7313]));
    assign layer1_outputs[8801] = ~(layer0_outputs[5917]);
    assign layer1_outputs[8802] = (layer0_outputs[3197]) & (layer0_outputs[5739]);
    assign layer1_outputs[8803] = ~((layer0_outputs[1388]) ^ (layer0_outputs[8043]));
    assign layer1_outputs[8804] = ~(layer0_outputs[9785]);
    assign layer1_outputs[8805] = layer0_outputs[12741];
    assign layer1_outputs[8806] = (layer0_outputs[7949]) ^ (layer0_outputs[1697]);
    assign layer1_outputs[8807] = (layer0_outputs[3129]) & ~(layer0_outputs[4632]);
    assign layer1_outputs[8808] = (layer0_outputs[5400]) | (layer0_outputs[10013]);
    assign layer1_outputs[8809] = (layer0_outputs[12547]) | (layer0_outputs[1006]);
    assign layer1_outputs[8810] = ~(layer0_outputs[2079]) | (layer0_outputs[4687]);
    assign layer1_outputs[8811] = (layer0_outputs[8339]) & ~(layer0_outputs[1705]);
    assign layer1_outputs[8812] = ~(layer0_outputs[3945]);
    assign layer1_outputs[8813] = ~((layer0_outputs[3634]) ^ (layer0_outputs[5338]));
    assign layer1_outputs[8814] = layer0_outputs[9997];
    assign layer1_outputs[8815] = (layer0_outputs[7290]) | (layer0_outputs[12368]);
    assign layer1_outputs[8816] = layer0_outputs[7835];
    assign layer1_outputs[8817] = ~((layer0_outputs[2472]) | (layer0_outputs[10744]));
    assign layer1_outputs[8818] = ~((layer0_outputs[1700]) | (layer0_outputs[704]));
    assign layer1_outputs[8819] = (layer0_outputs[3465]) | (layer0_outputs[5075]);
    assign layer1_outputs[8820] = ~((layer0_outputs[12506]) ^ (layer0_outputs[5943]));
    assign layer1_outputs[8821] = ~((layer0_outputs[7766]) ^ (layer0_outputs[8390]));
    assign layer1_outputs[8822] = (layer0_outputs[7812]) & ~(layer0_outputs[10908]);
    assign layer1_outputs[8823] = ~((layer0_outputs[1513]) & (layer0_outputs[6745]));
    assign layer1_outputs[8824] = ~(layer0_outputs[6569]);
    assign layer1_outputs[8825] = ~(layer0_outputs[4360]) | (layer0_outputs[3286]);
    assign layer1_outputs[8826] = layer0_outputs[3785];
    assign layer1_outputs[8827] = (layer0_outputs[1261]) & (layer0_outputs[2126]);
    assign layer1_outputs[8828] = ~((layer0_outputs[7753]) ^ (layer0_outputs[7484]));
    assign layer1_outputs[8829] = ~(layer0_outputs[6200]);
    assign layer1_outputs[8830] = ~(layer0_outputs[11166]);
    assign layer1_outputs[8831] = ~(layer0_outputs[5890]) | (layer0_outputs[12065]);
    assign layer1_outputs[8832] = layer0_outputs[8947];
    assign layer1_outputs[8833] = 1'b1;
    assign layer1_outputs[8834] = ~(layer0_outputs[8244]);
    assign layer1_outputs[8835] = (layer0_outputs[2217]) | (layer0_outputs[261]);
    assign layer1_outputs[8836] = (layer0_outputs[7884]) & ~(layer0_outputs[12240]);
    assign layer1_outputs[8837] = ~(layer0_outputs[7733]) | (layer0_outputs[10366]);
    assign layer1_outputs[8838] = (layer0_outputs[2454]) & ~(layer0_outputs[10752]);
    assign layer1_outputs[8839] = ~((layer0_outputs[8612]) ^ (layer0_outputs[10150]));
    assign layer1_outputs[8840] = 1'b0;
    assign layer1_outputs[8841] = layer0_outputs[8931];
    assign layer1_outputs[8842] = ~(layer0_outputs[6969]);
    assign layer1_outputs[8843] = ~(layer0_outputs[10097]) | (layer0_outputs[5671]);
    assign layer1_outputs[8844] = layer0_outputs[445];
    assign layer1_outputs[8845] = layer0_outputs[9223];
    assign layer1_outputs[8846] = (layer0_outputs[12224]) & ~(layer0_outputs[11498]);
    assign layer1_outputs[8847] = ~(layer0_outputs[5530]);
    assign layer1_outputs[8848] = ~(layer0_outputs[606]);
    assign layer1_outputs[8849] = ~(layer0_outputs[1427]) | (layer0_outputs[2706]);
    assign layer1_outputs[8850] = ~((layer0_outputs[9192]) & (layer0_outputs[7192]));
    assign layer1_outputs[8851] = ~((layer0_outputs[1920]) ^ (layer0_outputs[968]));
    assign layer1_outputs[8852] = (layer0_outputs[10229]) & ~(layer0_outputs[4641]);
    assign layer1_outputs[8853] = (layer0_outputs[3711]) & ~(layer0_outputs[3167]);
    assign layer1_outputs[8854] = ~(layer0_outputs[10031]) | (layer0_outputs[8076]);
    assign layer1_outputs[8855] = ~(layer0_outputs[184]);
    assign layer1_outputs[8856] = ~(layer0_outputs[5004]);
    assign layer1_outputs[8857] = (layer0_outputs[3748]) & ~(layer0_outputs[7638]);
    assign layer1_outputs[8858] = (layer0_outputs[10660]) & (layer0_outputs[10891]);
    assign layer1_outputs[8859] = layer0_outputs[7584];
    assign layer1_outputs[8860] = ~(layer0_outputs[5939]);
    assign layer1_outputs[8861] = (layer0_outputs[1624]) | (layer0_outputs[778]);
    assign layer1_outputs[8862] = (layer0_outputs[568]) & (layer0_outputs[12483]);
    assign layer1_outputs[8863] = ~(layer0_outputs[9242]) | (layer0_outputs[7044]);
    assign layer1_outputs[8864] = (layer0_outputs[523]) & ~(layer0_outputs[6346]);
    assign layer1_outputs[8865] = ~(layer0_outputs[11567]);
    assign layer1_outputs[8866] = ~(layer0_outputs[12397]);
    assign layer1_outputs[8867] = (layer0_outputs[2347]) & (layer0_outputs[3760]);
    assign layer1_outputs[8868] = ~((layer0_outputs[7979]) | (layer0_outputs[502]));
    assign layer1_outputs[8869] = (layer0_outputs[5523]) & ~(layer0_outputs[5099]);
    assign layer1_outputs[8870] = (layer0_outputs[4709]) & ~(layer0_outputs[9522]);
    assign layer1_outputs[8871] = 1'b0;
    assign layer1_outputs[8872] = (layer0_outputs[1895]) & ~(layer0_outputs[9666]);
    assign layer1_outputs[8873] = layer0_outputs[11602];
    assign layer1_outputs[8874] = (layer0_outputs[6450]) & ~(layer0_outputs[5345]);
    assign layer1_outputs[8875] = 1'b0;
    assign layer1_outputs[8876] = layer0_outputs[817];
    assign layer1_outputs[8877] = layer0_outputs[5187];
    assign layer1_outputs[8878] = ~(layer0_outputs[10976]);
    assign layer1_outputs[8879] = ~((layer0_outputs[79]) & (layer0_outputs[7380]));
    assign layer1_outputs[8880] = ~((layer0_outputs[1312]) & (layer0_outputs[5126]));
    assign layer1_outputs[8881] = (layer0_outputs[3674]) & ~(layer0_outputs[4769]);
    assign layer1_outputs[8882] = ~(layer0_outputs[8011]) | (layer0_outputs[12602]);
    assign layer1_outputs[8883] = ~(layer0_outputs[4174]);
    assign layer1_outputs[8884] = ~(layer0_outputs[6312]);
    assign layer1_outputs[8885] = (layer0_outputs[4525]) & ~(layer0_outputs[7872]);
    assign layer1_outputs[8886] = 1'b1;
    assign layer1_outputs[8887] = ~(layer0_outputs[3325]);
    assign layer1_outputs[8888] = ~((layer0_outputs[119]) ^ (layer0_outputs[6948]));
    assign layer1_outputs[8889] = 1'b1;
    assign layer1_outputs[8890] = ~(layer0_outputs[7555]) | (layer0_outputs[2958]);
    assign layer1_outputs[8891] = (layer0_outputs[7581]) & ~(layer0_outputs[9743]);
    assign layer1_outputs[8892] = ~(layer0_outputs[10084]) | (layer0_outputs[4119]);
    assign layer1_outputs[8893] = (layer0_outputs[7131]) & ~(layer0_outputs[5332]);
    assign layer1_outputs[8894] = (layer0_outputs[11892]) & ~(layer0_outputs[11744]);
    assign layer1_outputs[8895] = layer0_outputs[3152];
    assign layer1_outputs[8896] = 1'b0;
    assign layer1_outputs[8897] = (layer0_outputs[7005]) & ~(layer0_outputs[11576]);
    assign layer1_outputs[8898] = 1'b0;
    assign layer1_outputs[8899] = ~(layer0_outputs[11671]);
    assign layer1_outputs[8900] = ~(layer0_outputs[2676]);
    assign layer1_outputs[8901] = (layer0_outputs[6923]) & ~(layer0_outputs[1305]);
    assign layer1_outputs[8902] = layer0_outputs[11216];
    assign layer1_outputs[8903] = (layer0_outputs[11766]) | (layer0_outputs[9105]);
    assign layer1_outputs[8904] = ~(layer0_outputs[11931]) | (layer0_outputs[9245]);
    assign layer1_outputs[8905] = layer0_outputs[5337];
    assign layer1_outputs[8906] = 1'b1;
    assign layer1_outputs[8907] = ~(layer0_outputs[12487]);
    assign layer1_outputs[8908] = ~(layer0_outputs[8445]) | (layer0_outputs[2209]);
    assign layer1_outputs[8909] = layer0_outputs[1338];
    assign layer1_outputs[8910] = 1'b0;
    assign layer1_outputs[8911] = ~(layer0_outputs[9404]) | (layer0_outputs[11127]);
    assign layer1_outputs[8912] = (layer0_outputs[8058]) & (layer0_outputs[1386]);
    assign layer1_outputs[8913] = ~(layer0_outputs[7565]) | (layer0_outputs[3948]);
    assign layer1_outputs[8914] = ~(layer0_outputs[847]);
    assign layer1_outputs[8915] = ~(layer0_outputs[4126]);
    assign layer1_outputs[8916] = ~(layer0_outputs[4701]);
    assign layer1_outputs[8917] = ~((layer0_outputs[2683]) & (layer0_outputs[4233]));
    assign layer1_outputs[8918] = ~((layer0_outputs[5265]) & (layer0_outputs[12370]));
    assign layer1_outputs[8919] = layer0_outputs[8412];
    assign layer1_outputs[8920] = layer0_outputs[2018];
    assign layer1_outputs[8921] = (layer0_outputs[6937]) ^ (layer0_outputs[3475]);
    assign layer1_outputs[8922] = ~(layer0_outputs[3580]);
    assign layer1_outputs[8923] = layer0_outputs[124];
    assign layer1_outputs[8924] = layer0_outputs[8852];
    assign layer1_outputs[8925] = (layer0_outputs[11021]) & ~(layer0_outputs[7481]);
    assign layer1_outputs[8926] = ~((layer0_outputs[2257]) & (layer0_outputs[4621]));
    assign layer1_outputs[8927] = (layer0_outputs[5807]) & ~(layer0_outputs[3830]);
    assign layer1_outputs[8928] = (layer0_outputs[11713]) | (layer0_outputs[8148]);
    assign layer1_outputs[8929] = (layer0_outputs[1323]) & (layer0_outputs[10083]);
    assign layer1_outputs[8930] = ~(layer0_outputs[2841]) | (layer0_outputs[1878]);
    assign layer1_outputs[8931] = (layer0_outputs[975]) ^ (layer0_outputs[8079]);
    assign layer1_outputs[8932] = ~(layer0_outputs[7220]);
    assign layer1_outputs[8933] = ~((layer0_outputs[3329]) | (layer0_outputs[6271]));
    assign layer1_outputs[8934] = layer0_outputs[12623];
    assign layer1_outputs[8935] = (layer0_outputs[12138]) | (layer0_outputs[11201]);
    assign layer1_outputs[8936] = (layer0_outputs[246]) & ~(layer0_outputs[2323]);
    assign layer1_outputs[8937] = (layer0_outputs[4721]) & ~(layer0_outputs[3937]);
    assign layer1_outputs[8938] = (layer0_outputs[10291]) | (layer0_outputs[5765]);
    assign layer1_outputs[8939] = ~(layer0_outputs[1492]) | (layer0_outputs[2099]);
    assign layer1_outputs[8940] = (layer0_outputs[5346]) ^ (layer0_outputs[7600]);
    assign layer1_outputs[8941] = ~((layer0_outputs[2147]) & (layer0_outputs[4799]));
    assign layer1_outputs[8942] = ~(layer0_outputs[9597]) | (layer0_outputs[7710]);
    assign layer1_outputs[8943] = ~(layer0_outputs[3706]);
    assign layer1_outputs[8944] = 1'b0;
    assign layer1_outputs[8945] = layer0_outputs[2354];
    assign layer1_outputs[8946] = ~(layer0_outputs[8660]) | (layer0_outputs[9246]);
    assign layer1_outputs[8947] = ~(layer0_outputs[11715]) | (layer0_outputs[10816]);
    assign layer1_outputs[8948] = (layer0_outputs[1995]) | (layer0_outputs[4712]);
    assign layer1_outputs[8949] = ~((layer0_outputs[6062]) ^ (layer0_outputs[8833]));
    assign layer1_outputs[8950] = (layer0_outputs[8471]) & ~(layer0_outputs[10258]);
    assign layer1_outputs[8951] = ~(layer0_outputs[4113]);
    assign layer1_outputs[8952] = layer0_outputs[7506];
    assign layer1_outputs[8953] = ~(layer0_outputs[2428]) | (layer0_outputs[10723]);
    assign layer1_outputs[8954] = ~(layer0_outputs[7362]);
    assign layer1_outputs[8955] = layer0_outputs[11034];
    assign layer1_outputs[8956] = ~((layer0_outputs[3617]) & (layer0_outputs[6078]));
    assign layer1_outputs[8957] = ~(layer0_outputs[4920]);
    assign layer1_outputs[8958] = ~(layer0_outputs[8530]);
    assign layer1_outputs[8959] = ~(layer0_outputs[2844]);
    assign layer1_outputs[8960] = ~((layer0_outputs[3125]) ^ (layer0_outputs[3968]));
    assign layer1_outputs[8961] = (layer0_outputs[1352]) & ~(layer0_outputs[4089]);
    assign layer1_outputs[8962] = ~((layer0_outputs[12336]) | (layer0_outputs[3080]));
    assign layer1_outputs[8963] = ~((layer0_outputs[4226]) & (layer0_outputs[7590]));
    assign layer1_outputs[8964] = ~(layer0_outputs[2931]) | (layer0_outputs[4218]);
    assign layer1_outputs[8965] = ~(layer0_outputs[12776]) | (layer0_outputs[6165]);
    assign layer1_outputs[8966] = ~(layer0_outputs[4335]) | (layer0_outputs[12329]);
    assign layer1_outputs[8967] = ~(layer0_outputs[1835]);
    assign layer1_outputs[8968] = layer0_outputs[12665];
    assign layer1_outputs[8969] = ~((layer0_outputs[8353]) | (layer0_outputs[4109]));
    assign layer1_outputs[8970] = (layer0_outputs[4051]) | (layer0_outputs[8017]);
    assign layer1_outputs[8971] = (layer0_outputs[4575]) | (layer0_outputs[11139]);
    assign layer1_outputs[8972] = (layer0_outputs[9450]) & (layer0_outputs[12011]);
    assign layer1_outputs[8973] = layer0_outputs[5654];
    assign layer1_outputs[8974] = layer0_outputs[5436];
    assign layer1_outputs[8975] = (layer0_outputs[3192]) & ~(layer0_outputs[6568]);
    assign layer1_outputs[8976] = layer0_outputs[10973];
    assign layer1_outputs[8977] = ~(layer0_outputs[9576]) | (layer0_outputs[2135]);
    assign layer1_outputs[8978] = ~((layer0_outputs[6329]) ^ (layer0_outputs[6052]));
    assign layer1_outputs[8979] = ~(layer0_outputs[11334]) | (layer0_outputs[2185]);
    assign layer1_outputs[8980] = ~((layer0_outputs[10058]) ^ (layer0_outputs[3447]));
    assign layer1_outputs[8981] = layer0_outputs[2035];
    assign layer1_outputs[8982] = 1'b0;
    assign layer1_outputs[8983] = (layer0_outputs[6998]) & ~(layer0_outputs[3631]);
    assign layer1_outputs[8984] = (layer0_outputs[7444]) | (layer0_outputs[2020]);
    assign layer1_outputs[8985] = (layer0_outputs[3437]) & ~(layer0_outputs[10861]);
    assign layer1_outputs[8986] = (layer0_outputs[2151]) | (layer0_outputs[4148]);
    assign layer1_outputs[8987] = (layer0_outputs[1422]) & ~(layer0_outputs[5957]);
    assign layer1_outputs[8988] = ~(layer0_outputs[474]) | (layer0_outputs[8161]);
    assign layer1_outputs[8989] = ~(layer0_outputs[11724]) | (layer0_outputs[3630]);
    assign layer1_outputs[8990] = (layer0_outputs[10080]) & ~(layer0_outputs[3184]);
    assign layer1_outputs[8991] = ~(layer0_outputs[12191]);
    assign layer1_outputs[8992] = 1'b0;
    assign layer1_outputs[8993] = ~(layer0_outputs[10288]);
    assign layer1_outputs[8994] = layer0_outputs[10686];
    assign layer1_outputs[8995] = ~((layer0_outputs[6525]) & (layer0_outputs[11857]));
    assign layer1_outputs[8996] = ~(layer0_outputs[1197]);
    assign layer1_outputs[8997] = ~((layer0_outputs[2877]) & (layer0_outputs[9770]));
    assign layer1_outputs[8998] = ~(layer0_outputs[4155]) | (layer0_outputs[1252]);
    assign layer1_outputs[8999] = layer0_outputs[2075];
    assign layer1_outputs[9000] = ~(layer0_outputs[9243]);
    assign layer1_outputs[9001] = ~(layer0_outputs[1983]);
    assign layer1_outputs[9002] = layer0_outputs[11474];
    assign layer1_outputs[9003] = (layer0_outputs[3218]) & ~(layer0_outputs[3091]);
    assign layer1_outputs[9004] = layer0_outputs[5353];
    assign layer1_outputs[9005] = ~(layer0_outputs[1071]) | (layer0_outputs[12029]);
    assign layer1_outputs[9006] = ~(layer0_outputs[4735]);
    assign layer1_outputs[9007] = ~((layer0_outputs[608]) & (layer0_outputs[8260]));
    assign layer1_outputs[9008] = ~(layer0_outputs[5258]);
    assign layer1_outputs[9009] = (layer0_outputs[3177]) ^ (layer0_outputs[9107]);
    assign layer1_outputs[9010] = layer0_outputs[6377];
    assign layer1_outputs[9011] = (layer0_outputs[5103]) & (layer0_outputs[9946]);
    assign layer1_outputs[9012] = (layer0_outputs[11009]) ^ (layer0_outputs[578]);
    assign layer1_outputs[9013] = (layer0_outputs[6056]) ^ (layer0_outputs[7040]);
    assign layer1_outputs[9014] = (layer0_outputs[3110]) & (layer0_outputs[12394]);
    assign layer1_outputs[9015] = ~(layer0_outputs[11225]);
    assign layer1_outputs[9016] = ~((layer0_outputs[8708]) ^ (layer0_outputs[8604]));
    assign layer1_outputs[9017] = (layer0_outputs[1106]) ^ (layer0_outputs[3301]);
    assign layer1_outputs[9018] = layer0_outputs[1612];
    assign layer1_outputs[9019] = 1'b1;
    assign layer1_outputs[9020] = (layer0_outputs[2422]) ^ (layer0_outputs[8928]);
    assign layer1_outputs[9021] = ~(layer0_outputs[4898]);
    assign layer1_outputs[9022] = ~((layer0_outputs[7271]) & (layer0_outputs[50]));
    assign layer1_outputs[9023] = (layer0_outputs[7120]) & ~(layer0_outputs[6270]);
    assign layer1_outputs[9024] = layer0_outputs[10155];
    assign layer1_outputs[9025] = ~(layer0_outputs[663]) | (layer0_outputs[12476]);
    assign layer1_outputs[9026] = ~(layer0_outputs[3041]);
    assign layer1_outputs[9027] = ~(layer0_outputs[7279]);
    assign layer1_outputs[9028] = ~((layer0_outputs[2410]) & (layer0_outputs[10786]));
    assign layer1_outputs[9029] = (layer0_outputs[2329]) & (layer0_outputs[8448]);
    assign layer1_outputs[9030] = ~((layer0_outputs[5678]) | (layer0_outputs[2465]));
    assign layer1_outputs[9031] = layer0_outputs[12702];
    assign layer1_outputs[9032] = ~(layer0_outputs[8849]);
    assign layer1_outputs[9033] = ~(layer0_outputs[5299]) | (layer0_outputs[3375]);
    assign layer1_outputs[9034] = layer0_outputs[6813];
    assign layer1_outputs[9035] = ~((layer0_outputs[5143]) | (layer0_outputs[11023]));
    assign layer1_outputs[9036] = ~((layer0_outputs[10169]) | (layer0_outputs[11585]));
    assign layer1_outputs[9037] = ~(layer0_outputs[9220]);
    assign layer1_outputs[9038] = (layer0_outputs[28]) | (layer0_outputs[5649]);
    assign layer1_outputs[9039] = (layer0_outputs[7592]) ^ (layer0_outputs[7564]);
    assign layer1_outputs[9040] = layer0_outputs[9874];
    assign layer1_outputs[9041] = ~(layer0_outputs[12280]);
    assign layer1_outputs[9042] = layer0_outputs[10313];
    assign layer1_outputs[9043] = 1'b0;
    assign layer1_outputs[9044] = layer0_outputs[10580];
    assign layer1_outputs[9045] = ~(layer0_outputs[200]);
    assign layer1_outputs[9046] = ~(layer0_outputs[8201]);
    assign layer1_outputs[9047] = (layer0_outputs[1400]) & ~(layer0_outputs[9896]);
    assign layer1_outputs[9048] = layer0_outputs[9457];
    assign layer1_outputs[9049] = ~((layer0_outputs[195]) & (layer0_outputs[10204]));
    assign layer1_outputs[9050] = ~(layer0_outputs[7601]);
    assign layer1_outputs[9051] = (layer0_outputs[1976]) & ~(layer0_outputs[8179]);
    assign layer1_outputs[9052] = ~((layer0_outputs[7977]) | (layer0_outputs[7920]));
    assign layer1_outputs[9053] = (layer0_outputs[1886]) & ~(layer0_outputs[4124]);
    assign layer1_outputs[9054] = ~(layer0_outputs[1868]);
    assign layer1_outputs[9055] = (layer0_outputs[535]) & ~(layer0_outputs[1959]);
    assign layer1_outputs[9056] = 1'b1;
    assign layer1_outputs[9057] = ~(layer0_outputs[2539]);
    assign layer1_outputs[9058] = ~(layer0_outputs[260]) | (layer0_outputs[1842]);
    assign layer1_outputs[9059] = (layer0_outputs[310]) & (layer0_outputs[2925]);
    assign layer1_outputs[9060] = (layer0_outputs[4987]) & ~(layer0_outputs[5087]);
    assign layer1_outputs[9061] = ~(layer0_outputs[4126]) | (layer0_outputs[9790]);
    assign layer1_outputs[9062] = (layer0_outputs[7384]) & ~(layer0_outputs[1540]);
    assign layer1_outputs[9063] = 1'b0;
    assign layer1_outputs[9064] = ~(layer0_outputs[9290]) | (layer0_outputs[9087]);
    assign layer1_outputs[9065] = layer0_outputs[1532];
    assign layer1_outputs[9066] = ~(layer0_outputs[7622]) | (layer0_outputs[4332]);
    assign layer1_outputs[9067] = ~((layer0_outputs[7299]) & (layer0_outputs[8449]));
    assign layer1_outputs[9068] = 1'b0;
    assign layer1_outputs[9069] = layer0_outputs[1787];
    assign layer1_outputs[9070] = layer0_outputs[1378];
    assign layer1_outputs[9071] = (layer0_outputs[6756]) | (layer0_outputs[11780]);
    assign layer1_outputs[9072] = layer0_outputs[2609];
    assign layer1_outputs[9073] = (layer0_outputs[9880]) & (layer0_outputs[10812]);
    assign layer1_outputs[9074] = layer0_outputs[5926];
    assign layer1_outputs[9075] = ~((layer0_outputs[2778]) | (layer0_outputs[817]));
    assign layer1_outputs[9076] = ~((layer0_outputs[9084]) & (layer0_outputs[2206]));
    assign layer1_outputs[9077] = layer0_outputs[5330];
    assign layer1_outputs[9078] = ~(layer0_outputs[8499]);
    assign layer1_outputs[9079] = ~(layer0_outputs[3969]);
    assign layer1_outputs[9080] = ~(layer0_outputs[10507]);
    assign layer1_outputs[9081] = ~(layer0_outputs[9276]);
    assign layer1_outputs[9082] = ~((layer0_outputs[2482]) & (layer0_outputs[12567]));
    assign layer1_outputs[9083] = ~(layer0_outputs[12418]);
    assign layer1_outputs[9084] = ~((layer0_outputs[4573]) ^ (layer0_outputs[4889]));
    assign layer1_outputs[9085] = layer0_outputs[3470];
    assign layer1_outputs[9086] = (layer0_outputs[11269]) | (layer0_outputs[6831]);
    assign layer1_outputs[9087] = ~(layer0_outputs[9669]);
    assign layer1_outputs[9088] = ~((layer0_outputs[3426]) ^ (layer0_outputs[1217]));
    assign layer1_outputs[9089] = (layer0_outputs[10233]) ^ (layer0_outputs[7359]);
    assign layer1_outputs[9090] = ~((layer0_outputs[7418]) ^ (layer0_outputs[3645]));
    assign layer1_outputs[9091] = (layer0_outputs[11122]) & (layer0_outputs[7080]);
    assign layer1_outputs[9092] = (layer0_outputs[2594]) & ~(layer0_outputs[11148]);
    assign layer1_outputs[9093] = ~(layer0_outputs[5793]);
    assign layer1_outputs[9094] = ~((layer0_outputs[11815]) & (layer0_outputs[11681]));
    assign layer1_outputs[9095] = (layer0_outputs[1179]) ^ (layer0_outputs[12490]);
    assign layer1_outputs[9096] = ~(layer0_outputs[3808]);
    assign layer1_outputs[9097] = layer0_outputs[1519];
    assign layer1_outputs[9098] = layer0_outputs[4600];
    assign layer1_outputs[9099] = (layer0_outputs[5459]) ^ (layer0_outputs[536]);
    assign layer1_outputs[9100] = layer0_outputs[3937];
    assign layer1_outputs[9101] = layer0_outputs[12448];
    assign layer1_outputs[9102] = (layer0_outputs[2915]) | (layer0_outputs[7880]);
    assign layer1_outputs[9103] = ~(layer0_outputs[2816]) | (layer0_outputs[5983]);
    assign layer1_outputs[9104] = ~(layer0_outputs[10493]);
    assign layer1_outputs[9105] = (layer0_outputs[3985]) & ~(layer0_outputs[11859]);
    assign layer1_outputs[9106] = ~((layer0_outputs[5255]) ^ (layer0_outputs[5424]));
    assign layer1_outputs[9107] = (layer0_outputs[9869]) & (layer0_outputs[3992]);
    assign layer1_outputs[9108] = ~((layer0_outputs[3770]) & (layer0_outputs[5321]));
    assign layer1_outputs[9109] = (layer0_outputs[6201]) & ~(layer0_outputs[522]);
    assign layer1_outputs[9110] = ~(layer0_outputs[10429]);
    assign layer1_outputs[9111] = (layer0_outputs[176]) | (layer0_outputs[5054]);
    assign layer1_outputs[9112] = ~((layer0_outputs[7674]) | (layer0_outputs[8844]));
    assign layer1_outputs[9113] = ~(layer0_outputs[2626]) | (layer0_outputs[12736]);
    assign layer1_outputs[9114] = ~(layer0_outputs[5267]) | (layer0_outputs[6725]);
    assign layer1_outputs[9115] = ~(layer0_outputs[12782]);
    assign layer1_outputs[9116] = ~((layer0_outputs[12740]) | (layer0_outputs[8044]));
    assign layer1_outputs[9117] = 1'b1;
    assign layer1_outputs[9118] = ~(layer0_outputs[12505]) | (layer0_outputs[2662]);
    assign layer1_outputs[9119] = ~(layer0_outputs[12345]);
    assign layer1_outputs[9120] = ~(layer0_outputs[11740]);
    assign layer1_outputs[9121] = layer0_outputs[4890];
    assign layer1_outputs[9122] = (layer0_outputs[10255]) & ~(layer0_outputs[6535]);
    assign layer1_outputs[9123] = (layer0_outputs[11596]) ^ (layer0_outputs[11716]);
    assign layer1_outputs[9124] = ~((layer0_outputs[12652]) | (layer0_outputs[10296]));
    assign layer1_outputs[9125] = ~((layer0_outputs[11226]) & (layer0_outputs[9547]));
    assign layer1_outputs[9126] = ~(layer0_outputs[9132]);
    assign layer1_outputs[9127] = ~(layer0_outputs[2996]);
    assign layer1_outputs[9128] = ~(layer0_outputs[9581]) | (layer0_outputs[12239]);
    assign layer1_outputs[9129] = (layer0_outputs[3778]) ^ (layer0_outputs[8498]);
    assign layer1_outputs[9130] = ~(layer0_outputs[378]);
    assign layer1_outputs[9131] = ~(layer0_outputs[4810]) | (layer0_outputs[3570]);
    assign layer1_outputs[9132] = ~((layer0_outputs[5690]) ^ (layer0_outputs[9177]));
    assign layer1_outputs[9133] = ~(layer0_outputs[4356]);
    assign layer1_outputs[9134] = (layer0_outputs[5389]) & ~(layer0_outputs[3939]);
    assign layer1_outputs[9135] = (layer0_outputs[9632]) & ~(layer0_outputs[2063]);
    assign layer1_outputs[9136] = (layer0_outputs[7382]) | (layer0_outputs[8354]);
    assign layer1_outputs[9137] = (layer0_outputs[10082]) & ~(layer0_outputs[3728]);
    assign layer1_outputs[9138] = ~(layer0_outputs[5557]);
    assign layer1_outputs[9139] = layer0_outputs[3980];
    assign layer1_outputs[9140] = ~(layer0_outputs[7456]);
    assign layer1_outputs[9141] = (layer0_outputs[4387]) & ~(layer0_outputs[6665]);
    assign layer1_outputs[9142] = (layer0_outputs[3360]) & (layer0_outputs[3542]);
    assign layer1_outputs[9143] = ~(layer0_outputs[7222]);
    assign layer1_outputs[9144] = (layer0_outputs[12747]) | (layer0_outputs[7072]);
    assign layer1_outputs[9145] = ~(layer0_outputs[3658]);
    assign layer1_outputs[9146] = ~(layer0_outputs[9020]);
    assign layer1_outputs[9147] = layer0_outputs[8519];
    assign layer1_outputs[9148] = ~((layer0_outputs[12282]) | (layer0_outputs[9237]));
    assign layer1_outputs[9149] = ~(layer0_outputs[2916]);
    assign layer1_outputs[9150] = (layer0_outputs[11797]) & (layer0_outputs[854]);
    assign layer1_outputs[9151] = ~(layer0_outputs[11995]) | (layer0_outputs[12130]);
    assign layer1_outputs[9152] = layer0_outputs[4250];
    assign layer1_outputs[9153] = ~((layer0_outputs[4943]) | (layer0_outputs[6067]));
    assign layer1_outputs[9154] = ~(layer0_outputs[4879]);
    assign layer1_outputs[9155] = ~((layer0_outputs[8429]) | (layer0_outputs[4798]));
    assign layer1_outputs[9156] = layer0_outputs[2156];
    assign layer1_outputs[9157] = ~(layer0_outputs[11691]);
    assign layer1_outputs[9158] = layer0_outputs[4594];
    assign layer1_outputs[9159] = layer0_outputs[7765];
    assign layer1_outputs[9160] = ~((layer0_outputs[8059]) | (layer0_outputs[2057]));
    assign layer1_outputs[9161] = ~(layer0_outputs[4237]);
    assign layer1_outputs[9162] = layer0_outputs[4461];
    assign layer1_outputs[9163] = layer0_outputs[12491];
    assign layer1_outputs[9164] = ~(layer0_outputs[4470]) | (layer0_outputs[12528]);
    assign layer1_outputs[9165] = ~((layer0_outputs[1843]) | (layer0_outputs[1768]));
    assign layer1_outputs[9166] = ~(layer0_outputs[1776]) | (layer0_outputs[980]);
    assign layer1_outputs[9167] = (layer0_outputs[10396]) ^ (layer0_outputs[7084]);
    assign layer1_outputs[9168] = ~(layer0_outputs[10494]);
    assign layer1_outputs[9169] = ~(layer0_outputs[7397]) | (layer0_outputs[8049]);
    assign layer1_outputs[9170] = 1'b0;
    assign layer1_outputs[9171] = (layer0_outputs[10282]) & (layer0_outputs[9670]);
    assign layer1_outputs[9172] = ~((layer0_outputs[3309]) & (layer0_outputs[9406]));
    assign layer1_outputs[9173] = 1'b0;
    assign layer1_outputs[9174] = ~(layer0_outputs[8021]) | (layer0_outputs[7792]);
    assign layer1_outputs[9175] = ~((layer0_outputs[4480]) ^ (layer0_outputs[5574]));
    assign layer1_outputs[9176] = ~(layer0_outputs[3538]);
    assign layer1_outputs[9177] = ~((layer0_outputs[11297]) ^ (layer0_outputs[9005]));
    assign layer1_outputs[9178] = ~(layer0_outputs[3453]);
    assign layer1_outputs[9179] = ~(layer0_outputs[9283]);
    assign layer1_outputs[9180] = ~(layer0_outputs[12491]) | (layer0_outputs[9677]);
    assign layer1_outputs[9181] = layer0_outputs[8670];
    assign layer1_outputs[9182] = layer0_outputs[1320];
    assign layer1_outputs[9183] = ~(layer0_outputs[6420]);
    assign layer1_outputs[9184] = (layer0_outputs[1306]) & (layer0_outputs[2610]);
    assign layer1_outputs[9185] = layer0_outputs[163];
    assign layer1_outputs[9186] = ~((layer0_outputs[6938]) | (layer0_outputs[6218]));
    assign layer1_outputs[9187] = (layer0_outputs[9716]) | (layer0_outputs[857]);
    assign layer1_outputs[9188] = ~(layer0_outputs[7030]) | (layer0_outputs[7909]);
    assign layer1_outputs[9189] = layer0_outputs[8233];
    assign layer1_outputs[9190] = ~(layer0_outputs[1971]);
    assign layer1_outputs[9191] = ~(layer0_outputs[6862]);
    assign layer1_outputs[9192] = layer0_outputs[2760];
    assign layer1_outputs[9193] = (layer0_outputs[827]) & ~(layer0_outputs[987]);
    assign layer1_outputs[9194] = ~((layer0_outputs[1270]) | (layer0_outputs[4295]));
    assign layer1_outputs[9195] = (layer0_outputs[1056]) & ~(layer0_outputs[6569]);
    assign layer1_outputs[9196] = 1'b1;
    assign layer1_outputs[9197] = (layer0_outputs[10722]) ^ (layer0_outputs[6411]);
    assign layer1_outputs[9198] = layer0_outputs[12489];
    assign layer1_outputs[9199] = (layer0_outputs[8153]) & ~(layer0_outputs[11355]);
    assign layer1_outputs[9200] = (layer0_outputs[2483]) & ~(layer0_outputs[1627]);
    assign layer1_outputs[9201] = layer0_outputs[1849];
    assign layer1_outputs[9202] = ~(layer0_outputs[6944]);
    assign layer1_outputs[9203] = layer0_outputs[8552];
    assign layer1_outputs[9204] = layer0_outputs[11706];
    assign layer1_outputs[9205] = layer0_outputs[2144];
    assign layer1_outputs[9206] = ~((layer0_outputs[8314]) | (layer0_outputs[9052]));
    assign layer1_outputs[9207] = layer0_outputs[4528];
    assign layer1_outputs[9208] = (layer0_outputs[4380]) & ~(layer0_outputs[1885]);
    assign layer1_outputs[9209] = ~(layer0_outputs[3951]) | (layer0_outputs[2758]);
    assign layer1_outputs[9210] = ~(layer0_outputs[4078]);
    assign layer1_outputs[9211] = ~(layer0_outputs[9288]);
    assign layer1_outputs[9212] = ~(layer0_outputs[1863]);
    assign layer1_outputs[9213] = ~((layer0_outputs[9449]) | (layer0_outputs[1979]));
    assign layer1_outputs[9214] = ~((layer0_outputs[9340]) ^ (layer0_outputs[4144]));
    assign layer1_outputs[9215] = ~(layer0_outputs[8156]) | (layer0_outputs[3024]);
    assign layer1_outputs[9216] = (layer0_outputs[11890]) & ~(layer0_outputs[11302]);
    assign layer1_outputs[9217] = (layer0_outputs[4894]) & (layer0_outputs[12307]);
    assign layer1_outputs[9218] = layer0_outputs[9831];
    assign layer1_outputs[9219] = layer0_outputs[7775];
    assign layer1_outputs[9220] = layer0_outputs[12772];
    assign layer1_outputs[9221] = ~(layer0_outputs[3392]) | (layer0_outputs[11903]);
    assign layer1_outputs[9222] = ~(layer0_outputs[1987]);
    assign layer1_outputs[9223] = (layer0_outputs[3441]) | (layer0_outputs[109]);
    assign layer1_outputs[9224] = ~(layer0_outputs[10388]) | (layer0_outputs[9472]);
    assign layer1_outputs[9225] = ~(layer0_outputs[11306]);
    assign layer1_outputs[9226] = layer0_outputs[11871];
    assign layer1_outputs[9227] = (layer0_outputs[12458]) & (layer0_outputs[1213]);
    assign layer1_outputs[9228] = (layer0_outputs[5052]) & ~(layer0_outputs[10884]);
    assign layer1_outputs[9229] = (layer0_outputs[7712]) & ~(layer0_outputs[9814]);
    assign layer1_outputs[9230] = ~((layer0_outputs[9317]) | (layer0_outputs[146]));
    assign layer1_outputs[9231] = layer0_outputs[6207];
    assign layer1_outputs[9232] = ~(layer0_outputs[7922]) | (layer0_outputs[4365]);
    assign layer1_outputs[9233] = (layer0_outputs[485]) | (layer0_outputs[2971]);
    assign layer1_outputs[9234] = (layer0_outputs[10106]) | (layer0_outputs[619]);
    assign layer1_outputs[9235] = layer0_outputs[10459];
    assign layer1_outputs[9236] = ~((layer0_outputs[7945]) & (layer0_outputs[11071]));
    assign layer1_outputs[9237] = (layer0_outputs[8341]) ^ (layer0_outputs[3520]);
    assign layer1_outputs[9238] = (layer0_outputs[3123]) & (layer0_outputs[8982]);
    assign layer1_outputs[9239] = layer0_outputs[10619];
    assign layer1_outputs[9240] = (layer0_outputs[8745]) | (layer0_outputs[93]);
    assign layer1_outputs[9241] = ~(layer0_outputs[8077]);
    assign layer1_outputs[9242] = layer0_outputs[1738];
    assign layer1_outputs[9243] = ~(layer0_outputs[6598]);
    assign layer1_outputs[9244] = (layer0_outputs[1325]) | (layer0_outputs[9680]);
    assign layer1_outputs[9245] = ~((layer0_outputs[9411]) | (layer0_outputs[8872]));
    assign layer1_outputs[9246] = layer0_outputs[8690];
    assign layer1_outputs[9247] = ~((layer0_outputs[336]) | (layer0_outputs[11639]));
    assign layer1_outputs[9248] = layer0_outputs[930];
    assign layer1_outputs[9249] = ~(layer0_outputs[6294]) | (layer0_outputs[7400]);
    assign layer1_outputs[9250] = ~((layer0_outputs[7100]) ^ (layer0_outputs[8425]));
    assign layer1_outputs[9251] = ~(layer0_outputs[9985]);
    assign layer1_outputs[9252] = layer0_outputs[8588];
    assign layer1_outputs[9253] = ~(layer0_outputs[3130]);
    assign layer1_outputs[9254] = (layer0_outputs[4309]) ^ (layer0_outputs[11899]);
    assign layer1_outputs[9255] = ~(layer0_outputs[8607]);
    assign layer1_outputs[9256] = ~((layer0_outputs[6620]) | (layer0_outputs[4814]));
    assign layer1_outputs[9257] = layer0_outputs[4297];
    assign layer1_outputs[9258] = ~((layer0_outputs[4344]) ^ (layer0_outputs[12175]));
    assign layer1_outputs[9259] = ~(layer0_outputs[1945]);
    assign layer1_outputs[9260] = (layer0_outputs[4652]) & ~(layer0_outputs[5078]);
    assign layer1_outputs[9261] = ~(layer0_outputs[3138]);
    assign layer1_outputs[9262] = (layer0_outputs[4069]) ^ (layer0_outputs[11562]);
    assign layer1_outputs[9263] = ~((layer0_outputs[5068]) & (layer0_outputs[6931]));
    assign layer1_outputs[9264] = ~(layer0_outputs[4241]);
    assign layer1_outputs[9265] = (layer0_outputs[11202]) | (layer0_outputs[409]);
    assign layer1_outputs[9266] = ~(layer0_outputs[4480]);
    assign layer1_outputs[9267] = layer0_outputs[8303];
    assign layer1_outputs[9268] = ~(layer0_outputs[205]) | (layer0_outputs[9063]);
    assign layer1_outputs[9269] = (layer0_outputs[9995]) & ~(layer0_outputs[7854]);
    assign layer1_outputs[9270] = ~(layer0_outputs[73]) | (layer0_outputs[48]);
    assign layer1_outputs[9271] = ~(layer0_outputs[852]);
    assign layer1_outputs[9272] = layer0_outputs[6264];
    assign layer1_outputs[9273] = ~(layer0_outputs[9702]) | (layer0_outputs[3292]);
    assign layer1_outputs[9274] = layer0_outputs[1621];
    assign layer1_outputs[9275] = (layer0_outputs[8767]) | (layer0_outputs[3175]);
    assign layer1_outputs[9276] = ~((layer0_outputs[10730]) ^ (layer0_outputs[6715]));
    assign layer1_outputs[9277] = layer0_outputs[11068];
    assign layer1_outputs[9278] = ~(layer0_outputs[487]);
    assign layer1_outputs[9279] = layer0_outputs[12610];
    assign layer1_outputs[9280] = ~(layer0_outputs[6332]);
    assign layer1_outputs[9281] = ~(layer0_outputs[997]) | (layer0_outputs[12710]);
    assign layer1_outputs[9282] = (layer0_outputs[2432]) & (layer0_outputs[5322]);
    assign layer1_outputs[9283] = ~((layer0_outputs[12664]) ^ (layer0_outputs[181]));
    assign layer1_outputs[9284] = ~(layer0_outputs[7871]) | (layer0_outputs[5918]);
    assign layer1_outputs[9285] = (layer0_outputs[9309]) & (layer0_outputs[143]);
    assign layer1_outputs[9286] = layer0_outputs[12701];
    assign layer1_outputs[9287] = ~(layer0_outputs[630]);
    assign layer1_outputs[9288] = ~((layer0_outputs[10963]) ^ (layer0_outputs[10230]));
    assign layer1_outputs[9289] = ~(layer0_outputs[2573]);
    assign layer1_outputs[9290] = ~(layer0_outputs[6516]);
    assign layer1_outputs[9291] = layer0_outputs[7672];
    assign layer1_outputs[9292] = ~(layer0_outputs[3855]);
    assign layer1_outputs[9293] = 1'b1;
    assign layer1_outputs[9294] = (layer0_outputs[10176]) & (layer0_outputs[2988]);
    assign layer1_outputs[9295] = (layer0_outputs[7938]) ^ (layer0_outputs[11765]);
    assign layer1_outputs[9296] = ~(layer0_outputs[11025]);
    assign layer1_outputs[9297] = ~(layer0_outputs[8191]) | (layer0_outputs[6013]);
    assign layer1_outputs[9298] = (layer0_outputs[4612]) ^ (layer0_outputs[224]);
    assign layer1_outputs[9299] = (layer0_outputs[186]) & ~(layer0_outputs[5954]);
    assign layer1_outputs[9300] = (layer0_outputs[3355]) ^ (layer0_outputs[10269]);
    assign layer1_outputs[9301] = ~(layer0_outputs[3417]);
    assign layer1_outputs[9302] = ~(layer0_outputs[8206]);
    assign layer1_outputs[9303] = ~(layer0_outputs[9091]) | (layer0_outputs[353]);
    assign layer1_outputs[9304] = ~(layer0_outputs[5786]);
    assign layer1_outputs[9305] = (layer0_outputs[6428]) & ~(layer0_outputs[6416]);
    assign layer1_outputs[9306] = (layer0_outputs[3514]) & (layer0_outputs[10892]);
    assign layer1_outputs[9307] = layer0_outputs[11128];
    assign layer1_outputs[9308] = layer0_outputs[9000];
    assign layer1_outputs[9309] = ~(layer0_outputs[10557]);
    assign layer1_outputs[9310] = ~(layer0_outputs[12510]);
    assign layer1_outputs[9311] = ~((layer0_outputs[4559]) | (layer0_outputs[8981]));
    assign layer1_outputs[9312] = ~(layer0_outputs[2873]);
    assign layer1_outputs[9313] = layer0_outputs[10522];
    assign layer1_outputs[9314] = ~(layer0_outputs[7520]);
    assign layer1_outputs[9315] = ~(layer0_outputs[6704]);
    assign layer1_outputs[9316] = (layer0_outputs[1471]) & ~(layer0_outputs[434]);
    assign layer1_outputs[9317] = ~(layer0_outputs[4397]) | (layer0_outputs[4506]);
    assign layer1_outputs[9318] = (layer0_outputs[10341]) & ~(layer0_outputs[1493]);
    assign layer1_outputs[9319] = (layer0_outputs[8591]) | (layer0_outputs[5124]);
    assign layer1_outputs[9320] = (layer0_outputs[8911]) & (layer0_outputs[821]);
    assign layer1_outputs[9321] = ~(layer0_outputs[11541]) | (layer0_outputs[10756]);
    assign layer1_outputs[9322] = (layer0_outputs[11895]) | (layer0_outputs[11013]);
    assign layer1_outputs[9323] = 1'b1;
    assign layer1_outputs[9324] = layer0_outputs[2941];
    assign layer1_outputs[9325] = 1'b0;
    assign layer1_outputs[9326] = (layer0_outputs[6564]) & (layer0_outputs[5841]);
    assign layer1_outputs[9327] = (layer0_outputs[8023]) ^ (layer0_outputs[1312]);
    assign layer1_outputs[9328] = layer0_outputs[12496];
    assign layer1_outputs[9329] = ~(layer0_outputs[7383]);
    assign layer1_outputs[9330] = ~(layer0_outputs[10426]);
    assign layer1_outputs[9331] = (layer0_outputs[526]) | (layer0_outputs[6125]);
    assign layer1_outputs[9332] = ~((layer0_outputs[7751]) & (layer0_outputs[3118]));
    assign layer1_outputs[9333] = (layer0_outputs[4083]) & ~(layer0_outputs[8685]);
    assign layer1_outputs[9334] = layer0_outputs[12];
    assign layer1_outputs[9335] = (layer0_outputs[2043]) & ~(layer0_outputs[8198]);
    assign layer1_outputs[9336] = (layer0_outputs[2538]) & (layer0_outputs[9679]);
    assign layer1_outputs[9337] = ~(layer0_outputs[3261]) | (layer0_outputs[12393]);
    assign layer1_outputs[9338] = layer0_outputs[2325];
    assign layer1_outputs[9339] = ~(layer0_outputs[856]) | (layer0_outputs[12756]);
    assign layer1_outputs[9340] = ~(layer0_outputs[8996]);
    assign layer1_outputs[9341] = ~((layer0_outputs[3183]) ^ (layer0_outputs[4649]));
    assign layer1_outputs[9342] = ~(layer0_outputs[2484]);
    assign layer1_outputs[9343] = ~(layer0_outputs[243]) | (layer0_outputs[1456]);
    assign layer1_outputs[9344] = (layer0_outputs[5220]) ^ (layer0_outputs[9092]);
    assign layer1_outputs[9345] = (layer0_outputs[6170]) & ~(layer0_outputs[3483]);
    assign layer1_outputs[9346] = (layer0_outputs[6669]) & (layer0_outputs[8842]);
    assign layer1_outputs[9347] = ~(layer0_outputs[12093]);
    assign layer1_outputs[9348] = layer0_outputs[7968];
    assign layer1_outputs[9349] = ~(layer0_outputs[2436]);
    assign layer1_outputs[9350] = layer0_outputs[11787];
    assign layer1_outputs[9351] = ~(layer0_outputs[11573]);
    assign layer1_outputs[9352] = 1'b1;
    assign layer1_outputs[9353] = (layer0_outputs[6936]) | (layer0_outputs[377]);
    assign layer1_outputs[9354] = ~(layer0_outputs[3699]) | (layer0_outputs[8411]);
    assign layer1_outputs[9355] = (layer0_outputs[3981]) ^ (layer0_outputs[1884]);
    assign layer1_outputs[9356] = ~((layer0_outputs[10128]) & (layer0_outputs[12349]));
    assign layer1_outputs[9357] = layer0_outputs[3193];
    assign layer1_outputs[9358] = layer0_outputs[5819];
    assign layer1_outputs[9359] = ~((layer0_outputs[8903]) & (layer0_outputs[2264]));
    assign layer1_outputs[9360] = (layer0_outputs[10851]) & ~(layer0_outputs[8475]);
    assign layer1_outputs[9361] = ~(layer0_outputs[10656]) | (layer0_outputs[6692]);
    assign layer1_outputs[9362] = layer0_outputs[12760];
    assign layer1_outputs[9363] = (layer0_outputs[11276]) & ~(layer0_outputs[4002]);
    assign layer1_outputs[9364] = (layer0_outputs[3720]) | (layer0_outputs[11050]);
    assign layer1_outputs[9365] = ~(layer0_outputs[118]) | (layer0_outputs[2430]);
    assign layer1_outputs[9366] = (layer0_outputs[6680]) & (layer0_outputs[10641]);
    assign layer1_outputs[9367] = layer0_outputs[5896];
    assign layer1_outputs[9368] = ~(layer0_outputs[11822]);
    assign layer1_outputs[9369] = ~((layer0_outputs[10208]) & (layer0_outputs[2222]));
    assign layer1_outputs[9370] = (layer0_outputs[3125]) & ~(layer0_outputs[2494]);
    assign layer1_outputs[9371] = ~(layer0_outputs[8561]) | (layer0_outputs[4887]);
    assign layer1_outputs[9372] = ~(layer0_outputs[8322]);
    assign layer1_outputs[9373] = ~(layer0_outputs[2772]) | (layer0_outputs[2343]);
    assign layer1_outputs[9374] = (layer0_outputs[10446]) & (layer0_outputs[11763]);
    assign layer1_outputs[9375] = layer0_outputs[874];
    assign layer1_outputs[9376] = 1'b1;
    assign layer1_outputs[9377] = ~(layer0_outputs[8968]);
    assign layer1_outputs[9378] = ~((layer0_outputs[7781]) ^ (layer0_outputs[1584]));
    assign layer1_outputs[9379] = layer0_outputs[932];
    assign layer1_outputs[9380] = (layer0_outputs[11976]) | (layer0_outputs[6465]);
    assign layer1_outputs[9381] = layer0_outputs[6144];
    assign layer1_outputs[9382] = (layer0_outputs[6164]) & (layer0_outputs[8446]);
    assign layer1_outputs[9383] = ~(layer0_outputs[1429]);
    assign layer1_outputs[9384] = ~((layer0_outputs[7500]) ^ (layer0_outputs[155]));
    assign layer1_outputs[9385] = ~(layer0_outputs[4394]) | (layer0_outputs[12106]);
    assign layer1_outputs[9386] = ~((layer0_outputs[5402]) | (layer0_outputs[3015]));
    assign layer1_outputs[9387] = (layer0_outputs[10248]) & (layer0_outputs[4876]);
    assign layer1_outputs[9388] = (layer0_outputs[912]) & (layer0_outputs[8481]);
    assign layer1_outputs[9389] = ~((layer0_outputs[7246]) & (layer0_outputs[6904]));
    assign layer1_outputs[9390] = (layer0_outputs[2246]) & (layer0_outputs[4491]);
    assign layer1_outputs[9391] = layer0_outputs[9966];
    assign layer1_outputs[9392] = (layer0_outputs[9081]) | (layer0_outputs[7595]);
    assign layer1_outputs[9393] = layer0_outputs[6799];
    assign layer1_outputs[9394] = layer0_outputs[190];
    assign layer1_outputs[9395] = ~(layer0_outputs[9349]);
    assign layer1_outputs[9396] = ~(layer0_outputs[7604]) | (layer0_outputs[8172]);
    assign layer1_outputs[9397] = (layer0_outputs[10597]) | (layer0_outputs[7059]);
    assign layer1_outputs[9398] = ~((layer0_outputs[8347]) & (layer0_outputs[272]));
    assign layer1_outputs[9399] = ~(layer0_outputs[9649]) | (layer0_outputs[9449]);
    assign layer1_outputs[9400] = layer0_outputs[8913];
    assign layer1_outputs[9401] = (layer0_outputs[7823]) & (layer0_outputs[9156]);
    assign layer1_outputs[9402] = (layer0_outputs[6022]) | (layer0_outputs[4240]);
    assign layer1_outputs[9403] = layer0_outputs[6427];
    assign layer1_outputs[9404] = layer0_outputs[8307];
    assign layer1_outputs[9405] = (layer0_outputs[5997]) & ~(layer0_outputs[9108]);
    assign layer1_outputs[9406] = (layer0_outputs[23]) & ~(layer0_outputs[11400]);
    assign layer1_outputs[9407] = layer0_outputs[5466];
    assign layer1_outputs[9408] = ~(layer0_outputs[4086]);
    assign layer1_outputs[9409] = layer0_outputs[8843];
    assign layer1_outputs[9410] = ~((layer0_outputs[11849]) & (layer0_outputs[2016]));
    assign layer1_outputs[9411] = (layer0_outputs[10059]) | (layer0_outputs[2648]);
    assign layer1_outputs[9412] = ~(layer0_outputs[1267]);
    assign layer1_outputs[9413] = ~((layer0_outputs[3698]) | (layer0_outputs[3774]));
    assign layer1_outputs[9414] = (layer0_outputs[2079]) & (layer0_outputs[1234]);
    assign layer1_outputs[9415] = 1'b1;
    assign layer1_outputs[9416] = 1'b1;
    assign layer1_outputs[9417] = layer0_outputs[981];
    assign layer1_outputs[9418] = ~(layer0_outputs[5986]);
    assign layer1_outputs[9419] = (layer0_outputs[7392]) & ~(layer0_outputs[5579]);
    assign layer1_outputs[9420] = layer0_outputs[10456];
    assign layer1_outputs[9421] = ~(layer0_outputs[3659]) | (layer0_outputs[3636]);
    assign layer1_outputs[9422] = ~((layer0_outputs[8787]) | (layer0_outputs[2109]));
    assign layer1_outputs[9423] = (layer0_outputs[12081]) & ~(layer0_outputs[1620]);
    assign layer1_outputs[9424] = (layer0_outputs[8679]) | (layer0_outputs[6804]);
    assign layer1_outputs[9425] = ~(layer0_outputs[4361]);
    assign layer1_outputs[9426] = (layer0_outputs[10465]) & (layer0_outputs[10120]);
    assign layer1_outputs[9427] = (layer0_outputs[4330]) | (layer0_outputs[596]);
    assign layer1_outputs[9428] = (layer0_outputs[2668]) ^ (layer0_outputs[12314]);
    assign layer1_outputs[9429] = ~(layer0_outputs[869]) | (layer0_outputs[1940]);
    assign layer1_outputs[9430] = ~((layer0_outputs[11813]) | (layer0_outputs[6082]));
    assign layer1_outputs[9431] = ~(layer0_outputs[925]);
    assign layer1_outputs[9432] = layer0_outputs[10961];
    assign layer1_outputs[9433] = ~(layer0_outputs[9702]);
    assign layer1_outputs[9434] = ~(layer0_outputs[682]);
    assign layer1_outputs[9435] = 1'b1;
    assign layer1_outputs[9436] = (layer0_outputs[11536]) & (layer0_outputs[3661]);
    assign layer1_outputs[9437] = ~(layer0_outputs[6726]);
    assign layer1_outputs[9438] = ~((layer0_outputs[12785]) ^ (layer0_outputs[12786]));
    assign layer1_outputs[9439] = layer0_outputs[5426];
    assign layer1_outputs[9440] = (layer0_outputs[1483]) & ~(layer0_outputs[9202]);
    assign layer1_outputs[9441] = layer0_outputs[7885];
    assign layer1_outputs[9442] = ~(layer0_outputs[5625]);
    assign layer1_outputs[9443] = layer0_outputs[2492];
    assign layer1_outputs[9444] = ~(layer0_outputs[3698]);
    assign layer1_outputs[9445] = ~(layer0_outputs[12720]) | (layer0_outputs[8224]);
    assign layer1_outputs[9446] = ~(layer0_outputs[7687]) | (layer0_outputs[1067]);
    assign layer1_outputs[9447] = layer0_outputs[4939];
    assign layer1_outputs[9448] = (layer0_outputs[4323]) & ~(layer0_outputs[2924]);
    assign layer1_outputs[9449] = ~((layer0_outputs[11082]) & (layer0_outputs[12520]));
    assign layer1_outputs[9450] = (layer0_outputs[8460]) & ~(layer0_outputs[4149]);
    assign layer1_outputs[9451] = layer0_outputs[6168];
    assign layer1_outputs[9452] = (layer0_outputs[544]) | (layer0_outputs[3544]);
    assign layer1_outputs[9453] = (layer0_outputs[388]) & (layer0_outputs[435]);
    assign layer1_outputs[9454] = ~(layer0_outputs[9416]) | (layer0_outputs[8600]);
    assign layer1_outputs[9455] = ~(layer0_outputs[977]);
    assign layer1_outputs[9456] = (layer0_outputs[1981]) | (layer0_outputs[3930]);
    assign layer1_outputs[9457] = ~((layer0_outputs[3609]) ^ (layer0_outputs[2537]));
    assign layer1_outputs[9458] = ~(layer0_outputs[6151]) | (layer0_outputs[1239]);
    assign layer1_outputs[9459] = ~((layer0_outputs[11020]) ^ (layer0_outputs[8982]));
    assign layer1_outputs[9460] = (layer0_outputs[5165]) & ~(layer0_outputs[1294]);
    assign layer1_outputs[9461] = (layer0_outputs[10651]) & (layer0_outputs[3080]);
    assign layer1_outputs[9462] = ~((layer0_outputs[6367]) & (layer0_outputs[8480]));
    assign layer1_outputs[9463] = (layer0_outputs[3481]) ^ (layer0_outputs[6894]);
    assign layer1_outputs[9464] = ~(layer0_outputs[4736]) | (layer0_outputs[8313]);
    assign layer1_outputs[9465] = 1'b0;
    assign layer1_outputs[9466] = ~(layer0_outputs[9428]);
    assign layer1_outputs[9467] = (layer0_outputs[6004]) | (layer0_outputs[1377]);
    assign layer1_outputs[9468] = ~(layer0_outputs[8799]);
    assign layer1_outputs[9469] = (layer0_outputs[11123]) & ~(layer0_outputs[3425]);
    assign layer1_outputs[9470] = (layer0_outputs[11735]) & (layer0_outputs[410]);
    assign layer1_outputs[9471] = layer0_outputs[7731];
    assign layer1_outputs[9472] = ~(layer0_outputs[3916]) | (layer0_outputs[1317]);
    assign layer1_outputs[9473] = layer0_outputs[11047];
    assign layer1_outputs[9474] = ~(layer0_outputs[8464]) | (layer0_outputs[8463]);
    assign layer1_outputs[9475] = ~(layer0_outputs[12148]);
    assign layer1_outputs[9476] = ~(layer0_outputs[2655]) | (layer0_outputs[12171]);
    assign layer1_outputs[9477] = (layer0_outputs[4589]) ^ (layer0_outputs[3202]);
    assign layer1_outputs[9478] = ~(layer0_outputs[10197]) | (layer0_outputs[8256]);
    assign layer1_outputs[9479] = layer0_outputs[3798];
    assign layer1_outputs[9480] = (layer0_outputs[2407]) & ~(layer0_outputs[8441]);
    assign layer1_outputs[9481] = layer0_outputs[10899];
    assign layer1_outputs[9482] = ~(layer0_outputs[5734]) | (layer0_outputs[10312]);
    assign layer1_outputs[9483] = 1'b1;
    assign layer1_outputs[9484] = ~(layer0_outputs[1784]) | (layer0_outputs[9555]);
    assign layer1_outputs[9485] = ~(layer0_outputs[9132]);
    assign layer1_outputs[9486] = ~(layer0_outputs[2874]) | (layer0_outputs[8186]);
    assign layer1_outputs[9487] = ~((layer0_outputs[5756]) ^ (layer0_outputs[10905]));
    assign layer1_outputs[9488] = layer0_outputs[3092];
    assign layer1_outputs[9489] = (layer0_outputs[2455]) & ~(layer0_outputs[8715]);
    assign layer1_outputs[9490] = ~(layer0_outputs[6495]);
    assign layer1_outputs[9491] = layer0_outputs[10608];
    assign layer1_outputs[9492] = ~(layer0_outputs[2143]);
    assign layer1_outputs[9493] = ~(layer0_outputs[3359]) | (layer0_outputs[5432]);
    assign layer1_outputs[9494] = ~((layer0_outputs[1216]) | (layer0_outputs[4303]));
    assign layer1_outputs[9495] = ~((layer0_outputs[8655]) & (layer0_outputs[2552]));
    assign layer1_outputs[9496] = (layer0_outputs[8791]) | (layer0_outputs[11756]);
    assign layer1_outputs[9497] = ~((layer0_outputs[3405]) | (layer0_outputs[11764]));
    assign layer1_outputs[9498] = ~(layer0_outputs[7670]);
    assign layer1_outputs[9499] = (layer0_outputs[6510]) & ~(layer0_outputs[1965]);
    assign layer1_outputs[9500] = layer0_outputs[5489];
    assign layer1_outputs[9501] = (layer0_outputs[9572]) & ~(layer0_outputs[6388]);
    assign layer1_outputs[9502] = ~(layer0_outputs[10086]);
    assign layer1_outputs[9503] = ~(layer0_outputs[9403]);
    assign layer1_outputs[9504] = ~(layer0_outputs[10481]);
    assign layer1_outputs[9505] = ~((layer0_outputs[6866]) | (layer0_outputs[4376]));
    assign layer1_outputs[9506] = ~((layer0_outputs[1356]) | (layer0_outputs[9487]));
    assign layer1_outputs[9507] = 1'b0;
    assign layer1_outputs[9508] = ~(layer0_outputs[4390]);
    assign layer1_outputs[9509] = (layer0_outputs[1524]) | (layer0_outputs[9514]);
    assign layer1_outputs[9510] = ~(layer0_outputs[7329]) | (layer0_outputs[4524]);
    assign layer1_outputs[9511] = layer0_outputs[3912];
    assign layer1_outputs[9512] = (layer0_outputs[10828]) & ~(layer0_outputs[6973]);
    assign layer1_outputs[9513] = (layer0_outputs[563]) ^ (layer0_outputs[5053]);
    assign layer1_outputs[9514] = ~((layer0_outputs[6356]) & (layer0_outputs[3376]));
    assign layer1_outputs[9515] = ~((layer0_outputs[1949]) & (layer0_outputs[1810]));
    assign layer1_outputs[9516] = (layer0_outputs[4284]) ^ (layer0_outputs[7046]);
    assign layer1_outputs[9517] = ~(layer0_outputs[11951]);
    assign layer1_outputs[9518] = (layer0_outputs[3615]) | (layer0_outputs[3503]);
    assign layer1_outputs[9519] = ~((layer0_outputs[923]) | (layer0_outputs[109]));
    assign layer1_outputs[9520] = (layer0_outputs[3928]) | (layer0_outputs[9379]);
    assign layer1_outputs[9521] = 1'b0;
    assign layer1_outputs[9522] = 1'b1;
    assign layer1_outputs[9523] = ~((layer0_outputs[1926]) | (layer0_outputs[11606]));
    assign layer1_outputs[9524] = (layer0_outputs[2085]) ^ (layer0_outputs[6163]);
    assign layer1_outputs[9525] = ~(layer0_outputs[5459]) | (layer0_outputs[10789]);
    assign layer1_outputs[9526] = (layer0_outputs[3596]) & ~(layer0_outputs[5254]);
    assign layer1_outputs[9527] = layer0_outputs[3122];
    assign layer1_outputs[9528] = layer0_outputs[2917];
    assign layer1_outputs[9529] = (layer0_outputs[8560]) & ~(layer0_outputs[2155]);
    assign layer1_outputs[9530] = (layer0_outputs[7417]) & ~(layer0_outputs[9980]);
    assign layer1_outputs[9531] = ~((layer0_outputs[10068]) ^ (layer0_outputs[2093]));
    assign layer1_outputs[9532] = layer0_outputs[12753];
    assign layer1_outputs[9533] = (layer0_outputs[1282]) & ~(layer0_outputs[6034]);
    assign layer1_outputs[9534] = ~((layer0_outputs[7239]) & (layer0_outputs[37]));
    assign layer1_outputs[9535] = ~((layer0_outputs[8240]) & (layer0_outputs[5335]));
    assign layer1_outputs[9536] = ~(layer0_outputs[8054]);
    assign layer1_outputs[9537] = ~(layer0_outputs[11356]);
    assign layer1_outputs[9538] = (layer0_outputs[11195]) & ~(layer0_outputs[12478]);
    assign layer1_outputs[9539] = ~(layer0_outputs[6329]);
    assign layer1_outputs[9540] = ~((layer0_outputs[11288]) ^ (layer0_outputs[4997]));
    assign layer1_outputs[9541] = (layer0_outputs[1467]) & ~(layer0_outputs[3640]);
    assign layer1_outputs[9542] = ~(layer0_outputs[6790]) | (layer0_outputs[504]);
    assign layer1_outputs[9543] = ~((layer0_outputs[10035]) & (layer0_outputs[5974]));
    assign layer1_outputs[9544] = (layer0_outputs[5614]) | (layer0_outputs[6901]);
    assign layer1_outputs[9545] = ~((layer0_outputs[7752]) ^ (layer0_outputs[8811]));
    assign layer1_outputs[9546] = (layer0_outputs[4871]) & ~(layer0_outputs[10095]);
    assign layer1_outputs[9547] = layer0_outputs[6443];
    assign layer1_outputs[9548] = layer0_outputs[2058];
    assign layer1_outputs[9549] = (layer0_outputs[8096]) & (layer0_outputs[3521]);
    assign layer1_outputs[9550] = ~((layer0_outputs[5645]) ^ (layer0_outputs[542]));
    assign layer1_outputs[9551] = (layer0_outputs[5530]) & ~(layer0_outputs[4763]);
    assign layer1_outputs[9552] = (layer0_outputs[5649]) & ~(layer0_outputs[1435]);
    assign layer1_outputs[9553] = ~((layer0_outputs[7470]) & (layer0_outputs[6427]));
    assign layer1_outputs[9554] = 1'b0;
    assign layer1_outputs[9555] = ~((layer0_outputs[8413]) ^ (layer0_outputs[11726]));
    assign layer1_outputs[9556] = ~(layer0_outputs[9339]) | (layer0_outputs[3076]);
    assign layer1_outputs[9557] = (layer0_outputs[7778]) & ~(layer0_outputs[7297]);
    assign layer1_outputs[9558] = layer0_outputs[6330];
    assign layer1_outputs[9559] = (layer0_outputs[9192]) & ~(layer0_outputs[5691]);
    assign layer1_outputs[9560] = ~((layer0_outputs[1580]) | (layer0_outputs[9720]));
    assign layer1_outputs[9561] = (layer0_outputs[4517]) & ~(layer0_outputs[12698]);
    assign layer1_outputs[9562] = ~((layer0_outputs[5722]) | (layer0_outputs[6860]));
    assign layer1_outputs[9563] = ~((layer0_outputs[4483]) | (layer0_outputs[3745]));
    assign layer1_outputs[9564] = (layer0_outputs[2184]) & (layer0_outputs[4016]);
    assign layer1_outputs[9565] = ~(layer0_outputs[8929]) | (layer0_outputs[4911]);
    assign layer1_outputs[9566] = (layer0_outputs[8489]) & ~(layer0_outputs[11075]);
    assign layer1_outputs[9567] = ~(layer0_outputs[11469]) | (layer0_outputs[5168]);
    assign layer1_outputs[9568] = ~(layer0_outputs[12555]) | (layer0_outputs[4432]);
    assign layer1_outputs[9569] = ~(layer0_outputs[2782]) | (layer0_outputs[1388]);
    assign layer1_outputs[9570] = ~((layer0_outputs[12502]) | (layer0_outputs[12530]));
    assign layer1_outputs[9571] = (layer0_outputs[783]) ^ (layer0_outputs[1092]);
    assign layer1_outputs[9572] = ~((layer0_outputs[10947]) | (layer0_outputs[3995]));
    assign layer1_outputs[9573] = layer0_outputs[9387];
    assign layer1_outputs[9574] = (layer0_outputs[8470]) & (layer0_outputs[4963]);
    assign layer1_outputs[9575] = ~(layer0_outputs[68]) | (layer0_outputs[451]);
    assign layer1_outputs[9576] = (layer0_outputs[5869]) & ~(layer0_outputs[10021]);
    assign layer1_outputs[9577] = layer0_outputs[9675];
    assign layer1_outputs[9578] = ~(layer0_outputs[3269]) | (layer0_outputs[2716]);
    assign layer1_outputs[9579] = ~(layer0_outputs[10779]);
    assign layer1_outputs[9580] = layer0_outputs[2857];
    assign layer1_outputs[9581] = ~(layer0_outputs[4104]);
    assign layer1_outputs[9582] = (layer0_outputs[521]) ^ (layer0_outputs[7172]);
    assign layer1_outputs[9583] = (layer0_outputs[696]) & (layer0_outputs[10188]);
    assign layer1_outputs[9584] = ~(layer0_outputs[7438]) | (layer0_outputs[2025]);
    assign layer1_outputs[9585] = ~(layer0_outputs[3605]) | (layer0_outputs[3365]);
    assign layer1_outputs[9586] = (layer0_outputs[8997]) ^ (layer0_outputs[10071]);
    assign layer1_outputs[9587] = 1'b0;
    assign layer1_outputs[9588] = ~((layer0_outputs[7428]) | (layer0_outputs[649]));
    assign layer1_outputs[9589] = layer0_outputs[5413];
    assign layer1_outputs[9590] = ~(layer0_outputs[8683]) | (layer0_outputs[4011]);
    assign layer1_outputs[9591] = ~((layer0_outputs[3784]) | (layer0_outputs[9671]));
    assign layer1_outputs[9592] = ~(layer0_outputs[1457]);
    assign layer1_outputs[9593] = 1'b1;
    assign layer1_outputs[9594] = (layer0_outputs[8672]) ^ (layer0_outputs[8108]);
    assign layer1_outputs[9595] = layer0_outputs[3424];
    assign layer1_outputs[9596] = ~((layer0_outputs[1550]) & (layer0_outputs[1780]));
    assign layer1_outputs[9597] = ~(layer0_outputs[12583]);
    assign layer1_outputs[9598] = layer0_outputs[10007];
    assign layer1_outputs[9599] = (layer0_outputs[1276]) ^ (layer0_outputs[11328]);
    assign layer1_outputs[9600] = ~(layer0_outputs[4489]);
    assign layer1_outputs[9601] = (layer0_outputs[1399]) ^ (layer0_outputs[5882]);
    assign layer1_outputs[9602] = (layer0_outputs[3403]) & (layer0_outputs[3778]);
    assign layer1_outputs[9603] = ~((layer0_outputs[7906]) | (layer0_outputs[3885]));
    assign layer1_outputs[9604] = (layer0_outputs[7829]) ^ (layer0_outputs[3120]);
    assign layer1_outputs[9605] = (layer0_outputs[9951]) & (layer0_outputs[11926]);
    assign layer1_outputs[9606] = layer0_outputs[3708];
    assign layer1_outputs[9607] = ~((layer0_outputs[8129]) & (layer0_outputs[3653]));
    assign layer1_outputs[9608] = ~(layer0_outputs[8549]);
    assign layer1_outputs[9609] = ~(layer0_outputs[2490]);
    assign layer1_outputs[9610] = layer0_outputs[2203];
    assign layer1_outputs[9611] = ~(layer0_outputs[10345]);
    assign layer1_outputs[9612] = ~(layer0_outputs[534]) | (layer0_outputs[11402]);
    assign layer1_outputs[9613] = layer0_outputs[10786];
    assign layer1_outputs[9614] = (layer0_outputs[909]) ^ (layer0_outputs[4903]);
    assign layer1_outputs[9615] = ~(layer0_outputs[2746]);
    assign layer1_outputs[9616] = (layer0_outputs[7703]) & ~(layer0_outputs[7488]);
    assign layer1_outputs[9617] = ~(layer0_outputs[7074]);
    assign layer1_outputs[9618] = layer0_outputs[1389];
    assign layer1_outputs[9619] = layer0_outputs[3881];
    assign layer1_outputs[9620] = (layer0_outputs[10023]) & ~(layer0_outputs[3421]);
    assign layer1_outputs[9621] = (layer0_outputs[2656]) & ~(layer0_outputs[11065]);
    assign layer1_outputs[9622] = (layer0_outputs[10525]) & ~(layer0_outputs[2485]);
    assign layer1_outputs[9623] = (layer0_outputs[5143]) & ~(layer0_outputs[9150]);
    assign layer1_outputs[9624] = ~((layer0_outputs[430]) | (layer0_outputs[8681]));
    assign layer1_outputs[9625] = layer0_outputs[2341];
    assign layer1_outputs[9626] = ~((layer0_outputs[8897]) | (layer0_outputs[11142]));
    assign layer1_outputs[9627] = layer0_outputs[2222];
    assign layer1_outputs[9628] = ~((layer0_outputs[8181]) | (layer0_outputs[11805]));
    assign layer1_outputs[9629] = (layer0_outputs[7180]) | (layer0_outputs[1179]);
    assign layer1_outputs[9630] = layer0_outputs[2327];
    assign layer1_outputs[9631] = layer0_outputs[4916];
    assign layer1_outputs[9632] = ~((layer0_outputs[4221]) | (layer0_outputs[7122]));
    assign layer1_outputs[9633] = ~(layer0_outputs[5661]);
    assign layer1_outputs[9634] = (layer0_outputs[11204]) & ~(layer0_outputs[6894]);
    assign layer1_outputs[9635] = layer0_outputs[3256];
    assign layer1_outputs[9636] = ~(layer0_outputs[12176]);
    assign layer1_outputs[9637] = ~(layer0_outputs[838]);
    assign layer1_outputs[9638] = ~(layer0_outputs[5624]);
    assign layer1_outputs[9639] = ~(layer0_outputs[8097]) | (layer0_outputs[5379]);
    assign layer1_outputs[9640] = layer0_outputs[6261];
    assign layer1_outputs[9641] = layer0_outputs[7648];
    assign layer1_outputs[9642] = ~((layer0_outputs[3408]) | (layer0_outputs[5347]));
    assign layer1_outputs[9643] = ~(layer0_outputs[2687]) | (layer0_outputs[4907]);
    assign layer1_outputs[9644] = ~(layer0_outputs[10757]);
    assign layer1_outputs[9645] = ~((layer0_outputs[1712]) | (layer0_outputs[10444]));
    assign layer1_outputs[9646] = (layer0_outputs[1693]) & ~(layer0_outputs[6021]);
    assign layer1_outputs[9647] = (layer0_outputs[10895]) & ~(layer0_outputs[3572]);
    assign layer1_outputs[9648] = layer0_outputs[221];
    assign layer1_outputs[9649] = ~(layer0_outputs[2645]);
    assign layer1_outputs[9650] = ~((layer0_outputs[3274]) | (layer0_outputs[2767]));
    assign layer1_outputs[9651] = (layer0_outputs[3005]) ^ (layer0_outputs[8024]);
    assign layer1_outputs[9652] = (layer0_outputs[12788]) & (layer0_outputs[6086]);
    assign layer1_outputs[9653] = (layer0_outputs[12134]) & ~(layer0_outputs[2136]);
    assign layer1_outputs[9654] = ~(layer0_outputs[2370]);
    assign layer1_outputs[9655] = (layer0_outputs[12034]) & ~(layer0_outputs[12700]);
    assign layer1_outputs[9656] = layer0_outputs[5435];
    assign layer1_outputs[9657] = ~(layer0_outputs[3461]) | (layer0_outputs[11496]);
    assign layer1_outputs[9658] = (layer0_outputs[2177]) & ~(layer0_outputs[10695]);
    assign layer1_outputs[9659] = ~((layer0_outputs[11733]) ^ (layer0_outputs[6340]));
    assign layer1_outputs[9660] = ~(layer0_outputs[2976]) | (layer0_outputs[4962]);
    assign layer1_outputs[9661] = (layer0_outputs[8258]) ^ (layer0_outputs[2820]);
    assign layer1_outputs[9662] = ~(layer0_outputs[7734]);
    assign layer1_outputs[9663] = (layer0_outputs[668]) & ~(layer0_outputs[3535]);
    assign layer1_outputs[9664] = ~((layer0_outputs[9336]) ^ (layer0_outputs[5325]));
    assign layer1_outputs[9665] = ~(layer0_outputs[11310]) | (layer0_outputs[11376]);
    assign layer1_outputs[9666] = (layer0_outputs[5417]) & ~(layer0_outputs[10574]);
    assign layer1_outputs[9667] = ~(layer0_outputs[247]) | (layer0_outputs[1046]);
    assign layer1_outputs[9668] = 1'b1;
    assign layer1_outputs[9669] = layer0_outputs[11865];
    assign layer1_outputs[9670] = layer0_outputs[2123];
    assign layer1_outputs[9671] = ~((layer0_outputs[5194]) ^ (layer0_outputs[10450]));
    assign layer1_outputs[9672] = ~(layer0_outputs[1615]) | (layer0_outputs[9553]);
    assign layer1_outputs[9673] = (layer0_outputs[9214]) & ~(layer0_outputs[11794]);
    assign layer1_outputs[9674] = layer0_outputs[7318];
    assign layer1_outputs[9675] = (layer0_outputs[0]) & ~(layer0_outputs[10486]);
    assign layer1_outputs[9676] = layer0_outputs[10602];
    assign layer1_outputs[9677] = ~((layer0_outputs[3734]) | (layer0_outputs[8087]));
    assign layer1_outputs[9678] = ~((layer0_outputs[2560]) | (layer0_outputs[4179]));
    assign layer1_outputs[9679] = (layer0_outputs[5111]) | (layer0_outputs[8079]);
    assign layer1_outputs[9680] = (layer0_outputs[5341]) & (layer0_outputs[5364]);
    assign layer1_outputs[9681] = ~(layer0_outputs[6642]);
    assign layer1_outputs[9682] = ~(layer0_outputs[8012]);
    assign layer1_outputs[9683] = ~((layer0_outputs[3340]) ^ (layer0_outputs[7820]));
    assign layer1_outputs[9684] = (layer0_outputs[11468]) & ~(layer0_outputs[7137]);
    assign layer1_outputs[9685] = ~(layer0_outputs[9071]) | (layer0_outputs[8350]);
    assign layer1_outputs[9686] = ~(layer0_outputs[7900]);
    assign layer1_outputs[9687] = ~(layer0_outputs[8395]) | (layer0_outputs[10480]);
    assign layer1_outputs[9688] = ~(layer0_outputs[7888]);
    assign layer1_outputs[9689] = layer0_outputs[7447];
    assign layer1_outputs[9690] = ~(layer0_outputs[3367]);
    assign layer1_outputs[9691] = ~(layer0_outputs[7350]) | (layer0_outputs[4541]);
    assign layer1_outputs[9692] = (layer0_outputs[726]) & ~(layer0_outputs[8188]);
    assign layer1_outputs[9693] = (layer0_outputs[12354]) ^ (layer0_outputs[115]);
    assign layer1_outputs[9694] = ~((layer0_outputs[2029]) | (layer0_outputs[4304]));
    assign layer1_outputs[9695] = layer0_outputs[7330];
    assign layer1_outputs[9696] = ~((layer0_outputs[2798]) & (layer0_outputs[5552]));
    assign layer1_outputs[9697] = (layer0_outputs[7561]) & ~(layer0_outputs[4257]);
    assign layer1_outputs[9698] = ~(layer0_outputs[5904]);
    assign layer1_outputs[9699] = layer0_outputs[6852];
    assign layer1_outputs[9700] = ~(layer0_outputs[6935]) | (layer0_outputs[3207]);
    assign layer1_outputs[9701] = (layer0_outputs[623]) & ~(layer0_outputs[6017]);
    assign layer1_outputs[9702] = ~(layer0_outputs[9318]);
    assign layer1_outputs[9703] = ~((layer0_outputs[4154]) ^ (layer0_outputs[7116]));
    assign layer1_outputs[9704] = (layer0_outputs[7496]) ^ (layer0_outputs[2576]);
    assign layer1_outputs[9705] = (layer0_outputs[3833]) & ~(layer0_outputs[6289]);
    assign layer1_outputs[9706] = layer0_outputs[6637];
    assign layer1_outputs[9707] = (layer0_outputs[7847]) & ~(layer0_outputs[7797]);
    assign layer1_outputs[9708] = ~((layer0_outputs[9760]) & (layer0_outputs[9797]));
    assign layer1_outputs[9709] = ~((layer0_outputs[5866]) & (layer0_outputs[1487]));
    assign layer1_outputs[9710] = (layer0_outputs[9317]) | (layer0_outputs[2026]);
    assign layer1_outputs[9711] = 1'b1;
    assign layer1_outputs[9712] = ~(layer0_outputs[6161]);
    assign layer1_outputs[9713] = (layer0_outputs[10099]) & (layer0_outputs[11104]);
    assign layer1_outputs[9714] = ~((layer0_outputs[7801]) ^ (layer0_outputs[7777]));
    assign layer1_outputs[9715] = ~((layer0_outputs[8145]) ^ (layer0_outputs[994]));
    assign layer1_outputs[9716] = ~(layer0_outputs[5888]);
    assign layer1_outputs[9717] = ~((layer0_outputs[4048]) | (layer0_outputs[970]));
    assign layer1_outputs[9718] = ~(layer0_outputs[8379]);
    assign layer1_outputs[9719] = layer0_outputs[10517];
    assign layer1_outputs[9720] = ~(layer0_outputs[10506]) | (layer0_outputs[10295]);
    assign layer1_outputs[9721] = (layer0_outputs[10376]) & ~(layer0_outputs[5142]);
    assign layer1_outputs[9722] = layer0_outputs[5290];
    assign layer1_outputs[9723] = ~(layer0_outputs[2935]);
    assign layer1_outputs[9724] = ~(layer0_outputs[2327]);
    assign layer1_outputs[9725] = layer0_outputs[4375];
    assign layer1_outputs[9726] = layer0_outputs[3508];
    assign layer1_outputs[9727] = 1'b1;
    assign layer1_outputs[9728] = (layer0_outputs[7696]) & ~(layer0_outputs[5112]);
    assign layer1_outputs[9729] = ~((layer0_outputs[10094]) & (layer0_outputs[7014]));
    assign layer1_outputs[9730] = ~(layer0_outputs[774]) | (layer0_outputs[10399]);
    assign layer1_outputs[9731] = layer0_outputs[12730];
    assign layer1_outputs[9732] = ~(layer0_outputs[10390]);
    assign layer1_outputs[9733] = layer0_outputs[1663];
    assign layer1_outputs[9734] = ~(layer0_outputs[3038]);
    assign layer1_outputs[9735] = ~((layer0_outputs[4272]) ^ (layer0_outputs[4281]));
    assign layer1_outputs[9736] = ~(layer0_outputs[6005]);
    assign layer1_outputs[9737] = (layer0_outputs[202]) & (layer0_outputs[8793]);
    assign layer1_outputs[9738] = ~(layer0_outputs[10392]) | (layer0_outputs[12392]);
    assign layer1_outputs[9739] = (layer0_outputs[197]) & ~(layer0_outputs[4965]);
    assign layer1_outputs[9740] = layer0_outputs[4220];
    assign layer1_outputs[9741] = (layer0_outputs[3271]) & (layer0_outputs[2125]);
    assign layer1_outputs[9742] = ~(layer0_outputs[7923]);
    assign layer1_outputs[9743] = ~(layer0_outputs[9865]);
    assign layer1_outputs[9744] = layer0_outputs[6181];
    assign layer1_outputs[9745] = (layer0_outputs[9323]) & ~(layer0_outputs[4922]);
    assign layer1_outputs[9746] = ~((layer0_outputs[7021]) ^ (layer0_outputs[7795]));
    assign layer1_outputs[9747] = ~(layer0_outputs[3844]);
    assign layer1_outputs[9748] = ~(layer0_outputs[8893]) | (layer0_outputs[2208]);
    assign layer1_outputs[9749] = ~((layer0_outputs[4812]) & (layer0_outputs[9977]));
    assign layer1_outputs[9750] = layer0_outputs[11695];
    assign layer1_outputs[9751] = layer0_outputs[1861];
    assign layer1_outputs[9752] = (layer0_outputs[11490]) & (layer0_outputs[5085]);
    assign layer1_outputs[9753] = ~(layer0_outputs[9930]);
    assign layer1_outputs[9754] = ~(layer0_outputs[9698]) | (layer0_outputs[10011]);
    assign layer1_outputs[9755] = 1'b1;
    assign layer1_outputs[9756] = layer0_outputs[4228];
    assign layer1_outputs[9757] = (layer0_outputs[5017]) & (layer0_outputs[7890]);
    assign layer1_outputs[9758] = ~(layer0_outputs[5710]);
    assign layer1_outputs[9759] = layer0_outputs[4277];
    assign layer1_outputs[9760] = ~((layer0_outputs[9349]) ^ (layer0_outputs[319]));
    assign layer1_outputs[9761] = ~(layer0_outputs[11911]);
    assign layer1_outputs[9762] = (layer0_outputs[4827]) ^ (layer0_outputs[11007]);
    assign layer1_outputs[9763] = ~(layer0_outputs[1363]);
    assign layer1_outputs[9764] = ~(layer0_outputs[1291]);
    assign layer1_outputs[9765] = (layer0_outputs[12201]) | (layer0_outputs[3557]);
    assign layer1_outputs[9766] = (layer0_outputs[1906]) ^ (layer0_outputs[7861]);
    assign layer1_outputs[9767] = ~(layer0_outputs[6399]) | (layer0_outputs[5129]);
    assign layer1_outputs[9768] = (layer0_outputs[10162]) | (layer0_outputs[8465]);
    assign layer1_outputs[9769] = (layer0_outputs[2118]) & ~(layer0_outputs[4750]);
    assign layer1_outputs[9770] = (layer0_outputs[8899]) & ~(layer0_outputs[4627]);
    assign layer1_outputs[9771] = ~(layer0_outputs[4912]) | (layer0_outputs[658]);
    assign layer1_outputs[9772] = ~(layer0_outputs[8307]);
    assign layer1_outputs[9773] = layer0_outputs[6599];
    assign layer1_outputs[9774] = ~((layer0_outputs[11093]) | (layer0_outputs[1491]));
    assign layer1_outputs[9775] = ~(layer0_outputs[3857]) | (layer0_outputs[7645]);
    assign layer1_outputs[9776] = ~(layer0_outputs[6196]);
    assign layer1_outputs[9777] = (layer0_outputs[11954]) | (layer0_outputs[4424]);
    assign layer1_outputs[9778] = ~((layer0_outputs[10536]) & (layer0_outputs[8061]));
    assign layer1_outputs[9779] = (layer0_outputs[1141]) | (layer0_outputs[4863]);
    assign layer1_outputs[9780] = ~(layer0_outputs[12159]);
    assign layer1_outputs[9781] = ~((layer0_outputs[1852]) & (layer0_outputs[7363]));
    assign layer1_outputs[9782] = layer0_outputs[2302];
    assign layer1_outputs[9783] = layer0_outputs[10983];
    assign layer1_outputs[9784] = layer0_outputs[11018];
    assign layer1_outputs[9785] = (layer0_outputs[1577]) & (layer0_outputs[1369]);
    assign layer1_outputs[9786] = ~((layer0_outputs[2773]) ^ (layer0_outputs[10898]));
    assign layer1_outputs[9787] = ~(layer0_outputs[6627]);
    assign layer1_outputs[9788] = (layer0_outputs[8255]) ^ (layer0_outputs[2274]);
    assign layer1_outputs[9789] = 1'b0;
    assign layer1_outputs[9790] = layer0_outputs[5383];
    assign layer1_outputs[9791] = ~(layer0_outputs[4697]) | (layer0_outputs[8506]);
    assign layer1_outputs[9792] = layer0_outputs[10148];
    assign layer1_outputs[9793] = layer0_outputs[4473];
    assign layer1_outputs[9794] = (layer0_outputs[1032]) & ~(layer0_outputs[8952]);
    assign layer1_outputs[9795] = layer0_outputs[10780];
    assign layer1_outputs[9796] = (layer0_outputs[2044]) & (layer0_outputs[892]);
    assign layer1_outputs[9797] = layer0_outputs[2794];
    assign layer1_outputs[9798] = ~(layer0_outputs[10090]);
    assign layer1_outputs[9799] = ~((layer0_outputs[10099]) | (layer0_outputs[12238]));
    assign layer1_outputs[9800] = (layer0_outputs[10942]) & (layer0_outputs[6099]);
    assign layer1_outputs[9801] = ~(layer0_outputs[10387]) | (layer0_outputs[10018]);
    assign layer1_outputs[9802] = ~(layer0_outputs[12487]);
    assign layer1_outputs[9803] = layer0_outputs[6768];
    assign layer1_outputs[9804] = (layer0_outputs[2159]) & ~(layer0_outputs[5686]);
    assign layer1_outputs[9805] = (layer0_outputs[2564]) & ~(layer0_outputs[9056]);
    assign layer1_outputs[9806] = (layer0_outputs[946]) & ~(layer0_outputs[4170]);
    assign layer1_outputs[9807] = layer0_outputs[1187];
    assign layer1_outputs[9808] = ~((layer0_outputs[6180]) | (layer0_outputs[2975]));
    assign layer1_outputs[9809] = ~((layer0_outputs[2847]) & (layer0_outputs[105]));
    assign layer1_outputs[9810] = (layer0_outputs[11582]) & (layer0_outputs[1168]);
    assign layer1_outputs[9811] = (layer0_outputs[454]) & (layer0_outputs[5892]);
    assign layer1_outputs[9812] = ~(layer0_outputs[621]);
    assign layer1_outputs[9813] = ~(layer0_outputs[12335]);
    assign layer1_outputs[9814] = ~(layer0_outputs[8185]);
    assign layer1_outputs[9815] = ~(layer0_outputs[6403]) | (layer0_outputs[8061]);
    assign layer1_outputs[9816] = ~((layer0_outputs[755]) & (layer0_outputs[10368]));
    assign layer1_outputs[9817] = ~(layer0_outputs[10180]);
    assign layer1_outputs[9818] = ~(layer0_outputs[3397]);
    assign layer1_outputs[9819] = layer0_outputs[12729];
    assign layer1_outputs[9820] = ~(layer0_outputs[9039]) | (layer0_outputs[3294]);
    assign layer1_outputs[9821] = layer0_outputs[11560];
    assign layer1_outputs[9822] = layer0_outputs[788];
    assign layer1_outputs[9823] = ~(layer0_outputs[3085]) | (layer0_outputs[1854]);
    assign layer1_outputs[9824] = ~(layer0_outputs[6754]) | (layer0_outputs[2183]);
    assign layer1_outputs[9825] = layer0_outputs[11355];
    assign layer1_outputs[9826] = ~(layer0_outputs[4199]);
    assign layer1_outputs[9827] = ~((layer0_outputs[5039]) ^ (layer0_outputs[3527]));
    assign layer1_outputs[9828] = ~((layer0_outputs[7422]) ^ (layer0_outputs[7463]));
    assign layer1_outputs[9829] = layer0_outputs[9904];
    assign layer1_outputs[9830] = ~(layer0_outputs[6042]);
    assign layer1_outputs[9831] = (layer0_outputs[3298]) & ~(layer0_outputs[12367]);
    assign layer1_outputs[9832] = layer0_outputs[10424];
    assign layer1_outputs[9833] = (layer0_outputs[10813]) & (layer0_outputs[7742]);
    assign layer1_outputs[9834] = layer0_outputs[9843];
    assign layer1_outputs[9835] = layer0_outputs[7725];
    assign layer1_outputs[9836] = ~((layer0_outputs[5720]) ^ (layer0_outputs[7320]));
    assign layer1_outputs[9837] = layer0_outputs[9784];
    assign layer1_outputs[9838] = (layer0_outputs[9468]) & ~(layer0_outputs[8363]);
    assign layer1_outputs[9839] = (layer0_outputs[9973]) & ~(layer0_outputs[4589]);
    assign layer1_outputs[9840] = ~(layer0_outputs[9359]);
    assign layer1_outputs[9841] = ~(layer0_outputs[6503]) | (layer0_outputs[9393]);
    assign layer1_outputs[9842] = (layer0_outputs[1668]) ^ (layer0_outputs[11312]);
    assign layer1_outputs[9843] = layer0_outputs[7365];
    assign layer1_outputs[9844] = layer0_outputs[6247];
    assign layer1_outputs[9845] = ~(layer0_outputs[2934]);
    assign layer1_outputs[9846] = ~(layer0_outputs[2723]) | (layer0_outputs[7169]);
    assign layer1_outputs[9847] = layer0_outputs[11980];
    assign layer1_outputs[9848] = ~((layer0_outputs[11672]) & (layer0_outputs[1936]));
    assign layer1_outputs[9849] = layer0_outputs[10498];
    assign layer1_outputs[9850] = ~(layer0_outputs[1383]) | (layer0_outputs[3499]);
    assign layer1_outputs[9851] = ~(layer0_outputs[14]);
    assign layer1_outputs[9852] = 1'b0;
    assign layer1_outputs[9853] = ~((layer0_outputs[12511]) ^ (layer0_outputs[1256]));
    assign layer1_outputs[9854] = 1'b0;
    assign layer1_outputs[9855] = layer0_outputs[8280];
    assign layer1_outputs[9856] = layer0_outputs[3146];
    assign layer1_outputs[9857] = 1'b0;
    assign layer1_outputs[9858] = ~(layer0_outputs[7258]);
    assign layer1_outputs[9859] = (layer0_outputs[4383]) & ~(layer0_outputs[278]);
    assign layer1_outputs[9860] = ~((layer0_outputs[9585]) | (layer0_outputs[7942]));
    assign layer1_outputs[9861] = layer0_outputs[3801];
    assign layer1_outputs[9862] = layer0_outputs[7110];
    assign layer1_outputs[9863] = layer0_outputs[1974];
    assign layer1_outputs[9864] = (layer0_outputs[5756]) | (layer0_outputs[3215]);
    assign layer1_outputs[9865] = ~(layer0_outputs[8336]);
    assign layer1_outputs[9866] = (layer0_outputs[1731]) ^ (layer0_outputs[1537]);
    assign layer1_outputs[9867] = (layer0_outputs[10154]) ^ (layer0_outputs[8768]);
    assign layer1_outputs[9868] = ~(layer0_outputs[11796]) | (layer0_outputs[1835]);
    assign layer1_outputs[9869] = layer0_outputs[954];
    assign layer1_outputs[9870] = ~(layer0_outputs[3092]) | (layer0_outputs[2809]);
    assign layer1_outputs[9871] = layer0_outputs[8838];
    assign layer1_outputs[9872] = (layer0_outputs[7032]) & ~(layer0_outputs[7457]);
    assign layer1_outputs[9873] = ~(layer0_outputs[8882]) | (layer0_outputs[8427]);
    assign layer1_outputs[9874] = layer0_outputs[1548];
    assign layer1_outputs[9875] = (layer0_outputs[12583]) & (layer0_outputs[829]);
    assign layer1_outputs[9876] = layer0_outputs[1653];
    assign layer1_outputs[9877] = (layer0_outputs[2054]) & (layer0_outputs[4239]);
    assign layer1_outputs[9878] = ~(layer0_outputs[10253]);
    assign layer1_outputs[9879] = layer0_outputs[1918];
    assign layer1_outputs[9880] = layer0_outputs[2629];
    assign layer1_outputs[9881] = layer0_outputs[11896];
    assign layer1_outputs[9882] = layer0_outputs[4934];
    assign layer1_outputs[9883] = ~((layer0_outputs[3616]) | (layer0_outputs[88]));
    assign layer1_outputs[9884] = (layer0_outputs[12088]) ^ (layer0_outputs[10164]);
    assign layer1_outputs[9885] = (layer0_outputs[11660]) & ~(layer0_outputs[6803]);
    assign layer1_outputs[9886] = ~((layer0_outputs[2048]) | (layer0_outputs[7788]));
    assign layer1_outputs[9887] = ~(layer0_outputs[775]);
    assign layer1_outputs[9888] = ~(layer0_outputs[11441]);
    assign layer1_outputs[9889] = ~(layer0_outputs[4387]);
    assign layer1_outputs[9890] = layer0_outputs[7222];
    assign layer1_outputs[9891] = (layer0_outputs[11116]) & ~(layer0_outputs[2730]);
    assign layer1_outputs[9892] = ~(layer0_outputs[4808]);
    assign layer1_outputs[9893] = (layer0_outputs[1257]) & ~(layer0_outputs[9594]);
    assign layer1_outputs[9894] = ~(layer0_outputs[4761]) | (layer0_outputs[8028]);
    assign layer1_outputs[9895] = layer0_outputs[4552];
    assign layer1_outputs[9896] = layer0_outputs[3213];
    assign layer1_outputs[9897] = ~(layer0_outputs[11459]);
    assign layer1_outputs[9898] = ~((layer0_outputs[1020]) | (layer0_outputs[5713]));
    assign layer1_outputs[9899] = ~((layer0_outputs[10662]) | (layer0_outputs[6997]));
    assign layer1_outputs[9900] = layer0_outputs[866];
    assign layer1_outputs[9901] = ~(layer0_outputs[11618]);
    assign layer1_outputs[9902] = ~(layer0_outputs[12390]);
    assign layer1_outputs[9903] = ~((layer0_outputs[8298]) ^ (layer0_outputs[11793]));
    assign layer1_outputs[9904] = ~((layer0_outputs[1471]) ^ (layer0_outputs[11128]));
    assign layer1_outputs[9905] = (layer0_outputs[3039]) & ~(layer0_outputs[8417]);
    assign layer1_outputs[9906] = ~(layer0_outputs[3029]);
    assign layer1_outputs[9907] = ~(layer0_outputs[9242]);
    assign layer1_outputs[9908] = layer0_outputs[12698];
    assign layer1_outputs[9909] = ~(layer0_outputs[6833]);
    assign layer1_outputs[9910] = (layer0_outputs[1649]) & ~(layer0_outputs[1423]);
    assign layer1_outputs[9911] = layer0_outputs[9137];
    assign layer1_outputs[9912] = ~(layer0_outputs[10010]);
    assign layer1_outputs[9913] = layer0_outputs[5169];
    assign layer1_outputs[9914] = (layer0_outputs[7069]) & ~(layer0_outputs[482]);
    assign layer1_outputs[9915] = 1'b1;
    assign layer1_outputs[9916] = (layer0_outputs[6326]) ^ (layer0_outputs[3722]);
    assign layer1_outputs[9917] = layer0_outputs[2981];
    assign layer1_outputs[9918] = ~((layer0_outputs[11252]) | (layer0_outputs[1087]));
    assign layer1_outputs[9919] = ~((layer0_outputs[11176]) ^ (layer0_outputs[10160]));
    assign layer1_outputs[9920] = (layer0_outputs[6633]) & ~(layer0_outputs[2558]);
    assign layer1_outputs[9921] = (layer0_outputs[2068]) & ~(layer0_outputs[10797]);
    assign layer1_outputs[9922] = ~(layer0_outputs[2161]);
    assign layer1_outputs[9923] = ~(layer0_outputs[7598]);
    assign layer1_outputs[9924] = layer0_outputs[7379];
    assign layer1_outputs[9925] = ~(layer0_outputs[7693]);
    assign layer1_outputs[9926] = ~(layer0_outputs[11846]);
    assign layer1_outputs[9927] = (layer0_outputs[10043]) & ~(layer0_outputs[8872]);
    assign layer1_outputs[9928] = layer0_outputs[6240];
    assign layer1_outputs[9929] = ~(layer0_outputs[5301]);
    assign layer1_outputs[9930] = ~(layer0_outputs[976]) | (layer0_outputs[8762]);
    assign layer1_outputs[9931] = ~(layer0_outputs[3304]);
    assign layer1_outputs[9932] = 1'b0;
    assign layer1_outputs[9933] = (layer0_outputs[8173]) & (layer0_outputs[17]);
    assign layer1_outputs[9934] = (layer0_outputs[11463]) & (layer0_outputs[4965]);
    assign layer1_outputs[9935] = 1'b0;
    assign layer1_outputs[9936] = ~(layer0_outputs[3254]);
    assign layer1_outputs[9937] = layer0_outputs[5465];
    assign layer1_outputs[9938] = ~(layer0_outputs[1133]);
    assign layer1_outputs[9939] = layer0_outputs[12307];
    assign layer1_outputs[9940] = ~(layer0_outputs[1817]);
    assign layer1_outputs[9941] = (layer0_outputs[1436]) & (layer0_outputs[12495]);
    assign layer1_outputs[9942] = ~(layer0_outputs[4440]) | (layer0_outputs[10900]);
    assign layer1_outputs[9943] = ~((layer0_outputs[3376]) ^ (layer0_outputs[7415]));
    assign layer1_outputs[9944] = layer0_outputs[12450];
    assign layer1_outputs[9945] = ~(layer0_outputs[10718]) | (layer0_outputs[12475]);
    assign layer1_outputs[9946] = ~((layer0_outputs[1089]) | (layer0_outputs[3783]));
    assign layer1_outputs[9947] = ~((layer0_outputs[335]) ^ (layer0_outputs[6385]));
    assign layer1_outputs[9948] = layer0_outputs[6336];
    assign layer1_outputs[9949] = ~(layer0_outputs[6045]) | (layer0_outputs[4088]);
    assign layer1_outputs[9950] = layer0_outputs[341];
    assign layer1_outputs[9951] = (layer0_outputs[5973]) & ~(layer0_outputs[5901]);
    assign layer1_outputs[9952] = ~(layer0_outputs[5494]);
    assign layer1_outputs[9953] = layer0_outputs[3227];
    assign layer1_outputs[9954] = ~(layer0_outputs[5262]) | (layer0_outputs[1942]);
    assign layer1_outputs[9955] = (layer0_outputs[8075]) & (layer0_outputs[8975]);
    assign layer1_outputs[9956] = layer0_outputs[11627];
    assign layer1_outputs[9957] = (layer0_outputs[349]) & ~(layer0_outputs[1391]);
    assign layer1_outputs[9958] = ~(layer0_outputs[940]);
    assign layer1_outputs[9959] = (layer0_outputs[3089]) & (layer0_outputs[6423]);
    assign layer1_outputs[9960] = (layer0_outputs[6458]) ^ (layer0_outputs[2407]);
    assign layer1_outputs[9961] = ~((layer0_outputs[1379]) ^ (layer0_outputs[7309]));
    assign layer1_outputs[9962] = (layer0_outputs[3914]) ^ (layer0_outputs[5110]);
    assign layer1_outputs[9963] = ~(layer0_outputs[5862]) | (layer0_outputs[4768]);
    assign layer1_outputs[9964] = (layer0_outputs[8839]) & (layer0_outputs[1800]);
    assign layer1_outputs[9965] = (layer0_outputs[7062]) & (layer0_outputs[4933]);
    assign layer1_outputs[9966] = (layer0_outputs[12682]) ^ (layer0_outputs[10000]);
    assign layer1_outputs[9967] = ~((layer0_outputs[11018]) ^ (layer0_outputs[4481]));
    assign layer1_outputs[9968] = ~((layer0_outputs[1290]) | (layer0_outputs[11748]));
    assign layer1_outputs[9969] = ~(layer0_outputs[848]);
    assign layer1_outputs[9970] = (layer0_outputs[7078]) & (layer0_outputs[9992]);
    assign layer1_outputs[9971] = (layer0_outputs[7109]) & ~(layer0_outputs[10821]);
    assign layer1_outputs[9972] = layer0_outputs[5264];
    assign layer1_outputs[9973] = (layer0_outputs[6208]) & ~(layer0_outputs[4914]);
    assign layer1_outputs[9974] = ~(layer0_outputs[2618]);
    assign layer1_outputs[9975] = (layer0_outputs[5986]) | (layer0_outputs[5816]);
    assign layer1_outputs[9976] = ~(layer0_outputs[4708]);
    assign layer1_outputs[9977] = layer0_outputs[11386];
    assign layer1_outputs[9978] = ~(layer0_outputs[3140]) | (layer0_outputs[8272]);
    assign layer1_outputs[9979] = (layer0_outputs[4017]) & (layer0_outputs[6528]);
    assign layer1_outputs[9980] = ~(layer0_outputs[1134]);
    assign layer1_outputs[9981] = ~((layer0_outputs[3568]) ^ (layer0_outputs[5502]));
    assign layer1_outputs[9982] = layer0_outputs[9174];
    assign layer1_outputs[9983] = (layer0_outputs[10869]) & ~(layer0_outputs[4438]);
    assign layer1_outputs[9984] = ~((layer0_outputs[7287]) | (layer0_outputs[6650]));
    assign layer1_outputs[9985] = ~((layer0_outputs[2081]) & (layer0_outputs[9753]));
    assign layer1_outputs[9986] = ~((layer0_outputs[12664]) & (layer0_outputs[10178]));
    assign layer1_outputs[9987] = (layer0_outputs[12287]) & ~(layer0_outputs[11225]);
    assign layer1_outputs[9988] = ~(layer0_outputs[9552]);
    assign layer1_outputs[9989] = ~((layer0_outputs[734]) ^ (layer0_outputs[11546]));
    assign layer1_outputs[9990] = (layer0_outputs[3260]) | (layer0_outputs[6123]);
    assign layer1_outputs[9991] = layer0_outputs[4306];
    assign layer1_outputs[9992] = ~(layer0_outputs[9741]) | (layer0_outputs[4219]);
    assign layer1_outputs[9993] = (layer0_outputs[5216]) | (layer0_outputs[9372]);
    assign layer1_outputs[9994] = layer0_outputs[2588];
    assign layer1_outputs[9995] = ~((layer0_outputs[6686]) & (layer0_outputs[6913]));
    assign layer1_outputs[9996] = (layer0_outputs[12595]) & ~(layer0_outputs[4448]);
    assign layer1_outputs[9997] = ~(layer0_outputs[7892]);
    assign layer1_outputs[9998] = ~(layer0_outputs[2237]) | (layer0_outputs[5414]);
    assign layer1_outputs[9999] = ~(layer0_outputs[10657]) | (layer0_outputs[5448]);
    assign layer1_outputs[10000] = (layer0_outputs[1652]) & ~(layer0_outputs[5875]);
    assign layer1_outputs[10001] = layer0_outputs[7726];
    assign layer1_outputs[10002] = layer0_outputs[11667];
    assign layer1_outputs[10003] = (layer0_outputs[5955]) & ~(layer0_outputs[7505]);
    assign layer1_outputs[10004] = (layer0_outputs[9788]) & (layer0_outputs[11379]);
    assign layer1_outputs[10005] = ~((layer0_outputs[7347]) & (layer0_outputs[1678]));
    assign layer1_outputs[10006] = (layer0_outputs[10450]) | (layer0_outputs[2913]);
    assign layer1_outputs[10007] = ~((layer0_outputs[9806]) | (layer0_outputs[5800]));
    assign layer1_outputs[10008] = (layer0_outputs[11412]) | (layer0_outputs[7587]);
    assign layer1_outputs[10009] = ~(layer0_outputs[365]);
    assign layer1_outputs[10010] = (layer0_outputs[7263]) ^ (layer0_outputs[1537]);
    assign layer1_outputs[10011] = 1'b1;
    assign layer1_outputs[10012] = ~(layer0_outputs[8860]);
    assign layer1_outputs[10013] = ~((layer0_outputs[6342]) | (layer0_outputs[9230]));
    assign layer1_outputs[10014] = layer0_outputs[12479];
    assign layer1_outputs[10015] = ~(layer0_outputs[9190]);
    assign layer1_outputs[10016] = ~(layer0_outputs[4342]);
    assign layer1_outputs[10017] = layer0_outputs[4738];
    assign layer1_outputs[10018] = (layer0_outputs[997]) | (layer0_outputs[809]);
    assign layer1_outputs[10019] = ~(layer0_outputs[6901]);
    assign layer1_outputs[10020] = ~(layer0_outputs[10896]) | (layer0_outputs[2278]);
    assign layer1_outputs[10021] = ~(layer0_outputs[8456]) | (layer0_outputs[6687]);
    assign layer1_outputs[10022] = (layer0_outputs[8276]) & ~(layer0_outputs[10830]);
    assign layer1_outputs[10023] = layer0_outputs[10846];
    assign layer1_outputs[10024] = ~(layer0_outputs[6621]);
    assign layer1_outputs[10025] = (layer0_outputs[4892]) & ~(layer0_outputs[668]);
    assign layer1_outputs[10026] = ~(layer0_outputs[7244]) | (layer0_outputs[12787]);
    assign layer1_outputs[10027] = layer0_outputs[7982];
    assign layer1_outputs[10028] = layer0_outputs[12117];
    assign layer1_outputs[10029] = layer0_outputs[1608];
    assign layer1_outputs[10030] = (layer0_outputs[7056]) | (layer0_outputs[4058]);
    assign layer1_outputs[10031] = layer0_outputs[4519];
    assign layer1_outputs[10032] = ~(layer0_outputs[2108]);
    assign layer1_outputs[10033] = (layer0_outputs[3434]) & ~(layer0_outputs[11154]);
    assign layer1_outputs[10034] = 1'b1;
    assign layer1_outputs[10035] = 1'b1;
    assign layer1_outputs[10036] = (layer0_outputs[4223]) | (layer0_outputs[11853]);
    assign layer1_outputs[10037] = ~(layer0_outputs[8404]);
    assign layer1_outputs[10038] = layer0_outputs[2595];
    assign layer1_outputs[10039] = ~(layer0_outputs[11851]);
    assign layer1_outputs[10040] = ~((layer0_outputs[12758]) | (layer0_outputs[12119]));
    assign layer1_outputs[10041] = layer0_outputs[5063];
    assign layer1_outputs[10042] = ~(layer0_outputs[3357]) | (layer0_outputs[8311]);
    assign layer1_outputs[10043] = ~((layer0_outputs[12161]) | (layer0_outputs[7112]));
    assign layer1_outputs[10044] = 1'b0;
    assign layer1_outputs[10045] = ~(layer0_outputs[7036]);
    assign layer1_outputs[10046] = ~((layer0_outputs[676]) | (layer0_outputs[9102]));
    assign layer1_outputs[10047] = ~((layer0_outputs[8418]) ^ (layer0_outputs[5880]));
    assign layer1_outputs[10048] = ~(layer0_outputs[9425]) | (layer0_outputs[5983]);
    assign layer1_outputs[10049] = layer0_outputs[433];
    assign layer1_outputs[10050] = ~(layer0_outputs[8889]) | (layer0_outputs[8778]);
    assign layer1_outputs[10051] = ~((layer0_outputs[8182]) | (layer0_outputs[2567]));
    assign layer1_outputs[10052] = ~(layer0_outputs[9942]);
    assign layer1_outputs[10053] = ~(layer0_outputs[778]) | (layer0_outputs[11662]);
    assign layer1_outputs[10054] = (layer0_outputs[3629]) & ~(layer0_outputs[1155]);
    assign layer1_outputs[10055] = ~(layer0_outputs[10589]) | (layer0_outputs[4013]);
    assign layer1_outputs[10056] = ~(layer0_outputs[2423]);
    assign layer1_outputs[10057] = ~(layer0_outputs[6945]);
    assign layer1_outputs[10058] = 1'b0;
    assign layer1_outputs[10059] = ~(layer0_outputs[5855]) | (layer0_outputs[4757]);
    assign layer1_outputs[10060] = ~(layer0_outputs[3573]);
    assign layer1_outputs[10061] = (layer0_outputs[5407]) ^ (layer0_outputs[2199]);
    assign layer1_outputs[10062] = ~((layer0_outputs[7553]) & (layer0_outputs[7252]));
    assign layer1_outputs[10063] = ~(layer0_outputs[6809]);
    assign layer1_outputs[10064] = ~((layer0_outputs[8840]) | (layer0_outputs[3420]));
    assign layer1_outputs[10065] = layer0_outputs[7009];
    assign layer1_outputs[10066] = 1'b0;
    assign layer1_outputs[10067] = layer0_outputs[9347];
    assign layer1_outputs[10068] = layer0_outputs[1434];
    assign layer1_outputs[10069] = ~(layer0_outputs[4717]) | (layer0_outputs[3541]);
    assign layer1_outputs[10070] = ~((layer0_outputs[2191]) ^ (layer0_outputs[1765]));
    assign layer1_outputs[10071] = ~(layer0_outputs[5047]);
    assign layer1_outputs[10072] = ~((layer0_outputs[7875]) & (layer0_outputs[10170]));
    assign layer1_outputs[10073] = (layer0_outputs[625]) ^ (layer0_outputs[1485]);
    assign layer1_outputs[10074] = ~((layer0_outputs[2245]) & (layer0_outputs[6291]));
    assign layer1_outputs[10075] = ~((layer0_outputs[9559]) | (layer0_outputs[4806]));
    assign layer1_outputs[10076] = layer0_outputs[2391];
    assign layer1_outputs[10077] = ~((layer0_outputs[10159]) & (layer0_outputs[11812]));
    assign layer1_outputs[10078] = (layer0_outputs[2607]) & ~(layer0_outputs[7019]);
    assign layer1_outputs[10079] = layer0_outputs[3065];
    assign layer1_outputs[10080] = ~(layer0_outputs[5612]) | (layer0_outputs[7916]);
    assign layer1_outputs[10081] = (layer0_outputs[2364]) & (layer0_outputs[8240]);
    assign layer1_outputs[10082] = (layer0_outputs[7442]) & ~(layer0_outputs[9351]);
    assign layer1_outputs[10083] = ~(layer0_outputs[5131]);
    assign layer1_outputs[10084] = ~(layer0_outputs[10075]);
    assign layer1_outputs[10085] = ~(layer0_outputs[3753]) | (layer0_outputs[8768]);
    assign layer1_outputs[10086] = layer0_outputs[1906];
    assign layer1_outputs[10087] = ~(layer0_outputs[9074]) | (layer0_outputs[1303]);
    assign layer1_outputs[10088] = layer0_outputs[1128];
    assign layer1_outputs[10089] = layer0_outputs[12485];
    assign layer1_outputs[10090] = (layer0_outputs[12797]) & ~(layer0_outputs[4722]);
    assign layer1_outputs[10091] = (layer0_outputs[4930]) & (layer0_outputs[4613]);
    assign layer1_outputs[10092] = (layer0_outputs[843]) & ~(layer0_outputs[9494]);
    assign layer1_outputs[10093] = ~((layer0_outputs[5559]) | (layer0_outputs[701]));
    assign layer1_outputs[10094] = (layer0_outputs[5074]) ^ (layer0_outputs[1097]);
    assign layer1_outputs[10095] = ~(layer0_outputs[6698]);
    assign layer1_outputs[10096] = ~((layer0_outputs[12512]) & (layer0_outputs[6248]));
    assign layer1_outputs[10097] = ~(layer0_outputs[2662]) | (layer0_outputs[11338]);
    assign layer1_outputs[10098] = ~(layer0_outputs[12751]);
    assign layer1_outputs[10099] = (layer0_outputs[9138]) | (layer0_outputs[9158]);
    assign layer1_outputs[10100] = layer0_outputs[8545];
    assign layer1_outputs[10101] = (layer0_outputs[3506]) & ~(layer0_outputs[2724]);
    assign layer1_outputs[10102] = (layer0_outputs[9279]) & ~(layer0_outputs[6653]);
    assign layer1_outputs[10103] = ~((layer0_outputs[12618]) ^ (layer0_outputs[5321]));
    assign layer1_outputs[10104] = (layer0_outputs[1985]) & ~(layer0_outputs[7175]);
    assign layer1_outputs[10105] = layer0_outputs[4372];
    assign layer1_outputs[10106] = (layer0_outputs[1759]) & ~(layer0_outputs[10316]);
    assign layer1_outputs[10107] = ~((layer0_outputs[1578]) | (layer0_outputs[11945]));
    assign layer1_outputs[10108] = ~((layer0_outputs[7936]) ^ (layer0_outputs[12533]));
    assign layer1_outputs[10109] = ~(layer0_outputs[10497]);
    assign layer1_outputs[10110] = ~(layer0_outputs[9563]) | (layer0_outputs[182]);
    assign layer1_outputs[10111] = (layer0_outputs[7648]) ^ (layer0_outputs[8477]);
    assign layer1_outputs[10112] = (layer0_outputs[11781]) & (layer0_outputs[1696]);
    assign layer1_outputs[10113] = ~((layer0_outputs[10364]) & (layer0_outputs[11736]));
    assign layer1_outputs[10114] = ~(layer0_outputs[694]);
    assign layer1_outputs[10115] = ~(layer0_outputs[59]);
    assign layer1_outputs[10116] = (layer0_outputs[167]) ^ (layer0_outputs[9631]);
    assign layer1_outputs[10117] = ~((layer0_outputs[1629]) | (layer0_outputs[7243]));
    assign layer1_outputs[10118] = ~(layer0_outputs[3710]);
    assign layer1_outputs[10119] = (layer0_outputs[148]) & ~(layer0_outputs[6520]);
    assign layer1_outputs[10120] = ~(layer0_outputs[7952]);
    assign layer1_outputs[10121] = ~(layer0_outputs[1277]);
    assign layer1_outputs[10122] = 1'b1;
    assign layer1_outputs[10123] = ~((layer0_outputs[10957]) ^ (layer0_outputs[11170]));
    assign layer1_outputs[10124] = layer0_outputs[2874];
    assign layer1_outputs[10125] = layer0_outputs[6955];
    assign layer1_outputs[10126] = ~(layer0_outputs[6648]);
    assign layer1_outputs[10127] = (layer0_outputs[7704]) & ~(layer0_outputs[1330]);
    assign layer1_outputs[10128] = ~(layer0_outputs[12109]) | (layer0_outputs[9173]);
    assign layer1_outputs[10129] = ~((layer0_outputs[8159]) | (layer0_outputs[8438]));
    assign layer1_outputs[10130] = layer0_outputs[2168];
    assign layer1_outputs[10131] = ~((layer0_outputs[4171]) & (layer0_outputs[3623]));
    assign layer1_outputs[10132] = ~(layer0_outputs[11337]);
    assign layer1_outputs[10133] = ~((layer0_outputs[9180]) | (layer0_outputs[9397]));
    assign layer1_outputs[10134] = (layer0_outputs[7151]) & ~(layer0_outputs[2457]);
    assign layer1_outputs[10135] = ~((layer0_outputs[11605]) & (layer0_outputs[6865]));
    assign layer1_outputs[10136] = ~((layer0_outputs[10019]) & (layer0_outputs[5020]));
    assign layer1_outputs[10137] = (layer0_outputs[5830]) & ~(layer0_outputs[8035]);
    assign layer1_outputs[10138] = ~(layer0_outputs[1782]);
    assign layer1_outputs[10139] = (layer0_outputs[11527]) & ~(layer0_outputs[11720]);
    assign layer1_outputs[10140] = layer0_outputs[7487];
    assign layer1_outputs[10141] = layer0_outputs[4958];
    assign layer1_outputs[10142] = ~((layer0_outputs[10001]) | (layer0_outputs[4983]));
    assign layer1_outputs[10143] = ~(layer0_outputs[3088]);
    assign layer1_outputs[10144] = ~(layer0_outputs[3694]);
    assign layer1_outputs[10145] = layer0_outputs[6080];
    assign layer1_outputs[10146] = layer0_outputs[4188];
    assign layer1_outputs[10147] = (layer0_outputs[6094]) ^ (layer0_outputs[4865]);
    assign layer1_outputs[10148] = ~(layer0_outputs[6276]);
    assign layer1_outputs[10149] = ~(layer0_outputs[4700]);
    assign layer1_outputs[10150] = ~((layer0_outputs[1570]) & (layer0_outputs[11518]));
    assign layer1_outputs[10151] = ~(layer0_outputs[4781]);
    assign layer1_outputs[10152] = (layer0_outputs[7144]) ^ (layer0_outputs[264]);
    assign layer1_outputs[10153] = (layer0_outputs[11203]) ^ (layer0_outputs[2784]);
    assign layer1_outputs[10154] = ~((layer0_outputs[603]) | (layer0_outputs[10616]));
    assign layer1_outputs[10155] = ~((layer0_outputs[582]) & (layer0_outputs[7560]));
    assign layer1_outputs[10156] = layer0_outputs[4338];
    assign layer1_outputs[10157] = ~((layer0_outputs[12227]) ^ (layer0_outputs[855]));
    assign layer1_outputs[10158] = layer0_outputs[8964];
    assign layer1_outputs[10159] = (layer0_outputs[5179]) ^ (layer0_outputs[9790]);
    assign layer1_outputs[10160] = (layer0_outputs[2565]) | (layer0_outputs[6334]);
    assign layer1_outputs[10161] = ~((layer0_outputs[6233]) ^ (layer0_outputs[3556]));
    assign layer1_outputs[10162] = ~((layer0_outputs[11119]) & (layer0_outputs[2137]));
    assign layer1_outputs[10163] = layer0_outputs[8155];
    assign layer1_outputs[10164] = ~(layer0_outputs[7887]);
    assign layer1_outputs[10165] = (layer0_outputs[6881]) & ~(layer0_outputs[11968]);
    assign layer1_outputs[10166] = ~(layer0_outputs[4460]);
    assign layer1_outputs[10167] = ~(layer0_outputs[632]);
    assign layer1_outputs[10168] = layer0_outputs[11987];
    assign layer1_outputs[10169] = ~((layer0_outputs[4388]) & (layer0_outputs[3178]));
    assign layer1_outputs[10170] = layer0_outputs[3278];
    assign layer1_outputs[10171] = ~(layer0_outputs[11802]) | (layer0_outputs[12377]);
    assign layer1_outputs[10172] = layer0_outputs[7556];
    assign layer1_outputs[10173] = ~((layer0_outputs[9506]) | (layer0_outputs[6073]));
    assign layer1_outputs[10174] = layer0_outputs[11533];
    assign layer1_outputs[10175] = (layer0_outputs[3565]) | (layer0_outputs[6072]);
    assign layer1_outputs[10176] = (layer0_outputs[6132]) | (layer0_outputs[1628]);
    assign layer1_outputs[10177] = layer0_outputs[4442];
    assign layer1_outputs[10178] = ~((layer0_outputs[6058]) & (layer0_outputs[7229]));
    assign layer1_outputs[10179] = layer0_outputs[8859];
    assign layer1_outputs[10180] = ~((layer0_outputs[946]) & (layer0_outputs[7319]));
    assign layer1_outputs[10181] = (layer0_outputs[11577]) & ~(layer0_outputs[11491]);
    assign layer1_outputs[10182] = layer0_outputs[3412];
    assign layer1_outputs[10183] = (layer0_outputs[12007]) & ~(layer0_outputs[11369]);
    assign layer1_outputs[10184] = (layer0_outputs[412]) & (layer0_outputs[306]);
    assign layer1_outputs[10185] = ~(layer0_outputs[8971]) | (layer0_outputs[4141]);
    assign layer1_outputs[10186] = (layer0_outputs[5404]) ^ (layer0_outputs[10333]);
    assign layer1_outputs[10187] = ~(layer0_outputs[2833]);
    assign layer1_outputs[10188] = layer0_outputs[6764];
    assign layer1_outputs[10189] = (layer0_outputs[9093]) ^ (layer0_outputs[702]);
    assign layer1_outputs[10190] = (layer0_outputs[11491]) | (layer0_outputs[7399]);
    assign layer1_outputs[10191] = (layer0_outputs[6109]) & ~(layer0_outputs[7553]);
    assign layer1_outputs[10192] = ~((layer0_outputs[42]) & (layer0_outputs[7060]));
    assign layer1_outputs[10193] = ~(layer0_outputs[6028]) | (layer0_outputs[12726]);
    assign layer1_outputs[10194] = ~(layer0_outputs[156]);
    assign layer1_outputs[10195] = (layer0_outputs[7551]) & (layer0_outputs[9007]);
    assign layer1_outputs[10196] = layer0_outputs[4685];
    assign layer1_outputs[10197] = ~((layer0_outputs[4712]) & (layer0_outputs[1176]));
    assign layer1_outputs[10198] = (layer0_outputs[11708]) | (layer0_outputs[2539]);
    assign layer1_outputs[10199] = ~((layer0_outputs[2455]) ^ (layer0_outputs[4977]));
    assign layer1_outputs[10200] = ~(layer0_outputs[6153]);
    assign layer1_outputs[10201] = layer0_outputs[7872];
    assign layer1_outputs[10202] = (layer0_outputs[6022]) & (layer0_outputs[2763]);
    assign layer1_outputs[10203] = (layer0_outputs[126]) & ~(layer0_outputs[9062]);
    assign layer1_outputs[10204] = (layer0_outputs[7291]) & ~(layer0_outputs[692]);
    assign layer1_outputs[10205] = layer0_outputs[139];
    assign layer1_outputs[10206] = layer0_outputs[2317];
    assign layer1_outputs[10207] = ~(layer0_outputs[5655]);
    assign layer1_outputs[10208] = layer0_outputs[10205];
    assign layer1_outputs[10209] = 1'b1;
    assign layer1_outputs[10210] = ~((layer0_outputs[6225]) | (layer0_outputs[4765]));
    assign layer1_outputs[10211] = layer0_outputs[3726];
    assign layer1_outputs[10212] = 1'b1;
    assign layer1_outputs[10213] = (layer0_outputs[10249]) & ~(layer0_outputs[7550]);
    assign layer1_outputs[10214] = ~(layer0_outputs[9722]) | (layer0_outputs[8008]);
    assign layer1_outputs[10215] = ~(layer0_outputs[3824]);
    assign layer1_outputs[10216] = ~(layer0_outputs[7602]);
    assign layer1_outputs[10217] = (layer0_outputs[5438]) & (layer0_outputs[11169]);
    assign layer1_outputs[10218] = ~((layer0_outputs[687]) & (layer0_outputs[6386]));
    assign layer1_outputs[10219] = ~(layer0_outputs[7432]);
    assign layer1_outputs[10220] = layer0_outputs[12737];
    assign layer1_outputs[10221] = (layer0_outputs[4361]) | (layer0_outputs[10857]);
    assign layer1_outputs[10222] = layer0_outputs[490];
    assign layer1_outputs[10223] = ~(layer0_outputs[2015]);
    assign layer1_outputs[10224] = (layer0_outputs[4228]) ^ (layer0_outputs[3633]);
    assign layer1_outputs[10225] = (layer0_outputs[5985]) & ~(layer0_outputs[500]);
    assign layer1_outputs[10226] = (layer0_outputs[2630]) & ~(layer0_outputs[1130]);
    assign layer1_outputs[10227] = 1'b0;
    assign layer1_outputs[10228] = ~(layer0_outputs[9865]) | (layer0_outputs[861]);
    assign layer1_outputs[10229] = (layer0_outputs[2853]) ^ (layer0_outputs[8722]);
    assign layer1_outputs[10230] = ~(layer0_outputs[7377]) | (layer0_outputs[7004]);
    assign layer1_outputs[10231] = (layer0_outputs[5126]) & ~(layer0_outputs[10]);
    assign layer1_outputs[10232] = layer0_outputs[11657];
    assign layer1_outputs[10233] = ~(layer0_outputs[12582]) | (layer0_outputs[4696]);
    assign layer1_outputs[10234] = ~((layer0_outputs[11675]) | (layer0_outputs[3600]));
    assign layer1_outputs[10235] = ~((layer0_outputs[6110]) ^ (layer0_outputs[11454]));
    assign layer1_outputs[10236] = (layer0_outputs[2905]) ^ (layer0_outputs[4817]);
    assign layer1_outputs[10237] = ~(layer0_outputs[11346]);
    assign layer1_outputs[10238] = layer0_outputs[1468];
    assign layer1_outputs[10239] = ~(layer0_outputs[9284]);
    assign layer1_outputs[10240] = (layer0_outputs[5781]) & ~(layer0_outputs[11145]);
    assign layer1_outputs[10241] = layer0_outputs[12076];
    assign layer1_outputs[10242] = ~(layer0_outputs[3377]);
    assign layer1_outputs[10243] = ~(layer0_outputs[1311]) | (layer0_outputs[5688]);
    assign layer1_outputs[10244] = (layer0_outputs[1362]) & (layer0_outputs[11784]);
    assign layer1_outputs[10245] = layer0_outputs[12327];
    assign layer1_outputs[10246] = ~((layer0_outputs[5414]) | (layer0_outputs[851]));
    assign layer1_outputs[10247] = ~((layer0_outputs[8006]) ^ (layer0_outputs[3986]));
    assign layer1_outputs[10248] = (layer0_outputs[1086]) & ~(layer0_outputs[6372]);
    assign layer1_outputs[10249] = layer0_outputs[6266];
    assign layer1_outputs[10250] = (layer0_outputs[6512]) ^ (layer0_outputs[5957]);
    assign layer1_outputs[10251] = ~(layer0_outputs[3550]);
    assign layer1_outputs[10252] = ~((layer0_outputs[2411]) | (layer0_outputs[8619]));
    assign layer1_outputs[10253] = ~(layer0_outputs[6148]);
    assign layer1_outputs[10254] = ~(layer0_outputs[7748]);
    assign layer1_outputs[10255] = ~(layer0_outputs[10310]) | (layer0_outputs[9589]);
    assign layer1_outputs[10256] = ~((layer0_outputs[4421]) | (layer0_outputs[1019]));
    assign layer1_outputs[10257] = layer0_outputs[8712];
    assign layer1_outputs[10258] = ~(layer0_outputs[8574]) | (layer0_outputs[10935]);
    assign layer1_outputs[10259] = (layer0_outputs[3648]) & ~(layer0_outputs[1934]);
    assign layer1_outputs[10260] = ~(layer0_outputs[8554]);
    assign layer1_outputs[10261] = ~(layer0_outputs[3655]);
    assign layer1_outputs[10262] = (layer0_outputs[9958]) & ~(layer0_outputs[9528]);
    assign layer1_outputs[10263] = ~(layer0_outputs[9496]);
    assign layer1_outputs[10264] = (layer0_outputs[10874]) & ~(layer0_outputs[11687]);
    assign layer1_outputs[10265] = ~(layer0_outputs[1011]);
    assign layer1_outputs[10266] = (layer0_outputs[10264]) & ~(layer0_outputs[12369]);
    assign layer1_outputs[10267] = ~(layer0_outputs[1693]);
    assign layer1_outputs[10268] = ~((layer0_outputs[1837]) ^ (layer0_outputs[10587]));
    assign layer1_outputs[10269] = ~(layer0_outputs[703]);
    assign layer1_outputs[10270] = (layer0_outputs[5747]) & (layer0_outputs[2515]);
    assign layer1_outputs[10271] = (layer0_outputs[348]) | (layer0_outputs[6644]);
    assign layer1_outputs[10272] = ~(layer0_outputs[12252]);
    assign layer1_outputs[10273] = ~((layer0_outputs[8103]) & (layer0_outputs[2938]));
    assign layer1_outputs[10274] = ~(layer0_outputs[10465]) | (layer0_outputs[12073]);
    assign layer1_outputs[10275] = ~(layer0_outputs[4976]) | (layer0_outputs[4809]);
    assign layer1_outputs[10276] = 1'b1;
    assign layer1_outputs[10277] = (layer0_outputs[3871]) & ~(layer0_outputs[9988]);
    assign layer1_outputs[10278] = (layer0_outputs[7141]) & ~(layer0_outputs[5946]);
    assign layer1_outputs[10279] = ~((layer0_outputs[2243]) ^ (layer0_outputs[8749]));
    assign layer1_outputs[10280] = ~((layer0_outputs[10918]) & (layer0_outputs[11914]));
    assign layer1_outputs[10281] = (layer0_outputs[3891]) ^ (layer0_outputs[4227]);
    assign layer1_outputs[10282] = ~((layer0_outputs[11233]) ^ (layer0_outputs[2479]));
    assign layer1_outputs[10283] = layer0_outputs[7301];
    assign layer1_outputs[10284] = layer0_outputs[12551];
    assign layer1_outputs[10285] = layer0_outputs[3920];
    assign layer1_outputs[10286] = ~((layer0_outputs[8819]) | (layer0_outputs[6008]));
    assign layer1_outputs[10287] = (layer0_outputs[10626]) & ~(layer0_outputs[8491]);
    assign layer1_outputs[10288] = ~(layer0_outputs[6589]);
    assign layer1_outputs[10289] = ~((layer0_outputs[5990]) & (layer0_outputs[12674]));
    assign layer1_outputs[10290] = ~((layer0_outputs[7359]) ^ (layer0_outputs[7011]));
    assign layer1_outputs[10291] = (layer0_outputs[10926]) & ~(layer0_outputs[5189]);
    assign layer1_outputs[10292] = ~(layer0_outputs[6555]) | (layer0_outputs[2286]);
    assign layer1_outputs[10293] = (layer0_outputs[9444]) ^ (layer0_outputs[7361]);
    assign layer1_outputs[10294] = 1'b1;
    assign layer1_outputs[10295] = ~((layer0_outputs[7751]) | (layer0_outputs[1932]));
    assign layer1_outputs[10296] = ~((layer0_outputs[2032]) & (layer0_outputs[3208]));
    assign layer1_outputs[10297] = layer0_outputs[2167];
    assign layer1_outputs[10298] = layer0_outputs[8055];
    assign layer1_outputs[10299] = ~(layer0_outputs[1607]);
    assign layer1_outputs[10300] = (layer0_outputs[4476]) & ~(layer0_outputs[3027]);
    assign layer1_outputs[10301] = ~(layer0_outputs[11235]);
    assign layer1_outputs[10302] = ~((layer0_outputs[1813]) ^ (layer0_outputs[8533]));
    assign layer1_outputs[10303] = ~(layer0_outputs[9337]);
    assign layer1_outputs[10304] = layer0_outputs[10502];
    assign layer1_outputs[10305] = ~((layer0_outputs[2389]) | (layer0_outputs[844]));
    assign layer1_outputs[10306] = 1'b0;
    assign layer1_outputs[10307] = ~(layer0_outputs[61]);
    assign layer1_outputs[10308] = ~((layer0_outputs[4863]) & (layer0_outputs[2871]));
    assign layer1_outputs[10309] = ~(layer0_outputs[9367]);
    assign layer1_outputs[10310] = layer0_outputs[1646];
    assign layer1_outputs[10311] = ~((layer0_outputs[6814]) ^ (layer0_outputs[10700]));
    assign layer1_outputs[10312] = (layer0_outputs[10865]) & (layer0_outputs[196]);
    assign layer1_outputs[10313] = layer0_outputs[4737];
    assign layer1_outputs[10314] = ~(layer0_outputs[11928]);
    assign layer1_outputs[10315] = ~(layer0_outputs[5319]);
    assign layer1_outputs[10316] = (layer0_outputs[6214]) | (layer0_outputs[462]);
    assign layer1_outputs[10317] = ~(layer0_outputs[1331]) | (layer0_outputs[7875]);
    assign layer1_outputs[10318] = (layer0_outputs[658]) & ~(layer0_outputs[7125]);
    assign layer1_outputs[10319] = (layer0_outputs[329]) ^ (layer0_outputs[3453]);
    assign layer1_outputs[10320] = ~(layer0_outputs[4730]);
    assign layer1_outputs[10321] = (layer0_outputs[12475]) & (layer0_outputs[11166]);
    assign layer1_outputs[10322] = layer0_outputs[10969];
    assign layer1_outputs[10323] = ~(layer0_outputs[788]);
    assign layer1_outputs[10324] = (layer0_outputs[4741]) & ~(layer0_outputs[5750]);
    assign layer1_outputs[10325] = (layer0_outputs[12324]) & ~(layer0_outputs[10739]);
    assign layer1_outputs[10326] = layer0_outputs[379];
    assign layer1_outputs[10327] = layer0_outputs[7818];
    assign layer1_outputs[10328] = (layer0_outputs[4142]) & ~(layer0_outputs[6713]);
    assign layer1_outputs[10329] = (layer0_outputs[11503]) & (layer0_outputs[5206]);
    assign layer1_outputs[10330] = ~(layer0_outputs[7346]);
    assign layer1_outputs[10331] = ~(layer0_outputs[7961]);
    assign layer1_outputs[10332] = ~((layer0_outputs[10653]) ^ (layer0_outputs[11546]));
    assign layer1_outputs[10333] = ~((layer0_outputs[9072]) ^ (layer0_outputs[639]));
    assign layer1_outputs[10334] = ~((layer0_outputs[9297]) ^ (layer0_outputs[11213]));
    assign layer1_outputs[10335] = ~(layer0_outputs[3816]) | (layer0_outputs[12426]);
    assign layer1_outputs[10336] = layer0_outputs[8092];
    assign layer1_outputs[10337] = (layer0_outputs[6811]) & ~(layer0_outputs[1523]);
    assign layer1_outputs[10338] = (layer0_outputs[11405]) | (layer0_outputs[10308]);
    assign layer1_outputs[10339] = (layer0_outputs[285]) & ~(layer0_outputs[5695]);
    assign layer1_outputs[10340] = layer0_outputs[7851];
    assign layer1_outputs[10341] = ~(layer0_outputs[1472]) | (layer0_outputs[1476]);
    assign layer1_outputs[10342] = layer0_outputs[3446];
    assign layer1_outputs[10343] = (layer0_outputs[6465]) | (layer0_outputs[8378]);
    assign layer1_outputs[10344] = (layer0_outputs[1233]) & (layer0_outputs[8862]);
    assign layer1_outputs[10345] = ~((layer0_outputs[674]) | (layer0_outputs[7948]));
    assign layer1_outputs[10346] = ~(layer0_outputs[10672]);
    assign layer1_outputs[10347] = (layer0_outputs[9746]) ^ (layer0_outputs[2149]);
    assign layer1_outputs[10348] = layer0_outputs[7512];
    assign layer1_outputs[10349] = ~(layer0_outputs[12311]) | (layer0_outputs[3971]);
    assign layer1_outputs[10350] = (layer0_outputs[8218]) & ~(layer0_outputs[3233]);
    assign layer1_outputs[10351] = ~(layer0_outputs[6936]);
    assign layer1_outputs[10352] = ~(layer0_outputs[10617]);
    assign layer1_outputs[10353] = (layer0_outputs[4375]) & ~(layer0_outputs[8698]);
    assign layer1_outputs[10354] = ~(layer0_outputs[12228]) | (layer0_outputs[7469]);
    assign layer1_outputs[10355] = layer0_outputs[729];
    assign layer1_outputs[10356] = ~(layer0_outputs[9492]) | (layer0_outputs[7247]);
    assign layer1_outputs[10357] = (layer0_outputs[1217]) ^ (layer0_outputs[4604]);
    assign layer1_outputs[10358] = layer0_outputs[7472];
    assign layer1_outputs[10359] = layer0_outputs[802];
    assign layer1_outputs[10360] = ~(layer0_outputs[2065]) | (layer0_outputs[3310]);
    assign layer1_outputs[10361] = (layer0_outputs[3929]) ^ (layer0_outputs[2203]);
    assign layer1_outputs[10362] = layer0_outputs[9083];
    assign layer1_outputs[10363] = (layer0_outputs[3959]) & (layer0_outputs[10725]);
    assign layer1_outputs[10364] = (layer0_outputs[11005]) & (layer0_outputs[180]);
    assign layer1_outputs[10365] = 1'b0;
    assign layer1_outputs[10366] = (layer0_outputs[2958]) & (layer0_outputs[2672]);
    assign layer1_outputs[10367] = layer0_outputs[4582];
    assign layer1_outputs[10368] = (layer0_outputs[2725]) ^ (layer0_outputs[10772]);
    assign layer1_outputs[10369] = ~(layer0_outputs[5611]) | (layer0_outputs[7663]);
    assign layer1_outputs[10370] = ~(layer0_outputs[6793]);
    assign layer1_outputs[10371] = layer0_outputs[9338];
    assign layer1_outputs[10372] = ~((layer0_outputs[187]) & (layer0_outputs[1170]));
    assign layer1_outputs[10373] = layer0_outputs[10172];
    assign layer1_outputs[10374] = 1'b0;
    assign layer1_outputs[10375] = (layer0_outputs[11586]) ^ (layer0_outputs[263]);
    assign layer1_outputs[10376] = ~(layer0_outputs[892]) | (layer0_outputs[1704]);
    assign layer1_outputs[10377] = (layer0_outputs[6625]) & ~(layer0_outputs[9837]);
    assign layer1_outputs[10378] = ~(layer0_outputs[10663]);
    assign layer1_outputs[10379] = layer0_outputs[1740];
    assign layer1_outputs[10380] = ~((layer0_outputs[6066]) | (layer0_outputs[7671]));
    assign layer1_outputs[10381] = ~(layer0_outputs[7111]) | (layer0_outputs[9217]);
    assign layer1_outputs[10382] = layer0_outputs[1757];
    assign layer1_outputs[10383] = 1'b0;
    assign layer1_outputs[10384] = ~(layer0_outputs[12384]);
    assign layer1_outputs[10385] = ~(layer0_outputs[8960]);
    assign layer1_outputs[10386] = ~((layer0_outputs[10051]) | (layer0_outputs[12783]));
    assign layer1_outputs[10387] = layer0_outputs[685];
    assign layer1_outputs[10388] = layer0_outputs[3384];
    assign layer1_outputs[10389] = (layer0_outputs[10276]) & ~(layer0_outputs[1853]);
    assign layer1_outputs[10390] = (layer0_outputs[1604]) & ~(layer0_outputs[4498]);
    assign layer1_outputs[10391] = layer0_outputs[2283];
    assign layer1_outputs[10392] = (layer0_outputs[6137]) | (layer0_outputs[631]);
    assign layer1_outputs[10393] = (layer0_outputs[7749]) ^ (layer0_outputs[3710]);
    assign layer1_outputs[10394] = (layer0_outputs[1433]) & (layer0_outputs[3563]);
    assign layer1_outputs[10395] = ~(layer0_outputs[576]) | (layer0_outputs[10678]);
    assign layer1_outputs[10396] = (layer0_outputs[4283]) ^ (layer0_outputs[739]);
    assign layer1_outputs[10397] = (layer0_outputs[5867]) & ~(layer0_outputs[4278]);
    assign layer1_outputs[10398] = (layer0_outputs[5246]) | (layer0_outputs[12681]);
    assign layer1_outputs[10399] = layer0_outputs[9820];
    assign layer1_outputs[10400] = ~(layer0_outputs[4977]);
    assign layer1_outputs[10401] = (layer0_outputs[10033]) & (layer0_outputs[12337]);
    assign layer1_outputs[10402] = ~(layer0_outputs[9001]) | (layer0_outputs[7179]);
    assign layer1_outputs[10403] = ~(layer0_outputs[2829]) | (layer0_outputs[12618]);
    assign layer1_outputs[10404] = ~((layer0_outputs[11935]) ^ (layer0_outputs[10541]));
    assign layer1_outputs[10405] = (layer0_outputs[2741]) ^ (layer0_outputs[10197]);
    assign layer1_outputs[10406] = (layer0_outputs[12279]) | (layer0_outputs[3522]);
    assign layer1_outputs[10407] = ~(layer0_outputs[4466]) | (layer0_outputs[9750]);
    assign layer1_outputs[10408] = ~(layer0_outputs[10297]);
    assign layer1_outputs[10409] = (layer0_outputs[4788]) | (layer0_outputs[10935]);
    assign layer1_outputs[10410] = ~(layer0_outputs[4374]);
    assign layer1_outputs[10411] = (layer0_outputs[10328]) & ~(layer0_outputs[6971]);
    assign layer1_outputs[10412] = ~(layer0_outputs[11548]);
    assign layer1_outputs[10413] = ~(layer0_outputs[6917]) | (layer0_outputs[7664]);
    assign layer1_outputs[10414] = ~((layer0_outputs[11375]) & (layer0_outputs[3769]));
    assign layer1_outputs[10415] = (layer0_outputs[6093]) & ~(layer0_outputs[10637]);
    assign layer1_outputs[10416] = layer0_outputs[5346];
    assign layer1_outputs[10417] = ~((layer0_outputs[2258]) | (layer0_outputs[11337]));
    assign layer1_outputs[10418] = (layer0_outputs[12581]) ^ (layer0_outputs[12179]);
    assign layer1_outputs[10419] = ~(layer0_outputs[3236]) | (layer0_outputs[5698]);
    assign layer1_outputs[10420] = (layer0_outputs[9673]) & ~(layer0_outputs[3928]);
    assign layer1_outputs[10421] = layer0_outputs[3427];
    assign layer1_outputs[10422] = (layer0_outputs[1487]) & ~(layer0_outputs[12684]);
    assign layer1_outputs[10423] = ~((layer0_outputs[3294]) | (layer0_outputs[1260]));
    assign layer1_outputs[10424] = (layer0_outputs[5779]) ^ (layer0_outputs[7023]);
    assign layer1_outputs[10425] = ~(layer0_outputs[1155]) | (layer0_outputs[4546]);
    assign layer1_outputs[10426] = layer0_outputs[13];
    assign layer1_outputs[10427] = ~((layer0_outputs[4230]) | (layer0_outputs[7902]));
    assign layer1_outputs[10428] = ~(layer0_outputs[8175]);
    assign layer1_outputs[10429] = ~(layer0_outputs[11004]) | (layer0_outputs[2791]);
    assign layer1_outputs[10430] = ~(layer0_outputs[4758]) | (layer0_outputs[10070]);
    assign layer1_outputs[10431] = ~(layer0_outputs[5160]) | (layer0_outputs[7509]);
    assign layer1_outputs[10432] = (layer0_outputs[3474]) | (layer0_outputs[3022]);
    assign layer1_outputs[10433] = layer0_outputs[11689];
    assign layer1_outputs[10434] = ~((layer0_outputs[8292]) | (layer0_outputs[11589]));
    assign layer1_outputs[10435] = layer0_outputs[11406];
    assign layer1_outputs[10436] = ~(layer0_outputs[5764]);
    assign layer1_outputs[10437] = ~(layer0_outputs[2974]);
    assign layer1_outputs[10438] = ~(layer0_outputs[4940]);
    assign layer1_outputs[10439] = (layer0_outputs[10231]) | (layer0_outputs[7706]);
    assign layer1_outputs[10440] = ~((layer0_outputs[12178]) | (layer0_outputs[9573]));
    assign layer1_outputs[10441] = (layer0_outputs[4326]) & ~(layer0_outputs[2413]);
    assign layer1_outputs[10442] = layer0_outputs[10216];
    assign layer1_outputs[10443] = layer0_outputs[4561];
    assign layer1_outputs[10444] = ~(layer0_outputs[5178]) | (layer0_outputs[10184]);
    assign layer1_outputs[10445] = layer0_outputs[5022];
    assign layer1_outputs[10446] = layer0_outputs[2994];
    assign layer1_outputs[10447] = layer0_outputs[2887];
    assign layer1_outputs[10448] = ~((layer0_outputs[2342]) | (layer0_outputs[9010]));
    assign layer1_outputs[10449] = ~((layer0_outputs[5927]) | (layer0_outputs[5959]));
    assign layer1_outputs[10450] = 1'b0;
    assign layer1_outputs[10451] = (layer0_outputs[6841]) & (layer0_outputs[4494]);
    assign layer1_outputs[10452] = ~(layer0_outputs[231]);
    assign layer1_outputs[10453] = ~(layer0_outputs[9840]);
    assign layer1_outputs[10454] = (layer0_outputs[10553]) & ~(layer0_outputs[394]);
    assign layer1_outputs[10455] = ~(layer0_outputs[1492]) | (layer0_outputs[3348]);
    assign layer1_outputs[10456] = layer0_outputs[6176];
    assign layer1_outputs[10457] = ~(layer0_outputs[10466]) | (layer0_outputs[2052]);
    assign layer1_outputs[10458] = (layer0_outputs[2876]) | (layer0_outputs[1710]);
    assign layer1_outputs[10459] = ~(layer0_outputs[7319]);
    assign layer1_outputs[10460] = (layer0_outputs[12374]) & (layer0_outputs[1495]);
    assign layer1_outputs[10461] = (layer0_outputs[6912]) & ~(layer0_outputs[4877]);
    assign layer1_outputs[10462] = ~(layer0_outputs[6299]);
    assign layer1_outputs[10463] = layer0_outputs[8063];
    assign layer1_outputs[10464] = (layer0_outputs[9265]) ^ (layer0_outputs[9320]);
    assign layer1_outputs[10465] = ~((layer0_outputs[8833]) & (layer0_outputs[4253]));
    assign layer1_outputs[10466] = (layer0_outputs[3216]) | (layer0_outputs[8511]);
    assign layer1_outputs[10467] = (layer0_outputs[7578]) & ~(layer0_outputs[8370]);
    assign layer1_outputs[10468] = ~(layer0_outputs[7786]) | (layer0_outputs[10370]);
    assign layer1_outputs[10469] = ~((layer0_outputs[3465]) | (layer0_outputs[6629]));
    assign layer1_outputs[10470] = ~(layer0_outputs[9438]) | (layer0_outputs[8650]);
    assign layer1_outputs[10471] = layer0_outputs[247];
    assign layer1_outputs[10472] = ~(layer0_outputs[6394]);
    assign layer1_outputs[10473] = layer0_outputs[11854];
    assign layer1_outputs[10474] = layer0_outputs[10951];
    assign layer1_outputs[10475] = layer0_outputs[1662];
    assign layer1_outputs[10476] = layer0_outputs[11500];
    assign layer1_outputs[10477] = ~(layer0_outputs[8411]);
    assign layer1_outputs[10478] = 1'b0;
    assign layer1_outputs[10479] = ~((layer0_outputs[8107]) | (layer0_outputs[11247]));
    assign layer1_outputs[10480] = (layer0_outputs[2816]) & ~(layer0_outputs[9472]);
    assign layer1_outputs[10481] = 1'b0;
    assign layer1_outputs[10482] = layer0_outputs[8759];
    assign layer1_outputs[10483] = layer0_outputs[7254];
    assign layer1_outputs[10484] = (layer0_outputs[2218]) & (layer0_outputs[2908]);
    assign layer1_outputs[10485] = ~(layer0_outputs[12749]) | (layer0_outputs[8277]);
    assign layer1_outputs[10486] = ~((layer0_outputs[8014]) & (layer0_outputs[5929]));
    assign layer1_outputs[10487] = ~(layer0_outputs[11220]);
    assign layer1_outputs[10488] = ~(layer0_outputs[8461]);
    assign layer1_outputs[10489] = (layer0_outputs[172]) & ~(layer0_outputs[1966]);
    assign layer1_outputs[10490] = ~((layer0_outputs[485]) ^ (layer0_outputs[6755]));
    assign layer1_outputs[10491] = ~(layer0_outputs[600]) | (layer0_outputs[4705]);
    assign layer1_outputs[10492] = ~((layer0_outputs[577]) ^ (layer0_outputs[6002]));
    assign layer1_outputs[10493] = (layer0_outputs[5598]) ^ (layer0_outputs[9076]);
    assign layer1_outputs[10494] = ~(layer0_outputs[1538]);
    assign layer1_outputs[10495] = ~(layer0_outputs[1419]) | (layer0_outputs[10329]);
    assign layer1_outputs[10496] = ~(layer0_outputs[4177]);
    assign layer1_outputs[10497] = ~((layer0_outputs[11607]) | (layer0_outputs[3436]));
    assign layer1_outputs[10498] = ~(layer0_outputs[1563]);
    assign layer1_outputs[10499] = ~(layer0_outputs[675]) | (layer0_outputs[4384]);
    assign layer1_outputs[10500] = layer0_outputs[5576];
    assign layer1_outputs[10501] = ~(layer0_outputs[9035]);
    assign layer1_outputs[10502] = ~(layer0_outputs[6020]);
    assign layer1_outputs[10503] = ~(layer0_outputs[6453]) | (layer0_outputs[3657]);
    assign layer1_outputs[10504] = (layer0_outputs[2636]) & ~(layer0_outputs[5064]);
    assign layer1_outputs[10505] = ~(layer0_outputs[2043]);
    assign layer1_outputs[10506] = layer0_outputs[9937];
    assign layer1_outputs[10507] = (layer0_outputs[3737]) | (layer0_outputs[2466]);
    assign layer1_outputs[10508] = ~(layer0_outputs[7588]);
    assign layer1_outputs[10509] = layer0_outputs[6561];
    assign layer1_outputs[10510] = (layer0_outputs[7518]) & (layer0_outputs[563]);
    assign layer1_outputs[10511] = ~((layer0_outputs[7527]) | (layer0_outputs[2660]));
    assign layer1_outputs[10512] = 1'b1;
    assign layer1_outputs[10513] = (layer0_outputs[4982]) & ~(layer0_outputs[8266]);
    assign layer1_outputs[10514] = (layer0_outputs[5462]) & (layer0_outputs[6341]);
    assign layer1_outputs[10515] = ~(layer0_outputs[268]);
    assign layer1_outputs[10516] = ~(layer0_outputs[3201]) | (layer0_outputs[5247]);
    assign layer1_outputs[10517] = ~((layer0_outputs[7919]) | (layer0_outputs[1559]));
    assign layer1_outputs[10518] = (layer0_outputs[2334]) & ~(layer0_outputs[4437]);
    assign layer1_outputs[10519] = ~(layer0_outputs[2061]) | (layer0_outputs[9440]);
    assign layer1_outputs[10520] = ~(layer0_outputs[5819]);
    assign layer1_outputs[10521] = ~((layer0_outputs[11174]) & (layer0_outputs[7381]));
    assign layer1_outputs[10522] = (layer0_outputs[9292]) ^ (layer0_outputs[1348]);
    assign layer1_outputs[10523] = (layer0_outputs[8262]) & ~(layer0_outputs[1936]);
    assign layer1_outputs[10524] = ~((layer0_outputs[9126]) | (layer0_outputs[9845]));
    assign layer1_outputs[10525] = ~(layer0_outputs[9103]) | (layer0_outputs[6781]);
    assign layer1_outputs[10526] = (layer0_outputs[2286]) & ~(layer0_outputs[1731]);
    assign layer1_outputs[10527] = ~(layer0_outputs[7856]) | (layer0_outputs[3202]);
    assign layer1_outputs[10528] = layer0_outputs[11439];
    assign layer1_outputs[10529] = ~((layer0_outputs[12730]) & (layer0_outputs[10636]));
    assign layer1_outputs[10530] = layer0_outputs[1069];
    assign layer1_outputs[10531] = (layer0_outputs[3176]) ^ (layer0_outputs[9812]);
    assign layer1_outputs[10532] = ~((layer0_outputs[11952]) & (layer0_outputs[234]));
    assign layer1_outputs[10533] = (layer0_outputs[8896]) & ~(layer0_outputs[9715]);
    assign layer1_outputs[10534] = ~(layer0_outputs[8069]);
    assign layer1_outputs[10535] = ~(layer0_outputs[2013]);
    assign layer1_outputs[10536] = layer0_outputs[6828];
    assign layer1_outputs[10537] = ~((layer0_outputs[6008]) | (layer0_outputs[1758]));
    assign layer1_outputs[10538] = ~(layer0_outputs[9403]);
    assign layer1_outputs[10539] = (layer0_outputs[4111]) ^ (layer0_outputs[11652]);
    assign layer1_outputs[10540] = ~(layer0_outputs[9136]);
    assign layer1_outputs[10541] = 1'b1;
    assign layer1_outputs[10542] = ~((layer0_outputs[11798]) & (layer0_outputs[2196]));
    assign layer1_outputs[10543] = (layer0_outputs[9155]) | (layer0_outputs[1775]);
    assign layer1_outputs[10544] = ~((layer0_outputs[11300]) | (layer0_outputs[11456]));
    assign layer1_outputs[10545] = (layer0_outputs[3763]) ^ (layer0_outputs[9417]);
    assign layer1_outputs[10546] = layer0_outputs[5373];
    assign layer1_outputs[10547] = (layer0_outputs[11125]) ^ (layer0_outputs[270]);
    assign layer1_outputs[10548] = 1'b0;
    assign layer1_outputs[10549] = ~(layer0_outputs[7910]) | (layer0_outputs[702]);
    assign layer1_outputs[10550] = (layer0_outputs[8922]) | (layer0_outputs[10326]);
    assign layer1_outputs[10551] = (layer0_outputs[7162]) ^ (layer0_outputs[327]);
    assign layer1_outputs[10552] = (layer0_outputs[7236]) ^ (layer0_outputs[9123]);
    assign layer1_outputs[10553] = ~(layer0_outputs[11691]);
    assign layer1_outputs[10554] = ~((layer0_outputs[4508]) & (layer0_outputs[7452]));
    assign layer1_outputs[10555] = ~(layer0_outputs[5888]) | (layer0_outputs[11378]);
    assign layer1_outputs[10556] = ~(layer0_outputs[10794]) | (layer0_outputs[12701]);
    assign layer1_outputs[10557] = ~(layer0_outputs[1215]);
    assign layer1_outputs[10558] = 1'b0;
    assign layer1_outputs[10559] = ~((layer0_outputs[11443]) | (layer0_outputs[6068]));
    assign layer1_outputs[10560] = (layer0_outputs[12204]) & ~(layer0_outputs[2296]);
    assign layer1_outputs[10561] = (layer0_outputs[7260]) | (layer0_outputs[5780]);
    assign layer1_outputs[10562] = ~(layer0_outputs[7617]) | (layer0_outputs[5724]);
    assign layer1_outputs[10563] = ~(layer0_outputs[5123]);
    assign layer1_outputs[10564] = ~(layer0_outputs[6882]);
    assign layer1_outputs[10565] = layer0_outputs[2296];
    assign layer1_outputs[10566] = ~(layer0_outputs[11287]) | (layer0_outputs[11854]);
    assign layer1_outputs[10567] = layer0_outputs[5152];
    assign layer1_outputs[10568] = layer0_outputs[11345];
    assign layer1_outputs[10569] = layer0_outputs[7413];
    assign layer1_outputs[10570] = ~(layer0_outputs[958]);
    assign layer1_outputs[10571] = (layer0_outputs[10558]) & ~(layer0_outputs[3078]);
    assign layer1_outputs[10572] = (layer0_outputs[1025]) & ~(layer0_outputs[3235]);
    assign layer1_outputs[10573] = ~(layer0_outputs[10889]) | (layer0_outputs[7063]);
    assign layer1_outputs[10574] = ~(layer0_outputs[9727]) | (layer0_outputs[3971]);
    assign layer1_outputs[10575] = (layer0_outputs[4507]) & (layer0_outputs[37]);
    assign layer1_outputs[10576] = ~((layer0_outputs[11812]) & (layer0_outputs[8247]));
    assign layer1_outputs[10577] = (layer0_outputs[2643]) | (layer0_outputs[7143]);
    assign layer1_outputs[10578] = 1'b0;
    assign layer1_outputs[10579] = ~(layer0_outputs[12014]);
    assign layer1_outputs[10580] = layer0_outputs[3223];
    assign layer1_outputs[10581] = ~((layer0_outputs[3198]) & (layer0_outputs[3319]));
    assign layer1_outputs[10582] = ~(layer0_outputs[6584]);
    assign layer1_outputs[10583] = ~((layer0_outputs[7149]) | (layer0_outputs[8630]));
    assign layer1_outputs[10584] = ~((layer0_outputs[4290]) ^ (layer0_outputs[5362]));
    assign layer1_outputs[10585] = layer0_outputs[1227];
    assign layer1_outputs[10586] = layer0_outputs[3915];
    assign layer1_outputs[10587] = ~((layer0_outputs[3456]) ^ (layer0_outputs[3862]));
    assign layer1_outputs[10588] = layer0_outputs[1449];
    assign layer1_outputs[10589] = (layer0_outputs[5643]) & ~(layer0_outputs[7101]);
    assign layer1_outputs[10590] = ~((layer0_outputs[9881]) | (layer0_outputs[3537]));
    assign layer1_outputs[10591] = (layer0_outputs[7620]) ^ (layer0_outputs[3275]);
    assign layer1_outputs[10592] = ~((layer0_outputs[8465]) | (layer0_outputs[11769]));
    assign layer1_outputs[10593] = ~(layer0_outputs[7951]) | (layer0_outputs[8395]);
    assign layer1_outputs[10594] = ~(layer0_outputs[4572]);
    assign layer1_outputs[10595] = layer0_outputs[9209];
    assign layer1_outputs[10596] = ~((layer0_outputs[1642]) & (layer0_outputs[685]));
    assign layer1_outputs[10597] = ~((layer0_outputs[10610]) | (layer0_outputs[7043]));
    assign layer1_outputs[10598] = layer0_outputs[8305];
    assign layer1_outputs[10599] = ~(layer0_outputs[11755]);
    assign layer1_outputs[10600] = ~(layer0_outputs[7241]);
    assign layer1_outputs[10601] = (layer0_outputs[9377]) & ~(layer0_outputs[1406]);
    assign layer1_outputs[10602] = (layer0_outputs[1866]) & ~(layer0_outputs[9591]);
    assign layer1_outputs[10603] = ~(layer0_outputs[8281]);
    assign layer1_outputs[10604] = (layer0_outputs[10814]) & ~(layer0_outputs[11063]);
    assign layer1_outputs[10605] = (layer0_outputs[10766]) & (layer0_outputs[6298]);
    assign layer1_outputs[10606] = layer0_outputs[5120];
    assign layer1_outputs[10607] = ~((layer0_outputs[8338]) | (layer0_outputs[10863]));
    assign layer1_outputs[10608] = ~(layer0_outputs[4008]) | (layer0_outputs[3023]);
    assign layer1_outputs[10609] = layer0_outputs[6627];
    assign layer1_outputs[10610] = ~(layer0_outputs[500]);
    assign layer1_outputs[10611] = ~((layer0_outputs[4601]) ^ (layer0_outputs[2723]));
    assign layer1_outputs[10612] = layer0_outputs[5519];
    assign layer1_outputs[10613] = (layer0_outputs[5307]) ^ (layer0_outputs[4411]);
    assign layer1_outputs[10614] = layer0_outputs[10517];
    assign layer1_outputs[10615] = ~((layer0_outputs[5251]) | (layer0_outputs[1635]));
    assign layer1_outputs[10616] = (layer0_outputs[6897]) & ~(layer0_outputs[11331]);
    assign layer1_outputs[10617] = ~(layer0_outputs[6579]);
    assign layer1_outputs[10618] = (layer0_outputs[581]) | (layer0_outputs[1333]);
    assign layer1_outputs[10619] = (layer0_outputs[6147]) | (layer0_outputs[8419]);
    assign layer1_outputs[10620] = layer0_outputs[2263];
    assign layer1_outputs[10621] = layer0_outputs[4824];
    assign layer1_outputs[10622] = ~(layer0_outputs[9345]) | (layer0_outputs[6953]);
    assign layer1_outputs[10623] = (layer0_outputs[11289]) & ~(layer0_outputs[6241]);
    assign layer1_outputs[10624] = ~((layer0_outputs[1102]) | (layer0_outputs[4064]));
    assign layer1_outputs[10625] = layer0_outputs[5887];
    assign layer1_outputs[10626] = (layer0_outputs[2424]) ^ (layer0_outputs[4005]);
    assign layer1_outputs[10627] = ~((layer0_outputs[5363]) | (layer0_outputs[10074]));
    assign layer1_outputs[10628] = 1'b1;
    assign layer1_outputs[10629] = ~(layer0_outputs[8231]) | (layer0_outputs[1608]);
    assign layer1_outputs[10630] = (layer0_outputs[1786]) & ~(layer0_outputs[6718]);
    assign layer1_outputs[10631] = ~(layer0_outputs[220]);
    assign layer1_outputs[10632] = (layer0_outputs[2050]) ^ (layer0_outputs[1360]);
    assign layer1_outputs[10633] = ~((layer0_outputs[6001]) & (layer0_outputs[12275]));
    assign layer1_outputs[10634] = layer0_outputs[10443];
    assign layer1_outputs[10635] = ~(layer0_outputs[5585]);
    assign layer1_outputs[10636] = (layer0_outputs[7191]) ^ (layer0_outputs[5995]);
    assign layer1_outputs[10637] = layer0_outputs[12722];
    assign layer1_outputs[10638] = ~(layer0_outputs[4606]);
    assign layer1_outputs[10639] = ~(layer0_outputs[10367]);
    assign layer1_outputs[10640] = ~((layer0_outputs[9813]) ^ (layer0_outputs[8127]));
    assign layer1_outputs[10641] = ~(layer0_outputs[6960]) | (layer0_outputs[4624]);
    assign layer1_outputs[10642] = ~(layer0_outputs[1176]);
    assign layer1_outputs[10643] = ~((layer0_outputs[11656]) & (layer0_outputs[5623]));
    assign layer1_outputs[10644] = (layer0_outputs[12050]) & (layer0_outputs[9848]);
    assign layer1_outputs[10645] = ~(layer0_outputs[3984]);
    assign layer1_outputs[10646] = (layer0_outputs[10883]) | (layer0_outputs[4390]);
    assign layer1_outputs[10647] = ~(layer0_outputs[4216]) | (layer0_outputs[3832]);
    assign layer1_outputs[10648] = ~((layer0_outputs[5377]) | (layer0_outputs[1620]));
    assign layer1_outputs[10649] = ~(layer0_outputs[8913]);
    assign layer1_outputs[10650] = ~((layer0_outputs[11938]) | (layer0_outputs[10957]));
    assign layer1_outputs[10651] = layer0_outputs[11461];
    assign layer1_outputs[10652] = ~(layer0_outputs[4413]) | (layer0_outputs[2571]);
    assign layer1_outputs[10653] = ~(layer0_outputs[2165]);
    assign layer1_outputs[10654] = (layer0_outputs[6080]) ^ (layer0_outputs[6587]);
    assign layer1_outputs[10655] = 1'b0;
    assign layer1_outputs[10656] = ~(layer0_outputs[11582]);
    assign layer1_outputs[10657] = (layer0_outputs[4096]) & ~(layer0_outputs[8608]);
    assign layer1_outputs[10658] = (layer0_outputs[11754]) & ~(layer0_outputs[4423]);
    assign layer1_outputs[10659] = ~(layer0_outputs[11003]);
    assign layer1_outputs[10660] = (layer0_outputs[9970]) | (layer0_outputs[9380]);
    assign layer1_outputs[10661] = ~(layer0_outputs[3450]) | (layer0_outputs[7895]);
    assign layer1_outputs[10662] = ~((layer0_outputs[4590]) | (layer0_outputs[4046]));
    assign layer1_outputs[10663] = ~((layer0_outputs[11070]) & (layer0_outputs[12715]));
    assign layer1_outputs[10664] = ~(layer0_outputs[610]);
    assign layer1_outputs[10665] = (layer0_outputs[994]) & ~(layer0_outputs[679]);
    assign layer1_outputs[10666] = layer0_outputs[6516];
    assign layer1_outputs[10667] = (layer0_outputs[11813]) | (layer0_outputs[9421]);
    assign layer1_outputs[10668] = ~(layer0_outputs[7181]) | (layer0_outputs[6364]);
    assign layer1_outputs[10669] = ~(layer0_outputs[6545]);
    assign layer1_outputs[10670] = (layer0_outputs[3256]) & ~(layer0_outputs[4627]);
    assign layer1_outputs[10671] = (layer0_outputs[3198]) & ~(layer0_outputs[10226]);
    assign layer1_outputs[10672] = (layer0_outputs[9121]) | (layer0_outputs[3552]);
    assign layer1_outputs[10673] = (layer0_outputs[5295]) & ~(layer0_outputs[3894]);
    assign layer1_outputs[10674] = (layer0_outputs[8392]) ^ (layer0_outputs[1309]);
    assign layer1_outputs[10675] = ~(layer0_outputs[12612]) | (layer0_outputs[7743]);
    assign layer1_outputs[10676] = (layer0_outputs[3148]) & ~(layer0_outputs[10482]);
    assign layer1_outputs[10677] = ~((layer0_outputs[8196]) | (layer0_outputs[853]));
    assign layer1_outputs[10678] = (layer0_outputs[11429]) ^ (layer0_outputs[2998]);
    assign layer1_outputs[10679] = ~((layer0_outputs[2247]) & (layer0_outputs[6381]));
    assign layer1_outputs[10680] = (layer0_outputs[1151]) & ~(layer0_outputs[7796]);
    assign layer1_outputs[10681] = layer0_outputs[39];
    assign layer1_outputs[10682] = ~(layer0_outputs[10821]);
    assign layer1_outputs[10683] = layer0_outputs[4003];
    assign layer1_outputs[10684] = layer0_outputs[2141];
    assign layer1_outputs[10685] = ~(layer0_outputs[1335]) | (layer0_outputs[12649]);
    assign layer1_outputs[10686] = ~((layer0_outputs[4059]) | (layer0_outputs[9203]));
    assign layer1_outputs[10687] = ~(layer0_outputs[9350]);
    assign layer1_outputs[10688] = (layer0_outputs[4567]) ^ (layer0_outputs[11639]);
    assign layer1_outputs[10689] = ~((layer0_outputs[7317]) | (layer0_outputs[3829]));
    assign layer1_outputs[10690] = ~((layer0_outputs[3162]) ^ (layer0_outputs[7585]));
    assign layer1_outputs[10691] = layer0_outputs[10808];
    assign layer1_outputs[10692] = 1'b1;
    assign layer1_outputs[10693] = ~(layer0_outputs[9379]) | (layer0_outputs[11676]);
    assign layer1_outputs[10694] = ~(layer0_outputs[6638]);
    assign layer1_outputs[10695] = ~((layer0_outputs[11739]) & (layer0_outputs[9171]));
    assign layer1_outputs[10696] = ~(layer0_outputs[60]);
    assign layer1_outputs[10697] = ~(layer0_outputs[5358]);
    assign layer1_outputs[10698] = ~(layer0_outputs[2470]);
    assign layer1_outputs[10699] = ~((layer0_outputs[7673]) ^ (layer0_outputs[8141]));
    assign layer1_outputs[10700] = ~((layer0_outputs[7593]) | (layer0_outputs[5602]));
    assign layer1_outputs[10701] = (layer0_outputs[2526]) ^ (layer0_outputs[12179]);
    assign layer1_outputs[10702] = (layer0_outputs[3561]) ^ (layer0_outputs[8057]);
    assign layer1_outputs[10703] = (layer0_outputs[10801]) & (layer0_outputs[6960]);
    assign layer1_outputs[10704] = layer0_outputs[610];
    assign layer1_outputs[10705] = ~(layer0_outputs[11054]) | (layer0_outputs[11830]);
    assign layer1_outputs[10706] = ~((layer0_outputs[1501]) & (layer0_outputs[2207]));
    assign layer1_outputs[10707] = ~(layer0_outputs[10572]) | (layer0_outputs[4632]);
    assign layer1_outputs[10708] = layer0_outputs[11551];
    assign layer1_outputs[10709] = layer0_outputs[7340];
    assign layer1_outputs[10710] = (layer0_outputs[6169]) ^ (layer0_outputs[49]);
    assign layer1_outputs[10711] = (layer0_outputs[9644]) & ~(layer0_outputs[5271]);
    assign layer1_outputs[10712] = ~(layer0_outputs[1148]);
    assign layer1_outputs[10713] = layer0_outputs[9686];
    assign layer1_outputs[10714] = ~(layer0_outputs[10814]);
    assign layer1_outputs[10715] = ~(layer0_outputs[8607]);
    assign layer1_outputs[10716] = ~(layer0_outputs[12508]);
    assign layer1_outputs[10717] = ~(layer0_outputs[6078]);
    assign layer1_outputs[10718] = (layer0_outputs[11091]) ^ (layer0_outputs[12033]);
    assign layer1_outputs[10719] = ~(layer0_outputs[11278]);
    assign layer1_outputs[10720] = ~((layer0_outputs[2497]) & (layer0_outputs[7889]));
    assign layer1_outputs[10721] = 1'b0;
    assign layer1_outputs[10722] = (layer0_outputs[5568]) & ~(layer0_outputs[5868]);
    assign layer1_outputs[10723] = layer0_outputs[580];
    assign layer1_outputs[10724] = 1'b1;
    assign layer1_outputs[10725] = ~((layer0_outputs[1978]) | (layer0_outputs[11220]));
    assign layer1_outputs[10726] = ~((layer0_outputs[7236]) & (layer0_outputs[3589]));
    assign layer1_outputs[10727] = ~(layer0_outputs[11591]);
    assign layer1_outputs[10728] = ~((layer0_outputs[3560]) | (layer0_outputs[7257]));
    assign layer1_outputs[10729] = ~(layer0_outputs[12318]);
    assign layer1_outputs[10730] = ~(layer0_outputs[9249]);
    assign layer1_outputs[10731] = layer0_outputs[7574];
    assign layer1_outputs[10732] = ~(layer0_outputs[4519]);
    assign layer1_outputs[10733] = (layer0_outputs[10905]) & (layer0_outputs[6295]);
    assign layer1_outputs[10734] = layer0_outputs[1911];
    assign layer1_outputs[10735] = layer0_outputs[9410];
    assign layer1_outputs[10736] = ~((layer0_outputs[12083]) & (layer0_outputs[8231]));
    assign layer1_outputs[10737] = ~((layer0_outputs[2718]) & (layer0_outputs[1060]));
    assign layer1_outputs[10738] = (layer0_outputs[3280]) | (layer0_outputs[199]);
    assign layer1_outputs[10739] = ~(layer0_outputs[12761]);
    assign layer1_outputs[10740] = layer0_outputs[3651];
    assign layer1_outputs[10741] = ~(layer0_outputs[3032]);
    assign layer1_outputs[10742] = layer0_outputs[1017];
    assign layer1_outputs[10743] = (layer0_outputs[7388]) | (layer0_outputs[6840]);
    assign layer1_outputs[10744] = ~((layer0_outputs[6904]) ^ (layer0_outputs[5525]));
    assign layer1_outputs[10745] = ~((layer0_outputs[3422]) & (layer0_outputs[2928]));
    assign layer1_outputs[10746] = layer0_outputs[3419];
    assign layer1_outputs[10747] = layer0_outputs[11079];
    assign layer1_outputs[10748] = (layer0_outputs[5399]) ^ (layer0_outputs[1414]);
    assign layer1_outputs[10749] = (layer0_outputs[5407]) & (layer0_outputs[4986]);
    assign layer1_outputs[10750] = layer0_outputs[2105];
    assign layer1_outputs[10751] = layer0_outputs[3707];
    assign layer1_outputs[10752] = (layer0_outputs[3116]) & ~(layer0_outputs[2597]);
    assign layer1_outputs[10753] = ~(layer0_outputs[5145]);
    assign layer1_outputs[10754] = layer0_outputs[6378];
    assign layer1_outputs[10755] = (layer0_outputs[6544]) & ~(layer0_outputs[1202]);
    assign layer1_outputs[10756] = layer0_outputs[3831];
    assign layer1_outputs[10757] = ~(layer0_outputs[3059]) | (layer0_outputs[9255]);
    assign layer1_outputs[10758] = ~((layer0_outputs[777]) & (layer0_outputs[5491]));
    assign layer1_outputs[10759] = ~(layer0_outputs[6549]) | (layer0_outputs[8954]);
    assign layer1_outputs[10760] = (layer0_outputs[5698]) | (layer0_outputs[8299]);
    assign layer1_outputs[10761] = ~(layer0_outputs[11517]);
    assign layer1_outputs[10762] = ~((layer0_outputs[8810]) ^ (layer0_outputs[7546]));
    assign layer1_outputs[10763] = ~((layer0_outputs[1303]) | (layer0_outputs[8737]));
    assign layer1_outputs[10764] = layer0_outputs[3117];
    assign layer1_outputs[10765] = ~(layer0_outputs[3518]);
    assign layer1_outputs[10766] = ~((layer0_outputs[9215]) | (layer0_outputs[1875]));
    assign layer1_outputs[10767] = ~((layer0_outputs[9134]) ^ (layer0_outputs[8692]));
    assign layer1_outputs[10768] = 1'b0;
    assign layer1_outputs[10769] = ~(layer0_outputs[7061]);
    assign layer1_outputs[10770] = (layer0_outputs[2803]) & (layer0_outputs[1960]);
    assign layer1_outputs[10771] = (layer0_outputs[1671]) & ~(layer0_outputs[4279]);
    assign layer1_outputs[10772] = layer0_outputs[8548];
    assign layer1_outputs[10773] = layer0_outputs[12603];
    assign layer1_outputs[10774] = layer0_outputs[9514];
    assign layer1_outputs[10775] = (layer0_outputs[8044]) & ~(layer0_outputs[9376]);
    assign layer1_outputs[10776] = (layer0_outputs[11079]) | (layer0_outputs[8260]);
    assign layer1_outputs[10777] = ~(layer0_outputs[9894]) | (layer0_outputs[10533]);
    assign layer1_outputs[10778] = ~((layer0_outputs[8217]) & (layer0_outputs[10538]));
    assign layer1_outputs[10779] = layer0_outputs[3423];
    assign layer1_outputs[10780] = ~((layer0_outputs[1961]) | (layer0_outputs[6949]));
    assign layer1_outputs[10781] = (layer0_outputs[653]) & ~(layer0_outputs[6262]);
    assign layer1_outputs[10782] = ~(layer0_outputs[8204]);
    assign layer1_outputs[10783] = (layer0_outputs[10655]) & ~(layer0_outputs[8415]);
    assign layer1_outputs[10784] = ~(layer0_outputs[5778]) | (layer0_outputs[9043]);
    assign layer1_outputs[10785] = ~(layer0_outputs[428]);
    assign layer1_outputs[10786] = layer0_outputs[11860];
    assign layer1_outputs[10787] = (layer0_outputs[3505]) | (layer0_outputs[7257]);
    assign layer1_outputs[10788] = ~(layer0_outputs[1722]);
    assign layer1_outputs[10789] = ~(layer0_outputs[10255]) | (layer0_outputs[9422]);
    assign layer1_outputs[10790] = (layer0_outputs[3515]) & ~(layer0_outputs[3627]);
    assign layer1_outputs[10791] = (layer0_outputs[4484]) & ~(layer0_outputs[5600]);
    assign layer1_outputs[10792] = ~(layer0_outputs[4694]) | (layer0_outputs[2263]);
    assign layer1_outputs[10793] = (layer0_outputs[12250]) & ~(layer0_outputs[1220]);
    assign layer1_outputs[10794] = (layer0_outputs[7686]) & (layer0_outputs[1466]);
    assign layer1_outputs[10795] = (layer0_outputs[9401]) | (layer0_outputs[12338]);
    assign layer1_outputs[10796] = ~((layer0_outputs[4435]) ^ (layer0_outputs[10917]));
    assign layer1_outputs[10797] = (layer0_outputs[9310]) & (layer0_outputs[5641]);
    assign layer1_outputs[10798] = ~((layer0_outputs[7146]) ^ (layer0_outputs[4178]));
    assign layer1_outputs[10799] = layer0_outputs[3200];
    assign layer1_outputs[10800] = ~(layer0_outputs[10896]);
    assign layer1_outputs[10801] = (layer0_outputs[793]) | (layer0_outputs[3314]);
    assign layer1_outputs[10802] = layer0_outputs[1549];
    assign layer1_outputs[10803] = ~((layer0_outputs[6872]) | (layer0_outputs[9900]));
    assign layer1_outputs[10804] = layer0_outputs[11271];
    assign layer1_outputs[10805] = layer0_outputs[8791];
    assign layer1_outputs[10806] = layer0_outputs[4327];
    assign layer1_outputs[10807] = layer0_outputs[10898];
    assign layer1_outputs[10808] = ~(layer0_outputs[9414]) | (layer0_outputs[2251]);
    assign layer1_outputs[10809] = layer0_outputs[8639];
    assign layer1_outputs[10810] = (layer0_outputs[10829]) ^ (layer0_outputs[7325]);
    assign layer1_outputs[10811] = (layer0_outputs[5826]) & ~(layer0_outputs[7540]);
    assign layer1_outputs[10812] = ~(layer0_outputs[11874]);
    assign layer1_outputs[10813] = (layer0_outputs[10989]) ^ (layer0_outputs[7828]);
    assign layer1_outputs[10814] = ~(layer0_outputs[5371]);
    assign layer1_outputs[10815] = layer0_outputs[10370];
    assign layer1_outputs[10816] = ~((layer0_outputs[7050]) ^ (layer0_outputs[30]));
    assign layer1_outputs[10817] = ~(layer0_outputs[11392]);
    assign layer1_outputs[10818] = ~(layer0_outputs[7385]);
    assign layer1_outputs[10819] = ~(layer0_outputs[2330]) | (layer0_outputs[4219]);
    assign layer1_outputs[10820] = (layer0_outputs[10571]) & ~(layer0_outputs[6647]);
    assign layer1_outputs[10821] = ~((layer0_outputs[2709]) | (layer0_outputs[10474]));
    assign layer1_outputs[10822] = (layer0_outputs[1536]) ^ (layer0_outputs[10551]);
    assign layer1_outputs[10823] = (layer0_outputs[6336]) & ~(layer0_outputs[12599]);
    assign layer1_outputs[10824] = (layer0_outputs[637]) & ~(layer0_outputs[1792]);
    assign layer1_outputs[10825] = ~(layer0_outputs[589]);
    assign layer1_outputs[10826] = ~(layer0_outputs[4791]);
    assign layer1_outputs[10827] = ~(layer0_outputs[8178]);
    assign layer1_outputs[10828] = layer0_outputs[5648];
    assign layer1_outputs[10829] = (layer0_outputs[385]) & ~(layer0_outputs[992]);
    assign layer1_outputs[10830] = layer0_outputs[11229];
    assign layer1_outputs[10831] = ~(layer0_outputs[3546]) | (layer0_outputs[7283]);
    assign layer1_outputs[10832] = ~(layer0_outputs[6690]);
    assign layer1_outputs[10833] = (layer0_outputs[7721]) & ~(layer0_outputs[2137]);
    assign layer1_outputs[10834] = (layer0_outputs[11472]) & ~(layer0_outputs[8135]);
    assign layer1_outputs[10835] = (layer0_outputs[7170]) | (layer0_outputs[2245]);
    assign layer1_outputs[10836] = ~(layer0_outputs[11438]) | (layer0_outputs[6415]);
    assign layer1_outputs[10837] = ~(layer0_outputs[9208]);
    assign layer1_outputs[10838] = layer0_outputs[11883];
    assign layer1_outputs[10839] = ~(layer0_outputs[12564]) | (layer0_outputs[10857]);
    assign layer1_outputs[10840] = ~(layer0_outputs[4913]) | (layer0_outputs[1932]);
    assign layer1_outputs[10841] = (layer0_outputs[5391]) & ~(layer0_outputs[2661]);
    assign layer1_outputs[10842] = ~((layer0_outputs[9145]) & (layer0_outputs[7628]));
    assign layer1_outputs[10843] = (layer0_outputs[12640]) & (layer0_outputs[2382]);
    assign layer1_outputs[10844] = 1'b0;
    assign layer1_outputs[10845] = ~(layer0_outputs[7464]);
    assign layer1_outputs[10846] = ~((layer0_outputs[12160]) & (layer0_outputs[7992]));
    assign layer1_outputs[10847] = layer0_outputs[798];
    assign layer1_outputs[10848] = (layer0_outputs[11155]) & ~(layer0_outputs[406]);
    assign layer1_outputs[10849] = ~(layer0_outputs[8700]) | (layer0_outputs[1741]);
    assign layer1_outputs[10850] = ~(layer0_outputs[7097]);
    assign layer1_outputs[10851] = 1'b0;
    assign layer1_outputs[10852] = ~(layer0_outputs[3819]) | (layer0_outputs[3090]);
    assign layer1_outputs[10853] = ~(layer0_outputs[217]);
    assign layer1_outputs[10854] = ~(layer0_outputs[5632]);
    assign layer1_outputs[10855] = (layer0_outputs[6484]) & ~(layer0_outputs[2166]);
    assign layer1_outputs[10856] = ~((layer0_outputs[9378]) | (layer0_outputs[5036]));
    assign layer1_outputs[10857] = ~(layer0_outputs[5299]) | (layer0_outputs[363]);
    assign layer1_outputs[10858] = (layer0_outputs[8522]) & (layer0_outputs[971]);
    assign layer1_outputs[10859] = ~((layer0_outputs[11223]) & (layer0_outputs[12126]));
    assign layer1_outputs[10860] = (layer0_outputs[11298]) & (layer0_outputs[6562]);
    assign layer1_outputs[10861] = ~(layer0_outputs[5443]);
    assign layer1_outputs[10862] = ~((layer0_outputs[849]) & (layer0_outputs[5071]));
    assign layer1_outputs[10863] = (layer0_outputs[5162]) & (layer0_outputs[2082]);
    assign layer1_outputs[10864] = (layer0_outputs[2127]) & ~(layer0_outputs[7048]);
    assign layer1_outputs[10865] = ~(layer0_outputs[2783]) | (layer0_outputs[10518]);
    assign layer1_outputs[10866] = ~(layer0_outputs[5787]) | (layer0_outputs[9892]);
    assign layer1_outputs[10867] = (layer0_outputs[12383]) & (layer0_outputs[3519]);
    assign layer1_outputs[10868] = (layer0_outputs[8363]) | (layer0_outputs[9413]);
    assign layer1_outputs[10869] = ~(layer0_outputs[8899]) | (layer0_outputs[7992]);
    assign layer1_outputs[10870] = ~((layer0_outputs[6818]) & (layer0_outputs[2559]));
    assign layer1_outputs[10871] = (layer0_outputs[137]) | (layer0_outputs[7846]);
    assign layer1_outputs[10872] = 1'b1;
    assign layer1_outputs[10873] = ~(layer0_outputs[1967]);
    assign layer1_outputs[10874] = ~(layer0_outputs[5134]) | (layer0_outputs[8496]);
    assign layer1_outputs[10875] = ~(layer0_outputs[5418]);
    assign layer1_outputs[10876] = (layer0_outputs[8167]) & ~(layer0_outputs[4676]);
    assign layer1_outputs[10877] = ~(layer0_outputs[10279]) | (layer0_outputs[637]);
    assign layer1_outputs[10878] = ~(layer0_outputs[5956]);
    assign layer1_outputs[10879] = (layer0_outputs[3373]) & (layer0_outputs[7189]);
    assign layer1_outputs[10880] = (layer0_outputs[6665]) & ~(layer0_outputs[9934]);
    assign layer1_outputs[10881] = ~(layer0_outputs[10235]) | (layer0_outputs[3131]);
    assign layer1_outputs[10882] = (layer0_outputs[1750]) & ~(layer0_outputs[8209]);
    assign layer1_outputs[10883] = layer0_outputs[9551];
    assign layer1_outputs[10884] = ~((layer0_outputs[3727]) & (layer0_outputs[30]));
    assign layer1_outputs[10885] = layer0_outputs[1041];
    assign layer1_outputs[10886] = ~(layer0_outputs[4123]) | (layer0_outputs[1336]);
    assign layer1_outputs[10887] = (layer0_outputs[10530]) & ~(layer0_outputs[11750]);
    assign layer1_outputs[10888] = ~(layer0_outputs[11655]);
    assign layer1_outputs[10889] = ~((layer0_outputs[5706]) ^ (layer0_outputs[10146]));
    assign layer1_outputs[10890] = layer0_outputs[6159];
    assign layer1_outputs[10891] = ~(layer0_outputs[2774]) | (layer0_outputs[1485]);
    assign layer1_outputs[10892] = ~(layer0_outputs[10742]);
    assign layer1_outputs[10893] = ~(layer0_outputs[12436]) | (layer0_outputs[7607]);
    assign layer1_outputs[10894] = (layer0_outputs[10256]) | (layer0_outputs[1122]);
    assign layer1_outputs[10895] = layer0_outputs[3626];
    assign layer1_outputs[10896] = (layer0_outputs[2372]) & ~(layer0_outputs[6985]);
    assign layer1_outputs[10897] = (layer0_outputs[10777]) & (layer0_outputs[11672]);
    assign layer1_outputs[10898] = ~(layer0_outputs[7282]);
    assign layer1_outputs[10899] = ~((layer0_outputs[12073]) | (layer0_outputs[11055]));
    assign layer1_outputs[10900] = layer0_outputs[4378];
    assign layer1_outputs[10901] = layer0_outputs[9027];
    assign layer1_outputs[10902] = ~(layer0_outputs[8666]) | (layer0_outputs[7721]);
    assign layer1_outputs[10903] = ~((layer0_outputs[7195]) | (layer0_outputs[12771]));
    assign layer1_outputs[10904] = layer0_outputs[8352];
    assign layer1_outputs[10905] = ~(layer0_outputs[2331]) | (layer0_outputs[5682]);
    assign layer1_outputs[10906] = ~((layer0_outputs[2528]) ^ (layer0_outputs[5312]));
    assign layer1_outputs[10907] = ~(layer0_outputs[11989]);
    assign layer1_outputs[10908] = 1'b1;
    assign layer1_outputs[10909] = layer0_outputs[2826];
    assign layer1_outputs[10910] = ~((layer0_outputs[11365]) & (layer0_outputs[265]));
    assign layer1_outputs[10911] = ~(layer0_outputs[8662]);
    assign layer1_outputs[10912] = (layer0_outputs[6379]) | (layer0_outputs[9244]);
    assign layer1_outputs[10913] = layer0_outputs[1966];
    assign layer1_outputs[10914] = layer0_outputs[9124];
    assign layer1_outputs[10915] = ~((layer0_outputs[2139]) & (layer0_outputs[12577]));
    assign layer1_outputs[10916] = (layer0_outputs[11262]) & ~(layer0_outputs[3364]);
    assign layer1_outputs[10917] = (layer0_outputs[3190]) & (layer0_outputs[11511]);
    assign layer1_outputs[10918] = layer0_outputs[677];
    assign layer1_outputs[10919] = (layer0_outputs[2383]) & ~(layer0_outputs[5705]);
    assign layer1_outputs[10920] = layer0_outputs[5864];
    assign layer1_outputs[10921] = 1'b1;
    assign layer1_outputs[10922] = layer0_outputs[11502];
    assign layer1_outputs[10923] = (layer0_outputs[7712]) ^ (layer0_outputs[10840]);
    assign layer1_outputs[10924] = ~((layer0_outputs[5034]) & (layer0_outputs[4555]));
    assign layer1_outputs[10925] = ~(layer0_outputs[3136]);
    assign layer1_outputs[10926] = (layer0_outputs[10516]) & ~(layer0_outputs[9437]);
    assign layer1_outputs[10927] = (layer0_outputs[11697]) ^ (layer0_outputs[2461]);
    assign layer1_outputs[10928] = (layer0_outputs[4487]) ^ (layer0_outputs[10198]);
    assign layer1_outputs[10929] = layer0_outputs[5073];
    assign layer1_outputs[10930] = (layer0_outputs[12016]) & ~(layer0_outputs[3274]);
    assign layer1_outputs[10931] = (layer0_outputs[5590]) & ~(layer0_outputs[5359]);
    assign layer1_outputs[10932] = layer0_outputs[8183];
    assign layer1_outputs[10933] = layer0_outputs[5865];
    assign layer1_outputs[10934] = ~(layer0_outputs[8555]);
    assign layer1_outputs[10935] = (layer0_outputs[4423]) ^ (layer0_outputs[7203]);
    assign layer1_outputs[10936] = 1'b0;
    assign layer1_outputs[10937] = ~((layer0_outputs[6071]) ^ (layer0_outputs[3368]));
    assign layer1_outputs[10938] = (layer0_outputs[7956]) & ~(layer0_outputs[966]);
    assign layer1_outputs[10939] = (layer0_outputs[116]) | (layer0_outputs[5106]);
    assign layer1_outputs[10940] = layer0_outputs[2872];
    assign layer1_outputs[10941] = layer0_outputs[5172];
    assign layer1_outputs[10942] = (layer0_outputs[6631]) & ~(layer0_outputs[7528]);
    assign layer1_outputs[10943] = ~(layer0_outputs[11828]) | (layer0_outputs[2869]);
    assign layer1_outputs[10944] = (layer0_outputs[10974]) | (layer0_outputs[12213]);
    assign layer1_outputs[10945] = (layer0_outputs[12643]) | (layer0_outputs[1425]);
    assign layer1_outputs[10946] = ~(layer0_outputs[12743]);
    assign layer1_outputs[10947] = (layer0_outputs[11448]) ^ (layer0_outputs[6554]);
    assign layer1_outputs[10948] = layer0_outputs[1480];
    assign layer1_outputs[10949] = ~((layer0_outputs[4565]) & (layer0_outputs[9777]));
    assign layer1_outputs[10950] = layer0_outputs[11106];
    assign layer1_outputs[10951] = (layer0_outputs[10750]) | (layer0_outputs[11774]);
    assign layer1_outputs[10952] = (layer0_outputs[8099]) & (layer0_outputs[10308]);
    assign layer1_outputs[10953] = ~((layer0_outputs[6486]) & (layer0_outputs[10876]));
    assign layer1_outputs[10954] = ~((layer0_outputs[3313]) & (layer0_outputs[5967]));
    assign layer1_outputs[10955] = (layer0_outputs[10468]) & ~(layer0_outputs[12024]);
    assign layer1_outputs[10956] = ~(layer0_outputs[4620]) | (layer0_outputs[9633]);
    assign layer1_outputs[10957] = layer0_outputs[11962];
    assign layer1_outputs[10958] = ~(layer0_outputs[12403]) | (layer0_outputs[389]);
    assign layer1_outputs[10959] = (layer0_outputs[3400]) & ~(layer0_outputs[8117]);
    assign layer1_outputs[10960] = (layer0_outputs[10142]) & ~(layer0_outputs[10615]);
    assign layer1_outputs[10961] = layer0_outputs[8484];
    assign layer1_outputs[10962] = ~(layer0_outputs[4056]);
    assign layer1_outputs[10963] = 1'b1;
    assign layer1_outputs[10964] = layer0_outputs[7210];
    assign layer1_outputs[10965] = (layer0_outputs[219]) & (layer0_outputs[5583]);
    assign layer1_outputs[10966] = ~(layer0_outputs[8989]);
    assign layer1_outputs[10967] = ~(layer0_outputs[12225]);
    assign layer1_outputs[10968] = ~(layer0_outputs[7204]);
    assign layer1_outputs[10969] = ~((layer0_outputs[9376]) & (layer0_outputs[3503]));
    assign layer1_outputs[10970] = (layer0_outputs[5793]) | (layer0_outputs[8000]);
    assign layer1_outputs[10971] = ~(layer0_outputs[3369]);
    assign layer1_outputs[10972] = (layer0_outputs[2504]) ^ (layer0_outputs[9857]);
    assign layer1_outputs[10973] = ~(layer0_outputs[7560]);
    assign layer1_outputs[10974] = layer0_outputs[7715];
    assign layer1_outputs[10975] = layer0_outputs[688];
    assign layer1_outputs[10976] = layer0_outputs[10528];
    assign layer1_outputs[10977] = ~((layer0_outputs[8945]) & (layer0_outputs[6950]));
    assign layer1_outputs[10978] = (layer0_outputs[9863]) & (layer0_outputs[1788]);
    assign layer1_outputs[10979] = layer0_outputs[10532];
    assign layer1_outputs[10980] = (layer0_outputs[9473]) | (layer0_outputs[9037]);
    assign layer1_outputs[10981] = layer0_outputs[3902];
    assign layer1_outputs[10982] = (layer0_outputs[6811]) & ~(layer0_outputs[2743]);
    assign layer1_outputs[10983] = ~((layer0_outputs[6979]) ^ (layer0_outputs[8050]));
    assign layer1_outputs[10984] = ~(layer0_outputs[3157]);
    assign layer1_outputs[10985] = layer0_outputs[1357];
    assign layer1_outputs[10986] = ~(layer0_outputs[5972]);
    assign layer1_outputs[10987] = (layer0_outputs[1847]) & ~(layer0_outputs[5381]);
    assign layer1_outputs[10988] = ~(layer0_outputs[11014]);
    assign layer1_outputs[10989] = ~(layer0_outputs[1525]);
    assign layer1_outputs[10990] = (layer0_outputs[2860]) & (layer0_outputs[8549]);
    assign layer1_outputs[10991] = (layer0_outputs[4124]) & (layer0_outputs[8592]);
    assign layer1_outputs[10992] = layer0_outputs[1305];
    assign layer1_outputs[10993] = (layer0_outputs[1444]) & ~(layer0_outputs[11973]);
    assign layer1_outputs[10994] = ~(layer0_outputs[10219]);
    assign layer1_outputs[10995] = ~(layer0_outputs[9632]);
    assign layer1_outputs[10996] = ~(layer0_outputs[4197]) | (layer0_outputs[9402]);
    assign layer1_outputs[10997] = (layer0_outputs[9171]) & ~(layer0_outputs[4645]);
    assign layer1_outputs[10998] = ~((layer0_outputs[1316]) | (layer0_outputs[1639]));
    assign layer1_outputs[10999] = (layer0_outputs[2536]) & ~(layer0_outputs[990]);
    assign layer1_outputs[11000] = ~((layer0_outputs[5336]) ^ (layer0_outputs[4127]));
    assign layer1_outputs[11001] = ~((layer0_outputs[3293]) ^ (layer0_outputs[10094]));
    assign layer1_outputs[11002] = ~((layer0_outputs[5147]) ^ (layer0_outputs[794]));
    assign layer1_outputs[11003] = ~(layer0_outputs[5925]);
    assign layer1_outputs[11004] = layer0_outputs[8695];
    assign layer1_outputs[11005] = ~(layer0_outputs[7065]) | (layer0_outputs[12602]);
    assign layer1_outputs[11006] = ~((layer0_outputs[4844]) | (layer0_outputs[125]));
    assign layer1_outputs[11007] = 1'b1;
    assign layer1_outputs[11008] = ~((layer0_outputs[4190]) & (layer0_outputs[559]));
    assign layer1_outputs[11009] = ~(layer0_outputs[12562]) | (layer0_outputs[6541]);
    assign layer1_outputs[11010] = layer0_outputs[9736];
    assign layer1_outputs[11011] = ~((layer0_outputs[12786]) ^ (layer0_outputs[7194]));
    assign layer1_outputs[11012] = ~(layer0_outputs[6806]);
    assign layer1_outputs[11013] = ~((layer0_outputs[9518]) ^ (layer0_outputs[5535]));
    assign layer1_outputs[11014] = ~(layer0_outputs[4772]);
    assign layer1_outputs[11015] = ~((layer0_outputs[11819]) | (layer0_outputs[1129]));
    assign layer1_outputs[11016] = ~((layer0_outputs[12313]) & (layer0_outputs[5416]));
    assign layer1_outputs[11017] = ~(layer0_outputs[12343]);
    assign layer1_outputs[11018] = layer0_outputs[3714];
    assign layer1_outputs[11019] = (layer0_outputs[3155]) & ~(layer0_outputs[6244]);
    assign layer1_outputs[11020] = (layer0_outputs[6216]) & ~(layer0_outputs[1173]);
    assign layer1_outputs[11021] = (layer0_outputs[1024]) ^ (layer0_outputs[2762]);
    assign layer1_outputs[11022] = (layer0_outputs[6175]) | (layer0_outputs[3690]);
    assign layer1_outputs[11023] = (layer0_outputs[9086]) ^ (layer0_outputs[11705]);
    assign layer1_outputs[11024] = layer0_outputs[11260];
    assign layer1_outputs[11025] = 1'b1;
    assign layer1_outputs[11026] = ~(layer0_outputs[10781]);
    assign layer1_outputs[11027] = (layer0_outputs[11949]) & ~(layer0_outputs[5670]);
    assign layer1_outputs[11028] = (layer0_outputs[3510]) | (layer0_outputs[6532]);
    assign layer1_outputs[11029] = ~(layer0_outputs[3463]);
    assign layer1_outputs[11030] = layer0_outputs[10772];
    assign layer1_outputs[11031] = ~((layer0_outputs[223]) & (layer0_outputs[2350]));
    assign layer1_outputs[11032] = ~((layer0_outputs[955]) ^ (layer0_outputs[10386]));
    assign layer1_outputs[11033] = ~(layer0_outputs[3523]);
    assign layer1_outputs[11034] = (layer0_outputs[1403]) & (layer0_outputs[6839]);
    assign layer1_outputs[11035] = (layer0_outputs[7980]) & ~(layer0_outputs[5240]);
    assign layer1_outputs[11036] = ~((layer0_outputs[1374]) & (layer0_outputs[7398]));
    assign layer1_outputs[11037] = ~(layer0_outputs[339]);
    assign layer1_outputs[11038] = ~(layer0_outputs[3818]);
    assign layer1_outputs[11039] = 1'b1;
    assign layer1_outputs[11040] = ~(layer0_outputs[6469]);
    assign layer1_outputs[11041] = ~(layer0_outputs[6338]);
    assign layer1_outputs[11042] = (layer0_outputs[11684]) | (layer0_outputs[12310]);
    assign layer1_outputs[11043] = (layer0_outputs[5298]) ^ (layer0_outputs[3520]);
    assign layer1_outputs[11044] = ~(layer0_outputs[12705]);
    assign layer1_outputs[11045] = (layer0_outputs[1999]) & ~(layer0_outputs[11515]);
    assign layer1_outputs[11046] = (layer0_outputs[4629]) & (layer0_outputs[11392]);
    assign layer1_outputs[11047] = (layer0_outputs[5942]) & ~(layer0_outputs[6183]);
    assign layer1_outputs[11048] = ~(layer0_outputs[872]) | (layer0_outputs[10239]);
    assign layer1_outputs[11049] = layer0_outputs[7615];
    assign layer1_outputs[11050] = layer0_outputs[503];
    assign layer1_outputs[11051] = layer0_outputs[4321];
    assign layer1_outputs[11052] = layer0_outputs[6380];
    assign layer1_outputs[11053] = ~(layer0_outputs[2669]);
    assign layer1_outputs[11054] = layer0_outputs[12619];
    assign layer1_outputs[11055] = ~((layer0_outputs[8987]) & (layer0_outputs[5522]));
    assign layer1_outputs[11056] = ~(layer0_outputs[1799]);
    assign layer1_outputs[11057] = ~(layer0_outputs[10866]);
    assign layer1_outputs[11058] = (layer0_outputs[4026]) ^ (layer0_outputs[11716]);
    assign layer1_outputs[11059] = ~((layer0_outputs[3149]) | (layer0_outputs[4284]));
    assign layer1_outputs[11060] = ~(layer0_outputs[1018]);
    assign layer1_outputs[11061] = (layer0_outputs[3696]) ^ (layer0_outputs[6724]);
    assign layer1_outputs[11062] = ~(layer0_outputs[6582]);
    assign layer1_outputs[11063] = (layer0_outputs[2522]) | (layer0_outputs[10017]);
    assign layer1_outputs[11064] = (layer0_outputs[2444]) ^ (layer0_outputs[802]);
    assign layer1_outputs[11065] = ~(layer0_outputs[1584]) | (layer0_outputs[551]);
    assign layer1_outputs[11066] = (layer0_outputs[8739]) & ~(layer0_outputs[2508]);
    assign layer1_outputs[11067] = ~(layer0_outputs[4536]);
    assign layer1_outputs[11068] = ~((layer0_outputs[6616]) & (layer0_outputs[5259]));
    assign layer1_outputs[11069] = ~(layer0_outputs[11705]) | (layer0_outputs[5262]);
    assign layer1_outputs[11070] = (layer0_outputs[81]) ^ (layer0_outputs[8058]);
    assign layer1_outputs[11071] = (layer0_outputs[3845]) & (layer0_outputs[6595]);
    assign layer1_outputs[11072] = ~((layer0_outputs[6550]) & (layer0_outputs[7733]));
    assign layer1_outputs[11073] = ~(layer0_outputs[4263]);
    assign layer1_outputs[11074] = ~((layer0_outputs[11324]) ^ (layer0_outputs[9361]));
    assign layer1_outputs[11075] = (layer0_outputs[3832]) ^ (layer0_outputs[11397]);
    assign layer1_outputs[11076] = layer0_outputs[10806];
    assign layer1_outputs[11077] = (layer0_outputs[3885]) ^ (layer0_outputs[12531]);
    assign layer1_outputs[11078] = (layer0_outputs[6277]) ^ (layer0_outputs[8829]);
    assign layer1_outputs[11079] = ~(layer0_outputs[8996]);
    assign layer1_outputs[11080] = ~(layer0_outputs[3145]) | (layer0_outputs[7789]);
    assign layer1_outputs[11081] = (layer0_outputs[8113]) & ~(layer0_outputs[9236]);
    assign layer1_outputs[11082] = (layer0_outputs[11152]) & ~(layer0_outputs[8645]);
    assign layer1_outputs[11083] = ~(layer0_outputs[7135]);
    assign layer1_outputs[11084] = 1'b1;
    assign layer1_outputs[11085] = layer0_outputs[3231];
    assign layer1_outputs[11086] = ~((layer0_outputs[8275]) & (layer0_outputs[11665]));
    assign layer1_outputs[11087] = (layer0_outputs[10435]) & ~(layer0_outputs[9510]);
    assign layer1_outputs[11088] = ~(layer0_outputs[11408]) | (layer0_outputs[3009]);
    assign layer1_outputs[11089] = ~(layer0_outputs[1090]);
    assign layer1_outputs[11090] = (layer0_outputs[7760]) & ~(layer0_outputs[5732]);
    assign layer1_outputs[11091] = (layer0_outputs[10461]) & ~(layer0_outputs[3128]);
    assign layer1_outputs[11092] = (layer0_outputs[10141]) & ~(layer0_outputs[7432]);
    assign layer1_outputs[11093] = layer0_outputs[2045];
    assign layer1_outputs[11094] = layer0_outputs[11825];
    assign layer1_outputs[11095] = (layer0_outputs[1350]) ^ (layer0_outputs[5995]);
    assign layer1_outputs[11096] = layer0_outputs[2775];
    assign layer1_outputs[11097] = (layer0_outputs[10247]) ^ (layer0_outputs[2315]);
    assign layer1_outputs[11098] = ~(layer0_outputs[3088]) | (layer0_outputs[68]);
    assign layer1_outputs[11099] = layer0_outputs[10399];
    assign layer1_outputs[11100] = layer0_outputs[12285];
    assign layer1_outputs[11101] = layer0_outputs[5523];
    assign layer1_outputs[11102] = ~(layer0_outputs[7072]) | (layer0_outputs[11975]);
    assign layer1_outputs[11103] = (layer0_outputs[7079]) & ~(layer0_outputs[1737]);
    assign layer1_outputs[11104] = (layer0_outputs[2735]) ^ (layer0_outputs[4002]);
    assign layer1_outputs[11105] = ~(layer0_outputs[3501]);
    assign layer1_outputs[11106] = layer0_outputs[9888];
    assign layer1_outputs[11107] = layer0_outputs[10241];
    assign layer1_outputs[11108] = ~((layer0_outputs[2541]) ^ (layer0_outputs[3478]));
    assign layer1_outputs[11109] = ~(layer0_outputs[7624]) | (layer0_outputs[9622]);
    assign layer1_outputs[11110] = ~(layer0_outputs[8642]) | (layer0_outputs[10638]);
    assign layer1_outputs[11111] = ~(layer0_outputs[939]) | (layer0_outputs[1408]);
    assign layer1_outputs[11112] = ~(layer0_outputs[10042]) | (layer0_outputs[318]);
    assign layer1_outputs[11113] = (layer0_outputs[8351]) & (layer0_outputs[719]);
    assign layer1_outputs[11114] = ~((layer0_outputs[10107]) ^ (layer0_outputs[7435]));
    assign layer1_outputs[11115] = ~((layer0_outputs[3897]) ^ (layer0_outputs[11371]));
    assign layer1_outputs[11116] = ~((layer0_outputs[1691]) & (layer0_outputs[7880]));
    assign layer1_outputs[11117] = ~(layer0_outputs[10052]);
    assign layer1_outputs[11118] = ~(layer0_outputs[5551]);
    assign layer1_outputs[11119] = ~(layer0_outputs[8955]) | (layer0_outputs[1138]);
    assign layer1_outputs[11120] = ~((layer0_outputs[6052]) | (layer0_outputs[8511]));
    assign layer1_outputs[11121] = (layer0_outputs[8798]) & ~(layer0_outputs[9436]);
    assign layer1_outputs[11122] = (layer0_outputs[3860]) & ~(layer0_outputs[10513]);
    assign layer1_outputs[11123] = layer0_outputs[104];
    assign layer1_outputs[11124] = ~((layer0_outputs[2120]) ^ (layer0_outputs[7069]));
    assign layer1_outputs[11125] = layer0_outputs[9686];
    assign layer1_outputs[11126] = layer0_outputs[9537];
    assign layer1_outputs[11127] = (layer0_outputs[11257]) & ~(layer0_outputs[9060]);
    assign layer1_outputs[11128] = (layer0_outputs[2771]) & (layer0_outputs[10168]);
    assign layer1_outputs[11129] = ~((layer0_outputs[10208]) & (layer0_outputs[7741]));
    assign layer1_outputs[11130] = ~(layer0_outputs[2262]);
    assign layer1_outputs[11131] = layer0_outputs[6448];
    assign layer1_outputs[11132] = ~(layer0_outputs[12439]) | (layer0_outputs[11325]);
    assign layer1_outputs[11133] = (layer0_outputs[6044]) | (layer0_outputs[10690]);
    assign layer1_outputs[11134] = ~((layer0_outputs[292]) | (layer0_outputs[6097]));
    assign layer1_outputs[11135] = layer0_outputs[11239];
    assign layer1_outputs[11136] = (layer0_outputs[11202]) & (layer0_outputs[9723]);
    assign layer1_outputs[11137] = ~((layer0_outputs[4302]) | (layer0_outputs[8176]));
    assign layer1_outputs[11138] = ~(layer0_outputs[6279]) | (layer0_outputs[10805]);
    assign layer1_outputs[11139] = (layer0_outputs[8056]) ^ (layer0_outputs[4719]);
    assign layer1_outputs[11140] = (layer0_outputs[6677]) | (layer0_outputs[9986]);
    assign layer1_outputs[11141] = ~(layer0_outputs[7525]);
    assign layer1_outputs[11142] = ~(layer0_outputs[8504]);
    assign layer1_outputs[11143] = layer0_outputs[10210];
    assign layer1_outputs[11144] = ~(layer0_outputs[6029]);
    assign layer1_outputs[11145] = layer0_outputs[1013];
    assign layer1_outputs[11146] = ~((layer0_outputs[4979]) & (layer0_outputs[1557]));
    assign layer1_outputs[11147] = layer0_outputs[3893];
    assign layer1_outputs[11148] = (layer0_outputs[5233]) & ~(layer0_outputs[9961]);
    assign layer1_outputs[11149] = (layer0_outputs[1739]) & ~(layer0_outputs[2297]);
    assign layer1_outputs[11150] = ~(layer0_outputs[10003]);
    assign layer1_outputs[11151] = (layer0_outputs[4209]) & ~(layer0_outputs[10150]);
    assign layer1_outputs[11152] = (layer0_outputs[11109]) & ~(layer0_outputs[12742]);
    assign layer1_outputs[11153] = ~(layer0_outputs[3665]);
    assign layer1_outputs[11154] = (layer0_outputs[7202]) ^ (layer0_outputs[9507]);
    assign layer1_outputs[11155] = ~((layer0_outputs[9062]) ^ (layer0_outputs[7042]));
    assign layer1_outputs[11156] = layer0_outputs[8373];
    assign layer1_outputs[11157] = ~(layer0_outputs[6053]);
    assign layer1_outputs[11158] = ~(layer0_outputs[6324]);
    assign layer1_outputs[11159] = ~(layer0_outputs[8615]) | (layer0_outputs[10457]);
    assign layer1_outputs[11160] = (layer0_outputs[4493]) & (layer0_outputs[524]);
    assign layer1_outputs[11161] = layer0_outputs[2019];
    assign layer1_outputs[11162] = ~((layer0_outputs[10117]) | (layer0_outputs[8966]));
    assign layer1_outputs[11163] = ~(layer0_outputs[1977]) | (layer0_outputs[1482]);
    assign layer1_outputs[11164] = layer0_outputs[2542];
    assign layer1_outputs[11165] = (layer0_outputs[9258]) & ~(layer0_outputs[4881]);
    assign layer1_outputs[11166] = ~((layer0_outputs[7533]) & (layer0_outputs[43]));
    assign layer1_outputs[11167] = ~(layer0_outputs[12559]);
    assign layer1_outputs[11168] = (layer0_outputs[4755]) & ~(layer0_outputs[10830]);
    assign layer1_outputs[11169] = (layer0_outputs[11509]) & ~(layer0_outputs[2321]);
    assign layer1_outputs[11170] = (layer0_outputs[11264]) | (layer0_outputs[9002]);
    assign layer1_outputs[11171] = ~((layer0_outputs[1425]) & (layer0_outputs[3158]));
    assign layer1_outputs[11172] = layer0_outputs[4106];
    assign layer1_outputs[11173] = layer0_outputs[9730];
    assign layer1_outputs[11174] = ~(layer0_outputs[8454]);
    assign layer1_outputs[11175] = (layer0_outputs[12628]) & ~(layer0_outputs[7450]);
    assign layer1_outputs[11176] = ~(layer0_outputs[5329]);
    assign layer1_outputs[11177] = ~(layer0_outputs[1661]) | (layer0_outputs[9599]);
    assign layer1_outputs[11178] = ~((layer0_outputs[12212]) ^ (layer0_outputs[1482]));
    assign layer1_outputs[11179] = ~((layer0_outputs[6198]) & (layer0_outputs[9073]));
    assign layer1_outputs[11180] = layer0_outputs[3386];
    assign layer1_outputs[11181] = 1'b1;
    assign layer1_outputs[11182] = (layer0_outputs[270]) ^ (layer0_outputs[1308]);
    assign layer1_outputs[11183] = ~(layer0_outputs[11403]) | (layer0_outputs[10121]);
    assign layer1_outputs[11184] = (layer0_outputs[4130]) & ~(layer0_outputs[9496]);
    assign layer1_outputs[11185] = ~(layer0_outputs[3797]);
    assign layer1_outputs[11186] = ~(layer0_outputs[4838]) | (layer0_outputs[9273]);
    assign layer1_outputs[11187] = ~((layer0_outputs[1475]) ^ (layer0_outputs[9224]));
    assign layer1_outputs[11188] = layer0_outputs[1052];
    assign layer1_outputs[11189] = layer0_outputs[3471];
    assign layer1_outputs[11190] = (layer0_outputs[6381]) | (layer0_outputs[11523]);
    assign layer1_outputs[11191] = ~((layer0_outputs[12616]) | (layer0_outputs[11181]));
    assign layer1_outputs[11192] = 1'b0;
    assign layer1_outputs[11193] = 1'b1;
    assign layer1_outputs[11194] = ~((layer0_outputs[173]) ^ (layer0_outputs[7797]));
    assign layer1_outputs[11195] = ~((layer0_outputs[10928]) | (layer0_outputs[2467]));
    assign layer1_outputs[11196] = layer0_outputs[10447];
    assign layer1_outputs[11197] = ~((layer0_outputs[3063]) ^ (layer0_outputs[11920]));
    assign layer1_outputs[11198] = layer0_outputs[804];
    assign layer1_outputs[11199] = (layer0_outputs[11736]) ^ (layer0_outputs[4278]);
    assign layer1_outputs[11200] = (layer0_outputs[12251]) ^ (layer0_outputs[9398]);
    assign layer1_outputs[11201] = (layer0_outputs[5659]) & ~(layer0_outputs[12284]);
    assign layer1_outputs[11202] = ~(layer0_outputs[3533]) | (layer0_outputs[634]);
    assign layer1_outputs[11203] = layer0_outputs[5071];
    assign layer1_outputs[11204] = ~(layer0_outputs[7173]);
    assign layer1_outputs[11205] = (layer0_outputs[9971]) & (layer0_outputs[2821]);
    assign layer1_outputs[11206] = ~(layer0_outputs[1747]) | (layer0_outputs[4221]);
    assign layer1_outputs[11207] = 1'b0;
    assign layer1_outputs[11208] = ~(layer0_outputs[5430]);
    assign layer1_outputs[11209] = ~((layer0_outputs[2236]) ^ (layer0_outputs[12750]));
    assign layer1_outputs[11210] = ~(layer0_outputs[10425]);
    assign layer1_outputs[11211] = (layer0_outputs[3691]) | (layer0_outputs[4418]);
    assign layer1_outputs[11212] = ~((layer0_outputs[12764]) | (layer0_outputs[10839]));
    assign layer1_outputs[11213] = ~((layer0_outputs[6511]) | (layer0_outputs[8686]));
    assign layer1_outputs[11214] = (layer0_outputs[6471]) | (layer0_outputs[1092]);
    assign layer1_outputs[11215] = ~(layer0_outputs[8360]);
    assign layer1_outputs[11216] = layer0_outputs[4243];
    assign layer1_outputs[11217] = 1'b0;
    assign layer1_outputs[11218] = ~((layer0_outputs[3693]) & (layer0_outputs[11613]));
    assign layer1_outputs[11219] = (layer0_outputs[6183]) | (layer0_outputs[9225]);
    assign layer1_outputs[11220] = ~((layer0_outputs[4076]) & (layer0_outputs[7795]));
    assign layer1_outputs[11221] = layer0_outputs[1836];
    assign layer1_outputs[11222] = layer0_outputs[1420];
    assign layer1_outputs[11223] = (layer0_outputs[10849]) & ~(layer0_outputs[1744]);
    assign layer1_outputs[11224] = (layer0_outputs[2436]) | (layer0_outputs[5954]);
    assign layer1_outputs[11225] = ~(layer0_outputs[6510]);
    assign layer1_outputs[11226] = (layer0_outputs[4479]) & (layer0_outputs[11436]);
    assign layer1_outputs[11227] = ~((layer0_outputs[9931]) ^ (layer0_outputs[220]));
    assign layer1_outputs[11228] = 1'b1;
    assign layer1_outputs[11229] = (layer0_outputs[10088]) | (layer0_outputs[5175]);
    assign layer1_outputs[11230] = (layer0_outputs[2863]) ^ (layer0_outputs[4849]);
    assign layer1_outputs[11231] = ~(layer0_outputs[4744]);
    assign layer1_outputs[11232] = (layer0_outputs[7333]) & ~(layer0_outputs[7328]);
    assign layer1_outputs[11233] = ~(layer0_outputs[8975]) | (layer0_outputs[12164]);
    assign layer1_outputs[11234] = ~(layer0_outputs[2600]);
    assign layer1_outputs[11235] = ~(layer0_outputs[3736]);
    assign layer1_outputs[11236] = (layer0_outputs[1142]) & ~(layer0_outputs[4400]);
    assign layer1_outputs[11237] = ~(layer0_outputs[430]);
    assign layer1_outputs[11238] = ~(layer0_outputs[8756]) | (layer0_outputs[12677]);
    assign layer1_outputs[11239] = (layer0_outputs[10470]) & ~(layer0_outputs[7572]);
    assign layer1_outputs[11240] = layer0_outputs[11760];
    assign layer1_outputs[11241] = ~(layer0_outputs[6296]);
    assign layer1_outputs[11242] = ~((layer0_outputs[9483]) | (layer0_outputs[3925]));
    assign layer1_outputs[11243] = layer0_outputs[9984];
    assign layer1_outputs[11244] = ~(layer0_outputs[4340]) | (layer0_outputs[1295]);
    assign layer1_outputs[11245] = ~(layer0_outputs[7964]) | (layer0_outputs[8783]);
    assign layer1_outputs[11246] = ~((layer0_outputs[7700]) & (layer0_outputs[7448]));
    assign layer1_outputs[11247] = ~((layer0_outputs[8258]) | (layer0_outputs[2947]));
    assign layer1_outputs[11248] = (layer0_outputs[3042]) ^ (layer0_outputs[3901]);
    assign layer1_outputs[11249] = ~(layer0_outputs[2929]);
    assign layer1_outputs[11250] = ~(layer0_outputs[8941]);
    assign layer1_outputs[11251] = layer0_outputs[11316];
    assign layer1_outputs[11252] = ~(layer0_outputs[4870]) | (layer0_outputs[9845]);
    assign layer1_outputs[11253] = layer0_outputs[8208];
    assign layer1_outputs[11254] = (layer0_outputs[1003]) | (layer0_outputs[7790]);
    assign layer1_outputs[11255] = (layer0_outputs[3498]) & ~(layer0_outputs[12059]);
    assign layer1_outputs[11256] = layer0_outputs[8775];
    assign layer1_outputs[11257] = (layer0_outputs[5604]) & ~(layer0_outputs[11772]);
    assign layer1_outputs[11258] = layer0_outputs[2008];
    assign layer1_outputs[11259] = ~((layer0_outputs[9779]) & (layer0_outputs[8726]));
    assign layer1_outputs[11260] = 1'b1;
    assign layer1_outputs[11261] = 1'b0;
    assign layer1_outputs[11262] = 1'b1;
    assign layer1_outputs[11263] = 1'b0;
    assign layer1_outputs[11264] = ~(layer0_outputs[4250]);
    assign layer1_outputs[11265] = (layer0_outputs[11638]) | (layer0_outputs[8140]);
    assign layer1_outputs[11266] = ~(layer0_outputs[6796]);
    assign layer1_outputs[11267] = layer0_outputs[12006];
    assign layer1_outputs[11268] = ~(layer0_outputs[5827]) | (layer0_outputs[10232]);
    assign layer1_outputs[11269] = layer0_outputs[7385];
    assign layer1_outputs[11270] = (layer0_outputs[2440]) ^ (layer0_outputs[10831]);
    assign layer1_outputs[11271] = ~((layer0_outputs[419]) & (layer0_outputs[2429]));
    assign layer1_outputs[11272] = ~(layer0_outputs[3171]);
    assign layer1_outputs[11273] = (layer0_outputs[2344]) | (layer0_outputs[8868]);
    assign layer1_outputs[11274] = ~((layer0_outputs[4200]) & (layer0_outputs[8164]));
    assign layer1_outputs[11275] = (layer0_outputs[11943]) & ~(layer0_outputs[7452]);
    assign layer1_outputs[11276] = (layer0_outputs[5446]) & ~(layer0_outputs[7514]);
    assign layer1_outputs[11277] = (layer0_outputs[1951]) | (layer0_outputs[386]);
    assign layer1_outputs[11278] = ~(layer0_outputs[395]) | (layer0_outputs[3582]);
    assign layer1_outputs[11279] = ~(layer0_outputs[1520]);
    assign layer1_outputs[11280] = ~(layer0_outputs[3064]);
    assign layer1_outputs[11281] = layer0_outputs[8942];
    assign layer1_outputs[11282] = (layer0_outputs[10675]) & ~(layer0_outputs[6810]);
    assign layer1_outputs[11283] = ~(layer0_outputs[2572]);
    assign layer1_outputs[11284] = (layer0_outputs[1512]) ^ (layer0_outputs[11761]);
    assign layer1_outputs[11285] = (layer0_outputs[7029]) | (layer0_outputs[8251]);
    assign layer1_outputs[11286] = ~(layer0_outputs[7706]);
    assign layer1_outputs[11287] = ~((layer0_outputs[3827]) & (layer0_outputs[4870]));
    assign layer1_outputs[11288] = 1'b0;
    assign layer1_outputs[11289] = ~(layer0_outputs[12003]);
    assign layer1_outputs[11290] = (layer0_outputs[4426]) | (layer0_outputs[11866]);
    assign layer1_outputs[11291] = ~((layer0_outputs[616]) | (layer0_outputs[980]));
    assign layer1_outputs[11292] = layer0_outputs[10319];
    assign layer1_outputs[11293] = (layer0_outputs[3272]) & ~(layer0_outputs[4557]);
    assign layer1_outputs[11294] = ~((layer0_outputs[6716]) & (layer0_outputs[5889]));
    assign layer1_outputs[11295] = (layer0_outputs[3929]) & ~(layer0_outputs[5805]);
    assign layer1_outputs[11296] = (layer0_outputs[8602]) ^ (layer0_outputs[4024]);
    assign layer1_outputs[11297] = layer0_outputs[6331];
    assign layer1_outputs[11298] = (layer0_outputs[6084]) ^ (layer0_outputs[1128]);
    assign layer1_outputs[11299] = 1'b1;
    assign layer1_outputs[11300] = ~(layer0_outputs[1463]) | (layer0_outputs[2098]);
    assign layer1_outputs[11301] = ~((layer0_outputs[383]) | (layer0_outputs[12143]));
    assign layer1_outputs[11302] = 1'b0;
    assign layer1_outputs[11303] = ~((layer0_outputs[8502]) ^ (layer0_outputs[7850]));
    assign layer1_outputs[11304] = (layer0_outputs[555]) | (layer0_outputs[10339]);
    assign layer1_outputs[11305] = (layer0_outputs[1118]) & ~(layer0_outputs[3267]);
    assign layer1_outputs[11306] = ~((layer0_outputs[7265]) & (layer0_outputs[8576]));
    assign layer1_outputs[11307] = layer0_outputs[12216];
    assign layer1_outputs[11308] = ~((layer0_outputs[10858]) ^ (layer0_outputs[10161]));
    assign layer1_outputs[11309] = ~((layer0_outputs[10704]) & (layer0_outputs[11078]));
    assign layer1_outputs[11310] = ~(layer0_outputs[10677]);
    assign layer1_outputs[11311] = (layer0_outputs[12513]) | (layer0_outputs[6216]);
    assign layer1_outputs[11312] = ~(layer0_outputs[236]) | (layer0_outputs[7103]);
    assign layer1_outputs[11313] = (layer0_outputs[3095]) & ~(layer0_outputs[1934]);
    assign layer1_outputs[11314] = (layer0_outputs[3199]) ^ (layer0_outputs[2230]);
    assign layer1_outputs[11315] = (layer0_outputs[3219]) & ~(layer0_outputs[1602]);
    assign layer1_outputs[11316] = (layer0_outputs[10919]) & ~(layer0_outputs[10891]);
    assign layer1_outputs[11317] = ~((layer0_outputs[11721]) | (layer0_outputs[1751]));
    assign layer1_outputs[11318] = ~(layer0_outputs[2092]) | (layer0_outputs[6661]);
    assign layer1_outputs[11319] = ~(layer0_outputs[11051]);
    assign layer1_outputs[11320] = ~((layer0_outputs[6081]) ^ (layer0_outputs[9732]));
    assign layer1_outputs[11321] = ~(layer0_outputs[2129]);
    assign layer1_outputs[11322] = ~(layer0_outputs[10749]);
    assign layer1_outputs[11323] = ~((layer0_outputs[6849]) ^ (layer0_outputs[8095]));
    assign layer1_outputs[11324] = (layer0_outputs[3436]) ^ (layer0_outputs[11275]);
    assign layer1_outputs[11325] = ~(layer0_outputs[10954]);
    assign layer1_outputs[11326] = ~(layer0_outputs[1235]) | (layer0_outputs[4185]);
    assign layer1_outputs[11327] = ~(layer0_outputs[11011]) | (layer0_outputs[4947]);
    assign layer1_outputs[11328] = ~(layer0_outputs[11980]);
    assign layer1_outputs[11329] = ~((layer0_outputs[5961]) & (layer0_outputs[12588]));
    assign layer1_outputs[11330] = layer0_outputs[9499];
    assign layer1_outputs[11331] = (layer0_outputs[4148]) & ~(layer0_outputs[9475]);
    assign layer1_outputs[11332] = ~((layer0_outputs[9980]) | (layer0_outputs[3528]));
    assign layer1_outputs[11333] = layer0_outputs[11887];
    assign layer1_outputs[11334] = ~(layer0_outputs[9776]) | (layer0_outputs[1078]);
    assign layer1_outputs[11335] = ~((layer0_outputs[6405]) & (layer0_outputs[9655]));
    assign layer1_outputs[11336] = (layer0_outputs[9061]) & ~(layer0_outputs[1956]);
    assign layer1_outputs[11337] = ~(layer0_outputs[2953]);
    assign layer1_outputs[11338] = (layer0_outputs[8455]) | (layer0_outputs[4014]);
    assign layer1_outputs[11339] = (layer0_outputs[6192]) & ~(layer0_outputs[4463]);
    assign layer1_outputs[11340] = (layer0_outputs[2487]) & (layer0_outputs[11095]);
    assign layer1_outputs[11341] = layer0_outputs[5951];
    assign layer1_outputs[11342] = layer0_outputs[8287];
    assign layer1_outputs[11343] = (layer0_outputs[23]) & ~(layer0_outputs[7753]);
    assign layer1_outputs[11344] = (layer0_outputs[8365]) & ~(layer0_outputs[4312]);
    assign layer1_outputs[11345] = ~((layer0_outputs[4131]) & (layer0_outputs[5536]));
    assign layer1_outputs[11346] = layer0_outputs[3635];
    assign layer1_outputs[11347] = ~((layer0_outputs[4568]) | (layer0_outputs[8226]));
    assign layer1_outputs[11348] = ~(layer0_outputs[8230]);
    assign layer1_outputs[11349] = layer0_outputs[4796];
    assign layer1_outputs[11350] = ~(layer0_outputs[3331]);
    assign layer1_outputs[11351] = layer0_outputs[6989];
    assign layer1_outputs[11352] = (layer0_outputs[1238]) | (layer0_outputs[8316]);
    assign layer1_outputs[11353] = ~((layer0_outputs[9404]) & (layer0_outputs[4827]));
    assign layer1_outputs[11354] = ~((layer0_outputs[7436]) & (layer0_outputs[8069]));
    assign layer1_outputs[11355] = ~(layer0_outputs[7393]);
    assign layer1_outputs[11356] = ~(layer0_outputs[301]);
    assign layer1_outputs[11357] = (layer0_outputs[10001]) ^ (layer0_outputs[333]);
    assign layer1_outputs[11358] = (layer0_outputs[10038]) & ~(layer0_outputs[5965]);
    assign layer1_outputs[11359] = layer0_outputs[10380];
    assign layer1_outputs[11360] = ~(layer0_outputs[2801]);
    assign layer1_outputs[11361] = ~(layer0_outputs[738]);
    assign layer1_outputs[11362] = (layer0_outputs[9891]) ^ (layer0_outputs[9965]);
    assign layer1_outputs[11363] = ~((layer0_outputs[8406]) | (layer0_outputs[3817]));
    assign layer1_outputs[11364] = layer0_outputs[6222];
    assign layer1_outputs[11365] = 1'b1;
    assign layer1_outputs[11366] = (layer0_outputs[10651]) & ~(layer0_outputs[4634]);
    assign layer1_outputs[11367] = (layer0_outputs[10643]) ^ (layer0_outputs[9454]);
    assign layer1_outputs[11368] = (layer0_outputs[12473]) | (layer0_outputs[10925]);
    assign layer1_outputs[11369] = layer0_outputs[3318];
    assign layer1_outputs[11370] = (layer0_outputs[11227]) & ~(layer0_outputs[5130]);
    assign layer1_outputs[11371] = (layer0_outputs[10690]) ^ (layer0_outputs[7221]);
    assign layer1_outputs[11372] = layer0_outputs[4510];
    assign layer1_outputs[11373] = (layer0_outputs[4981]) ^ (layer0_outputs[12116]);
    assign layer1_outputs[11374] = ~(layer0_outputs[10614]);
    assign layer1_outputs[11375] = ~(layer0_outputs[5886]);
    assign layer1_outputs[11376] = layer0_outputs[4260];
    assign layer1_outputs[11377] = layer0_outputs[7125];
    assign layer1_outputs[11378] = ~(layer0_outputs[6922]) | (layer0_outputs[2890]);
    assign layer1_outputs[11379] = ~(layer0_outputs[4083]);
    assign layer1_outputs[11380] = ~(layer0_outputs[8066]) | (layer0_outputs[9168]);
    assign layer1_outputs[11381] = layer0_outputs[1822];
    assign layer1_outputs[11382] = ~(layer0_outputs[1567]) | (layer0_outputs[8500]);
    assign layer1_outputs[11383] = ~((layer0_outputs[5606]) & (layer0_outputs[4128]));
    assign layer1_outputs[11384] = (layer0_outputs[560]) & ~(layer0_outputs[7551]);
    assign layer1_outputs[11385] = ~(layer0_outputs[11027]) | (layer0_outputs[1974]);
    assign layer1_outputs[11386] = (layer0_outputs[6916]) & ~(layer0_outputs[8978]);
    assign layer1_outputs[11387] = ~(layer0_outputs[267]) | (layer0_outputs[10351]);
    assign layer1_outputs[11388] = (layer0_outputs[4319]) & ~(layer0_outputs[8571]);
    assign layer1_outputs[11389] = 1'b0;
    assign layer1_outputs[11390] = (layer0_outputs[531]) & ~(layer0_outputs[3594]);
    assign layer1_outputs[11391] = ~((layer0_outputs[3846]) & (layer0_outputs[6253]));
    assign layer1_outputs[11392] = ~((layer0_outputs[6117]) | (layer0_outputs[3983]));
    assign layer1_outputs[11393] = (layer0_outputs[4273]) | (layer0_outputs[6344]);
    assign layer1_outputs[11394] = layer0_outputs[8296];
    assign layer1_outputs[11395] = 1'b0;
    assign layer1_outputs[11396] = ~(layer0_outputs[6831]);
    assign layer1_outputs[11397] = (layer0_outputs[214]) & ~(layer0_outputs[3083]);
    assign layer1_outputs[11398] = ~((layer0_outputs[6174]) & (layer0_outputs[10801]));
    assign layer1_outputs[11399] = layer0_outputs[12474];
    assign layer1_outputs[11400] = (layer0_outputs[684]) & (layer0_outputs[8414]);
    assign layer1_outputs[11401] = layer0_outputs[11076];
    assign layer1_outputs[11402] = (layer0_outputs[4757]) | (layer0_outputs[3366]);
    assign layer1_outputs[11403] = ~((layer0_outputs[9176]) & (layer0_outputs[10044]));
    assign layer1_outputs[11404] = layer0_outputs[7439];
    assign layer1_outputs[11405] = ~(layer0_outputs[1982]);
    assign layer1_outputs[11406] = 1'b0;
    assign layer1_outputs[11407] = layer0_outputs[8492];
    assign layer1_outputs[11408] = ~(layer0_outputs[8171]) | (layer0_outputs[12676]);
    assign layer1_outputs[11409] = ~(layer0_outputs[11410]) | (layer0_outputs[11046]);
    assign layer1_outputs[11410] = ~(layer0_outputs[7681]);
    assign layer1_outputs[11411] = layer0_outputs[5531];
    assign layer1_outputs[11412] = (layer0_outputs[312]) & ~(layer0_outputs[7570]);
    assign layer1_outputs[11413] = ~(layer0_outputs[11181]) | (layer0_outputs[3790]);
    assign layer1_outputs[11414] = (layer0_outputs[216]) & ~(layer0_outputs[4129]);
    assign layer1_outputs[11415] = ~(layer0_outputs[8011]) | (layer0_outputs[3507]);
    assign layer1_outputs[11416] = (layer0_outputs[11569]) & ~(layer0_outputs[12434]);
    assign layer1_outputs[11417] = ~((layer0_outputs[6970]) ^ (layer0_outputs[5481]));
    assign layer1_outputs[11418] = (layer0_outputs[4601]) | (layer0_outputs[11628]);
    assign layer1_outputs[11419] = (layer0_outputs[3213]) & ~(layer0_outputs[3470]);
    assign layer1_outputs[11420] = layer0_outputs[12114];
    assign layer1_outputs[11421] = layer0_outputs[588];
    assign layer1_outputs[11422] = ~(layer0_outputs[2831]);
    assign layer1_outputs[11423] = (layer0_outputs[2300]) | (layer0_outputs[5709]);
    assign layer1_outputs[11424] = layer0_outputs[3079];
    assign layer1_outputs[11425] = ~(layer0_outputs[2573]);
    assign layer1_outputs[11426] = layer0_outputs[10157];
    assign layer1_outputs[11427] = ~((layer0_outputs[10336]) ^ (layer0_outputs[4445]));
    assign layer1_outputs[11428] = layer0_outputs[1219];
    assign layer1_outputs[11429] = (layer0_outputs[143]) & ~(layer0_outputs[11273]);
    assign layer1_outputs[11430] = layer0_outputs[4610];
    assign layer1_outputs[11431] = ~(layer0_outputs[7111]) | (layer0_outputs[12243]);
    assign layer1_outputs[11432] = (layer0_outputs[2899]) | (layer0_outputs[1453]);
    assign layer1_outputs[11433] = 1'b0;
    assign layer1_outputs[11434] = (layer0_outputs[11670]) & ~(layer0_outputs[9875]);
    assign layer1_outputs[11435] = (layer0_outputs[3049]) & ~(layer0_outputs[11349]);
    assign layer1_outputs[11436] = 1'b1;
    assign layer1_outputs[11437] = ~(layer0_outputs[10455]) | (layer0_outputs[5064]);
    assign layer1_outputs[11438] = (layer0_outputs[4471]) ^ (layer0_outputs[12342]);
    assign layer1_outputs[11439] = layer0_outputs[2562];
    assign layer1_outputs[11440] = (layer0_outputs[10025]) & (layer0_outputs[5927]);
    assign layer1_outputs[11441] = layer0_outputs[2429];
    assign layer1_outputs[11442] = layer0_outputs[752];
    assign layer1_outputs[11443] = ~((layer0_outputs[1234]) & (layer0_outputs[832]));
    assign layer1_outputs[11444] = ~(layer0_outputs[3548]);
    assign layer1_outputs[11445] = ~(layer0_outputs[5107]) | (layer0_outputs[10670]);
    assign layer1_outputs[11446] = layer0_outputs[11972];
    assign layer1_outputs[11447] = ~(layer0_outputs[7168]);
    assign layer1_outputs[11448] = ~(layer0_outputs[2547]);
    assign layer1_outputs[11449] = ~(layer0_outputs[2425]);
    assign layer1_outputs[11450] = ~(layer0_outputs[11506]) | (layer0_outputs[8787]);
    assign layer1_outputs[11451] = layer0_outputs[6105];
    assign layer1_outputs[11452] = 1'b0;
    assign layer1_outputs[11453] = (layer0_outputs[6055]) & ~(layer0_outputs[3961]);
    assign layer1_outputs[11454] = (layer0_outputs[10975]) & ~(layer0_outputs[2918]);
    assign layer1_outputs[11455] = ~(layer0_outputs[2529]);
    assign layer1_outputs[11456] = (layer0_outputs[4669]) | (layer0_outputs[6909]);
    assign layer1_outputs[11457] = 1'b1;
    assign layer1_outputs[11458] = (layer0_outputs[10046]) ^ (layer0_outputs[3361]);
    assign layer1_outputs[11459] = ~(layer0_outputs[11111]);
    assign layer1_outputs[11460] = ~(layer0_outputs[1465]) | (layer0_outputs[10055]);
    assign layer1_outputs[11461] = ~((layer0_outputs[11653]) | (layer0_outputs[5467]));
    assign layer1_outputs[11462] = ~((layer0_outputs[7673]) & (layer0_outputs[2940]));
    assign layer1_outputs[11463] = ~(layer0_outputs[1035]) | (layer0_outputs[7635]);
    assign layer1_outputs[11464] = (layer0_outputs[11983]) ^ (layer0_outputs[8233]);
    assign layer1_outputs[11465] = ~(layer0_outputs[10092]);
    assign layer1_outputs[11466] = (layer0_outputs[8116]) & ~(layer0_outputs[4054]);
    assign layer1_outputs[11467] = ~(layer0_outputs[7938]) | (layer0_outputs[12234]);
    assign layer1_outputs[11468] = ~(layer0_outputs[6654]);
    assign layer1_outputs[11469] = (layer0_outputs[9319]) | (layer0_outputs[9084]);
    assign layer1_outputs[11470] = layer0_outputs[8976];
    assign layer1_outputs[11471] = (layer0_outputs[4957]) & ~(layer0_outputs[8862]);
    assign layer1_outputs[11472] = layer0_outputs[9572];
    assign layer1_outputs[11473] = (layer0_outputs[4544]) ^ (layer0_outputs[1862]);
    assign layer1_outputs[11474] = ~(layer0_outputs[10800]) | (layer0_outputs[153]);
    assign layer1_outputs[11475] = ~((layer0_outputs[12196]) ^ (layer0_outputs[9294]));
    assign layer1_outputs[11476] = layer0_outputs[5589];
    assign layer1_outputs[11477] = layer0_outputs[6242];
    assign layer1_outputs[11478] = layer0_outputs[1249];
    assign layer1_outputs[11479] = (layer0_outputs[11723]) ^ (layer0_outputs[8301]);
    assign layer1_outputs[11480] = ~(layer0_outputs[6253]);
    assign layer1_outputs[11481] = ~(layer0_outputs[922]) | (layer0_outputs[9950]);
    assign layer1_outputs[11482] = layer0_outputs[7658];
    assign layer1_outputs[11483] = layer0_outputs[786];
    assign layer1_outputs[11484] = (layer0_outputs[10879]) ^ (layer0_outputs[9930]);
    assign layer1_outputs[11485] = (layer0_outputs[1042]) ^ (layer0_outputs[8323]);
    assign layer1_outputs[11486] = ~((layer0_outputs[4210]) & (layer0_outputs[8101]));
    assign layer1_outputs[11487] = layer0_outputs[2410];
    assign layer1_outputs[11488] = ~(layer0_outputs[7147]) | (layer0_outputs[11614]);
    assign layer1_outputs[11489] = layer0_outputs[2517];
    assign layer1_outputs[11490] = ~((layer0_outputs[5802]) ^ (layer0_outputs[2951]));
    assign layer1_outputs[11491] = ~(layer0_outputs[12075]);
    assign layer1_outputs[11492] = (layer0_outputs[9962]) & ~(layer0_outputs[7745]);
    assign layer1_outputs[11493] = ~(layer0_outputs[6764]) | (layer0_outputs[982]);
    assign layer1_outputs[11494] = ~(layer0_outputs[4447]);
    assign layer1_outputs[11495] = ~((layer0_outputs[1659]) ^ (layer0_outputs[12687]));
    assign layer1_outputs[11496] = (layer0_outputs[11782]) ^ (layer0_outputs[467]);
    assign layer1_outputs[11497] = (layer0_outputs[1057]) & ~(layer0_outputs[7331]);
    assign layer1_outputs[11498] = ~(layer0_outputs[11234]);
    assign layer1_outputs[11499] = layer0_outputs[11354];
    assign layer1_outputs[11500] = layer0_outputs[6234];
    assign layer1_outputs[11501] = ~((layer0_outputs[334]) ^ (layer0_outputs[5498]));
    assign layer1_outputs[11502] = ~(layer0_outputs[7755]) | (layer0_outputs[835]);
    assign layer1_outputs[11503] = ~(layer0_outputs[7489]);
    assign layer1_outputs[11504] = ~(layer0_outputs[2738]) | (layer0_outputs[2989]);
    assign layer1_outputs[11505] = layer0_outputs[11382];
    assign layer1_outputs[11506] = layer0_outputs[12291];
    assign layer1_outputs[11507] = ~(layer0_outputs[7062]);
    assign layer1_outputs[11508] = layer0_outputs[6670];
    assign layer1_outputs[11509] = ~(layer0_outputs[12378]);
    assign layer1_outputs[11510] = ~((layer0_outputs[11293]) & (layer0_outputs[6370]));
    assign layer1_outputs[11511] = (layer0_outputs[12764]) & ~(layer0_outputs[3557]);
    assign layer1_outputs[11512] = (layer0_outputs[1157]) & (layer0_outputs[9918]);
    assign layer1_outputs[11513] = (layer0_outputs[12490]) ^ (layer0_outputs[2314]);
    assign layer1_outputs[11514] = ~(layer0_outputs[305]) | (layer0_outputs[9154]);
    assign layer1_outputs[11515] = (layer0_outputs[6509]) & ~(layer0_outputs[12552]);
    assign layer1_outputs[11516] = layer0_outputs[7800];
    assign layer1_outputs[11517] = 1'b1;
    assign layer1_outputs[11518] = 1'b0;
    assign layer1_outputs[11519] = (layer0_outputs[9698]) & ~(layer0_outputs[11563]);
    assign layer1_outputs[11520] = layer0_outputs[2578];
    assign layer1_outputs[11521] = ~(layer0_outputs[1554]);
    assign layer1_outputs[11522] = (layer0_outputs[12033]) | (layer0_outputs[2304]);
    assign layer1_outputs[11523] = (layer0_outputs[4385]) & ~(layer0_outputs[2527]);
    assign layer1_outputs[11524] = ~((layer0_outputs[9668]) ^ (layer0_outputs[1838]));
    assign layer1_outputs[11525] = ~(layer0_outputs[8359]);
    assign layer1_outputs[11526] = layer0_outputs[3323];
    assign layer1_outputs[11527] = ~(layer0_outputs[2195]);
    assign layer1_outputs[11528] = layer0_outputs[6064];
    assign layer1_outputs[11529] = (layer0_outputs[1431]) | (layer0_outputs[7303]);
    assign layer1_outputs[11530] = (layer0_outputs[9808]) & ~(layer0_outputs[859]);
    assign layer1_outputs[11531] = ~(layer0_outputs[8389]);
    assign layer1_outputs[11532] = (layer0_outputs[2911]) | (layer0_outputs[5947]);
    assign layer1_outputs[11533] = ~((layer0_outputs[810]) & (layer0_outputs[514]));
    assign layer1_outputs[11534] = ~(layer0_outputs[615]) | (layer0_outputs[2976]);
    assign layer1_outputs[11535] = ~((layer0_outputs[1272]) & (layer0_outputs[12488]));
    assign layer1_outputs[11536] = ~((layer0_outputs[5736]) ^ (layer0_outputs[5543]));
    assign layer1_outputs[11537] = ~((layer0_outputs[12732]) & (layer0_outputs[8444]));
    assign layer1_outputs[11538] = ~(layer0_outputs[8709]);
    assign layer1_outputs[11539] = ~(layer0_outputs[9907]) | (layer0_outputs[9009]);
    assign layer1_outputs[11540] = ~(layer0_outputs[169]) | (layer0_outputs[4000]);
    assign layer1_outputs[11541] = ~(layer0_outputs[2830]);
    assign layer1_outputs[11542] = ~((layer0_outputs[1684]) & (layer0_outputs[7182]));
    assign layer1_outputs[11543] = layer0_outputs[9920];
    assign layer1_outputs[11544] = ~(layer0_outputs[7003]) | (layer0_outputs[9939]);
    assign layer1_outputs[11545] = ~((layer0_outputs[320]) | (layer0_outputs[11780]));
    assign layer1_outputs[11546] = layer0_outputs[7256];
    assign layer1_outputs[11547] = ~(layer0_outputs[8165]);
    assign layer1_outputs[11548] = layer0_outputs[669];
    assign layer1_outputs[11549] = ~((layer0_outputs[6009]) & (layer0_outputs[4966]));
    assign layer1_outputs[11550] = ~(layer0_outputs[5393]);
    assign layer1_outputs[11551] = ~(layer0_outputs[5073]);
    assign layer1_outputs[11552] = ~(layer0_outputs[8654]);
    assign layer1_outputs[11553] = ~(layer0_outputs[4553]);
    assign layer1_outputs[11554] = (layer0_outputs[1745]) & ~(layer0_outputs[9206]);
    assign layer1_outputs[11555] = layer0_outputs[6456];
    assign layer1_outputs[11556] = ~((layer0_outputs[1435]) ^ (layer0_outputs[1970]));
    assign layer1_outputs[11557] = ~(layer0_outputs[5356]) | (layer0_outputs[9917]);
    assign layer1_outputs[11558] = (layer0_outputs[4181]) ^ (layer0_outputs[6065]);
    assign layer1_outputs[11559] = ~(layer0_outputs[4872]);
    assign layer1_outputs[11560] = layer0_outputs[11811];
    assign layer1_outputs[11561] = ~((layer0_outputs[3913]) & (layer0_outputs[1785]));
    assign layer1_outputs[11562] = layer0_outputs[7404];
    assign layer1_outputs[11563] = (layer0_outputs[4500]) | (layer0_outputs[8944]);
    assign layer1_outputs[11564] = ~(layer0_outputs[1409]);
    assign layer1_outputs[11565] = (layer0_outputs[879]) | (layer0_outputs[3808]);
    assign layer1_outputs[11566] = (layer0_outputs[2221]) ^ (layer0_outputs[7802]);
    assign layer1_outputs[11567] = (layer0_outputs[885]) & ~(layer0_outputs[10061]);
    assign layer1_outputs[11568] = layer0_outputs[3303];
    assign layer1_outputs[11569] = ~((layer0_outputs[1558]) | (layer0_outputs[11732]));
    assign layer1_outputs[11570] = ~(layer0_outputs[1915]) | (layer0_outputs[12198]);
    assign layer1_outputs[11571] = ~((layer0_outputs[6374]) | (layer0_outputs[8419]));
    assign layer1_outputs[11572] = layer0_outputs[5881];
    assign layer1_outputs[11573] = 1'b0;
    assign layer1_outputs[11574] = layer0_outputs[5482];
    assign layer1_outputs[11575] = ~((layer0_outputs[85]) ^ (layer0_outputs[7789]));
    assign layer1_outputs[11576] = layer0_outputs[7475];
    assign layer1_outputs[11577] = (layer0_outputs[7150]) & (layer0_outputs[7973]);
    assign layer1_outputs[11578] = layer0_outputs[6113];
    assign layer1_outputs[11579] = (layer0_outputs[10165]) | (layer0_outputs[11084]);
    assign layer1_outputs[11580] = layer0_outputs[6785];
    assign layer1_outputs[11581] = (layer0_outputs[9330]) & (layer0_outputs[11293]);
    assign layer1_outputs[11582] = ~((layer0_outputs[3933]) & (layer0_outputs[1714]));
    assign layer1_outputs[11583] = ~(layer0_outputs[5119]);
    assign layer1_outputs[11584] = ~(layer0_outputs[7946]);
    assign layer1_outputs[11585] = (layer0_outputs[3545]) ^ (layer0_outputs[5549]);
    assign layer1_outputs[11586] = (layer0_outputs[9721]) & (layer0_outputs[4118]);
    assign layer1_outputs[11587] = ~((layer0_outputs[5979]) | (layer0_outputs[5660]));
    assign layer1_outputs[11588] = layer0_outputs[929];
    assign layer1_outputs[11589] = ~(layer0_outputs[12555]) | (layer0_outputs[10671]);
    assign layer1_outputs[11590] = layer0_outputs[11408];
    assign layer1_outputs[11591] = ~(layer0_outputs[2076]);
    assign layer1_outputs[11592] = ~((layer0_outputs[953]) | (layer0_outputs[7921]));
    assign layer1_outputs[11593] = layer0_outputs[1696];
    assign layer1_outputs[11594] = (layer0_outputs[4970]) & (layer0_outputs[12399]);
    assign layer1_outputs[11595] = ~(layer0_outputs[1762]);
    assign layer1_outputs[11596] = (layer0_outputs[9272]) | (layer0_outputs[3966]);
    assign layer1_outputs[11597] = (layer0_outputs[10624]) ^ (layer0_outputs[5943]);
    assign layer1_outputs[11598] = 1'b0;
    assign layer1_outputs[11599] = ~((layer0_outputs[6074]) & (layer0_outputs[9484]));
    assign layer1_outputs[11600] = (layer0_outputs[7242]) ^ (layer0_outputs[10799]);
    assign layer1_outputs[11601] = (layer0_outputs[12532]) & (layer0_outputs[7793]);
    assign layer1_outputs[11602] = ~((layer0_outputs[5463]) & (layer0_outputs[5592]));
    assign layer1_outputs[11603] = layer0_outputs[3697];
    assign layer1_outputs[11604] = ~(layer0_outputs[3856]) | (layer0_outputs[5472]);
    assign layer1_outputs[11605] = (layer0_outputs[9503]) ^ (layer0_outputs[8062]);
    assign layer1_outputs[11606] = (layer0_outputs[6102]) & ~(layer0_outputs[2386]);
    assign layer1_outputs[11607] = (layer0_outputs[132]) & ~(layer0_outputs[2585]);
    assign layer1_outputs[11608] = layer0_outputs[10492];
    assign layer1_outputs[11609] = ~((layer0_outputs[5695]) ^ (layer0_outputs[4305]));
    assign layer1_outputs[11610] = (layer0_outputs[10646]) & ~(layer0_outputs[9581]);
    assign layer1_outputs[11611] = ~(layer0_outputs[4404]);
    assign layer1_outputs[11612] = layer0_outputs[7346];
    assign layer1_outputs[11613] = (layer0_outputs[12046]) ^ (layer0_outputs[372]);
    assign layer1_outputs[11614] = (layer0_outputs[7314]) ^ (layer0_outputs[12345]);
    assign layer1_outputs[11615] = ~((layer0_outputs[5100]) ^ (layer0_outputs[3063]));
    assign layer1_outputs[11616] = layer0_outputs[1183];
    assign layer1_outputs[11617] = (layer0_outputs[12671]) & ~(layer0_outputs[6509]);
    assign layer1_outputs[11618] = ~(layer0_outputs[3241]);
    assign layer1_outputs[11619] = ~(layer0_outputs[8119]);
    assign layer1_outputs[11620] = ~(layer0_outputs[10885]);
    assign layer1_outputs[11621] = (layer0_outputs[11089]) & ~(layer0_outputs[6604]);
    assign layer1_outputs[11622] = ~((layer0_outputs[1591]) & (layer0_outputs[233]));
    assign layer1_outputs[11623] = ~(layer0_outputs[10124]);
    assign layer1_outputs[11624] = ~(layer0_outputs[709]);
    assign layer1_outputs[11625] = ~((layer0_outputs[9489]) ^ (layer0_outputs[10421]));
    assign layer1_outputs[11626] = layer0_outputs[9079];
    assign layer1_outputs[11627] = ~((layer0_outputs[6692]) & (layer0_outputs[2053]));
    assign layer1_outputs[11628] = layer0_outputs[4811];
    assign layer1_outputs[11629] = layer0_outputs[11661];
    assign layer1_outputs[11630] = ~(layer0_outputs[6313]);
    assign layer1_outputs[11631] = layer0_outputs[8267];
    assign layer1_outputs[11632] = layer0_outputs[1748];
    assign layer1_outputs[11633] = (layer0_outputs[8723]) & ~(layer0_outputs[4334]);
    assign layer1_outputs[11634] = (layer0_outputs[8918]) & ~(layer0_outputs[11484]);
    assign layer1_outputs[11635] = ~((layer0_outputs[6296]) | (layer0_outputs[6089]));
    assign layer1_outputs[11636] = ~(layer0_outputs[1795]);
    assign layer1_outputs[11637] = (layer0_outputs[3259]) & (layer0_outputs[5403]);
    assign layer1_outputs[11638] = (layer0_outputs[10266]) & ~(layer0_outputs[8449]);
    assign layer1_outputs[11639] = layer0_outputs[3518];
    assign layer1_outputs[11640] = ~((layer0_outputs[4596]) ^ (layer0_outputs[2733]));
    assign layer1_outputs[11641] = (layer0_outputs[8147]) | (layer0_outputs[8963]);
    assign layer1_outputs[11642] = layer0_outputs[5978];
    assign layer1_outputs[11643] = ~(layer0_outputs[7459]);
    assign layer1_outputs[11644] = ~(layer0_outputs[5199]);
    assign layer1_outputs[11645] = layer0_outputs[5789];
    assign layer1_outputs[11646] = ~((layer0_outputs[11396]) ^ (layer0_outputs[4719]));
    assign layer1_outputs[11647] = 1'b0;
    assign layer1_outputs[11648] = ~(layer0_outputs[6392]) | (layer0_outputs[4511]);
    assign layer1_outputs[11649] = ~(layer0_outputs[2157]);
    assign layer1_outputs[11650] = ~(layer0_outputs[6457]);
    assign layer1_outputs[11651] = layer0_outputs[10406];
    assign layer1_outputs[11652] = ~((layer0_outputs[2337]) | (layer0_outputs[1551]));
    assign layer1_outputs[11653] = ~(layer0_outputs[3245]);
    assign layer1_outputs[11654] = ~(layer0_outputs[14]);
    assign layer1_outputs[11655] = ~(layer0_outputs[258]);
    assign layer1_outputs[11656] = ~((layer0_outputs[343]) & (layer0_outputs[2689]));
    assign layer1_outputs[11657] = ~(layer0_outputs[2694]);
    assign layer1_outputs[11658] = ~((layer0_outputs[11026]) ^ (layer0_outputs[11422]));
    assign layer1_outputs[11659] = layer0_outputs[1858];
    assign layer1_outputs[11660] = layer0_outputs[1703];
    assign layer1_outputs[11661] = ~((layer0_outputs[5707]) & (layer0_outputs[4961]));
    assign layer1_outputs[11662] = (layer0_outputs[8856]) ^ (layer0_outputs[6982]);
    assign layer1_outputs[11663] = ~(layer0_outputs[12042]);
    assign layer1_outputs[11664] = ~(layer0_outputs[11579]);
    assign layer1_outputs[11665] = ~((layer0_outputs[3777]) ^ (layer0_outputs[12773]));
    assign layer1_outputs[11666] = ~(layer0_outputs[2771]);
    assign layer1_outputs[11667] = ~(layer0_outputs[5365]);
    assign layer1_outputs[11668] = ~(layer0_outputs[4935]) | (layer0_outputs[5343]);
    assign layer1_outputs[11669] = layer0_outputs[1421];
    assign layer1_outputs[11670] = (layer0_outputs[12458]) & ~(layer0_outputs[8878]);
    assign layer1_outputs[11671] = ~((layer0_outputs[4626]) & (layer0_outputs[974]));
    assign layer1_outputs[11672] = layer0_outputs[756];
    assign layer1_outputs[11673] = ~(layer0_outputs[1474]);
    assign layer1_outputs[11674] = layer0_outputs[2959];
    assign layer1_outputs[11675] = layer0_outputs[11929];
    assign layer1_outputs[11676] = layer0_outputs[1917];
    assign layer1_outputs[11677] = ~((layer0_outputs[7862]) | (layer0_outputs[2581]));
    assign layer1_outputs[11678] = (layer0_outputs[9431]) & (layer0_outputs[1824]);
    assign layer1_outputs[11679] = ~(layer0_outputs[141]) | (layer0_outputs[727]);
    assign layer1_outputs[11680] = ~(layer0_outputs[2498]);
    assign layer1_outputs[11681] = (layer0_outputs[9588]) & (layer0_outputs[8169]);
    assign layer1_outputs[11682] = layer0_outputs[6747];
    assign layer1_outputs[11683] = ~((layer0_outputs[9131]) ^ (layer0_outputs[2636]));
    assign layer1_outputs[11684] = ~(layer0_outputs[3850]);
    assign layer1_outputs[11685] = ~((layer0_outputs[9227]) & (layer0_outputs[12250]));
    assign layer1_outputs[11686] = (layer0_outputs[12450]) & ~(layer0_outputs[8358]);
    assign layer1_outputs[11687] = ~((layer0_outputs[10250]) & (layer0_outputs[9287]));
    assign layer1_outputs[11688] = layer0_outputs[12036];
    assign layer1_outputs[11689] = ~(layer0_outputs[5285]);
    assign layer1_outputs[11690] = layer0_outputs[12551];
    assign layer1_outputs[11691] = ~(layer0_outputs[5311]);
    assign layer1_outputs[11692] = (layer0_outputs[2735]) | (layer0_outputs[2012]);
    assign layer1_outputs[11693] = layer0_outputs[8306];
    assign layer1_outputs[11694] = ~((layer0_outputs[4179]) ^ (layer0_outputs[7351]));
    assign layer1_outputs[11695] = (layer0_outputs[5245]) & (layer0_outputs[6421]);
    assign layer1_outputs[11696] = ~(layer0_outputs[1597]) | (layer0_outputs[4750]);
    assign layer1_outputs[11697] = layer0_outputs[10495];
    assign layer1_outputs[11698] = ~(layer0_outputs[6309]) | (layer0_outputs[7833]);
    assign layer1_outputs[11699] = (layer0_outputs[4867]) | (layer0_outputs[5668]);
    assign layer1_outputs[11700] = (layer0_outputs[3896]) | (layer0_outputs[616]);
    assign layer1_outputs[11701] = ~(layer0_outputs[1367]);
    assign layer1_outputs[11702] = layer0_outputs[12082];
    assign layer1_outputs[11703] = ~(layer0_outputs[9375]);
    assign layer1_outputs[11704] = ~(layer0_outputs[9046]) | (layer0_outputs[2204]);
    assign layer1_outputs[11705] = ~(layer0_outputs[11351]);
    assign layer1_outputs[11706] = layer0_outputs[7777];
    assign layer1_outputs[11707] = ~(layer0_outputs[455]);
    assign layer1_outputs[11708] = ~(layer0_outputs[7356]);
    assign layer1_outputs[11709] = layer0_outputs[9760];
    assign layer1_outputs[11710] = (layer0_outputs[11725]) & ~(layer0_outputs[5380]);
    assign layer1_outputs[11711] = ~(layer0_outputs[5786]);
    assign layer1_outputs[11712] = layer0_outputs[10965];
    assign layer1_outputs[11713] = (layer0_outputs[9237]) & ~(layer0_outputs[8617]);
    assign layer1_outputs[11714] = layer0_outputs[11641];
    assign layer1_outputs[11715] = (layer0_outputs[8232]) ^ (layer0_outputs[6712]);
    assign layer1_outputs[11716] = ~((layer0_outputs[9897]) ^ (layer0_outputs[9048]));
    assign layer1_outputs[11717] = ~(layer0_outputs[5366]);
    assign layer1_outputs[11718] = (layer0_outputs[6850]) & ~(layer0_outputs[4227]);
    assign layer1_outputs[11719] = layer0_outputs[3334];
    assign layer1_outputs[11720] = (layer0_outputs[5215]) & ~(layer0_outputs[5541]);
    assign layer1_outputs[11721] = ~(layer0_outputs[1597]) | (layer0_outputs[7817]);
    assign layer1_outputs[11722] = ~((layer0_outputs[12402]) | (layer0_outputs[808]));
    assign layer1_outputs[11723] = ~(layer0_outputs[10511]);
    assign layer1_outputs[11724] = (layer0_outputs[3766]) & (layer0_outputs[2601]);
    assign layer1_outputs[11725] = layer0_outputs[2619];
    assign layer1_outputs[11726] = (layer0_outputs[11416]) & ~(layer0_outputs[3464]);
    assign layer1_outputs[11727] = layer0_outputs[4311];
    assign layer1_outputs[11728] = (layer0_outputs[3522]) & ~(layer0_outputs[8828]);
    assign layer1_outputs[11729] = layer0_outputs[12673];
    assign layer1_outputs[11730] = (layer0_outputs[2279]) & (layer0_outputs[2834]);
    assign layer1_outputs[11731] = ~(layer0_outputs[2589]);
    assign layer1_outputs[11732] = ~(layer0_outputs[7232]) | (layer0_outputs[1114]);
    assign layer1_outputs[11733] = ~((layer0_outputs[1137]) & (layer0_outputs[7022]));
    assign layer1_outputs[11734] = ~(layer0_outputs[3838]) | (layer0_outputs[1783]);
    assign layer1_outputs[11735] = ~(layer0_outputs[1764]) | (layer0_outputs[8998]);
    assign layer1_outputs[11736] = layer0_outputs[10329];
    assign layer1_outputs[11737] = ~(layer0_outputs[3129]) | (layer0_outputs[876]);
    assign layer1_outputs[11738] = (layer0_outputs[11859]) | (layer0_outputs[4368]);
    assign layer1_outputs[11739] = ~((layer0_outputs[4008]) ^ (layer0_outputs[4721]));
    assign layer1_outputs[11740] = (layer0_outputs[3315]) ^ (layer0_outputs[8545]);
    assign layer1_outputs[11741] = (layer0_outputs[8578]) & (layer0_outputs[12333]);
    assign layer1_outputs[11742] = ~((layer0_outputs[373]) ^ (layer0_outputs[6804]));
    assign layer1_outputs[11743] = (layer0_outputs[1351]) & ~(layer0_outputs[8442]);
    assign layer1_outputs[11744] = ~(layer0_outputs[8741]);
    assign layer1_outputs[11745] = layer0_outputs[4963];
    assign layer1_outputs[11746] = (layer0_outputs[9251]) & ~(layer0_outputs[5609]);
    assign layer1_outputs[11747] = ~(layer0_outputs[3430]) | (layer0_outputs[3454]);
    assign layer1_outputs[11748] = layer0_outputs[8567];
    assign layer1_outputs[11749] = ~((layer0_outputs[12785]) ^ (layer0_outputs[7744]));
    assign layer1_outputs[11750] = (layer0_outputs[5173]) & (layer0_outputs[3605]);
    assign layer1_outputs[11751] = ~(layer0_outputs[7407]);
    assign layer1_outputs[11752] = layer0_outputs[215];
    assign layer1_outputs[11753] = ~(layer0_outputs[8441]) | (layer0_outputs[5852]);
    assign layer1_outputs[11754] = ~(layer0_outputs[6211]);
    assign layer1_outputs[11755] = ~(layer0_outputs[9360]) | (layer0_outputs[7689]);
    assign layer1_outputs[11756] = ~(layer0_outputs[10537]) | (layer0_outputs[3056]);
    assign layer1_outputs[11757] = ~((layer0_outputs[2836]) ^ (layer0_outputs[11576]));
    assign layer1_outputs[11758] = ~((layer0_outputs[2151]) | (layer0_outputs[6097]));
    assign layer1_outputs[11759] = (layer0_outputs[1976]) & (layer0_outputs[2736]);
    assign layer1_outputs[11760] = 1'b1;
    assign layer1_outputs[11761] = ~(layer0_outputs[11906]) | (layer0_outputs[6258]);
    assign layer1_outputs[11762] = layer0_outputs[3457];
    assign layer1_outputs[11763] = ~(layer0_outputs[3350]);
    assign layer1_outputs[11764] = layer0_outputs[11559];
    assign layer1_outputs[11765] = ~((layer0_outputs[5736]) & (layer0_outputs[86]));
    assign layer1_outputs[11766] = ~((layer0_outputs[1109]) ^ (layer0_outputs[6077]));
    assign layer1_outputs[11767] = layer0_outputs[10166];
    assign layer1_outputs[11768] = ~(layer0_outputs[4997]);
    assign layer1_outputs[11769] = ~(layer0_outputs[5547]) | (layer0_outputs[7279]);
    assign layer1_outputs[11770] = ~(layer0_outputs[9341]);
    assign layer1_outputs[11771] = ~((layer0_outputs[8554]) | (layer0_outputs[7839]));
    assign layer1_outputs[11772] = ~(layer0_outputs[2805]);
    assign layer1_outputs[11773] = (layer0_outputs[6925]) & ~(layer0_outputs[2796]);
    assign layer1_outputs[11774] = layer0_outputs[4975];
    assign layer1_outputs[11775] = layer0_outputs[272];
    assign layer1_outputs[11776] = layer0_outputs[10522];
    assign layer1_outputs[11777] = 1'b0;
    assign layer1_outputs[11778] = (layer0_outputs[4556]) ^ (layer0_outputs[4018]);
    assign layer1_outputs[11779] = layer0_outputs[7286];
    assign layer1_outputs[11780] = ~(layer0_outputs[7167]) | (layer0_outputs[2290]);
    assign layer1_outputs[11781] = layer0_outputs[9634];
    assign layer1_outputs[11782] = (layer0_outputs[2763]) & ~(layer0_outputs[10419]);
    assign layer1_outputs[11783] = ~(layer0_outputs[11401]);
    assign layer1_outputs[11784] = (layer0_outputs[1254]) & ~(layer0_outputs[346]);
    assign layer1_outputs[11785] = (layer0_outputs[11428]) ^ (layer0_outputs[8885]);
    assign layer1_outputs[11786] = (layer0_outputs[8356]) & ~(layer0_outputs[3457]);
    assign layer1_outputs[11787] = ~(layer0_outputs[4675]);
    assign layer1_outputs[11788] = layer0_outputs[5008];
    assign layer1_outputs[11789] = (layer0_outputs[10105]) & (layer0_outputs[64]);
    assign layer1_outputs[11790] = (layer0_outputs[4834]) | (layer0_outputs[12385]);
    assign layer1_outputs[11791] = ~((layer0_outputs[7647]) ^ (layer0_outputs[8573]));
    assign layer1_outputs[11792] = (layer0_outputs[6318]) ^ (layer0_outputs[11327]);
    assign layer1_outputs[11793] = (layer0_outputs[6226]) & ~(layer0_outputs[4806]);
    assign layer1_outputs[11794] = (layer0_outputs[9974]) | (layer0_outputs[1925]);
    assign layer1_outputs[11795] = 1'b1;
    assign layer1_outputs[11796] = ~((layer0_outputs[3054]) & (layer0_outputs[11021]));
    assign layer1_outputs[11797] = layer0_outputs[6440];
    assign layer1_outputs[11798] = (layer0_outputs[18]) & (layer0_outputs[8271]);
    assign layer1_outputs[11799] = layer0_outputs[4731];
    assign layer1_outputs[11800] = ~((layer0_outputs[8811]) | (layer0_outputs[5811]));
    assign layer1_outputs[11801] = ~(layer0_outputs[2033]);
    assign layer1_outputs[11802] = (layer0_outputs[7502]) | (layer0_outputs[8830]);
    assign layer1_outputs[11803] = ~(layer0_outputs[7403]);
    assign layer1_outputs[11804] = layer0_outputs[1989];
    assign layer1_outputs[11805] = (layer0_outputs[2857]) ^ (layer0_outputs[122]);
    assign layer1_outputs[11806] = layer0_outputs[2228];
    assign layer1_outputs[11807] = layer0_outputs[6271];
    assign layer1_outputs[11808] = ~((layer0_outputs[7199]) | (layer0_outputs[11653]));
    assign layer1_outputs[11809] = layer0_outputs[12222];
    assign layer1_outputs[11810] = ~(layer0_outputs[11347]);
    assign layer1_outputs[11811] = ~(layer0_outputs[9153]) | (layer0_outputs[2207]);
    assign layer1_outputs[11812] = ~(layer0_outputs[6667]) | (layer0_outputs[2714]);
    assign layer1_outputs[11813] = layer0_outputs[7];
    assign layer1_outputs[11814] = ~((layer0_outputs[4405]) | (layer0_outputs[8281]));
    assign layer1_outputs[11815] = (layer0_outputs[8467]) & ~(layer0_outputs[10693]);
    assign layer1_outputs[11816] = ~(layer0_outputs[9803]) | (layer0_outputs[4074]);
    assign layer1_outputs[11817] = ~(layer0_outputs[7931]);
    assign layer1_outputs[11818] = ~((layer0_outputs[3308]) ^ (layer0_outputs[3871]));
    assign layer1_outputs[11819] = ~(layer0_outputs[9388]);
    assign layer1_outputs[11820] = (layer0_outputs[9270]) & ~(layer0_outputs[10627]);
    assign layer1_outputs[11821] = ~(layer0_outputs[803]) | (layer0_outputs[10332]);
    assign layer1_outputs[11822] = (layer0_outputs[1080]) | (layer0_outputs[3381]);
    assign layer1_outputs[11823] = layer0_outputs[4639];
    assign layer1_outputs[11824] = ~((layer0_outputs[9034]) | (layer0_outputs[309]));
    assign layer1_outputs[11825] = (layer0_outputs[10669]) & ~(layer0_outputs[2139]);
    assign layer1_outputs[11826] = (layer0_outputs[8764]) & ~(layer0_outputs[6508]);
    assign layer1_outputs[11827] = layer0_outputs[5353];
    assign layer1_outputs[11828] = layer0_outputs[225];
    assign layer1_outputs[11829] = ~((layer0_outputs[6150]) ^ (layer0_outputs[11377]));
    assign layer1_outputs[11830] = ~(layer0_outputs[11976]) | (layer0_outputs[8779]);
    assign layer1_outputs[11831] = ~(layer0_outputs[4595]) | (layer0_outputs[7482]);
    assign layer1_outputs[11832] = (layer0_outputs[12034]) & ~(layer0_outputs[2734]);
    assign layer1_outputs[11833] = (layer0_outputs[10378]) & ~(layer0_outputs[547]);
    assign layer1_outputs[11834] = ~((layer0_outputs[548]) | (layer0_outputs[10108]));
    assign layer1_outputs[11835] = 1'b1;
    assign layer1_outputs[11836] = ~((layer0_outputs[4978]) | (layer0_outputs[12301]));
    assign layer1_outputs[11837] = (layer0_outputs[114]) | (layer0_outputs[3679]);
    assign layer1_outputs[11838] = (layer0_outputs[6346]) & (layer0_outputs[9045]);
    assign layer1_outputs[11839] = (layer0_outputs[2519]) & ~(layer0_outputs[10539]);
    assign layer1_outputs[11840] = ~((layer0_outputs[10118]) | (layer0_outputs[1162]));
    assign layer1_outputs[11841] = ~((layer0_outputs[12541]) | (layer0_outputs[12408]));
    assign layer1_outputs[11842] = ~(layer0_outputs[4351]) | (layer0_outputs[2228]);
    assign layer1_outputs[11843] = ~((layer0_outputs[6387]) & (layer0_outputs[8366]));
    assign layer1_outputs[11844] = layer0_outputs[5015];
    assign layer1_outputs[11845] = ~((layer0_outputs[6233]) & (layer0_outputs[10510]));
    assign layer1_outputs[11846] = ~(layer0_outputs[11333]);
    assign layer1_outputs[11847] = layer0_outputs[5374];
    assign layer1_outputs[11848] = layer0_outputs[2178];
    assign layer1_outputs[11849] = (layer0_outputs[8407]) & ~(layer0_outputs[8476]);
    assign layer1_outputs[11850] = (layer0_outputs[9384]) | (layer0_outputs[6567]);
    assign layer1_outputs[11851] = ~(layer0_outputs[6175]);
    assign layer1_outputs[11852] = ~((layer0_outputs[7760]) ^ (layer0_outputs[5993]));
    assign layer1_outputs[11853] = (layer0_outputs[4846]) & ~(layer0_outputs[5621]);
    assign layer1_outputs[11854] = ~((layer0_outputs[4502]) | (layer0_outputs[9028]));
    assign layer1_outputs[11855] = ~((layer0_outputs[7402]) & (layer0_outputs[6723]));
    assign layer1_outputs[11856] = (layer0_outputs[6310]) | (layer0_outputs[10566]);
    assign layer1_outputs[11857] = ~((layer0_outputs[4555]) & (layer0_outputs[5428]));
    assign layer1_outputs[11858] = ~(layer0_outputs[12175]) | (layer0_outputs[6783]);
    assign layer1_outputs[11859] = ~(layer0_outputs[8951]);
    assign layer1_outputs[11860] = ~((layer0_outputs[541]) | (layer0_outputs[3410]));
    assign layer1_outputs[11861] = ~((layer0_outputs[7074]) ^ (layer0_outputs[1998]));
    assign layer1_outputs[11862] = ~((layer0_outputs[8905]) | (layer0_outputs[7559]));
    assign layer1_outputs[11863] = (layer0_outputs[2710]) & (layer0_outputs[10715]);
    assign layer1_outputs[11864] = ~(layer0_outputs[4080]);
    assign layer1_outputs[11865] = layer0_outputs[886];
    assign layer1_outputs[11866] = (layer0_outputs[12062]) ^ (layer0_outputs[6683]);
    assign layer1_outputs[11867] = ~(layer0_outputs[712]) | (layer0_outputs[7780]);
    assign layer1_outputs[11868] = ~(layer0_outputs[11060]) | (layer0_outputs[11670]);
    assign layer1_outputs[11869] = ~((layer0_outputs[10997]) ^ (layer0_outputs[8137]));
    assign layer1_outputs[11870] = ~(layer0_outputs[231]) | (layer0_outputs[2181]);
    assign layer1_outputs[11871] = (layer0_outputs[12172]) & (layer0_outputs[12152]);
    assign layer1_outputs[11872] = (layer0_outputs[3987]) | (layer0_outputs[10819]);
    assign layer1_outputs[11873] = (layer0_outputs[7530]) & ~(layer0_outputs[1876]);
    assign layer1_outputs[11874] = layer0_outputs[634];
    assign layer1_outputs[11875] = ~((layer0_outputs[6597]) ^ (layer0_outputs[5618]));
    assign layer1_outputs[11876] = (layer0_outputs[3106]) | (layer0_outputs[5127]);
    assign layer1_outputs[11877] = ~(layer0_outputs[296]);
    assign layer1_outputs[11878] = ~(layer0_outputs[4603]) | (layer0_outputs[9580]);
    assign layer1_outputs[11879] = ~((layer0_outputs[3022]) | (layer0_outputs[1452]));
    assign layer1_outputs[11880] = ~(layer0_outputs[9493]);
    assign layer1_outputs[11881] = ~((layer0_outputs[3731]) & (layer0_outputs[3408]));
    assign layer1_outputs[11882] = ~(layer0_outputs[4286]);
    assign layer1_outputs[11883] = ~(layer0_outputs[7413]);
    assign layer1_outputs[11884] = layer0_outputs[4316];
    assign layer1_outputs[11885] = ~(layer0_outputs[9433]);
    assign layer1_outputs[11886] = layer0_outputs[8815];
    assign layer1_outputs[11887] = ~((layer0_outputs[6972]) | (layer0_outputs[3754]));
    assign layer1_outputs[11888] = layer0_outputs[11996];
    assign layer1_outputs[11889] = ~(layer0_outputs[11513]);
    assign layer1_outputs[11890] = layer0_outputs[7806];
    assign layer1_outputs[11891] = ~(layer0_outputs[4741]) | (layer0_outputs[6847]);
    assign layer1_outputs[11892] = (layer0_outputs[9927]) | (layer0_outputs[829]);
    assign layer1_outputs[11893] = ~((layer0_outputs[6850]) ^ (layer0_outputs[4584]));
    assign layer1_outputs[11894] = (layer0_outputs[10691]) ^ (layer0_outputs[546]);
    assign layer1_outputs[11895] = layer0_outputs[8515];
    assign layer1_outputs[11896] = ~(layer0_outputs[8410]);
    assign layer1_outputs[11897] = (layer0_outputs[5810]) | (layer0_outputs[5124]);
    assign layer1_outputs[11898] = (layer0_outputs[2356]) & ~(layer0_outputs[5599]);
    assign layer1_outputs[11899] = (layer0_outputs[952]) & (layer0_outputs[8782]);
    assign layer1_outputs[11900] = (layer0_outputs[125]) & ~(layer0_outputs[2435]);
    assign layer1_outputs[11901] = layer0_outputs[469];
    assign layer1_outputs[11902] = layer0_outputs[11284];
    assign layer1_outputs[11903] = ~((layer0_outputs[8221]) & (layer0_outputs[79]));
    assign layer1_outputs[11904] = layer0_outputs[1281];
    assign layer1_outputs[11905] = ~(layer0_outputs[10159]);
    assign layer1_outputs[11906] = ~(layer0_outputs[4891]);
    assign layer1_outputs[11907] = ~((layer0_outputs[12341]) | (layer0_outputs[9374]));
    assign layer1_outputs[11908] = (layer0_outputs[8706]) & (layer0_outputs[12160]);
    assign layer1_outputs[11909] = (layer0_outputs[5968]) & ~(layer0_outputs[5532]);
    assign layer1_outputs[11910] = ~(layer0_outputs[940]);
    assign layer1_outputs[11911] = ~(layer0_outputs[845]);
    assign layer1_outputs[11912] = ~((layer0_outputs[7865]) | (layer0_outputs[6173]));
    assign layer1_outputs[11913] = ~(layer0_outputs[499]);
    assign layer1_outputs[11914] = layer0_outputs[11844];
    assign layer1_outputs[11915] = (layer0_outputs[3449]) & ~(layer0_outputs[1665]);
    assign layer1_outputs[11916] = layer0_outputs[10745];
    assign layer1_outputs[11917] = ~(layer0_outputs[9532]);
    assign layer1_outputs[11918] = ~((layer0_outputs[3312]) ^ (layer0_outputs[2089]));
    assign layer1_outputs[11919] = ~(layer0_outputs[9458]);
    assign layer1_outputs[11920] = ~(layer0_outputs[4720]) | (layer0_outputs[6074]);
    assign layer1_outputs[11921] = ~((layer0_outputs[9519]) & (layer0_outputs[1593]));
    assign layer1_outputs[11922] = (layer0_outputs[6177]) & ~(layer0_outputs[7367]);
    assign layer1_outputs[11923] = ~(layer0_outputs[12524]);
    assign layer1_outputs[11924] = ~(layer0_outputs[135]) | (layer0_outputs[8524]);
    assign layer1_outputs[11925] = layer0_outputs[2659];
    assign layer1_outputs[11926] = (layer0_outputs[6389]) ^ (layer0_outputs[3907]);
    assign layer1_outputs[11927] = ~(layer0_outputs[827]);
    assign layer1_outputs[11928] = ~(layer0_outputs[11754]);
    assign layer1_outputs[11929] = ~((layer0_outputs[11475]) ^ (layer0_outputs[5471]));
    assign layer1_outputs[11930] = ~(layer0_outputs[3354]) | (layer0_outputs[2134]);
    assign layer1_outputs[11931] = ~(layer0_outputs[10032]);
    assign layer1_outputs[11932] = (layer0_outputs[5849]) ^ (layer0_outputs[9138]);
    assign layer1_outputs[11933] = ~(layer0_outputs[5919]);
    assign layer1_outputs[11934] = (layer0_outputs[465]) & ~(layer0_outputs[7852]);
    assign layer1_outputs[11935] = ~(layer0_outputs[1759]) | (layer0_outputs[8604]);
    assign layer1_outputs[11936] = 1'b1;
    assign layer1_outputs[11937] = ~(layer0_outputs[4178]);
    assign layer1_outputs[11938] = ~((layer0_outputs[7631]) & (layer0_outputs[12763]));
    assign layer1_outputs[11939] = ~((layer0_outputs[12114]) & (layer0_outputs[11114]));
    assign layer1_outputs[11940] = ~(layer0_outputs[6195]);
    assign layer1_outputs[11941] = (layer0_outputs[1477]) & ~(layer0_outputs[8520]);
    assign layer1_outputs[11942] = ~((layer0_outputs[1919]) & (layer0_outputs[11470]));
    assign layer1_outputs[11943] = ~(layer0_outputs[393]);
    assign layer1_outputs[11944] = layer0_outputs[10912];
    assign layer1_outputs[11945] = (layer0_outputs[2269]) & ~(layer0_outputs[8009]);
    assign layer1_outputs[11946] = layer0_outputs[2510];
    assign layer1_outputs[11947] = (layer0_outputs[9587]) & ~(layer0_outputs[7493]);
    assign layer1_outputs[11948] = ~(layer0_outputs[3733]);
    assign layer1_outputs[11949] = layer0_outputs[8540];
    assign layer1_outputs[11950] = ~((layer0_outputs[9728]) | (layer0_outputs[3835]));
    assign layer1_outputs[11951] = (layer0_outputs[469]) & ~(layer0_outputs[1000]);
    assign layer1_outputs[11952] = (layer0_outputs[2449]) & ~(layer0_outputs[4935]);
    assign layer1_outputs[11953] = layer0_outputs[11610];
    assign layer1_outputs[11954] = (layer0_outputs[4732]) | (layer0_outputs[1047]);
    assign layer1_outputs[11955] = (layer0_outputs[11212]) & ~(layer0_outputs[4635]);
    assign layer1_outputs[11956] = (layer0_outputs[1393]) & ~(layer0_outputs[5331]);
    assign layer1_outputs[11957] = ~((layer0_outputs[301]) | (layer0_outputs[7464]));
    assign layer1_outputs[11958] = ~(layer0_outputs[1169]) | (layer0_outputs[5435]);
    assign layer1_outputs[11959] = ~(layer0_outputs[4251]) | (layer0_outputs[7656]);
    assign layer1_outputs[11960] = layer0_outputs[5558];
    assign layer1_outputs[11961] = 1'b0;
    assign layer1_outputs[11962] = layer0_outputs[8403];
    assign layer1_outputs[11963] = ~(layer0_outputs[11688]) | (layer0_outputs[6685]);
    assign layer1_outputs[11964] = layer0_outputs[9414];
    assign layer1_outputs[11965] = ~(layer0_outputs[3981]) | (layer0_outputs[4012]);
    assign layer1_outputs[11966] = (layer0_outputs[771]) & ~(layer0_outputs[8755]);
    assign layer1_outputs[11967] = layer0_outputs[11734];
    assign layer1_outputs[11968] = ~((layer0_outputs[735]) | (layer0_outputs[2895]));
    assign layer1_outputs[11969] = ~((layer0_outputs[1766]) | (layer0_outputs[5272]));
    assign layer1_outputs[11970] = ~(layer0_outputs[5672]);
    assign layer1_outputs[11971] = ~((layer0_outputs[3926]) & (layer0_outputs[6352]));
    assign layer1_outputs[11972] = (layer0_outputs[4677]) ^ (layer0_outputs[156]);
    assign layer1_outputs[11973] = (layer0_outputs[5229]) & ~(layer0_outputs[3570]);
    assign layer1_outputs[11974] = layer0_outputs[4504];
    assign layer1_outputs[11975] = ~((layer0_outputs[9077]) & (layer0_outputs[1565]));
    assign layer1_outputs[11976] = ~(layer0_outputs[12526]);
    assign layer1_outputs[11977] = layer0_outputs[1014];
    assign layer1_outputs[11978] = ~(layer0_outputs[6277]);
    assign layer1_outputs[11979] = layer0_outputs[7189];
    assign layer1_outputs[11980] = layer0_outputs[1510];
    assign layer1_outputs[11981] = layer0_outputs[12633];
    assign layer1_outputs[11982] = ~((layer0_outputs[3730]) | (layer0_outputs[5874]));
    assign layer1_outputs[11983] = (layer0_outputs[3730]) | (layer0_outputs[9575]);
    assign layer1_outputs[11984] = (layer0_outputs[3497]) | (layer0_outputs[3993]);
    assign layer1_outputs[11985] = (layer0_outputs[1735]) & ~(layer0_outputs[4708]);
    assign layer1_outputs[11986] = (layer0_outputs[2093]) & ~(layer0_outputs[10642]);
    assign layer1_outputs[11987] = (layer0_outputs[3650]) & ~(layer0_outputs[10826]);
    assign layer1_outputs[11988] = ~((layer0_outputs[1922]) | (layer0_outputs[7627]));
    assign layer1_outputs[11989] = layer0_outputs[9752];
    assign layer1_outputs[11990] = ~(layer0_outputs[9818]) | (layer0_outputs[2679]);
    assign layer1_outputs[11991] = ~(layer0_outputs[11615]);
    assign layer1_outputs[11992] = ~(layer0_outputs[10473]) | (layer0_outputs[10344]);
    assign layer1_outputs[11993] = ~(layer0_outputs[279]);
    assign layer1_outputs[11994] = ~(layer0_outputs[5403]);
    assign layer1_outputs[11995] = (layer0_outputs[11718]) & ~(layer0_outputs[9119]);
    assign layer1_outputs[11996] = (layer0_outputs[5450]) & (layer0_outputs[1613]);
    assign layer1_outputs[11997] = (layer0_outputs[11846]) & (layer0_outputs[10661]);
    assign layer1_outputs[11998] = (layer0_outputs[9588]) & ~(layer0_outputs[4885]);
    assign layer1_outputs[11999] = layer0_outputs[6967];
    assign layer1_outputs[12000] = (layer0_outputs[7416]) & (layer0_outputs[719]);
    assign layer1_outputs[12001] = (layer0_outputs[12292]) & (layer0_outputs[5394]);
    assign layer1_outputs[12002] = ~(layer0_outputs[12446]);
    assign layer1_outputs[12003] = (layer0_outputs[8556]) | (layer0_outputs[12439]);
    assign layer1_outputs[12004] = (layer0_outputs[12514]) & ~(layer0_outputs[5513]);
    assign layer1_outputs[12005] = ~((layer0_outputs[5507]) & (layer0_outputs[720]));
    assign layer1_outputs[12006] = (layer0_outputs[12607]) ^ (layer0_outputs[9853]);
    assign layer1_outputs[12007] = 1'b1;
    assign layer1_outputs[12008] = ~(layer0_outputs[12477]);
    assign layer1_outputs[12009] = (layer0_outputs[10537]) & (layer0_outputs[806]);
    assign layer1_outputs[12010] = (layer0_outputs[6281]) ^ (layer0_outputs[4917]);
    assign layer1_outputs[12011] = ~(layer0_outputs[11240]) | (layer0_outputs[9738]);
    assign layer1_outputs[12012] = ~((layer0_outputs[11521]) & (layer0_outputs[3027]));
    assign layer1_outputs[12013] = ~(layer0_outputs[10485]);
    assign layer1_outputs[12014] = ~(layer0_outputs[6348]);
    assign layer1_outputs[12015] = ~((layer0_outputs[8481]) | (layer0_outputs[7450]));
    assign layer1_outputs[12016] = (layer0_outputs[4950]) | (layer0_outputs[7109]);
    assign layer1_outputs[12017] = (layer0_outputs[9661]) & ~(layer0_outputs[11973]);
    assign layer1_outputs[12018] = ~(layer0_outputs[6339]);
    assign layer1_outputs[12019] = ~(layer0_outputs[11759]) | (layer0_outputs[10709]);
    assign layer1_outputs[12020] = ~(layer0_outputs[3545]) | (layer0_outputs[2039]);
    assign layer1_outputs[12021] = ~((layer0_outputs[536]) & (layer0_outputs[4120]));
    assign layer1_outputs[12022] = 1'b1;
    assign layer1_outputs[12023] = layer0_outputs[1588];
    assign layer1_outputs[12024] = ~(layer0_outputs[12395]);
    assign layer1_outputs[12025] = ~(layer0_outputs[4451]);
    assign layer1_outputs[12026] = ~(layer0_outputs[7332]);
    assign layer1_outputs[12027] = ~(layer0_outputs[10733]);
    assign layer1_outputs[12028] = 1'b0;
    assign layer1_outputs[12029] = layer0_outputs[12685];
    assign layer1_outputs[12030] = (layer0_outputs[1354]) & ~(layer0_outputs[12217]);
    assign layer1_outputs[12031] = ~(layer0_outputs[11251]);
    assign layer1_outputs[12032] = (layer0_outputs[1545]) & ~(layer0_outputs[6586]);
    assign layer1_outputs[12033] = (layer0_outputs[9495]) & ~(layer0_outputs[9229]);
    assign layer1_outputs[12034] = layer0_outputs[9285];
    assign layer1_outputs[12035] = layer0_outputs[12565];
    assign layer1_outputs[12036] = layer0_outputs[2580];
    assign layer1_outputs[12037] = (layer0_outputs[5334]) & ~(layer0_outputs[6802]);
    assign layer1_outputs[12038] = (layer0_outputs[1616]) & ~(layer0_outputs[7371]);
    assign layer1_outputs[12039] = (layer0_outputs[7611]) & (layer0_outputs[636]);
    assign layer1_outputs[12040] = (layer0_outputs[10133]) & ~(layer0_outputs[10856]);
    assign layer1_outputs[12041] = layer0_outputs[3918];
    assign layer1_outputs[12042] = ~(layer0_outputs[881]);
    assign layer1_outputs[12043] = layer0_outputs[1135];
    assign layer1_outputs[12044] = ~(layer0_outputs[3406]) | (layer0_outputs[9831]);
    assign layer1_outputs[12045] = (layer0_outputs[517]) & ~(layer0_outputs[5573]);
    assign layer1_outputs[12046] = (layer0_outputs[10388]) | (layer0_outputs[8936]);
    assign layer1_outputs[12047] = (layer0_outputs[3369]) & (layer0_outputs[11211]);
    assign layer1_outputs[12048] = ~((layer0_outputs[7043]) & (layer0_outputs[9683]));
    assign layer1_outputs[12049] = ~(layer0_outputs[8750]) | (layer0_outputs[2501]);
    assign layer1_outputs[12050] = layer0_outputs[1094];
    assign layer1_outputs[12051] = layer0_outputs[1372];
    assign layer1_outputs[12052] = ~(layer0_outputs[4804]);
    assign layer1_outputs[12053] = ~((layer0_outputs[391]) | (layer0_outputs[5920]));
    assign layer1_outputs[12054] = layer0_outputs[11789];
    assign layer1_outputs[12055] = ~(layer0_outputs[704]);
    assign layer1_outputs[12056] = ~(layer0_outputs[11988]);
    assign layer1_outputs[12057] = ~(layer0_outputs[12773]);
    assign layer1_outputs[12058] = ~(layer0_outputs[8818]);
    assign layer1_outputs[12059] = ~((layer0_outputs[2986]) & (layer0_outputs[509]));
    assign layer1_outputs[12060] = ~((layer0_outputs[11263]) ^ (layer0_outputs[5238]));
    assign layer1_outputs[12061] = layer0_outputs[10996];
    assign layer1_outputs[12062] = ~(layer0_outputs[3169]) | (layer0_outputs[11045]);
    assign layer1_outputs[12063] = ~(layer0_outputs[2647]);
    assign layer1_outputs[12064] = ~((layer0_outputs[8945]) & (layer0_outputs[7563]));
    assign layer1_outputs[12065] = (layer0_outputs[2502]) | (layer0_outputs[6931]);
    assign layer1_outputs[12066] = (layer0_outputs[9710]) | (layer0_outputs[1538]);
    assign layer1_outputs[12067] = (layer0_outputs[5580]) & ~(layer0_outputs[10049]);
    assign layer1_outputs[12068] = ~((layer0_outputs[9814]) ^ (layer0_outputs[11520]));
    assign layer1_outputs[12069] = (layer0_outputs[25]) | (layer0_outputs[2917]);
    assign layer1_outputs[12070] = (layer0_outputs[4186]) ^ (layer0_outputs[5141]);
    assign layer1_outputs[12071] = ~(layer0_outputs[12140]);
    assign layer1_outputs[12072] = (layer0_outputs[4329]) & ~(layer0_outputs[8130]);
    assign layer1_outputs[12073] = (layer0_outputs[6411]) | (layer0_outputs[10790]);
    assign layer1_outputs[12074] = (layer0_outputs[11782]) | (layer0_outputs[1470]);
    assign layer1_outputs[12075] = layer0_outputs[4398];
    assign layer1_outputs[12076] = ~(layer0_outputs[4516]);
    assign layer1_outputs[12077] = (layer0_outputs[362]) | (layer0_outputs[323]);
    assign layer1_outputs[12078] = (layer0_outputs[6734]) & (layer0_outputs[2941]);
    assign layer1_outputs[12079] = (layer0_outputs[6128]) ^ (layer0_outputs[1159]);
    assign layer1_outputs[12080] = (layer0_outputs[3999]) ^ (layer0_outputs[1651]);
    assign layer1_outputs[12081] = ~(layer0_outputs[8201]);
    assign layer1_outputs[12082] = layer0_outputs[5940];
    assign layer1_outputs[12083] = 1'b1;
    assign layer1_outputs[12084] = layer0_outputs[1869];
    assign layer1_outputs[12085] = ~((layer0_outputs[11346]) | (layer0_outputs[7814]));
    assign layer1_outputs[12086] = layer0_outputs[11451];
    assign layer1_outputs[12087] = ~((layer0_outputs[12047]) ^ (layer0_outputs[6101]));
    assign layer1_outputs[12088] = ~((layer0_outputs[314]) | (layer0_outputs[2101]));
    assign layer1_outputs[12089] = ~(layer0_outputs[11019]) | (layer0_outputs[2346]);
    assign layer1_outputs[12090] = (layer0_outputs[8937]) & ~(layer0_outputs[7731]);
    assign layer1_outputs[12091] = 1'b1;
    assign layer1_outputs[12092] = (layer0_outputs[9566]) & ~(layer0_outputs[760]);
    assign layer1_outputs[12093] = (layer0_outputs[11489]) & ~(layer0_outputs[10110]);
    assign layer1_outputs[12094] = (layer0_outputs[5729]) & ~(layer0_outputs[5715]);
    assign layer1_outputs[12095] = ~((layer0_outputs[6630]) | (layer0_outputs[3224]));
    assign layer1_outputs[12096] = layer0_outputs[8868];
    assign layer1_outputs[12097] = ~((layer0_outputs[2359]) | (layer0_outputs[7684]));
    assign layer1_outputs[12098] = ~(layer0_outputs[7329]);
    assign layer1_outputs[12099] = layer0_outputs[11173];
    assign layer1_outputs[12100] = (layer0_outputs[482]) | (layer0_outputs[9063]);
    assign layer1_outputs[12101] = layer0_outputs[7078];
    assign layer1_outputs[12102] = layer0_outputs[7788];
    assign layer1_outputs[12103] = layer0_outputs[10734];
    assign layer1_outputs[12104] = (layer0_outputs[1070]) | (layer0_outputs[5421]);
    assign layer1_outputs[12105] = layer0_outputs[7662];
    assign layer1_outputs[12106] = (layer0_outputs[1533]) & ~(layer0_outputs[5627]);
    assign layer1_outputs[12107] = layer0_outputs[5217];
    assign layer1_outputs[12108] = (layer0_outputs[11350]) ^ (layer0_outputs[10293]);
    assign layer1_outputs[12109] = layer0_outputs[6880];
    assign layer1_outputs[12110] = ~(layer0_outputs[1754]) | (layer0_outputs[7974]);
    assign layer1_outputs[12111] = (layer0_outputs[8533]) ^ (layer0_outputs[9430]);
    assign layer1_outputs[12112] = 1'b1;
    assign layer1_outputs[12113] = ~(layer0_outputs[8188]);
    assign layer1_outputs[12114] = (layer0_outputs[5038]) | (layer0_outputs[11015]);
    assign layer1_outputs[12115] = ~(layer0_outputs[2034]);
    assign layer1_outputs[12116] = layer0_outputs[3241];
    assign layer1_outputs[12117] = (layer0_outputs[5477]) & (layer0_outputs[5441]);
    assign layer1_outputs[12118] = ~(layer0_outputs[8962]);
    assign layer1_outputs[12119] = ~(layer0_outputs[4061]) | (layer0_outputs[4932]);
    assign layer1_outputs[12120] = ~(layer0_outputs[12389]);
    assign layer1_outputs[12121] = ~(layer0_outputs[10412]);
    assign layer1_outputs[12122] = layer0_outputs[4129];
    assign layer1_outputs[12123] = ~(layer0_outputs[4873]);
    assign layer1_outputs[12124] = ~((layer0_outputs[12673]) ^ (layer0_outputs[11581]));
    assign layer1_outputs[12125] = ~(layer0_outputs[8352]);
    assign layer1_outputs[12126] = (layer0_outputs[5184]) & (layer0_outputs[10647]);
    assign layer1_outputs[12127] = (layer0_outputs[7066]) & ~(layer0_outputs[11492]);
    assign layer1_outputs[12128] = (layer0_outputs[4371]) | (layer0_outputs[5987]);
    assign layer1_outputs[12129] = layer0_outputs[2755];
    assign layer1_outputs[12130] = (layer0_outputs[1780]) | (layer0_outputs[4889]);
    assign layer1_outputs[12131] = (layer0_outputs[6759]) & (layer0_outputs[8611]);
    assign layer1_outputs[12132] = (layer0_outputs[8063]) ^ (layer0_outputs[11838]);
    assign layer1_outputs[12133] = layer0_outputs[1931];
    assign layer1_outputs[12134] = ~(layer0_outputs[12219]) | (layer0_outputs[7934]);
    assign layer1_outputs[12135] = (layer0_outputs[3221]) ^ (layer0_outputs[2631]);
    assign layer1_outputs[12136] = ~((layer0_outputs[2351]) & (layer0_outputs[6534]));
    assign layer1_outputs[12137] = ~(layer0_outputs[11650]);
    assign layer1_outputs[12138] = ~((layer0_outputs[11953]) | (layer0_outputs[4996]));
    assign layer1_outputs[12139] = layer0_outputs[1318];
    assign layer1_outputs[12140] = ~(layer0_outputs[12659]);
    assign layer1_outputs[12141] = ~(layer0_outputs[9022]);
    assign layer1_outputs[12142] = ~(layer0_outputs[4153]);
    assign layer1_outputs[12143] = ~(layer0_outputs[8257]) | (layer0_outputs[4871]);
    assign layer1_outputs[12144] = ~((layer0_outputs[3541]) ^ (layer0_outputs[10110]));
    assign layer1_outputs[12145] = layer0_outputs[783];
    assign layer1_outputs[12146] = ~((layer0_outputs[11885]) & (layer0_outputs[10688]));
    assign layer1_outputs[12147] = (layer0_outputs[1330]) ^ (layer0_outputs[11964]);
    assign layer1_outputs[12148] = (layer0_outputs[5492]) & ~(layer0_outputs[6865]);
    assign layer1_outputs[12149] = layer0_outputs[7921];
    assign layer1_outputs[12150] = (layer0_outputs[12163]) ^ (layer0_outputs[10751]);
    assign layer1_outputs[12151] = ~(layer0_outputs[7182]) | (layer0_outputs[961]);
    assign layer1_outputs[12152] = layer0_outputs[1969];
    assign layer1_outputs[12153] = (layer0_outputs[6929]) & ~(layer0_outputs[12376]);
    assign layer1_outputs[12154] = ~((layer0_outputs[10378]) & (layer0_outputs[9893]));
    assign layer1_outputs[12155] = ~((layer0_outputs[10397]) & (layer0_outputs[3753]));
    assign layer1_outputs[12156] = ~(layer0_outputs[4016]);
    assign layer1_outputs[12157] = ~(layer0_outputs[12580]);
    assign layer1_outputs[12158] = (layer0_outputs[12087]) ^ (layer0_outputs[11010]);
    assign layer1_outputs[12159] = ~(layer0_outputs[7904]);
    assign layer1_outputs[12160] = layer0_outputs[2768];
    assign layer1_outputs[12161] = layer0_outputs[1621];
    assign layer1_outputs[12162] = ~((layer0_outputs[5065]) | (layer0_outputs[1667]));
    assign layer1_outputs[12163] = (layer0_outputs[8684]) | (layer0_outputs[9176]);
    assign layer1_outputs[12164] = ~(layer0_outputs[8219]);
    assign layer1_outputs[12165] = (layer0_outputs[6604]) & (layer0_outputs[10609]);
    assign layer1_outputs[12166] = ~(layer0_outputs[11725]);
    assign layer1_outputs[12167] = layer0_outputs[8778];
    assign layer1_outputs[12168] = layer0_outputs[3998];
    assign layer1_outputs[12169] = ~(layer0_outputs[8115]);
    assign layer1_outputs[12170] = (layer0_outputs[2792]) ^ (layer0_outputs[8306]);
    assign layer1_outputs[12171] = 1'b0;
    assign layer1_outputs[12172] = (layer0_outputs[3820]) ^ (layer0_outputs[7602]);
    assign layer1_outputs[12173] = (layer0_outputs[7224]) & ~(layer0_outputs[11282]);
    assign layer1_outputs[12174] = ~((layer0_outputs[10019]) & (layer0_outputs[1569]));
    assign layer1_outputs[12175] = ~((layer0_outputs[8631]) | (layer0_outputs[3533]));
    assign layer1_outputs[12176] = (layer0_outputs[12669]) ^ (layer0_outputs[2737]);
    assign layer1_outputs[12177] = ~(layer0_outputs[5556]) | (layer0_outputs[2644]);
    assign layer1_outputs[12178] = ~(layer0_outputs[7031]);
    assign layer1_outputs[12179] = ~(layer0_outputs[5561]);
    assign layer1_outputs[12180] = layer0_outputs[2884];
    assign layer1_outputs[12181] = ~((layer0_outputs[11751]) & (layer0_outputs[12398]));
    assign layer1_outputs[12182] = layer0_outputs[303];
    assign layer1_outputs[12183] = ~((layer0_outputs[2961]) & (layer0_outputs[1398]));
    assign layer1_outputs[12184] = layer0_outputs[11196];
    assign layer1_outputs[12185] = (layer0_outputs[608]) & (layer0_outputs[4291]);
    assign layer1_outputs[12186] = ~(layer0_outputs[7684]);
    assign layer1_outputs[12187] = ~(layer0_outputs[819]) | (layer0_outputs[8644]);
    assign layer1_outputs[12188] = layer0_outputs[5309];
    assign layer1_outputs[12189] = layer0_outputs[2392];
    assign layer1_outputs[12190] = (layer0_outputs[8435]) & (layer0_outputs[3338]);
    assign layer1_outputs[12191] = ~(layer0_outputs[4452]) | (layer0_outputs[728]);
    assign layer1_outputs[12192] = layer0_outputs[11707];
    assign layer1_outputs[12193] = ~((layer0_outputs[1875]) ^ (layer0_outputs[8963]));
    assign layer1_outputs[12194] = (layer0_outputs[7352]) & (layer0_outputs[4259]);
    assign layer1_outputs[12195] = ~(layer0_outputs[9419]);
    assign layer1_outputs[12196] = layer0_outputs[2637];
    assign layer1_outputs[12197] = ~((layer0_outputs[5860]) ^ (layer0_outputs[8558]));
    assign layer1_outputs[12198] = (layer0_outputs[2471]) & (layer0_outputs[8858]);
    assign layer1_outputs[12199] = (layer0_outputs[7883]) & ~(layer0_outputs[7596]);
    assign layer1_outputs[12200] = (layer0_outputs[10599]) ^ (layer0_outputs[5139]);
    assign layer1_outputs[12201] = ~((layer0_outputs[7176]) & (layer0_outputs[3106]));
    assign layer1_outputs[12202] = layer0_outputs[4534];
    assign layer1_outputs[12203] = layer0_outputs[10160];
    assign layer1_outputs[12204] = (layer0_outputs[9929]) | (layer0_outputs[4643]);
    assign layer1_outputs[12205] = ~(layer0_outputs[4901]);
    assign layer1_outputs[12206] = ~(layer0_outputs[10999]);
    assign layer1_outputs[12207] = ~(layer0_outputs[9527]);
    assign layer1_outputs[12208] = (layer0_outputs[8319]) & (layer0_outputs[1029]);
    assign layer1_outputs[12209] = ~((layer0_outputs[6893]) | (layer0_outputs[5629]));
    assign layer1_outputs[12210] = ~(layer0_outputs[82]);
    assign layer1_outputs[12211] = ~((layer0_outputs[10798]) | (layer0_outputs[7153]));
    assign layer1_outputs[12212] = ~(layer0_outputs[3066]);
    assign layer1_outputs[12213] = ~(layer0_outputs[421]) | (layer0_outputs[8742]);
    assign layer1_outputs[12214] = ~((layer0_outputs[4896]) | (layer0_outputs[5230]));
    assign layer1_outputs[12215] = ~(layer0_outputs[3697]);
    assign layer1_outputs[12216] = ~((layer0_outputs[4156]) | (layer0_outputs[9471]));
    assign layer1_outputs[12217] = (layer0_outputs[11270]) & ~(layer0_outputs[11965]);
    assign layer1_outputs[12218] = layer0_outputs[3569];
    assign layer1_outputs[12219] = ~(layer0_outputs[5675]) | (layer0_outputs[9019]);
    assign layer1_outputs[12220] = ~(layer0_outputs[1888]);
    assign layer1_outputs[12221] = (layer0_outputs[12494]) | (layer0_outputs[4291]);
    assign layer1_outputs[12222] = ~(layer0_outputs[3473]);
    assign layer1_outputs[12223] = ~(layer0_outputs[8714]) | (layer0_outputs[1461]);
    assign layer1_outputs[12224] = ~(layer0_outputs[6206]);
    assign layer1_outputs[12225] = ~(layer0_outputs[320]) | (layer0_outputs[8015]);
    assign layer1_outputs[12226] = ~(layer0_outputs[12243]);
    assign layer1_outputs[12227] = ~(layer0_outputs[2821]) | (layer0_outputs[8316]);
    assign layer1_outputs[12228] = ~(layer0_outputs[12145]) | (layer0_outputs[9654]);
    assign layer1_outputs[12229] = (layer0_outputs[571]) | (layer0_outputs[5286]);
    assign layer1_outputs[12230] = ~(layer0_outputs[2756]);
    assign layer1_outputs[12231] = ~(layer0_outputs[8040]) | (layer0_outputs[2385]);
    assign layer1_outputs[12232] = (layer0_outputs[4908]) | (layer0_outputs[1843]);
    assign layer1_outputs[12233] = ~(layer0_outputs[12093]) | (layer0_outputs[4629]);
    assign layer1_outputs[12234] = layer0_outputs[8300];
    assign layer1_outputs[12235] = ~((layer0_outputs[4060]) | (layer0_outputs[6003]));
    assign layer1_outputs[12236] = (layer0_outputs[11424]) ^ (layer0_outputs[7495]);
    assign layer1_outputs[12237] = (layer0_outputs[8605]) ^ (layer0_outputs[7889]);
    assign layer1_outputs[12238] = layer0_outputs[2936];
    assign layer1_outputs[12239] = ~((layer0_outputs[4461]) & (layer0_outputs[2133]));
    assign layer1_outputs[12240] = (layer0_outputs[3446]) & (layer0_outputs[476]);
    assign layer1_outputs[12241] = ~(layer0_outputs[12453]);
    assign layer1_outputs[12242] = (layer0_outputs[4868]) & (layer0_outputs[8754]);
    assign layer1_outputs[12243] = ~(layer0_outputs[11666]) | (layer0_outputs[4487]);
    assign layer1_outputs[12244] = ~(layer0_outputs[9240]) | (layer0_outputs[12199]);
    assign layer1_outputs[12245] = (layer0_outputs[5994]) | (layer0_outputs[6642]);
    assign layer1_outputs[12246] = (layer0_outputs[6657]) & (layer0_outputs[4402]);
    assign layer1_outputs[12247] = ~((layer0_outputs[11878]) ^ (layer0_outputs[7562]));
    assign layer1_outputs[12248] = ~(layer0_outputs[11172]);
    assign layer1_outputs[12249] = (layer0_outputs[386]) & (layer0_outputs[10141]);
    assign layer1_outputs[12250] = (layer0_outputs[9743]) & (layer0_outputs[2258]);
    assign layer1_outputs[12251] = layer0_outputs[9744];
    assign layer1_outputs[12252] = ~(layer0_outputs[6348]);
    assign layer1_outputs[12253] = ~(layer0_outputs[5625]);
    assign layer1_outputs[12254] = (layer0_outputs[10837]) ^ (layer0_outputs[4429]);
    assign layer1_outputs[12255] = ~(layer0_outputs[3792]);
    assign layer1_outputs[12256] = 1'b0;
    assign layer1_outputs[12257] = (layer0_outputs[9167]) & (layer0_outputs[7093]);
    assign layer1_outputs[12258] = (layer0_outputs[9810]) & (layer0_outputs[10214]);
    assign layer1_outputs[12259] = ~(layer0_outputs[6230]);
    assign layer1_outputs[12260] = ~((layer0_outputs[377]) ^ (layer0_outputs[9899]));
    assign layer1_outputs[12261] = ~(layer0_outputs[7386]);
    assign layer1_outputs[12262] = ~(layer0_outputs[1466]);
    assign layer1_outputs[12263] = layer0_outputs[2088];
    assign layer1_outputs[12264] = (layer0_outputs[3870]) & ~(layer0_outputs[7573]);
    assign layer1_outputs[12265] = ~(layer0_outputs[8817]);
    assign layer1_outputs[12266] = (layer0_outputs[4180]) ^ (layer0_outputs[2667]);
    assign layer1_outputs[12267] = ~(layer0_outputs[1134]) | (layer0_outputs[8150]);
    assign layer1_outputs[12268] = (layer0_outputs[11066]) | (layer0_outputs[3278]);
    assign layer1_outputs[12269] = (layer0_outputs[11023]) | (layer0_outputs[7047]);
    assign layer1_outputs[12270] = ~(layer0_outputs[8744]);
    assign layer1_outputs[12271] = ~(layer0_outputs[1636]) | (layer0_outputs[4581]);
    assign layer1_outputs[12272] = layer0_outputs[8114];
    assign layer1_outputs[12273] = (layer0_outputs[8813]) | (layer0_outputs[7599]);
    assign layer1_outputs[12274] = ~((layer0_outputs[1360]) ^ (layer0_outputs[3390]));
    assign layer1_outputs[12275] = (layer0_outputs[1860]) ^ (layer0_outputs[6280]);
    assign layer1_outputs[12276] = (layer0_outputs[10000]) | (layer0_outputs[9068]);
    assign layer1_outputs[12277] = layer0_outputs[3716];
    assign layer1_outputs[12278] = ~(layer0_outputs[1946]);
    assign layer1_outputs[12279] = (layer0_outputs[11282]) & ~(layer0_outputs[6635]);
    assign layer1_outputs[12280] = ~((layer0_outputs[12546]) ^ (layer0_outputs[305]));
    assign layer1_outputs[12281] = layer0_outputs[4110];
    assign layer1_outputs[12282] = layer0_outputs[149];
    assign layer1_outputs[12283] = layer0_outputs[12553];
    assign layer1_outputs[12284] = ~(layer0_outputs[8728]);
    assign layer1_outputs[12285] = layer0_outputs[2201];
    assign layer1_outputs[12286] = (layer0_outputs[10652]) | (layer0_outputs[11567]);
    assign layer1_outputs[12287] = ~(layer0_outputs[3896]);
    assign layer1_outputs[12288] = (layer0_outputs[10078]) | (layer0_outputs[3267]);
    assign layer1_outputs[12289] = ~(layer0_outputs[4773]);
    assign layer1_outputs[12290] = layer0_outputs[7152];
    assign layer1_outputs[12291] = layer0_outputs[629];
    assign layer1_outputs[12292] = ~(layer0_outputs[501]);
    assign layer1_outputs[12293] = ~(layer0_outputs[12600]) | (layer0_outputs[674]);
    assign layer1_outputs[12294] = layer0_outputs[2914];
    assign layer1_outputs[12295] = (layer0_outputs[7479]) | (layer0_outputs[5093]);
    assign layer1_outputs[12296] = ~((layer0_outputs[122]) & (layer0_outputs[4564]));
    assign layer1_outputs[12297] = ~(layer0_outputs[4263]);
    assign layer1_outputs[12298] = 1'b0;
    assign layer1_outputs[12299] = 1'b1;
    assign layer1_outputs[12300] = ~((layer0_outputs[9725]) & (layer0_outputs[436]));
    assign layer1_outputs[12301] = layer0_outputs[8537];
    assign layer1_outputs[12302] = ~(layer0_outputs[9605]) | (layer0_outputs[10710]);
    assign layer1_outputs[12303] = ~(layer0_outputs[8134]);
    assign layer1_outputs[12304] = ~((layer0_outputs[2335]) ^ (layer0_outputs[11900]));
    assign layer1_outputs[12305] = ~(layer0_outputs[7172]);
    assign layer1_outputs[12306] = layer0_outputs[7348];
    assign layer1_outputs[12307] = ~(layer0_outputs[4936]);
    assign layer1_outputs[12308] = layer0_outputs[4872];
    assign layer1_outputs[12309] = ~(layer0_outputs[3116]);
    assign layer1_outputs[12310] = layer0_outputs[5592];
    assign layer1_outputs[12311] = ~(layer0_outputs[4915]);
    assign layer1_outputs[12312] = (layer0_outputs[3906]) ^ (layer0_outputs[11199]);
    assign layer1_outputs[12313] = ~(layer0_outputs[8852]) | (layer0_outputs[5918]);
    assign layer1_outputs[12314] = (layer0_outputs[1398]) ^ (layer0_outputs[1214]);
    assign layer1_outputs[12315] = ~((layer0_outputs[12143]) & (layer0_outputs[5730]));
    assign layer1_outputs[12316] = layer0_outputs[1727];
    assign layer1_outputs[12317] = ~(layer0_outputs[5454]) | (layer0_outputs[4318]);
    assign layer1_outputs[12318] = ~(layer0_outputs[8961]);
    assign layer1_outputs[12319] = layer0_outputs[1654];
    assign layer1_outputs[12320] = ~(layer0_outputs[6066]);
    assign layer1_outputs[12321] = (layer0_outputs[9638]) & ~(layer0_outputs[7272]);
    assign layer1_outputs[12322] = (layer0_outputs[6856]) | (layer0_outputs[2906]);
    assign layer1_outputs[12323] = 1'b1;
    assign layer1_outputs[12324] = layer0_outputs[3048];
    assign layer1_outputs[12325] = layer0_outputs[6565];
    assign layer1_outputs[12326] = ~(layer0_outputs[4021]);
    assign layer1_outputs[12327] = (layer0_outputs[7979]) & ~(layer0_outputs[3923]);
    assign layer1_outputs[12328] = ~(layer0_outputs[3561]) | (layer0_outputs[11329]);
    assign layer1_outputs[12329] = ~(layer0_outputs[2264]) | (layer0_outputs[6820]);
    assign layer1_outputs[12330] = (layer0_outputs[3986]) & (layer0_outputs[4890]);
    assign layer1_outputs[12331] = ~(layer0_outputs[8022]);
    assign layer1_outputs[12332] = (layer0_outputs[12582]) & (layer0_outputs[9465]);
    assign layer1_outputs[12333] = ~((layer0_outputs[6488]) ^ (layer0_outputs[7435]));
    assign layer1_outputs[12334] = (layer0_outputs[12510]) | (layer0_outputs[10827]);
    assign layer1_outputs[12335] = (layer0_outputs[273]) | (layer0_outputs[4455]);
    assign layer1_outputs[12336] = (layer0_outputs[660]) & ~(layer0_outputs[10859]);
    assign layer1_outputs[12337] = ~((layer0_outputs[7782]) & (layer0_outputs[6318]));
    assign layer1_outputs[12338] = layer0_outputs[248];
    assign layer1_outputs[12339] = ~(layer0_outputs[3255]) | (layer0_outputs[9886]);
    assign layer1_outputs[12340] = layer0_outputs[6649];
    assign layer1_outputs[12341] = (layer0_outputs[2507]) & ~(layer0_outputs[9878]);
    assign layer1_outputs[12342] = (layer0_outputs[10119]) | (layer0_outputs[9747]);
    assign layer1_outputs[12343] = ~(layer0_outputs[8848]);
    assign layer1_outputs[12344] = ~(layer0_outputs[2097]) | (layer0_outputs[5505]);
    assign layer1_outputs[12345] = ~((layer0_outputs[12799]) & (layer0_outputs[4044]));
    assign layer1_outputs[12346] = (layer0_outputs[7658]) & ~(layer0_outputs[5326]);
    assign layer1_outputs[12347] = ~(layer0_outputs[1072]);
    assign layer1_outputs[12348] = (layer0_outputs[7910]) & ~(layer0_outputs[6115]);
    assign layer1_outputs[12349] = ~(layer0_outputs[12080]);
    assign layer1_outputs[12350] = ~((layer0_outputs[6076]) | (layer0_outputs[1990]));
    assign layer1_outputs[12351] = ~(layer0_outputs[1314]) | (layer0_outputs[10888]);
    assign layer1_outputs[12352] = ~((layer0_outputs[9781]) | (layer0_outputs[10524]));
    assign layer1_outputs[12353] = (layer0_outputs[901]) | (layer0_outputs[10175]);
    assign layer1_outputs[12354] = ~(layer0_outputs[6954]) | (layer0_outputs[7864]);
    assign layer1_outputs[12355] = ~(layer0_outputs[1304]) | (layer0_outputs[12343]);
    assign layer1_outputs[12356] = ~(layer0_outputs[4672]);
    assign layer1_outputs[12357] = layer0_outputs[5547];
    assign layer1_outputs[12358] = ~(layer0_outputs[11358]);
    assign layer1_outputs[12359] = layer0_outputs[3934];
    assign layer1_outputs[12360] = ~(layer0_outputs[4466]);
    assign layer1_outputs[12361] = ~((layer0_outputs[12759]) | (layer0_outputs[9066]));
    assign layer1_outputs[12362] = (layer0_outputs[10515]) & ~(layer0_outputs[863]);
    assign layer1_outputs[12363] = ~(layer0_outputs[5855]);
    assign layer1_outputs[12364] = ~(layer0_outputs[3759]) | (layer0_outputs[9816]);
    assign layer1_outputs[12365] = ~(layer0_outputs[9751]);
    assign layer1_outputs[12366] = ~((layer0_outputs[10125]) ^ (layer0_outputs[4981]));
    assign layer1_outputs[12367] = ~(layer0_outputs[10335]) | (layer0_outputs[12188]);
    assign layer1_outputs[12368] = ~(layer0_outputs[6616]) | (layer0_outputs[1342]);
    assign layer1_outputs[12369] = layer0_outputs[5521];
    assign layer1_outputs[12370] = layer0_outputs[7313];
    assign layer1_outputs[12371] = ~(layer0_outputs[12053]);
    assign layer1_outputs[12372] = (layer0_outputs[12336]) | (layer0_outputs[402]);
    assign layer1_outputs[12373] = ~((layer0_outputs[5913]) ^ (layer0_outputs[3109]));
    assign layer1_outputs[12374] = ~(layer0_outputs[2244]);
    assign layer1_outputs[12375] = ~(layer0_outputs[11838]);
    assign layer1_outputs[12376] = ~(layer0_outputs[5042]);
    assign layer1_outputs[12377] = ~(layer0_outputs[8023]);
    assign layer1_outputs[12378] = ~(layer0_outputs[404]);
    assign layer1_outputs[12379] = ~(layer0_outputs[10502]);
    assign layer1_outputs[12380] = layer0_outputs[9911];
    assign layer1_outputs[12381] = ~((layer0_outputs[12387]) ^ (layer0_outputs[12552]));
    assign layer1_outputs[12382] = (layer0_outputs[6480]) ^ (layer0_outputs[5368]);
    assign layer1_outputs[12383] = ~(layer0_outputs[730]) | (layer0_outputs[1947]);
    assign layer1_outputs[12384] = (layer0_outputs[1442]) & (layer0_outputs[2339]);
    assign layer1_outputs[12385] = ~(layer0_outputs[7425]);
    assign layer1_outputs[12386] = layer0_outputs[5848];
    assign layer1_outputs[12387] = ~(layer0_outputs[6218]) | (layer0_outputs[922]);
    assign layer1_outputs[12388] = 1'b0;
    assign layer1_outputs[12389] = ~((layer0_outputs[6178]) & (layer0_outputs[6324]));
    assign layer1_outputs[12390] = ~(layer0_outputs[11040]) | (layer0_outputs[2524]);
    assign layer1_outputs[12391] = ~(layer0_outputs[10148]);
    assign layer1_outputs[12392] = ~(layer0_outputs[5040]);
    assign layer1_outputs[12393] = layer0_outputs[5357];
    assign layer1_outputs[12394] = (layer0_outputs[1702]) | (layer0_outputs[9661]);
    assign layer1_outputs[12395] = layer0_outputs[5515];
    assign layer1_outputs[12396] = ~(layer0_outputs[6815]);
    assign layer1_outputs[12397] = ~(layer0_outputs[8478]);
    assign layer1_outputs[12398] = layer0_outputs[6431];
    assign layer1_outputs[12399] = ~((layer0_outputs[3310]) | (layer0_outputs[1548]));
    assign layer1_outputs[12400] = layer0_outputs[10327];
    assign layer1_outputs[12401] = (layer0_outputs[10608]) | (layer0_outputs[6599]);
    assign layer1_outputs[12402] = ~(layer0_outputs[5216]) | (layer0_outputs[11799]);
    assign layer1_outputs[12403] = (layer0_outputs[8083]) & ~(layer0_outputs[6484]);
    assign layer1_outputs[12404] = ~(layer0_outputs[8095]);
    assign layer1_outputs[12405] = (layer0_outputs[11621]) & (layer0_outputs[11448]);
    assign layer1_outputs[12406] = ~((layer0_outputs[2757]) ^ (layer0_outputs[928]));
    assign layer1_outputs[12407] = (layer0_outputs[8451]) | (layer0_outputs[5820]);
    assign layer1_outputs[12408] = (layer0_outputs[7461]) & ~(layer0_outputs[12288]);
    assign layer1_outputs[12409] = (layer0_outputs[5897]) ^ (layer0_outputs[12462]);
    assign layer1_outputs[12410] = ~(layer0_outputs[5917]);
    assign layer1_outputs[12411] = (layer0_outputs[8952]) ^ (layer0_outputs[8113]);
    assign layer1_outputs[12412] = ~(layer0_outputs[3492]);
    assign layer1_outputs[12413] = ~(layer0_outputs[6526]);
    assign layer1_outputs[12414] = (layer0_outputs[2680]) | (layer0_outputs[7448]);
    assign layer1_outputs[12415] = ~(layer0_outputs[12170]);
    assign layer1_outputs[12416] = ~(layer0_outputs[10251]);
    assign layer1_outputs[12417] = ~((layer0_outputs[5116]) & (layer0_outputs[12139]));
    assign layer1_outputs[12418] = 1'b1;
    assign layer1_outputs[12419] = ~(layer0_outputs[11869]);
    assign layer1_outputs[12420] = ~(layer0_outputs[8098]);
    assign layer1_outputs[12421] = 1'b0;
    assign layer1_outputs[12422] = (layer0_outputs[8589]) & ~(layer0_outputs[3985]);
    assign layer1_outputs[12423] = (layer0_outputs[3416]) & (layer0_outputs[3217]);
    assign layer1_outputs[12424] = layer0_outputs[8349];
    assign layer1_outputs[12425] = ~(layer0_outputs[4764]);
    assign layer1_outputs[12426] = ~(layer0_outputs[10956]) | (layer0_outputs[4190]);
    assign layer1_outputs[12427] = (layer0_outputs[3302]) & ~(layer0_outputs[10521]);
    assign layer1_outputs[12428] = layer0_outputs[12645];
    assign layer1_outputs[12429] = (layer0_outputs[8534]) & ~(layer0_outputs[3160]);
    assign layer1_outputs[12430] = (layer0_outputs[6037]) & ~(layer0_outputs[10966]);
    assign layer1_outputs[12431] = ~((layer0_outputs[1837]) & (layer0_outputs[602]));
    assign layer1_outputs[12432] = ~(layer0_outputs[965]);
    assign layer1_outputs[12433] = (layer0_outputs[8139]) ^ (layer0_outputs[2451]);
    assign layer1_outputs[12434] = (layer0_outputs[3587]) & ~(layer0_outputs[2047]);
    assign layer1_outputs[12435] = layer0_outputs[662];
    assign layer1_outputs[12436] = ~(layer0_outputs[712]);
    assign layer1_outputs[12437] = ~(layer0_outputs[2732]) | (layer0_outputs[11818]);
    assign layer1_outputs[12438] = (layer0_outputs[2954]) & (layer0_outputs[5314]);
    assign layer1_outputs[12439] = layer0_outputs[11152];
    assign layer1_outputs[12440] = layer0_outputs[12113];
    assign layer1_outputs[12441] = ~(layer0_outputs[8858]) | (layer0_outputs[2849]);
    assign layer1_outputs[12442] = ~((layer0_outputs[4072]) ^ (layer0_outputs[2750]));
    assign layer1_outputs[12443] = (layer0_outputs[5041]) & (layer0_outputs[2037]);
    assign layer1_outputs[12444] = (layer0_outputs[9208]) ^ (layer0_outputs[1769]);
    assign layer1_outputs[12445] = layer0_outputs[3195];
    assign layer1_outputs[12446] = (layer0_outputs[3709]) ^ (layer0_outputs[5650]);
    assign layer1_outputs[12447] = ~(layer0_outputs[7293]) | (layer0_outputs[11383]);
    assign layer1_outputs[12448] = (layer0_outputs[10067]) & (layer0_outputs[12219]);
    assign layer1_outputs[12449] = ~((layer0_outputs[4175]) & (layer0_outputs[7554]));
    assign layer1_outputs[12450] = ~(layer0_outputs[9327]);
    assign layer1_outputs[12451] = layer0_outputs[598];
    assign layer1_outputs[12452] = layer0_outputs[2865];
    assign layer1_outputs[12453] = (layer0_outputs[12081]) & ~(layer0_outputs[9201]);
    assign layer1_outputs[12454] = (layer0_outputs[302]) | (layer0_outputs[106]);
    assign layer1_outputs[12455] = (layer0_outputs[12104]) & (layer0_outputs[6374]);
    assign layer1_outputs[12456] = ~(layer0_outputs[1872]);
    assign layer1_outputs[12457] = layer0_outputs[11108];
    assign layer1_outputs[12458] = layer0_outputs[4097];
    assign layer1_outputs[12459] = layer0_outputs[10893];
    assign layer1_outputs[12460] = layer0_outputs[2196];
    assign layer1_outputs[12461] = (layer0_outputs[8208]) & ~(layer0_outputs[2974]);
    assign layer1_outputs[12462] = layer0_outputs[1437];
    assign layer1_outputs[12463] = layer0_outputs[5889];
    assign layer1_outputs[12464] = (layer0_outputs[7747]) & ~(layer0_outputs[2353]);
    assign layer1_outputs[12465] = ~((layer0_outputs[12167]) | (layer0_outputs[9343]));
    assign layer1_outputs[12466] = ~(layer0_outputs[5213]);
    assign layer1_outputs[12467] = ~(layer0_outputs[415]);
    assign layer1_outputs[12468] = (layer0_outputs[629]) & (layer0_outputs[4929]);
    assign layer1_outputs[12469] = ~(layer0_outputs[9139]) | (layer0_outputs[6797]);
    assign layer1_outputs[12470] = layer0_outputs[5824];
    assign layer1_outputs[12471] = ~((layer0_outputs[12351]) ^ (layer0_outputs[12755]));
    assign layer1_outputs[12472] = (layer0_outputs[3487]) & ~(layer0_outputs[2170]);
    assign layer1_outputs[12473] = layer0_outputs[3030];
    assign layer1_outputs[12474] = (layer0_outputs[9365]) & ~(layer0_outputs[6855]);
    assign layer1_outputs[12475] = layer0_outputs[3132];
    assign layer1_outputs[12476] = layer0_outputs[6112];
    assign layer1_outputs[12477] = ~(layer0_outputs[1108]);
    assign layer1_outputs[12478] = ~((layer0_outputs[4887]) | (layer0_outputs[1093]));
    assign layer1_outputs[12479] = layer0_outputs[440];
    assign layer1_outputs[12480] = ~(layer0_outputs[8442]) | (layer0_outputs[2584]);
    assign layer1_outputs[12481] = layer0_outputs[7542];
    assign layer1_outputs[12482] = ~(layer0_outputs[12042]);
    assign layer1_outputs[12483] = (layer0_outputs[210]) & ~(layer0_outputs[11900]);
    assign layer1_outputs[12484] = (layer0_outputs[11696]) | (layer0_outputs[9461]);
    assign layer1_outputs[12485] = ~(layer0_outputs[11475]);
    assign layer1_outputs[12486] = (layer0_outputs[6487]) ^ (layer0_outputs[8324]);
    assign layer1_outputs[12487] = (layer0_outputs[5189]) & ~(layer0_outputs[8143]);
    assign layer1_outputs[12488] = (layer0_outputs[1891]) & ~(layer0_outputs[4203]);
    assign layer1_outputs[12489] = (layer0_outputs[4748]) ^ (layer0_outputs[10914]);
    assign layer1_outputs[12490] = layer0_outputs[4331];
    assign layer1_outputs[12491] = ~((layer0_outputs[7000]) & (layer0_outputs[12188]));
    assign layer1_outputs[12492] = layer0_outputs[6559];
    assign layer1_outputs[12493] = (layer0_outputs[7983]) | (layer0_outputs[11391]);
    assign layer1_outputs[12494] = ~(layer0_outputs[8724]);
    assign layer1_outputs[12495] = ~(layer0_outputs[11005]);
    assign layer1_outputs[12496] = 1'b1;
    assign layer1_outputs[12497] = ~(layer0_outputs[4040]);
    assign layer1_outputs[12498] = layer0_outputs[3309];
    assign layer1_outputs[12499] = (layer0_outputs[4473]) & ~(layer0_outputs[3374]);
    assign layer1_outputs[12500] = (layer0_outputs[10269]) & ~(layer0_outputs[8782]);
    assign layer1_outputs[12501] = layer0_outputs[8107];
    assign layer1_outputs[12502] = ~((layer0_outputs[3604]) & (layer0_outputs[11554]));
    assign layer1_outputs[12503] = ~(layer0_outputs[4212]);
    assign layer1_outputs[12504] = (layer0_outputs[12574]) ^ (layer0_outputs[8550]);
    assign layer1_outputs[12505] = ~((layer0_outputs[11065]) & (layer0_outputs[2444]));
    assign layer1_outputs[12506] = (layer0_outputs[9714]) & ~(layer0_outputs[4792]);
    assign layer1_outputs[12507] = ~(layer0_outputs[11791]);
    assign layer1_outputs[12508] = (layer0_outputs[9399]) & ~(layer0_outputs[2231]);
    assign layer1_outputs[12509] = ~(layer0_outputs[10062]);
    assign layer1_outputs[12510] = ~((layer0_outputs[6775]) | (layer0_outputs[2367]));
    assign layer1_outputs[12511] = (layer0_outputs[2509]) ^ (layer0_outputs[3877]);
    assign layer1_outputs[12512] = ~((layer0_outputs[12263]) & (layer0_outputs[9338]));
    assign layer1_outputs[12513] = ~(layer0_outputs[2074]) | (layer0_outputs[11941]);
    assign layer1_outputs[12514] = (layer0_outputs[6574]) & (layer0_outputs[9773]);
    assign layer1_outputs[12515] = (layer0_outputs[8701]) | (layer0_outputs[10096]);
    assign layer1_outputs[12516] = (layer0_outputs[7186]) ^ (layer0_outputs[11701]);
    assign layer1_outputs[12517] = ~((layer0_outputs[2898]) ^ (layer0_outputs[8901]));
    assign layer1_outputs[12518] = ~(layer0_outputs[3612]);
    assign layer1_outputs[12519] = ~(layer0_outputs[6605]);
    assign layer1_outputs[12520] = ~((layer0_outputs[2825]) | (layer0_outputs[9729]));
    assign layer1_outputs[12521] = (layer0_outputs[816]) & (layer0_outputs[3719]);
    assign layer1_outputs[12522] = ~(layer0_outputs[5105]);
    assign layer1_outputs[12523] = ~(layer0_outputs[9813]);
    assign layer1_outputs[12524] = layer0_outputs[12460];
    assign layer1_outputs[12525] = ~((layer0_outputs[10585]) ^ (layer0_outputs[2063]));
    assign layer1_outputs[12526] = ~(layer0_outputs[5226]);
    assign layer1_outputs[12527] = ~(layer0_outputs[10540]);
    assign layer1_outputs[12528] = ~(layer0_outputs[9061]) | (layer0_outputs[8237]);
    assign layer1_outputs[12529] = ~((layer0_outputs[7527]) & (layer0_outputs[1904]));
    assign layer1_outputs[12530] = ~(layer0_outputs[12638]);
    assign layer1_outputs[12531] = ~((layer0_outputs[7915]) ^ (layer0_outputs[7248]));
    assign layer1_outputs[12532] = ~((layer0_outputs[10627]) & (layer0_outputs[6060]));
    assign layer1_outputs[12533] = layer0_outputs[8323];
    assign layer1_outputs[12534] = layer0_outputs[3359];
    assign layer1_outputs[12535] = ~(layer0_outputs[3045]) | (layer0_outputs[3185]);
    assign layer1_outputs[12536] = layer0_outputs[10212];
    assign layer1_outputs[12537] = ~(layer0_outputs[5444]) | (layer0_outputs[11437]);
    assign layer1_outputs[12538] = (layer0_outputs[11557]) ^ (layer0_outputs[6476]);
    assign layer1_outputs[12539] = ~((layer0_outputs[2719]) & (layer0_outputs[10970]));
    assign layer1_outputs[12540] = (layer0_outputs[9609]) & ~(layer0_outputs[12156]);
    assign layer1_outputs[12541] = ~(layer0_outputs[12030]) | (layer0_outputs[12305]);
    assign layer1_outputs[12542] = (layer0_outputs[12348]) ^ (layer0_outputs[1328]);
    assign layer1_outputs[12543] = layer0_outputs[9397];
    assign layer1_outputs[12544] = ~((layer0_outputs[4687]) & (layer0_outputs[8522]));
    assign layer1_outputs[12545] = ~(layer0_outputs[2181]) | (layer0_outputs[6107]);
    assign layer1_outputs[12546] = ~(layer0_outputs[12443]);
    assign layer1_outputs[12547] = layer0_outputs[9555];
    assign layer1_outputs[12548] = ~((layer0_outputs[7548]) & (layer0_outputs[3970]));
    assign layer1_outputs[12549] = layer0_outputs[895];
    assign layer1_outputs[12550] = ~((layer0_outputs[3458]) ^ (layer0_outputs[9278]));
    assign layer1_outputs[12551] = layer0_outputs[7341];
    assign layer1_outputs[12552] = ~((layer0_outputs[7267]) | (layer0_outputs[808]));
    assign layer1_outputs[12553] = ~(layer0_outputs[8790]) | (layer0_outputs[809]);
    assign layer1_outputs[12554] = (layer0_outputs[3771]) ^ (layer0_outputs[12278]);
    assign layer1_outputs[12555] = (layer0_outputs[3734]) & (layer0_outputs[3671]);
    assign layer1_outputs[12556] = layer0_outputs[6751];
    assign layer1_outputs[12557] = (layer0_outputs[11788]) ^ (layer0_outputs[12493]);
    assign layer1_outputs[12558] = (layer0_outputs[12233]) & ~(layer0_outputs[5857]);
    assign layer1_outputs[12559] = ~(layer0_outputs[4558]) | (layer0_outputs[44]);
    assign layer1_outputs[12560] = 1'b0;
    assign layer1_outputs[12561] = layer0_outputs[12262];
    assign layer1_outputs[12562] = ~(layer0_outputs[11981]);
    assign layer1_outputs[12563] = 1'b0;
    assign layer1_outputs[12564] = ~(layer0_outputs[11427]) | (layer0_outputs[10952]);
    assign layer1_outputs[12565] = ~(layer0_outputs[3499]) | (layer0_outputs[7310]);
    assign layer1_outputs[12566] = (layer0_outputs[34]) & ~(layer0_outputs[8317]);
    assign layer1_outputs[12567] = ~((layer0_outputs[8027]) ^ (layer0_outputs[8857]));
    assign layer1_outputs[12568] = layer0_outputs[111];
    assign layer1_outputs[12569] = (layer0_outputs[100]) & ~(layer0_outputs[6390]);
    assign layer1_outputs[12570] = ~(layer0_outputs[12283]);
    assign layer1_outputs[12571] = (layer0_outputs[12316]) | (layer0_outputs[2385]);
    assign layer1_outputs[12572] = ~((layer0_outputs[3489]) & (layer0_outputs[8674]));
    assign layer1_outputs[12573] = (layer0_outputs[6980]) & ~(layer0_outputs[4684]);
    assign layer1_outputs[12574] = ~(layer0_outputs[11643]);
    assign layer1_outputs[12575] = layer0_outputs[8564];
    assign layer1_outputs[12576] = ~(layer0_outputs[10982]);
    assign layer1_outputs[12577] = ~(layer0_outputs[4019]);
    assign layer1_outputs[12578] = ~((layer0_outputs[8988]) & (layer0_outputs[5908]));
    assign layer1_outputs[12579] = (layer0_outputs[8452]) ^ (layer0_outputs[2747]);
    assign layer1_outputs[12580] = (layer0_outputs[1460]) & (layer0_outputs[1495]);
    assign layer1_outputs[12581] = ~(layer0_outputs[8688]);
    assign layer1_outputs[12582] = (layer0_outputs[4386]) & ~(layer0_outputs[6741]);
    assign layer1_outputs[12583] = ~((layer0_outputs[7322]) | (layer0_outputs[8910]));
    assign layer1_outputs[12584] = layer0_outputs[12721];
    assign layer1_outputs[12585] = (layer0_outputs[5410]) | (layer0_outputs[357]);
    assign layer1_outputs[12586] = ~(layer0_outputs[12190]);
    assign layer1_outputs[12587] = ~(layer0_outputs[5076]) | (layer0_outputs[6542]);
    assign layer1_outputs[12588] = (layer0_outputs[3950]) & ~(layer0_outputs[3800]);
    assign layer1_outputs[12589] = ~((layer0_outputs[7905]) ^ (layer0_outputs[3722]));
    assign layer1_outputs[12590] = (layer0_outputs[9293]) & ~(layer0_outputs[9695]);
    assign layer1_outputs[12591] = (layer0_outputs[1657]) ^ (layer0_outputs[2622]);
    assign layer1_outputs[12592] = (layer0_outputs[9767]) & (layer0_outputs[9493]);
    assign layer1_outputs[12593] = ~((layer0_outputs[5560]) & (layer0_outputs[10566]));
    assign layer1_outputs[12594] = ~(layer0_outputs[7858]);
    assign layer1_outputs[12595] = (layer0_outputs[6873]) & ~(layer0_outputs[8972]);
    assign layer1_outputs[12596] = (layer0_outputs[1027]) | (layer0_outputs[6923]);
    assign layer1_outputs[12597] = ~(layer0_outputs[8315]) | (layer0_outputs[6863]);
    assign layer1_outputs[12598] = ~((layer0_outputs[1496]) | (layer0_outputs[5575]));
    assign layer1_outputs[12599] = ~(layer0_outputs[6300]);
    assign layer1_outputs[12600] = ~(layer0_outputs[4585]) | (layer0_outputs[9273]);
    assign layer1_outputs[12601] = ~((layer0_outputs[6426]) & (layer0_outputs[11009]));
    assign layer1_outputs[12602] = (layer0_outputs[11238]) | (layer0_outputs[5992]);
    assign layer1_outputs[12603] = ~(layer0_outputs[3695]) | (layer0_outputs[11651]);
    assign layer1_outputs[12604] = layer0_outputs[877];
    assign layer1_outputs[12605] = ~(layer0_outputs[10546]);
    assign layer1_outputs[12606] = (layer0_outputs[11164]) | (layer0_outputs[177]);
    assign layer1_outputs[12607] = (layer0_outputs[7081]) ^ (layer0_outputs[5704]);
    assign layer1_outputs[12608] = layer0_outputs[8275];
    assign layer1_outputs[12609] = ~(layer0_outputs[4785]) | (layer0_outputs[5067]);
    assign layer1_outputs[12610] = ~((layer0_outputs[9200]) & (layer0_outputs[4039]));
    assign layer1_outputs[12611] = (layer0_outputs[1988]) ^ (layer0_outputs[7769]);
    assign layer1_outputs[12612] = (layer0_outputs[7285]) & ~(layer0_outputs[8813]);
    assign layer1_outputs[12613] = ~((layer0_outputs[1264]) | (layer0_outputs[2610]));
    assign layer1_outputs[12614] = ~((layer0_outputs[11875]) | (layer0_outputs[11431]));
    assign layer1_outputs[12615] = ~(layer0_outputs[2521]);
    assign layer1_outputs[12616] = (layer0_outputs[10441]) ^ (layer0_outputs[3512]);
    assign layer1_outputs[12617] = (layer0_outputs[5909]) & ~(layer0_outputs[6337]);
    assign layer1_outputs[12618] = ~((layer0_outputs[780]) & (layer0_outputs[1364]));
    assign layer1_outputs[12619] = layer0_outputs[5737];
    assign layer1_outputs[12620] = ~(layer0_outputs[10245]);
    assign layer1_outputs[12621] = (layer0_outputs[7430]) & ~(layer0_outputs[579]);
    assign layer1_outputs[12622] = (layer0_outputs[7707]) & ~(layer0_outputs[11186]);
    assign layer1_outputs[12623] = ~((layer0_outputs[8788]) & (layer0_outputs[1718]));
    assign layer1_outputs[12624] = layer0_outputs[7027];
    assign layer1_outputs[12625] = (layer0_outputs[8145]) & ~(layer0_outputs[11664]);
    assign layer1_outputs[12626] = ~(layer0_outputs[3568]);
    assign layer1_outputs[12627] = ~(layer0_outputs[12325]) | (layer0_outputs[4047]);
    assign layer1_outputs[12628] = ~(layer0_outputs[8206]);
    assign layer1_outputs[12629] = layer0_outputs[3355];
    assign layer1_outputs[12630] = (layer0_outputs[9923]) & ~(layer0_outputs[10259]);
    assign layer1_outputs[12631] = ~(layer0_outputs[8940]) | (layer0_outputs[7666]);
    assign layer1_outputs[12632] = ~(layer0_outputs[8995]) | (layer0_outputs[9362]);
    assign layer1_outputs[12633] = ~(layer0_outputs[9670]);
    assign layer1_outputs[12634] = (layer0_outputs[1341]) | (layer0_outputs[8560]);
    assign layer1_outputs[12635] = layer0_outputs[9520];
    assign layer1_outputs[12636] = layer0_outputs[1638];
    assign layer1_outputs[12637] = (layer0_outputs[5839]) & ~(layer0_outputs[3487]);
    assign layer1_outputs[12638] = ~(layer0_outputs[1053]);
    assign layer1_outputs[12639] = ~(layer0_outputs[8189]);
    assign layer1_outputs[12640] = ~(layer0_outputs[6504]);
    assign layer1_outputs[12641] = ~(layer0_outputs[9983]) | (layer0_outputs[11528]);
    assign layer1_outputs[12642] = ~((layer0_outputs[1823]) & (layer0_outputs[7321]));
    assign layer1_outputs[12643] = (layer0_outputs[8369]) ^ (layer0_outputs[3931]);
    assign layer1_outputs[12644] = ~(layer0_outputs[12561]);
    assign layer1_outputs[12645] = ~(layer0_outputs[10831]) | (layer0_outputs[4276]);
    assign layer1_outputs[12646] = ~(layer0_outputs[11540]) | (layer0_outputs[8064]);
    assign layer1_outputs[12647] = ~((layer0_outputs[11059]) & (layer0_outputs[4888]));
    assign layer1_outputs[12648] = (layer0_outputs[872]) & ~(layer0_outputs[5291]);
    assign layer1_outputs[12649] = layer0_outputs[4431];
    assign layer1_outputs[12650] = ~((layer0_outputs[7578]) & (layer0_outputs[5616]));
    assign layer1_outputs[12651] = layer0_outputs[11096];
    assign layer1_outputs[12652] = ~(layer0_outputs[2790]);
    assign layer1_outputs[12653] = ~((layer0_outputs[12686]) ^ (layer0_outputs[5349]));
    assign layer1_outputs[12654] = ~(layer0_outputs[5531]);
    assign layer1_outputs[12655] = ~(layer0_outputs[8656]) | (layer0_outputs[10319]);
    assign layer1_outputs[12656] = ~(layer0_outputs[5870]);
    assign layer1_outputs[12657] = ~((layer0_outputs[10028]) ^ (layer0_outputs[12455]));
    assign layer1_outputs[12658] = layer0_outputs[7739];
    assign layer1_outputs[12659] = ~(layer0_outputs[170]);
    assign layer1_outputs[12660] = layer0_outputs[6422];
    assign layer1_outputs[12661] = ~((layer0_outputs[2458]) & (layer0_outputs[4518]));
    assign layer1_outputs[12662] = layer0_outputs[5453];
    assign layer1_outputs[12663] = ~(layer0_outputs[1066]) | (layer0_outputs[4439]);
    assign layer1_outputs[12664] = (layer0_outputs[10783]) & ~(layer0_outputs[2398]);
    assign layer1_outputs[12665] = ~(layer0_outputs[6981]);
    assign layer1_outputs[12666] = ~((layer0_outputs[7381]) & (layer0_outputs[12550]));
    assign layer1_outputs[12667] = (layer0_outputs[12644]) & ~(layer0_outputs[10012]);
    assign layer1_outputs[12668] = ~(layer0_outputs[5755]);
    assign layer1_outputs[12669] = (layer0_outputs[6937]) & (layer0_outputs[11234]);
    assign layer1_outputs[12670] = ~((layer0_outputs[9763]) | (layer0_outputs[10737]));
    assign layer1_outputs[12671] = ~((layer0_outputs[1707]) & (layer0_outputs[7119]));
    assign layer1_outputs[12672] = ~(layer0_outputs[10963]);
    assign layer1_outputs[12673] = ~(layer0_outputs[3953]) | (layer0_outputs[3906]);
    assign layer1_outputs[12674] = (layer0_outputs[10733]) ^ (layer0_outputs[5316]);
    assign layer1_outputs[12675] = ~(layer0_outputs[12121]);
    assign layer1_outputs[12676] = layer0_outputs[4837];
    assign layer1_outputs[12677] = layer0_outputs[7959];
    assign layer1_outputs[12678] = layer0_outputs[10131];
    assign layer1_outputs[12679] = (layer0_outputs[3721]) & ~(layer0_outputs[9528]);
    assign layer1_outputs[12680] = layer0_outputs[2851];
    assign layer1_outputs[12681] = layer0_outputs[4071];
    assign layer1_outputs[12682] = ~(layer0_outputs[12500]);
    assign layer1_outputs[12683] = layer0_outputs[2028];
    assign layer1_outputs[12684] = ~(layer0_outputs[10827]) | (layer0_outputs[4151]);
    assign layer1_outputs[12685] = (layer0_outputs[11499]) & ~(layer0_outputs[1126]);
    assign layer1_outputs[12686] = (layer0_outputs[8786]) ^ (layer0_outputs[8836]);
    assign layer1_outputs[12687] = ~((layer0_outputs[7838]) | (layer0_outputs[8636]));
    assign layer1_outputs[12688] = layer0_outputs[9896];
    assign layer1_outputs[12689] = ~(layer0_outputs[4092]);
    assign layer1_outputs[12690] = layer0_outputs[174];
    assign layer1_outputs[12691] = ~(layer0_outputs[5879]);
    assign layer1_outputs[12692] = layer0_outputs[11764];
    assign layer1_outputs[12693] = ~((layer0_outputs[280]) ^ (layer0_outputs[9558]));
    assign layer1_outputs[12694] = ~((layer0_outputs[9279]) | (layer0_outputs[6682]));
    assign layer1_outputs[12695] = ~(layer0_outputs[10736]) | (layer0_outputs[2121]);
    assign layer1_outputs[12696] = (layer0_outputs[1486]) & (layer0_outputs[1772]);
    assign layer1_outputs[12697] = ~((layer0_outputs[7246]) & (layer0_outputs[11850]));
    assign layer1_outputs[12698] = (layer0_outputs[2033]) | (layer0_outputs[11795]);
    assign layer1_outputs[12699] = ~((layer0_outputs[5581]) & (layer0_outputs[11738]));
    assign layer1_outputs[12700] = layer0_outputs[4808];
    assign layer1_outputs[12701] = (layer0_outputs[49]) & (layer0_outputs[11920]);
    assign layer1_outputs[12702] = 1'b0;
    assign layer1_outputs[12703] = layer0_outputs[4851];
    assign layer1_outputs[12704] = ~(layer0_outputs[479]);
    assign layer1_outputs[12705] = ~((layer0_outputs[5651]) ^ (layer0_outputs[10983]));
    assign layer1_outputs[12706] = ~(layer0_outputs[4611]);
    assign layer1_outputs[12707] = layer0_outputs[12413];
    assign layer1_outputs[12708] = ~(layer0_outputs[8673]);
    assign layer1_outputs[12709] = ~(layer0_outputs[6475]) | (layer0_outputs[3182]);
    assign layer1_outputs[12710] = ~((layer0_outputs[1691]) | (layer0_outputs[7821]));
    assign layer1_outputs[12711] = ~(layer0_outputs[5788]) | (layer0_outputs[6213]);
    assign layer1_outputs[12712] = (layer0_outputs[2002]) & (layer0_outputs[10855]);
    assign layer1_outputs[12713] = (layer0_outputs[11591]) & (layer0_outputs[4300]);
    assign layer1_outputs[12714] = ~(layer0_outputs[3653]);
    assign layer1_outputs[12715] = ~((layer0_outputs[11368]) & (layer0_outputs[11022]));
    assign layer1_outputs[12716] = layer0_outputs[10236];
    assign layer1_outputs[12717] = ~(layer0_outputs[542]) | (layer0_outputs[6501]);
    assign layer1_outputs[12718] = (layer0_outputs[1349]) & ~(layer0_outputs[4784]);
    assign layer1_outputs[12719] = layer0_outputs[2130];
    assign layer1_outputs[12720] = ~((layer0_outputs[11150]) & (layer0_outputs[2677]));
    assign layer1_outputs[12721] = ~((layer0_outputs[7173]) & (layer0_outputs[9737]));
    assign layer1_outputs[12722] = ~(layer0_outputs[7250]);
    assign layer1_outputs[12723] = (layer0_outputs[7251]) & ~(layer0_outputs[9759]);
    assign layer1_outputs[12724] = ~((layer0_outputs[11294]) & (layer0_outputs[4143]));
    assign layer1_outputs[12725] = (layer0_outputs[10837]) & ~(layer0_outputs[11862]);
    assign layer1_outputs[12726] = (layer0_outputs[10762]) & ~(layer0_outputs[7389]);
    assign layer1_outputs[12727] = layer0_outputs[12493];
    assign layer1_outputs[12728] = ~((layer0_outputs[2474]) & (layer0_outputs[1265]));
    assign layer1_outputs[12729] = 1'b1;
    assign layer1_outputs[12730] = ~(layer0_outputs[10457]) | (layer0_outputs[3316]);
    assign layer1_outputs[12731] = 1'b0;
    assign layer1_outputs[12732] = ~((layer0_outputs[6361]) | (layer0_outputs[8939]));
    assign layer1_outputs[12733] = layer0_outputs[5697];
    assign layer1_outputs[12734] = (layer0_outputs[6721]) ^ (layer0_outputs[187]);
    assign layer1_outputs[12735] = layer0_outputs[578];
    assign layer1_outputs[12736] = (layer0_outputs[9328]) & ~(layer0_outputs[11505]);
    assign layer1_outputs[12737] = layer0_outputs[8190];
    assign layer1_outputs[12738] = (layer0_outputs[5428]) & (layer0_outputs[10593]);
    assign layer1_outputs[12739] = ~((layer0_outputs[4578]) & (layer0_outputs[1254]));
    assign layer1_outputs[12740] = layer0_outputs[9025];
    assign layer1_outputs[12741] = ~((layer0_outputs[205]) & (layer0_outputs[4680]));
    assign layer1_outputs[12742] = layer0_outputs[5626];
    assign layer1_outputs[12743] = 1'b0;
    assign layer1_outputs[12744] = (layer0_outputs[12187]) & (layer0_outputs[4647]);
    assign layer1_outputs[12745] = (layer0_outputs[2096]) & ~(layer0_outputs[3949]);
    assign layer1_outputs[12746] = layer0_outputs[1135];
    assign layer1_outputs[12747] = ~((layer0_outputs[10060]) & (layer0_outputs[7845]));
    assign layer1_outputs[12748] = ~(layer0_outputs[7253]);
    assign layer1_outputs[12749] = (layer0_outputs[12277]) ^ (layer0_outputs[9971]);
    assign layer1_outputs[12750] = (layer0_outputs[4991]) & ~(layer0_outputs[10947]);
    assign layer1_outputs[12751] = 1'b1;
    assign layer1_outputs[12752] = ~(layer0_outputs[9426]) | (layer0_outputs[12321]);
    assign layer1_outputs[12753] = layer0_outputs[2955];
    assign layer1_outputs[12754] = (layer0_outputs[6670]) & ~(layer0_outputs[6302]);
    assign layer1_outputs[12755] = ~(layer0_outputs[8823]);
    assign layer1_outputs[12756] = ~(layer0_outputs[3263]) | (layer0_outputs[943]);
    assign layer1_outputs[12757] = (layer0_outputs[4693]) ^ (layer0_outputs[257]);
    assign layer1_outputs[12758] = (layer0_outputs[539]) & ~(layer0_outputs[2645]);
    assign layer1_outputs[12759] = (layer0_outputs[2361]) & (layer0_outputs[10091]);
    assign layer1_outputs[12760] = ~(layer0_outputs[10416]);
    assign layer1_outputs[12761] = (layer0_outputs[855]) & ~(layer0_outputs[7264]);
    assign layer1_outputs[12762] = (layer0_outputs[9198]) & ~(layer0_outputs[2048]);
    assign layer1_outputs[12763] = (layer0_outputs[2360]) & ~(layer0_outputs[11873]);
    assign layer1_outputs[12764] = ~((layer0_outputs[6454]) ^ (layer0_outputs[11228]));
    assign layer1_outputs[12765] = ~((layer0_outputs[8341]) | (layer0_outputs[2060]));
    assign layer1_outputs[12766] = ~(layer0_outputs[10283]);
    assign layer1_outputs[12767] = ~((layer0_outputs[9662]) ^ (layer0_outputs[5733]));
    assign layer1_outputs[12768] = layer0_outputs[11515];
    assign layer1_outputs[12769] = ~(layer0_outputs[7277]);
    assign layer1_outputs[12770] = (layer0_outputs[47]) & ~(layer0_outputs[8810]);
    assign layer1_outputs[12771] = (layer0_outputs[937]) & ~(layer0_outputs[6007]);
    assign layer1_outputs[12772] = (layer0_outputs[4970]) & ~(layer0_outputs[8726]);
    assign layer1_outputs[12773] = (layer0_outputs[10499]) | (layer0_outputs[12434]);
    assign layer1_outputs[12774] = ~(layer0_outputs[7914]) | (layer0_outputs[11862]);
    assign layer1_outputs[12775] = ~((layer0_outputs[10136]) & (layer0_outputs[258]));
    assign layer1_outputs[12776] = ~(layer0_outputs[11553]) | (layer0_outputs[9023]);
    assign layer1_outputs[12777] = layer0_outputs[7984];
    assign layer1_outputs[12778] = ~(layer0_outputs[5066]);
    assign layer1_outputs[12779] = layer0_outputs[3252];
    assign layer1_outputs[12780] = ~(layer0_outputs[11309]);
    assign layer1_outputs[12781] = (layer0_outputs[5408]) | (layer0_outputs[3271]);
    assign layer1_outputs[12782] = (layer0_outputs[12111]) & (layer0_outputs[3934]);
    assign layer1_outputs[12783] = ~(layer0_outputs[2120]);
    assign layer1_outputs[12784] = ~(layer0_outputs[2638]);
    assign layer1_outputs[12785] = ~(layer0_outputs[8205]);
    assign layer1_outputs[12786] = ~(layer0_outputs[10234]);
    assign layer1_outputs[12787] = (layer0_outputs[554]) & ~(layer0_outputs[9366]);
    assign layer1_outputs[12788] = ~(layer0_outputs[5016]);
    assign layer1_outputs[12789] = layer0_outputs[5770];
    assign layer1_outputs[12790] = ~((layer0_outputs[3768]) | (layer0_outputs[8586]));
    assign layer1_outputs[12791] = ~((layer0_outputs[11340]) | (layer0_outputs[1034]));
    assign layer1_outputs[12792] = ~(layer0_outputs[5310]);
    assign layer1_outputs[12793] = ~(layer0_outputs[1490]) | (layer0_outputs[3625]);
    assign layer1_outputs[12794] = ~(layer0_outputs[9211]);
    assign layer1_outputs[12795] = ~(layer0_outputs[257]);
    assign layer1_outputs[12796] = (layer0_outputs[6331]) & ~(layer0_outputs[1827]);
    assign layer1_outputs[12797] = layer0_outputs[10215];
    assign layer1_outputs[12798] = ~(layer0_outputs[1767]) | (layer0_outputs[7127]);
    assign layer1_outputs[12799] = ~(layer0_outputs[12524]);
    assign layer2_outputs[0] = layer1_outputs[5610];
    assign layer2_outputs[1] = ~((layer1_outputs[6367]) & (layer1_outputs[8112]));
    assign layer2_outputs[2] = layer1_outputs[2629];
    assign layer2_outputs[3] = layer1_outputs[4634];
    assign layer2_outputs[4] = ~(layer1_outputs[723]);
    assign layer2_outputs[5] = ~(layer1_outputs[3399]);
    assign layer2_outputs[6] = (layer1_outputs[8317]) & ~(layer1_outputs[7366]);
    assign layer2_outputs[7] = ~(layer1_outputs[3896]);
    assign layer2_outputs[8] = (layer1_outputs[3767]) & ~(layer1_outputs[2774]);
    assign layer2_outputs[9] = ~(layer1_outputs[12121]);
    assign layer2_outputs[10] = ~((layer1_outputs[3344]) | (layer1_outputs[8473]));
    assign layer2_outputs[11] = layer1_outputs[451];
    assign layer2_outputs[12] = layer1_outputs[1371];
    assign layer2_outputs[13] = ~((layer1_outputs[8428]) ^ (layer1_outputs[9939]));
    assign layer2_outputs[14] = ~(layer1_outputs[3952]);
    assign layer2_outputs[15] = layer1_outputs[5963];
    assign layer2_outputs[16] = ~(layer1_outputs[8704]);
    assign layer2_outputs[17] = ~((layer1_outputs[4949]) ^ (layer1_outputs[10257]));
    assign layer2_outputs[18] = (layer1_outputs[8497]) & (layer1_outputs[4733]);
    assign layer2_outputs[19] = ~((layer1_outputs[2730]) & (layer1_outputs[1542]));
    assign layer2_outputs[20] = (layer1_outputs[4342]) & ~(layer1_outputs[6110]);
    assign layer2_outputs[21] = layer1_outputs[6504];
    assign layer2_outputs[22] = ~(layer1_outputs[3606]);
    assign layer2_outputs[23] = ~(layer1_outputs[4936]);
    assign layer2_outputs[24] = ~(layer1_outputs[6315]) | (layer1_outputs[7331]);
    assign layer2_outputs[25] = ~(layer1_outputs[9918]);
    assign layer2_outputs[26] = layer1_outputs[6206];
    assign layer2_outputs[27] = ~((layer1_outputs[257]) ^ (layer1_outputs[12126]));
    assign layer2_outputs[28] = layer1_outputs[181];
    assign layer2_outputs[29] = layer1_outputs[7604];
    assign layer2_outputs[30] = ~(layer1_outputs[1409]);
    assign layer2_outputs[31] = ~(layer1_outputs[8576]);
    assign layer2_outputs[32] = layer1_outputs[6177];
    assign layer2_outputs[33] = layer1_outputs[1632];
    assign layer2_outputs[34] = layer1_outputs[221];
    assign layer2_outputs[35] = ~(layer1_outputs[11843]);
    assign layer2_outputs[36] = (layer1_outputs[5418]) & ~(layer1_outputs[10480]);
    assign layer2_outputs[37] = ~(layer1_outputs[10531]);
    assign layer2_outputs[38] = (layer1_outputs[8550]) ^ (layer1_outputs[5982]);
    assign layer2_outputs[39] = ~(layer1_outputs[11333]) | (layer1_outputs[7826]);
    assign layer2_outputs[40] = layer1_outputs[10407];
    assign layer2_outputs[41] = ~((layer1_outputs[4961]) ^ (layer1_outputs[3056]));
    assign layer2_outputs[42] = ~(layer1_outputs[10796]);
    assign layer2_outputs[43] = ~(layer1_outputs[2538]);
    assign layer2_outputs[44] = ~((layer1_outputs[5492]) | (layer1_outputs[4718]));
    assign layer2_outputs[45] = layer1_outputs[4305];
    assign layer2_outputs[46] = ~(layer1_outputs[12014]);
    assign layer2_outputs[47] = (layer1_outputs[9920]) | (layer1_outputs[4331]);
    assign layer2_outputs[48] = ~(layer1_outputs[4857]);
    assign layer2_outputs[49] = ~((layer1_outputs[2856]) & (layer1_outputs[10446]));
    assign layer2_outputs[50] = (layer1_outputs[12591]) & (layer1_outputs[8933]);
    assign layer2_outputs[51] = layer1_outputs[3506];
    assign layer2_outputs[52] = layer1_outputs[8440];
    assign layer2_outputs[53] = (layer1_outputs[1724]) ^ (layer1_outputs[8664]);
    assign layer2_outputs[54] = ~(layer1_outputs[476]);
    assign layer2_outputs[55] = ~(layer1_outputs[11468]) | (layer1_outputs[2203]);
    assign layer2_outputs[56] = layer1_outputs[8432];
    assign layer2_outputs[57] = layer1_outputs[10703];
    assign layer2_outputs[58] = ~(layer1_outputs[4870]) | (layer1_outputs[4894]);
    assign layer2_outputs[59] = layer1_outputs[7237];
    assign layer2_outputs[60] = (layer1_outputs[9579]) ^ (layer1_outputs[12155]);
    assign layer2_outputs[61] = ~(layer1_outputs[8347]);
    assign layer2_outputs[62] = ~(layer1_outputs[4974]);
    assign layer2_outputs[63] = (layer1_outputs[12306]) & (layer1_outputs[10069]);
    assign layer2_outputs[64] = (layer1_outputs[5810]) & ~(layer1_outputs[5795]);
    assign layer2_outputs[65] = layer1_outputs[11013];
    assign layer2_outputs[66] = layer1_outputs[12480];
    assign layer2_outputs[67] = ~(layer1_outputs[4008]);
    assign layer2_outputs[68] = ~(layer1_outputs[1482]);
    assign layer2_outputs[69] = ~(layer1_outputs[7308]);
    assign layer2_outputs[70] = ~((layer1_outputs[7502]) ^ (layer1_outputs[6941]));
    assign layer2_outputs[71] = ~((layer1_outputs[9242]) & (layer1_outputs[5398]));
    assign layer2_outputs[72] = layer1_outputs[1379];
    assign layer2_outputs[73] = layer1_outputs[7412];
    assign layer2_outputs[74] = layer1_outputs[1016];
    assign layer2_outputs[75] = layer1_outputs[6561];
    assign layer2_outputs[76] = (layer1_outputs[2846]) & ~(layer1_outputs[9105]);
    assign layer2_outputs[77] = ~(layer1_outputs[5417]);
    assign layer2_outputs[78] = (layer1_outputs[9820]) & (layer1_outputs[12729]);
    assign layer2_outputs[79] = (layer1_outputs[3071]) & ~(layer1_outputs[11888]);
    assign layer2_outputs[80] = (layer1_outputs[4735]) | (layer1_outputs[10739]);
    assign layer2_outputs[81] = ~((layer1_outputs[10866]) ^ (layer1_outputs[8041]));
    assign layer2_outputs[82] = ~(layer1_outputs[3111]);
    assign layer2_outputs[83] = ~((layer1_outputs[1860]) | (layer1_outputs[12558]));
    assign layer2_outputs[84] = (layer1_outputs[8007]) & ~(layer1_outputs[9099]);
    assign layer2_outputs[85] = ~(layer1_outputs[5386]);
    assign layer2_outputs[86] = 1'b1;
    assign layer2_outputs[87] = ~((layer1_outputs[10462]) ^ (layer1_outputs[2095]));
    assign layer2_outputs[88] = ~((layer1_outputs[10147]) ^ (layer1_outputs[9515]));
    assign layer2_outputs[89] = ~((layer1_outputs[11632]) ^ (layer1_outputs[0]));
    assign layer2_outputs[90] = (layer1_outputs[5848]) ^ (layer1_outputs[9677]);
    assign layer2_outputs[91] = ~(layer1_outputs[1807]);
    assign layer2_outputs[92] = (layer1_outputs[2932]) & (layer1_outputs[12716]);
    assign layer2_outputs[93] = layer1_outputs[4432];
    assign layer2_outputs[94] = ~(layer1_outputs[5301]);
    assign layer2_outputs[95] = (layer1_outputs[2849]) | (layer1_outputs[7745]);
    assign layer2_outputs[96] = layer1_outputs[2034];
    assign layer2_outputs[97] = ~(layer1_outputs[12291]) | (layer1_outputs[10882]);
    assign layer2_outputs[98] = (layer1_outputs[3243]) & ~(layer1_outputs[12700]);
    assign layer2_outputs[99] = ~(layer1_outputs[7212]);
    assign layer2_outputs[100] = (layer1_outputs[2669]) | (layer1_outputs[875]);
    assign layer2_outputs[101] = (layer1_outputs[6695]) | (layer1_outputs[6401]);
    assign layer2_outputs[102] = (layer1_outputs[6564]) ^ (layer1_outputs[11673]);
    assign layer2_outputs[103] = ~((layer1_outputs[12775]) | (layer1_outputs[2918]));
    assign layer2_outputs[104] = (layer1_outputs[9414]) & ~(layer1_outputs[8274]);
    assign layer2_outputs[105] = ~((layer1_outputs[2423]) | (layer1_outputs[6733]));
    assign layer2_outputs[106] = ~(layer1_outputs[12652]);
    assign layer2_outputs[107] = layer1_outputs[10492];
    assign layer2_outputs[108] = layer1_outputs[5412];
    assign layer2_outputs[109] = (layer1_outputs[6459]) | (layer1_outputs[7526]);
    assign layer2_outputs[110] = (layer1_outputs[3368]) ^ (layer1_outputs[3345]);
    assign layer2_outputs[111] = ~((layer1_outputs[6106]) ^ (layer1_outputs[173]));
    assign layer2_outputs[112] = layer1_outputs[762];
    assign layer2_outputs[113] = ~(layer1_outputs[1745]) | (layer1_outputs[9651]);
    assign layer2_outputs[114] = (layer1_outputs[3802]) & ~(layer1_outputs[3800]);
    assign layer2_outputs[115] = (layer1_outputs[1118]) & ~(layer1_outputs[12721]);
    assign layer2_outputs[116] = layer1_outputs[8645];
    assign layer2_outputs[117] = (layer1_outputs[8731]) & ~(layer1_outputs[4135]);
    assign layer2_outputs[118] = (layer1_outputs[11456]) & (layer1_outputs[18]);
    assign layer2_outputs[119] = ~(layer1_outputs[1771]);
    assign layer2_outputs[120] = ~(layer1_outputs[3239]);
    assign layer2_outputs[121] = layer1_outputs[10856];
    assign layer2_outputs[122] = ~((layer1_outputs[11235]) & (layer1_outputs[11993]));
    assign layer2_outputs[123] = ~(layer1_outputs[2942]);
    assign layer2_outputs[124] = (layer1_outputs[2154]) & ~(layer1_outputs[1760]);
    assign layer2_outputs[125] = ~(layer1_outputs[11778]) | (layer1_outputs[2448]);
    assign layer2_outputs[126] = layer1_outputs[2078];
    assign layer2_outputs[127] = ~((layer1_outputs[11825]) | (layer1_outputs[4267]));
    assign layer2_outputs[128] = ~(layer1_outputs[8325]) | (layer1_outputs[1013]);
    assign layer2_outputs[129] = (layer1_outputs[8489]) & ~(layer1_outputs[529]);
    assign layer2_outputs[130] = (layer1_outputs[6834]) | (layer1_outputs[4653]);
    assign layer2_outputs[131] = layer1_outputs[8737];
    assign layer2_outputs[132] = ~(layer1_outputs[10337]);
    assign layer2_outputs[133] = ~(layer1_outputs[4618]);
    assign layer2_outputs[134] = ~(layer1_outputs[10490]);
    assign layer2_outputs[135] = layer1_outputs[1668];
    assign layer2_outputs[136] = ~((layer1_outputs[1987]) & (layer1_outputs[10625]));
    assign layer2_outputs[137] = layer1_outputs[11850];
    assign layer2_outputs[138] = (layer1_outputs[1743]) | (layer1_outputs[4885]);
    assign layer2_outputs[139] = ~(layer1_outputs[10997]);
    assign layer2_outputs[140] = ~(layer1_outputs[788]) | (layer1_outputs[2350]);
    assign layer2_outputs[141] = (layer1_outputs[12252]) & (layer1_outputs[12616]);
    assign layer2_outputs[142] = (layer1_outputs[11757]) ^ (layer1_outputs[4696]);
    assign layer2_outputs[143] = layer1_outputs[7533];
    assign layer2_outputs[144] = layer1_outputs[5047];
    assign layer2_outputs[145] = layer1_outputs[8617];
    assign layer2_outputs[146] = ~(layer1_outputs[12686]);
    assign layer2_outputs[147] = ~((layer1_outputs[4803]) ^ (layer1_outputs[4770]));
    assign layer2_outputs[148] = (layer1_outputs[4284]) & ~(layer1_outputs[8164]);
    assign layer2_outputs[149] = ~(layer1_outputs[2931]);
    assign layer2_outputs[150] = layer1_outputs[3066];
    assign layer2_outputs[151] = ~(layer1_outputs[1183]);
    assign layer2_outputs[152] = layer1_outputs[12296];
    assign layer2_outputs[153] = layer1_outputs[8310];
    assign layer2_outputs[154] = layer1_outputs[8028];
    assign layer2_outputs[155] = ~(layer1_outputs[6698]);
    assign layer2_outputs[156] = ~(layer1_outputs[6400]);
    assign layer2_outputs[157] = ~(layer1_outputs[10976]);
    assign layer2_outputs[158] = ~((layer1_outputs[12519]) ^ (layer1_outputs[9527]));
    assign layer2_outputs[159] = ~(layer1_outputs[6922]);
    assign layer2_outputs[160] = (layer1_outputs[3957]) ^ (layer1_outputs[11907]);
    assign layer2_outputs[161] = 1'b0;
    assign layer2_outputs[162] = layer1_outputs[3387];
    assign layer2_outputs[163] = ~(layer1_outputs[8214]);
    assign layer2_outputs[164] = ~((layer1_outputs[693]) ^ (layer1_outputs[2534]));
    assign layer2_outputs[165] = (layer1_outputs[4079]) & ~(layer1_outputs[1820]);
    assign layer2_outputs[166] = (layer1_outputs[3470]) & ~(layer1_outputs[10289]);
    assign layer2_outputs[167] = layer1_outputs[5426];
    assign layer2_outputs[168] = layer1_outputs[1400];
    assign layer2_outputs[169] = (layer1_outputs[7134]) | (layer1_outputs[5555]);
    assign layer2_outputs[170] = ~(layer1_outputs[3648]);
    assign layer2_outputs[171] = ~(layer1_outputs[10343]) | (layer1_outputs[4676]);
    assign layer2_outputs[172] = (layer1_outputs[10339]) & (layer1_outputs[3915]);
    assign layer2_outputs[173] = (layer1_outputs[10829]) | (layer1_outputs[7176]);
    assign layer2_outputs[174] = ~(layer1_outputs[5370]);
    assign layer2_outputs[175] = ~(layer1_outputs[11798]);
    assign layer2_outputs[176] = ~((layer1_outputs[6391]) & (layer1_outputs[12771]));
    assign layer2_outputs[177] = ~(layer1_outputs[7217]);
    assign layer2_outputs[178] = ~(layer1_outputs[12188]) | (layer1_outputs[495]);
    assign layer2_outputs[179] = ~(layer1_outputs[10342]) | (layer1_outputs[9448]);
    assign layer2_outputs[180] = layer1_outputs[9410];
    assign layer2_outputs[181] = ~(layer1_outputs[2542]);
    assign layer2_outputs[182] = ~((layer1_outputs[9700]) & (layer1_outputs[4363]));
    assign layer2_outputs[183] = ~(layer1_outputs[11232]);
    assign layer2_outputs[184] = ~(layer1_outputs[2522]) | (layer1_outputs[5374]);
    assign layer2_outputs[185] = layer1_outputs[12508];
    assign layer2_outputs[186] = ~(layer1_outputs[7148]) | (layer1_outputs[2123]);
    assign layer2_outputs[187] = ~((layer1_outputs[8242]) | (layer1_outputs[1283]));
    assign layer2_outputs[188] = ~(layer1_outputs[6452]) | (layer1_outputs[8725]);
    assign layer2_outputs[189] = ~(layer1_outputs[10160]);
    assign layer2_outputs[190] = (layer1_outputs[2021]) & ~(layer1_outputs[6175]);
    assign layer2_outputs[191] = ~(layer1_outputs[7164]);
    assign layer2_outputs[192] = layer1_outputs[1930];
    assign layer2_outputs[193] = layer1_outputs[7260];
    assign layer2_outputs[194] = ~(layer1_outputs[9271]);
    assign layer2_outputs[195] = (layer1_outputs[71]) ^ (layer1_outputs[3466]);
    assign layer2_outputs[196] = layer1_outputs[4539];
    assign layer2_outputs[197] = layer1_outputs[7285];
    assign layer2_outputs[198] = (layer1_outputs[605]) & ~(layer1_outputs[6226]);
    assign layer2_outputs[199] = layer1_outputs[3313];
    assign layer2_outputs[200] = ~(layer1_outputs[10915]);
    assign layer2_outputs[201] = layer1_outputs[6156];
    assign layer2_outputs[202] = layer1_outputs[8585];
    assign layer2_outputs[203] = (layer1_outputs[2824]) | (layer1_outputs[4225]);
    assign layer2_outputs[204] = layer1_outputs[390];
    assign layer2_outputs[205] = layer1_outputs[5988];
    assign layer2_outputs[206] = layer1_outputs[2694];
    assign layer2_outputs[207] = ~(layer1_outputs[2725]);
    assign layer2_outputs[208] = layer1_outputs[8453];
    assign layer2_outputs[209] = ~(layer1_outputs[5412]);
    assign layer2_outputs[210] = ~((layer1_outputs[1619]) & (layer1_outputs[6741]));
    assign layer2_outputs[211] = ~(layer1_outputs[10500]) | (layer1_outputs[8635]);
    assign layer2_outputs[212] = ~((layer1_outputs[8299]) ^ (layer1_outputs[5922]));
    assign layer2_outputs[213] = (layer1_outputs[10053]) & ~(layer1_outputs[6859]);
    assign layer2_outputs[214] = ~(layer1_outputs[9252]);
    assign layer2_outputs[215] = ~((layer1_outputs[9394]) ^ (layer1_outputs[4593]));
    assign layer2_outputs[216] = layer1_outputs[11972];
    assign layer2_outputs[217] = (layer1_outputs[4968]) | (layer1_outputs[11270]);
    assign layer2_outputs[218] = ~(layer1_outputs[12445]);
    assign layer2_outputs[219] = ~(layer1_outputs[3914]);
    assign layer2_outputs[220] = ~(layer1_outputs[361]);
    assign layer2_outputs[221] = (layer1_outputs[2557]) & ~(layer1_outputs[7005]);
    assign layer2_outputs[222] = layer1_outputs[4812];
    assign layer2_outputs[223] = ~(layer1_outputs[11243]);
    assign layer2_outputs[224] = (layer1_outputs[5153]) | (layer1_outputs[5293]);
    assign layer2_outputs[225] = ~(layer1_outputs[8494]) | (layer1_outputs[6899]);
    assign layer2_outputs[226] = 1'b1;
    assign layer2_outputs[227] = layer1_outputs[1064];
    assign layer2_outputs[228] = layer1_outputs[3827];
    assign layer2_outputs[229] = layer1_outputs[97];
    assign layer2_outputs[230] = (layer1_outputs[607]) ^ (layer1_outputs[1933]);
    assign layer2_outputs[231] = ~(layer1_outputs[9991]);
    assign layer2_outputs[232] = ~((layer1_outputs[7291]) & (layer1_outputs[9567]));
    assign layer2_outputs[233] = ~((layer1_outputs[3098]) | (layer1_outputs[8548]));
    assign layer2_outputs[234] = ~(layer1_outputs[7274]) | (layer1_outputs[10986]);
    assign layer2_outputs[235] = layer1_outputs[6664];
    assign layer2_outputs[236] = ~(layer1_outputs[2274]);
    assign layer2_outputs[237] = ~(layer1_outputs[6080]);
    assign layer2_outputs[238] = ~(layer1_outputs[4185]) | (layer1_outputs[11221]);
    assign layer2_outputs[239] = (layer1_outputs[8160]) ^ (layer1_outputs[9248]);
    assign layer2_outputs[240] = ~(layer1_outputs[3361]);
    assign layer2_outputs[241] = ~((layer1_outputs[12345]) | (layer1_outputs[9152]));
    assign layer2_outputs[242] = ~(layer1_outputs[8193]);
    assign layer2_outputs[243] = ~((layer1_outputs[5727]) ^ (layer1_outputs[11261]));
    assign layer2_outputs[244] = (layer1_outputs[8919]) & ~(layer1_outputs[2131]);
    assign layer2_outputs[245] = layer1_outputs[4564];
    assign layer2_outputs[246] = ~((layer1_outputs[3705]) & (layer1_outputs[9784]));
    assign layer2_outputs[247] = ~(layer1_outputs[5724]);
    assign layer2_outputs[248] = ~(layer1_outputs[9906]);
    assign layer2_outputs[249] = layer1_outputs[10733];
    assign layer2_outputs[250] = (layer1_outputs[2986]) & (layer1_outputs[7425]);
    assign layer2_outputs[251] = (layer1_outputs[5564]) & ~(layer1_outputs[8619]);
    assign layer2_outputs[252] = (layer1_outputs[11757]) & ~(layer1_outputs[2863]);
    assign layer2_outputs[253] = ~(layer1_outputs[10073]);
    assign layer2_outputs[254] = ~(layer1_outputs[8541]);
    assign layer2_outputs[255] = layer1_outputs[2324];
    assign layer2_outputs[256] = (layer1_outputs[8988]) & (layer1_outputs[7]);
    assign layer2_outputs[257] = (layer1_outputs[6891]) & (layer1_outputs[4498]);
    assign layer2_outputs[258] = (layer1_outputs[8382]) & ~(layer1_outputs[4405]);
    assign layer2_outputs[259] = layer1_outputs[3021];
    assign layer2_outputs[260] = (layer1_outputs[1740]) & ~(layer1_outputs[3437]);
    assign layer2_outputs[261] = layer1_outputs[7417];
    assign layer2_outputs[262] = layer1_outputs[10785];
    assign layer2_outputs[263] = layer1_outputs[11809];
    assign layer2_outputs[264] = ~(layer1_outputs[12368]);
    assign layer2_outputs[265] = layer1_outputs[2941];
    assign layer2_outputs[266] = (layer1_outputs[9233]) ^ (layer1_outputs[80]);
    assign layer2_outputs[267] = ~(layer1_outputs[7991]) | (layer1_outputs[1686]);
    assign layer2_outputs[268] = layer1_outputs[10357];
    assign layer2_outputs[269] = 1'b0;
    assign layer2_outputs[270] = (layer1_outputs[2457]) ^ (layer1_outputs[1121]);
    assign layer2_outputs[271] = ~((layer1_outputs[642]) & (layer1_outputs[10830]));
    assign layer2_outputs[272] = 1'b0;
    assign layer2_outputs[273] = layer1_outputs[8803];
    assign layer2_outputs[274] = layer1_outputs[2949];
    assign layer2_outputs[275] = (layer1_outputs[7125]) ^ (layer1_outputs[5268]);
    assign layer2_outputs[276] = ~(layer1_outputs[2705]);
    assign layer2_outputs[277] = layer1_outputs[5435];
    assign layer2_outputs[278] = layer1_outputs[12626];
    assign layer2_outputs[279] = layer1_outputs[3183];
    assign layer2_outputs[280] = ~((layer1_outputs[8615]) ^ (layer1_outputs[11856]));
    assign layer2_outputs[281] = (layer1_outputs[2292]) | (layer1_outputs[485]);
    assign layer2_outputs[282] = ~((layer1_outputs[1736]) ^ (layer1_outputs[4479]));
    assign layer2_outputs[283] = ~(layer1_outputs[7882]) | (layer1_outputs[12263]);
    assign layer2_outputs[284] = layer1_outputs[3223];
    assign layer2_outputs[285] = ~(layer1_outputs[2412]);
    assign layer2_outputs[286] = (layer1_outputs[4222]) & ~(layer1_outputs[9678]);
    assign layer2_outputs[287] = (layer1_outputs[12128]) | (layer1_outputs[1681]);
    assign layer2_outputs[288] = ~((layer1_outputs[11021]) ^ (layer1_outputs[11290]));
    assign layer2_outputs[289] = layer1_outputs[3123];
    assign layer2_outputs[290] = ~((layer1_outputs[7334]) ^ (layer1_outputs[4615]));
    assign layer2_outputs[291] = layer1_outputs[12591];
    assign layer2_outputs[292] = (layer1_outputs[5424]) & (layer1_outputs[4173]);
    assign layer2_outputs[293] = ~(layer1_outputs[6902]);
    assign layer2_outputs[294] = ~((layer1_outputs[8289]) ^ (layer1_outputs[7907]));
    assign layer2_outputs[295] = layer1_outputs[7460];
    assign layer2_outputs[296] = (layer1_outputs[2744]) & ~(layer1_outputs[3727]);
    assign layer2_outputs[297] = ~(layer1_outputs[10444]);
    assign layer2_outputs[298] = ~(layer1_outputs[3445]);
    assign layer2_outputs[299] = ~(layer1_outputs[3391]);
    assign layer2_outputs[300] = ~(layer1_outputs[5871]);
    assign layer2_outputs[301] = layer1_outputs[2783];
    assign layer2_outputs[302] = ~((layer1_outputs[1030]) ^ (layer1_outputs[10278]));
    assign layer2_outputs[303] = ~(layer1_outputs[3102]) | (layer1_outputs[27]);
    assign layer2_outputs[304] = ~(layer1_outputs[3115]);
    assign layer2_outputs[305] = ~(layer1_outputs[11245]);
    assign layer2_outputs[306] = ~(layer1_outputs[5691]) | (layer1_outputs[4851]);
    assign layer2_outputs[307] = ~(layer1_outputs[2754]);
    assign layer2_outputs[308] = ~((layer1_outputs[9833]) | (layer1_outputs[2]));
    assign layer2_outputs[309] = ~(layer1_outputs[7424]);
    assign layer2_outputs[310] = (layer1_outputs[10527]) | (layer1_outputs[11941]);
    assign layer2_outputs[311] = ~(layer1_outputs[3330]);
    assign layer2_outputs[312] = ~(layer1_outputs[7624]);
    assign layer2_outputs[313] = layer1_outputs[8322];
    assign layer2_outputs[314] = ~(layer1_outputs[8532]);
    assign layer2_outputs[315] = layer1_outputs[1390];
    assign layer2_outputs[316] = (layer1_outputs[8857]) & (layer1_outputs[5726]);
    assign layer2_outputs[317] = ~((layer1_outputs[3481]) & (layer1_outputs[10119]));
    assign layer2_outputs[318] = (layer1_outputs[8831]) ^ (layer1_outputs[7219]);
    assign layer2_outputs[319] = (layer1_outputs[10944]) & ~(layer1_outputs[11429]);
    assign layer2_outputs[320] = layer1_outputs[6969];
    assign layer2_outputs[321] = ~(layer1_outputs[6735]);
    assign layer2_outputs[322] = (layer1_outputs[2944]) | (layer1_outputs[4632]);
    assign layer2_outputs[323] = ~(layer1_outputs[3675]);
    assign layer2_outputs[324] = layer1_outputs[6514];
    assign layer2_outputs[325] = ~(layer1_outputs[1367]);
    assign layer2_outputs[326] = layer1_outputs[8727];
    assign layer2_outputs[327] = ~((layer1_outputs[1092]) & (layer1_outputs[10522]));
    assign layer2_outputs[328] = ~(layer1_outputs[1026]);
    assign layer2_outputs[329] = (layer1_outputs[6961]) ^ (layer1_outputs[2217]);
    assign layer2_outputs[330] = (layer1_outputs[10641]) & ~(layer1_outputs[2022]);
    assign layer2_outputs[331] = (layer1_outputs[6455]) & (layer1_outputs[10734]);
    assign layer2_outputs[332] = (layer1_outputs[9086]) & ~(layer1_outputs[1296]);
    assign layer2_outputs[333] = ~(layer1_outputs[8801]);
    assign layer2_outputs[334] = (layer1_outputs[4645]) & ~(layer1_outputs[10674]);
    assign layer2_outputs[335] = ~((layer1_outputs[9769]) ^ (layer1_outputs[11820]));
    assign layer2_outputs[336] = ~(layer1_outputs[5392]) | (layer1_outputs[5999]);
    assign layer2_outputs[337] = ~(layer1_outputs[10623]) | (layer1_outputs[11024]);
    assign layer2_outputs[338] = ~(layer1_outputs[280]) | (layer1_outputs[3785]);
    assign layer2_outputs[339] = ~(layer1_outputs[794]) | (layer1_outputs[7185]);
    assign layer2_outputs[340] = (layer1_outputs[1588]) ^ (layer1_outputs[8597]);
    assign layer2_outputs[341] = ~(layer1_outputs[10678]);
    assign layer2_outputs[342] = ~(layer1_outputs[6772]);
    assign layer2_outputs[343] = (layer1_outputs[5601]) & ~(layer1_outputs[8435]);
    assign layer2_outputs[344] = ~(layer1_outputs[10832]);
    assign layer2_outputs[345] = ~(layer1_outputs[4137]);
    assign layer2_outputs[346] = layer1_outputs[12690];
    assign layer2_outputs[347] = ~(layer1_outputs[7663]) | (layer1_outputs[11239]);
    assign layer2_outputs[348] = ~(layer1_outputs[12263]);
    assign layer2_outputs[349] = (layer1_outputs[11587]) & ~(layer1_outputs[3045]);
    assign layer2_outputs[350] = ~(layer1_outputs[3253]) | (layer1_outputs[7875]);
    assign layer2_outputs[351] = (layer1_outputs[10313]) ^ (layer1_outputs[7754]);
    assign layer2_outputs[352] = ~((layer1_outputs[6593]) ^ (layer1_outputs[1701]));
    assign layer2_outputs[353] = layer1_outputs[9066];
    assign layer2_outputs[354] = ~(layer1_outputs[8725]);
    assign layer2_outputs[355] = ~(layer1_outputs[5777]);
    assign layer2_outputs[356] = layer1_outputs[7771];
    assign layer2_outputs[357] = (layer1_outputs[11285]) & ~(layer1_outputs[7065]);
    assign layer2_outputs[358] = (layer1_outputs[11223]) ^ (layer1_outputs[11833]);
    assign layer2_outputs[359] = layer1_outputs[6039];
    assign layer2_outputs[360] = layer1_outputs[8451];
    assign layer2_outputs[361] = (layer1_outputs[6110]) | (layer1_outputs[4327]);
    assign layer2_outputs[362] = layer1_outputs[2451];
    assign layer2_outputs[363] = layer1_outputs[473];
    assign layer2_outputs[364] = layer1_outputs[6298];
    assign layer2_outputs[365] = layer1_outputs[5433];
    assign layer2_outputs[366] = ~((layer1_outputs[3882]) ^ (layer1_outputs[10539]));
    assign layer2_outputs[367] = layer1_outputs[5297];
    assign layer2_outputs[368] = layer1_outputs[2170];
    assign layer2_outputs[369] = (layer1_outputs[12460]) | (layer1_outputs[7840]);
    assign layer2_outputs[370] = (layer1_outputs[3603]) & ~(layer1_outputs[603]);
    assign layer2_outputs[371] = layer1_outputs[6359];
    assign layer2_outputs[372] = ~(layer1_outputs[12099]) | (layer1_outputs[8533]);
    assign layer2_outputs[373] = layer1_outputs[4677];
    assign layer2_outputs[374] = ~((layer1_outputs[2732]) | (layer1_outputs[10321]));
    assign layer2_outputs[375] = layer1_outputs[4319];
    assign layer2_outputs[376] = (layer1_outputs[2995]) | (layer1_outputs[3673]);
    assign layer2_outputs[377] = ~((layer1_outputs[6123]) | (layer1_outputs[5307]));
    assign layer2_outputs[378] = (layer1_outputs[4076]) & ~(layer1_outputs[1245]);
    assign layer2_outputs[379] = ~((layer1_outputs[9811]) ^ (layer1_outputs[8008]));
    assign layer2_outputs[380] = layer1_outputs[8314];
    assign layer2_outputs[381] = ~((layer1_outputs[6877]) | (layer1_outputs[2287]));
    assign layer2_outputs[382] = ~(layer1_outputs[11226]) | (layer1_outputs[1486]);
    assign layer2_outputs[383] = layer1_outputs[1463];
    assign layer2_outputs[384] = (layer1_outputs[11803]) | (layer1_outputs[1166]);
    assign layer2_outputs[385] = ~(layer1_outputs[12603]) | (layer1_outputs[6527]);
    assign layer2_outputs[386] = ~(layer1_outputs[6861]);
    assign layer2_outputs[387] = ~((layer1_outputs[10181]) ^ (layer1_outputs[9169]));
    assign layer2_outputs[388] = (layer1_outputs[11256]) ^ (layer1_outputs[4860]);
    assign layer2_outputs[389] = layer1_outputs[4911];
    assign layer2_outputs[390] = layer1_outputs[10400];
    assign layer2_outputs[391] = ~(layer1_outputs[8364]);
    assign layer2_outputs[392] = ~(layer1_outputs[11451]);
    assign layer2_outputs[393] = ~(layer1_outputs[9458]) | (layer1_outputs[6511]);
    assign layer2_outputs[394] = ~(layer1_outputs[5851]);
    assign layer2_outputs[395] = layer1_outputs[12283];
    assign layer2_outputs[396] = (layer1_outputs[5371]) | (layer1_outputs[5036]);
    assign layer2_outputs[397] = ~((layer1_outputs[922]) ^ (layer1_outputs[288]));
    assign layer2_outputs[398] = ~(layer1_outputs[5136]) | (layer1_outputs[1286]);
    assign layer2_outputs[399] = layer1_outputs[3203];
    assign layer2_outputs[400] = layer1_outputs[3543];
    assign layer2_outputs[401] = ~((layer1_outputs[2481]) & (layer1_outputs[6893]));
    assign layer2_outputs[402] = ~(layer1_outputs[10529]);
    assign layer2_outputs[403] = ~((layer1_outputs[2495]) & (layer1_outputs[1366]));
    assign layer2_outputs[404] = (layer1_outputs[7429]) & ~(layer1_outputs[7923]);
    assign layer2_outputs[405] = 1'b0;
    assign layer2_outputs[406] = layer1_outputs[3305];
    assign layer2_outputs[407] = (layer1_outputs[4666]) & (layer1_outputs[8413]);
    assign layer2_outputs[408] = (layer1_outputs[1426]) | (layer1_outputs[11549]);
    assign layer2_outputs[409] = (layer1_outputs[6512]) & ~(layer1_outputs[6546]);
    assign layer2_outputs[410] = (layer1_outputs[11471]) & (layer1_outputs[5567]);
    assign layer2_outputs[411] = layer1_outputs[9649];
    assign layer2_outputs[412] = (layer1_outputs[9063]) | (layer1_outputs[91]);
    assign layer2_outputs[413] = (layer1_outputs[2274]) | (layer1_outputs[7493]);
    assign layer2_outputs[414] = (layer1_outputs[3256]) | (layer1_outputs[5175]);
    assign layer2_outputs[415] = ~(layer1_outputs[745]);
    assign layer2_outputs[416] = (layer1_outputs[10850]) & ~(layer1_outputs[3]);
    assign layer2_outputs[417] = layer1_outputs[6191];
    assign layer2_outputs[418] = ~(layer1_outputs[3537]);
    assign layer2_outputs[419] = ~((layer1_outputs[9272]) & (layer1_outputs[9522]));
    assign layer2_outputs[420] = ~((layer1_outputs[3614]) & (layer1_outputs[4775]));
    assign layer2_outputs[421] = ~(layer1_outputs[8309]);
    assign layer2_outputs[422] = (layer1_outputs[9284]) & (layer1_outputs[4165]);
    assign layer2_outputs[423] = (layer1_outputs[10531]) & (layer1_outputs[6224]);
    assign layer2_outputs[424] = layer1_outputs[9939];
    assign layer2_outputs[425] = layer1_outputs[6160];
    assign layer2_outputs[426] = layer1_outputs[7047];
    assign layer2_outputs[427] = (layer1_outputs[3506]) ^ (layer1_outputs[4212]);
    assign layer2_outputs[428] = ~((layer1_outputs[4491]) | (layer1_outputs[5397]));
    assign layer2_outputs[429] = layer1_outputs[1373];
    assign layer2_outputs[430] = (layer1_outputs[1658]) ^ (layer1_outputs[10123]);
    assign layer2_outputs[431] = layer1_outputs[7223];
    assign layer2_outputs[432] = layer1_outputs[11627];
    assign layer2_outputs[433] = ~(layer1_outputs[2919]) | (layer1_outputs[6426]);
    assign layer2_outputs[434] = layer1_outputs[3854];
    assign layer2_outputs[435] = layer1_outputs[6757];
    assign layer2_outputs[436] = ~(layer1_outputs[12047]);
    assign layer2_outputs[437] = layer1_outputs[8139];
    assign layer2_outputs[438] = layer1_outputs[4319];
    assign layer2_outputs[439] = layer1_outputs[8569];
    assign layer2_outputs[440] = ~(layer1_outputs[7757]);
    assign layer2_outputs[441] = 1'b1;
    assign layer2_outputs[442] = (layer1_outputs[5715]) & ~(layer1_outputs[11250]);
    assign layer2_outputs[443] = ~(layer1_outputs[3763]) | (layer1_outputs[10569]);
    assign layer2_outputs[444] = (layer1_outputs[4665]) & ~(layer1_outputs[1528]);
    assign layer2_outputs[445] = (layer1_outputs[7488]) & ~(layer1_outputs[376]);
    assign layer2_outputs[446] = ~((layer1_outputs[4793]) | (layer1_outputs[4416]));
    assign layer2_outputs[447] = layer1_outputs[11677];
    assign layer2_outputs[448] = (layer1_outputs[7815]) & ~(layer1_outputs[7774]);
    assign layer2_outputs[449] = ~((layer1_outputs[5473]) & (layer1_outputs[11383]));
    assign layer2_outputs[450] = ~(layer1_outputs[11512]);
    assign layer2_outputs[451] = (layer1_outputs[10285]) & (layer1_outputs[4848]);
    assign layer2_outputs[452] = layer1_outputs[9052];
    assign layer2_outputs[453] = ~((layer1_outputs[8060]) ^ (layer1_outputs[5257]));
    assign layer2_outputs[454] = ~(layer1_outputs[10978]);
    assign layer2_outputs[455] = ~(layer1_outputs[10463]);
    assign layer2_outputs[456] = ~(layer1_outputs[6167]) | (layer1_outputs[7027]);
    assign layer2_outputs[457] = ~((layer1_outputs[903]) ^ (layer1_outputs[5932]));
    assign layer2_outputs[458] = ~((layer1_outputs[10048]) ^ (layer1_outputs[5672]));
    assign layer2_outputs[459] = (layer1_outputs[6558]) & ~(layer1_outputs[9847]);
    assign layer2_outputs[460] = ~(layer1_outputs[7453]);
    assign layer2_outputs[461] = ~(layer1_outputs[12391]);
    assign layer2_outputs[462] = layer1_outputs[2745];
    assign layer2_outputs[463] = (layer1_outputs[10901]) & ~(layer1_outputs[10445]);
    assign layer2_outputs[464] = layer1_outputs[10638];
    assign layer2_outputs[465] = ~(layer1_outputs[3576]) | (layer1_outputs[12138]);
    assign layer2_outputs[466] = ~(layer1_outputs[11681]);
    assign layer2_outputs[467] = ~((layer1_outputs[12433]) ^ (layer1_outputs[4579]));
    assign layer2_outputs[468] = ~((layer1_outputs[6257]) | (layer1_outputs[7912]));
    assign layer2_outputs[469] = ~((layer1_outputs[10187]) & (layer1_outputs[4810]));
    assign layer2_outputs[470] = ~(layer1_outputs[8763]) | (layer1_outputs[10635]);
    assign layer2_outputs[471] = ~((layer1_outputs[233]) ^ (layer1_outputs[382]));
    assign layer2_outputs[472] = ~(layer1_outputs[3961]);
    assign layer2_outputs[473] = ~(layer1_outputs[10437]);
    assign layer2_outputs[474] = ~(layer1_outputs[2256]);
    assign layer2_outputs[475] = ~(layer1_outputs[473]);
    assign layer2_outputs[476] = layer1_outputs[1379];
    assign layer2_outputs[477] = ~(layer1_outputs[9350]) | (layer1_outputs[4489]);
    assign layer2_outputs[478] = (layer1_outputs[6287]) & ~(layer1_outputs[9876]);
    assign layer2_outputs[479] = 1'b0;
    assign layer2_outputs[480] = ~(layer1_outputs[11362]);
    assign layer2_outputs[481] = layer1_outputs[4847];
    assign layer2_outputs[482] = (layer1_outputs[7484]) ^ (layer1_outputs[8534]);
    assign layer2_outputs[483] = layer1_outputs[9562];
    assign layer2_outputs[484] = ~((layer1_outputs[9513]) ^ (layer1_outputs[728]));
    assign layer2_outputs[485] = layer1_outputs[3352];
    assign layer2_outputs[486] = ~(layer1_outputs[3757]);
    assign layer2_outputs[487] = ~(layer1_outputs[7976]);
    assign layer2_outputs[488] = ~((layer1_outputs[4120]) | (layer1_outputs[10768]));
    assign layer2_outputs[489] = ~(layer1_outputs[2476]) | (layer1_outputs[1538]);
    assign layer2_outputs[490] = ~((layer1_outputs[1431]) | (layer1_outputs[7721]));
    assign layer2_outputs[491] = (layer1_outputs[7143]) & (layer1_outputs[996]);
    assign layer2_outputs[492] = ~((layer1_outputs[9625]) & (layer1_outputs[5611]));
    assign layer2_outputs[493] = ~(layer1_outputs[11533]);
    assign layer2_outputs[494] = ~(layer1_outputs[10984]) | (layer1_outputs[3508]);
    assign layer2_outputs[495] = ~(layer1_outputs[3981]);
    assign layer2_outputs[496] = ~(layer1_outputs[8387]);
    assign layer2_outputs[497] = ~(layer1_outputs[4774]) | (layer1_outputs[10792]);
    assign layer2_outputs[498] = 1'b1;
    assign layer2_outputs[499] = ~((layer1_outputs[3831]) ^ (layer1_outputs[7805]));
    assign layer2_outputs[500] = (layer1_outputs[8108]) & ~(layer1_outputs[1816]);
    assign layer2_outputs[501] = layer1_outputs[10962];
    assign layer2_outputs[502] = (layer1_outputs[9192]) & ~(layer1_outputs[6089]);
    assign layer2_outputs[503] = layer1_outputs[12303];
    assign layer2_outputs[504] = (layer1_outputs[4332]) & (layer1_outputs[8952]);
    assign layer2_outputs[505] = layer1_outputs[10961];
    assign layer2_outputs[506] = (layer1_outputs[2510]) & ~(layer1_outputs[1679]);
    assign layer2_outputs[507] = ~((layer1_outputs[3925]) ^ (layer1_outputs[100]));
    assign layer2_outputs[508] = ~((layer1_outputs[730]) | (layer1_outputs[9572]));
    assign layer2_outputs[509] = ~(layer1_outputs[91]);
    assign layer2_outputs[510] = (layer1_outputs[11482]) ^ (layer1_outputs[9709]);
    assign layer2_outputs[511] = ~((layer1_outputs[987]) & (layer1_outputs[12330]));
    assign layer2_outputs[512] = (layer1_outputs[9073]) ^ (layer1_outputs[8189]);
    assign layer2_outputs[513] = (layer1_outputs[12603]) & (layer1_outputs[11930]);
    assign layer2_outputs[514] = ~((layer1_outputs[10627]) ^ (layer1_outputs[2707]));
    assign layer2_outputs[515] = 1'b0;
    assign layer2_outputs[516] = ~(layer1_outputs[2677]) | (layer1_outputs[7294]);
    assign layer2_outputs[517] = layer1_outputs[12762];
    assign layer2_outputs[518] = layer1_outputs[6998];
    assign layer2_outputs[519] = (layer1_outputs[4182]) & ~(layer1_outputs[10089]);
    assign layer2_outputs[520] = layer1_outputs[11140];
    assign layer2_outputs[521] = (layer1_outputs[7261]) ^ (layer1_outputs[1573]);
    assign layer2_outputs[522] = (layer1_outputs[6078]) ^ (layer1_outputs[8799]);
    assign layer2_outputs[523] = ~((layer1_outputs[4924]) & (layer1_outputs[11673]));
    assign layer2_outputs[524] = ~(layer1_outputs[8222]);
    assign layer2_outputs[525] = ~(layer1_outputs[7502]);
    assign layer2_outputs[526] = ~((layer1_outputs[4275]) ^ (layer1_outputs[2822]));
    assign layer2_outputs[527] = layer1_outputs[9622];
    assign layer2_outputs[528] = (layer1_outputs[10717]) | (layer1_outputs[5148]);
    assign layer2_outputs[529] = ~(layer1_outputs[5007]) | (layer1_outputs[5476]);
    assign layer2_outputs[530] = ~(layer1_outputs[4024]);
    assign layer2_outputs[531] = ~(layer1_outputs[12298]) | (layer1_outputs[1560]);
    assign layer2_outputs[532] = layer1_outputs[9328];
    assign layer2_outputs[533] = layer1_outputs[10320];
    assign layer2_outputs[534] = (layer1_outputs[12609]) | (layer1_outputs[8665]);
    assign layer2_outputs[535] = ~(layer1_outputs[9834]);
    assign layer2_outputs[536] = (layer1_outputs[5009]) ^ (layer1_outputs[876]);
    assign layer2_outputs[537] = ~((layer1_outputs[10059]) & (layer1_outputs[933]));
    assign layer2_outputs[538] = layer1_outputs[2440];
    assign layer2_outputs[539] = (layer1_outputs[10348]) | (layer1_outputs[9260]);
    assign layer2_outputs[540] = layer1_outputs[1667];
    assign layer2_outputs[541] = (layer1_outputs[11008]) & ~(layer1_outputs[947]);
    assign layer2_outputs[542] = layer1_outputs[9259];
    assign layer2_outputs[543] = (layer1_outputs[8867]) | (layer1_outputs[12310]);
    assign layer2_outputs[544] = ~((layer1_outputs[10775]) | (layer1_outputs[1270]));
    assign layer2_outputs[545] = (layer1_outputs[10513]) & (layer1_outputs[11918]);
    assign layer2_outputs[546] = layer1_outputs[7377];
    assign layer2_outputs[547] = (layer1_outputs[3306]) & ~(layer1_outputs[8808]);
    assign layer2_outputs[548] = ~(layer1_outputs[1962]);
    assign layer2_outputs[549] = (layer1_outputs[7642]) ^ (layer1_outputs[5539]);
    assign layer2_outputs[550] = ~((layer1_outputs[10518]) ^ (layer1_outputs[6156]));
    assign layer2_outputs[551] = ~(layer1_outputs[7004]);
    assign layer2_outputs[552] = ~(layer1_outputs[2992]);
    assign layer2_outputs[553] = ~(layer1_outputs[10322]);
    assign layer2_outputs[554] = (layer1_outputs[9843]) & (layer1_outputs[12090]);
    assign layer2_outputs[555] = ~(layer1_outputs[12158]);
    assign layer2_outputs[556] = ~(layer1_outputs[5974]);
    assign layer2_outputs[557] = (layer1_outputs[7470]) & (layer1_outputs[8411]);
    assign layer2_outputs[558] = ~(layer1_outputs[4139]);
    assign layer2_outputs[559] = ~((layer1_outputs[12375]) ^ (layer1_outputs[6747]));
    assign layer2_outputs[560] = layer1_outputs[5261];
    assign layer2_outputs[561] = ~(layer1_outputs[8930]);
    assign layer2_outputs[562] = ~((layer1_outputs[8279]) | (layer1_outputs[2865]));
    assign layer2_outputs[563] = layer1_outputs[7594];
    assign layer2_outputs[564] = (layer1_outputs[11933]) & (layer1_outputs[9679]);
    assign layer2_outputs[565] = ~(layer1_outputs[11660]);
    assign layer2_outputs[566] = layer1_outputs[12365];
    assign layer2_outputs[567] = ~(layer1_outputs[4772]);
    assign layer2_outputs[568] = layer1_outputs[5409];
    assign layer2_outputs[569] = (layer1_outputs[10102]) ^ (layer1_outputs[9583]);
    assign layer2_outputs[570] = (layer1_outputs[5773]) | (layer1_outputs[8506]);
    assign layer2_outputs[571] = ~((layer1_outputs[7521]) ^ (layer1_outputs[5511]));
    assign layer2_outputs[572] = layer1_outputs[4090];
    assign layer2_outputs[573] = ~(layer1_outputs[8462]);
    assign layer2_outputs[574] = ~(layer1_outputs[665]);
    assign layer2_outputs[575] = ~((layer1_outputs[3547]) | (layer1_outputs[7288]));
    assign layer2_outputs[576] = (layer1_outputs[8040]) | (layer1_outputs[12505]);
    assign layer2_outputs[577] = ~(layer1_outputs[2864]);
    assign layer2_outputs[578] = ~(layer1_outputs[347]);
    assign layer2_outputs[579] = layer1_outputs[6491];
    assign layer2_outputs[580] = ~((layer1_outputs[2712]) | (layer1_outputs[2626]));
    assign layer2_outputs[581] = (layer1_outputs[12547]) ^ (layer1_outputs[2209]);
    assign layer2_outputs[582] = layer1_outputs[9756];
    assign layer2_outputs[583] = (layer1_outputs[5991]) & ~(layer1_outputs[6799]);
    assign layer2_outputs[584] = (layer1_outputs[3451]) | (layer1_outputs[11434]);
    assign layer2_outputs[585] = layer1_outputs[5684];
    assign layer2_outputs[586] = layer1_outputs[7889];
    assign layer2_outputs[587] = ~(layer1_outputs[1908]);
    assign layer2_outputs[588] = ~(layer1_outputs[10492]) | (layer1_outputs[527]);
    assign layer2_outputs[589] = ~(layer1_outputs[5990]);
    assign layer2_outputs[590] = ~(layer1_outputs[5456]);
    assign layer2_outputs[591] = (layer1_outputs[472]) ^ (layer1_outputs[2784]);
    assign layer2_outputs[592] = (layer1_outputs[1469]) & (layer1_outputs[3993]);
    assign layer2_outputs[593] = (layer1_outputs[8957]) & (layer1_outputs[1640]);
    assign layer2_outputs[594] = ~(layer1_outputs[10280]);
    assign layer2_outputs[595] = ~(layer1_outputs[5234]);
    assign layer2_outputs[596] = layer1_outputs[2998];
    assign layer2_outputs[597] = layer1_outputs[3332];
    assign layer2_outputs[598] = layer1_outputs[10967];
    assign layer2_outputs[599] = layer1_outputs[10267];
    assign layer2_outputs[600] = layer1_outputs[1089];
    assign layer2_outputs[601] = layer1_outputs[4637];
    assign layer2_outputs[602] = (layer1_outputs[12739]) ^ (layer1_outputs[2413]);
    assign layer2_outputs[603] = (layer1_outputs[6130]) & ~(layer1_outputs[4180]);
    assign layer2_outputs[604] = layer1_outputs[6896];
    assign layer2_outputs[605] = layer1_outputs[530];
    assign layer2_outputs[606] = ~(layer1_outputs[3840]);
    assign layer2_outputs[607] = ~(layer1_outputs[4250]);
    assign layer2_outputs[608] = ~(layer1_outputs[6196]);
    assign layer2_outputs[609] = (layer1_outputs[3606]) | (layer1_outputs[6625]);
    assign layer2_outputs[610] = (layer1_outputs[9373]) ^ (layer1_outputs[4904]);
    assign layer2_outputs[611] = (layer1_outputs[9699]) & ~(layer1_outputs[1947]);
    assign layer2_outputs[612] = ~(layer1_outputs[5573]) | (layer1_outputs[10504]);
    assign layer2_outputs[613] = ~(layer1_outputs[12779]) | (layer1_outputs[1225]);
    assign layer2_outputs[614] = layer1_outputs[6714];
    assign layer2_outputs[615] = layer1_outputs[481];
    assign layer2_outputs[616] = (layer1_outputs[11989]) ^ (layer1_outputs[11771]);
    assign layer2_outputs[617] = layer1_outputs[10776];
    assign layer2_outputs[618] = ~(layer1_outputs[2397]);
    assign layer2_outputs[619] = (layer1_outputs[4057]) | (layer1_outputs[11102]);
    assign layer2_outputs[620] = (layer1_outputs[2363]) ^ (layer1_outputs[3385]);
    assign layer2_outputs[621] = (layer1_outputs[4357]) ^ (layer1_outputs[9275]);
    assign layer2_outputs[622] = ~(layer1_outputs[6541]) | (layer1_outputs[11233]);
    assign layer2_outputs[623] = ~((layer1_outputs[6813]) | (layer1_outputs[12754]));
    assign layer2_outputs[624] = ~(layer1_outputs[12718]);
    assign layer2_outputs[625] = ~(layer1_outputs[10704]) | (layer1_outputs[11216]);
    assign layer2_outputs[626] = (layer1_outputs[2706]) & (layer1_outputs[10126]);
    assign layer2_outputs[627] = layer1_outputs[2039];
    assign layer2_outputs[628] = ~(layer1_outputs[3500]);
    assign layer2_outputs[629] = ~(layer1_outputs[1173]);
    assign layer2_outputs[630] = ~(layer1_outputs[10688]);
    assign layer2_outputs[631] = (layer1_outputs[3918]) ^ (layer1_outputs[11278]);
    assign layer2_outputs[632] = 1'b1;
    assign layer2_outputs[633] = ~(layer1_outputs[2077]);
    assign layer2_outputs[634] = ~(layer1_outputs[1708]);
    assign layer2_outputs[635] = ~(layer1_outputs[4148]);
    assign layer2_outputs[636] = layer1_outputs[5606];
    assign layer2_outputs[637] = ~(layer1_outputs[12328]) | (layer1_outputs[8137]);
    assign layer2_outputs[638] = layer1_outputs[5396];
    assign layer2_outputs[639] = (layer1_outputs[11110]) & ~(layer1_outputs[3668]);
    assign layer2_outputs[640] = layer1_outputs[4510];
    assign layer2_outputs[641] = ~((layer1_outputs[861]) | (layer1_outputs[10904]));
    assign layer2_outputs[642] = layer1_outputs[6737];
    assign layer2_outputs[643] = layer1_outputs[4680];
    assign layer2_outputs[644] = ~(layer1_outputs[4433]);
    assign layer2_outputs[645] = ~((layer1_outputs[10049]) ^ (layer1_outputs[11444]));
    assign layer2_outputs[646] = ~(layer1_outputs[5127]);
    assign layer2_outputs[647] = ~(layer1_outputs[12314]) | (layer1_outputs[2592]);
    assign layer2_outputs[648] = (layer1_outputs[5809]) & (layer1_outputs[9316]);
    assign layer2_outputs[649] = ~(layer1_outputs[12778]);
    assign layer2_outputs[650] = ~(layer1_outputs[4405]);
    assign layer2_outputs[651] = layer1_outputs[8329];
    assign layer2_outputs[652] = (layer1_outputs[5523]) & (layer1_outputs[9877]);
    assign layer2_outputs[653] = (layer1_outputs[3106]) & ~(layer1_outputs[9452]);
    assign layer2_outputs[654] = ~(layer1_outputs[7977]) | (layer1_outputs[2400]);
    assign layer2_outputs[655] = layer1_outputs[11583];
    assign layer2_outputs[656] = ~(layer1_outputs[4011]);
    assign layer2_outputs[657] = ~(layer1_outputs[6952]);
    assign layer2_outputs[658] = (layer1_outputs[7315]) & (layer1_outputs[5254]);
    assign layer2_outputs[659] = ~((layer1_outputs[9069]) & (layer1_outputs[5254]));
    assign layer2_outputs[660] = ~(layer1_outputs[3059]);
    assign layer2_outputs[661] = (layer1_outputs[10940]) & ~(layer1_outputs[4402]);
    assign layer2_outputs[662] = ~(layer1_outputs[11469]) | (layer1_outputs[3850]);
    assign layer2_outputs[663] = layer1_outputs[4516];
    assign layer2_outputs[664] = ~(layer1_outputs[9154]);
    assign layer2_outputs[665] = ~(layer1_outputs[2279]);
    assign layer2_outputs[666] = ~((layer1_outputs[4440]) ^ (layer1_outputs[5954]));
    assign layer2_outputs[667] = layer1_outputs[748];
    assign layer2_outputs[668] = (layer1_outputs[3442]) | (layer1_outputs[3188]);
    assign layer2_outputs[669] = (layer1_outputs[6181]) & ~(layer1_outputs[7968]);
    assign layer2_outputs[670] = ~((layer1_outputs[4884]) | (layer1_outputs[6904]));
    assign layer2_outputs[671] = ~((layer1_outputs[8709]) ^ (layer1_outputs[42]));
    assign layer2_outputs[672] = (layer1_outputs[10158]) & (layer1_outputs[667]);
    assign layer2_outputs[673] = layer1_outputs[6850];
    assign layer2_outputs[674] = ~((layer1_outputs[12495]) | (layer1_outputs[4473]));
    assign layer2_outputs[675] = layer1_outputs[11643];
    assign layer2_outputs[676] = ~(layer1_outputs[10433]);
    assign layer2_outputs[677] = (layer1_outputs[11810]) & ~(layer1_outputs[8165]);
    assign layer2_outputs[678] = ~((layer1_outputs[4158]) & (layer1_outputs[12510]));
    assign layer2_outputs[679] = ~(layer1_outputs[4604]) | (layer1_outputs[2161]);
    assign layer2_outputs[680] = ~((layer1_outputs[9981]) & (layer1_outputs[8637]));
    assign layer2_outputs[681] = ~(layer1_outputs[2175]) | (layer1_outputs[11957]);
    assign layer2_outputs[682] = layer1_outputs[6872];
    assign layer2_outputs[683] = ~((layer1_outputs[1682]) | (layer1_outputs[3650]));
    assign layer2_outputs[684] = (layer1_outputs[5745]) & ~(layer1_outputs[4597]);
    assign layer2_outputs[685] = ~(layer1_outputs[10095]);
    assign layer2_outputs[686] = ~(layer1_outputs[8945]);
    assign layer2_outputs[687] = layer1_outputs[4226];
    assign layer2_outputs[688] = (layer1_outputs[5496]) | (layer1_outputs[3727]);
    assign layer2_outputs[689] = ~(layer1_outputs[7616]) | (layer1_outputs[668]);
    assign layer2_outputs[690] = ~(layer1_outputs[4516]);
    assign layer2_outputs[691] = (layer1_outputs[11558]) & ~(layer1_outputs[11003]);
    assign layer2_outputs[692] = ~((layer1_outputs[948]) & (layer1_outputs[6233]));
    assign layer2_outputs[693] = ~(layer1_outputs[9724]);
    assign layer2_outputs[694] = layer1_outputs[2332];
    assign layer2_outputs[695] = layer1_outputs[5575];
    assign layer2_outputs[696] = layer1_outputs[4123];
    assign layer2_outputs[697] = ~(layer1_outputs[6449]) | (layer1_outputs[3894]);
    assign layer2_outputs[698] = ~((layer1_outputs[12193]) ^ (layer1_outputs[4871]));
    assign layer2_outputs[699] = ~(layer1_outputs[6341]);
    assign layer2_outputs[700] = layer1_outputs[6251];
    assign layer2_outputs[701] = ~((layer1_outputs[7657]) | (layer1_outputs[1076]));
    assign layer2_outputs[702] = ~(layer1_outputs[9772]) | (layer1_outputs[6666]);
    assign layer2_outputs[703] = (layer1_outputs[1282]) ^ (layer1_outputs[6727]);
    assign layer2_outputs[704] = layer1_outputs[9474];
    assign layer2_outputs[705] = (layer1_outputs[10315]) ^ (layer1_outputs[8505]);
    assign layer2_outputs[706] = ~((layer1_outputs[3760]) ^ (layer1_outputs[9567]));
    assign layer2_outputs[707] = 1'b0;
    assign layer2_outputs[708] = layer1_outputs[1074];
    assign layer2_outputs[709] = ~(layer1_outputs[12600]);
    assign layer2_outputs[710] = ~(layer1_outputs[11575]);
    assign layer2_outputs[711] = ~(layer1_outputs[771]);
    assign layer2_outputs[712] = layer1_outputs[4865];
    assign layer2_outputs[713] = (layer1_outputs[7974]) ^ (layer1_outputs[9345]);
    assign layer2_outputs[714] = (layer1_outputs[9932]) | (layer1_outputs[7398]);
    assign layer2_outputs[715] = layer1_outputs[8859];
    assign layer2_outputs[716] = ~((layer1_outputs[3826]) & (layer1_outputs[5674]));
    assign layer2_outputs[717] = (layer1_outputs[12095]) & (layer1_outputs[3052]);
    assign layer2_outputs[718] = ~((layer1_outputs[11881]) & (layer1_outputs[7791]));
    assign layer2_outputs[719] = (layer1_outputs[5902]) & (layer1_outputs[5010]);
    assign layer2_outputs[720] = (layer1_outputs[9013]) | (layer1_outputs[11664]);
    assign layer2_outputs[721] = layer1_outputs[9158];
    assign layer2_outputs[722] = layer1_outputs[1146];
    assign layer2_outputs[723] = layer1_outputs[6366];
    assign layer2_outputs[724] = (layer1_outputs[6595]) ^ (layer1_outputs[2093]);
    assign layer2_outputs[725] = (layer1_outputs[3929]) & ~(layer1_outputs[7882]);
    assign layer2_outputs[726] = (layer1_outputs[8623]) & (layer1_outputs[8093]);
    assign layer2_outputs[727] = layer1_outputs[6915];
    assign layer2_outputs[728] = ~(layer1_outputs[11590]);
    assign layer2_outputs[729] = 1'b0;
    assign layer2_outputs[730] = (layer1_outputs[2491]) & (layer1_outputs[477]);
    assign layer2_outputs[731] = ~(layer1_outputs[2717]) | (layer1_outputs[1014]);
    assign layer2_outputs[732] = ~(layer1_outputs[1764]) | (layer1_outputs[232]);
    assign layer2_outputs[733] = ~(layer1_outputs[3878]);
    assign layer2_outputs[734] = ~(layer1_outputs[2399]);
    assign layer2_outputs[735] = (layer1_outputs[1142]) ^ (layer1_outputs[7750]);
    assign layer2_outputs[736] = (layer1_outputs[1763]) ^ (layer1_outputs[8949]);
    assign layer2_outputs[737] = ~(layer1_outputs[3903]);
    assign layer2_outputs[738] = (layer1_outputs[1828]) & ~(layer1_outputs[12731]);
    assign layer2_outputs[739] = layer1_outputs[7999];
    assign layer2_outputs[740] = (layer1_outputs[2465]) & (layer1_outputs[5420]);
    assign layer2_outputs[741] = layer1_outputs[3050];
    assign layer2_outputs[742] = ~((layer1_outputs[5351]) & (layer1_outputs[2572]));
    assign layer2_outputs[743] = ~(layer1_outputs[3533]);
    assign layer2_outputs[744] = layer1_outputs[1782];
    assign layer2_outputs[745] = layer1_outputs[6949];
    assign layer2_outputs[746] = ~(layer1_outputs[1182]) | (layer1_outputs[6494]);
    assign layer2_outputs[747] = ~((layer1_outputs[37]) ^ (layer1_outputs[7287]));
    assign layer2_outputs[748] = ~(layer1_outputs[8367]) | (layer1_outputs[6203]);
    assign layer2_outputs[749] = ~((layer1_outputs[11867]) & (layer1_outputs[3844]));
    assign layer2_outputs[750] = (layer1_outputs[6346]) | (layer1_outputs[8547]);
    assign layer2_outputs[751] = ~(layer1_outputs[1996]);
    assign layer2_outputs[752] = ~(layer1_outputs[9449]);
    assign layer2_outputs[753] = (layer1_outputs[12675]) | (layer1_outputs[4916]);
    assign layer2_outputs[754] = ~(layer1_outputs[1287]) | (layer1_outputs[703]);
    assign layer2_outputs[755] = ~(layer1_outputs[566]) | (layer1_outputs[8452]);
    assign layer2_outputs[756] = layer1_outputs[488];
    assign layer2_outputs[757] = ~(layer1_outputs[12615]) | (layer1_outputs[10816]);
    assign layer2_outputs[758] = (layer1_outputs[9753]) ^ (layer1_outputs[9049]);
    assign layer2_outputs[759] = layer1_outputs[487];
    assign layer2_outputs[760] = ~((layer1_outputs[8051]) | (layer1_outputs[10824]));
    assign layer2_outputs[761] = ~((layer1_outputs[6863]) ^ (layer1_outputs[4650]));
    assign layer2_outputs[762] = layer1_outputs[1866];
    assign layer2_outputs[763] = ~((layer1_outputs[5055]) | (layer1_outputs[3755]));
    assign layer2_outputs[764] = ~(layer1_outputs[757]);
    assign layer2_outputs[765] = ~(layer1_outputs[2330]) | (layer1_outputs[12098]);
    assign layer2_outputs[766] = (layer1_outputs[6031]) | (layer1_outputs[11758]);
    assign layer2_outputs[767] = ~((layer1_outputs[10722]) & (layer1_outputs[10985]));
    assign layer2_outputs[768] = layer1_outputs[1249];
    assign layer2_outputs[769] = ~((layer1_outputs[124]) & (layer1_outputs[3181]));
    assign layer2_outputs[770] = ~(layer1_outputs[2641]) | (layer1_outputs[1846]);
    assign layer2_outputs[771] = 1'b0;
    assign layer2_outputs[772] = layer1_outputs[7918];
    assign layer2_outputs[773] = ~(layer1_outputs[413]);
    assign layer2_outputs[774] = ~((layer1_outputs[3697]) | (layer1_outputs[365]));
    assign layer2_outputs[775] = ~(layer1_outputs[4497]);
    assign layer2_outputs[776] = (layer1_outputs[2543]) ^ (layer1_outputs[7894]);
    assign layer2_outputs[777] = layer1_outputs[10726];
    assign layer2_outputs[778] = layer1_outputs[1900];
    assign layer2_outputs[779] = (layer1_outputs[2532]) ^ (layer1_outputs[110]);
    assign layer2_outputs[780] = ~((layer1_outputs[2838]) & (layer1_outputs[2873]));
    assign layer2_outputs[781] = ~(layer1_outputs[46]) | (layer1_outputs[4331]);
    assign layer2_outputs[782] = (layer1_outputs[10532]) & ~(layer1_outputs[8994]);
    assign layer2_outputs[783] = layer1_outputs[2253];
    assign layer2_outputs[784] = ~(layer1_outputs[9633]);
    assign layer2_outputs[785] = (layer1_outputs[5073]) & (layer1_outputs[12273]);
    assign layer2_outputs[786] = layer1_outputs[9620];
    assign layer2_outputs[787] = layer1_outputs[4972];
    assign layer2_outputs[788] = layer1_outputs[8814];
    assign layer2_outputs[789] = ~(layer1_outputs[2530]) | (layer1_outputs[1049]);
    assign layer2_outputs[790] = layer1_outputs[303];
    assign layer2_outputs[791] = ~(layer1_outputs[11643]);
    assign layer2_outputs[792] = (layer1_outputs[9807]) & ~(layer1_outputs[2321]);
    assign layer2_outputs[793] = (layer1_outputs[11266]) ^ (layer1_outputs[958]);
    assign layer2_outputs[794] = ~((layer1_outputs[7970]) & (layer1_outputs[1296]));
    assign layer2_outputs[795] = layer1_outputs[11001];
    assign layer2_outputs[796] = (layer1_outputs[4262]) & ~(layer1_outputs[11650]);
    assign layer2_outputs[797] = ~((layer1_outputs[11766]) ^ (layer1_outputs[145]));
    assign layer2_outputs[798] = ~((layer1_outputs[5978]) ^ (layer1_outputs[10926]));
    assign layer2_outputs[799] = (layer1_outputs[9882]) ^ (layer1_outputs[6510]);
    assign layer2_outputs[800] = ~(layer1_outputs[8075]);
    assign layer2_outputs[801] = ~(layer1_outputs[8645]);
    assign layer2_outputs[802] = 1'b1;
    assign layer2_outputs[803] = ~((layer1_outputs[9642]) & (layer1_outputs[4131]));
    assign layer2_outputs[804] = layer1_outputs[10638];
    assign layer2_outputs[805] = ~((layer1_outputs[12796]) ^ (layer1_outputs[8980]));
    assign layer2_outputs[806] = ~((layer1_outputs[5377]) ^ (layer1_outputs[10869]));
    assign layer2_outputs[807] = ~((layer1_outputs[6974]) & (layer1_outputs[760]));
    assign layer2_outputs[808] = ~(layer1_outputs[3568]);
    assign layer2_outputs[809] = layer1_outputs[11031];
    assign layer2_outputs[810] = ~(layer1_outputs[3685]);
    assign layer2_outputs[811] = (layer1_outputs[9320]) | (layer1_outputs[3340]);
    assign layer2_outputs[812] = layer1_outputs[6051];
    assign layer2_outputs[813] = ~(layer1_outputs[9161]) | (layer1_outputs[6623]);
    assign layer2_outputs[814] = (layer1_outputs[1688]) & ~(layer1_outputs[1764]);
    assign layer2_outputs[815] = ~((layer1_outputs[2634]) ^ (layer1_outputs[7197]));
    assign layer2_outputs[816] = layer1_outputs[5790];
    assign layer2_outputs[817] = ~(layer1_outputs[8991]);
    assign layer2_outputs[818] = ~((layer1_outputs[1246]) ^ (layer1_outputs[4077]));
    assign layer2_outputs[819] = ~((layer1_outputs[10992]) | (layer1_outputs[12518]));
    assign layer2_outputs[820] = (layer1_outputs[6241]) & ~(layer1_outputs[1317]);
    assign layer2_outputs[821] = ~((layer1_outputs[8931]) ^ (layer1_outputs[11900]));
    assign layer2_outputs[822] = layer1_outputs[784];
    assign layer2_outputs[823] = ~(layer1_outputs[7265]) | (layer1_outputs[3257]);
    assign layer2_outputs[824] = layer1_outputs[1699];
    assign layer2_outputs[825] = ~(layer1_outputs[2580]) | (layer1_outputs[3014]);
    assign layer2_outputs[826] = (layer1_outputs[3274]) ^ (layer1_outputs[2281]);
    assign layer2_outputs[827] = ~(layer1_outputs[11366]) | (layer1_outputs[8029]);
    assign layer2_outputs[828] = layer1_outputs[7554];
    assign layer2_outputs[829] = layer1_outputs[7680];
    assign layer2_outputs[830] = (layer1_outputs[10566]) & ~(layer1_outputs[4055]);
    assign layer2_outputs[831] = ~(layer1_outputs[4632]) | (layer1_outputs[1632]);
    assign layer2_outputs[832] = (layer1_outputs[1050]) & ~(layer1_outputs[8389]);
    assign layer2_outputs[833] = ~((layer1_outputs[2541]) | (layer1_outputs[6047]));
    assign layer2_outputs[834] = 1'b1;
    assign layer2_outputs[835] = layer1_outputs[7011];
    assign layer2_outputs[836] = ~(layer1_outputs[1061]);
    assign layer2_outputs[837] = layer1_outputs[11730];
    assign layer2_outputs[838] = layer1_outputs[2883];
    assign layer2_outputs[839] = layer1_outputs[8186];
    assign layer2_outputs[840] = layer1_outputs[7733];
    assign layer2_outputs[841] = ~(layer1_outputs[10912]);
    assign layer2_outputs[842] = layer1_outputs[7639];
    assign layer2_outputs[843] = layer1_outputs[2458];
    assign layer2_outputs[844] = layer1_outputs[5289];
    assign layer2_outputs[845] = ~((layer1_outputs[9332]) ^ (layer1_outputs[12191]));
    assign layer2_outputs[846] = (layer1_outputs[4665]) & ~(layer1_outputs[3000]);
    assign layer2_outputs[847] = ~((layer1_outputs[8917]) ^ (layer1_outputs[9259]));
    assign layer2_outputs[848] = ~((layer1_outputs[5568]) | (layer1_outputs[402]));
    assign layer2_outputs[849] = ~(layer1_outputs[3990]);
    assign layer2_outputs[850] = ~(layer1_outputs[12127]);
    assign layer2_outputs[851] = ~((layer1_outputs[12411]) & (layer1_outputs[9296]));
    assign layer2_outputs[852] = layer1_outputs[10705];
    assign layer2_outputs[853] = layer1_outputs[8413];
    assign layer2_outputs[854] = layer1_outputs[2561];
    assign layer2_outputs[855] = ~(layer1_outputs[1947]);
    assign layer2_outputs[856] = layer1_outputs[1124];
    assign layer2_outputs[857] = (layer1_outputs[10252]) | (layer1_outputs[2771]);
    assign layer2_outputs[858] = (layer1_outputs[10067]) & ~(layer1_outputs[7226]);
    assign layer2_outputs[859] = ~(layer1_outputs[12281]);
    assign layer2_outputs[860] = ~(layer1_outputs[9747]);
    assign layer2_outputs[861] = 1'b0;
    assign layer2_outputs[862] = ~((layer1_outputs[2613]) | (layer1_outputs[3160]));
    assign layer2_outputs[863] = layer1_outputs[8555];
    assign layer2_outputs[864] = ~(layer1_outputs[5441]);
    assign layer2_outputs[865] = layer1_outputs[1498];
    assign layer2_outputs[866] = (layer1_outputs[4647]) ^ (layer1_outputs[8741]);
    assign layer2_outputs[867] = layer1_outputs[12406];
    assign layer2_outputs[868] = ~(layer1_outputs[6777]);
    assign layer2_outputs[869] = ~((layer1_outputs[9735]) | (layer1_outputs[5915]));
    assign layer2_outputs[870] = ~(layer1_outputs[11172]);
    assign layer2_outputs[871] = ~(layer1_outputs[9056]);
    assign layer2_outputs[872] = ~(layer1_outputs[6741]);
    assign layer2_outputs[873] = (layer1_outputs[12079]) & ~(layer1_outputs[4051]);
    assign layer2_outputs[874] = (layer1_outputs[1943]) & ~(layer1_outputs[11432]);
    assign layer2_outputs[875] = ~((layer1_outputs[9730]) | (layer1_outputs[6999]));
    assign layer2_outputs[876] = (layer1_outputs[9274]) & (layer1_outputs[9956]);
    assign layer2_outputs[877] = ~((layer1_outputs[5622]) | (layer1_outputs[8351]));
    assign layer2_outputs[878] = ~((layer1_outputs[6413]) ^ (layer1_outputs[25]));
    assign layer2_outputs[879] = ~(layer1_outputs[7560]);
    assign layer2_outputs[880] = ~(layer1_outputs[5083]);
    assign layer2_outputs[881] = layer1_outputs[6340];
    assign layer2_outputs[882] = ~((layer1_outputs[812]) & (layer1_outputs[5849]));
    assign layer2_outputs[883] = ~((layer1_outputs[2403]) ^ (layer1_outputs[7281]));
    assign layer2_outputs[884] = ~(layer1_outputs[1797]) | (layer1_outputs[3198]);
    assign layer2_outputs[885] = layer1_outputs[64];
    assign layer2_outputs[886] = layer1_outputs[4914];
    assign layer2_outputs[887] = (layer1_outputs[8431]) & (layer1_outputs[11488]);
    assign layer2_outputs[888] = (layer1_outputs[11826]) & (layer1_outputs[6683]);
    assign layer2_outputs[889] = layer1_outputs[7906];
    assign layer2_outputs[890] = (layer1_outputs[3913]) & ~(layer1_outputs[546]);
    assign layer2_outputs[891] = ~((layer1_outputs[3793]) ^ (layer1_outputs[9860]));
    assign layer2_outputs[892] = layer1_outputs[2875];
    assign layer2_outputs[893] = (layer1_outputs[10955]) & ~(layer1_outputs[3080]);
    assign layer2_outputs[894] = (layer1_outputs[12324]) & ~(layer1_outputs[7036]);
    assign layer2_outputs[895] = ~(layer1_outputs[1514]);
    assign layer2_outputs[896] = ~(layer1_outputs[8759]);
    assign layer2_outputs[897] = ~(layer1_outputs[5280]);
    assign layer2_outputs[898] = layer1_outputs[985];
    assign layer2_outputs[899] = ~((layer1_outputs[6505]) & (layer1_outputs[5193]));
    assign layer2_outputs[900] = ~((layer1_outputs[2381]) ^ (layer1_outputs[810]));
    assign layer2_outputs[901] = (layer1_outputs[11780]) & ~(layer1_outputs[5091]);
    assign layer2_outputs[902] = ~(layer1_outputs[2212]);
    assign layer2_outputs[903] = (layer1_outputs[5808]) & ~(layer1_outputs[4817]);
    assign layer2_outputs[904] = layer1_outputs[12562];
    assign layer2_outputs[905] = layer1_outputs[8026];
    assign layer2_outputs[906] = (layer1_outputs[1192]) & ~(layer1_outputs[6903]);
    assign layer2_outputs[907] = ~(layer1_outputs[3042]);
    assign layer2_outputs[908] = (layer1_outputs[5223]) & (layer1_outputs[8774]);
    assign layer2_outputs[909] = ~(layer1_outputs[11454]) | (layer1_outputs[3485]);
    assign layer2_outputs[910] = (layer1_outputs[11817]) ^ (layer1_outputs[9733]);
    assign layer2_outputs[911] = (layer1_outputs[8553]) & ~(layer1_outputs[10301]);
    assign layer2_outputs[912] = ~(layer1_outputs[8283]);
    assign layer2_outputs[913] = layer1_outputs[11430];
    assign layer2_outputs[914] = (layer1_outputs[4562]) ^ (layer1_outputs[3524]);
    assign layer2_outputs[915] = ~(layer1_outputs[4407]);
    assign layer2_outputs[916] = ~((layer1_outputs[1719]) & (layer1_outputs[6588]));
    assign layer2_outputs[917] = ~(layer1_outputs[1702]) | (layer1_outputs[11577]);
    assign layer2_outputs[918] = layer1_outputs[8915];
    assign layer2_outputs[919] = ~((layer1_outputs[5992]) | (layer1_outputs[6396]));
    assign layer2_outputs[920] = ~(layer1_outputs[6584]);
    assign layer2_outputs[921] = ~(layer1_outputs[4915]);
    assign layer2_outputs[922] = (layer1_outputs[4030]) | (layer1_outputs[11371]);
    assign layer2_outputs[923] = (layer1_outputs[888]) ^ (layer1_outputs[2686]);
    assign layer2_outputs[924] = ~(layer1_outputs[8066]);
    assign layer2_outputs[925] = (layer1_outputs[5649]) & ~(layer1_outputs[12486]);
    assign layer2_outputs[926] = ~((layer1_outputs[3743]) ^ (layer1_outputs[12227]));
    assign layer2_outputs[927] = (layer1_outputs[5703]) & ~(layer1_outputs[7324]);
    assign layer2_outputs[928] = ~(layer1_outputs[1991]) | (layer1_outputs[7772]);
    assign layer2_outputs[929] = ~(layer1_outputs[7547]);
    assign layer2_outputs[930] = ~(layer1_outputs[2576]);
    assign layer2_outputs[931] = layer1_outputs[10412];
    assign layer2_outputs[932] = ~(layer1_outputs[763]) | (layer1_outputs[12075]);
    assign layer2_outputs[933] = ~((layer1_outputs[7790]) ^ (layer1_outputs[1524]));
    assign layer2_outputs[934] = layer1_outputs[10829];
    assign layer2_outputs[935] = 1'b0;
    assign layer2_outputs[936] = (layer1_outputs[4743]) & (layer1_outputs[10057]);
    assign layer2_outputs[937] = ~(layer1_outputs[136]) | (layer1_outputs[9135]);
    assign layer2_outputs[938] = layer1_outputs[6665];
    assign layer2_outputs[939] = ~(layer1_outputs[1158]);
    assign layer2_outputs[940] = ~(layer1_outputs[7016]);
    assign layer2_outputs[941] = (layer1_outputs[12276]) | (layer1_outputs[8001]);
    assign layer2_outputs[942] = (layer1_outputs[6817]) ^ (layer1_outputs[550]);
    assign layer2_outputs[943] = (layer1_outputs[3848]) & ~(layer1_outputs[2074]);
    assign layer2_outputs[944] = ~(layer1_outputs[669]);
    assign layer2_outputs[945] = layer1_outputs[6831];
    assign layer2_outputs[946] = ~(layer1_outputs[8315]);
    assign layer2_outputs[947] = (layer1_outputs[5355]) & ~(layer1_outputs[4704]);
    assign layer2_outputs[948] = layer1_outputs[2188];
    assign layer2_outputs[949] = 1'b0;
    assign layer2_outputs[950] = (layer1_outputs[294]) | (layer1_outputs[12759]);
    assign layer2_outputs[951] = ~(layer1_outputs[8813]);
    assign layer2_outputs[952] = ~(layer1_outputs[10063]) | (layer1_outputs[6070]);
    assign layer2_outputs[953] = ~((layer1_outputs[337]) ^ (layer1_outputs[6084]));
    assign layer2_outputs[954] = ~(layer1_outputs[8132]);
    assign layer2_outputs[955] = (layer1_outputs[2749]) & (layer1_outputs[5520]);
    assign layer2_outputs[956] = layer1_outputs[646];
    assign layer2_outputs[957] = layer1_outputs[482];
    assign layer2_outputs[958] = layer1_outputs[10366];
    assign layer2_outputs[959] = ~((layer1_outputs[6477]) ^ (layer1_outputs[5393]));
    assign layer2_outputs[960] = layer1_outputs[11280];
    assign layer2_outputs[961] = (layer1_outputs[11291]) & ~(layer1_outputs[2271]);
    assign layer2_outputs[962] = ~(layer1_outputs[8519]);
    assign layer2_outputs[963] = (layer1_outputs[9466]) & ~(layer1_outputs[7227]);
    assign layer2_outputs[964] = layer1_outputs[11370];
    assign layer2_outputs[965] = ~((layer1_outputs[7723]) ^ (layer1_outputs[4004]));
    assign layer2_outputs[966] = ~((layer1_outputs[3170]) & (layer1_outputs[12088]));
    assign layer2_outputs[967] = layer1_outputs[7857];
    assign layer2_outputs[968] = (layer1_outputs[4942]) & (layer1_outputs[3005]);
    assign layer2_outputs[969] = (layer1_outputs[2967]) & ~(layer1_outputs[5367]);
    assign layer2_outputs[970] = (layer1_outputs[7900]) ^ (layer1_outputs[4550]);
    assign layer2_outputs[971] = ~(layer1_outputs[10766]);
    assign layer2_outputs[972] = layer1_outputs[12284];
    assign layer2_outputs[973] = (layer1_outputs[4998]) & ~(layer1_outputs[10794]);
    assign layer2_outputs[974] = ~((layer1_outputs[10255]) ^ (layer1_outputs[582]));
    assign layer2_outputs[975] = layer1_outputs[713];
    assign layer2_outputs[976] = ~((layer1_outputs[5444]) ^ (layer1_outputs[5901]));
    assign layer2_outputs[977] = ~(layer1_outputs[241]);
    assign layer2_outputs[978] = layer1_outputs[9104];
    assign layer2_outputs[979] = ~(layer1_outputs[11283]) | (layer1_outputs[4058]);
    assign layer2_outputs[980] = 1'b0;
    assign layer2_outputs[981] = layer1_outputs[6041];
    assign layer2_outputs[982] = ~(layer1_outputs[11969]);
    assign layer2_outputs[983] = (layer1_outputs[7031]) ^ (layer1_outputs[2968]);
    assign layer2_outputs[984] = (layer1_outputs[10136]) ^ (layer1_outputs[7597]);
    assign layer2_outputs[985] = layer1_outputs[2076];
    assign layer2_outputs[986] = ~(layer1_outputs[9961]) | (layer1_outputs[4773]);
    assign layer2_outputs[987] = (layer1_outputs[1313]) ^ (layer1_outputs[610]);
    assign layer2_outputs[988] = ~((layer1_outputs[6130]) | (layer1_outputs[3483]));
    assign layer2_outputs[989] = (layer1_outputs[2074]) ^ (layer1_outputs[11830]);
    assign layer2_outputs[990] = ~(layer1_outputs[9342]);
    assign layer2_outputs[991] = ~(layer1_outputs[4434]) | (layer1_outputs[1946]);
    assign layer2_outputs[992] = (layer1_outputs[7487]) & ~(layer1_outputs[5898]);
    assign layer2_outputs[993] = layer1_outputs[9646];
    assign layer2_outputs[994] = layer1_outputs[7481];
    assign layer2_outputs[995] = (layer1_outputs[3224]) ^ (layer1_outputs[8711]);
    assign layer2_outputs[996] = (layer1_outputs[11710]) ^ (layer1_outputs[10085]);
    assign layer2_outputs[997] = layer1_outputs[10787];
    assign layer2_outputs[998] = ~(layer1_outputs[3665]) | (layer1_outputs[7171]);
    assign layer2_outputs[999] = layer1_outputs[3710];
    assign layer2_outputs[1000] = ~(layer1_outputs[4608]);
    assign layer2_outputs[1001] = ~(layer1_outputs[10543]);
    assign layer2_outputs[1002] = (layer1_outputs[6868]) ^ (layer1_outputs[2369]);
    assign layer2_outputs[1003] = (layer1_outputs[12443]) | (layer1_outputs[10293]);
    assign layer2_outputs[1004] = ~((layer1_outputs[10735]) | (layer1_outputs[9770]));
    assign layer2_outputs[1005] = ~((layer1_outputs[1062]) | (layer1_outputs[10413]));
    assign layer2_outputs[1006] = ~(layer1_outputs[3196]);
    assign layer2_outputs[1007] = ~(layer1_outputs[11334]) | (layer1_outputs[3146]);
    assign layer2_outputs[1008] = (layer1_outputs[11737]) ^ (layer1_outputs[3001]);
    assign layer2_outputs[1009] = layer1_outputs[5947];
    assign layer2_outputs[1010] = ~(layer1_outputs[2791]);
    assign layer2_outputs[1011] = (layer1_outputs[3857]) & ~(layer1_outputs[5473]);
    assign layer2_outputs[1012] = ~(layer1_outputs[11350]);
    assign layer2_outputs[1013] = layer1_outputs[11806];
    assign layer2_outputs[1014] = layer1_outputs[9741];
    assign layer2_outputs[1015] = (layer1_outputs[8575]) ^ (layer1_outputs[10786]);
    assign layer2_outputs[1016] = layer1_outputs[9930];
    assign layer2_outputs[1017] = layer1_outputs[11222];
    assign layer2_outputs[1018] = ~(layer1_outputs[5467]);
    assign layer2_outputs[1019] = layer1_outputs[9837];
    assign layer2_outputs[1020] = ~(layer1_outputs[5179]);
    assign layer2_outputs[1021] = ~(layer1_outputs[3703]);
    assign layer2_outputs[1022] = (layer1_outputs[10221]) & ~(layer1_outputs[10034]);
    assign layer2_outputs[1023] = layer1_outputs[1583];
    assign layer2_outputs[1024] = ~(layer1_outputs[12082]);
    assign layer2_outputs[1025] = ~(layer1_outputs[1417]);
    assign layer2_outputs[1026] = layer1_outputs[8053];
    assign layer2_outputs[1027] = ~(layer1_outputs[3300]);
    assign layer2_outputs[1028] = ~(layer1_outputs[4856]) | (layer1_outputs[12049]);
    assign layer2_outputs[1029] = ~(layer1_outputs[8074]);
    assign layer2_outputs[1030] = layer1_outputs[11987];
    assign layer2_outputs[1031] = layer1_outputs[250];
    assign layer2_outputs[1032] = (layer1_outputs[12574]) & ~(layer1_outputs[7397]);
    assign layer2_outputs[1033] = ~(layer1_outputs[9106]);
    assign layer2_outputs[1034] = (layer1_outputs[6006]) | (layer1_outputs[1246]);
    assign layer2_outputs[1035] = ~(layer1_outputs[5070]) | (layer1_outputs[12195]);
    assign layer2_outputs[1036] = (layer1_outputs[3749]) | (layer1_outputs[4660]);
    assign layer2_outputs[1037] = (layer1_outputs[5981]) | (layer1_outputs[2102]);
    assign layer2_outputs[1038] = (layer1_outputs[3803]) ^ (layer1_outputs[8492]);
    assign layer2_outputs[1039] = (layer1_outputs[7403]) | (layer1_outputs[204]);
    assign layer2_outputs[1040] = layer1_outputs[1695];
    assign layer2_outputs[1041] = (layer1_outputs[617]) & ~(layer1_outputs[5510]);
    assign layer2_outputs[1042] = ~((layer1_outputs[10403]) | (layer1_outputs[9812]));
    assign layer2_outputs[1043] = (layer1_outputs[144]) & (layer1_outputs[7580]);
    assign layer2_outputs[1044] = ~((layer1_outputs[10935]) | (layer1_outputs[1289]));
    assign layer2_outputs[1045] = ~((layer1_outputs[10671]) ^ (layer1_outputs[5932]));
    assign layer2_outputs[1046] = ~((layer1_outputs[7885]) ^ (layer1_outputs[412]));
    assign layer2_outputs[1047] = (layer1_outputs[4941]) | (layer1_outputs[6580]);
    assign layer2_outputs[1048] = ~((layer1_outputs[12327]) & (layer1_outputs[4207]));
    assign layer2_outputs[1049] = ~(layer1_outputs[10606]);
    assign layer2_outputs[1050] = ~(layer1_outputs[4404]);
    assign layer2_outputs[1051] = ~(layer1_outputs[4766]);
    assign layer2_outputs[1052] = layer1_outputs[10330];
    assign layer2_outputs[1053] = ~((layer1_outputs[8533]) | (layer1_outputs[1229]));
    assign layer2_outputs[1054] = ~(layer1_outputs[10282]) | (layer1_outputs[5489]);
    assign layer2_outputs[1055] = layer1_outputs[2593];
    assign layer2_outputs[1056] = ~(layer1_outputs[790]);
    assign layer2_outputs[1057] = ~(layer1_outputs[10980]);
    assign layer2_outputs[1058] = ~(layer1_outputs[913]);
    assign layer2_outputs[1059] = (layer1_outputs[166]) & ~(layer1_outputs[5829]);
    assign layer2_outputs[1060] = ~(layer1_outputs[1388]);
    assign layer2_outputs[1061] = ~(layer1_outputs[11940]);
    assign layer2_outputs[1062] = ~((layer1_outputs[6542]) & (layer1_outputs[12659]));
    assign layer2_outputs[1063] = layer1_outputs[9273];
    assign layer2_outputs[1064] = ~(layer1_outputs[121]);
    assign layer2_outputs[1065] = (layer1_outputs[3019]) & ~(layer1_outputs[2137]);
    assign layer2_outputs[1066] = layer1_outputs[10876];
    assign layer2_outputs[1067] = ~(layer1_outputs[6907]);
    assign layer2_outputs[1068] = ~(layer1_outputs[11842]) | (layer1_outputs[3870]);
    assign layer2_outputs[1069] = (layer1_outputs[10540]) & ~(layer1_outputs[7365]);
    assign layer2_outputs[1070] = ~(layer1_outputs[5140]) | (layer1_outputs[11761]);
    assign layer2_outputs[1071] = ~(layer1_outputs[2667]);
    assign layer2_outputs[1072] = (layer1_outputs[5451]) & ~(layer1_outputs[3398]);
    assign layer2_outputs[1073] = layer1_outputs[102];
    assign layer2_outputs[1074] = (layer1_outputs[9163]) & (layer1_outputs[9706]);
    assign layer2_outputs[1075] = (layer1_outputs[11314]) & ~(layer1_outputs[8241]);
    assign layer2_outputs[1076] = ~(layer1_outputs[7603]);
    assign layer2_outputs[1077] = layer1_outputs[1188];
    assign layer2_outputs[1078] = layer1_outputs[6200];
    assign layer2_outputs[1079] = ~((layer1_outputs[61]) & (layer1_outputs[598]));
    assign layer2_outputs[1080] = layer1_outputs[5846];
    assign layer2_outputs[1081] = ~(layer1_outputs[9536]);
    assign layer2_outputs[1082] = ~(layer1_outputs[6501]);
    assign layer2_outputs[1083] = 1'b1;
    assign layer2_outputs[1084] = ~(layer1_outputs[8762]) | (layer1_outputs[8101]);
    assign layer2_outputs[1085] = ~(layer1_outputs[6418]);
    assign layer2_outputs[1086] = ~(layer1_outputs[7454]);
    assign layer2_outputs[1087] = ~(layer1_outputs[6819]);
    assign layer2_outputs[1088] = ~(layer1_outputs[8581]);
    assign layer2_outputs[1089] = ~(layer1_outputs[2098]);
    assign layer2_outputs[1090] = layer1_outputs[2027];
    assign layer2_outputs[1091] = (layer1_outputs[8828]) | (layer1_outputs[7784]);
    assign layer2_outputs[1092] = layer1_outputs[2006];
    assign layer2_outputs[1093] = (layer1_outputs[10971]) ^ (layer1_outputs[7560]);
    assign layer2_outputs[1094] = ~(layer1_outputs[1826]);
    assign layer2_outputs[1095] = (layer1_outputs[9554]) ^ (layer1_outputs[11601]);
    assign layer2_outputs[1096] = ~(layer1_outputs[11571]);
    assign layer2_outputs[1097] = ~((layer1_outputs[6149]) ^ (layer1_outputs[9759]));
    assign layer2_outputs[1098] = (layer1_outputs[7490]) ^ (layer1_outputs[11706]);
    assign layer2_outputs[1099] = 1'b1;
    assign layer2_outputs[1100] = ~((layer1_outputs[12648]) ^ (layer1_outputs[7114]));
    assign layer2_outputs[1101] = ~(layer1_outputs[8733]) | (layer1_outputs[8749]);
    assign layer2_outputs[1102] = layer1_outputs[10236];
    assign layer2_outputs[1103] = ~(layer1_outputs[1215]);
    assign layer2_outputs[1104] = ~(layer1_outputs[946]);
    assign layer2_outputs[1105] = layer1_outputs[11984];
    assign layer2_outputs[1106] = (layer1_outputs[7267]) ^ (layer1_outputs[10369]);
    assign layer2_outputs[1107] = ~(layer1_outputs[11416]);
    assign layer2_outputs[1108] = ~((layer1_outputs[10515]) ^ (layer1_outputs[2191]));
    assign layer2_outputs[1109] = (layer1_outputs[3280]) | (layer1_outputs[2142]);
    assign layer2_outputs[1110] = (layer1_outputs[1302]) & ~(layer1_outputs[7070]);
    assign layer2_outputs[1111] = (layer1_outputs[2055]) & ~(layer1_outputs[8434]);
    assign layer2_outputs[1112] = layer1_outputs[10805];
    assign layer2_outputs[1113] = ~((layer1_outputs[956]) ^ (layer1_outputs[10141]));
    assign layer2_outputs[1114] = (layer1_outputs[2403]) & (layer1_outputs[1230]);
    assign layer2_outputs[1115] = ~((layer1_outputs[2388]) ^ (layer1_outputs[11181]));
    assign layer2_outputs[1116] = ~((layer1_outputs[1193]) & (layer1_outputs[4834]));
    assign layer2_outputs[1117] = ~(layer1_outputs[10396]);
    assign layer2_outputs[1118] = ~(layer1_outputs[7175]);
    assign layer2_outputs[1119] = ~(layer1_outputs[309]);
    assign layer2_outputs[1120] = ~(layer1_outputs[4468]);
    assign layer2_outputs[1121] = layer1_outputs[1484];
    assign layer2_outputs[1122] = (layer1_outputs[2987]) & (layer1_outputs[10055]);
    assign layer2_outputs[1123] = (layer1_outputs[7008]) & (layer1_outputs[8273]);
    assign layer2_outputs[1124] = ~(layer1_outputs[4966]);
    assign layer2_outputs[1125] = (layer1_outputs[6712]) & (layer1_outputs[6824]);
    assign layer2_outputs[1126] = layer1_outputs[165];
    assign layer2_outputs[1127] = ~(layer1_outputs[4277]);
    assign layer2_outputs[1128] = ~(layer1_outputs[1159]);
    assign layer2_outputs[1129] = (layer1_outputs[6872]) | (layer1_outputs[8032]);
    assign layer2_outputs[1130] = ~(layer1_outputs[12017]);
    assign layer2_outputs[1131] = ~(layer1_outputs[773]);
    assign layer2_outputs[1132] = (layer1_outputs[6195]) ^ (layer1_outputs[8769]);
    assign layer2_outputs[1133] = ~(layer1_outputs[9730]);
    assign layer2_outputs[1134] = ~(layer1_outputs[5840]);
    assign layer2_outputs[1135] = ~(layer1_outputs[6081]);
    assign layer2_outputs[1136] = ~(layer1_outputs[6597]) | (layer1_outputs[11132]);
    assign layer2_outputs[1137] = ~((layer1_outputs[11878]) & (layer1_outputs[9897]));
    assign layer2_outputs[1138] = (layer1_outputs[8120]) & (layer1_outputs[497]);
    assign layer2_outputs[1139] = layer1_outputs[9577];
    assign layer2_outputs[1140] = ~(layer1_outputs[12469]);
    assign layer2_outputs[1141] = ~(layer1_outputs[7907]) | (layer1_outputs[10125]);
    assign layer2_outputs[1142] = ~(layer1_outputs[11158]);
    assign layer2_outputs[1143] = (layer1_outputs[8349]) & ~(layer1_outputs[1872]);
    assign layer2_outputs[1144] = (layer1_outputs[8722]) & ~(layer1_outputs[3718]);
    assign layer2_outputs[1145] = ~((layer1_outputs[6029]) & (layer1_outputs[4866]));
    assign layer2_outputs[1146] = ~((layer1_outputs[1295]) & (layer1_outputs[4365]));
    assign layer2_outputs[1147] = ~(layer1_outputs[11550]) | (layer1_outputs[9390]);
    assign layer2_outputs[1148] = ~(layer1_outputs[489]);
    assign layer2_outputs[1149] = ~(layer1_outputs[9676]);
    assign layer2_outputs[1150] = ~((layer1_outputs[1647]) | (layer1_outputs[7324]));
    assign layer2_outputs[1151] = ~((layer1_outputs[4421]) ^ (layer1_outputs[10906]));
    assign layer2_outputs[1152] = ~(layer1_outputs[5]);
    assign layer2_outputs[1153] = ~(layer1_outputs[159]) | (layer1_outputs[8827]);
    assign layer2_outputs[1154] = ~((layer1_outputs[10605]) ^ (layer1_outputs[3472]));
    assign layer2_outputs[1155] = (layer1_outputs[6119]) & ~(layer1_outputs[671]);
    assign layer2_outputs[1156] = (layer1_outputs[11800]) | (layer1_outputs[1564]);
    assign layer2_outputs[1157] = ~(layer1_outputs[8085]);
    assign layer2_outputs[1158] = (layer1_outputs[1515]) ^ (layer1_outputs[2805]);
    assign layer2_outputs[1159] = ~(layer1_outputs[5872]);
    assign layer2_outputs[1160] = ~((layer1_outputs[10412]) & (layer1_outputs[10567]));
    assign layer2_outputs[1161] = (layer1_outputs[4996]) | (layer1_outputs[6723]);
    assign layer2_outputs[1162] = ~(layer1_outputs[5973]);
    assign layer2_outputs[1163] = (layer1_outputs[4834]) ^ (layer1_outputs[4663]);
    assign layer2_outputs[1164] = layer1_outputs[11029];
    assign layer2_outputs[1165] = (layer1_outputs[12398]) | (layer1_outputs[6995]);
    assign layer2_outputs[1166] = (layer1_outputs[7651]) & (layer1_outputs[4195]);
    assign layer2_outputs[1167] = layer1_outputs[2588];
    assign layer2_outputs[1168] = layer1_outputs[10976];
    assign layer2_outputs[1169] = (layer1_outputs[9507]) ^ (layer1_outputs[3380]);
    assign layer2_outputs[1170] = ~((layer1_outputs[7167]) | (layer1_outputs[8158]));
    assign layer2_outputs[1171] = (layer1_outputs[12312]) ^ (layer1_outputs[5353]);
    assign layer2_outputs[1172] = ~(layer1_outputs[2657]);
    assign layer2_outputs[1173] = ~((layer1_outputs[7642]) ^ (layer1_outputs[11075]));
    assign layer2_outputs[1174] = ~(layer1_outputs[7545]);
    assign layer2_outputs[1175] = (layer1_outputs[7798]) ^ (layer1_outputs[5088]);
    assign layer2_outputs[1176] = (layer1_outputs[8846]) ^ (layer1_outputs[5199]);
    assign layer2_outputs[1177] = ~((layer1_outputs[9234]) ^ (layer1_outputs[8017]));
    assign layer2_outputs[1178] = layer1_outputs[6773];
    assign layer2_outputs[1179] = ~(layer1_outputs[4755]) | (layer1_outputs[2340]);
    assign layer2_outputs[1180] = ~(layer1_outputs[10631]) | (layer1_outputs[6215]);
    assign layer2_outputs[1181] = layer1_outputs[7835];
    assign layer2_outputs[1182] = ~(layer1_outputs[8952]);
    assign layer2_outputs[1183] = ~((layer1_outputs[9674]) | (layer1_outputs[12250]));
    assign layer2_outputs[1184] = ~((layer1_outputs[6190]) | (layer1_outputs[918]));
    assign layer2_outputs[1185] = ~(layer1_outputs[6954]);
    assign layer2_outputs[1186] = ~(layer1_outputs[8149]);
    assign layer2_outputs[1187] = layer1_outputs[10269];
    assign layer2_outputs[1188] = (layer1_outputs[7801]) | (layer1_outputs[6990]);
    assign layer2_outputs[1189] = layer1_outputs[3745];
    assign layer2_outputs[1190] = ~((layer1_outputs[2454]) | (layer1_outputs[1531]));
    assign layer2_outputs[1191] = ~((layer1_outputs[1232]) | (layer1_outputs[10510]));
    assign layer2_outputs[1192] = ~(layer1_outputs[967]);
    assign layer2_outputs[1193] = ~(layer1_outputs[1698]);
    assign layer2_outputs[1194] = ~(layer1_outputs[1907]);
    assign layer2_outputs[1195] = ~(layer1_outputs[12317]);
    assign layer2_outputs[1196] = layer1_outputs[11271];
    assign layer2_outputs[1197] = ~(layer1_outputs[2823]);
    assign layer2_outputs[1198] = (layer1_outputs[11388]) & ~(layer1_outputs[2901]);
    assign layer2_outputs[1199] = (layer1_outputs[10345]) ^ (layer1_outputs[6192]);
    assign layer2_outputs[1200] = (layer1_outputs[1544]) & ~(layer1_outputs[8014]);
    assign layer2_outputs[1201] = (layer1_outputs[11035]) & ~(layer1_outputs[1553]);
    assign layer2_outputs[1202] = (layer1_outputs[11897]) ^ (layer1_outputs[2656]);
    assign layer2_outputs[1203] = (layer1_outputs[6634]) & (layer1_outputs[7621]);
    assign layer2_outputs[1204] = layer1_outputs[7499];
    assign layer2_outputs[1205] = ~(layer1_outputs[9734]);
    assign layer2_outputs[1206] = layer1_outputs[7654];
    assign layer2_outputs[1207] = layer1_outputs[10177];
    assign layer2_outputs[1208] = (layer1_outputs[1125]) & ~(layer1_outputs[7111]);
    assign layer2_outputs[1209] = layer1_outputs[3463];
    assign layer2_outputs[1210] = ~(layer1_outputs[9964]) | (layer1_outputs[2073]);
    assign layer2_outputs[1211] = ~((layer1_outputs[8926]) | (layer1_outputs[6675]));
    assign layer2_outputs[1212] = ~(layer1_outputs[7034]) | (layer1_outputs[9341]);
    assign layer2_outputs[1213] = ~(layer1_outputs[10951]);
    assign layer2_outputs[1214] = (layer1_outputs[5969]) & ~(layer1_outputs[8873]);
    assign layer2_outputs[1215] = (layer1_outputs[823]) ^ (layer1_outputs[2534]);
    assign layer2_outputs[1216] = layer1_outputs[2934];
    assign layer2_outputs[1217] = ~(layer1_outputs[766]);
    assign layer2_outputs[1218] = layer1_outputs[2101];
    assign layer2_outputs[1219] = ~(layer1_outputs[9780]) | (layer1_outputs[4352]);
    assign layer2_outputs[1220] = ~(layer1_outputs[10089]);
    assign layer2_outputs[1221] = layer1_outputs[10841];
    assign layer2_outputs[1222] = (layer1_outputs[6831]) & ~(layer1_outputs[4172]);
    assign layer2_outputs[1223] = ~(layer1_outputs[8383]);
    assign layer2_outputs[1224] = layer1_outputs[3658];
    assign layer2_outputs[1225] = ~((layer1_outputs[3205]) & (layer1_outputs[12754]));
    assign layer2_outputs[1226] = 1'b0;
    assign layer2_outputs[1227] = ~(layer1_outputs[6988]);
    assign layer2_outputs[1228] = (layer1_outputs[8291]) & (layer1_outputs[281]);
    assign layer2_outputs[1229] = (layer1_outputs[2925]) | (layer1_outputs[11363]);
    assign layer2_outputs[1230] = (layer1_outputs[11533]) | (layer1_outputs[8372]);
    assign layer2_outputs[1231] = layer1_outputs[7127];
    assign layer2_outputs[1232] = layer1_outputs[12285];
    assign layer2_outputs[1233] = (layer1_outputs[81]) ^ (layer1_outputs[12576]);
    assign layer2_outputs[1234] = (layer1_outputs[5059]) ^ (layer1_outputs[8312]);
    assign layer2_outputs[1235] = layer1_outputs[10265];
    assign layer2_outputs[1236] = ~(layer1_outputs[2179]) | (layer1_outputs[7576]);
    assign layer2_outputs[1237] = layer1_outputs[5243];
    assign layer2_outputs[1238] = layer1_outputs[7621];
    assign layer2_outputs[1239] = (layer1_outputs[8652]) & (layer1_outputs[2836]);
    assign layer2_outputs[1240] = ~(layer1_outputs[5255]);
    assign layer2_outputs[1241] = (layer1_outputs[27]) & ~(layer1_outputs[10582]);
    assign layer2_outputs[1242] = (layer1_outputs[4256]) ^ (layer1_outputs[3022]);
    assign layer2_outputs[1243] = ~(layer1_outputs[10687]);
    assign layer2_outputs[1244] = (layer1_outputs[11985]) ^ (layer1_outputs[9476]);
    assign layer2_outputs[1245] = ~(layer1_outputs[395]);
    assign layer2_outputs[1246] = layer1_outputs[7168];
    assign layer2_outputs[1247] = ~((layer1_outputs[3013]) ^ (layer1_outputs[8220]));
    assign layer2_outputs[1248] = layer1_outputs[8777];
    assign layer2_outputs[1249] = ~((layer1_outputs[2819]) & (layer1_outputs[1815]));
    assign layer2_outputs[1250] = ~(layer1_outputs[1604]);
    assign layer2_outputs[1251] = ~((layer1_outputs[6508]) | (layer1_outputs[7312]));
    assign layer2_outputs[1252] = (layer1_outputs[11313]) ^ (layer1_outputs[7678]);
    assign layer2_outputs[1253] = (layer1_outputs[12383]) & ~(layer1_outputs[1065]);
    assign layer2_outputs[1254] = (layer1_outputs[10344]) ^ (layer1_outputs[7693]);
    assign layer2_outputs[1255] = ~(layer1_outputs[12043]);
    assign layer2_outputs[1256] = ~((layer1_outputs[8278]) ^ (layer1_outputs[3101]));
    assign layer2_outputs[1257] = layer1_outputs[8259];
    assign layer2_outputs[1258] = ~(layer1_outputs[9096]) | (layer1_outputs[2430]);
    assign layer2_outputs[1259] = (layer1_outputs[8791]) & (layer1_outputs[11923]);
    assign layer2_outputs[1260] = layer1_outputs[940];
    assign layer2_outputs[1261] = (layer1_outputs[8921]) & (layer1_outputs[1595]);
    assign layer2_outputs[1262] = (layer1_outputs[2375]) | (layer1_outputs[18]);
    assign layer2_outputs[1263] = ~((layer1_outputs[6135]) | (layer1_outputs[11922]));
    assign layer2_outputs[1264] = (layer1_outputs[2485]) ^ (layer1_outputs[9200]);
    assign layer2_outputs[1265] = ~(layer1_outputs[2279]) | (layer1_outputs[1006]);
    assign layer2_outputs[1266] = (layer1_outputs[2540]) & (layer1_outputs[4674]);
    assign layer2_outputs[1267] = (layer1_outputs[10008]) ^ (layer1_outputs[10127]);
    assign layer2_outputs[1268] = layer1_outputs[3294];
    assign layer2_outputs[1269] = 1'b1;
    assign layer2_outputs[1270] = ~(layer1_outputs[9125]) | (layer1_outputs[11497]);
    assign layer2_outputs[1271] = ~(layer1_outputs[6062]);
    assign layer2_outputs[1272] = ~((layer1_outputs[6022]) & (layer1_outputs[12234]));
    assign layer2_outputs[1273] = (layer1_outputs[5278]) & (layer1_outputs[4517]);
    assign layer2_outputs[1274] = layer1_outputs[5752];
    assign layer2_outputs[1275] = (layer1_outputs[330]) & ~(layer1_outputs[1986]);
    assign layer2_outputs[1276] = ~((layer1_outputs[10364]) ^ (layer1_outputs[1168]));
    assign layer2_outputs[1277] = ~(layer1_outputs[5847]) | (layer1_outputs[9141]);
    assign layer2_outputs[1278] = layer1_outputs[7608];
    assign layer2_outputs[1279] = layer1_outputs[1159];
    assign layer2_outputs[1280] = ~(layer1_outputs[5167]) | (layer1_outputs[10114]);
    assign layer2_outputs[1281] = ~(layer1_outputs[11326]);
    assign layer2_outputs[1282] = layer1_outputs[8233];
    assign layer2_outputs[1283] = ~(layer1_outputs[7220]);
    assign layer2_outputs[1284] = ~(layer1_outputs[9791]);
    assign layer2_outputs[1285] = (layer1_outputs[10459]) & (layer1_outputs[12266]);
    assign layer2_outputs[1286] = (layer1_outputs[9944]) & ~(layer1_outputs[3070]);
    assign layer2_outputs[1287] = (layer1_outputs[11290]) | (layer1_outputs[12758]);
    assign layer2_outputs[1288] = layer1_outputs[12068];
    assign layer2_outputs[1289] = ~((layer1_outputs[12210]) | (layer1_outputs[10088]));
    assign layer2_outputs[1290] = (layer1_outputs[3946]) & (layer1_outputs[6889]);
    assign layer2_outputs[1291] = ~(layer1_outputs[6749]);
    assign layer2_outputs[1292] = ~((layer1_outputs[3779]) ^ (layer1_outputs[3377]));
    assign layer2_outputs[1293] = ~((layer1_outputs[7957]) | (layer1_outputs[584]));
    assign layer2_outputs[1294] = layer1_outputs[826];
    assign layer2_outputs[1295] = layer1_outputs[5111];
    assign layer2_outputs[1296] = ~(layer1_outputs[7349]);
    assign layer2_outputs[1297] = ~(layer1_outputs[3151]) | (layer1_outputs[10460]);
    assign layer2_outputs[1298] = layer1_outputs[3545];
    assign layer2_outputs[1299] = ~(layer1_outputs[10484]);
    assign layer2_outputs[1300] = (layer1_outputs[2800]) ^ (layer1_outputs[2704]);
    assign layer2_outputs[1301] = layer1_outputs[8834];
    assign layer2_outputs[1302] = (layer1_outputs[11508]) & ~(layer1_outputs[4655]);
    assign layer2_outputs[1303] = ~(layer1_outputs[5549]);
    assign layer2_outputs[1304] = (layer1_outputs[2818]) ^ (layer1_outputs[4640]);
    assign layer2_outputs[1305] = ~((layer1_outputs[2749]) & (layer1_outputs[9630]));
    assign layer2_outputs[1306] = layer1_outputs[4369];
    assign layer2_outputs[1307] = (layer1_outputs[4316]) ^ (layer1_outputs[10246]);
    assign layer2_outputs[1308] = ~(layer1_outputs[3079]);
    assign layer2_outputs[1309] = layer1_outputs[10830];
    assign layer2_outputs[1310] = ~((layer1_outputs[6232]) & (layer1_outputs[3752]));
    assign layer2_outputs[1311] = ~(layer1_outputs[5891]);
    assign layer2_outputs[1312] = ~(layer1_outputs[10678]);
    assign layer2_outputs[1313] = layer1_outputs[5627];
    assign layer2_outputs[1314] = layer1_outputs[3676];
    assign layer2_outputs[1315] = layer1_outputs[10148];
    assign layer2_outputs[1316] = ~(layer1_outputs[9384]);
    assign layer2_outputs[1317] = ~(layer1_outputs[8854]);
    assign layer2_outputs[1318] = layer1_outputs[4485];
    assign layer2_outputs[1319] = ~(layer1_outputs[9868]) | (layer1_outputs[5381]);
    assign layer2_outputs[1320] = ~(layer1_outputs[3166]);
    assign layer2_outputs[1321] = ~(layer1_outputs[8476]) | (layer1_outputs[8734]);
    assign layer2_outputs[1322] = (layer1_outputs[8656]) & (layer1_outputs[724]);
    assign layer2_outputs[1323] = layer1_outputs[5045];
    assign layer2_outputs[1324] = ~(layer1_outputs[3697]);
    assign layer2_outputs[1325] = ~(layer1_outputs[2027]) | (layer1_outputs[10848]);
    assign layer2_outputs[1326] = ~(layer1_outputs[7707]) | (layer1_outputs[1515]);
    assign layer2_outputs[1327] = ~(layer1_outputs[10663]);
    assign layer2_outputs[1328] = layer1_outputs[2394];
    assign layer2_outputs[1329] = layer1_outputs[4490];
    assign layer2_outputs[1330] = (layer1_outputs[9585]) & ~(layer1_outputs[1214]);
    assign layer2_outputs[1331] = ~((layer1_outputs[5798]) | (layer1_outputs[9955]));
    assign layer2_outputs[1332] = ~(layer1_outputs[8003]) | (layer1_outputs[21]);
    assign layer2_outputs[1333] = (layer1_outputs[5753]) ^ (layer1_outputs[9493]);
    assign layer2_outputs[1334] = (layer1_outputs[5125]) & ~(layer1_outputs[10619]);
    assign layer2_outputs[1335] = ~(layer1_outputs[9501]);
    assign layer2_outputs[1336] = layer1_outputs[4536];
    assign layer2_outputs[1337] = layer1_outputs[11085];
    assign layer2_outputs[1338] = ~((layer1_outputs[6540]) | (layer1_outputs[1620]));
    assign layer2_outputs[1339] = ~(layer1_outputs[1082]);
    assign layer2_outputs[1340] = (layer1_outputs[6274]) ^ (layer1_outputs[8157]);
    assign layer2_outputs[1341] = layer1_outputs[2974];
    assign layer2_outputs[1342] = (layer1_outputs[9782]) & (layer1_outputs[5839]);
    assign layer2_outputs[1343] = 1'b0;
    assign layer2_outputs[1344] = ~((layer1_outputs[3780]) | (layer1_outputs[12020]));
    assign layer2_outputs[1345] = ~((layer1_outputs[1248]) | (layer1_outputs[10102]));
    assign layer2_outputs[1346] = layer1_outputs[3003];
    assign layer2_outputs[1347] = ~(layer1_outputs[9738]) | (layer1_outputs[8806]);
    assign layer2_outputs[1348] = 1'b1;
    assign layer2_outputs[1349] = layer1_outputs[9042];
    assign layer2_outputs[1350] = ~(layer1_outputs[10802]) | (layer1_outputs[11262]);
    assign layer2_outputs[1351] = layer1_outputs[10894];
    assign layer2_outputs[1352] = (layer1_outputs[7971]) ^ (layer1_outputs[8603]);
    assign layer2_outputs[1353] = layer1_outputs[9651];
    assign layer2_outputs[1354] = ~(layer1_outputs[3234]);
    assign layer2_outputs[1355] = layer1_outputs[1992];
    assign layer2_outputs[1356] = 1'b1;
    assign layer2_outputs[1357] = (layer1_outputs[5514]) | (layer1_outputs[12062]);
    assign layer2_outputs[1358] = ~(layer1_outputs[12252]);
    assign layer2_outputs[1359] = ~(layer1_outputs[7773]);
    assign layer2_outputs[1360] = ~(layer1_outputs[11764]);
    assign layer2_outputs[1361] = ~((layer1_outputs[6205]) ^ (layer1_outputs[4430]));
    assign layer2_outputs[1362] = layer1_outputs[1067];
    assign layer2_outputs[1363] = (layer1_outputs[571]) & ~(layer1_outputs[2744]);
    assign layer2_outputs[1364] = ~(layer1_outputs[11853]) | (layer1_outputs[8425]);
    assign layer2_outputs[1365] = (layer1_outputs[12703]) & ~(layer1_outputs[10138]);
    assign layer2_outputs[1366] = (layer1_outputs[10950]) | (layer1_outputs[8136]);
    assign layer2_outputs[1367] = layer1_outputs[3861];
    assign layer2_outputs[1368] = ~((layer1_outputs[1346]) ^ (layer1_outputs[496]));
    assign layer2_outputs[1369] = layer1_outputs[1978];
    assign layer2_outputs[1370] = ~(layer1_outputs[11905]);
    assign layer2_outputs[1371] = ~((layer1_outputs[12492]) ^ (layer1_outputs[2058]));
    assign layer2_outputs[1372] = ~((layer1_outputs[1572]) ^ (layer1_outputs[9995]));
    assign layer2_outputs[1373] = (layer1_outputs[4039]) & ~(layer1_outputs[2468]);
    assign layer2_outputs[1374] = ~((layer1_outputs[639]) | (layer1_outputs[1570]));
    assign layer2_outputs[1375] = ~(layer1_outputs[8642]);
    assign layer2_outputs[1376] = ~(layer1_outputs[6332]) | (layer1_outputs[8679]);
    assign layer2_outputs[1377] = ~((layer1_outputs[3605]) | (layer1_outputs[6969]));
    assign layer2_outputs[1378] = ~((layer1_outputs[5782]) ^ (layer1_outputs[100]));
    assign layer2_outputs[1379] = ~(layer1_outputs[1502]);
    assign layer2_outputs[1380] = layer1_outputs[3525];
    assign layer2_outputs[1381] = ~((layer1_outputs[8520]) ^ (layer1_outputs[3865]));
    assign layer2_outputs[1382] = (layer1_outputs[4600]) ^ (layer1_outputs[1459]);
    assign layer2_outputs[1383] = ~(layer1_outputs[11974]);
    assign layer2_outputs[1384] = (layer1_outputs[2987]) ^ (layer1_outputs[8465]);
    assign layer2_outputs[1385] = ~(layer1_outputs[4049]);
    assign layer2_outputs[1386] = (layer1_outputs[9510]) & (layer1_outputs[3372]);
    assign layer2_outputs[1387] = ~(layer1_outputs[7133]) | (layer1_outputs[1793]);
    assign layer2_outputs[1388] = (layer1_outputs[9975]) | (layer1_outputs[9692]);
    assign layer2_outputs[1389] = layer1_outputs[11605];
    assign layer2_outputs[1390] = ~((layer1_outputs[784]) ^ (layer1_outputs[7643]));
    assign layer2_outputs[1391] = layer1_outputs[6756];
    assign layer2_outputs[1392] = ~((layer1_outputs[7017]) & (layer1_outputs[11268]));
    assign layer2_outputs[1393] = (layer1_outputs[7018]) & (layer1_outputs[5203]);
    assign layer2_outputs[1394] = ~((layer1_outputs[6719]) & (layer1_outputs[1184]));
    assign layer2_outputs[1395] = (layer1_outputs[8621]) | (layer1_outputs[10845]);
    assign layer2_outputs[1396] = ~((layer1_outputs[3947]) & (layer1_outputs[1517]));
    assign layer2_outputs[1397] = (layer1_outputs[595]) & (layer1_outputs[938]);
    assign layer2_outputs[1398] = ~((layer1_outputs[9185]) ^ (layer1_outputs[3484]));
    assign layer2_outputs[1399] = layer1_outputs[10063];
    assign layer2_outputs[1400] = layer1_outputs[2185];
    assign layer2_outputs[1401] = ~(layer1_outputs[11756]);
    assign layer2_outputs[1402] = layer1_outputs[11067];
    assign layer2_outputs[1403] = (layer1_outputs[5769]) | (layer1_outputs[9733]);
    assign layer2_outputs[1404] = ~(layer1_outputs[5228]);
    assign layer2_outputs[1405] = (layer1_outputs[7194]) | (layer1_outputs[5013]);
    assign layer2_outputs[1406] = ~(layer1_outputs[6651]) | (layer1_outputs[7121]);
    assign layer2_outputs[1407] = (layer1_outputs[9860]) ^ (layer1_outputs[1382]);
    assign layer2_outputs[1408] = ~(layer1_outputs[12430]);
    assign layer2_outputs[1409] = (layer1_outputs[11115]) ^ (layer1_outputs[11820]);
    assign layer2_outputs[1410] = (layer1_outputs[6906]) | (layer1_outputs[4527]);
    assign layer2_outputs[1411] = (layer1_outputs[9383]) ^ (layer1_outputs[5664]);
    assign layer2_outputs[1412] = (layer1_outputs[10519]) & ~(layer1_outputs[7866]);
    assign layer2_outputs[1413] = ~(layer1_outputs[4777]);
    assign layer2_outputs[1414] = ~((layer1_outputs[8435]) ^ (layer1_outputs[6072]));
    assign layer2_outputs[1415] = (layer1_outputs[724]) & ~(layer1_outputs[9879]);
    assign layer2_outputs[1416] = layer1_outputs[2761];
    assign layer2_outputs[1417] = ~(layer1_outputs[1841]);
    assign layer2_outputs[1418] = ~(layer1_outputs[11770]);
    assign layer2_outputs[1419] = ~((layer1_outputs[6060]) ^ (layer1_outputs[3842]));
    assign layer2_outputs[1420] = ~(layer1_outputs[2012]) | (layer1_outputs[6524]);
    assign layer2_outputs[1421] = ~(layer1_outputs[4126]);
    assign layer2_outputs[1422] = ~(layer1_outputs[1858]);
    assign layer2_outputs[1423] = (layer1_outputs[8768]) & ~(layer1_outputs[10394]);
    assign layer2_outputs[1424] = ~(layer1_outputs[273]);
    assign layer2_outputs[1425] = (layer1_outputs[7744]) & ~(layer1_outputs[7174]);
    assign layer2_outputs[1426] = ~((layer1_outputs[8625]) | (layer1_outputs[6194]));
    assign layer2_outputs[1427] = (layer1_outputs[12154]) & ~(layer1_outputs[8744]);
    assign layer2_outputs[1428] = ~((layer1_outputs[7023]) & (layer1_outputs[5617]));
    assign layer2_outputs[1429] = (layer1_outputs[2096]) | (layer1_outputs[1639]);
    assign layer2_outputs[1430] = (layer1_outputs[6701]) & ~(layer1_outputs[3347]);
    assign layer2_outputs[1431] = (layer1_outputs[7665]) ^ (layer1_outputs[5501]);
    assign layer2_outputs[1432] = layer1_outputs[5908];
    assign layer2_outputs[1433] = layer1_outputs[8464];
    assign layer2_outputs[1434] = layer1_outputs[4638];
    assign layer2_outputs[1435] = layer1_outputs[10194];
    assign layer2_outputs[1436] = ~(layer1_outputs[1032]);
    assign layer2_outputs[1437] = ~((layer1_outputs[4228]) ^ (layer1_outputs[11016]));
    assign layer2_outputs[1438] = layer1_outputs[11338];
    assign layer2_outputs[1439] = (layer1_outputs[7327]) & (layer1_outputs[102]);
    assign layer2_outputs[1440] = ~(layer1_outputs[4287]);
    assign layer2_outputs[1441] = (layer1_outputs[2779]) & ~(layer1_outputs[11958]);
    assign layer2_outputs[1442] = ~(layer1_outputs[8836]);
    assign layer2_outputs[1443] = layer1_outputs[12417];
    assign layer2_outputs[1444] = ~(layer1_outputs[1794]);
    assign layer2_outputs[1445] = ~(layer1_outputs[9835]);
    assign layer2_outputs[1446] = (layer1_outputs[10285]) ^ (layer1_outputs[11999]);
    assign layer2_outputs[1447] = layer1_outputs[5625];
    assign layer2_outputs[1448] = (layer1_outputs[3992]) | (layer1_outputs[441]);
    assign layer2_outputs[1449] = ~((layer1_outputs[4026]) & (layer1_outputs[11138]));
    assign layer2_outputs[1450] = (layer1_outputs[3111]) ^ (layer1_outputs[10069]);
    assign layer2_outputs[1451] = layer1_outputs[3891];
    assign layer2_outputs[1452] = ~(layer1_outputs[4125]);
    assign layer2_outputs[1453] = (layer1_outputs[64]) & ~(layer1_outputs[7083]);
    assign layer2_outputs[1454] = ~(layer1_outputs[6116]) | (layer1_outputs[6920]);
    assign layer2_outputs[1455] = layer1_outputs[8338];
    assign layer2_outputs[1456] = layer1_outputs[253];
    assign layer2_outputs[1457] = ~(layer1_outputs[3097]);
    assign layer2_outputs[1458] = ~(layer1_outputs[125]);
    assign layer2_outputs[1459] = (layer1_outputs[1137]) | (layer1_outputs[956]);
    assign layer2_outputs[1460] = ~(layer1_outputs[2416]);
    assign layer2_outputs[1461] = ~((layer1_outputs[9611]) & (layer1_outputs[345]));
    assign layer2_outputs[1462] = ~((layer1_outputs[9954]) ^ (layer1_outputs[3031]));
    assign layer2_outputs[1463] = ~((layer1_outputs[8558]) & (layer1_outputs[6222]));
    assign layer2_outputs[1464] = (layer1_outputs[85]) & (layer1_outputs[6888]);
    assign layer2_outputs[1465] = (layer1_outputs[8339]) & ~(layer1_outputs[12675]);
    assign layer2_outputs[1466] = (layer1_outputs[4073]) & ~(layer1_outputs[5340]);
    assign layer2_outputs[1467] = ~((layer1_outputs[142]) ^ (layer1_outputs[11440]));
    assign layer2_outputs[1468] = layer1_outputs[5476];
    assign layer2_outputs[1469] = ~((layer1_outputs[4211]) | (layer1_outputs[3144]));
    assign layer2_outputs[1470] = ~(layer1_outputs[9298]);
    assign layer2_outputs[1471] = ~((layer1_outputs[3731]) ^ (layer1_outputs[1094]));
    assign layer2_outputs[1472] = (layer1_outputs[8539]) | (layer1_outputs[12327]);
    assign layer2_outputs[1473] = (layer1_outputs[10811]) & ~(layer1_outputs[5150]);
    assign layer2_outputs[1474] = layer1_outputs[8945];
    assign layer2_outputs[1475] = ~(layer1_outputs[11112]);
    assign layer2_outputs[1476] = ~(layer1_outputs[835]) | (layer1_outputs[40]);
    assign layer2_outputs[1477] = layer1_outputs[524];
    assign layer2_outputs[1478] = (layer1_outputs[12477]) & ~(layer1_outputs[9508]);
    assign layer2_outputs[1479] = (layer1_outputs[2742]) & ~(layer1_outputs[5207]);
    assign layer2_outputs[1480] = ~(layer1_outputs[2395]);
    assign layer2_outputs[1481] = (layer1_outputs[8383]) & (layer1_outputs[12544]);
    assign layer2_outputs[1482] = layer1_outputs[3652];
    assign layer2_outputs[1483] = layer1_outputs[10410];
    assign layer2_outputs[1484] = layer1_outputs[5493];
    assign layer2_outputs[1485] = (layer1_outputs[3103]) ^ (layer1_outputs[7234]);
    assign layer2_outputs[1486] = (layer1_outputs[10635]) & (layer1_outputs[2225]);
    assign layer2_outputs[1487] = (layer1_outputs[11805]) & (layer1_outputs[10273]);
    assign layer2_outputs[1488] = ~(layer1_outputs[3302]);
    assign layer2_outputs[1489] = layer1_outputs[10153];
    assign layer2_outputs[1490] = (layer1_outputs[3886]) & ~(layer1_outputs[6038]);
    assign layer2_outputs[1491] = (layer1_outputs[12696]) & ~(layer1_outputs[7268]);
    assign layer2_outputs[1492] = ~((layer1_outputs[4480]) ^ (layer1_outputs[7422]));
    assign layer2_outputs[1493] = ~((layer1_outputs[11495]) ^ (layer1_outputs[7320]));
    assign layer2_outputs[1494] = (layer1_outputs[8273]) | (layer1_outputs[6567]);
    assign layer2_outputs[1495] = layer1_outputs[289];
    assign layer2_outputs[1496] = 1'b0;
    assign layer2_outputs[1497] = ~((layer1_outputs[6608]) & (layer1_outputs[8355]));
    assign layer2_outputs[1498] = ~((layer1_outputs[4369]) | (layer1_outputs[8238]));
    assign layer2_outputs[1499] = ~((layer1_outputs[11839]) ^ (layer1_outputs[1195]));
    assign layer2_outputs[1500] = layer1_outputs[6740];
    assign layer2_outputs[1501] = (layer1_outputs[9788]) ^ (layer1_outputs[5046]);
    assign layer2_outputs[1502] = (layer1_outputs[3439]) & ~(layer1_outputs[9494]);
    assign layer2_outputs[1503] = (layer1_outputs[5690]) & ~(layer1_outputs[2907]);
    assign layer2_outputs[1504] = (layer1_outputs[12506]) & ~(layer1_outputs[3668]);
    assign layer2_outputs[1505] = (layer1_outputs[9312]) ^ (layer1_outputs[10222]);
    assign layer2_outputs[1506] = ~((layer1_outputs[9720]) ^ (layer1_outputs[9813]));
    assign layer2_outputs[1507] = layer1_outputs[11358];
    assign layer2_outputs[1508] = ~(layer1_outputs[2477]);
    assign layer2_outputs[1509] = ~(layer1_outputs[4006]);
    assign layer2_outputs[1510] = ~(layer1_outputs[605]) | (layer1_outputs[645]);
    assign layer2_outputs[1511] = ~((layer1_outputs[1691]) | (layer1_outputs[4997]));
    assign layer2_outputs[1512] = ~(layer1_outputs[12018]);
    assign layer2_outputs[1513] = (layer1_outputs[5432]) & ~(layer1_outputs[1518]);
    assign layer2_outputs[1514] = layer1_outputs[10415];
    assign layer2_outputs[1515] = ~((layer1_outputs[6564]) ^ (layer1_outputs[5195]));
    assign layer2_outputs[1516] = ~(layer1_outputs[6403]);
    assign layer2_outputs[1517] = layer1_outputs[4926];
    assign layer2_outputs[1518] = ~(layer1_outputs[301]);
    assign layer2_outputs[1519] = (layer1_outputs[6197]) & ~(layer1_outputs[9336]);
    assign layer2_outputs[1520] = (layer1_outputs[3099]) ^ (layer1_outputs[12044]);
    assign layer2_outputs[1521] = ~(layer1_outputs[3837]);
    assign layer2_outputs[1522] = ~(layer1_outputs[5363]);
    assign layer2_outputs[1523] = layer1_outputs[3522];
    assign layer2_outputs[1524] = ~(layer1_outputs[3422]);
    assign layer2_outputs[1525] = (layer1_outputs[1209]) & ~(layer1_outputs[11720]);
    assign layer2_outputs[1526] = (layer1_outputs[11772]) & (layer1_outputs[4098]);
    assign layer2_outputs[1527] = ~(layer1_outputs[7897]);
    assign layer2_outputs[1528] = ~(layer1_outputs[7992]) | (layer1_outputs[5260]);
    assign layer2_outputs[1529] = (layer1_outputs[11589]) ^ (layer1_outputs[8666]);
    assign layer2_outputs[1530] = ~(layer1_outputs[10681]);
    assign layer2_outputs[1531] = ~(layer1_outputs[969]) | (layer1_outputs[9149]);
    assign layer2_outputs[1532] = (layer1_outputs[8479]) ^ (layer1_outputs[2386]);
    assign layer2_outputs[1533] = (layer1_outputs[12171]) ^ (layer1_outputs[11225]);
    assign layer2_outputs[1534] = layer1_outputs[3671];
    assign layer2_outputs[1535] = ~(layer1_outputs[2678]) | (layer1_outputs[1699]);
    assign layer2_outputs[1536] = (layer1_outputs[2280]) | (layer1_outputs[7233]);
    assign layer2_outputs[1537] = ~(layer1_outputs[10871]);
    assign layer2_outputs[1538] = ~((layer1_outputs[887]) ^ (layer1_outputs[4738]));
    assign layer2_outputs[1539] = ~(layer1_outputs[7212]);
    assign layer2_outputs[1540] = ~(layer1_outputs[1103]);
    assign layer2_outputs[1541] = ~(layer1_outputs[5022]) | (layer1_outputs[7536]);
    assign layer2_outputs[1542] = ~((layer1_outputs[6015]) ^ (layer1_outputs[12294]));
    assign layer2_outputs[1543] = layer1_outputs[2924];
    assign layer2_outputs[1544] = layer1_outputs[7458];
    assign layer2_outputs[1545] = (layer1_outputs[1519]) | (layer1_outputs[9809]);
    assign layer2_outputs[1546] = ~(layer1_outputs[9044]);
    assign layer2_outputs[1547] = (layer1_outputs[12136]) ^ (layer1_outputs[12216]);
    assign layer2_outputs[1548] = ~(layer1_outputs[4455]);
    assign layer2_outputs[1549] = ~(layer1_outputs[9788]);
    assign layer2_outputs[1550] = (layer1_outputs[6490]) ^ (layer1_outputs[8226]);
    assign layer2_outputs[1551] = ~((layer1_outputs[10103]) ^ (layer1_outputs[7536]));
    assign layer2_outputs[1552] = layer1_outputs[7153];
    assign layer2_outputs[1553] = ~(layer1_outputs[11460]) | (layer1_outputs[11153]);
    assign layer2_outputs[1554] = layer1_outputs[9909];
    assign layer2_outputs[1555] = layer1_outputs[1467];
    assign layer2_outputs[1556] = (layer1_outputs[2387]) | (layer1_outputs[6995]);
    assign layer2_outputs[1557] = ~(layer1_outputs[8460]) | (layer1_outputs[10518]);
    assign layer2_outputs[1558] = (layer1_outputs[12783]) & ~(layer1_outputs[10653]);
    assign layer2_outputs[1559] = layer1_outputs[2157];
    assign layer2_outputs[1560] = layer1_outputs[5715];
    assign layer2_outputs[1561] = ~(layer1_outputs[9017]);
    assign layer2_outputs[1562] = ~(layer1_outputs[3572]) | (layer1_outputs[6006]);
    assign layer2_outputs[1563] = ~((layer1_outputs[1221]) ^ (layer1_outputs[9927]));
    assign layer2_outputs[1564] = layer1_outputs[5506];
    assign layer2_outputs[1565] = (layer1_outputs[3711]) & ~(layer1_outputs[1097]);
    assign layer2_outputs[1566] = (layer1_outputs[3]) | (layer1_outputs[9219]);
    assign layer2_outputs[1567] = layer1_outputs[7902];
    assign layer2_outputs[1568] = ~(layer1_outputs[8237]) | (layer1_outputs[8143]);
    assign layer2_outputs[1569] = ~(layer1_outputs[2255]);
    assign layer2_outputs[1570] = ~(layer1_outputs[2637]);
    assign layer2_outputs[1571] = ~((layer1_outputs[842]) & (layer1_outputs[1575]));
    assign layer2_outputs[1572] = layer1_outputs[5544];
    assign layer2_outputs[1573] = ~(layer1_outputs[11458]);
    assign layer2_outputs[1574] = ~((layer1_outputs[5700]) | (layer1_outputs[7803]));
    assign layer2_outputs[1575] = (layer1_outputs[3973]) ^ (layer1_outputs[3557]);
    assign layer2_outputs[1576] = ~(layer1_outputs[4620]);
    assign layer2_outputs[1577] = (layer1_outputs[2437]) | (layer1_outputs[5182]);
    assign layer2_outputs[1578] = layer1_outputs[8791];
    assign layer2_outputs[1579] = ~((layer1_outputs[12651]) ^ (layer1_outputs[521]));
    assign layer2_outputs[1580] = ~(layer1_outputs[630]);
    assign layer2_outputs[1581] = layer1_outputs[4255];
    assign layer2_outputs[1582] = layer1_outputs[909];
    assign layer2_outputs[1583] = layer1_outputs[10828];
    assign layer2_outputs[1584] = layer1_outputs[1311];
    assign layer2_outputs[1585] = ~(layer1_outputs[2152]) | (layer1_outputs[1261]);
    assign layer2_outputs[1586] = (layer1_outputs[11306]) ^ (layer1_outputs[1173]);
    assign layer2_outputs[1587] = ~(layer1_outputs[10728]) | (layer1_outputs[4031]);
    assign layer2_outputs[1588] = (layer1_outputs[5274]) | (layer1_outputs[2233]);
    assign layer2_outputs[1589] = ~(layer1_outputs[4675]) | (layer1_outputs[6076]);
    assign layer2_outputs[1590] = ~((layer1_outputs[3624]) ^ (layer1_outputs[3588]));
    assign layer2_outputs[1591] = layer1_outputs[7269];
    assign layer2_outputs[1592] = layer1_outputs[2840];
    assign layer2_outputs[1593] = layer1_outputs[1665];
    assign layer2_outputs[1594] = (layer1_outputs[7235]) & ~(layer1_outputs[4355]);
    assign layer2_outputs[1595] = layer1_outputs[4681];
    assign layer2_outputs[1596] = (layer1_outputs[10280]) ^ (layer1_outputs[96]);
    assign layer2_outputs[1597] = layer1_outputs[1549];
    assign layer2_outputs[1598] = ~(layer1_outputs[6162]);
    assign layer2_outputs[1599] = ~(layer1_outputs[4617]);
    assign layer2_outputs[1600] = ~(layer1_outputs[10652]) | (layer1_outputs[10948]);
    assign layer2_outputs[1601] = (layer1_outputs[7961]) & ~(layer1_outputs[4146]);
    assign layer2_outputs[1602] = ~(layer1_outputs[3084]);
    assign layer2_outputs[1603] = ~(layer1_outputs[5707]);
    assign layer2_outputs[1604] = ~((layer1_outputs[2943]) ^ (layer1_outputs[4475]));
    assign layer2_outputs[1605] = ~(layer1_outputs[4220]);
    assign layer2_outputs[1606] = (layer1_outputs[8312]) & ~(layer1_outputs[4983]);
    assign layer2_outputs[1607] = layer1_outputs[12377];
    assign layer2_outputs[1608] = ~(layer1_outputs[4037]);
    assign layer2_outputs[1609] = (layer1_outputs[2083]) ^ (layer1_outputs[8597]);
    assign layer2_outputs[1610] = (layer1_outputs[2603]) & (layer1_outputs[3255]);
    assign layer2_outputs[1611] = ~((layer1_outputs[12119]) | (layer1_outputs[8946]));
    assign layer2_outputs[1612] = (layer1_outputs[9869]) | (layer1_outputs[7176]);
    assign layer2_outputs[1613] = ~(layer1_outputs[2721]);
    assign layer2_outputs[1614] = layer1_outputs[4184];
    assign layer2_outputs[1615] = (layer1_outputs[5259]) ^ (layer1_outputs[6430]);
    assign layer2_outputs[1616] = ~(layer1_outputs[7434]);
    assign layer2_outputs[1617] = layer1_outputs[3742];
    assign layer2_outputs[1618] = ~(layer1_outputs[8717]);
    assign layer2_outputs[1619] = layer1_outputs[5187];
    assign layer2_outputs[1620] = (layer1_outputs[1074]) & ~(layer1_outputs[4904]);
    assign layer2_outputs[1621] = (layer1_outputs[11686]) | (layer1_outputs[5135]);
    assign layer2_outputs[1622] = ~(layer1_outputs[11319]) | (layer1_outputs[6276]);
    assign layer2_outputs[1623] = layer1_outputs[3417];
    assign layer2_outputs[1624] = layer1_outputs[10942];
    assign layer2_outputs[1625] = ~((layer1_outputs[2035]) & (layer1_outputs[4317]));
    assign layer2_outputs[1626] = (layer1_outputs[8315]) & ~(layer1_outputs[9549]);
    assign layer2_outputs[1627] = ~(layer1_outputs[9148]);
    assign layer2_outputs[1628] = layer1_outputs[12338];
    assign layer2_outputs[1629] = ~(layer1_outputs[2856]) | (layer1_outputs[12010]);
    assign layer2_outputs[1630] = ~(layer1_outputs[5003]);
    assign layer2_outputs[1631] = ~(layer1_outputs[3478]);
    assign layer2_outputs[1632] = layer1_outputs[1119];
    assign layer2_outputs[1633] = ~(layer1_outputs[270]);
    assign layer2_outputs[1634] = ~((layer1_outputs[3968]) ^ (layer1_outputs[11721]));
    assign layer2_outputs[1635] = ~(layer1_outputs[7474]);
    assign layer2_outputs[1636] = ~(layer1_outputs[768]);
    assign layer2_outputs[1637] = ~(layer1_outputs[5105]);
    assign layer2_outputs[1638] = layer1_outputs[4574];
    assign layer2_outputs[1639] = ~((layer1_outputs[9451]) | (layer1_outputs[11595]));
    assign layer2_outputs[1640] = layer1_outputs[12222];
    assign layer2_outputs[1641] = layer1_outputs[1120];
    assign layer2_outputs[1642] = (layer1_outputs[11378]) ^ (layer1_outputs[7169]);
    assign layer2_outputs[1643] = (layer1_outputs[5408]) & ~(layer1_outputs[5461]);
    assign layer2_outputs[1644] = layer1_outputs[747];
    assign layer2_outputs[1645] = (layer1_outputs[9314]) & ~(layer1_outputs[6365]);
    assign layer2_outputs[1646] = 1'b1;
    assign layer2_outputs[1647] = (layer1_outputs[5907]) & ~(layer1_outputs[297]);
    assign layer2_outputs[1648] = layer1_outputs[6196];
    assign layer2_outputs[1649] = ~(layer1_outputs[132]);
    assign layer2_outputs[1650] = layer1_outputs[803];
    assign layer2_outputs[1651] = ~((layer1_outputs[6330]) & (layer1_outputs[697]));
    assign layer2_outputs[1652] = layer1_outputs[9353];
    assign layer2_outputs[1653] = ~(layer1_outputs[3193]);
    assign layer2_outputs[1654] = ~(layer1_outputs[2845]);
    assign layer2_outputs[1655] = layer1_outputs[4417];
    assign layer2_outputs[1656] = (layer1_outputs[1536]) & ~(layer1_outputs[6589]);
    assign layer2_outputs[1657] = ~((layer1_outputs[3930]) ^ (layer1_outputs[115]));
    assign layer2_outputs[1658] = (layer1_outputs[8667]) & (layer1_outputs[5889]);
    assign layer2_outputs[1659] = ~(layer1_outputs[12307]);
    assign layer2_outputs[1660] = ~(layer1_outputs[7100]);
    assign layer2_outputs[1661] = layer1_outputs[2695];
    assign layer2_outputs[1662] = ~((layer1_outputs[7144]) | (layer1_outputs[5944]));
    assign layer2_outputs[1663] = (layer1_outputs[8426]) | (layer1_outputs[2615]);
    assign layer2_outputs[1664] = (layer1_outputs[12672]) ^ (layer1_outputs[9130]);
    assign layer2_outputs[1665] = layer1_outputs[2516];
    assign layer2_outputs[1666] = ~(layer1_outputs[11089]) | (layer1_outputs[5444]);
    assign layer2_outputs[1667] = ~(layer1_outputs[11521]) | (layer1_outputs[10478]);
    assign layer2_outputs[1668] = layer1_outputs[9617];
    assign layer2_outputs[1669] = (layer1_outputs[12517]) | (layer1_outputs[5983]);
    assign layer2_outputs[1670] = layer1_outputs[11562];
    assign layer2_outputs[1671] = layer1_outputs[4565];
    assign layer2_outputs[1672] = ~(layer1_outputs[10547]);
    assign layer2_outputs[1673] = layer1_outputs[8993];
    assign layer2_outputs[1674] = (layer1_outputs[7347]) ^ (layer1_outputs[8876]);
    assign layer2_outputs[1675] = (layer1_outputs[3681]) | (layer1_outputs[8480]);
    assign layer2_outputs[1676] = (layer1_outputs[9121]) | (layer1_outputs[11825]);
    assign layer2_outputs[1677] = (layer1_outputs[5575]) | (layer1_outputs[11263]);
    assign layer2_outputs[1678] = (layer1_outputs[12139]) | (layer1_outputs[1903]);
    assign layer2_outputs[1679] = ~(layer1_outputs[159]);
    assign layer2_outputs[1680] = layer1_outputs[8069];
    assign layer2_outputs[1681] = layer1_outputs[12305];
    assign layer2_outputs[1682] = layer1_outputs[10505];
    assign layer2_outputs[1683] = ~((layer1_outputs[6589]) ^ (layer1_outputs[8928]));
    assign layer2_outputs[1684] = ~(layer1_outputs[9935]);
    assign layer2_outputs[1685] = ~((layer1_outputs[3536]) ^ (layer1_outputs[10530]));
    assign layer2_outputs[1686] = ~((layer1_outputs[3578]) | (layer1_outputs[119]));
    assign layer2_outputs[1687] = ~((layer1_outputs[12225]) ^ (layer1_outputs[4392]));
    assign layer2_outputs[1688] = layer1_outputs[1899];
    assign layer2_outputs[1689] = (layer1_outputs[6884]) ^ (layer1_outputs[12315]);
    assign layer2_outputs[1690] = layer1_outputs[7820];
    assign layer2_outputs[1691] = layer1_outputs[6220];
    assign layer2_outputs[1692] = ~(layer1_outputs[11147]);
    assign layer2_outputs[1693] = 1'b0;
    assign layer2_outputs[1694] = (layer1_outputs[4387]) & (layer1_outputs[4377]);
    assign layer2_outputs[1695] = ~(layer1_outputs[6161]);
    assign layer2_outputs[1696] = (layer1_outputs[11033]) ^ (layer1_outputs[671]);
    assign layer2_outputs[1697] = ~(layer1_outputs[12269]);
    assign layer2_outputs[1698] = (layer1_outputs[49]) & ~(layer1_outputs[6708]);
    assign layer2_outputs[1699] = layer1_outputs[5533];
    assign layer2_outputs[1700] = ~((layer1_outputs[116]) & (layer1_outputs[3709]));
    assign layer2_outputs[1701] = ~((layer1_outputs[3590]) | (layer1_outputs[33]));
    assign layer2_outputs[1702] = ~(layer1_outputs[2899]);
    assign layer2_outputs[1703] = (layer1_outputs[12411]) & ~(layer1_outputs[8659]);
    assign layer2_outputs[1704] = layer1_outputs[323];
    assign layer2_outputs[1705] = ~((layer1_outputs[2880]) | (layer1_outputs[9195]));
    assign layer2_outputs[1706] = (layer1_outputs[12481]) ^ (layer1_outputs[4360]);
    assign layer2_outputs[1707] = layer1_outputs[2514];
    assign layer2_outputs[1708] = (layer1_outputs[9262]) ^ (layer1_outputs[11173]);
    assign layer2_outputs[1709] = ~((layer1_outputs[5552]) ^ (layer1_outputs[7726]));
    assign layer2_outputs[1710] = ~(layer1_outputs[11725]) | (layer1_outputs[571]);
    assign layer2_outputs[1711] = ~(layer1_outputs[11185]);
    assign layer2_outputs[1712] = layer1_outputs[9906];
    assign layer2_outputs[1713] = layer1_outputs[10242];
    assign layer2_outputs[1714] = (layer1_outputs[4999]) & ~(layer1_outputs[5466]);
    assign layer2_outputs[1715] = ~(layer1_outputs[4979]) | (layer1_outputs[12202]);
    assign layer2_outputs[1716] = ~(layer1_outputs[5052]);
    assign layer2_outputs[1717] = (layer1_outputs[1734]) | (layer1_outputs[4494]);
    assign layer2_outputs[1718] = ~((layer1_outputs[11443]) ^ (layer1_outputs[7115]));
    assign layer2_outputs[1719] = layer1_outputs[9095];
    assign layer2_outputs[1720] = ~(layer1_outputs[11040]);
    assign layer2_outputs[1721] = layer1_outputs[7092];
    assign layer2_outputs[1722] = (layer1_outputs[5862]) | (layer1_outputs[5906]);
    assign layer2_outputs[1723] = layer1_outputs[1512];
    assign layer2_outputs[1724] = ~(layer1_outputs[3460]);
    assign layer2_outputs[1725] = layer1_outputs[4351];
    assign layer2_outputs[1726] = ~(layer1_outputs[4721]);
    assign layer2_outputs[1727] = ~(layer1_outputs[8508]);
    assign layer2_outputs[1728] = layer1_outputs[11563];
    assign layer2_outputs[1729] = layer1_outputs[5069];
    assign layer2_outputs[1730] = layer1_outputs[7667];
    assign layer2_outputs[1731] = ~((layer1_outputs[4094]) ^ (layer1_outputs[4928]));
    assign layer2_outputs[1732] = ~(layer1_outputs[8698]);
    assign layer2_outputs[1733] = (layer1_outputs[8654]) ^ (layer1_outputs[5738]);
    assign layer2_outputs[1734] = ~(layer1_outputs[12690]);
    assign layer2_outputs[1735] = ~(layer1_outputs[9620]);
    assign layer2_outputs[1736] = 1'b0;
    assign layer2_outputs[1737] = ~(layer1_outputs[1454]) | (layer1_outputs[3825]);
    assign layer2_outputs[1738] = layer1_outputs[3556];
    assign layer2_outputs[1739] = ~(layer1_outputs[9071]) | (layer1_outputs[6266]);
    assign layer2_outputs[1740] = ~(layer1_outputs[12069]) | (layer1_outputs[7437]);
    assign layer2_outputs[1741] = ~((layer1_outputs[1873]) & (layer1_outputs[5012]));
    assign layer2_outputs[1742] = layer1_outputs[5263];
    assign layer2_outputs[1743] = ~((layer1_outputs[10114]) ^ (layer1_outputs[12152]));
    assign layer2_outputs[1744] = 1'b1;
    assign layer2_outputs[1745] = ~(layer1_outputs[4377]);
    assign layer2_outputs[1746] = layer1_outputs[8866];
    assign layer2_outputs[1747] = ~(layer1_outputs[5736]);
    assign layer2_outputs[1748] = ~((layer1_outputs[9525]) | (layer1_outputs[11938]));
    assign layer2_outputs[1749] = ~((layer1_outputs[12047]) ^ (layer1_outputs[3024]));
    assign layer2_outputs[1750] = layer1_outputs[8792];
    assign layer2_outputs[1751] = ~(layer1_outputs[4056]) | (layer1_outputs[328]);
    assign layer2_outputs[1752] = layer1_outputs[9474];
    assign layer2_outputs[1753] = layer1_outputs[4964];
    assign layer2_outputs[1754] = ~(layer1_outputs[10135]) | (layer1_outputs[2176]);
    assign layer2_outputs[1755] = ~(layer1_outputs[4448]);
    assign layer2_outputs[1756] = (layer1_outputs[2410]) & ~(layer1_outputs[3398]);
    assign layer2_outputs[1757] = ~(layer1_outputs[1495]);
    assign layer2_outputs[1758] = ~((layer1_outputs[7318]) & (layer1_outputs[8887]));
    assign layer2_outputs[1759] = ~(layer1_outputs[1802]);
    assign layer2_outputs[1760] = layer1_outputs[7468];
    assign layer2_outputs[1761] = ~((layer1_outputs[11879]) ^ (layer1_outputs[6769]));
    assign layer2_outputs[1762] = ~((layer1_outputs[4075]) | (layer1_outputs[10527]));
    assign layer2_outputs[1763] = (layer1_outputs[5092]) & (layer1_outputs[9656]);
    assign layer2_outputs[1764] = (layer1_outputs[5865]) | (layer1_outputs[409]);
    assign layer2_outputs[1765] = layer1_outputs[5625];
    assign layer2_outputs[1766] = layer1_outputs[2813];
    assign layer2_outputs[1767] = ~(layer1_outputs[3775]);
    assign layer2_outputs[1768] = ~(layer1_outputs[9952]);
    assign layer2_outputs[1769] = ~(layer1_outputs[9685]);
    assign layer2_outputs[1770] = layer1_outputs[313];
    assign layer2_outputs[1771] = ~((layer1_outputs[11069]) ^ (layer1_outputs[10956]));
    assign layer2_outputs[1772] = ~((layer1_outputs[11687]) ^ (layer1_outputs[11774]));
    assign layer2_outputs[1773] = layer1_outputs[7025];
    assign layer2_outputs[1774] = (layer1_outputs[427]) & (layer1_outputs[11527]);
    assign layer2_outputs[1775] = (layer1_outputs[4576]) | (layer1_outputs[6082]);
    assign layer2_outputs[1776] = ~(layer1_outputs[8200]) | (layer1_outputs[9968]);
    assign layer2_outputs[1777] = ~(layer1_outputs[7472]);
    assign layer2_outputs[1778] = ~(layer1_outputs[10070]);
    assign layer2_outputs[1779] = ~(layer1_outputs[7142]);
    assign layer2_outputs[1780] = ~((layer1_outputs[2786]) ^ (layer1_outputs[2361]));
    assign layer2_outputs[1781] = layer1_outputs[9090];
    assign layer2_outputs[1782] = layer1_outputs[2862];
    assign layer2_outputs[1783] = ~(layer1_outputs[9644]);
    assign layer2_outputs[1784] = ~((layer1_outputs[5126]) ^ (layer1_outputs[836]));
    assign layer2_outputs[1785] = ~(layer1_outputs[6766]);
    assign layer2_outputs[1786] = (layer1_outputs[10848]) & ~(layer1_outputs[9480]);
    assign layer2_outputs[1787] = ~(layer1_outputs[8977]);
    assign layer2_outputs[1788] = ~((layer1_outputs[9756]) & (layer1_outputs[6909]));
    assign layer2_outputs[1789] = ~(layer1_outputs[1436]);
    assign layer2_outputs[1790] = layer1_outputs[7102];
    assign layer2_outputs[1791] = ~((layer1_outputs[8275]) | (layer1_outputs[1304]));
    assign layer2_outputs[1792] = ~(layer1_outputs[4310]) | (layer1_outputs[3078]);
    assign layer2_outputs[1793] = ~((layer1_outputs[1789]) | (layer1_outputs[5024]));
    assign layer2_outputs[1794] = ~((layer1_outputs[11402]) ^ (layer1_outputs[6081]));
    assign layer2_outputs[1795] = ~((layer1_outputs[2442]) ^ (layer1_outputs[2663]));
    assign layer2_outputs[1796] = (layer1_outputs[7082]) & ~(layer1_outputs[10738]);
    assign layer2_outputs[1797] = layer1_outputs[10762];
    assign layer2_outputs[1798] = ~(layer1_outputs[11546]) | (layer1_outputs[8648]);
    assign layer2_outputs[1799] = ~((layer1_outputs[12686]) & (layer1_outputs[11716]));
    assign layer2_outputs[1800] = ~((layer1_outputs[4980]) ^ (layer1_outputs[9636]));
    assign layer2_outputs[1801] = ~(layer1_outputs[4934]);
    assign layer2_outputs[1802] = ~(layer1_outputs[3846]);
    assign layer2_outputs[1803] = ~((layer1_outputs[10760]) ^ (layer1_outputs[9377]));
    assign layer2_outputs[1804] = (layer1_outputs[6594]) & (layer1_outputs[7208]);
    assign layer2_outputs[1805] = layer1_outputs[1469];
    assign layer2_outputs[1806] = (layer1_outputs[113]) & (layer1_outputs[2952]);
    assign layer2_outputs[1807] = (layer1_outputs[3450]) ^ (layer1_outputs[8936]);
    assign layer2_outputs[1808] = layer1_outputs[7123];
    assign layer2_outputs[1809] = ~((layer1_outputs[499]) ^ (layer1_outputs[10043]));
    assign layer2_outputs[1810] = (layer1_outputs[4788]) ^ (layer1_outputs[7238]);
    assign layer2_outputs[1811] = ~(layer1_outputs[12371]) | (layer1_outputs[3286]);
    assign layer2_outputs[1812] = (layer1_outputs[3538]) & (layer1_outputs[8681]);
    assign layer2_outputs[1813] = layer1_outputs[3745];
    assign layer2_outputs[1814] = layer1_outputs[5143];
    assign layer2_outputs[1815] = layer1_outputs[6172];
    assign layer2_outputs[1816] = (layer1_outputs[1525]) ^ (layer1_outputs[5032]);
    assign layer2_outputs[1817] = layer1_outputs[10193];
    assign layer2_outputs[1818] = ~((layer1_outputs[1364]) & (layer1_outputs[643]));
    assign layer2_outputs[1819] = ~(layer1_outputs[11153]);
    assign layer2_outputs[1820] = 1'b0;
    assign layer2_outputs[1821] = layer1_outputs[11561];
    assign layer2_outputs[1822] = (layer1_outputs[9007]) & ~(layer1_outputs[4763]);
    assign layer2_outputs[1823] = ~(layer1_outputs[7629]);
    assign layer2_outputs[1824] = (layer1_outputs[10870]) & ~(layer1_outputs[7485]);
    assign layer2_outputs[1825] = (layer1_outputs[7690]) & (layer1_outputs[3302]);
    assign layer2_outputs[1826] = ~(layer1_outputs[10251]);
    assign layer2_outputs[1827] = (layer1_outputs[7258]) & (layer1_outputs[8564]);
    assign layer2_outputs[1828] = ~(layer1_outputs[4217]);
    assign layer2_outputs[1829] = (layer1_outputs[1530]) & ~(layer1_outputs[7224]);
    assign layer2_outputs[1830] = ~((layer1_outputs[3295]) ^ (layer1_outputs[6271]));
    assign layer2_outputs[1831] = layer1_outputs[8737];
    assign layer2_outputs[1832] = ~((layer1_outputs[3356]) & (layer1_outputs[7321]));
    assign layer2_outputs[1833] = 1'b1;
    assign layer2_outputs[1834] = ~(layer1_outputs[11159]);
    assign layer2_outputs[1835] = ~(layer1_outputs[7222]) | (layer1_outputs[9727]);
    assign layer2_outputs[1836] = ~(layer1_outputs[6443]) | (layer1_outputs[4129]);
    assign layer2_outputs[1837] = ~(layer1_outputs[3182]) | (layer1_outputs[5490]);
    assign layer2_outputs[1838] = ~(layer1_outputs[242]);
    assign layer2_outputs[1839] = ~((layer1_outputs[2060]) & (layer1_outputs[4661]));
    assign layer2_outputs[1840] = ~(layer1_outputs[410]);
    assign layer2_outputs[1841] = layer1_outputs[6894];
    assign layer2_outputs[1842] = layer1_outputs[8849];
    assign layer2_outputs[1843] = (layer1_outputs[11971]) & (layer1_outputs[8938]);
    assign layer2_outputs[1844] = layer1_outputs[6294];
    assign layer2_outputs[1845] = layer1_outputs[3892];
    assign layer2_outputs[1846] = ~(layer1_outputs[4215]);
    assign layer2_outputs[1847] = (layer1_outputs[11512]) & ~(layer1_outputs[11965]);
    assign layer2_outputs[1848] = (layer1_outputs[11262]) & ~(layer1_outputs[678]);
    assign layer2_outputs[1849] = ~((layer1_outputs[11327]) ^ (layer1_outputs[7035]));
    assign layer2_outputs[1850] = ~((layer1_outputs[4631]) ^ (layer1_outputs[5093]));
    assign layer2_outputs[1851] = ~((layer1_outputs[10734]) & (layer1_outputs[3567]));
    assign layer2_outputs[1852] = ~(layer1_outputs[12051]) | (layer1_outputs[3736]);
    assign layer2_outputs[1853] = layer1_outputs[6769];
    assign layer2_outputs[1854] = (layer1_outputs[11591]) & (layer1_outputs[2579]);
    assign layer2_outputs[1855] = ~(layer1_outputs[620]);
    assign layer2_outputs[1856] = (layer1_outputs[9072]) ^ (layer1_outputs[10788]);
    assign layer2_outputs[1857] = ~(layer1_outputs[12483]);
    assign layer2_outputs[1858] = 1'b1;
    assign layer2_outputs[1859] = ~((layer1_outputs[12336]) ^ (layer1_outputs[10099]));
    assign layer2_outputs[1860] = ~(layer1_outputs[6218]) | (layer1_outputs[11335]);
    assign layer2_outputs[1861] = layer1_outputs[217];
    assign layer2_outputs[1862] = ~((layer1_outputs[12617]) | (layer1_outputs[9781]));
    assign layer2_outputs[1863] = layer1_outputs[4783];
    assign layer2_outputs[1864] = layer1_outputs[8501];
    assign layer2_outputs[1865] = (layer1_outputs[1243]) & ~(layer1_outputs[9166]);
    assign layer2_outputs[1866] = (layer1_outputs[4740]) ^ (layer1_outputs[447]);
    assign layer2_outputs[1867] = ~(layer1_outputs[6514]) | (layer1_outputs[7205]);
    assign layer2_outputs[1868] = layer1_outputs[1829];
    assign layer2_outputs[1869] = ~(layer1_outputs[12688]);
    assign layer2_outputs[1870] = ~(layer1_outputs[5589]);
    assign layer2_outputs[1871] = layer1_outputs[2134];
    assign layer2_outputs[1872] = ~(layer1_outputs[9439]);
    assign layer2_outputs[1873] = layer1_outputs[10555];
    assign layer2_outputs[1874] = (layer1_outputs[7856]) ^ (layer1_outputs[1172]);
    assign layer2_outputs[1875] = ~(layer1_outputs[7435]) | (layer1_outputs[4417]);
    assign layer2_outputs[1876] = ~((layer1_outputs[4406]) | (layer1_outputs[380]));
    assign layer2_outputs[1877] = (layer1_outputs[1844]) & ~(layer1_outputs[4547]);
    assign layer2_outputs[1878] = layer1_outputs[11679];
    assign layer2_outputs[1879] = ~((layer1_outputs[3252]) & (layer1_outputs[3589]));
    assign layer2_outputs[1880] = (layer1_outputs[9232]) & ~(layer1_outputs[6561]);
    assign layer2_outputs[1881] = layer1_outputs[6395];
    assign layer2_outputs[1882] = (layer1_outputs[10909]) | (layer1_outputs[12676]);
    assign layer2_outputs[1883] = (layer1_outputs[9164]) & ~(layer1_outputs[10597]);
    assign layer2_outputs[1884] = (layer1_outputs[5615]) ^ (layer1_outputs[1619]);
    assign layer2_outputs[1885] = ~(layer1_outputs[1332]);
    assign layer2_outputs[1886] = layer1_outputs[3694];
    assign layer2_outputs[1887] = (layer1_outputs[3983]) & ~(layer1_outputs[2332]);
    assign layer2_outputs[1888] = (layer1_outputs[3114]) ^ (layer1_outputs[9039]);
    assign layer2_outputs[1889] = ~(layer1_outputs[3684]);
    assign layer2_outputs[1890] = layer1_outputs[12158];
    assign layer2_outputs[1891] = ~(layer1_outputs[6614]);
    assign layer2_outputs[1892] = ~(layer1_outputs[8186]) | (layer1_outputs[4192]);
    assign layer2_outputs[1893] = ~((layer1_outputs[7921]) | (layer1_outputs[3129]));
    assign layer2_outputs[1894] = ~((layer1_outputs[9367]) ^ (layer1_outputs[9272]));
    assign layer2_outputs[1895] = ~(layer1_outputs[7751]);
    assign layer2_outputs[1896] = layer1_outputs[3577];
    assign layer2_outputs[1897] = layer1_outputs[3258];
    assign layer2_outputs[1898] = ~((layer1_outputs[7058]) ^ (layer1_outputs[3241]));
    assign layer2_outputs[1899] = ~(layer1_outputs[1408]) | (layer1_outputs[11656]);
    assign layer2_outputs[1900] = (layer1_outputs[9972]) & ~(layer1_outputs[10858]);
    assign layer2_outputs[1901] = (layer1_outputs[6131]) ^ (layer1_outputs[4770]);
    assign layer2_outputs[1902] = ~(layer1_outputs[11519]);
    assign layer2_outputs[1903] = ~(layer1_outputs[11551]);
    assign layer2_outputs[1904] = layer1_outputs[12261];
    assign layer2_outputs[1905] = (layer1_outputs[9590]) & ~(layer1_outputs[2319]);
    assign layer2_outputs[1906] = (layer1_outputs[5393]) ^ (layer1_outputs[8892]);
    assign layer2_outputs[1907] = layer1_outputs[7270];
    assign layer2_outputs[1908] = layer1_outputs[8897];
    assign layer2_outputs[1909] = ~((layer1_outputs[487]) | (layer1_outputs[1800]));
    assign layer2_outputs[1910] = ~((layer1_outputs[11453]) & (layer1_outputs[10573]));
    assign layer2_outputs[1911] = ~(layer1_outputs[4622]);
    assign layer2_outputs[1912] = ~(layer1_outputs[6918]);
    assign layer2_outputs[1913] = layer1_outputs[2164];
    assign layer2_outputs[1914] = layer1_outputs[5669];
    assign layer2_outputs[1915] = ~(layer1_outputs[9161]);
    assign layer2_outputs[1916] = 1'b1;
    assign layer2_outputs[1917] = (layer1_outputs[10020]) & ~(layer1_outputs[2231]);
    assign layer2_outputs[1918] = ~(layer1_outputs[10278]);
    assign layer2_outputs[1919] = ~(layer1_outputs[267]);
    assign layer2_outputs[1920] = ~(layer1_outputs[11114]) | (layer1_outputs[6898]);
    assign layer2_outputs[1921] = layer1_outputs[4174];
    assign layer2_outputs[1922] = layer1_outputs[6862];
    assign layer2_outputs[1923] = layer1_outputs[559];
    assign layer2_outputs[1924] = (layer1_outputs[2616]) ^ (layer1_outputs[354]);
    assign layer2_outputs[1925] = layer1_outputs[1053];
    assign layer2_outputs[1926] = ~((layer1_outputs[9299]) & (layer1_outputs[3206]));
    assign layer2_outputs[1927] = layer1_outputs[2037];
    assign layer2_outputs[1928] = layer1_outputs[10894];
    assign layer2_outputs[1929] = layer1_outputs[12241];
    assign layer2_outputs[1930] = ~((layer1_outputs[5927]) | (layer1_outputs[2018]));
    assign layer2_outputs[1931] = (layer1_outputs[6276]) & (layer1_outputs[3502]);
    assign layer2_outputs[1932] = (layer1_outputs[8448]) & ~(layer1_outputs[7404]);
    assign layer2_outputs[1933] = (layer1_outputs[2134]) & ~(layer1_outputs[8118]);
    assign layer2_outputs[1934] = ~(layer1_outputs[1004]);
    assign layer2_outputs[1935] = ~(layer1_outputs[3270]);
    assign layer2_outputs[1936] = (layer1_outputs[6038]) & ~(layer1_outputs[4564]);
    assign layer2_outputs[1937] = layer1_outputs[1101];
    assign layer2_outputs[1938] = (layer1_outputs[3083]) & ~(layer1_outputs[4941]);
    assign layer2_outputs[1939] = ~(layer1_outputs[4220]);
    assign layer2_outputs[1940] = ~(layer1_outputs[6469]);
    assign layer2_outputs[1941] = layer1_outputs[2596];
    assign layer2_outputs[1942] = layer1_outputs[5942];
    assign layer2_outputs[1943] = (layer1_outputs[871]) & ~(layer1_outputs[10997]);
    assign layer2_outputs[1944] = ~(layer1_outputs[2305]) | (layer1_outputs[11788]);
    assign layer2_outputs[1945] = layer1_outputs[1255];
    assign layer2_outputs[1946] = ~(layer1_outputs[11215]) | (layer1_outputs[8177]);
    assign layer2_outputs[1947] = (layer1_outputs[4002]) | (layer1_outputs[8378]);
    assign layer2_outputs[1948] = ~((layer1_outputs[9222]) ^ (layer1_outputs[720]));
    assign layer2_outputs[1949] = layer1_outputs[8036];
    assign layer2_outputs[1950] = (layer1_outputs[8483]) & ~(layer1_outputs[3662]);
    assign layer2_outputs[1951] = ~(layer1_outputs[4165]);
    assign layer2_outputs[1952] = ~((layer1_outputs[3808]) ^ (layer1_outputs[2460]));
    assign layer2_outputs[1953] = ~((layer1_outputs[3048]) | (layer1_outputs[5453]));
    assign layer2_outputs[1954] = (layer1_outputs[5292]) & ~(layer1_outputs[3762]);
    assign layer2_outputs[1955] = ~(layer1_outputs[10577]);
    assign layer2_outputs[1956] = layer1_outputs[2116];
    assign layer2_outputs[1957] = ~(layer1_outputs[8761]);
    assign layer2_outputs[1958] = ~(layer1_outputs[4382]) | (layer1_outputs[12357]);
    assign layer2_outputs[1959] = (layer1_outputs[2890]) & (layer1_outputs[2527]);
    assign layer2_outputs[1960] = (layer1_outputs[8604]) & ~(layer1_outputs[2591]);
    assign layer2_outputs[1961] = ~(layer1_outputs[10216]);
    assign layer2_outputs[1962] = ~(layer1_outputs[4947]);
    assign layer2_outputs[1963] = ~(layer1_outputs[12345]);
    assign layer2_outputs[1964] = layer1_outputs[2895];
    assign layer2_outputs[1965] = ~(layer1_outputs[8579]);
    assign layer2_outputs[1966] = ~(layer1_outputs[2254]);
    assign layer2_outputs[1967] = (layer1_outputs[3810]) & ~(layer1_outputs[5110]);
    assign layer2_outputs[1968] = layer1_outputs[106];
    assign layer2_outputs[1969] = ~(layer1_outputs[4359]);
    assign layer2_outputs[1970] = ~((layer1_outputs[4818]) | (layer1_outputs[11069]));
    assign layer2_outputs[1971] = layer1_outputs[9538];
    assign layer2_outputs[1972] = (layer1_outputs[1280]) & ~(layer1_outputs[4549]);
    assign layer2_outputs[1973] = ~(layer1_outputs[7751]);
    assign layer2_outputs[1974] = ~(layer1_outputs[4759]) | (layer1_outputs[6451]);
    assign layer2_outputs[1975] = (layer1_outputs[731]) & (layer1_outputs[12767]);
    assign layer2_outputs[1976] = layer1_outputs[11682];
    assign layer2_outputs[1977] = ~(layer1_outputs[3214]);
    assign layer2_outputs[1978] = ~(layer1_outputs[6289]);
    assign layer2_outputs[1979] = ~((layer1_outputs[270]) & (layer1_outputs[8360]));
    assign layer2_outputs[1980] = ~(layer1_outputs[3900]);
    assign layer2_outputs[1981] = layer1_outputs[4337];
    assign layer2_outputs[1982] = layer1_outputs[8347];
    assign layer2_outputs[1983] = ~(layer1_outputs[7719]);
    assign layer2_outputs[1984] = ~((layer1_outputs[2183]) | (layer1_outputs[5264]));
    assign layer2_outputs[1985] = ~(layer1_outputs[1313]);
    assign layer2_outputs[1986] = ~(layer1_outputs[12177]);
    assign layer2_outputs[1987] = layer1_outputs[9395];
    assign layer2_outputs[1988] = layer1_outputs[7162];
    assign layer2_outputs[1989] = layer1_outputs[5106];
    assign layer2_outputs[1990] = layer1_outputs[9369];
    assign layer2_outputs[1991] = (layer1_outputs[4392]) | (layer1_outputs[2449]);
    assign layer2_outputs[1992] = ~((layer1_outputs[3839]) & (layer1_outputs[12785]));
    assign layer2_outputs[1993] = ~(layer1_outputs[12130]);
    assign layer2_outputs[1994] = layer1_outputs[5962];
    assign layer2_outputs[1995] = layer1_outputs[1558];
    assign layer2_outputs[1996] = ~((layer1_outputs[5331]) | (layer1_outputs[2959]));
    assign layer2_outputs[1997] = ~((layer1_outputs[2383]) & (layer1_outputs[8348]));
    assign layer2_outputs[1998] = (layer1_outputs[1856]) & ~(layer1_outputs[9920]);
    assign layer2_outputs[1999] = ~(layer1_outputs[6643]);
    assign layer2_outputs[2000] = (layer1_outputs[3972]) | (layer1_outputs[12405]);
    assign layer2_outputs[2001] = ~((layer1_outputs[7330]) ^ (layer1_outputs[8851]));
    assign layer2_outputs[2002] = ~(layer1_outputs[8049]);
    assign layer2_outputs[2003] = ~((layer1_outputs[7477]) ^ (layer1_outputs[2396]));
    assign layer2_outputs[2004] = (layer1_outputs[5695]) ^ (layer1_outputs[5422]);
    assign layer2_outputs[2005] = layer1_outputs[10998];
    assign layer2_outputs[2006] = ~((layer1_outputs[11041]) | (layer1_outputs[187]));
    assign layer2_outputs[2007] = ~((layer1_outputs[4122]) ^ (layer1_outputs[7819]));
    assign layer2_outputs[2008] = (layer1_outputs[9080]) ^ (layer1_outputs[3145]);
    assign layer2_outputs[2009] = layer1_outputs[2457];
    assign layer2_outputs[2010] = layer1_outputs[107];
    assign layer2_outputs[2011] = (layer1_outputs[4824]) ^ (layer1_outputs[7142]);
    assign layer2_outputs[2012] = (layer1_outputs[9904]) | (layer1_outputs[6973]);
    assign layer2_outputs[2013] = ~(layer1_outputs[4294]) | (layer1_outputs[2689]);
    assign layer2_outputs[2014] = ~((layer1_outputs[7606]) | (layer1_outputs[7634]));
    assign layer2_outputs[2015] = (layer1_outputs[5637]) & ~(layer1_outputs[161]);
    assign layer2_outputs[2016] = ~((layer1_outputs[3459]) ^ (layer1_outputs[11057]));
    assign layer2_outputs[2017] = ~((layer1_outputs[2049]) ^ (layer1_outputs[7851]));
    assign layer2_outputs[2018] = 1'b1;
    assign layer2_outputs[2019] = ~(layer1_outputs[548]);
    assign layer2_outputs[2020] = (layer1_outputs[4881]) ^ (layer1_outputs[333]);
    assign layer2_outputs[2021] = ~(layer1_outputs[6940]);
    assign layer2_outputs[2022] = ~(layer1_outputs[1051]);
    assign layer2_outputs[2023] = ~((layer1_outputs[3316]) | (layer1_outputs[4401]));
    assign layer2_outputs[2024] = ~((layer1_outputs[555]) | (layer1_outputs[209]));
    assign layer2_outputs[2025] = layer1_outputs[6024];
    assign layer2_outputs[2026] = layer1_outputs[1920];
    assign layer2_outputs[2027] = (layer1_outputs[3523]) ^ (layer1_outputs[258]);
    assign layer2_outputs[2028] = ~(layer1_outputs[4020]);
    assign layer2_outputs[2029] = (layer1_outputs[8116]) & ~(layer1_outputs[5654]);
    assign layer2_outputs[2030] = (layer1_outputs[5701]) & ~(layer1_outputs[9147]);
    assign layer2_outputs[2031] = ~(layer1_outputs[350]);
    assign layer2_outputs[2032] = ~(layer1_outputs[6951]);
    assign layer2_outputs[2033] = layer1_outputs[5073];
    assign layer2_outputs[2034] = ~(layer1_outputs[10378]) | (layer1_outputs[1959]);
    assign layer2_outputs[2035] = layer1_outputs[1046];
    assign layer2_outputs[2036] = layer1_outputs[3586];
    assign layer2_outputs[2037] = layer1_outputs[94];
    assign layer2_outputs[2038] = ~((layer1_outputs[2178]) & (layer1_outputs[2292]));
    assign layer2_outputs[2039] = layer1_outputs[8915];
    assign layer2_outputs[2040] = ~(layer1_outputs[9439]);
    assign layer2_outputs[2041] = (layer1_outputs[5690]) & ~(layer1_outputs[9176]);
    assign layer2_outputs[2042] = (layer1_outputs[3024]) ^ (layer1_outputs[10006]);
    assign layer2_outputs[2043] = ~(layer1_outputs[12409]);
    assign layer2_outputs[2044] = ~(layer1_outputs[5881]) | (layer1_outputs[3600]);
    assign layer2_outputs[2045] = (layer1_outputs[1175]) & ~(layer1_outputs[4290]);
    assign layer2_outputs[2046] = layer1_outputs[6310];
    assign layer2_outputs[2047] = ~(layer1_outputs[8480]) | (layer1_outputs[10250]);
    assign layer2_outputs[2048] = layer1_outputs[12685];
    assign layer2_outputs[2049] = layer1_outputs[3552];
    assign layer2_outputs[2050] = layer1_outputs[4599];
    assign layer2_outputs[2051] = ~(layer1_outputs[12194]);
    assign layer2_outputs[2052] = layer1_outputs[7281];
    assign layer2_outputs[2053] = (layer1_outputs[10712]) & ~(layer1_outputs[442]);
    assign layer2_outputs[2054] = ~(layer1_outputs[8071]);
    assign layer2_outputs[2055] = (layer1_outputs[7057]) ^ (layer1_outputs[2548]);
    assign layer2_outputs[2056] = layer1_outputs[5987];
    assign layer2_outputs[2057] = ~(layer1_outputs[3291]);
    assign layer2_outputs[2058] = (layer1_outputs[12280]) | (layer1_outputs[10961]);
    assign layer2_outputs[2059] = ~(layer1_outputs[11121]);
    assign layer2_outputs[2060] = (layer1_outputs[3947]) & ~(layer1_outputs[3260]);
    assign layer2_outputs[2061] = layer1_outputs[10698];
    assign layer2_outputs[2062] = ~(layer1_outputs[6708]);
    assign layer2_outputs[2063] = ~(layer1_outputs[11614]);
    assign layer2_outputs[2064] = ~(layer1_outputs[5680]);
    assign layer2_outputs[2065] = ~(layer1_outputs[6221]);
    assign layer2_outputs[2066] = (layer1_outputs[6945]) | (layer1_outputs[5707]);
    assign layer2_outputs[2067] = (layer1_outputs[6978]) ^ (layer1_outputs[6604]);
    assign layer2_outputs[2068] = layer1_outputs[3910];
    assign layer2_outputs[2069] = ~(layer1_outputs[2758]);
    assign layer2_outputs[2070] = ~((layer1_outputs[1464]) ^ (layer1_outputs[2533]));
    assign layer2_outputs[2071] = (layer1_outputs[6198]) ^ (layer1_outputs[8540]);
    assign layer2_outputs[2072] = ~(layer1_outputs[8462]);
    assign layer2_outputs[2073] = layer1_outputs[11356];
    assign layer2_outputs[2074] = ~(layer1_outputs[3144]);
    assign layer2_outputs[2075] = layer1_outputs[11850];
    assign layer2_outputs[2076] = layer1_outputs[7656];
    assign layer2_outputs[2077] = layer1_outputs[12341];
    assign layer2_outputs[2078] = ~((layer1_outputs[9790]) & (layer1_outputs[875]));
    assign layer2_outputs[2079] = (layer1_outputs[7819]) & ~(layer1_outputs[916]);
    assign layer2_outputs[2080] = layer1_outputs[9101];
    assign layer2_outputs[2081] = layer1_outputs[8918];
    assign layer2_outputs[2082] = ~(layer1_outputs[4858]);
    assign layer2_outputs[2083] = layer1_outputs[2182];
    assign layer2_outputs[2084] = (layer1_outputs[5385]) | (layer1_outputs[652]);
    assign layer2_outputs[2085] = layer1_outputs[3288];
    assign layer2_outputs[2086] = (layer1_outputs[5032]) & ~(layer1_outputs[7762]);
    assign layer2_outputs[2087] = ~(layer1_outputs[3772]);
    assign layer2_outputs[2088] = ~(layer1_outputs[902]);
    assign layer2_outputs[2089] = ~((layer1_outputs[10108]) & (layer1_outputs[11277]));
    assign layer2_outputs[2090] = ~(layer1_outputs[5418]);
    assign layer2_outputs[2091] = ~((layer1_outputs[2743]) ^ (layer1_outputs[10474]));
    assign layer2_outputs[2092] = ~(layer1_outputs[9515]) | (layer1_outputs[6543]);
    assign layer2_outputs[2093] = ~(layer1_outputs[3130]);
    assign layer2_outputs[2094] = ~((layer1_outputs[4141]) & (layer1_outputs[231]));
    assign layer2_outputs[2095] = 1'b1;
    assign layer2_outputs[2096] = layer1_outputs[1339];
    assign layer2_outputs[2097] = ~((layer1_outputs[8946]) ^ (layer1_outputs[6209]));
    assign layer2_outputs[2098] = (layer1_outputs[12221]) & ~(layer1_outputs[10507]);
    assign layer2_outputs[2099] = (layer1_outputs[2221]) ^ (layer1_outputs[6573]);
    assign layer2_outputs[2100] = ~((layer1_outputs[8221]) ^ (layer1_outputs[3527]));
    assign layer2_outputs[2101] = ~(layer1_outputs[5047]);
    assign layer2_outputs[2102] = ~((layer1_outputs[4766]) ^ (layer1_outputs[1671]));
    assign layer2_outputs[2103] = layer1_outputs[6356];
    assign layer2_outputs[2104] = ~((layer1_outputs[9278]) & (layer1_outputs[6811]));
    assign layer2_outputs[2105] = ~(layer1_outputs[5313]) | (layer1_outputs[3924]);
    assign layer2_outputs[2106] = layer1_outputs[2318];
    assign layer2_outputs[2107] = layer1_outputs[1385];
    assign layer2_outputs[2108] = (layer1_outputs[4624]) & (layer1_outputs[9739]);
    assign layer2_outputs[2109] = layer1_outputs[11177];
    assign layer2_outputs[2110] = (layer1_outputs[10464]) & ~(layer1_outputs[6009]);
    assign layer2_outputs[2111] = ~(layer1_outputs[5498]) | (layer1_outputs[2625]);
    assign layer2_outputs[2112] = layer1_outputs[6744];
    assign layer2_outputs[2113] = ~(layer1_outputs[4301]);
    assign layer2_outputs[2114] = ~(layer1_outputs[12691]) | (layer1_outputs[10991]);
    assign layer2_outputs[2115] = (layer1_outputs[1443]) & ~(layer1_outputs[5366]);
    assign layer2_outputs[2116] = ~((layer1_outputs[9717]) ^ (layer1_outputs[7965]));
    assign layer2_outputs[2117] = layer1_outputs[11399];
    assign layer2_outputs[2118] = ~(layer1_outputs[8913]) | (layer1_outputs[4933]);
    assign layer2_outputs[2119] = ~((layer1_outputs[7879]) | (layer1_outputs[1722]));
    assign layer2_outputs[2120] = layer1_outputs[241];
    assign layer2_outputs[2121] = layer1_outputs[464];
    assign layer2_outputs[2122] = layer1_outputs[4005];
    assign layer2_outputs[2123] = 1'b1;
    assign layer2_outputs[2124] = ~(layer1_outputs[10319]);
    assign layer2_outputs[2125] = ~((layer1_outputs[10896]) | (layer1_outputs[456]));
    assign layer2_outputs[2126] = ~((layer1_outputs[4198]) ^ (layer1_outputs[6219]));
    assign layer2_outputs[2127] = (layer1_outputs[6542]) | (layer1_outputs[7953]);
    assign layer2_outputs[2128] = (layer1_outputs[9794]) & (layer1_outputs[5832]);
    assign layer2_outputs[2129] = ~(layer1_outputs[2555]);
    assign layer2_outputs[2130] = layer1_outputs[12124];
    assign layer2_outputs[2131] = ~((layer1_outputs[1684]) ^ (layer1_outputs[998]));
    assign layer2_outputs[2132] = ~((layer1_outputs[9366]) | (layer1_outputs[12530]));
    assign layer2_outputs[2133] = (layer1_outputs[10831]) & ~(layer1_outputs[10496]);
    assign layer2_outputs[2134] = ~((layer1_outputs[9657]) & (layer1_outputs[4843]));
    assign layer2_outputs[2135] = (layer1_outputs[5454]) & ~(layer1_outputs[5579]);
    assign layer2_outputs[2136] = layer1_outputs[8074];
    assign layer2_outputs[2137] = layer1_outputs[8970];
    assign layer2_outputs[2138] = ~(layer1_outputs[9885]);
    assign layer2_outputs[2139] = layer1_outputs[2737];
    assign layer2_outputs[2140] = (layer1_outputs[6913]) & ~(layer1_outputs[8872]);
    assign layer2_outputs[2141] = ~(layer1_outputs[5164]) | (layer1_outputs[8349]);
    assign layer2_outputs[2142] = ~((layer1_outputs[10899]) & (layer1_outputs[4816]));
    assign layer2_outputs[2143] = ~((layer1_outputs[6305]) ^ (layer1_outputs[9205]));
    assign layer2_outputs[2144] = ~((layer1_outputs[5513]) & (layer1_outputs[384]));
    assign layer2_outputs[2145] = ~(layer1_outputs[10996]);
    assign layer2_outputs[2146] = ~((layer1_outputs[9776]) ^ (layer1_outputs[3734]));
    assign layer2_outputs[2147] = (layer1_outputs[6028]) ^ (layer1_outputs[10364]);
    assign layer2_outputs[2148] = (layer1_outputs[8262]) | (layer1_outputs[7768]);
    assign layer2_outputs[2149] = layer1_outputs[12635];
    assign layer2_outputs[2150] = ~(layer1_outputs[7525]);
    assign layer2_outputs[2151] = layer1_outputs[11124];
    assign layer2_outputs[2152] = ~(layer1_outputs[8035]);
    assign layer2_outputs[2153] = ~(layer1_outputs[3500]) | (layer1_outputs[4128]);
    assign layer2_outputs[2154] = ~(layer1_outputs[12579]);
    assign layer2_outputs[2155] = ~((layer1_outputs[2936]) ^ (layer1_outputs[7371]));
    assign layer2_outputs[2156] = (layer1_outputs[8154]) ^ (layer1_outputs[9962]);
    assign layer2_outputs[2157] = ~(layer1_outputs[11082]);
    assign layer2_outputs[2158] = ~(layer1_outputs[8172]);
    assign layer2_outputs[2159] = ~(layer1_outputs[10662]) | (layer1_outputs[2490]);
    assign layer2_outputs[2160] = layer1_outputs[11593];
    assign layer2_outputs[2161] = ~((layer1_outputs[5563]) ^ (layer1_outputs[1216]));
    assign layer2_outputs[2162] = ~(layer1_outputs[4986]);
    assign layer2_outputs[2163] = layer1_outputs[9360];
    assign layer2_outputs[2164] = ~(layer1_outputs[1487]);
    assign layer2_outputs[2165] = (layer1_outputs[11531]) ^ (layer1_outputs[5137]);
    assign layer2_outputs[2166] = ~(layer1_outputs[1206]);
    assign layer2_outputs[2167] = ~((layer1_outputs[2384]) | (layer1_outputs[3883]));
    assign layer2_outputs[2168] = layer1_outputs[11652];
    assign layer2_outputs[2169] = layer1_outputs[7972];
    assign layer2_outputs[2170] = (layer1_outputs[10780]) & ~(layer1_outputs[151]);
    assign layer2_outputs[2171] = (layer1_outputs[445]) & (layer1_outputs[4833]);
    assign layer2_outputs[2172] = layer1_outputs[1865];
    assign layer2_outputs[2173] = layer1_outputs[12795];
    assign layer2_outputs[2174] = ~(layer1_outputs[5325]) | (layer1_outputs[4427]);
    assign layer2_outputs[2175] = ~(layer1_outputs[7019]) | (layer1_outputs[9958]);
    assign layer2_outputs[2176] = ~((layer1_outputs[12381]) | (layer1_outputs[4508]));
    assign layer2_outputs[2177] = (layer1_outputs[579]) & ~(layer1_outputs[672]);
    assign layer2_outputs[2178] = ~(layer1_outputs[1372]);
    assign layer2_outputs[2179] = ~((layer1_outputs[9048]) & (layer1_outputs[2668]));
    assign layer2_outputs[2180] = (layer1_outputs[2301]) & ~(layer1_outputs[5828]);
    assign layer2_outputs[2181] = ~((layer1_outputs[7576]) ^ (layer1_outputs[8687]));
    assign layer2_outputs[2182] = ~(layer1_outputs[12544]);
    assign layer2_outputs[2183] = ~(layer1_outputs[6048]) | (layer1_outputs[10196]);
    assign layer2_outputs[2184] = ~(layer1_outputs[11396]);
    assign layer2_outputs[2185] = (layer1_outputs[2110]) ^ (layer1_outputs[10528]);
    assign layer2_outputs[2186] = ~(layer1_outputs[2195]) | (layer1_outputs[8166]);
    assign layer2_outputs[2187] = (layer1_outputs[8587]) ^ (layer1_outputs[9372]);
    assign layer2_outputs[2188] = layer1_outputs[5864];
    assign layer2_outputs[2189] = ~((layer1_outputs[8730]) & (layer1_outputs[624]));
    assign layer2_outputs[2190] = ~(layer1_outputs[9680]);
    assign layer2_outputs[2191] = (layer1_outputs[2265]) | (layer1_outputs[1132]);
    assign layer2_outputs[2192] = ~(layer1_outputs[12375]);
    assign layer2_outputs[2193] = (layer1_outputs[1331]) ^ (layer1_outputs[10811]);
    assign layer2_outputs[2194] = (layer1_outputs[12077]) & ~(layer1_outputs[7818]);
    assign layer2_outputs[2195] = layer1_outputs[9819];
    assign layer2_outputs[2196] = layer1_outputs[12084];
    assign layer2_outputs[2197] = (layer1_outputs[4189]) & ~(layer1_outputs[12589]);
    assign layer2_outputs[2198] = ~(layer1_outputs[2032]);
    assign layer2_outputs[2199] = (layer1_outputs[5326]) ^ (layer1_outputs[10807]);
    assign layer2_outputs[2200] = ~(layer1_outputs[7997]);
    assign layer2_outputs[2201] = (layer1_outputs[7780]) ^ (layer1_outputs[635]);
    assign layer2_outputs[2202] = ~((layer1_outputs[6104]) ^ (layer1_outputs[9420]));
    assign layer2_outputs[2203] = ~(layer1_outputs[4657]);
    assign layer2_outputs[2204] = ~(layer1_outputs[1890]);
    assign layer2_outputs[2205] = (layer1_outputs[1753]) & ~(layer1_outputs[6303]);
    assign layer2_outputs[2206] = (layer1_outputs[6490]) ^ (layer1_outputs[7436]);
    assign layer2_outputs[2207] = layer1_outputs[4936];
    assign layer2_outputs[2208] = (layer1_outputs[7619]) & (layer1_outputs[1718]);
    assign layer2_outputs[2209] = ~(layer1_outputs[6599]);
    assign layer2_outputs[2210] = layer1_outputs[7475];
    assign layer2_outputs[2211] = ~(layer1_outputs[4382]) | (layer1_outputs[8011]);
    assign layer2_outputs[2212] = ~(layer1_outputs[6341]);
    assign layer2_outputs[2213] = ~(layer1_outputs[2933]);
    assign layer2_outputs[2214] = ~(layer1_outputs[6164]);
    assign layer2_outputs[2215] = (layer1_outputs[10402]) ^ (layer1_outputs[4619]);
    assign layer2_outputs[2216] = (layer1_outputs[7077]) ^ (layer1_outputs[3521]);
    assign layer2_outputs[2217] = layer1_outputs[10858];
    assign layer2_outputs[2218] = ~((layer1_outputs[5739]) | (layer1_outputs[8877]));
    assign layer2_outputs[2219] = ~(layer1_outputs[5087]);
    assign layer2_outputs[2220] = layer1_outputs[6441];
    assign layer2_outputs[2221] = layer1_outputs[7420];
    assign layer2_outputs[2222] = layer1_outputs[8779];
    assign layer2_outputs[2223] = layer1_outputs[452];
    assign layer2_outputs[2224] = layer1_outputs[12135];
    assign layer2_outputs[2225] = ~(layer1_outputs[10479]);
    assign layer2_outputs[2226] = (layer1_outputs[5589]) ^ (layer1_outputs[3304]);
    assign layer2_outputs[2227] = layer1_outputs[2851];
    assign layer2_outputs[2228] = (layer1_outputs[8292]) ^ (layer1_outputs[11118]);
    assign layer2_outputs[2229] = ~(layer1_outputs[2205]);
    assign layer2_outputs[2230] = layer1_outputs[3635];
    assign layer2_outputs[2231] = ~((layer1_outputs[8350]) | (layer1_outputs[5861]));
    assign layer2_outputs[2232] = ~(layer1_outputs[1181]);
    assign layer2_outputs[2233] = layer1_outputs[10397];
    assign layer2_outputs[2234] = layer1_outputs[5324];
    assign layer2_outputs[2235] = (layer1_outputs[52]) & ~(layer1_outputs[1648]);
    assign layer2_outputs[2236] = layer1_outputs[1264];
    assign layer2_outputs[2237] = ~(layer1_outputs[7177]);
    assign layer2_outputs[2238] = ~(layer1_outputs[7590]);
    assign layer2_outputs[2239] = ~(layer1_outputs[7392]) | (layer1_outputs[1220]);
    assign layer2_outputs[2240] = (layer1_outputs[5373]) & (layer1_outputs[6173]);
    assign layer2_outputs[2241] = (layer1_outputs[11693]) & ~(layer1_outputs[11807]);
    assign layer2_outputs[2242] = ~(layer1_outputs[9967]);
    assign layer2_outputs[2243] = 1'b0;
    assign layer2_outputs[2244] = (layer1_outputs[4103]) | (layer1_outputs[9748]);
    assign layer2_outputs[2245] = ~(layer1_outputs[8257]);
    assign layer2_outputs[2246] = ~(layer1_outputs[960]);
    assign layer2_outputs[2247] = ~((layer1_outputs[9352]) | (layer1_outputs[10897]));
    assign layer2_outputs[2248] = layer1_outputs[3926];
    assign layer2_outputs[2249] = layer1_outputs[11170];
    assign layer2_outputs[2250] = layer1_outputs[11550];
    assign layer2_outputs[2251] = ~((layer1_outputs[8581]) & (layer1_outputs[8157]));
    assign layer2_outputs[2252] = layer1_outputs[12356];
    assign layer2_outputs[2253] = layer1_outputs[10546];
    assign layer2_outputs[2254] = layer1_outputs[1239];
    assign layer2_outputs[2255] = ~(layer1_outputs[6610]);
    assign layer2_outputs[2256] = (layer1_outputs[4411]) & ~(layer1_outputs[7630]);
    assign layer2_outputs[2257] = 1'b1;
    assign layer2_outputs[2258] = layer1_outputs[5925];
    assign layer2_outputs[2259] = (layer1_outputs[5936]) & (layer1_outputs[5878]);
    assign layer2_outputs[2260] = (layer1_outputs[3541]) & ~(layer1_outputs[11390]);
    assign layer2_outputs[2261] = ~(layer1_outputs[6441]);
    assign layer2_outputs[2262] = layer1_outputs[4451];
    assign layer2_outputs[2263] = layer1_outputs[4586];
    assign layer2_outputs[2264] = ~((layer1_outputs[519]) ^ (layer1_outputs[12097]));
    assign layer2_outputs[2265] = (layer1_outputs[6713]) | (layer1_outputs[2141]);
    assign layer2_outputs[2266] = ~(layer1_outputs[9896]);
    assign layer2_outputs[2267] = ~((layer1_outputs[6684]) ^ (layer1_outputs[9775]));
    assign layer2_outputs[2268] = ~(layer1_outputs[5812]) | (layer1_outputs[4101]);
    assign layer2_outputs[2269] = layer1_outputs[7013];
    assign layer2_outputs[2270] = (layer1_outputs[4310]) & (layer1_outputs[8269]);
    assign layer2_outputs[2271] = (layer1_outputs[3828]) & ~(layer1_outputs[3416]);
    assign layer2_outputs[2272] = layer1_outputs[1153];
    assign layer2_outputs[2273] = ~(layer1_outputs[6558]);
    assign layer2_outputs[2274] = layer1_outputs[248];
    assign layer2_outputs[2275] = ~(layer1_outputs[3168]) | (layer1_outputs[6600]);
    assign layer2_outputs[2276] = ~(layer1_outputs[11017]) | (layer1_outputs[3855]);
    assign layer2_outputs[2277] = ~((layer1_outputs[3698]) | (layer1_outputs[9188]));
    assign layer2_outputs[2278] = ~(layer1_outputs[5731]) | (layer1_outputs[3764]);
    assign layer2_outputs[2279] = layer1_outputs[9893];
    assign layer2_outputs[2280] = ~(layer1_outputs[10551]);
    assign layer2_outputs[2281] = layer1_outputs[4238];
    assign layer2_outputs[2282] = layer1_outputs[11699];
    assign layer2_outputs[2283] = layer1_outputs[9189];
    assign layer2_outputs[2284] = ~((layer1_outputs[8755]) ^ (layer1_outputs[4493]));
    assign layer2_outputs[2285] = (layer1_outputs[6670]) ^ (layer1_outputs[11777]);
    assign layer2_outputs[2286] = layer1_outputs[7557];
    assign layer2_outputs[2287] = ~(layer1_outputs[8690]);
    assign layer2_outputs[2288] = ~(layer1_outputs[9767]) | (layer1_outputs[2287]);
    assign layer2_outputs[2289] = ~((layer1_outputs[4780]) & (layer1_outputs[4254]));
    assign layer2_outputs[2290] = ~(layer1_outputs[5184]);
    assign layer2_outputs[2291] = ~(layer1_outputs[10711]);
    assign layer2_outputs[2292] = ~(layer1_outputs[5077]);
    assign layer2_outputs[2293] = ~((layer1_outputs[6671]) ^ (layer1_outputs[12253]));
    assign layer2_outputs[2294] = (layer1_outputs[11555]) & (layer1_outputs[8388]);
    assign layer2_outputs[2295] = layer1_outputs[8128];
    assign layer2_outputs[2296] = ~(layer1_outputs[6853]);
    assign layer2_outputs[2297] = (layer1_outputs[3860]) | (layer1_outputs[3709]);
    assign layer2_outputs[2298] = layer1_outputs[12297];
    assign layer2_outputs[2299] = ~((layer1_outputs[1187]) & (layer1_outputs[2687]));
    assign layer2_outputs[2300] = (layer1_outputs[9433]) | (layer1_outputs[10776]);
    assign layer2_outputs[2301] = (layer1_outputs[3215]) & (layer1_outputs[3377]);
    assign layer2_outputs[2302] = ~(layer1_outputs[10491]);
    assign layer2_outputs[2303] = (layer1_outputs[4658]) | (layer1_outputs[1212]);
    assign layer2_outputs[2304] = ~(layer1_outputs[564]);
    assign layer2_outputs[2305] = ~(layer1_outputs[3409]);
    assign layer2_outputs[2306] = ~((layer1_outputs[3453]) | (layer1_outputs[11322]));
    assign layer2_outputs[2307] = (layer1_outputs[3507]) & ~(layer1_outputs[2380]);
    assign layer2_outputs[2308] = ~((layer1_outputs[4707]) ^ (layer1_outputs[5019]));
    assign layer2_outputs[2309] = layer1_outputs[1554];
    assign layer2_outputs[2310] = ~(layer1_outputs[7994]);
    assign layer2_outputs[2311] = ~(layer1_outputs[7575]);
    assign layer2_outputs[2312] = ~(layer1_outputs[184]) | (layer1_outputs[8406]);
    assign layer2_outputs[2313] = ~((layer1_outputs[226]) & (layer1_outputs[2327]));
    assign layer2_outputs[2314] = layer1_outputs[912];
    assign layer2_outputs[2315] = ~(layer1_outputs[1427]);
    assign layer2_outputs[2316] = layer1_outputs[10696];
    assign layer2_outputs[2317] = (layer1_outputs[399]) | (layer1_outputs[9037]);
    assign layer2_outputs[2318] = ~((layer1_outputs[10170]) ^ (layer1_outputs[12789]));
    assign layer2_outputs[2319] = ~((layer1_outputs[9138]) & (layer1_outputs[398]));
    assign layer2_outputs[2320] = layer1_outputs[11966];
    assign layer2_outputs[2321] = layer1_outputs[5456];
    assign layer2_outputs[2322] = 1'b1;
    assign layer2_outputs[2323] = (layer1_outputs[1596]) & ~(layer1_outputs[10509]);
    assign layer2_outputs[2324] = (layer1_outputs[3766]) & (layer1_outputs[11061]);
    assign layer2_outputs[2325] = layer1_outputs[580];
    assign layer2_outputs[2326] = (layer1_outputs[1502]) & (layer1_outputs[6565]);
    assign layer2_outputs[2327] = layer1_outputs[10884];
    assign layer2_outputs[2328] = ~(layer1_outputs[4761]);
    assign layer2_outputs[2329] = (layer1_outputs[3582]) & ~(layer1_outputs[12149]);
    assign layer2_outputs[2330] = ~(layer1_outputs[3534]) | (layer1_outputs[9551]);
    assign layer2_outputs[2331] = ~(layer1_outputs[3532]);
    assign layer2_outputs[2332] = layer1_outputs[1659];
    assign layer2_outputs[2333] = ~(layer1_outputs[422]);
    assign layer2_outputs[2334] = layer1_outputs[10477];
    assign layer2_outputs[2335] = (layer1_outputs[12735]) & ~(layer1_outputs[9213]);
    assign layer2_outputs[2336] = ~(layer1_outputs[2098]);
    assign layer2_outputs[2337] = (layer1_outputs[6055]) | (layer1_outputs[508]);
    assign layer2_outputs[2338] = ~(layer1_outputs[10077]);
    assign layer2_outputs[2339] = ~(layer1_outputs[11984]) | (layer1_outputs[8844]);
    assign layer2_outputs[2340] = (layer1_outputs[8344]) & (layer1_outputs[4375]);
    assign layer2_outputs[2341] = (layer1_outputs[7154]) & (layer1_outputs[5622]);
    assign layer2_outputs[2342] = ~(layer1_outputs[8960]) | (layer1_outputs[4689]);
    assign layer2_outputs[2343] = (layer1_outputs[6296]) ^ (layer1_outputs[6445]);
    assign layer2_outputs[2344] = ~(layer1_outputs[1836]);
    assign layer2_outputs[2345] = ~(layer1_outputs[11774]);
    assign layer2_outputs[2346] = ~((layer1_outputs[12414]) | (layer1_outputs[12379]));
    assign layer2_outputs[2347] = ~(layer1_outputs[10033]);
    assign layer2_outputs[2348] = ~((layer1_outputs[5795]) & (layer1_outputs[5156]));
    assign layer2_outputs[2349] = layer1_outputs[1561];
    assign layer2_outputs[2350] = ~((layer1_outputs[9249]) & (layer1_outputs[675]));
    assign layer2_outputs[2351] = layer1_outputs[5153];
    assign layer2_outputs[2352] = layer1_outputs[4757];
    assign layer2_outputs[2353] = (layer1_outputs[5450]) & (layer1_outputs[2762]);
    assign layer2_outputs[2354] = (layer1_outputs[824]) ^ (layer1_outputs[6582]);
    assign layer2_outputs[2355] = layer1_outputs[9573];
    assign layer2_outputs[2356] = layer1_outputs[9039];
    assign layer2_outputs[2357] = ~(layer1_outputs[2739]) | (layer1_outputs[1126]);
    assign layer2_outputs[2358] = ~(layer1_outputs[3879]) | (layer1_outputs[5362]);
    assign layer2_outputs[2359] = layer1_outputs[7550];
    assign layer2_outputs[2360] = (layer1_outputs[8018]) | (layer1_outputs[9190]);
    assign layer2_outputs[2361] = ~(layer1_outputs[1170]);
    assign layer2_outputs[2362] = ~((layer1_outputs[1129]) & (layer1_outputs[4726]));
    assign layer2_outputs[2363] = ~((layer1_outputs[5870]) | (layer1_outputs[5762]));
    assign layer2_outputs[2364] = ~((layer1_outputs[9476]) & (layer1_outputs[10944]));
    assign layer2_outputs[2365] = layer1_outputs[1762];
    assign layer2_outputs[2366] = layer1_outputs[7518];
    assign layer2_outputs[2367] = layer1_outputs[11098];
    assign layer2_outputs[2368] = (layer1_outputs[10684]) ^ (layer1_outputs[11548]);
    assign layer2_outputs[2369] = 1'b1;
    assign layer2_outputs[2370] = ~(layer1_outputs[839]);
    assign layer2_outputs[2371] = (layer1_outputs[12503]) | (layer1_outputs[9346]);
    assign layer2_outputs[2372] = ~((layer1_outputs[389]) ^ (layer1_outputs[9356]));
    assign layer2_outputs[2373] = ~(layer1_outputs[8956]) | (layer1_outputs[11414]);
    assign layer2_outputs[2374] = (layer1_outputs[5376]) ^ (layer1_outputs[8543]);
    assign layer2_outputs[2375] = layer1_outputs[1869];
    assign layer2_outputs[2376] = layer1_outputs[7089];
    assign layer2_outputs[2377] = ~((layer1_outputs[12159]) & (layer1_outputs[4298]));
    assign layer2_outputs[2378] = (layer1_outputs[12641]) & ~(layer1_outputs[4113]);
    assign layer2_outputs[2379] = layer1_outputs[1078];
    assign layer2_outputs[2380] = layer1_outputs[12692];
    assign layer2_outputs[2381] = ~((layer1_outputs[174]) | (layer1_outputs[5178]));
    assign layer2_outputs[2382] = (layer1_outputs[268]) ^ (layer1_outputs[7595]);
    assign layer2_outputs[2383] = layer1_outputs[9874];
    assign layer2_outputs[2384] = layer1_outputs[12320];
    assign layer2_outputs[2385] = ~(layer1_outputs[11753]);
    assign layer2_outputs[2386] = (layer1_outputs[10087]) ^ (layer1_outputs[4558]);
    assign layer2_outputs[2387] = (layer1_outputs[3770]) & (layer1_outputs[11962]);
    assign layer2_outputs[2388] = (layer1_outputs[12029]) | (layer1_outputs[6730]);
    assign layer2_outputs[2389] = ~((layer1_outputs[3806]) ^ (layer1_outputs[2390]));
    assign layer2_outputs[2390] = ~(layer1_outputs[1603]) | (layer1_outputs[2822]);
    assign layer2_outputs[2391] = ~((layer1_outputs[5048]) ^ (layer1_outputs[8998]));
    assign layer2_outputs[2392] = ~(layer1_outputs[10881]);
    assign layer2_outputs[2393] = (layer1_outputs[6460]) & (layer1_outputs[5789]);
    assign layer2_outputs[2394] = layer1_outputs[6379];
    assign layer2_outputs[2395] = ~(layer1_outputs[8286]) | (layer1_outputs[10764]);
    assign layer2_outputs[2396] = ~((layer1_outputs[3915]) ^ (layer1_outputs[795]));
    assign layer2_outputs[2397] = ~((layer1_outputs[11354]) & (layer1_outputs[5599]));
    assign layer2_outputs[2398] = (layer1_outputs[5280]) & (layer1_outputs[3539]);
    assign layer2_outputs[2399] = ~(layer1_outputs[3863]) | (layer1_outputs[6742]);
    assign layer2_outputs[2400] = ~((layer1_outputs[11808]) & (layer1_outputs[10927]));
    assign layer2_outputs[2401] = ~(layer1_outputs[2440]);
    assign layer2_outputs[2402] = ~((layer1_outputs[6386]) | (layer1_outputs[9993]));
    assign layer2_outputs[2403] = layer1_outputs[11866];
    assign layer2_outputs[2404] = ~(layer1_outputs[11907]);
    assign layer2_outputs[2405] = (layer1_outputs[7859]) & ~(layer1_outputs[5878]);
    assign layer2_outputs[2406] = layer1_outputs[3219];
    assign layer2_outputs[2407] = layer1_outputs[10899];
    assign layer2_outputs[2408] = ~(layer1_outputs[9689]);
    assign layer2_outputs[2409] = ~((layer1_outputs[6506]) | (layer1_outputs[3876]));
    assign layer2_outputs[2410] = layer1_outputs[12363];
    assign layer2_outputs[2411] = layer1_outputs[788];
    assign layer2_outputs[2412] = ~((layer1_outputs[1170]) & (layer1_outputs[7224]));
    assign layer2_outputs[2413] = (layer1_outputs[759]) | (layer1_outputs[6027]);
    assign layer2_outputs[2414] = ~((layer1_outputs[188]) ^ (layer1_outputs[3804]));
    assign layer2_outputs[2415] = (layer1_outputs[4184]) | (layer1_outputs[9612]);
    assign layer2_outputs[2416] = layer1_outputs[11267];
    assign layer2_outputs[2417] = ~(layer1_outputs[2267]);
    assign layer2_outputs[2418] = layer1_outputs[1935];
    assign layer2_outputs[2419] = ~(layer1_outputs[2223]);
    assign layer2_outputs[2420] = ~(layer1_outputs[2109]);
    assign layer2_outputs[2421] = layer1_outputs[3100];
    assign layer2_outputs[2422] = ~((layer1_outputs[6830]) ^ (layer1_outputs[4018]));
    assign layer2_outputs[2423] = ~((layer1_outputs[10173]) ^ (layer1_outputs[8140]));
    assign layer2_outputs[2424] = ~(layer1_outputs[596]);
    assign layer2_outputs[2425] = layer1_outputs[5504];
    assign layer2_outputs[2426] = ~(layer1_outputs[8551]);
    assign layer2_outputs[2427] = layer1_outputs[431];
    assign layer2_outputs[2428] = ~(layer1_outputs[8180]);
    assign layer2_outputs[2429] = layer1_outputs[11455];
    assign layer2_outputs[2430] = ~(layer1_outputs[11886]) | (layer1_outputs[7955]);
    assign layer2_outputs[2431] = ~(layer1_outputs[8969]);
    assign layer2_outputs[2432] = ~((layer1_outputs[12203]) ^ (layer1_outputs[1197]));
    assign layer2_outputs[2433] = ~(layer1_outputs[8484]);
    assign layer2_outputs[2434] = (layer1_outputs[4897]) | (layer1_outputs[4623]);
    assign layer2_outputs[2435] = layer1_outputs[2631];
    assign layer2_outputs[2436] = ~(layer1_outputs[10772]) | (layer1_outputs[3339]);
    assign layer2_outputs[2437] = (layer1_outputs[6636]) ^ (layer1_outputs[8794]);
    assign layer2_outputs[2438] = ~(layer1_outputs[5191]);
    assign layer2_outputs[2439] = ~(layer1_outputs[4149]);
    assign layer2_outputs[2440] = ~(layer1_outputs[1850]);
    assign layer2_outputs[2441] = (layer1_outputs[2299]) & ~(layer1_outputs[4446]);
    assign layer2_outputs[2442] = (layer1_outputs[1418]) ^ (layer1_outputs[10682]);
    assign layer2_outputs[2443] = (layer1_outputs[7117]) & (layer1_outputs[1042]);
    assign layer2_outputs[2444] = (layer1_outputs[7306]) | (layer1_outputs[5081]);
    assign layer2_outputs[2445] = layer1_outputs[3515];
    assign layer2_outputs[2446] = ~(layer1_outputs[3903]);
    assign layer2_outputs[2447] = ~(layer1_outputs[2312]) | (layer1_outputs[12108]);
    assign layer2_outputs[2448] = ~((layer1_outputs[3837]) | (layer1_outputs[3477]));
    assign layer2_outputs[2449] = (layer1_outputs[1912]) ^ (layer1_outputs[11616]);
    assign layer2_outputs[2450] = layer1_outputs[11294];
    assign layer2_outputs[2451] = (layer1_outputs[469]) & ~(layer1_outputs[12174]);
    assign layer2_outputs[2452] = layer1_outputs[3616];
    assign layer2_outputs[2453] = ~(layer1_outputs[901]);
    assign layer2_outputs[2454] = ~(layer1_outputs[2341]);
    assign layer2_outputs[2455] = ~(layer1_outputs[7951]) | (layer1_outputs[3753]);
    assign layer2_outputs[2456] = (layer1_outputs[9662]) ^ (layer1_outputs[3284]);
    assign layer2_outputs[2457] = ~(layer1_outputs[3125]);
    assign layer2_outputs[2458] = (layer1_outputs[4078]) ^ (layer1_outputs[508]);
    assign layer2_outputs[2459] = ~(layer1_outputs[9428]);
    assign layer2_outputs[2460] = layer1_outputs[6523];
    assign layer2_outputs[2461] = layer1_outputs[3153];
    assign layer2_outputs[2462] = ~(layer1_outputs[498]);
    assign layer2_outputs[2463] = (layer1_outputs[5582]) & ~(layer1_outputs[6353]);
    assign layer2_outputs[2464] = ~((layer1_outputs[5964]) | (layer1_outputs[10949]));
    assign layer2_outputs[2465] = (layer1_outputs[2692]) & ~(layer1_outputs[9006]);
    assign layer2_outputs[2466] = layer1_outputs[6608];
    assign layer2_outputs[2467] = ~(layer1_outputs[3461]);
    assign layer2_outputs[2468] = ~(layer1_outputs[6371]);
    assign layer2_outputs[2469] = ~(layer1_outputs[4913]);
    assign layer2_outputs[2470] = ~((layer1_outputs[6122]) & (layer1_outputs[8091]));
    assign layer2_outputs[2471] = ~(layer1_outputs[9012]) | (layer1_outputs[6008]);
    assign layer2_outputs[2472] = ~((layer1_outputs[10179]) & (layer1_outputs[6467]));
    assign layer2_outputs[2473] = ~(layer1_outputs[8396]) | (layer1_outputs[3358]);
    assign layer2_outputs[2474] = layer1_outputs[1592];
    assign layer2_outputs[2475] = (layer1_outputs[12525]) & (layer1_outputs[5916]);
    assign layer2_outputs[2476] = layer1_outputs[2183];
    assign layer2_outputs[2477] = (layer1_outputs[4060]) & (layer1_outputs[5480]);
    assign layer2_outputs[2478] = ~((layer1_outputs[11960]) & (layer1_outputs[7172]));
    assign layer2_outputs[2479] = ~((layer1_outputs[4391]) ^ (layer1_outputs[10661]));
    assign layer2_outputs[2480] = (layer1_outputs[105]) & (layer1_outputs[2046]);
    assign layer2_outputs[2481] = ~(layer1_outputs[2769]);
    assign layer2_outputs[2482] = ~(layer1_outputs[6376]);
    assign layer2_outputs[2483] = layer1_outputs[5348];
    assign layer2_outputs[2484] = ~((layer1_outputs[2247]) & (layer1_outputs[123]));
    assign layer2_outputs[2485] = layer1_outputs[3751];
    assign layer2_outputs[2486] = (layer1_outputs[11591]) & (layer1_outputs[11623]);
    assign layer2_outputs[2487] = ~(layer1_outputs[2455]);
    assign layer2_outputs[2488] = ~((layer1_outputs[1520]) & (layer1_outputs[10741]));
    assign layer2_outputs[2489] = layer1_outputs[2792];
    assign layer2_outputs[2490] = ~(layer1_outputs[8266]) | (layer1_outputs[56]);
    assign layer2_outputs[2491] = (layer1_outputs[5720]) | (layer1_outputs[9320]);
    assign layer2_outputs[2492] = (layer1_outputs[11777]) | (layer1_outputs[11814]);
    assign layer2_outputs[2493] = ~(layer1_outputs[5340]);
    assign layer2_outputs[2494] = ~((layer1_outputs[8359]) & (layer1_outputs[9565]));
    assign layer2_outputs[2495] = ~(layer1_outputs[3436]);
    assign layer2_outputs[2496] = layer1_outputs[2503];
    assign layer2_outputs[2497] = ~(layer1_outputs[3701]);
    assign layer2_outputs[2498] = ~(layer1_outputs[12364]);
    assign layer2_outputs[2499] = ~(layer1_outputs[5913]);
    assign layer2_outputs[2500] = ~(layer1_outputs[4378]);
    assign layer2_outputs[2501] = ~(layer1_outputs[8765]) | (layer1_outputs[72]);
    assign layer2_outputs[2502] = (layer1_outputs[12693]) | (layer1_outputs[8925]);
    assign layer2_outputs[2503] = (layer1_outputs[6679]) & ~(layer1_outputs[1344]);
    assign layer2_outputs[2504] = (layer1_outputs[10259]) ^ (layer1_outputs[3494]);
    assign layer2_outputs[2505] = (layer1_outputs[3677]) & (layer1_outputs[5411]);
    assign layer2_outputs[2506] = ~(layer1_outputs[12130]) | (layer1_outputs[10504]);
    assign layer2_outputs[2507] = ~(layer1_outputs[191]);
    assign layer2_outputs[2508] = (layer1_outputs[12070]) & (layer1_outputs[7146]);
    assign layer2_outputs[2509] = layer1_outputs[2171];
    assign layer2_outputs[2510] = layer1_outputs[4902];
    assign layer2_outputs[2511] = layer1_outputs[5467];
    assign layer2_outputs[2512] = (layer1_outputs[3672]) ^ (layer1_outputs[6431]);
    assign layer2_outputs[2513] = ~(layer1_outputs[2536]) | (layer1_outputs[5892]);
    assign layer2_outputs[2514] = ~(layer1_outputs[2828]);
    assign layer2_outputs[2515] = layer1_outputs[945];
    assign layer2_outputs[2516] = ~(layer1_outputs[11649]);
    assign layer2_outputs[2517] = layer1_outputs[6270];
    assign layer2_outputs[2518] = (layer1_outputs[3853]) & ~(layer1_outputs[9381]);
    assign layer2_outputs[2519] = ~(layer1_outputs[8826]) | (layer1_outputs[3054]);
    assign layer2_outputs[2520] = ~((layer1_outputs[1569]) ^ (layer1_outputs[9913]));
    assign layer2_outputs[2521] = ~(layer1_outputs[5315]) | (layer1_outputs[12709]);
    assign layer2_outputs[2522] = ~(layer1_outputs[7381]) | (layer1_outputs[9583]);
    assign layer2_outputs[2523] = layer1_outputs[10207];
    assign layer2_outputs[2524] = layer1_outputs[10181];
    assign layer2_outputs[2525] = ~((layer1_outputs[3540]) ^ (layer1_outputs[7191]));
    assign layer2_outputs[2526] = ~(layer1_outputs[5484]);
    assign layer2_outputs[2527] = layer1_outputs[7];
    assign layer2_outputs[2528] = ~((layer1_outputs[8669]) & (layer1_outputs[1063]));
    assign layer2_outputs[2529] = layer1_outputs[9946];
    assign layer2_outputs[2530] = ~(layer1_outputs[8948]);
    assign layer2_outputs[2531] = ~((layer1_outputs[6221]) & (layer1_outputs[6327]));
    assign layer2_outputs[2532] = (layer1_outputs[3058]) & ~(layer1_outputs[2037]);
    assign layer2_outputs[2533] = ~(layer1_outputs[910]);
    assign layer2_outputs[2534] = (layer1_outputs[10284]) & ~(layer1_outputs[4950]);
    assign layer2_outputs[2535] = layer1_outputs[12409];
    assign layer2_outputs[2536] = ~(layer1_outputs[8255]) | (layer1_outputs[11487]);
    assign layer2_outputs[2537] = (layer1_outputs[9307]) & (layer1_outputs[8539]);
    assign layer2_outputs[2538] = (layer1_outputs[11959]) | (layer1_outputs[8099]);
    assign layer2_outputs[2539] = layer1_outputs[6246];
    assign layer2_outputs[2540] = ~(layer1_outputs[7345]);
    assign layer2_outputs[2541] = layer1_outputs[7371];
    assign layer2_outputs[2542] = (layer1_outputs[5763]) & (layer1_outputs[10615]);
    assign layer2_outputs[2543] = layer1_outputs[7228];
    assign layer2_outputs[2544] = (layer1_outputs[1433]) | (layer1_outputs[10622]);
    assign layer2_outputs[2545] = ~((layer1_outputs[2229]) ^ (layer1_outputs[8096]));
    assign layer2_outputs[2546] = ~(layer1_outputs[12176]) | (layer1_outputs[10549]);
    assign layer2_outputs[2547] = (layer1_outputs[824]) ^ (layer1_outputs[5702]);
    assign layer2_outputs[2548] = layer1_outputs[2912];
    assign layer2_outputs[2549] = ~((layer1_outputs[294]) ^ (layer1_outputs[3425]));
    assign layer2_outputs[2550] = ~(layer1_outputs[6260]) | (layer1_outputs[3325]);
    assign layer2_outputs[2551] = (layer1_outputs[9790]) & (layer1_outputs[4813]);
    assign layer2_outputs[2552] = ~(layer1_outputs[5322]);
    assign layer2_outputs[2553] = (layer1_outputs[11222]) ^ (layer1_outputs[8796]);
    assign layer2_outputs[2554] = ~(layer1_outputs[5893]);
    assign layer2_outputs[2555] = ~(layer1_outputs[12144]);
    assign layer2_outputs[2556] = (layer1_outputs[7650]) & ~(layer1_outputs[195]);
    assign layer2_outputs[2557] = ~((layer1_outputs[1114]) ^ (layer1_outputs[11728]));
    assign layer2_outputs[2558] = ~(layer1_outputs[10740]);
    assign layer2_outputs[2559] = 1'b1;
    assign layer2_outputs[2560] = (layer1_outputs[6555]) ^ (layer1_outputs[82]);
    assign layer2_outputs[2561] = (layer1_outputs[2990]) & ~(layer1_outputs[11648]);
    assign layer2_outputs[2562] = (layer1_outputs[4597]) | (layer1_outputs[12251]);
    assign layer2_outputs[2563] = ~(layer1_outputs[8460]);
    assign layer2_outputs[2564] = layer1_outputs[12392];
    assign layer2_outputs[2565] = layer1_outputs[12516];
    assign layer2_outputs[2566] = (layer1_outputs[10647]) & ~(layer1_outputs[7967]);
    assign layer2_outputs[2567] = (layer1_outputs[945]) | (layer1_outputs[8210]);
    assign layer2_outputs[2568] = (layer1_outputs[4636]) & ~(layer1_outputs[9631]);
    assign layer2_outputs[2569] = ~((layer1_outputs[7787]) | (layer1_outputs[8647]));
    assign layer2_outputs[2570] = layer1_outputs[9490];
    assign layer2_outputs[2571] = ~(layer1_outputs[7409]);
    assign layer2_outputs[2572] = layer1_outputs[9613];
    assign layer2_outputs[2573] = ~(layer1_outputs[7682]);
    assign layer2_outputs[2574] = layer1_outputs[8543];
    assign layer2_outputs[2575] = ~(layer1_outputs[9919]);
    assign layer2_outputs[2576] = ~((layer1_outputs[6356]) | (layer1_outputs[5106]));
    assign layer2_outputs[2577] = layer1_outputs[10990];
    assign layer2_outputs[2578] = (layer1_outputs[3604]) & ~(layer1_outputs[4701]);
    assign layer2_outputs[2579] = ~((layer1_outputs[11132]) & (layer1_outputs[6936]));
    assign layer2_outputs[2580] = layer1_outputs[9804];
    assign layer2_outputs[2581] = (layer1_outputs[2257]) & ~(layer1_outputs[11368]);
    assign layer2_outputs[2582] = layer1_outputs[9261];
    assign layer2_outputs[2583] = ~((layer1_outputs[1152]) & (layer1_outputs[3176]));
    assign layer2_outputs[2584] = (layer1_outputs[1116]) & ~(layer1_outputs[656]);
    assign layer2_outputs[2585] = ~(layer1_outputs[6642]) | (layer1_outputs[11961]);
    assign layer2_outputs[2586] = layer1_outputs[1994];
    assign layer2_outputs[2587] = layer1_outputs[4328];
    assign layer2_outputs[2588] = (layer1_outputs[10093]) & ~(layer1_outputs[4204]);
    assign layer2_outputs[2589] = ~((layer1_outputs[12172]) & (layer1_outputs[7086]));
    assign layer2_outputs[2590] = ~((layer1_outputs[8572]) & (layer1_outputs[9961]));
    assign layer2_outputs[2591] = ~((layer1_outputs[2587]) | (layer1_outputs[9023]));
    assign layer2_outputs[2592] = layer1_outputs[11745];
    assign layer2_outputs[2593] = (layer1_outputs[5837]) & (layer1_outputs[10214]);
    assign layer2_outputs[2594] = layer1_outputs[4792];
    assign layer2_outputs[2595] = (layer1_outputs[11159]) ^ (layer1_outputs[9499]);
    assign layer2_outputs[2596] = ~(layer1_outputs[5391]);
    assign layer2_outputs[2597] = layer1_outputs[4556];
    assign layer2_outputs[2598] = (layer1_outputs[9548]) & ~(layer1_outputs[368]);
    assign layer2_outputs[2599] = (layer1_outputs[10096]) ^ (layer1_outputs[3859]);
    assign layer2_outputs[2600] = ~(layer1_outputs[12561]) | (layer1_outputs[10142]);
    assign layer2_outputs[2601] = layer1_outputs[8275];
    assign layer2_outputs[2602] = ~(layer1_outputs[1382]);
    assign layer2_outputs[2603] = ~(layer1_outputs[117]) | (layer1_outputs[1233]);
    assign layer2_outputs[2604] = ~(layer1_outputs[5137]);
    assign layer2_outputs[2605] = ~((layer1_outputs[1300]) & (layer1_outputs[11343]));
    assign layer2_outputs[2606] = ~(layer1_outputs[11678]);
    assign layer2_outputs[2607] = layer1_outputs[10584];
    assign layer2_outputs[2608] = layer1_outputs[7243];
    assign layer2_outputs[2609] = (layer1_outputs[9938]) ^ (layer1_outputs[2754]);
    assign layer2_outputs[2610] = ~(layer1_outputs[10403]) | (layer1_outputs[9680]);
    assign layer2_outputs[2611] = ~(layer1_outputs[2281]) | (layer1_outputs[3303]);
    assign layer2_outputs[2612] = layer1_outputs[12077];
    assign layer2_outputs[2613] = ~(layer1_outputs[8082]);
    assign layer2_outputs[2614] = ~(layer1_outputs[9109]);
    assign layer2_outputs[2615] = ~(layer1_outputs[12404]) | (layer1_outputs[9062]);
    assign layer2_outputs[2616] = ~((layer1_outputs[748]) | (layer1_outputs[3746]));
    assign layer2_outputs[2617] = layer1_outputs[11322];
    assign layer2_outputs[2618] = layer1_outputs[4368];
    assign layer2_outputs[2619] = (layer1_outputs[7073]) ^ (layer1_outputs[4824]);
    assign layer2_outputs[2620] = (layer1_outputs[11452]) & ~(layer1_outputs[10790]);
    assign layer2_outputs[2621] = layer1_outputs[7203];
    assign layer2_outputs[2622] = (layer1_outputs[1766]) ^ (layer1_outputs[12432]);
    assign layer2_outputs[2623] = ~(layer1_outputs[12336]);
    assign layer2_outputs[2624] = ~(layer1_outputs[2723]);
    assign layer2_outputs[2625] = ~(layer1_outputs[8517]);
    assign layer2_outputs[2626] = ~(layer1_outputs[6457]);
    assign layer2_outputs[2627] = ~(layer1_outputs[1090]);
    assign layer2_outputs[2628] = ~((layer1_outputs[2216]) | (layer1_outputs[69]));
    assign layer2_outputs[2629] = ~(layer1_outputs[32]);
    assign layer2_outputs[2630] = (layer1_outputs[9045]) | (layer1_outputs[4486]);
    assign layer2_outputs[2631] = ~(layer1_outputs[6382]);
    assign layer2_outputs[2632] = layer1_outputs[1588];
    assign layer2_outputs[2633] = (layer1_outputs[6533]) & ~(layer1_outputs[11449]);
    assign layer2_outputs[2634] = layer1_outputs[214];
    assign layer2_outputs[2635] = ~(layer1_outputs[9590]) | (layer1_outputs[7460]);
    assign layer2_outputs[2636] = ~(layer1_outputs[12032]);
    assign layer2_outputs[2637] = layer1_outputs[5900];
    assign layer2_outputs[2638] = (layer1_outputs[693]) | (layer1_outputs[11168]);
    assign layer2_outputs[2639] = ~((layer1_outputs[2989]) ^ (layer1_outputs[4612]));
    assign layer2_outputs[2640] = layer1_outputs[1541];
    assign layer2_outputs[2641] = (layer1_outputs[7498]) ^ (layer1_outputs[12329]);
    assign layer2_outputs[2642] = layer1_outputs[3916];
    assign layer2_outputs[2643] = ~((layer1_outputs[5415]) ^ (layer1_outputs[10569]));
    assign layer2_outputs[2644] = (layer1_outputs[6867]) & (layer1_outputs[4020]);
    assign layer2_outputs[2645] = ~((layer1_outputs[11012]) | (layer1_outputs[7121]));
    assign layer2_outputs[2646] = (layer1_outputs[6516]) & ~(layer1_outputs[5095]);
    assign layer2_outputs[2647] = layer1_outputs[10279];
    assign layer2_outputs[2648] = ~(layer1_outputs[11784]) | (layer1_outputs[6743]);
    assign layer2_outputs[2649] = ~(layer1_outputs[2950]) | (layer1_outputs[3654]);
    assign layer2_outputs[2650] = (layer1_outputs[1261]) ^ (layer1_outputs[7359]);
    assign layer2_outputs[2651] = (layer1_outputs[2570]) & ~(layer1_outputs[11697]);
    assign layer2_outputs[2652] = ~(layer1_outputs[6099]);
    assign layer2_outputs[2653] = ~(layer1_outputs[11500]) | (layer1_outputs[5236]);
    assign layer2_outputs[2654] = ~((layer1_outputs[3712]) | (layer1_outputs[1247]));
    assign layer2_outputs[2655] = ~(layer1_outputs[8333]);
    assign layer2_outputs[2656] = ~(layer1_outputs[6191]) | (layer1_outputs[8369]);
    assign layer2_outputs[2657] = (layer1_outputs[502]) & ~(layer1_outputs[2331]);
    assign layer2_outputs[2658] = ~((layer1_outputs[4140]) ^ (layer1_outputs[7786]));
    assign layer2_outputs[2659] = ~(layer1_outputs[304]);
    assign layer2_outputs[2660] = ~(layer1_outputs[1477]);
    assign layer2_outputs[2661] = ~(layer1_outputs[1694]);
    assign layer2_outputs[2662] = ~(layer1_outputs[1924]);
    assign layer2_outputs[2663] = ~(layer1_outputs[1713]);
    assign layer2_outputs[2664] = layer1_outputs[1946];
    assign layer2_outputs[2665] = ~(layer1_outputs[8878]);
    assign layer2_outputs[2666] = layer1_outputs[397];
    assign layer2_outputs[2667] = (layer1_outputs[11755]) & ~(layer1_outputs[5535]);
    assign layer2_outputs[2668] = ~(layer1_outputs[1018]);
    assign layer2_outputs[2669] = ~(layer1_outputs[6428]);
    assign layer2_outputs[2670] = ~((layer1_outputs[9975]) ^ (layer1_outputs[12243]));
    assign layer2_outputs[2671] = (layer1_outputs[2112]) | (layer1_outputs[6135]);
    assign layer2_outputs[2672] = ~((layer1_outputs[5399]) ^ (layer1_outputs[420]));
    assign layer2_outputs[2673] = (layer1_outputs[9879]) & (layer1_outputs[9978]);
    assign layer2_outputs[2674] = layer1_outputs[8938];
    assign layer2_outputs[2675] = layer1_outputs[505];
    assign layer2_outputs[2676] = layer1_outputs[1845];
    assign layer2_outputs[2677] = layer1_outputs[8271];
    assign layer2_outputs[2678] = ~((layer1_outputs[6362]) | (layer1_outputs[602]));
    assign layer2_outputs[2679] = ~(layer1_outputs[12173]) | (layer1_outputs[5486]);
    assign layer2_outputs[2680] = (layer1_outputs[4442]) | (layer1_outputs[9672]);
    assign layer2_outputs[2681] = ~(layer1_outputs[3729]);
    assign layer2_outputs[2682] = ~(layer1_outputs[1389]);
    assign layer2_outputs[2683] = (layer1_outputs[10519]) & ~(layer1_outputs[8105]);
    assign layer2_outputs[2684] = ~(layer1_outputs[3287]);
    assign layer2_outputs[2685] = (layer1_outputs[2372]) & ~(layer1_outputs[10250]);
    assign layer2_outputs[2686] = (layer1_outputs[7651]) & (layer1_outputs[8728]);
    assign layer2_outputs[2687] = layer1_outputs[8839];
    assign layer2_outputs[2688] = (layer1_outputs[10971]) & ~(layer1_outputs[12284]);
    assign layer2_outputs[2689] = ~((layer1_outputs[4898]) ^ (layer1_outputs[3904]));
    assign layer2_outputs[2690] = ~(layer1_outputs[1439]);
    assign layer2_outputs[2691] = (layer1_outputs[12704]) ^ (layer1_outputs[9581]);
    assign layer2_outputs[2692] = (layer1_outputs[4937]) | (layer1_outputs[2389]);
    assign layer2_outputs[2693] = (layer1_outputs[8023]) & ~(layer1_outputs[2801]);
    assign layer2_outputs[2694] = ~(layer1_outputs[10691]);
    assign layer2_outputs[2695] = ~(layer1_outputs[1999]);
    assign layer2_outputs[2696] = ~((layer1_outputs[9690]) ^ (layer1_outputs[9276]));
    assign layer2_outputs[2697] = layer1_outputs[4567];
    assign layer2_outputs[2698] = ~((layer1_outputs[1735]) & (layer1_outputs[4010]));
    assign layer2_outputs[2699] = ~((layer1_outputs[10384]) | (layer1_outputs[10448]));
    assign layer2_outputs[2700] = ~(layer1_outputs[1802]);
    assign layer2_outputs[2701] = (layer1_outputs[11249]) | (layer1_outputs[3184]);
    assign layer2_outputs[2702] = layer1_outputs[2888];
    assign layer2_outputs[2703] = layer1_outputs[8334];
    assign layer2_outputs[2704] = (layer1_outputs[11994]) ^ (layer1_outputs[1254]);
    assign layer2_outputs[2705] = ~(layer1_outputs[11844]);
    assign layer2_outputs[2706] = ~((layer1_outputs[2651]) & (layer1_outputs[9060]));
    assign layer2_outputs[2707] = ~(layer1_outputs[7746]);
    assign layer2_outputs[2708] = ~(layer1_outputs[6113]);
    assign layer2_outputs[2709] = layer1_outputs[2266];
    assign layer2_outputs[2710] = ~((layer1_outputs[7296]) ^ (layer1_outputs[7913]));
    assign layer2_outputs[2711] = (layer1_outputs[7077]) & ~(layer1_outputs[11631]);
    assign layer2_outputs[2712] = ~(layer1_outputs[8067]);
    assign layer2_outputs[2713] = ~((layer1_outputs[661]) ^ (layer1_outputs[9413]));
    assign layer2_outputs[2714] = (layer1_outputs[1892]) & (layer1_outputs[12184]);
    assign layer2_outputs[2715] = layer1_outputs[3560];
    assign layer2_outputs[2716] = layer1_outputs[10769];
    assign layer2_outputs[2717] = ~((layer1_outputs[4686]) ^ (layer1_outputs[10171]));
    assign layer2_outputs[2718] = (layer1_outputs[10710]) ^ (layer1_outputs[7517]);
    assign layer2_outputs[2719] = ~(layer1_outputs[4082]);
    assign layer2_outputs[2720] = (layer1_outputs[7504]) & ~(layer1_outputs[2793]);
    assign layer2_outputs[2721] = ~(layer1_outputs[9492]);
    assign layer2_outputs[2722] = (layer1_outputs[10435]) & (layer1_outputs[10079]);
    assign layer2_outputs[2723] = layer1_outputs[11156];
    assign layer2_outputs[2724] = ~((layer1_outputs[10483]) & (layer1_outputs[10697]));
    assign layer2_outputs[2725] = (layer1_outputs[3637]) & ~(layer1_outputs[1500]);
    assign layer2_outputs[2726] = ~(layer1_outputs[7736]);
    assign layer2_outputs[2727] = ~(layer1_outputs[243]) | (layer1_outputs[6940]);
    assign layer2_outputs[2728] = ~(layer1_outputs[12040]);
    assign layer2_outputs[2729] = ~(layer1_outputs[5979]) | (layer1_outputs[8863]);
    assign layer2_outputs[2730] = (layer1_outputs[12656]) & ~(layer1_outputs[7699]);
    assign layer2_outputs[2731] = (layer1_outputs[10959]) ^ (layer1_outputs[10274]);
    assign layer2_outputs[2732] = layer1_outputs[7173];
    assign layer2_outputs[2733] = layer1_outputs[10937];
    assign layer2_outputs[2734] = ~((layer1_outputs[6057]) | (layer1_outputs[12321]));
    assign layer2_outputs[2735] = layer1_outputs[3444];
    assign layer2_outputs[2736] = layer1_outputs[7369];
    assign layer2_outputs[2737] = layer1_outputs[8393];
    assign layer2_outputs[2738] = ~(layer1_outputs[12190]);
    assign layer2_outputs[2739] = (layer1_outputs[11319]) & (layer1_outputs[7149]);
    assign layer2_outputs[2740] = ~((layer1_outputs[8115]) | (layer1_outputs[408]));
    assign layer2_outputs[2741] = layer1_outputs[2025];
    assign layer2_outputs[2742] = layer1_outputs[3520];
    assign layer2_outputs[2743] = layer1_outputs[6435];
    assign layer2_outputs[2744] = 1'b1;
    assign layer2_outputs[2745] = layer1_outputs[12512];
    assign layer2_outputs[2746] = ~(layer1_outputs[1369]);
    assign layer2_outputs[2747] = layer1_outputs[2972];
    assign layer2_outputs[2748] = ~(layer1_outputs[3293]);
    assign layer2_outputs[2749] = (layer1_outputs[6745]) & ~(layer1_outputs[5465]);
    assign layer2_outputs[2750] = layer1_outputs[6323];
    assign layer2_outputs[2751] = (layer1_outputs[8064]) ^ (layer1_outputs[1135]);
    assign layer2_outputs[2752] = layer1_outputs[7070];
    assign layer2_outputs[2753] = ~((layer1_outputs[3912]) & (layer1_outputs[4858]));
    assign layer2_outputs[2754] = layer1_outputs[9045];
    assign layer2_outputs[2755] = layer1_outputs[5547];
    assign layer2_outputs[2756] = ~((layer1_outputs[60]) & (layer1_outputs[274]));
    assign layer2_outputs[2757] = layer1_outputs[6220];
    assign layer2_outputs[2758] = ~(layer1_outputs[10914]) | (layer1_outputs[2854]);
    assign layer2_outputs[2759] = layer1_outputs[2601];
    assign layer2_outputs[2760] = (layer1_outputs[7857]) & ~(layer1_outputs[10896]);
    assign layer2_outputs[2761] = ~(layer1_outputs[1590]) | (layer1_outputs[6476]);
    assign layer2_outputs[2762] = ~(layer1_outputs[4240]) | (layer1_outputs[674]);
    assign layer2_outputs[2763] = ~(layer1_outputs[10535]);
    assign layer2_outputs[2764] = ~(layer1_outputs[11600]) | (layer1_outputs[1979]);
    assign layer2_outputs[2765] = 1'b0;
    assign layer2_outputs[2766] = layer1_outputs[10892];
    assign layer2_outputs[2767] = ~((layer1_outputs[7861]) & (layer1_outputs[5157]));
    assign layer2_outputs[2768] = layer1_outputs[3595];
    assign layer2_outputs[2769] = ~(layer1_outputs[10928]);
    assign layer2_outputs[2770] = ~(layer1_outputs[8691]) | (layer1_outputs[1529]);
    assign layer2_outputs[2771] = layer1_outputs[2825];
    assign layer2_outputs[2772] = ~((layer1_outputs[2478]) ^ (layer1_outputs[9891]));
    assign layer2_outputs[2773] = ~(layer1_outputs[289]);
    assign layer2_outputs[2774] = (layer1_outputs[1552]) & ~(layer1_outputs[66]);
    assign layer2_outputs[2775] = ~(layer1_outputs[8044]) | (layer1_outputs[9682]);
    assign layer2_outputs[2776] = layer1_outputs[8298];
    assign layer2_outputs[2777] = ~(layer1_outputs[11408]);
    assign layer2_outputs[2778] = layer1_outputs[12466];
    assign layer2_outputs[2779] = (layer1_outputs[11045]) | (layer1_outputs[3732]);
    assign layer2_outputs[2780] = (layer1_outputs[2523]) ^ (layer1_outputs[1524]);
    assign layer2_outputs[2781] = ~(layer1_outputs[2054]);
    assign layer2_outputs[2782] = layer1_outputs[9726];
    assign layer2_outputs[2783] = ~((layer1_outputs[11738]) ^ (layer1_outputs[8296]));
    assign layer2_outputs[2784] = ~((layer1_outputs[11085]) ^ (layer1_outputs[3623]));
    assign layer2_outputs[2785] = ~(layer1_outputs[353]);
    assign layer2_outputs[2786] = ~(layer1_outputs[9209]) | (layer1_outputs[707]);
    assign layer2_outputs[2787] = ~((layer1_outputs[9533]) | (layer1_outputs[9011]));
    assign layer2_outputs[2788] = (layer1_outputs[9401]) | (layer1_outputs[1972]);
    assign layer2_outputs[2789] = layer1_outputs[3895];
    assign layer2_outputs[2790] = ~((layer1_outputs[9296]) ^ (layer1_outputs[2670]));
    assign layer2_outputs[2791] = ~((layer1_outputs[1984]) ^ (layer1_outputs[5398]));
    assign layer2_outputs[2792] = (layer1_outputs[11298]) & (layer1_outputs[12620]);
    assign layer2_outputs[2793] = ~((layer1_outputs[3841]) & (layer1_outputs[9800]));
    assign layer2_outputs[2794] = ~(layer1_outputs[4841]);
    assign layer2_outputs[2795] = layer1_outputs[8613];
    assign layer2_outputs[2796] = ~(layer1_outputs[8975]);
    assign layer2_outputs[2797] = ~(layer1_outputs[105]);
    assign layer2_outputs[2798] = (layer1_outputs[4296]) | (layer1_outputs[11926]);
    assign layer2_outputs[2799] = (layer1_outputs[8439]) & ~(layer1_outputs[9009]);
    assign layer2_outputs[2800] = layer1_outputs[4512];
    assign layer2_outputs[2801] = layer1_outputs[1653];
    assign layer2_outputs[2802] = ~((layer1_outputs[5305]) & (layer1_outputs[11578]));
    assign layer2_outputs[2803] = (layer1_outputs[1995]) ^ (layer1_outputs[10664]);
    assign layer2_outputs[2804] = layer1_outputs[8813];
    assign layer2_outputs[2805] = (layer1_outputs[317]) & ~(layer1_outputs[9726]);
    assign layer2_outputs[2806] = ~(layer1_outputs[9631]) | (layer1_outputs[10904]);
    assign layer2_outputs[2807] = ~(layer1_outputs[8775]);
    assign layer2_outputs[2808] = ~(layer1_outputs[5166]);
    assign layer2_outputs[2809] = layer1_outputs[7523];
    assign layer2_outputs[2810] = layer1_outputs[9351];
    assign layer2_outputs[2811] = (layer1_outputs[3430]) & ~(layer1_outputs[8280]);
    assign layer2_outputs[2812] = ~(layer1_outputs[3609]) | (layer1_outputs[10003]);
    assign layer2_outputs[2813] = (layer1_outputs[8947]) & (layer1_outputs[9901]);
    assign layer2_outputs[2814] = ~(layer1_outputs[5068]);
    assign layer2_outputs[2815] = ~(layer1_outputs[6888]);
    assign layer2_outputs[2816] = (layer1_outputs[11357]) | (layer1_outputs[8222]);
    assign layer2_outputs[2817] = (layer1_outputs[6847]) ^ (layer1_outputs[6389]);
    assign layer2_outputs[2818] = ~((layer1_outputs[2803]) | (layer1_outputs[10184]));
    assign layer2_outputs[2819] = layer1_outputs[3613];
    assign layer2_outputs[2820] = ~((layer1_outputs[3204]) & (layer1_outputs[8874]));
    assign layer2_outputs[2821] = layer1_outputs[1662];
    assign layer2_outputs[2822] = layer1_outputs[3028];
    assign layer2_outputs[2823] = ~(layer1_outputs[1015]);
    assign layer2_outputs[2824] = ~(layer1_outputs[341]);
    assign layer2_outputs[2825] = (layer1_outputs[3967]) & ~(layer1_outputs[967]);
    assign layer2_outputs[2826] = (layer1_outputs[11145]) & ~(layer1_outputs[4426]);
    assign layer2_outputs[2827] = ~((layer1_outputs[1205]) ^ (layer1_outputs[1881]));
    assign layer2_outputs[2828] = layer1_outputs[5910];
    assign layer2_outputs[2829] = ~(layer1_outputs[10572]);
    assign layer2_outputs[2830] = ~((layer1_outputs[181]) ^ (layer1_outputs[11635]));
    assign layer2_outputs[2831] = layer1_outputs[4047];
    assign layer2_outputs[2832] = ~(layer1_outputs[1673]);
    assign layer2_outputs[2833] = ~((layer1_outputs[8899]) & (layer1_outputs[6767]));
    assign layer2_outputs[2834] = ~((layer1_outputs[8326]) ^ (layer1_outputs[10130]));
    assign layer2_outputs[2835] = layer1_outputs[4748];
    assign layer2_outputs[2836] = (layer1_outputs[8552]) & (layer1_outputs[9663]);
    assign layer2_outputs[2837] = (layer1_outputs[7605]) & ~(layer1_outputs[3138]);
    assign layer2_outputs[2838] = layer1_outputs[8149];
    assign layer2_outputs[2839] = ~((layer1_outputs[9252]) & (layer1_outputs[9308]));
    assign layer2_outputs[2840] = layer1_outputs[5539];
    assign layer2_outputs[2841] = layer1_outputs[5440];
    assign layer2_outputs[2842] = ~(layer1_outputs[11358]);
    assign layer2_outputs[2843] = layer1_outputs[3182];
    assign layer2_outputs[2844] = ~(layer1_outputs[10190]);
    assign layer2_outputs[2845] = (layer1_outputs[1489]) & ~(layer1_outputs[8430]);
    assign layer2_outputs[2846] = ~(layer1_outputs[2808]);
    assign layer2_outputs[2847] = ~(layer1_outputs[4445]);
    assign layer2_outputs[2848] = (layer1_outputs[4402]) & ~(layer1_outputs[7210]);
    assign layer2_outputs[2849] = layer1_outputs[1191];
    assign layer2_outputs[2850] = ~((layer1_outputs[6487]) ^ (layer1_outputs[12205]));
    assign layer2_outputs[2851] = layer1_outputs[12589];
    assign layer2_outputs[2852] = ~(layer1_outputs[381]) | (layer1_outputs[6688]);
    assign layer2_outputs[2853] = layer1_outputs[11079];
    assign layer2_outputs[2854] = layer1_outputs[11394];
    assign layer2_outputs[2855] = ~(layer1_outputs[1623]) | (layer1_outputs[779]);
    assign layer2_outputs[2856] = ~((layer1_outputs[10939]) | (layer1_outputs[8212]));
    assign layer2_outputs[2857] = 1'b0;
    assign layer2_outputs[2858] = ~(layer1_outputs[1010]);
    assign layer2_outputs[2859] = ~(layer1_outputs[3796]);
    assign layer2_outputs[2860] = ~((layer1_outputs[12318]) | (layer1_outputs[12289]));
    assign layer2_outputs[2861] = ~(layer1_outputs[2233]) | (layer1_outputs[1760]);
    assign layer2_outputs[2862] = layer1_outputs[12663];
    assign layer2_outputs[2863] = layer1_outputs[6066];
    assign layer2_outputs[2864] = layer1_outputs[11371];
    assign layer2_outputs[2865] = layer1_outputs[7055];
    assign layer2_outputs[2866] = ~(layer1_outputs[507]);
    assign layer2_outputs[2867] = layer1_outputs[1030];
    assign layer2_outputs[2868] = ~(layer1_outputs[9462]) | (layer1_outputs[11827]);
    assign layer2_outputs[2869] = ~(layer1_outputs[1705]) | (layer1_outputs[2283]);
    assign layer2_outputs[2870] = ~(layer1_outputs[11139]) | (layer1_outputs[2994]);
    assign layer2_outputs[2871] = ~(layer1_outputs[756]);
    assign layer2_outputs[2872] = ~(layer1_outputs[11328]) | (layer1_outputs[1681]);
    assign layer2_outputs[2873] = ~(layer1_outputs[3379]);
    assign layer2_outputs[2874] = layer1_outputs[1101];
    assign layer2_outputs[2875] = layer1_outputs[4183];
    assign layer2_outputs[2876] = layer1_outputs[5154];
    assign layer2_outputs[2877] = layer1_outputs[3544];
    assign layer2_outputs[2878] = layer1_outputs[9097];
    assign layer2_outputs[2879] = ~(layer1_outputs[5705]);
    assign layer2_outputs[2880] = ~(layer1_outputs[7676]);
    assign layer2_outputs[2881] = layer1_outputs[5855];
    assign layer2_outputs[2882] = (layer1_outputs[10623]) ^ (layer1_outputs[4239]);
    assign layer2_outputs[2883] = ~(layer1_outputs[2015]);
    assign layer2_outputs[2884] = (layer1_outputs[1203]) & ~(layer1_outputs[4812]);
    assign layer2_outputs[2885] = (layer1_outputs[9774]) | (layer1_outputs[6000]);
    assign layer2_outputs[2886] = ~(layer1_outputs[10234]);
    assign layer2_outputs[2887] = ~(layer1_outputs[12008]);
    assign layer2_outputs[2888] = layer1_outputs[6697];
    assign layer2_outputs[2889] = ~(layer1_outputs[5634]);
    assign layer2_outputs[2890] = (layer1_outputs[8724]) | (layer1_outputs[1405]);
    assign layer2_outputs[2891] = layer1_outputs[2501];
    assign layer2_outputs[2892] = (layer1_outputs[3803]) ^ (layer1_outputs[4182]);
    assign layer2_outputs[2893] = (layer1_outputs[2270]) & ~(layer1_outputs[12033]);
    assign layer2_outputs[2894] = layer1_outputs[10449];
    assign layer2_outputs[2895] = ~(layer1_outputs[6655]);
    assign layer2_outputs[2896] = layer1_outputs[3870];
    assign layer2_outputs[2897] = ~((layer1_outputs[238]) | (layer1_outputs[6685]));
    assign layer2_outputs[2898] = ~(layer1_outputs[12328]);
    assign layer2_outputs[2899] = (layer1_outputs[3423]) | (layer1_outputs[5925]);
    assign layer2_outputs[2900] = (layer1_outputs[6615]) | (layer1_outputs[7984]);
    assign layer2_outputs[2901] = 1'b1;
    assign layer2_outputs[2902] = (layer1_outputs[5769]) ^ (layer1_outputs[6920]);
    assign layer2_outputs[2903] = ~(layer1_outputs[5996]);
    assign layer2_outputs[2904] = ~((layer1_outputs[7315]) ^ (layer1_outputs[11128]));
    assign layer2_outputs[2905] = layer1_outputs[1786];
    assign layer2_outputs[2906] = layer1_outputs[12147];
    assign layer2_outputs[2907] = ~(layer1_outputs[10002]);
    assign layer2_outputs[2908] = (layer1_outputs[5214]) & ~(layer1_outputs[3965]);
    assign layer2_outputs[2909] = (layer1_outputs[3511]) & ~(layer1_outputs[9645]);
    assign layer2_outputs[2910] = (layer1_outputs[2629]) ^ (layer1_outputs[9062]);
    assign layer2_outputs[2911] = layer1_outputs[3579];
    assign layer2_outputs[2912] = (layer1_outputs[3807]) | (layer1_outputs[3165]);
    assign layer2_outputs[2913] = ~(layer1_outputs[2213]) | (layer1_outputs[12456]);
    assign layer2_outputs[2914] = (layer1_outputs[5343]) ^ (layer1_outputs[2997]);
    assign layer2_outputs[2915] = layer1_outputs[9531];
    assign layer2_outputs[2916] = ~(layer1_outputs[3890]);
    assign layer2_outputs[2917] = layer1_outputs[11205];
    assign layer2_outputs[2918] = (layer1_outputs[6453]) & (layer1_outputs[1434]);
    assign layer2_outputs[2919] = ~((layer1_outputs[5176]) ^ (layer1_outputs[3610]));
    assign layer2_outputs[2920] = ~(layer1_outputs[4162]);
    assign layer2_outputs[2921] = layer1_outputs[303];
    assign layer2_outputs[2922] = ~((layer1_outputs[6802]) | (layer1_outputs[6304]));
    assign layer2_outputs[2923] = (layer1_outputs[2147]) | (layer1_outputs[23]);
    assign layer2_outputs[2924] = ~((layer1_outputs[2714]) | (layer1_outputs[2196]));
    assign layer2_outputs[2925] = (layer1_outputs[5375]) | (layer1_outputs[7883]);
    assign layer2_outputs[2926] = layer1_outputs[9300];
    assign layer2_outputs[2927] = ~(layer1_outputs[2193]) | (layer1_outputs[5160]);
    assign layer2_outputs[2928] = ~(layer1_outputs[11105]);
    assign layer2_outputs[2929] = layer1_outputs[12156];
    assign layer2_outputs[2930] = ~((layer1_outputs[10735]) ^ (layer1_outputs[4160]));
    assign layer2_outputs[2931] = layer1_outputs[5300];
    assign layer2_outputs[2932] = layer1_outputs[11880];
    assign layer2_outputs[2933] = (layer1_outputs[2944]) | (layer1_outputs[7289]);
    assign layer2_outputs[2934] = ~(layer1_outputs[9638]);
    assign layer2_outputs[2935] = ~(layer1_outputs[9817]);
    assign layer2_outputs[2936] = ~(layer1_outputs[2863]);
    assign layer2_outputs[2937] = layer1_outputs[7036];
    assign layer2_outputs[2938] = ~((layer1_outputs[7286]) & (layer1_outputs[9640]));
    assign layer2_outputs[2939] = layer1_outputs[6582];
    assign layer2_outputs[2940] = (layer1_outputs[6079]) | (layer1_outputs[1395]);
    assign layer2_outputs[2941] = ~((layer1_outputs[10892]) ^ (layer1_outputs[716]));
    assign layer2_outputs[2942] = ~(layer1_outputs[3756]);
    assign layer2_outputs[2943] = layer1_outputs[2443];
    assign layer2_outputs[2944] = (layer1_outputs[8823]) ^ (layer1_outputs[7538]);
    assign layer2_outputs[2945] = layer1_outputs[8374];
    assign layer2_outputs[2946] = ~(layer1_outputs[9925]);
    assign layer2_outputs[2947] = layer1_outputs[7972];
    assign layer2_outputs[2948] = layer1_outputs[5497];
    assign layer2_outputs[2949] = (layer1_outputs[4910]) | (layer1_outputs[2644]);
    assign layer2_outputs[2950] = ~(layer1_outputs[10142]);
    assign layer2_outputs[2951] = ~(layer1_outputs[11219]) | (layer1_outputs[943]);
    assign layer2_outputs[2952] = ~((layer1_outputs[10083]) | (layer1_outputs[7647]));
    assign layer2_outputs[2953] = layer1_outputs[8653];
    assign layer2_outputs[2954] = ~(layer1_outputs[5591]);
    assign layer2_outputs[2955] = (layer1_outputs[6507]) ^ (layer1_outputs[5372]);
    assign layer2_outputs[2956] = ~((layer1_outputs[6985]) | (layer1_outputs[5076]));
    assign layer2_outputs[2957] = ~(layer1_outputs[4029]) | (layer1_outputs[11540]);
    assign layer2_outputs[2958] = 1'b0;
    assign layer2_outputs[2959] = ~((layer1_outputs[4348]) ^ (layer1_outputs[867]));
    assign layer2_outputs[2960] = layer1_outputs[5727];
    assign layer2_outputs[2961] = ~(layer1_outputs[7046]) | (layer1_outputs[7807]);
    assign layer2_outputs[2962] = layer1_outputs[6696];
    assign layer2_outputs[2963] = (layer1_outputs[9885]) | (layer1_outputs[11426]);
    assign layer2_outputs[2964] = (layer1_outputs[12192]) & ~(layer1_outputs[11510]);
    assign layer2_outputs[2965] = (layer1_outputs[12382]) & (layer1_outputs[5823]);
    assign layer2_outputs[2966] = layer1_outputs[11696];
    assign layer2_outputs[2967] = ~(layer1_outputs[9535]);
    assign layer2_outputs[2968] = ~(layer1_outputs[7804]) | (layer1_outputs[11187]);
    assign layer2_outputs[2969] = layer1_outputs[11640];
    assign layer2_outputs[2970] = (layer1_outputs[4320]) | (layer1_outputs[1867]);
    assign layer2_outputs[2971] = layer1_outputs[2072];
    assign layer2_outputs[2972] = ~((layer1_outputs[4424]) & (layer1_outputs[6493]));
    assign layer2_outputs[2973] = layer1_outputs[2167];
    assign layer2_outputs[2974] = layer1_outputs[8090];
    assign layer2_outputs[2975] = ~(layer1_outputs[9199]) | (layer1_outputs[4841]);
    assign layer2_outputs[2976] = ~((layer1_outputs[4560]) | (layer1_outputs[10781]));
    assign layer2_outputs[2977] = ~(layer1_outputs[5687]) | (layer1_outputs[5879]);
    assign layer2_outputs[2978] = ~(layer1_outputs[2886]);
    assign layer2_outputs[2979] = layer1_outputs[4040];
    assign layer2_outputs[2980] = ~((layer1_outputs[2422]) ^ (layer1_outputs[1818]));
    assign layer2_outputs[2981] = ~((layer1_outputs[9882]) | (layer1_outputs[3460]));
    assign layer2_outputs[2982] = layer1_outputs[1597];
    assign layer2_outputs[2983] = (layer1_outputs[2024]) & ~(layer1_outputs[8016]);
    assign layer2_outputs[2984] = (layer1_outputs[3767]) & ~(layer1_outputs[10624]);
    assign layer2_outputs[2985] = (layer1_outputs[7110]) | (layer1_outputs[662]);
    assign layer2_outputs[2986] = ~(layer1_outputs[11822]);
    assign layer2_outputs[2987] = (layer1_outputs[4581]) ^ (layer1_outputs[3331]);
    assign layer2_outputs[2988] = ~(layer1_outputs[6689]);
    assign layer2_outputs[2989] = (layer1_outputs[2334]) & ~(layer1_outputs[10113]);
    assign layer2_outputs[2990] = ~(layer1_outputs[8245]);
    assign layer2_outputs[2991] = layer1_outputs[7520];
    assign layer2_outputs[2992] = ~(layer1_outputs[10455]) | (layer1_outputs[4618]);
    assign layer2_outputs[2993] = ~(layer1_outputs[8973]) | (layer1_outputs[6211]);
    assign layer2_outputs[2994] = ~(layer1_outputs[732]);
    assign layer2_outputs[2995] = ~(layer1_outputs[4419]);
    assign layer2_outputs[2996] = ~(layer1_outputs[7136]);
    assign layer2_outputs[2997] = layer1_outputs[4778];
    assign layer2_outputs[2998] = (layer1_outputs[10593]) ^ (layer1_outputs[4554]);
    assign layer2_outputs[2999] = ~(layer1_outputs[5128]);
    assign layer2_outputs[3000] = ~((layer1_outputs[6682]) ^ (layer1_outputs[6887]));
    assign layer2_outputs[3001] = ~(layer1_outputs[6311]);
    assign layer2_outputs[3002] = ~((layer1_outputs[11230]) | (layer1_outputs[6930]));
    assign layer2_outputs[3003] = (layer1_outputs[10426]) & ~(layer1_outputs[3354]);
    assign layer2_outputs[3004] = ~((layer1_outputs[3561]) & (layer1_outputs[11939]));
    assign layer2_outputs[3005] = ~(layer1_outputs[3936]);
    assign layer2_outputs[3006] = (layer1_outputs[8864]) ^ (layer1_outputs[733]);
    assign layer2_outputs[3007] = (layer1_outputs[2456]) | (layer1_outputs[11994]);
    assign layer2_outputs[3008] = ~(layer1_outputs[11149]);
    assign layer2_outputs[3009] = ~(layer1_outputs[10178]);
    assign layer2_outputs[3010] = ~((layer1_outputs[3029]) & (layer1_outputs[11278]));
    assign layer2_outputs[3011] = ~(layer1_outputs[9870]) | (layer1_outputs[3725]);
    assign layer2_outputs[3012] = ~((layer1_outputs[4298]) & (layer1_outputs[6538]));
    assign layer2_outputs[3013] = ~(layer1_outputs[8257]);
    assign layer2_outputs[3014] = (layer1_outputs[568]) & ~(layer1_outputs[7442]);
    assign layer2_outputs[3015] = layer1_outputs[10256];
    assign layer2_outputs[3016] = ~((layer1_outputs[6201]) ^ (layer1_outputs[8039]));
    assign layer2_outputs[3017] = ~((layer1_outputs[1581]) ^ (layer1_outputs[9254]));
    assign layer2_outputs[3018] = ~(layer1_outputs[10930]);
    assign layer2_outputs[3019] = (layer1_outputs[7638]) & (layer1_outputs[8258]);
    assign layer2_outputs[3020] = (layer1_outputs[9945]) & ~(layer1_outputs[11641]);
    assign layer2_outputs[3021] = ~(layer1_outputs[1587]);
    assign layer2_outputs[3022] = layer1_outputs[6098];
    assign layer2_outputs[3023] = layer1_outputs[1109];
    assign layer2_outputs[3024] = ~(layer1_outputs[4994]);
    assign layer2_outputs[3025] = ~(layer1_outputs[3003]);
    assign layer2_outputs[3026] = (layer1_outputs[8621]) ^ (layer1_outputs[2473]);
    assign layer2_outputs[3027] = ~(layer1_outputs[11499]);
    assign layer2_outputs[3028] = ~(layer1_outputs[12070]);
    assign layer2_outputs[3029] = layer1_outputs[4479];
    assign layer2_outputs[3030] = ~(layer1_outputs[3465]);
    assign layer2_outputs[3031] = ~(layer1_outputs[1326]);
    assign layer2_outputs[3032] = (layer1_outputs[7026]) & ~(layer1_outputs[4635]);
    assign layer2_outputs[3033] = ~((layer1_outputs[5225]) & (layer1_outputs[2303]));
    assign layer2_outputs[3034] = layer1_outputs[2067];
    assign layer2_outputs[3035] = 1'b1;
    assign layer2_outputs[3036] = (layer1_outputs[8194]) ^ (layer1_outputs[7130]);
    assign layer2_outputs[3037] = layer1_outputs[3577];
    assign layer2_outputs[3038] = layer1_outputs[8225];
    assign layer2_outputs[3039] = ~(layer1_outputs[9324]);
    assign layer2_outputs[3040] = ~(layer1_outputs[9949]);
    assign layer2_outputs[3041] = (layer1_outputs[563]) & (layer1_outputs[7649]);
    assign layer2_outputs[3042] = (layer1_outputs[7939]) | (layer1_outputs[10401]);
    assign layer2_outputs[3043] = (layer1_outputs[6990]) ^ (layer1_outputs[8170]);
    assign layer2_outputs[3044] = (layer1_outputs[5317]) & ~(layer1_outputs[11743]);
    assign layer2_outputs[3045] = ~((layer1_outputs[10021]) & (layer1_outputs[1832]));
    assign layer2_outputs[3046] = ~(layer1_outputs[1970]);
    assign layer2_outputs[3047] = (layer1_outputs[1228]) | (layer1_outputs[7032]);
    assign layer2_outputs[3048] = ~((layer1_outputs[517]) & (layer1_outputs[11741]));
    assign layer2_outputs[3049] = layer1_outputs[1835];
    assign layer2_outputs[3050] = layer1_outputs[2925];
    assign layer2_outputs[3051] = (layer1_outputs[3770]) & ~(layer1_outputs[12275]);
    assign layer2_outputs[3052] = layer1_outputs[9840];
    assign layer2_outputs[3053] = (layer1_outputs[5267]) & ~(layer1_outputs[11768]);
    assign layer2_outputs[3054] = (layer1_outputs[8449]) | (layer1_outputs[2234]);
    assign layer2_outputs[3055] = ~((layer1_outputs[3113]) ^ (layer1_outputs[2455]));
    assign layer2_outputs[3056] = (layer1_outputs[1128]) | (layer1_outputs[10462]);
    assign layer2_outputs[3057] = (layer1_outputs[8311]) | (layer1_outputs[5529]);
    assign layer2_outputs[3058] = ~((layer1_outputs[4038]) & (layer1_outputs[2229]));
    assign layer2_outputs[3059] = ~(layer1_outputs[9694]);
    assign layer2_outputs[3060] = ~((layer1_outputs[10603]) | (layer1_outputs[67]));
    assign layer2_outputs[3061] = ~((layer1_outputs[526]) & (layer1_outputs[1742]));
    assign layer2_outputs[3062] = ~((layer1_outputs[10336]) ^ (layer1_outputs[7551]));
    assign layer2_outputs[3063] = ~(layer1_outputs[7107]);
    assign layer2_outputs[3064] = layer1_outputs[8162];
    assign layer2_outputs[3065] = (layer1_outputs[4219]) & ~(layer1_outputs[12140]);
    assign layer2_outputs[3066] = 1'b1;
    assign layer2_outputs[3067] = (layer1_outputs[9547]) ^ (layer1_outputs[11421]);
    assign layer2_outputs[3068] = ~((layer1_outputs[821]) | (layer1_outputs[2336]));
    assign layer2_outputs[3069] = ~((layer1_outputs[1509]) ^ (layer1_outputs[10335]));
    assign layer2_outputs[3070] = ~((layer1_outputs[7045]) ^ (layer1_outputs[5930]));
    assign layer2_outputs[3071] = layer1_outputs[4276];
    assign layer2_outputs[3072] = ~((layer1_outputs[49]) & (layer1_outputs[6405]));
    assign layer2_outputs[3073] = ~(layer1_outputs[3456]);
    assign layer2_outputs[3074] = ~(layer1_outputs[205]);
    assign layer2_outputs[3075] = ~(layer1_outputs[9265]);
    assign layer2_outputs[3076] = (layer1_outputs[7610]) | (layer1_outputs[10475]);
    assign layer2_outputs[3077] = ~(layer1_outputs[3504]);
    assign layer2_outputs[3078] = layer1_outputs[9278];
    assign layer2_outputs[3079] = (layer1_outputs[8126]) & (layer1_outputs[8344]);
    assign layer2_outputs[3080] = ~(layer1_outputs[10929]);
    assign layer2_outputs[3081] = (layer1_outputs[3066]) ^ (layer1_outputs[2127]);
    assign layer2_outputs[3082] = ~(layer1_outputs[4054]);
    assign layer2_outputs[3083] = ~((layer1_outputs[911]) | (layer1_outputs[9970]));
    assign layer2_outputs[3084] = ~(layer1_outputs[710]);
    assign layer2_outputs[3085] = ~(layer1_outputs[10215]);
    assign layer2_outputs[3086] = ~(layer1_outputs[9184]);
    assign layer2_outputs[3087] = (layer1_outputs[4294]) & (layer1_outputs[2715]);
    assign layer2_outputs[3088] = layer1_outputs[9679];
    assign layer2_outputs[3089] = layer1_outputs[6911];
    assign layer2_outputs[3090] = ~(layer1_outputs[6816]);
    assign layer2_outputs[3091] = layer1_outputs[1747];
    assign layer2_outputs[3092] = ~(layer1_outputs[10991]);
    assign layer2_outputs[3093] = ~(layer1_outputs[11951]) | (layer1_outputs[10497]);
    assign layer2_outputs[3094] = ~(layer1_outputs[3874]) | (layer1_outputs[2836]);
    assign layer2_outputs[3095] = ~((layer1_outputs[9347]) ^ (layer1_outputs[11385]));
    assign layer2_outputs[3096] = ~(layer1_outputs[6459]);
    assign layer2_outputs[3097] = layer1_outputs[11499];
    assign layer2_outputs[3098] = ~(layer1_outputs[5480]);
    assign layer2_outputs[3099] = layer1_outputs[10132];
    assign layer2_outputs[3100] = (layer1_outputs[3064]) & (layer1_outputs[6058]);
    assign layer2_outputs[3101] = ~(layer1_outputs[2590]);
    assign layer2_outputs[3102] = (layer1_outputs[3643]) ^ (layer1_outputs[6828]);
    assign layer2_outputs[3103] = ~((layer1_outputs[9118]) ^ (layer1_outputs[9545]));
    assign layer2_outputs[3104] = (layer1_outputs[11584]) ^ (layer1_outputs[7119]);
    assign layer2_outputs[3105] = ~(layer1_outputs[1184]);
    assign layer2_outputs[3106] = (layer1_outputs[6463]) | (layer1_outputs[7310]);
    assign layer2_outputs[3107] = (layer1_outputs[7908]) & (layer1_outputs[225]);
    assign layer2_outputs[3108] = ~(layer1_outputs[1732]);
    assign layer2_outputs[3109] = layer1_outputs[786];
    assign layer2_outputs[3110] = (layer1_outputs[1831]) | (layer1_outputs[12385]);
    assign layer2_outputs[3111] = ~((layer1_outputs[6439]) ^ (layer1_outputs[7414]));
    assign layer2_outputs[3112] = layer1_outputs[3554];
    assign layer2_outputs[3113] = (layer1_outputs[6394]) & ~(layer1_outputs[630]);
    assign layer2_outputs[3114] = ~(layer1_outputs[1089]);
    assign layer2_outputs[3115] = (layer1_outputs[1021]) & ~(layer1_outputs[14]);
    assign layer2_outputs[3116] = ~(layer1_outputs[2062]);
    assign layer2_outputs[3117] = layer1_outputs[9297];
    assign layer2_outputs[3118] = ~(layer1_outputs[5085]);
    assign layer2_outputs[3119] = ~((layer1_outputs[7753]) ^ (layer1_outputs[11903]));
    assign layer2_outputs[3120] = layer1_outputs[198];
    assign layer2_outputs[3121] = ~((layer1_outputs[5919]) | (layer1_outputs[4075]));
    assign layer2_outputs[3122] = layer1_outputs[5144];
    assign layer2_outputs[3123] = (layer1_outputs[11062]) & (layer1_outputs[5595]);
    assign layer2_outputs[3124] = ~((layer1_outputs[4364]) ^ (layer1_outputs[10653]));
    assign layer2_outputs[3125] = ~((layer1_outputs[10817]) ^ (layer1_outputs[11877]));
    assign layer2_outputs[3126] = (layer1_outputs[158]) ^ (layer1_outputs[9621]);
    assign layer2_outputs[3127] = layer1_outputs[4649];
    assign layer2_outputs[3128] = ~(layer1_outputs[10781]);
    assign layer2_outputs[3129] = layer1_outputs[7490];
    assign layer2_outputs[3130] = layer1_outputs[8147];
    assign layer2_outputs[3131] = ~(layer1_outputs[4203]);
    assign layer2_outputs[3132] = (layer1_outputs[1141]) & ~(layer1_outputs[3009]);
    assign layer2_outputs[3133] = ~(layer1_outputs[3997]);
    assign layer2_outputs[3134] = (layer1_outputs[11466]) | (layer1_outputs[1808]);
    assign layer2_outputs[3135] = layer1_outputs[8790];
    assign layer2_outputs[3136] = layer1_outputs[9129];
    assign layer2_outputs[3137] = ~((layer1_outputs[7700]) ^ (layer1_outputs[4694]));
    assign layer2_outputs[3138] = ~((layer1_outputs[2703]) & (layer1_outputs[9859]));
    assign layer2_outputs[3139] = layer1_outputs[12039];
    assign layer2_outputs[3140] = (layer1_outputs[12021]) & ~(layer1_outputs[10968]);
    assign layer2_outputs[3141] = layer1_outputs[7858];
    assign layer2_outputs[3142] = ~(layer1_outputs[8075]) | (layer1_outputs[4697]);
    assign layer2_outputs[3143] = (layer1_outputs[11017]) & ~(layer1_outputs[3471]);
    assign layer2_outputs[3144] = ~(layer1_outputs[3715]) | (layer1_outputs[10155]);
    assign layer2_outputs[3145] = ~(layer1_outputs[6539]);
    assign layer2_outputs[3146] = ~((layer1_outputs[10466]) ^ (layer1_outputs[4514]));
    assign layer2_outputs[3147] = (layer1_outputs[4257]) & ~(layer1_outputs[5843]);
    assign layer2_outputs[3148] = layer1_outputs[5367];
    assign layer2_outputs[3149] = layer1_outputs[2677];
    assign layer2_outputs[3150] = ~(layer1_outputs[12727]);
    assign layer2_outputs[3151] = (layer1_outputs[5820]) & ~(layer1_outputs[2401]);
    assign layer2_outputs[3152] = layer1_outputs[8107];
    assign layer2_outputs[3153] = ~((layer1_outputs[1630]) ^ (layer1_outputs[12757]));
    assign layer2_outputs[3154] = 1'b1;
    assign layer2_outputs[3155] = ~(layer1_outputs[2884]);
    assign layer2_outputs[3156] = layer1_outputs[12064];
    assign layer2_outputs[3157] = ~((layer1_outputs[2224]) ^ (layer1_outputs[4731]));
    assign layer2_outputs[3158] = ~((layer1_outputs[9536]) & (layer1_outputs[4989]));
    assign layer2_outputs[3159] = ~(layer1_outputs[6301]);
    assign layer2_outputs[3160] = layer1_outputs[1277];
    assign layer2_outputs[3161] = ~(layer1_outputs[6828]) | (layer1_outputs[889]);
    assign layer2_outputs[3162] = ~(layer1_outputs[5271]);
    assign layer2_outputs[3163] = ~(layer1_outputs[36]);
    assign layer2_outputs[3164] = (layer1_outputs[12293]) ^ (layer1_outputs[5748]);
    assign layer2_outputs[3165] = ~(layer1_outputs[10795]) | (layer1_outputs[2273]);
    assign layer2_outputs[3166] = ~((layer1_outputs[12712]) ^ (layer1_outputs[542]));
    assign layer2_outputs[3167] = (layer1_outputs[7654]) & ~(layer1_outputs[5129]);
    assign layer2_outputs[3168] = ~((layer1_outputs[8316]) | (layer1_outputs[806]));
    assign layer2_outputs[3169] = ~((layer1_outputs[12403]) ^ (layer1_outputs[1917]));
    assign layer2_outputs[3170] = (layer1_outputs[3575]) | (layer1_outputs[9089]);
    assign layer2_outputs[3171] = layer1_outputs[2657];
    assign layer2_outputs[3172] = layer1_outputs[1247];
    assign layer2_outputs[3173] = (layer1_outputs[129]) | (layer1_outputs[5835]);
    assign layer2_outputs[3174] = (layer1_outputs[4115]) | (layer1_outputs[8113]);
    assign layer2_outputs[3175] = ~(layer1_outputs[8241]);
    assign layer2_outputs[3176] = ~(layer1_outputs[5760]) | (layer1_outputs[11978]);
    assign layer2_outputs[3177] = ~(layer1_outputs[5883]);
    assign layer2_outputs[3178] = (layer1_outputs[239]) | (layer1_outputs[1488]);
    assign layer2_outputs[3179] = ~(layer1_outputs[9454]);
    assign layer2_outputs[3180] = (layer1_outputs[7727]) | (layer1_outputs[1231]);
    assign layer2_outputs[3181] = ~((layer1_outputs[7740]) & (layer1_outputs[10172]));
    assign layer2_outputs[3182] = ~((layer1_outputs[11303]) ^ (layer1_outputs[10405]));
    assign layer2_outputs[3183] = ~(layer1_outputs[476]);
    assign layer2_outputs[3184] = (layer1_outputs[4337]) & (layer1_outputs[6676]);
    assign layer2_outputs[3185] = ~(layer1_outputs[5869]);
    assign layer2_outputs[3186] = (layer1_outputs[9354]) & ~(layer1_outputs[6380]);
    assign layer2_outputs[3187] = ~(layer1_outputs[4116]);
    assign layer2_outputs[3188] = ~(layer1_outputs[6357]) | (layer1_outputs[11634]);
    assign layer2_outputs[3189] = ~((layer1_outputs[11250]) | (layer1_outputs[12246]));
    assign layer2_outputs[3190] = ~(layer1_outputs[8622]);
    assign layer2_outputs[3191] = layer1_outputs[11435];
    assign layer2_outputs[3192] = ~((layer1_outputs[4720]) | (layer1_outputs[5405]));
    assign layer2_outputs[3193] = ~(layer1_outputs[8139]);
    assign layer2_outputs[3194] = (layer1_outputs[9240]) ^ (layer1_outputs[6446]);
    assign layer2_outputs[3195] = ~(layer1_outputs[5834]);
    assign layer2_outputs[3196] = ~((layer1_outputs[2605]) ^ (layer1_outputs[4080]));
    assign layer2_outputs[3197] = (layer1_outputs[6155]) & ~(layer1_outputs[8375]);
    assign layer2_outputs[3198] = (layer1_outputs[4260]) & ~(layer1_outputs[8346]);
    assign layer2_outputs[3199] = ~((layer1_outputs[2238]) ^ (layer1_outputs[6740]));
    assign layer2_outputs[3200] = ~(layer1_outputs[2411]);
    assign layer2_outputs[3201] = ~((layer1_outputs[2910]) | (layer1_outputs[9417]));
    assign layer2_outputs[3202] = ~(layer1_outputs[3847]) | (layer1_outputs[8950]);
    assign layer2_outputs[3203] = ~(layer1_outputs[3126]);
    assign layer2_outputs[3204] = ~(layer1_outputs[2954]) | (layer1_outputs[1523]);
    assign layer2_outputs[3205] = layer1_outputs[462];
    assign layer2_outputs[3206] = ~((layer1_outputs[4076]) | (layer1_outputs[3622]));
    assign layer2_outputs[3207] = ~((layer1_outputs[5260]) & (layer1_outputs[2963]));
    assign layer2_outputs[3208] = layer1_outputs[3384];
    assign layer2_outputs[3209] = ~(layer1_outputs[9542]);
    assign layer2_outputs[3210] = ~(layer1_outputs[12474]) | (layer1_outputs[5039]);
    assign layer2_outputs[3211] = ~((layer1_outputs[11916]) & (layer1_outputs[7928]));
    assign layer2_outputs[3212] = ~(layer1_outputs[6288]);
    assign layer2_outputs[3213] = layer1_outputs[3789];
    assign layer2_outputs[3214] = ~(layer1_outputs[1536]);
    assign layer2_outputs[3215] = ~(layer1_outputs[1349]);
    assign layer2_outputs[3216] = ~(layer1_outputs[10509]);
    assign layer2_outputs[3217] = ~(layer1_outputs[12055]);
    assign layer2_outputs[3218] = (layer1_outputs[2802]) ^ (layer1_outputs[7302]);
    assign layer2_outputs[3219] = (layer1_outputs[2406]) & (layer1_outputs[10225]);
    assign layer2_outputs[3220] = 1'b1;
    assign layer2_outputs[3221] = ~(layer1_outputs[8885]);
    assign layer2_outputs[3222] = ~((layer1_outputs[8579]) & (layer1_outputs[10062]));
    assign layer2_outputs[3223] = ~(layer1_outputs[9142]);
    assign layer2_outputs[3224] = 1'b0;
    assign layer2_outputs[3225] = ~(layer1_outputs[649]);
    assign layer2_outputs[3226] = (layer1_outputs[5115]) & ~(layer1_outputs[6218]);
    assign layer2_outputs[3227] = ~(layer1_outputs[3049]) | (layer1_outputs[7855]);
    assign layer2_outputs[3228] = ~((layer1_outputs[1559]) & (layer1_outputs[2737]));
    assign layer2_outputs[3229] = layer1_outputs[9494];
    assign layer2_outputs[3230] = ~((layer1_outputs[4728]) ^ (layer1_outputs[11119]));
    assign layer2_outputs[3231] = layer1_outputs[10129];
    assign layer2_outputs[3232] = ~(layer1_outputs[2695]);
    assign layer2_outputs[3233] = layer1_outputs[12514];
    assign layer2_outputs[3234] = (layer1_outputs[5696]) & ~(layer1_outputs[494]);
    assign layer2_outputs[3235] = ~(layer1_outputs[1741]) | (layer1_outputs[2980]);
    assign layer2_outputs[3236] = ~(layer1_outputs[12749]);
    assign layer2_outputs[3237] = layer1_outputs[11404];
    assign layer2_outputs[3238] = layer1_outputs[616];
    assign layer2_outputs[3239] = ~((layer1_outputs[5821]) | (layer1_outputs[9217]));
    assign layer2_outputs[3240] = ~(layer1_outputs[7245]);
    assign layer2_outputs[3241] = ~(layer1_outputs[8819]);
    assign layer2_outputs[3242] = (layer1_outputs[804]) & ~(layer1_outputs[426]);
    assign layer2_outputs[3243] = (layer1_outputs[3376]) | (layer1_outputs[11473]);
    assign layer2_outputs[3244] = layer1_outputs[2346];
    assign layer2_outputs[3245] = ~(layer1_outputs[11670]);
    assign layer2_outputs[3246] = ~((layer1_outputs[10442]) ^ (layer1_outputs[2950]));
    assign layer2_outputs[3247] = ~((layer1_outputs[9080]) | (layer1_outputs[6529]));
    assign layer2_outputs[3248] = (layer1_outputs[8914]) ^ (layer1_outputs[3419]);
    assign layer2_outputs[3249] = layer1_outputs[4159];
    assign layer2_outputs[3250] = (layer1_outputs[4953]) ^ (layer1_outputs[10419]);
    assign layer2_outputs[3251] = ~((layer1_outputs[2064]) ^ (layer1_outputs[9565]));
    assign layer2_outputs[3252] = ~(layer1_outputs[8216]);
    assign layer2_outputs[3253] = (layer1_outputs[921]) & ~(layer1_outputs[6351]);
    assign layer2_outputs[3254] = ~(layer1_outputs[7265]) | (layer1_outputs[10658]);
    assign layer2_outputs[3255] = ~(layer1_outputs[9840]);
    assign layer2_outputs[3256] = layer1_outputs[11399];
    assign layer2_outputs[3257] = (layer1_outputs[189]) & ~(layer1_outputs[9830]);
    assign layer2_outputs[3258] = ~((layer1_outputs[8663]) | (layer1_outputs[9588]));
    assign layer2_outputs[3259] = layer1_outputs[158];
    assign layer2_outputs[3260] = ~(layer1_outputs[3876]);
    assign layer2_outputs[3261] = ~((layer1_outputs[11400]) | (layer1_outputs[6258]));
    assign layer2_outputs[3262] = ~(layer1_outputs[10277]);
    assign layer2_outputs[3263] = layer1_outputs[11662];
    assign layer2_outputs[3264] = layer1_outputs[5618];
    assign layer2_outputs[3265] = (layer1_outputs[11559]) & ~(layer1_outputs[11254]);
    assign layer2_outputs[3266] = ~(layer1_outputs[5431]);
    assign layer2_outputs[3267] = layer1_outputs[1398];
    assign layer2_outputs[3268] = ~((layer1_outputs[4063]) & (layer1_outputs[11588]));
    assign layer2_outputs[3269] = (layer1_outputs[1607]) | (layer1_outputs[10296]);
    assign layer2_outputs[3270] = ~(layer1_outputs[1939]);
    assign layer2_outputs[3271] = (layer1_outputs[6729]) & (layer1_outputs[5677]);
    assign layer2_outputs[3272] = (layer1_outputs[10502]) & ~(layer1_outputs[5054]);
    assign layer2_outputs[3273] = layer1_outputs[10245];
    assign layer2_outputs[3274] = layer1_outputs[8058];
    assign layer2_outputs[3275] = ~((layer1_outputs[2807]) | (layer1_outputs[2624]));
    assign layer2_outputs[3276] = ~(layer1_outputs[12655]);
    assign layer2_outputs[3277] = layer1_outputs[9422];
    assign layer2_outputs[3278] = ~((layer1_outputs[10511]) ^ (layer1_outputs[9495]));
    assign layer2_outputs[3279] = ~((layer1_outputs[9817]) & (layer1_outputs[3773]));
    assign layer2_outputs[3280] = (layer1_outputs[12389]) | (layer1_outputs[3540]);
    assign layer2_outputs[3281] = ~((layer1_outputs[11021]) ^ (layer1_outputs[7801]));
    assign layer2_outputs[3282] = (layer1_outputs[2023]) ^ (layer1_outputs[10331]);
    assign layer2_outputs[3283] = layer1_outputs[4521];
    assign layer2_outputs[3284] = layer1_outputs[6344];
    assign layer2_outputs[3285] = (layer1_outputs[6630]) ^ (layer1_outputs[8602]);
    assign layer2_outputs[3286] = (layer1_outputs[1367]) | (layer1_outputs[7778]);
    assign layer2_outputs[3287] = ~(layer1_outputs[4878]);
    assign layer2_outputs[3288] = layer1_outputs[873];
    assign layer2_outputs[3289] = ~((layer1_outputs[179]) ^ (layer1_outputs[4318]));
    assign layer2_outputs[3290] = (layer1_outputs[7909]) & ~(layer1_outputs[7668]);
    assign layer2_outputs[3291] = layer1_outputs[2841];
    assign layer2_outputs[3292] = ~(layer1_outputs[2316]) | (layer1_outputs[9752]);
    assign layer2_outputs[3293] = layer1_outputs[5093];
    assign layer2_outputs[3294] = ~((layer1_outputs[12785]) & (layer1_outputs[3907]));
    assign layer2_outputs[3295] = layer1_outputs[10027];
    assign layer2_outputs[3296] = ~(layer1_outputs[9721]);
    assign layer2_outputs[3297] = ~(layer1_outputs[8470]);
    assign layer2_outputs[3298] = ~(layer1_outputs[7454]) | (layer1_outputs[11440]);
    assign layer2_outputs[3299] = layer1_outputs[8827];
    assign layer2_outputs[3300] = ~((layer1_outputs[5095]) ^ (layer1_outputs[10756]));
    assign layer2_outputs[3301] = layer1_outputs[11146];
    assign layer2_outputs[3302] = ~(layer1_outputs[11791]);
    assign layer2_outputs[3303] = (layer1_outputs[8366]) | (layer1_outputs[7744]);
    assign layer2_outputs[3304] = ~(layer1_outputs[12467]);
    assign layer2_outputs[3305] = ~(layer1_outputs[12621]);
    assign layer2_outputs[3306] = (layer1_outputs[10442]) ^ (layer1_outputs[9966]);
    assign layer2_outputs[3307] = ~(layer1_outputs[12763]);
    assign layer2_outputs[3308] = layer1_outputs[9134];
    assign layer2_outputs[3309] = ~(layer1_outputs[9677]);
    assign layer2_outputs[3310] = ~(layer1_outputs[8109]);
    assign layer2_outputs[3311] = layer1_outputs[9934];
    assign layer2_outputs[3312] = (layer1_outputs[10308]) & (layer1_outputs[11137]);
    assign layer2_outputs[3313] = ~(layer1_outputs[8235]);
    assign layer2_outputs[3314] = (layer1_outputs[5197]) & ~(layer1_outputs[3361]);
    assign layer2_outputs[3315] = ~(layer1_outputs[4603]) | (layer1_outputs[12558]);
    assign layer2_outputs[3316] = ~(layer1_outputs[6406]);
    assign layer2_outputs[3317] = layer1_outputs[1900];
    assign layer2_outputs[3318] = (layer1_outputs[11626]) & ~(layer1_outputs[7161]);
    assign layer2_outputs[3319] = layer1_outputs[6999];
    assign layer2_outputs[3320] = layer1_outputs[9953];
    assign layer2_outputs[3321] = (layer1_outputs[8384]) & ~(layer1_outputs[12114]);
    assign layer2_outputs[3322] = layer1_outputs[6738];
    assign layer2_outputs[3323] = ~(layer1_outputs[2125]);
    assign layer2_outputs[3324] = (layer1_outputs[3277]) ^ (layer1_outputs[10350]);
    assign layer2_outputs[3325] = ~(layer1_outputs[10297]);
    assign layer2_outputs[3326] = layer1_outputs[4642];
    assign layer2_outputs[3327] = (layer1_outputs[5232]) ^ (layer1_outputs[2113]);
    assign layer2_outputs[3328] = ~(layer1_outputs[1054]) | (layer1_outputs[1161]);
    assign layer2_outputs[3329] = ~((layer1_outputs[9446]) | (layer1_outputs[11716]));
    assign layer2_outputs[3330] = (layer1_outputs[7332]) ^ (layer1_outputs[12655]);
    assign layer2_outputs[3331] = (layer1_outputs[2805]) & ~(layer1_outputs[10616]);
    assign layer2_outputs[3332] = (layer1_outputs[1451]) & (layer1_outputs[9501]);
    assign layer2_outputs[3333] = ~(layer1_outputs[5230]) | (layer1_outputs[7065]);
    assign layer2_outputs[3334] = ~(layer1_outputs[7507]);
    assign layer2_outputs[3335] = layer1_outputs[11067];
    assign layer2_outputs[3336] = layer1_outputs[5952];
    assign layer2_outputs[3337] = ~(layer1_outputs[6645]);
    assign layer2_outputs[3338] = ~((layer1_outputs[11981]) | (layer1_outputs[1201]));
    assign layer2_outputs[3339] = (layer1_outputs[6592]) ^ (layer1_outputs[11648]);
    assign layer2_outputs[3340] = ~((layer1_outputs[360]) & (layer1_outputs[5936]));
    assign layer2_outputs[3341] = (layer1_outputs[9319]) | (layer1_outputs[8683]);
    assign layer2_outputs[3342] = ~(layer1_outputs[6516]);
    assign layer2_outputs[3343] = ~(layer1_outputs[1000]) | (layer1_outputs[1965]);
    assign layer2_outputs[3344] = (layer1_outputs[7343]) & ~(layer1_outputs[4804]);
    assign layer2_outputs[3345] = ~(layer1_outputs[9047]);
    assign layer2_outputs[3346] = layer1_outputs[5502];
    assign layer2_outputs[3347] = (layer1_outputs[3557]) & ~(layer1_outputs[4264]);
    assign layer2_outputs[3348] = ~(layer1_outputs[5318]) | (layer1_outputs[7516]);
    assign layer2_outputs[3349] = (layer1_outputs[2756]) | (layer1_outputs[4549]);
    assign layer2_outputs[3350] = layer1_outputs[4509];
    assign layer2_outputs[3351] = layer1_outputs[2969];
    assign layer2_outputs[3352] = layer1_outputs[6147];
    assign layer2_outputs[3353] = ~((layer1_outputs[3655]) ^ (layer1_outputs[839]));
    assign layer2_outputs[3354] = layer1_outputs[3678];
    assign layer2_outputs[3355] = layer1_outputs[101];
    assign layer2_outputs[3356] = ~((layer1_outputs[7704]) ^ (layer1_outputs[11840]));
    assign layer2_outputs[3357] = ~(layer1_outputs[9028]);
    assign layer2_outputs[3358] = layer1_outputs[12628];
    assign layer2_outputs[3359] = ~((layer1_outputs[7747]) ^ (layer1_outputs[364]));
    assign layer2_outputs[3360] = layer1_outputs[6528];
    assign layer2_outputs[3361] = ~(layer1_outputs[1437]);
    assign layer2_outputs[3362] = ~(layer1_outputs[93]) | (layer1_outputs[5205]);
    assign layer2_outputs[3363] = layer1_outputs[6137];
    assign layer2_outputs[3364] = (layer1_outputs[8025]) | (layer1_outputs[6570]);
    assign layer2_outputs[3365] = (layer1_outputs[11197]) & ~(layer1_outputs[2180]);
    assign layer2_outputs[3366] = (layer1_outputs[2575]) & ~(layer1_outputs[4112]);
    assign layer2_outputs[3367] = layer1_outputs[2760];
    assign layer2_outputs[3368] = layer1_outputs[5896];
    assign layer2_outputs[3369] = layer1_outputs[7895];
    assign layer2_outputs[3370] = ~(layer1_outputs[2663]);
    assign layer2_outputs[3371] = ~(layer1_outputs[5037]);
    assign layer2_outputs[3372] = ~(layer1_outputs[4531]);
    assign layer2_outputs[3373] = layer1_outputs[7354];
    assign layer2_outputs[3374] = ~(layer1_outputs[388]);
    assign layer2_outputs[3375] = (layer1_outputs[11308]) & ~(layer1_outputs[8605]);
    assign layer2_outputs[3376] = layer1_outputs[1710];
    assign layer2_outputs[3377] = layer1_outputs[247];
    assign layer2_outputs[3378] = 1'b0;
    assign layer2_outputs[3379] = ~(layer1_outputs[5840]);
    assign layer2_outputs[3380] = ~((layer1_outputs[6918]) & (layer1_outputs[10030]));
    assign layer2_outputs[3381] = (layer1_outputs[10979]) & ~(layer1_outputs[5805]);
    assign layer2_outputs[3382] = layer1_outputs[2482];
    assign layer2_outputs[3383] = ~(layer1_outputs[4463]) | (layer1_outputs[7852]);
    assign layer2_outputs[3384] = ~(layer1_outputs[2586]);
    assign layer2_outputs[3385] = ~((layer1_outputs[1781]) ^ (layer1_outputs[9795]));
    assign layer2_outputs[3386] = (layer1_outputs[1667]) & (layer1_outputs[3705]);
    assign layer2_outputs[3387] = ~(layer1_outputs[3462]);
    assign layer2_outputs[3388] = ~(layer1_outputs[5124]);
    assign layer2_outputs[3389] = layer1_outputs[11333];
    assign layer2_outputs[3390] = (layer1_outputs[9219]) ^ (layer1_outputs[5545]);
    assign layer2_outputs[3391] = (layer1_outputs[10547]) | (layer1_outputs[4875]);
    assign layer2_outputs[3392] = layer1_outputs[9004];
    assign layer2_outputs[3393] = layer1_outputs[7570];
    assign layer2_outputs[3394] = (layer1_outputs[4990]) & (layer1_outputs[5907]);
    assign layer2_outputs[3395] = ~((layer1_outputs[6132]) & (layer1_outputs[7540]));
    assign layer2_outputs[3396] = layer1_outputs[10163];
    assign layer2_outputs[3397] = ~(layer1_outputs[1806]);
    assign layer2_outputs[3398] = layer1_outputs[7128];
    assign layer2_outputs[3399] = ~(layer1_outputs[11932]);
    assign layer2_outputs[3400] = ~((layer1_outputs[4206]) | (layer1_outputs[9698]));
    assign layer2_outputs[3401] = ~((layer1_outputs[8668]) ^ (layer1_outputs[2673]));
    assign layer2_outputs[3402] = ~(layer1_outputs[4685]) | (layer1_outputs[11226]);
    assign layer2_outputs[3403] = layer1_outputs[5429];
    assign layer2_outputs[3404] = layer1_outputs[1521];
    assign layer2_outputs[3405] = ~(layer1_outputs[6734]);
    assign layer2_outputs[3406] = ~(layer1_outputs[2350]);
    assign layer2_outputs[3407] = ~(layer1_outputs[12784]) | (layer1_outputs[10263]);
    assign layer2_outputs[3408] = ~((layer1_outputs[7904]) & (layer1_outputs[1366]));
    assign layer2_outputs[3409] = layer1_outputs[9523];
    assign layer2_outputs[3410] = ~(layer1_outputs[2433]) | (layer1_outputs[2622]);
    assign layer2_outputs[3411] = ~(layer1_outputs[1094]) | (layer1_outputs[930]);
    assign layer2_outputs[3412] = layer1_outputs[9302];
    assign layer2_outputs[3413] = layer1_outputs[10468];
    assign layer2_outputs[3414] = layer1_outputs[3012];
    assign layer2_outputs[3415] = layer1_outputs[10064];
    assign layer2_outputs[3416] = layer1_outputs[2899];
    assign layer2_outputs[3417] = (layer1_outputs[532]) | (layer1_outputs[9223]);
    assign layer2_outputs[3418] = ~(layer1_outputs[8373]) | (layer1_outputs[2525]);
    assign layer2_outputs[3419] = (layer1_outputs[10167]) & ~(layer1_outputs[5911]);
    assign layer2_outputs[3420] = layer1_outputs[1971];
    assign layer2_outputs[3421] = (layer1_outputs[8772]) ^ (layer1_outputs[1775]);
    assign layer2_outputs[3422] = ~((layer1_outputs[8130]) & (layer1_outputs[8656]));
    assign layer2_outputs[3423] = layer1_outputs[4694];
    assign layer2_outputs[3424] = (layer1_outputs[6434]) ^ (layer1_outputs[10774]);
    assign layer2_outputs[3425] = ~(layer1_outputs[11238]);
    assign layer2_outputs[3426] = (layer1_outputs[9001]) ^ (layer1_outputs[4700]);
    assign layer2_outputs[3427] = ~(layer1_outputs[8343]) | (layer1_outputs[3355]);
    assign layer2_outputs[3428] = ~(layer1_outputs[1974]);
    assign layer2_outputs[3429] = ~((layer1_outputs[9569]) ^ (layer1_outputs[11179]));
    assign layer2_outputs[3430] = (layer1_outputs[802]) & ~(layer1_outputs[7334]);
    assign layer2_outputs[3431] = (layer1_outputs[9739]) & ~(layer1_outputs[11486]);
    assign layer2_outputs[3432] = ~(layer1_outputs[4291]) | (layer1_outputs[767]);
    assign layer2_outputs[3433] = ~(layer1_outputs[11594]);
    assign layer2_outputs[3434] = ~((layer1_outputs[5891]) | (layer1_outputs[6693]));
    assign layer2_outputs[3435] = ~(layer1_outputs[9507]);
    assign layer2_outputs[3436] = layer1_outputs[11880];
    assign layer2_outputs[3437] = (layer1_outputs[7892]) ^ (layer1_outputs[11859]);
    assign layer2_outputs[3438] = layer1_outputs[5039];
    assign layer2_outputs[3439] = layer1_outputs[10177];
    assign layer2_outputs[3440] = ~((layer1_outputs[4533]) ^ (layer1_outputs[10880]));
    assign layer2_outputs[3441] = (layer1_outputs[5388]) & (layer1_outputs[5169]);
    assign layer2_outputs[3442] = layer1_outputs[10047];
    assign layer2_outputs[3443] = ~(layer1_outputs[7838]) | (layer1_outputs[9216]);
    assign layer2_outputs[3444] = ~(layer1_outputs[3271]) | (layer1_outputs[11202]);
    assign layer2_outputs[3445] = ~(layer1_outputs[8374]);
    assign layer2_outputs[3446] = (layer1_outputs[8644]) & ~(layer1_outputs[6143]);
    assign layer2_outputs[3447] = layer1_outputs[1720];
    assign layer2_outputs[3448] = ~(layer1_outputs[11332]) | (layer1_outputs[718]);
    assign layer2_outputs[3449] = ~((layer1_outputs[1951]) & (layer1_outputs[7064]));
    assign layer2_outputs[3450] = (layer1_outputs[3656]) & ~(layer1_outputs[12595]);
    assign layer2_outputs[3451] = layer1_outputs[1687];
    assign layer2_outputs[3452] = (layer1_outputs[2390]) ^ (layer1_outputs[12488]);
    assign layer2_outputs[3453] = ~(layer1_outputs[4155]);
    assign layer2_outputs[3454] = ~((layer1_outputs[5605]) | (layer1_outputs[12710]));
    assign layer2_outputs[3455] = ~((layer1_outputs[8747]) & (layer1_outputs[12204]));
    assign layer2_outputs[3456] = (layer1_outputs[3863]) | (layer1_outputs[3438]);
    assign layer2_outputs[3457] = ~(layer1_outputs[7809]);
    assign layer2_outputs[3458] = ~(layer1_outputs[9002]);
    assign layer2_outputs[3459] = ~(layer1_outputs[9520]);
    assign layer2_outputs[3460] = (layer1_outputs[6502]) ^ (layer1_outputs[1941]);
    assign layer2_outputs[3461] = ~(layer1_outputs[261]) | (layer1_outputs[8407]);
    assign layer2_outputs[3462] = layer1_outputs[589];
    assign layer2_outputs[3463] = ~(layer1_outputs[10241]);
    assign layer2_outputs[3464] = (layer1_outputs[10889]) & ~(layer1_outputs[10540]);
    assign layer2_outputs[3465] = ~(layer1_outputs[10745]);
    assign layer2_outputs[3466] = layer1_outputs[6772];
    assign layer2_outputs[3467] = layer1_outputs[1811];
    assign layer2_outputs[3468] = ~((layer1_outputs[2814]) & (layer1_outputs[8868]));
    assign layer2_outputs[3469] = ~((layer1_outputs[8420]) | (layer1_outputs[3678]));
    assign layer2_outputs[3470] = ~(layer1_outputs[2857]);
    assign layer2_outputs[3471] = layer1_outputs[2724];
    assign layer2_outputs[3472] = ~(layer1_outputs[12493]);
    assign layer2_outputs[3473] = layer1_outputs[10970];
    assign layer2_outputs[3474] = layer1_outputs[845];
    assign layer2_outputs[3475] = ~(layer1_outputs[9082]);
    assign layer2_outputs[3476] = ~(layer1_outputs[261]);
    assign layer2_outputs[3477] = ~(layer1_outputs[10587]) | (layer1_outputs[5029]);
    assign layer2_outputs[3478] = ~(layer1_outputs[4334]);
    assign layer2_outputs[3479] = ~(layer1_outputs[8750]) | (layer1_outputs[12514]);
    assign layer2_outputs[3480] = (layer1_outputs[9714]) | (layer1_outputs[3447]);
    assign layer2_outputs[3481] = (layer1_outputs[8368]) & ~(layer1_outputs[9598]);
    assign layer2_outputs[3482] = layer1_outputs[3387];
    assign layer2_outputs[3483] = (layer1_outputs[29]) ^ (layer1_outputs[9073]);
    assign layer2_outputs[3484] = ~(layer1_outputs[10855]);
    assign layer2_outputs[3485] = layer1_outputs[3026];
    assign layer2_outputs[3486] = (layer1_outputs[10286]) & ~(layer1_outputs[12177]);
    assign layer2_outputs[3487] = 1'b0;
    assign layer2_outputs[3488] = layer1_outputs[4579];
    assign layer2_outputs[3489] = ~(layer1_outputs[6060]);
    assign layer2_outputs[3490] = ~(layer1_outputs[10576]);
    assign layer2_outputs[3491] = layer1_outputs[8635];
    assign layer2_outputs[3492] = ~(layer1_outputs[8507]);
    assign layer2_outputs[3493] = ~(layer1_outputs[10404]);
    assign layer2_outputs[3494] = ~(layer1_outputs[12541]);
    assign layer2_outputs[3495] = layer1_outputs[12627];
    assign layer2_outputs[3496] = ~(layer1_outputs[3882]);
    assign layer2_outputs[3497] = ~(layer1_outputs[8451]);
    assign layer2_outputs[3498] = ~(layer1_outputs[5321]);
    assign layer2_outputs[3499] = ~(layer1_outputs[4339]);
    assign layer2_outputs[3500] = ~(layer1_outputs[10618]);
    assign layer2_outputs[3501] = ~((layer1_outputs[7299]) & (layer1_outputs[11536]));
    assign layer2_outputs[3502] = layer1_outputs[7491];
    assign layer2_outputs[3503] = (layer1_outputs[9516]) | (layer1_outputs[9124]);
    assign layer2_outputs[3504] = ~(layer1_outputs[2165]) | (layer1_outputs[11198]);
    assign layer2_outputs[3505] = layer1_outputs[979];
    assign layer2_outputs[3506] = ~((layer1_outputs[11736]) ^ (layer1_outputs[3674]));
    assign layer2_outputs[3507] = ~(layer1_outputs[9115]) | (layer1_outputs[7441]);
    assign layer2_outputs[3508] = ~(layer1_outputs[596]);
    assign layer2_outputs[3509] = ~(layer1_outputs[10342]);
    assign layer2_outputs[3510] = layer1_outputs[7157];
    assign layer2_outputs[3511] = ~(layer1_outputs[2707]);
    assign layer2_outputs[3512] = layer1_outputs[6363];
    assign layer2_outputs[3513] = ~(layer1_outputs[6063]);
    assign layer2_outputs[3514] = ~(layer1_outputs[4054]);
    assign layer2_outputs[3515] = ~(layer1_outputs[7319]);
    assign layer2_outputs[3516] = layer1_outputs[5221];
    assign layer2_outputs[3517] = layer1_outputs[2227];
    assign layer2_outputs[3518] = ~(layer1_outputs[7124]);
    assign layer2_outputs[3519] = ~(layer1_outputs[8692]) | (layer1_outputs[7627]);
    assign layer2_outputs[3520] = layer1_outputs[12781];
    assign layer2_outputs[3521] = ~((layer1_outputs[8243]) & (layer1_outputs[12634]));
    assign layer2_outputs[3522] = layer1_outputs[7332];
    assign layer2_outputs[3523] = layer1_outputs[7558];
    assign layer2_outputs[3524] = ~(layer1_outputs[2709]) | (layer1_outputs[12399]);
    assign layer2_outputs[3525] = ~(layer1_outputs[12596]);
    assign layer2_outputs[3526] = ~((layer1_outputs[1559]) ^ (layer1_outputs[12163]));
    assign layer2_outputs[3527] = ~((layer1_outputs[8524]) | (layer1_outputs[12797]));
    assign layer2_outputs[3528] = ~(layer1_outputs[9329]);
    assign layer2_outputs[3529] = layer1_outputs[6900];
    assign layer2_outputs[3530] = ~((layer1_outputs[6267]) ^ (layer1_outputs[6331]));
    assign layer2_outputs[3531] = layer1_outputs[4613];
    assign layer2_outputs[3532] = ~(layer1_outputs[10847]);
    assign layer2_outputs[3533] = ~(layer1_outputs[7322]);
    assign layer2_outputs[3534] = layer1_outputs[9477];
    assign layer2_outputs[3535] = ~(layer1_outputs[7132]) | (layer1_outputs[1683]);
    assign layer2_outputs[3536] = (layer1_outputs[898]) & ~(layer1_outputs[5926]);
    assign layer2_outputs[3537] = ~((layer1_outputs[11167]) ^ (layer1_outputs[12755]));
    assign layer2_outputs[3538] = ~(layer1_outputs[461]) | (layer1_outputs[11723]);
    assign layer2_outputs[3539] = ~(layer1_outputs[781]);
    assign layer2_outputs[3540] = ~(layer1_outputs[6656]);
    assign layer2_outputs[3541] = ~(layer1_outputs[4889]) | (layer1_outputs[7940]);
    assign layer2_outputs[3542] = (layer1_outputs[7463]) & ~(layer1_outputs[2607]);
    assign layer2_outputs[3543] = layer1_outputs[1909];
    assign layer2_outputs[3544] = 1'b0;
    assign layer2_outputs[3545] = (layer1_outputs[3919]) & (layer1_outputs[2650]);
    assign layer2_outputs[3546] = ~((layer1_outputs[4162]) | (layer1_outputs[11046]));
    assign layer2_outputs[3547] = 1'b0;
    assign layer2_outputs[3548] = ~(layer1_outputs[2136]) | (layer1_outputs[7652]);
    assign layer2_outputs[3549] = ~(layer1_outputs[377]) | (layer1_outputs[4938]);
    assign layer2_outputs[3550] = ~(layer1_outputs[3447]);
    assign layer2_outputs[3551] = layer1_outputs[244];
    assign layer2_outputs[3552] = layer1_outputs[8843];
    assign layer2_outputs[3553] = ~(layer1_outputs[6323]);
    assign layer2_outputs[3554] = ~(layer1_outputs[2619]);
    assign layer2_outputs[3555] = layer1_outputs[8528];
    assign layer2_outputs[3556] = layer1_outputs[6576];
    assign layer2_outputs[3557] = (layer1_outputs[838]) | (layer1_outputs[6164]);
    assign layer2_outputs[3558] = layer1_outputs[11469];
    assign layer2_outputs[3559] = ~(layer1_outputs[5520]);
    assign layer2_outputs[3560] = (layer1_outputs[830]) | (layer1_outputs[2515]);
    assign layer2_outputs[3561] = (layer1_outputs[7743]) | (layer1_outputs[4536]);
    assign layer2_outputs[3562] = ~(layer1_outputs[11320]);
    assign layer2_outputs[3563] = layer1_outputs[2740];
    assign layer2_outputs[3564] = layer1_outputs[11514];
    assign layer2_outputs[3565] = ~(layer1_outputs[6059]);
    assign layer2_outputs[3566] = ~(layer1_outputs[5004]);
    assign layer2_outputs[3567] = layer1_outputs[1651];
    assign layer2_outputs[3568] = layer1_outputs[5186];
    assign layer2_outputs[3569] = ~(layer1_outputs[7562]);
    assign layer2_outputs[3570] = layer1_outputs[5765];
    assign layer2_outputs[3571] = (layer1_outputs[10893]) ^ (layer1_outputs[1546]);
    assign layer2_outputs[3572] = ~(layer1_outputs[167]);
    assign layer2_outputs[3573] = ~(layer1_outputs[8465]);
    assign layer2_outputs[3574] = ~(layer1_outputs[8521]);
    assign layer2_outputs[3575] = ~(layer1_outputs[3565]);
    assign layer2_outputs[3576] = layer1_outputs[12147];
    assign layer2_outputs[3577] = (layer1_outputs[74]) & (layer1_outputs[11424]);
    assign layer2_outputs[3578] = layer1_outputs[8442];
    assign layer2_outputs[3579] = (layer1_outputs[6752]) & (layer1_outputs[1165]);
    assign layer2_outputs[3580] = (layer1_outputs[7509]) | (layer1_outputs[5617]);
    assign layer2_outputs[3581] = ~(layer1_outputs[2487]);
    assign layer2_outputs[3582] = layer1_outputs[8671];
    assign layer2_outputs[3583] = ~((layer1_outputs[1422]) & (layer1_outputs[5519]));
    assign layer2_outputs[3584] = ~((layer1_outputs[7302]) | (layer1_outputs[391]));
    assign layer2_outputs[3585] = ~((layer1_outputs[129]) ^ (layer1_outputs[1351]));
    assign layer2_outputs[3586] = ~(layer1_outputs[7736]);
    assign layer2_outputs[3587] = layer1_outputs[3136];
    assign layer2_outputs[3588] = ~((layer1_outputs[12232]) & (layer1_outputs[6244]));
    assign layer2_outputs[3589] = ~(layer1_outputs[6537]) | (layer1_outputs[2711]);
    assign layer2_outputs[3590] = (layer1_outputs[6630]) & (layer1_outputs[10963]);
    assign layer2_outputs[3591] = layer1_outputs[2595];
    assign layer2_outputs[3592] = ~(layer1_outputs[7241]);
    assign layer2_outputs[3593] = ~(layer1_outputs[6320]);
    assign layer2_outputs[3594] = layer1_outputs[10297];
    assign layer2_outputs[3595] = (layer1_outputs[9464]) & ~(layer1_outputs[410]);
    assign layer2_outputs[3596] = layer1_outputs[12507];
    assign layer2_outputs[3597] = ~(layer1_outputs[9971]);
    assign layer2_outputs[3598] = layer1_outputs[8511];
    assign layer2_outputs[3599] = ~(layer1_outputs[4692]) | (layer1_outputs[7230]);
    assign layer2_outputs[3600] = ~(layer1_outputs[701]) | (layer1_outputs[9854]);
    assign layer2_outputs[3601] = (layer1_outputs[9456]) & ~(layer1_outputs[2788]);
    assign layer2_outputs[3602] = (layer1_outputs[4515]) | (layer1_outputs[2910]);
    assign layer2_outputs[3603] = ~(layer1_outputs[4634]);
    assign layer2_outputs[3604] = ~(layer1_outputs[9962]);
    assign layer2_outputs[3605] = ~(layer1_outputs[9684]);
    assign layer2_outputs[3606] = layer1_outputs[11338];
    assign layer2_outputs[3607] = ~((layer1_outputs[1047]) ^ (layer1_outputs[218]));
    assign layer2_outputs[3608] = ~((layer1_outputs[331]) | (layer1_outputs[5155]));
    assign layer2_outputs[3609] = (layer1_outputs[8681]) & (layer1_outputs[10414]);
    assign layer2_outputs[3610] = (layer1_outputs[8456]) & ~(layer1_outputs[5395]);
    assign layer2_outputs[3611] = (layer1_outputs[5071]) & ~(layer1_outputs[10785]);
    assign layer2_outputs[3612] = (layer1_outputs[4658]) & ~(layer1_outputs[11627]);
    assign layer2_outputs[3613] = ~(layer1_outputs[2343]);
    assign layer2_outputs[3614] = layer1_outputs[1210];
    assign layer2_outputs[3615] = (layer1_outputs[10846]) & ~(layer1_outputs[7025]);
    assign layer2_outputs[3616] = (layer1_outputs[3210]) | (layer1_outputs[4897]);
    assign layer2_outputs[3617] = (layer1_outputs[10686]) & ~(layer1_outputs[10150]);
    assign layer2_outputs[3618] = layer1_outputs[5233];
    assign layer2_outputs[3619] = (layer1_outputs[8570]) | (layer1_outputs[11592]);
    assign layer2_outputs[3620] = ~(layer1_outputs[982]);
    assign layer2_outputs[3621] = ~((layer1_outputs[11018]) ^ (layer1_outputs[5329]));
    assign layer2_outputs[3622] = layer1_outputs[5166];
    assign layer2_outputs[3623] = ~((layer1_outputs[12371]) | (layer1_outputs[5211]));
    assign layer2_outputs[3624] = (layer1_outputs[966]) & (layer1_outputs[1351]);
    assign layer2_outputs[3625] = (layer1_outputs[7673]) & (layer1_outputs[5062]);
    assign layer2_outputs[3626] = (layer1_outputs[11493]) ^ (layer1_outputs[8117]);
    assign layer2_outputs[3627] = ~(layer1_outputs[5983]);
    assign layer2_outputs[3628] = ~((layer1_outputs[4385]) ^ (layer1_outputs[10333]));
    assign layer2_outputs[3629] = ~(layer1_outputs[12215]);
    assign layer2_outputs[3630] = layer1_outputs[6055];
    assign layer2_outputs[3631] = ~(layer1_outputs[9492]);
    assign layer2_outputs[3632] = ~((layer1_outputs[7854]) & (layer1_outputs[5424]));
    assign layer2_outputs[3633] = layer1_outputs[5018];
    assign layer2_outputs[3634] = (layer1_outputs[12056]) | (layer1_outputs[8591]);
    assign layer2_outputs[3635] = layer1_outputs[8986];
    assign layer2_outputs[3636] = ~(layer1_outputs[11253]);
    assign layer2_outputs[3637] = ~((layer1_outputs[8657]) | (layer1_outputs[7622]));
    assign layer2_outputs[3638] = layer1_outputs[5149];
    assign layer2_outputs[3639] = layer1_outputs[2249];
    assign layer2_outputs[3640] = ~((layer1_outputs[4918]) & (layer1_outputs[10083]));
    assign layer2_outputs[3641] = (layer1_outputs[10261]) & (layer1_outputs[10878]);
    assign layer2_outputs[3642] = layer1_outputs[392];
    assign layer2_outputs[3643] = ~(layer1_outputs[7501]);
    assign layer2_outputs[3644] = ~((layer1_outputs[3360]) & (layer1_outputs[5569]));
    assign layer2_outputs[3645] = ~(layer1_outputs[4828]);
    assign layer2_outputs[3646] = ~(layer1_outputs[1114]) | (layer1_outputs[6883]);
    assign layer2_outputs[3647] = layer1_outputs[4326];
    assign layer2_outputs[3648] = layer1_outputs[10836];
    assign layer2_outputs[3649] = ~(layer1_outputs[4526]);
    assign layer2_outputs[3650] = layer1_outputs[1503];
    assign layer2_outputs[3651] = ~(layer1_outputs[8610]);
    assign layer2_outputs[3652] = layer1_outputs[9407];
    assign layer2_outputs[3653] = (layer1_outputs[11199]) ^ (layer1_outputs[10925]);
    assign layer2_outputs[3654] = layer1_outputs[44];
    assign layer2_outputs[3655] = ~(layer1_outputs[960]);
    assign layer2_outputs[3656] = ~(layer1_outputs[10398]);
    assign layer2_outputs[3657] = ~(layer1_outputs[255]);
    assign layer2_outputs[3658] = ~(layer1_outputs[5299]);
    assign layer2_outputs[3659] = layer1_outputs[48];
    assign layer2_outputs[3660] = (layer1_outputs[7540]) & ~(layer1_outputs[8265]);
    assign layer2_outputs[3661] = ~(layer1_outputs[12025]);
    assign layer2_outputs[3662] = (layer1_outputs[3967]) & ~(layer1_outputs[192]);
    assign layer2_outputs[3663] = ~((layer1_outputs[5698]) & (layer1_outputs[5161]));
    assign layer2_outputs[3664] = ~((layer1_outputs[1825]) | (layer1_outputs[8523]));
    assign layer2_outputs[3665] = (layer1_outputs[9430]) & ~(layer1_outputs[1793]);
    assign layer2_outputs[3666] = (layer1_outputs[3412]) | (layer1_outputs[7340]);
    assign layer2_outputs[3667] = layer1_outputs[7346];
    assign layer2_outputs[3668] = ~((layer1_outputs[8307]) ^ (layer1_outputs[5227]));
    assign layer2_outputs[3669] = layer1_outputs[10884];
    assign layer2_outputs[3670] = ~((layer1_outputs[5601]) & (layer1_outputs[5860]));
    assign layer2_outputs[3671] = ~((layer1_outputs[9487]) ^ (layer1_outputs[10974]));
    assign layer2_outputs[3672] = ~((layer1_outputs[11748]) | (layer1_outputs[4957]));
    assign layer2_outputs[3673] = layer1_outputs[9867];
    assign layer2_outputs[3674] = ~(layer1_outputs[4797]) | (layer1_outputs[891]);
    assign layer2_outputs[3675] = ~(layer1_outputs[8376]) | (layer1_outputs[5614]);
    assign layer2_outputs[3676] = ~((layer1_outputs[10554]) & (layer1_outputs[8237]));
    assign layer2_outputs[3677] = 1'b0;
    assign layer2_outputs[3678] = layer1_outputs[10441];
    assign layer2_outputs[3679] = (layer1_outputs[10514]) & ~(layer1_outputs[506]);
    assign layer2_outputs[3680] = layer1_outputs[7273];
    assign layer2_outputs[3681] = layer1_outputs[5955];
    assign layer2_outputs[3682] = (layer1_outputs[12311]) & (layer1_outputs[11056]);
    assign layer2_outputs[3683] = (layer1_outputs[3766]) ^ (layer1_outputs[4251]);
    assign layer2_outputs[3684] = layer1_outputs[3432];
    assign layer2_outputs[3685] = (layer1_outputs[10254]) & (layer1_outputs[1938]);
    assign layer2_outputs[3686] = ~(layer1_outputs[6268]);
    assign layer2_outputs[3687] = ~(layer1_outputs[10727]);
    assign layer2_outputs[3688] = ~(layer1_outputs[6287]);
    assign layer2_outputs[3689] = (layer1_outputs[10863]) | (layer1_outputs[12772]);
    assign layer2_outputs[3690] = ~(layer1_outputs[10696]) | (layer1_outputs[2879]);
    assign layer2_outputs[3691] = ~(layer1_outputs[1925]);
    assign layer2_outputs[3692] = ~(layer1_outputs[3431]);
    assign layer2_outputs[3693] = ~(layer1_outputs[3687]);
    assign layer2_outputs[3694] = ~(layer1_outputs[6547]);
    assign layer2_outputs[3695] = layer1_outputs[4773];
    assign layer2_outputs[3696] = layer1_outputs[11913];
    assign layer2_outputs[3697] = layer1_outputs[8511];
    assign layer2_outputs[3698] = ~(layer1_outputs[12206]);
    assign layer2_outputs[3699] = ~(layer1_outputs[484]);
    assign layer2_outputs[3700] = layer1_outputs[2902];
    assign layer2_outputs[3701] = ~((layer1_outputs[11885]) ^ (layer1_outputs[1242]));
    assign layer2_outputs[3702] = (layer1_outputs[692]) | (layer1_outputs[4710]);
    assign layer2_outputs[3703] = (layer1_outputs[11356]) & ~(layer1_outputs[1913]);
    assign layer2_outputs[3704] = layer1_outputs[5926];
    assign layer2_outputs[3705] = ~(layer1_outputs[4964]);
    assign layer2_outputs[3706] = ~((layer1_outputs[470]) | (layer1_outputs[3181]));
    assign layer2_outputs[3707] = layer1_outputs[9315];
    assign layer2_outputs[3708] = ~(layer1_outputs[10544]);
    assign layer2_outputs[3709] = layer1_outputs[4601];
    assign layer2_outputs[3710] = (layer1_outputs[6308]) & ~(layer1_outputs[3137]);
    assign layer2_outputs[3711] = ~(layer1_outputs[425]) | (layer1_outputs[3692]);
    assign layer2_outputs[3712] = ~((layer1_outputs[1526]) | (layer1_outputs[7084]));
    assign layer2_outputs[3713] = layer1_outputs[9405];
    assign layer2_outputs[3714] = ~((layer1_outputs[7588]) | (layer1_outputs[12784]));
    assign layer2_outputs[3715] = ~(layer1_outputs[1821]);
    assign layer2_outputs[3716] = (layer1_outputs[5455]) ^ (layer1_outputs[12668]);
    assign layer2_outputs[3717] = (layer1_outputs[6043]) ^ (layer1_outputs[259]);
    assign layer2_outputs[3718] = (layer1_outputs[4754]) & (layer1_outputs[7844]);
    assign layer2_outputs[3719] = (layer1_outputs[4850]) | (layer1_outputs[7655]);
    assign layer2_outputs[3720] = ~((layer1_outputs[5201]) ^ (layer1_outputs[6027]));
    assign layer2_outputs[3721] = ~((layer1_outputs[8684]) & (layer1_outputs[5957]));
    assign layer2_outputs[3722] = ~(layer1_outputs[2030]);
    assign layer2_outputs[3723] = layer1_outputs[4739];
    assign layer2_outputs[3724] = ~(layer1_outputs[7079]);
    assign layer2_outputs[3725] = (layer1_outputs[275]) & ~(layer1_outputs[8385]);
    assign layer2_outputs[3726] = (layer1_outputs[10158]) ^ (layer1_outputs[11403]);
    assign layer2_outputs[3727] = ~(layer1_outputs[10013]);
    assign layer2_outputs[3728] = ~(layer1_outputs[4808]);
    assign layer2_outputs[3729] = layer1_outputs[2559];
    assign layer2_outputs[3730] = ~((layer1_outputs[10375]) ^ (layer1_outputs[9156]));
    assign layer2_outputs[3731] = layer1_outputs[4033];
    assign layer2_outputs[3732] = layer1_outputs[8414];
    assign layer2_outputs[3733] = (layer1_outputs[646]) & ~(layer1_outputs[5287]);
    assign layer2_outputs[3734] = ~((layer1_outputs[12200]) ^ (layer1_outputs[5297]));
    assign layer2_outputs[3735] = (layer1_outputs[3443]) & (layer1_outputs[1948]);
    assign layer2_outputs[3736] = (layer1_outputs[2155]) & ~(layer1_outputs[4795]);
    assign layer2_outputs[3737] = ~((layer1_outputs[7959]) | (layer1_outputs[3027]));
    assign layer2_outputs[3738] = ~(layer1_outputs[3832]);
    assign layer2_outputs[3739] = (layer1_outputs[10477]) ^ (layer1_outputs[7193]);
    assign layer2_outputs[3740] = ~(layer1_outputs[3554]);
    assign layer2_outputs[3741] = ~((layer1_outputs[10337]) & (layer1_outputs[11446]));
    assign layer2_outputs[3742] = layer1_outputs[7532];
    assign layer2_outputs[3743] = layer1_outputs[3119];
    assign layer2_outputs[3744] = (layer1_outputs[11874]) | (layer1_outputs[916]);
    assign layer2_outputs[3745] = ~(layer1_outputs[2364]);
    assign layer2_outputs[3746] = (layer1_outputs[2347]) & ~(layer1_outputs[137]);
    assign layer2_outputs[3747] = ~(layer1_outputs[2566]);
    assign layer2_outputs[3748] = ~((layer1_outputs[9000]) ^ (layer1_outputs[6694]));
    assign layer2_outputs[3749] = (layer1_outputs[2915]) & ~(layer1_outputs[10629]);
    assign layer2_outputs[3750] = layer1_outputs[6254];
    assign layer2_outputs[3751] = ~(layer1_outputs[7802]) | (layer1_outputs[6057]);
    assign layer2_outputs[3752] = (layer1_outputs[3838]) ^ (layer1_outputs[4955]);
    assign layer2_outputs[3753] = (layer1_outputs[1814]) | (layer1_outputs[11050]);
    assign layer2_outputs[3754] = ~(layer1_outputs[1024]);
    assign layer2_outputs[3755] = (layer1_outputs[5796]) & ~(layer1_outputs[9973]);
    assign layer2_outputs[3756] = ~((layer1_outputs[814]) | (layer1_outputs[11686]));
    assign layer2_outputs[3757] = (layer1_outputs[5627]) & ~(layer1_outputs[1761]);
    assign layer2_outputs[3758] = layer1_outputs[10755];
    assign layer2_outputs[3759] = (layer1_outputs[3983]) ^ (layer1_outputs[2269]);
    assign layer2_outputs[3760] = ~(layer1_outputs[1924]);
    assign layer2_outputs[3761] = ~(layer1_outputs[11131]) | (layer1_outputs[11388]);
    assign layer2_outputs[3762] = (layer1_outputs[4870]) & (layer1_outputs[5824]);
    assign layer2_outputs[3763] = ~(layer1_outputs[8693]);
    assign layer2_outputs[3764] = (layer1_outputs[8702]) | (layer1_outputs[3848]);
    assign layer2_outputs[3765] = ~(layer1_outputs[6748]);
    assign layer2_outputs[3766] = (layer1_outputs[534]) & ~(layer1_outputs[5468]);
    assign layer2_outputs[3767] = layer1_outputs[8589];
    assign layer2_outputs[3768] = ~((layer1_outputs[7081]) ^ (layer1_outputs[10239]));
    assign layer2_outputs[3769] = ~(layer1_outputs[5146]) | (layer1_outputs[2624]);
    assign layer2_outputs[3770] = layer1_outputs[6981];
    assign layer2_outputs[3771] = layer1_outputs[10821];
    assign layer2_outputs[3772] = (layer1_outputs[5295]) ^ (layer1_outputs[11813]);
    assign layer2_outputs[3773] = layer1_outputs[10176];
    assign layer2_outputs[3774] = layer1_outputs[1085];
    assign layer2_outputs[3775] = (layer1_outputs[8148]) & (layer1_outputs[12480]);
    assign layer2_outputs[3776] = (layer1_outputs[9098]) ^ (layer1_outputs[5811]);
    assign layer2_outputs[3777] = layer1_outputs[7386];
    assign layer2_outputs[3778] = (layer1_outputs[1652]) & ~(layer1_outputs[6471]);
    assign layer2_outputs[3779] = ~(layer1_outputs[11382]) | (layer1_outputs[8345]);
    assign layer2_outputs[3780] = ~((layer1_outputs[9534]) | (layer1_outputs[3579]));
    assign layer2_outputs[3781] = layer1_outputs[6659];
    assign layer2_outputs[3782] = layer1_outputs[1140];
    assign layer2_outputs[3783] = ~(layer1_outputs[8884]);
    assign layer2_outputs[3784] = (layer1_outputs[7451]) & (layer1_outputs[1744]);
    assign layer2_outputs[3785] = ~(layer1_outputs[6830]);
    assign layer2_outputs[3786] = layer1_outputs[9331];
    assign layer2_outputs[3787] = layer1_outputs[4876];
    assign layer2_outputs[3788] = ~(layer1_outputs[11256]);
    assign layer2_outputs[3789] = (layer1_outputs[3127]) & ~(layer1_outputs[5089]);
    assign layer2_outputs[3790] = (layer1_outputs[6431]) ^ (layer1_outputs[7541]);
    assign layer2_outputs[3791] = (layer1_outputs[3777]) & (layer1_outputs[9750]);
    assign layer2_outputs[3792] = ~((layer1_outputs[8228]) ^ (layer1_outputs[11949]));
    assign layer2_outputs[3793] = ~(layer1_outputs[10679]) | (layer1_outputs[9952]);
    assign layer2_outputs[3794] = ~(layer1_outputs[12613]);
    assign layer2_outputs[3795] = ~((layer1_outputs[5938]) & (layer1_outputs[3807]));
    assign layer2_outputs[3796] = ~(layer1_outputs[10549]);
    assign layer2_outputs[3797] = ~(layer1_outputs[2547]);
    assign layer2_outputs[3798] = ~(layer1_outputs[7555]);
    assign layer2_outputs[3799] = layer1_outputs[4570];
    assign layer2_outputs[3800] = layer1_outputs[10431];
    assign layer2_outputs[3801] = layer1_outputs[11808];
    assign layer2_outputs[3802] = layer1_outputs[6572];
    assign layer2_outputs[3803] = ~(layer1_outputs[3040]);
    assign layer2_outputs[3804] = layer1_outputs[10038];
    assign layer2_outputs[3805] = ~((layer1_outputs[3818]) ^ (layer1_outputs[10130]));
    assign layer2_outputs[3806] = ~((layer1_outputs[1582]) | (layer1_outputs[5103]));
    assign layer2_outputs[3807] = ~(layer1_outputs[4575]) | (layer1_outputs[5970]);
    assign layer2_outputs[3808] = (layer1_outputs[2163]) & (layer1_outputs[7815]);
    assign layer2_outputs[3809] = (layer1_outputs[3541]) ^ (layer1_outputs[10510]);
    assign layer2_outputs[3810] = ~(layer1_outputs[10538]);
    assign layer2_outputs[3811] = ~((layer1_outputs[9368]) | (layer1_outputs[466]));
    assign layer2_outputs[3812] = ~(layer1_outputs[1044]) | (layer1_outputs[6069]);
    assign layer2_outputs[3813] = ~((layer1_outputs[12170]) & (layer1_outputs[7269]));
    assign layer2_outputs[3814] = ~(layer1_outputs[85]);
    assign layer2_outputs[3815] = (layer1_outputs[2118]) & ~(layer1_outputs[8188]);
    assign layer2_outputs[3816] = (layer1_outputs[6217]) & ~(layer1_outputs[11529]);
    assign layer2_outputs[3817] = layer1_outputs[3864];
    assign layer2_outputs[3818] = layer1_outputs[7086];
    assign layer2_outputs[3819] = layer1_outputs[8673];
    assign layer2_outputs[3820] = ~((layer1_outputs[11037]) ^ (layer1_outputs[2625]));
    assign layer2_outputs[3821] = layer1_outputs[3937];
    assign layer2_outputs[3822] = layer1_outputs[12532];
    assign layer2_outputs[3823] = (layer1_outputs[10709]) & ~(layer1_outputs[2909]);
    assign layer2_outputs[3824] = ~(layer1_outputs[6437]) | (layer1_outputs[7200]);
    assign layer2_outputs[3825] = ~(layer1_outputs[586]);
    assign layer2_outputs[3826] = ~(layer1_outputs[2710]) | (layer1_outputs[6591]);
    assign layer2_outputs[3827] = ~(layer1_outputs[1040]) | (layer1_outputs[9412]);
    assign layer2_outputs[3828] = ~((layer1_outputs[11769]) | (layer1_outputs[9848]));
    assign layer2_outputs[3829] = ~(layer1_outputs[4525]) | (layer1_outputs[11883]);
    assign layer2_outputs[3830] = (layer1_outputs[11734]) ^ (layer1_outputs[4079]);
    assign layer2_outputs[3831] = 1'b0;
    assign layer2_outputs[3832] = (layer1_outputs[2445]) & (layer1_outputs[9661]);
    assign layer2_outputs[3833] = ~(layer1_outputs[6793]);
    assign layer2_outputs[3834] = ~(layer1_outputs[10290]);
    assign layer2_outputs[3835] = layer1_outputs[1031];
    assign layer2_outputs[3836] = ~(layer1_outputs[11341]);
    assign layer2_outputs[3837] = ~((layer1_outputs[2344]) & (layer1_outputs[2613]));
    assign layer2_outputs[3838] = ~(layer1_outputs[11441]);
    assign layer2_outputs[3839] = layer1_outputs[10715];
    assign layer2_outputs[3840] = (layer1_outputs[2352]) & ~(layer1_outputs[4066]);
    assign layer2_outputs[3841] = (layer1_outputs[5427]) ^ (layer1_outputs[7387]);
    assign layer2_outputs[3842] = ~(layer1_outputs[8246]);
    assign layer2_outputs[3843] = ~(layer1_outputs[3644]);
    assign layer2_outputs[3844] = layer1_outputs[12000];
    assign layer2_outputs[3845] = (layer1_outputs[5754]) ^ (layer1_outputs[5968]);
    assign layer2_outputs[3846] = ~(layer1_outputs[9826]);
    assign layer2_outputs[3847] = 1'b1;
    assign layer2_outputs[3848] = (layer1_outputs[4132]) ^ (layer1_outputs[10145]);
    assign layer2_outputs[3849] = ~(layer1_outputs[920]);
    assign layer2_outputs[3850] = (layer1_outputs[4198]) & (layer1_outputs[7057]);
    assign layer2_outputs[3851] = ~(layer1_outputs[7873]) | (layer1_outputs[1737]);
    assign layer2_outputs[3852] = ~(layer1_outputs[10911]);
    assign layer2_outputs[3853] = ~((layer1_outputs[8736]) | (layer1_outputs[11987]));
    assign layer2_outputs[3854] = ~((layer1_outputs[2832]) ^ (layer1_outputs[4803]));
    assign layer2_outputs[3855] = (layer1_outputs[1799]) | (layer1_outputs[10307]);
    assign layer2_outputs[3856] = ~(layer1_outputs[2531]);
    assign layer2_outputs[3857] = layer1_outputs[10762];
    assign layer2_outputs[3858] = ~(layer1_outputs[7952]);
    assign layer2_outputs[3859] = ~(layer1_outputs[6489]);
    assign layer2_outputs[3860] = ~(layer1_outputs[1456]);
    assign layer2_outputs[3861] = ~((layer1_outputs[5827]) & (layer1_outputs[12398]));
    assign layer2_outputs[3862] = ~(layer1_outputs[10760]);
    assign layer2_outputs[3863] = layer1_outputs[5214];
    assign layer2_outputs[3864] = layer1_outputs[9306];
    assign layer2_outputs[3865] = layer1_outputs[9613];
    assign layer2_outputs[3866] = (layer1_outputs[12458]) | (layer1_outputs[6825]);
    assign layer2_outputs[3867] = layer1_outputs[4289];
    assign layer2_outputs[3868] = ~(layer1_outputs[3700]);
    assign layer2_outputs[3869] = ~(layer1_outputs[12680]);
    assign layer2_outputs[3870] = ~((layer1_outputs[6032]) ^ (layer1_outputs[11248]));
    assign layer2_outputs[3871] = ~((layer1_outputs[3263]) ^ (layer1_outputs[7167]));
    assign layer2_outputs[3872] = ~(layer1_outputs[11]);
    assign layer2_outputs[3873] = ~(layer1_outputs[9284]);
    assign layer2_outputs[3874] = ~(layer1_outputs[9036]);
    assign layer2_outputs[3875] = ~((layer1_outputs[8819]) | (layer1_outputs[6526]));
    assign layer2_outputs[3876] = (layer1_outputs[6971]) ^ (layer1_outputs[3683]);
    assign layer2_outputs[3877] = (layer1_outputs[3433]) ^ (layer1_outputs[2266]);
    assign layer2_outputs[3878] = ~(layer1_outputs[973]);
    assign layer2_outputs[3879] = (layer1_outputs[1117]) | (layer1_outputs[1125]);
    assign layer2_outputs[3880] = ~((layer1_outputs[3383]) ^ (layer1_outputs[5924]));
    assign layer2_outputs[3881] = (layer1_outputs[4940]) & ~(layer1_outputs[4303]);
    assign layer2_outputs[3882] = layer1_outputs[10088];
    assign layer2_outputs[3883] = layer1_outputs[155];
    assign layer2_outputs[3884] = ~((layer1_outputs[4292]) & (layer1_outputs[8614]));
    assign layer2_outputs[3885] = ~((layer1_outputs[4862]) & (layer1_outputs[4526]));
    assign layer2_outputs[3886] = ~(layer1_outputs[7847]);
    assign layer2_outputs[3887] = ~((layer1_outputs[7641]) | (layer1_outputs[3569]));
    assign layer2_outputs[3888] = (layer1_outputs[5355]) ^ (layer1_outputs[5027]);
    assign layer2_outputs[3889] = ~(layer1_outputs[7566]) | (layer1_outputs[1263]);
    assign layer2_outputs[3890] = layer1_outputs[5721];
    assign layer2_outputs[3891] = ~((layer1_outputs[4734]) | (layer1_outputs[3667]));
    assign layer2_outputs[3892] = ~(layer1_outputs[2316]);
    assign layer2_outputs[3893] = (layer1_outputs[5057]) & ~(layer1_outputs[4806]);
    assign layer2_outputs[3894] = layer1_outputs[7043];
    assign layer2_outputs[3895] = layer1_outputs[10266];
    assign layer2_outputs[3896] = (layer1_outputs[9969]) ^ (layer1_outputs[2853]);
    assign layer2_outputs[3897] = ~(layer1_outputs[3649]);
    assign layer2_outputs[3898] = ~(layer1_outputs[768]);
    assign layer2_outputs[3899] = ~((layer1_outputs[11545]) ^ (layer1_outputs[9856]));
    assign layer2_outputs[3900] = (layer1_outputs[9250]) | (layer1_outputs[947]);
    assign layer2_outputs[3901] = ~(layer1_outputs[4531]);
    assign layer2_outputs[3902] = ~((layer1_outputs[4193]) ^ (layer1_outputs[6105]));
    assign layer2_outputs[3903] = ~(layer1_outputs[4414]);
    assign layer2_outputs[3904] = ~(layer1_outputs[9378]);
    assign layer2_outputs[3905] = ~((layer1_outputs[9610]) ^ (layer1_outputs[2979]));
    assign layer2_outputs[3906] = ~(layer1_outputs[12453]);
    assign layer2_outputs[3907] = ~((layer1_outputs[3655]) ^ (layer1_outputs[10229]));
    assign layer2_outputs[3908] = ~(layer1_outputs[8421]) | (layer1_outputs[5802]);
    assign layer2_outputs[3909] = (layer1_outputs[4017]) | (layer1_outputs[11524]);
    assign layer2_outputs[3910] = ~((layer1_outputs[5842]) ^ (layer1_outputs[4264]));
    assign layer2_outputs[3911] = ~(layer1_outputs[397]);
    assign layer2_outputs[3912] = 1'b1;
    assign layer2_outputs[3913] = (layer1_outputs[8436]) ^ (layer1_outputs[532]);
    assign layer2_outputs[3914] = layer1_outputs[10591];
    assign layer2_outputs[3915] = ~(layer1_outputs[9842]);
    assign layer2_outputs[3916] = layer1_outputs[9532];
    assign layer2_outputs[3917] = ~(layer1_outputs[1735]);
    assign layer2_outputs[3918] = ~(layer1_outputs[4308]) | (layer1_outputs[5065]);
    assign layer2_outputs[3919] = ~(layer1_outputs[541]) | (layer1_outputs[10476]);
    assign layer2_outputs[3920] = layer1_outputs[682];
    assign layer2_outputs[3921] = (layer1_outputs[8133]) & (layer1_outputs[4472]);
    assign layer2_outputs[3922] = ~(layer1_outputs[12207]);
    assign layer2_outputs[3923] = ~(layer1_outputs[9653]);
    assign layer2_outputs[3924] = ~(layer1_outputs[7509]);
    assign layer2_outputs[3925] = ~(layer1_outputs[12715]);
    assign layer2_outputs[3926] = ~((layer1_outputs[12725]) | (layer1_outputs[9376]));
    assign layer2_outputs[3927] = ~(layer1_outputs[12641]);
    assign layer2_outputs[3928] = layer1_outputs[5050];
    assign layer2_outputs[3929] = (layer1_outputs[8051]) | (layer1_outputs[7790]);
    assign layer2_outputs[3930] = ~((layer1_outputs[930]) ^ (layer1_outputs[12076]));
    assign layer2_outputs[3931] = ~((layer1_outputs[10019]) | (layer1_outputs[4678]));
    assign layer2_outputs[3932] = ~(layer1_outputs[9078]);
    assign layer2_outputs[3933] = layer1_outputs[4003];
    assign layer2_outputs[3934] = ~(layer1_outputs[2963]) | (layer1_outputs[11337]);
    assign layer2_outputs[3935] = (layer1_outputs[2391]) & ~(layer1_outputs[5272]);
    assign layer2_outputs[3936] = layer1_outputs[983];
    assign layer2_outputs[3937] = (layer1_outputs[6205]) & ~(layer1_outputs[3707]);
    assign layer2_outputs[3938] = ~((layer1_outputs[3510]) | (layer1_outputs[7287]));
    assign layer2_outputs[3939] = layer1_outputs[199];
    assign layer2_outputs[3940] = ~((layer1_outputs[5374]) & (layer1_outputs[152]));
    assign layer2_outputs[3941] = ~(layer1_outputs[2482]);
    assign layer2_outputs[3942] = ~((layer1_outputs[2587]) ^ (layer1_outputs[3784]));
    assign layer2_outputs[3943] = ~(layer1_outputs[2919]);
    assign layer2_outputs[3944] = ~(layer1_outputs[1576]);
    assign layer2_outputs[3945] = layer1_outputs[4206];
    assign layer2_outputs[3946] = ~(layer1_outputs[10103]);
    assign layer2_outputs[3947] = layer1_outputs[927];
    assign layer2_outputs[3948] = ~(layer1_outputs[2405]);
    assign layer2_outputs[3949] = ~(layer1_outputs[2324]) | (layer1_outputs[638]);
    assign layer2_outputs[3950] = 1'b1;
    assign layer2_outputs[3951] = 1'b0;
    assign layer2_outputs[3952] = ~(layer1_outputs[4682]);
    assign layer2_outputs[3953] = ~(layer1_outputs[5025]) | (layer1_outputs[5584]);
    assign layer2_outputs[3954] = ~(layer1_outputs[4459]) | (layer1_outputs[5438]);
    assign layer2_outputs[3955] = ~((layer1_outputs[8000]) | (layer1_outputs[9500]));
    assign layer2_outputs[3956] = ~((layer1_outputs[98]) ^ (layer1_outputs[10198]));
    assign layer2_outputs[3957] = ~(layer1_outputs[1203]);
    assign layer2_outputs[3958] = ~(layer1_outputs[8829]);
    assign layer2_outputs[3959] = ~(layer1_outputs[10427]) | (layer1_outputs[5211]);
    assign layer2_outputs[3960] = ~((layer1_outputs[322]) | (layer1_outputs[9795]));
    assign layer2_outputs[3961] = (layer1_outputs[1887]) ^ (layer1_outputs[11567]);
    assign layer2_outputs[3962] = ~(layer1_outputs[362]) | (layer1_outputs[3275]);
    assign layer2_outputs[3963] = (layer1_outputs[3107]) & ~(layer1_outputs[886]);
    assign layer2_outputs[3964] = (layer1_outputs[11810]) & ~(layer1_outputs[2143]);
    assign layer2_outputs[3965] = ~((layer1_outputs[10624]) ^ (layer1_outputs[6833]));
    assign layer2_outputs[3966] = ~((layer1_outputs[11117]) ^ (layer1_outputs[11238]));
    assign layer2_outputs[3967] = ~(layer1_outputs[5581]) | (layer1_outputs[7753]);
    assign layer2_outputs[3968] = (layer1_outputs[1748]) | (layer1_outputs[4450]);
    assign layer2_outputs[3969] = ~(layer1_outputs[4409]);
    assign layer2_outputs[3970] = (layer1_outputs[2119]) & (layer1_outputs[1813]);
    assign layer2_outputs[3971] = (layer1_outputs[202]) & ~(layer1_outputs[9067]);
    assign layer2_outputs[3972] = ~(layer1_outputs[12044]);
    assign layer2_outputs[3973] = layer1_outputs[7124];
    assign layer2_outputs[3974] = (layer1_outputs[7979]) & ~(layer1_outputs[1488]);
    assign layer2_outputs[3975] = ~(layer1_outputs[10336]);
    assign layer2_outputs[3976] = ~(layer1_outputs[8130]);
    assign layer2_outputs[3977] = layer1_outputs[5644];
    assign layer2_outputs[3978] = ~(layer1_outputs[3754]) | (layer1_outputs[822]);
    assign layer2_outputs[3979] = ~(layer1_outputs[10416]);
    assign layer2_outputs[3980] = ~((layer1_outputs[12376]) & (layer1_outputs[5559]));
    assign layer2_outputs[3981] = layer1_outputs[293];
    assign layer2_outputs[3982] = layer1_outputs[8807];
    assign layer2_outputs[3983] = layer1_outputs[6214];
    assign layer2_outputs[3984] = layer1_outputs[5656];
    assign layer2_outputs[3985] = ~((layer1_outputs[3627]) ^ (layer1_outputs[2865]));
    assign layer2_outputs[3986] = layer1_outputs[7443];
    assign layer2_outputs[3987] = ~((layer1_outputs[6942]) ^ (layer1_outputs[12734]));
    assign layer2_outputs[3988] = (layer1_outputs[5266]) ^ (layer1_outputs[6260]);
    assign layer2_outputs[3989] = ~(layer1_outputs[10487]);
    assign layer2_outputs[3990] = (layer1_outputs[8544]) | (layer1_outputs[2149]);
    assign layer2_outputs[3991] = ~(layer1_outputs[10467]);
    assign layer2_outputs[3992] = layer1_outputs[5967];
    assign layer2_outputs[3993] = (layer1_outputs[1886]) ^ (layer1_outputs[5880]);
    assign layer2_outputs[3994] = ~(layer1_outputs[263]);
    assign layer2_outputs[3995] = (layer1_outputs[10012]) ^ (layer1_outputs[1599]);
    assign layer2_outputs[3996] = ~(layer1_outputs[1375]) | (layer1_outputs[3131]);
    assign layer2_outputs[3997] = layer1_outputs[2891];
    assign layer2_outputs[3998] = ~(layer1_outputs[10574]);
    assign layer2_outputs[3999] = layer1_outputs[6841];
    assign layer2_outputs[4000] = ~(layer1_outputs[1387]) | (layer1_outputs[5107]);
    assign layer2_outputs[4001] = ~(layer1_outputs[808]);
    assign layer2_outputs[4002] = layer1_outputs[8920];
    assign layer2_outputs[4003] = (layer1_outputs[1570]) | (layer1_outputs[7677]);
    assign layer2_outputs[4004] = layer1_outputs[3382];
    assign layer2_outputs[4005] = ~(layer1_outputs[2468]);
    assign layer2_outputs[4006] = ~((layer1_outputs[9477]) & (layer1_outputs[2878]));
    assign layer2_outputs[4007] = ~(layer1_outputs[8745]);
    assign layer2_outputs[4008] = layer1_outputs[8356];
    assign layer2_outputs[4009] = layer1_outputs[2546];
    assign layer2_outputs[4010] = layer1_outputs[1036];
    assign layer2_outputs[4011] = ~(layer1_outputs[3899]);
    assign layer2_outputs[4012] = ~(layer1_outputs[764]);
    assign layer2_outputs[4013] = (layer1_outputs[7915]) ^ (layer1_outputs[2079]);
    assign layer2_outputs[4014] = ~(layer1_outputs[5656]) | (layer1_outputs[6183]);
    assign layer2_outputs[4015] = ~(layer1_outputs[6757]) | (layer1_outputs[4998]);
    assign layer2_outputs[4016] = ~((layer1_outputs[10875]) ^ (layer1_outputs[1077]));
    assign layer2_outputs[4017] = ~((layer1_outputs[1369]) & (layer1_outputs[8616]));
    assign layer2_outputs[4018] = ~(layer1_outputs[9370]);
    assign layer2_outputs[4019] = (layer1_outputs[10018]) & (layer1_outputs[511]);
    assign layer2_outputs[4020] = ~(layer1_outputs[3671]);
    assign layer2_outputs[4021] = ~(layer1_outputs[2385]);
    assign layer2_outputs[4022] = ~(layer1_outputs[6866]);
    assign layer2_outputs[4023] = ~((layer1_outputs[4197]) ^ (layer1_outputs[5792]));
    assign layer2_outputs[4024] = layer1_outputs[6648];
    assign layer2_outputs[4025] = ~((layer1_outputs[738]) & (layer1_outputs[12339]));
    assign layer2_outputs[4026] = layer1_outputs[3278];
    assign layer2_outputs[4027] = ~(layer1_outputs[1630]);
    assign layer2_outputs[4028] = layer1_outputs[892];
    assign layer2_outputs[4029] = layer1_outputs[10033];
    assign layer2_outputs[4030] = ~(layer1_outputs[1569]);
    assign layer2_outputs[4031] = (layer1_outputs[5903]) | (layer1_outputs[1025]);
    assign layer2_outputs[4032] = (layer1_outputs[9442]) & ~(layer1_outputs[12554]);
    assign layer2_outputs[4033] = ~(layer1_outputs[4872]);
    assign layer2_outputs[4034] = ~(layer1_outputs[1822]);
    assign layer2_outputs[4035] = layer1_outputs[722];
    assign layer2_outputs[4036] = (layer1_outputs[795]) & (layer1_outputs[8571]);
    assign layer2_outputs[4037] = layer1_outputs[435];
    assign layer2_outputs[4038] = ~(layer1_outputs[11031]) | (layer1_outputs[1381]);
    assign layer2_outputs[4039] = ~(layer1_outputs[10328]);
    assign layer2_outputs[4040] = (layer1_outputs[1292]) ^ (layer1_outputs[2083]);
    assign layer2_outputs[4041] = ~(layer1_outputs[4730]);
    assign layer2_outputs[4042] = ~((layer1_outputs[11999]) & (layer1_outputs[7821]));
    assign layer2_outputs[4043] = ~(layer1_outputs[9693]) | (layer1_outputs[11911]);
    assign layer2_outputs[4044] = layer1_outputs[4695];
    assign layer2_outputs[4045] = (layer1_outputs[9414]) ^ (layer1_outputs[3110]);
    assign layer2_outputs[4046] = (layer1_outputs[6178]) | (layer1_outputs[1819]);
    assign layer2_outputs[4047] = (layer1_outputs[6125]) ^ (layer1_outputs[9844]);
    assign layer2_outputs[4048] = ~((layer1_outputs[428]) & (layer1_outputs[9623]));
    assign layer2_outputs[4049] = ~(layer1_outputs[3115]);
    assign layer2_outputs[4050] = ~(layer1_outputs[4532]);
    assign layer2_outputs[4051] = (layer1_outputs[11006]) & ~(layer1_outputs[4681]);
    assign layer2_outputs[4052] = ~(layer1_outputs[10857]);
    assign layer2_outputs[4053] = (layer1_outputs[12247]) | (layer1_outputs[9114]);
    assign layer2_outputs[4054] = ~(layer1_outputs[8458]);
    assign layer2_outputs[4055] = ~((layer1_outputs[3353]) | (layer1_outputs[11331]));
    assign layer2_outputs[4056] = ~(layer1_outputs[12619]) | (layer1_outputs[6413]);
    assign layer2_outputs[4057] = layer1_outputs[1451];
    assign layer2_outputs[4058] = ~(layer1_outputs[10578]);
    assign layer2_outputs[4059] = ~(layer1_outputs[9175]);
    assign layer2_outputs[4060] = ~(layer1_outputs[2660]);
    assign layer2_outputs[4061] = ~((layer1_outputs[9615]) ^ (layer1_outputs[11225]));
    assign layer2_outputs[4062] = ~(layer1_outputs[5570]);
    assign layer2_outputs[4063] = ~(layer1_outputs[11572]);
    assign layer2_outputs[4064] = ~(layer1_outputs[7639]) | (layer1_outputs[8450]);
    assign layer2_outputs[4065] = (layer1_outputs[7507]) & ~(layer1_outputs[1755]);
    assign layer2_outputs[4066] = ~((layer1_outputs[9298]) | (layer1_outputs[12713]));
    assign layer2_outputs[4067] = (layer1_outputs[9132]) ^ (layer1_outputs[11717]);
    assign layer2_outputs[4068] = (layer1_outputs[1059]) | (layer1_outputs[6087]);
    assign layer2_outputs[4069] = layer1_outputs[8481];
    assign layer2_outputs[4070] = layer1_outputs[229];
    assign layer2_outputs[4071] = ~((layer1_outputs[974]) | (layer1_outputs[10007]));
    assign layer2_outputs[4072] = ~(layer1_outputs[8118]);
    assign layer2_outputs[4073] = ~(layer1_outputs[5580]);
    assign layer2_outputs[4074] = ~((layer1_outputs[12380]) ^ (layer1_outputs[12227]));
    assign layer2_outputs[4075] = (layer1_outputs[5788]) | (layer1_outputs[8301]);
    assign layer2_outputs[4076] = layer1_outputs[2775];
    assign layer2_outputs[4077] = layer1_outputs[840];
    assign layer2_outputs[4078] = (layer1_outputs[6127]) & (layer1_outputs[2033]);
    assign layer2_outputs[4079] = (layer1_outputs[1155]) ^ (layer1_outputs[12143]);
    assign layer2_outputs[4080] = ~((layer1_outputs[1316]) ^ (layer1_outputs[1468]));
    assign layer2_outputs[4081] = (layer1_outputs[8213]) & (layer1_outputs[3725]);
    assign layer2_outputs[4082] = ~((layer1_outputs[47]) & (layer1_outputs[3200]));
    assign layer2_outputs[4083] = (layer1_outputs[2921]) & ~(layer1_outputs[7763]);
    assign layer2_outputs[4084] = ~(layer1_outputs[5780]) | (layer1_outputs[9361]);
    assign layer2_outputs[4085] = ~((layer1_outputs[11]) | (layer1_outputs[8283]));
    assign layer2_outputs[4086] = (layer1_outputs[8438]) ^ (layer1_outputs[10744]);
    assign layer2_outputs[4087] = ~(layer1_outputs[8682]);
    assign layer2_outputs[4088] = layer1_outputs[1011];
    assign layer2_outputs[4089] = layer1_outputs[5204];
    assign layer2_outputs[4090] = ~((layer1_outputs[2003]) ^ (layer1_outputs[3758]));
    assign layer2_outputs[4091] = ~((layer1_outputs[9300]) & (layer1_outputs[11839]));
    assign layer2_outputs[4092] = ~(layer1_outputs[4275]);
    assign layer2_outputs[4093] = 1'b0;
    assign layer2_outputs[4094] = ~(layer1_outputs[6211]);
    assign layer2_outputs[4095] = layer1_outputs[3519];
    assign layer2_outputs[4096] = ~(layer1_outputs[11265]) | (layer1_outputs[4508]);
    assign layer2_outputs[4097] = ~(layer1_outputs[8850]);
    assign layer2_outputs[4098] = layer1_outputs[4673];
    assign layer2_outputs[4099] = ~((layer1_outputs[1016]) & (layer1_outputs[12295]));
    assign layer2_outputs[4100] = (layer1_outputs[2376]) & ~(layer1_outputs[8577]);
    assign layer2_outputs[4101] = ~((layer1_outputs[7231]) ^ (layer1_outputs[4193]));
    assign layer2_outputs[4102] = ~(layer1_outputs[7277]);
    assign layer2_outputs[4103] = (layer1_outputs[3064]) & ~(layer1_outputs[3718]);
    assign layer2_outputs[4104] = (layer1_outputs[2833]) ^ (layer1_outputs[1862]);
    assign layer2_outputs[4105] = layer1_outputs[6786];
    assign layer2_outputs[4106] = ~(layer1_outputs[4170]);
    assign layer2_outputs[4107] = ~(layer1_outputs[8340]);
    assign layer2_outputs[4108] = layer1_outputs[8324];
    assign layer2_outputs[4109] = ~((layer1_outputs[9615]) | (layer1_outputs[1834]));
    assign layer2_outputs[4110] = ~((layer1_outputs[12460]) & (layer1_outputs[2102]));
    assign layer2_outputs[4111] = layer1_outputs[1333];
    assign layer2_outputs[4112] = ~(layer1_outputs[334]) | (layer1_outputs[512]);
    assign layer2_outputs[4113] = ~((layer1_outputs[4862]) & (layer1_outputs[53]));
    assign layer2_outputs[4114] = layer1_outputs[3717];
    assign layer2_outputs[4115] = layer1_outputs[6732];
    assign layer2_outputs[4116] = layer1_outputs[5172];
    assign layer2_outputs[4117] = ~(layer1_outputs[12744]) | (layer1_outputs[5940]);
    assign layer2_outputs[4118] = layer1_outputs[4323];
    assign layer2_outputs[4119] = (layer1_outputs[5671]) ^ (layer1_outputs[2814]);
    assign layer2_outputs[4120] = layer1_outputs[8096];
    assign layer2_outputs[4121] = ~(layer1_outputs[1019]) | (layer1_outputs[7966]);
    assign layer2_outputs[4122] = (layer1_outputs[11794]) & ~(layer1_outputs[5361]);
    assign layer2_outputs[4123] = ~((layer1_outputs[6534]) | (layer1_outputs[5359]));
    assign layer2_outputs[4124] = 1'b0;
    assign layer2_outputs[4125] = (layer1_outputs[7056]) ^ (layer1_outputs[1145]);
    assign layer2_outputs[4126] = ~(layer1_outputs[470]);
    assign layer2_outputs[4127] = layer1_outputs[7880];
    assign layer2_outputs[4128] = layer1_outputs[6402];
    assign layer2_outputs[4129] = ~(layer1_outputs[9697]);
    assign layer2_outputs[4130] = ~(layer1_outputs[5291]);
    assign layer2_outputs[4131] = ~(layer1_outputs[8018]);
    assign layer2_outputs[4132] = ~((layer1_outputs[327]) ^ (layer1_outputs[4835]));
    assign layer2_outputs[4133] = layer1_outputs[2031];
    assign layer2_outputs[4134] = layer1_outputs[3764];
    assign layer2_outputs[4135] = ~(layer1_outputs[3216]);
    assign layer2_outputs[4136] = ~((layer1_outputs[114]) & (layer1_outputs[10810]));
    assign layer2_outputs[4137] = ~(layer1_outputs[50]);
    assign layer2_outputs[4138] = (layer1_outputs[4826]) ^ (layer1_outputs[764]);
    assign layer2_outputs[4139] = (layer1_outputs[3558]) | (layer1_outputs[2688]);
    assign layer2_outputs[4140] = ~(layer1_outputs[5854]) | (layer1_outputs[11980]);
    assign layer2_outputs[4141] = ~((layer1_outputs[6704]) | (layer1_outputs[1400]));
    assign layer2_outputs[4142] = ~(layer1_outputs[2308]) | (layer1_outputs[3666]);
    assign layer2_outputs[4143] = ~((layer1_outputs[1703]) & (layer1_outputs[2977]));
    assign layer2_outputs[4144] = ~((layer1_outputs[12681]) | (layer1_outputs[7770]));
    assign layer2_outputs[4145] = (layer1_outputs[893]) | (layer1_outputs[234]);
    assign layer2_outputs[4146] = ~((layer1_outputs[3143]) | (layer1_outputs[4993]));
    assign layer2_outputs[4147] = ~(layer1_outputs[8542]) | (layer1_outputs[1663]);
    assign layer2_outputs[4148] = (layer1_outputs[8745]) & (layer1_outputs[9888]);
    assign layer2_outputs[4149] = (layer1_outputs[1323]) | (layer1_outputs[7160]);
    assign layer2_outputs[4150] = layer1_outputs[10840];
    assign layer2_outputs[4151] = layer1_outputs[208];
    assign layer2_outputs[4152] = ~(layer1_outputs[10367]);
    assign layer2_outputs[4153] = (layer1_outputs[10115]) | (layer1_outputs[1617]);
    assign layer2_outputs[4154] = ~(layer1_outputs[9006]);
    assign layer2_outputs[4155] = layer1_outputs[1340];
    assign layer2_outputs[4156] = ~(layer1_outputs[10929]);
    assign layer2_outputs[4157] = layer1_outputs[2116];
    assign layer2_outputs[4158] = ~(layer1_outputs[12076]);
    assign layer2_outputs[4159] = ~(layer1_outputs[1243]) | (layer1_outputs[5980]);
    assign layer2_outputs[4160] = ~(layer1_outputs[9464]);
    assign layer2_outputs[4161] = ~((layer1_outputs[11969]) | (layer1_outputs[4884]));
    assign layer2_outputs[4162] = ~(layer1_outputs[11315]);
    assign layer2_outputs[4163] = ~(layer1_outputs[12026]);
    assign layer2_outputs[4164] = ~(layer1_outputs[9854]) | (layer1_outputs[9024]);
    assign layer2_outputs[4165] = ~(layer1_outputs[1007]);
    assign layer2_outputs[4166] = layer1_outputs[414];
    assign layer2_outputs[4167] = (layer1_outputs[7023]) ^ (layer1_outputs[265]);
    assign layer2_outputs[4168] = ~(layer1_outputs[3065]);
    assign layer2_outputs[4169] = (layer1_outputs[1859]) & ~(layer1_outputs[4671]);
    assign layer2_outputs[4170] = ~((layer1_outputs[5574]) | (layer1_outputs[6633]));
    assign layer2_outputs[4171] = ~((layer1_outputs[9951]) | (layer1_outputs[6926]));
    assign layer2_outputs[4172] = (layer1_outputs[28]) ^ (layer1_outputs[5847]);
    assign layer2_outputs[4173] = layer1_outputs[11646];
    assign layer2_outputs[4174] = ~((layer1_outputs[3543]) ^ (layer1_outputs[8713]));
    assign layer2_outputs[4175] = ~((layer1_outputs[3177]) ^ (layer1_outputs[11228]));
    assign layer2_outputs[4176] = (layer1_outputs[10367]) | (layer1_outputs[7005]);
    assign layer2_outputs[4177] = ~(layer1_outputs[6465]);
    assign layer2_outputs[4178] = ~(layer1_outputs[11786]);
    assign layer2_outputs[4179] = layer1_outputs[3830];
    assign layer2_outputs[4180] = layer1_outputs[10804];
    assign layer2_outputs[4181] = ~((layer1_outputs[6611]) & (layer1_outputs[5076]));
    assign layer2_outputs[4182] = (layer1_outputs[9815]) & (layer1_outputs[11848]);
    assign layer2_outputs[4183] = ~(layer1_outputs[12211]);
    assign layer2_outputs[4184] = layer1_outputs[5984];
    assign layer2_outputs[4185] = layer1_outputs[11633];
    assign layer2_outputs[4186] = ~(layer1_outputs[8602]);
    assign layer2_outputs[4187] = layer1_outputs[12384];
    assign layer2_outputs[4188] = ~(layer1_outputs[2404]);
    assign layer2_outputs[4189] = ~(layer1_outputs[7545]);
    assign layer2_outputs[4190] = (layer1_outputs[4668]) ^ (layer1_outputs[1845]);
    assign layer2_outputs[4191] = ~(layer1_outputs[73]);
    assign layer2_outputs[4192] = (layer1_outputs[6753]) & (layer1_outputs[3503]);
    assign layer2_outputs[4193] = (layer1_outputs[3670]) & (layer1_outputs[11522]);
    assign layer2_outputs[4194] = ~((layer1_outputs[7581]) & (layer1_outputs[8190]));
    assign layer2_outputs[4195] = (layer1_outputs[4227]) & (layer1_outputs[10050]);
    assign layer2_outputs[4196] = (layer1_outputs[10302]) & (layer1_outputs[7081]);
    assign layer2_outputs[4197] = ~(layer1_outputs[1412]) | (layer1_outputs[9859]);
    assign layer2_outputs[4198] = ~(layer1_outputs[4336]) | (layer1_outputs[4896]);
    assign layer2_outputs[4199] = (layer1_outputs[8288]) & ~(layer1_outputs[5409]);
    assign layer2_outputs[4200] = ~(layer1_outputs[10494]);
    assign layer2_outputs[4201] = ~(layer1_outputs[876]) | (layer1_outputs[11300]);
    assign layer2_outputs[4202] = ~(layer1_outputs[5917]);
    assign layer2_outputs[4203] = layer1_outputs[11702];
    assign layer2_outputs[4204] = layer1_outputs[2381];
    assign layer2_outputs[4205] = layer1_outputs[1874];
    assign layer2_outputs[4206] = layer1_outputs[12094];
    assign layer2_outputs[4207] = ~(layer1_outputs[2474]);
    assign layer2_outputs[4208] = (layer1_outputs[2653]) ^ (layer1_outputs[8943]);
    assign layer2_outputs[4209] = (layer1_outputs[11367]) & ~(layer1_outputs[4898]);
    assign layer2_outputs[4210] = layer1_outputs[306];
    assign layer2_outputs[4211] = layer1_outputs[9383];
    assign layer2_outputs[4212] = (layer1_outputs[4566]) & (layer1_outputs[4015]);
    assign layer2_outputs[4213] = ~(layer1_outputs[11015]) | (layer1_outputs[9759]);
    assign layer2_outputs[4214] = layer1_outputs[9301];
    assign layer2_outputs[4215] = (layer1_outputs[11210]) & (layer1_outputs[6031]);
    assign layer2_outputs[4216] = layer1_outputs[7985];
    assign layer2_outputs[4217] = (layer1_outputs[11554]) & (layer1_outputs[658]);
    assign layer2_outputs[4218] = ~(layer1_outputs[11321]);
    assign layer2_outputs[4219] = layer1_outputs[1029];
    assign layer2_outputs[4220] = (layer1_outputs[7905]) | (layer1_outputs[9213]);
    assign layer2_outputs[4221] = layer1_outputs[6116];
    assign layer2_outputs[4222] = ~((layer1_outputs[8675]) ^ (layer1_outputs[8904]));
    assign layer2_outputs[4223] = ~(layer1_outputs[8935]);
    assign layer2_outputs[4224] = layer1_outputs[12190];
    assign layer2_outputs[4225] = ~(layer1_outputs[12773]) | (layer1_outputs[5964]);
    assign layer2_outputs[4226] = (layer1_outputs[12106]) & ~(layer1_outputs[12658]);
    assign layer2_outputs[4227] = layer1_outputs[6470];
    assign layer2_outputs[4228] = ~((layer1_outputs[10006]) ^ (layer1_outputs[7164]));
    assign layer2_outputs[4229] = layer1_outputs[9100];
    assign layer2_outputs[4230] = ~(layer1_outputs[11677]);
    assign layer2_outputs[4231] = (layer1_outputs[374]) | (layer1_outputs[6605]);
    assign layer2_outputs[4232] = layer1_outputs[7059];
    assign layer2_outputs[4233] = layer1_outputs[1419];
    assign layer2_outputs[4234] = ~(layer1_outputs[3644]);
    assign layer2_outputs[4235] = (layer1_outputs[10397]) & ~(layer1_outputs[6312]);
    assign layer2_outputs[4236] = layer1_outputs[5704];
    assign layer2_outputs[4237] = ~(layer1_outputs[9475]) | (layer1_outputs[6548]);
    assign layer2_outputs[4238] = ~((layer1_outputs[11896]) ^ (layer1_outputs[9051]));
    assign layer2_outputs[4239] = ~((layer1_outputs[7172]) ^ (layer1_outputs[4429]));
    assign layer2_outputs[4240] = (layer1_outputs[12166]) & (layer1_outputs[11690]);
    assign layer2_outputs[4241] = ~(layer1_outputs[1127]) | (layer1_outputs[7162]);
    assign layer2_outputs[4242] = ~(layer1_outputs[11730]);
    assign layer2_outputs[4243] = ~(layer1_outputs[10116]) | (layer1_outputs[12346]);
    assign layer2_outputs[4244] = (layer1_outputs[11532]) ^ (layer1_outputs[12134]);
    assign layer2_outputs[4245] = (layer1_outputs[4948]) | (layer1_outputs[12350]);
    assign layer2_outputs[4246] = (layer1_outputs[2159]) | (layer1_outputs[12191]);
    assign layer2_outputs[4247] = ~(layer1_outputs[312]) | (layer1_outputs[8239]);
    assign layer2_outputs[4248] = ~(layer1_outputs[3780]);
    assign layer2_outputs[4249] = (layer1_outputs[10726]) & (layer1_outputs[2068]);
    assign layer2_outputs[4250] = ~(layer1_outputs[407]) | (layer1_outputs[10864]);
    assign layer2_outputs[4251] = ~(layer1_outputs[5726]) | (layer1_outputs[4444]);
    assign layer2_outputs[4252] = (layer1_outputs[7980]) ^ (layer1_outputs[1238]);
    assign layer2_outputs[4253] = ~((layer1_outputs[3357]) & (layer1_outputs[12733]));
    assign layer2_outputs[4254] = ~((layer1_outputs[12706]) ^ (layer1_outputs[828]));
    assign layer2_outputs[4255] = ~(layer1_outputs[12456]);
    assign layer2_outputs[4256] = ~(layer1_outputs[8526]);
    assign layer2_outputs[4257] = (layer1_outputs[8643]) & ~(layer1_outputs[11195]);
    assign layer2_outputs[4258] = ~(layer1_outputs[6355]) | (layer1_outputs[6283]);
    assign layer2_outputs[4259] = (layer1_outputs[984]) & ~(layer1_outputs[7800]);
    assign layer2_outputs[4260] = ~((layer1_outputs[4083]) & (layer1_outputs[12713]));
    assign layer2_outputs[4261] = (layer1_outputs[3203]) | (layer1_outputs[9578]);
    assign layer2_outputs[4262] = ~(layer1_outputs[10030]);
    assign layer2_outputs[4263] = layer1_outputs[8473];
    assign layer2_outputs[4264] = ~((layer1_outputs[8377]) | (layer1_outputs[4081]));
    assign layer2_outputs[4265] = layer1_outputs[10701];
    assign layer2_outputs[4266] = ~((layer1_outputs[6215]) | (layer1_outputs[8573]));
    assign layer2_outputs[4267] = ~((layer1_outputs[6662]) & (layer1_outputs[868]));
    assign layer2_outputs[4268] = (layer1_outputs[7105]) & (layer1_outputs[10855]);
    assign layer2_outputs[4269] = ~((layer1_outputs[7342]) ^ (layer1_outputs[8651]));
    assign layer2_outputs[4270] = layer1_outputs[436];
    assign layer2_outputs[4271] = layer1_outputs[4538];
    assign layer2_outputs[4272] = layer1_outputs[6876];
    assign layer2_outputs[4273] = ~(layer1_outputs[8743]) | (layer1_outputs[4576]);
    assign layer2_outputs[4274] = ~((layer1_outputs[10533]) ^ (layer1_outputs[2793]));
    assign layer2_outputs[4275] = layer1_outputs[6954];
    assign layer2_outputs[4276] = ~((layer1_outputs[5912]) ^ (layer1_outputs[5177]));
    assign layer2_outputs[4277] = layer1_outputs[10];
    assign layer2_outputs[4278] = (layer1_outputs[12305]) & ~(layer1_outputs[2835]);
    assign layer2_outputs[4279] = layer1_outputs[6633];
    assign layer2_outputs[4280] = layer1_outputs[1585];
    assign layer2_outputs[4281] = ~(layer1_outputs[4416]);
    assign layer2_outputs[4282] = layer1_outputs[8365];
    assign layer2_outputs[4283] = ~(layer1_outputs[11051]);
    assign layer2_outputs[4284] = ~(layer1_outputs[1918]);
    assign layer2_outputs[4285] = (layer1_outputs[12612]) & ~(layer1_outputs[5987]);
    assign layer2_outputs[4286] = (layer1_outputs[4373]) ^ (layer1_outputs[1095]);
    assign layer2_outputs[4287] = ~(layer1_outputs[9589]);
    assign layer2_outputs[4288] = layer1_outputs[3750];
    assign layer2_outputs[4289] = layer1_outputs[2201];
    assign layer2_outputs[4290] = (layer1_outputs[8160]) | (layer1_outputs[7030]);
    assign layer2_outputs[4291] = (layer1_outputs[1356]) | (layer1_outputs[9030]);
    assign layer2_outputs[4292] = ~(layer1_outputs[6854]) | (layer1_outputs[6371]);
    assign layer2_outputs[4293] = ~((layer1_outputs[6236]) | (layer1_outputs[6794]));
    assign layer2_outputs[4294] = ~((layer1_outputs[8985]) | (layer1_outputs[6924]));
    assign layer2_outputs[4295] = layer1_outputs[6825];
    assign layer2_outputs[4296] = ~(layer1_outputs[12467]) | (layer1_outputs[12428]);
    assign layer2_outputs[4297] = ~(layer1_outputs[3368]) | (layer1_outputs[357]);
    assign layer2_outputs[4298] = (layer1_outputs[12698]) ^ (layer1_outputs[6455]);
    assign layer2_outputs[4299] = layer1_outputs[433];
    assign layer2_outputs[4300] = ~(layer1_outputs[10608]);
    assign layer2_outputs[4301] = ~(layer1_outputs[1343]);
    assign layer2_outputs[4302] = (layer1_outputs[4023]) & ~(layer1_outputs[7627]);
    assign layer2_outputs[4303] = ~(layer1_outputs[1784]) | (layer1_outputs[7346]);
    assign layer2_outputs[4304] = ~(layer1_outputs[9089]) | (layer1_outputs[9563]);
    assign layer2_outputs[4305] = layer1_outputs[825];
    assign layer2_outputs[4306] = layer1_outputs[1891];
    assign layer2_outputs[4307] = (layer1_outputs[6826]) & ~(layer1_outputs[9029]);
    assign layer2_outputs[4308] = (layer1_outputs[3771]) & (layer1_outputs[11217]);
    assign layer2_outputs[4309] = ~((layer1_outputs[8299]) & (layer1_outputs[9015]));
    assign layer2_outputs[4310] = ~((layer1_outputs[4714]) & (layer1_outputs[1391]));
    assign layer2_outputs[4311] = ~(layer1_outputs[440]);
    assign layer2_outputs[4312] = ~(layer1_outputs[3680]);
    assign layer2_outputs[4313] = ~(layer1_outputs[11537]);
    assign layer2_outputs[4314] = ~((layer1_outputs[388]) ^ (layer1_outputs[1882]));
    assign layer2_outputs[4315] = layer1_outputs[7750];
    assign layer2_outputs[4316] = ~(layer1_outputs[12504]);
    assign layer2_outputs[4317] = layer1_outputs[7527];
    assign layer2_outputs[4318] = layer1_outputs[11655];
    assign layer2_outputs[4319] = ~(layer1_outputs[10538]) | (layer1_outputs[2309]);
    assign layer2_outputs[4320] = ~((layer1_outputs[12552]) ^ (layer1_outputs[7198]));
    assign layer2_outputs[4321] = (layer1_outputs[3948]) ^ (layer1_outputs[4648]);
    assign layer2_outputs[4322] = ~((layer1_outputs[4188]) & (layer1_outputs[11846]));
    assign layer2_outputs[4323] = (layer1_outputs[5512]) & (layer1_outputs[10298]);
    assign layer2_outputs[4324] = ~((layer1_outputs[4873]) | (layer1_outputs[1894]));
    assign layer2_outputs[4325] = (layer1_outputs[6472]) | (layer1_outputs[3951]);
    assign layer2_outputs[4326] = ~(layer1_outputs[11000]);
    assign layer2_outputs[4327] = ~(layer1_outputs[12761]);
    assign layer2_outputs[4328] = ~(layer1_outputs[6796]);
    assign layer2_outputs[4329] = ~((layer1_outputs[9595]) & (layer1_outputs[6286]));
    assign layer2_outputs[4330] = ~(layer1_outputs[8366]);
    assign layer2_outputs[4331] = ~(layer1_outputs[10582]);
    assign layer2_outputs[4332] = (layer1_outputs[9635]) | (layer1_outputs[9841]);
    assign layer2_outputs[4333] = ~((layer1_outputs[570]) & (layer1_outputs[5750]));
    assign layer2_outputs[4334] = ~(layer1_outputs[5314]) | (layer1_outputs[7891]);
    assign layer2_outputs[4335] = (layer1_outputs[7481]) & (layer1_outputs[9864]);
    assign layer2_outputs[4336] = ~(layer1_outputs[63]);
    assign layer2_outputs[4337] = ~((layer1_outputs[8818]) | (layer1_outputs[10190]));
    assign layer2_outputs[4338] = ~(layer1_outputs[9612]);
    assign layer2_outputs[4339] = layer1_outputs[7831];
    assign layer2_outputs[4340] = (layer1_outputs[2196]) & ~(layer1_outputs[2799]);
    assign layer2_outputs[4341] = (layer1_outputs[1356]) & (layer1_outputs[12330]);
    assign layer2_outputs[4342] = (layer1_outputs[1952]) ^ (layer1_outputs[7189]);
    assign layer2_outputs[4343] = (layer1_outputs[1557]) | (layer1_outputs[1210]);
    assign layer2_outputs[4344] = (layer1_outputs[153]) & ~(layer1_outputs[11763]);
    assign layer2_outputs[4345] = (layer1_outputs[11164]) ^ (layer1_outputs[1466]);
    assign layer2_outputs[4346] = (layer1_outputs[4169]) & (layer1_outputs[5198]);
    assign layer2_outputs[4347] = ~(layer1_outputs[11472]);
    assign layer2_outputs[4348] = ~((layer1_outputs[12116]) & (layer1_outputs[4362]));
    assign layer2_outputs[4349] = layer1_outputs[7500];
    assign layer2_outputs[4350] = layer1_outputs[1782];
    assign layer2_outputs[4351] = (layer1_outputs[266]) ^ (layer1_outputs[12423]);
    assign layer2_outputs[4352] = ~(layer1_outputs[6747]);
    assign layer2_outputs[4353] = ~(layer1_outputs[5091]);
    assign layer2_outputs[4354] = ~(layer1_outputs[6397]) | (layer1_outputs[1723]);
    assign layer2_outputs[4355] = ~((layer1_outputs[10598]) ^ (layer1_outputs[10996]));
    assign layer2_outputs[4356] = ~((layer1_outputs[8787]) | (layer1_outputs[296]));
    assign layer2_outputs[4357] = layer1_outputs[11911];
    assign layer2_outputs[4358] = layer1_outputs[11864];
    assign layer2_outputs[4359] = ~(layer1_outputs[8562]);
    assign layer2_outputs[4360] = layer1_outputs[4519];
    assign layer2_outputs[4361] = ~((layer1_outputs[10391]) | (layer1_outputs[7591]));
    assign layer2_outputs[4362] = ~((layer1_outputs[12016]) ^ (layer1_outputs[11309]));
    assign layer2_outputs[4363] = ~((layer1_outputs[5391]) ^ (layer1_outputs[399]));
    assign layer2_outputs[4364] = ~(layer1_outputs[10694]) | (layer1_outputs[11887]);
    assign layer2_outputs[4365] = layer1_outputs[8069];
    assign layer2_outputs[4366] = ~(layer1_outputs[11894]);
    assign layer2_outputs[4367] = ~((layer1_outputs[10373]) | (layer1_outputs[3805]));
    assign layer2_outputs[4368] = (layer1_outputs[794]) ^ (layer1_outputs[8606]);
    assign layer2_outputs[4369] = (layer1_outputs[4393]) & ~(layer1_outputs[11184]);
    assign layer2_outputs[4370] = ~(layer1_outputs[9303]);
    assign layer2_outputs[4371] = (layer1_outputs[8869]) | (layer1_outputs[7118]);
    assign layer2_outputs[4372] = ~(layer1_outputs[2130]);
    assign layer2_outputs[4373] = ~((layer1_outputs[1527]) ^ (layer1_outputs[1302]));
    assign layer2_outputs[4374] = layer1_outputs[9732];
    assign layer2_outputs[4375] = ~(layer1_outputs[2796]) | (layer1_outputs[12079]);
    assign layer2_outputs[4376] = layer1_outputs[9283];
    assign layer2_outputs[4377] = (layer1_outputs[10599]) | (layer1_outputs[8471]);
    assign layer2_outputs[4378] = layer1_outputs[7782];
    assign layer2_outputs[4379] = ~(layer1_outputs[9970]);
    assign layer2_outputs[4380] = (layer1_outputs[886]) | (layer1_outputs[9327]);
    assign layer2_outputs[4381] = layer1_outputs[483];
    assign layer2_outputs[4382] = ~(layer1_outputs[5537]);
    assign layer2_outputs[4383] = layer1_outputs[2355];
    assign layer2_outputs[4384] = (layer1_outputs[11683]) & (layer1_outputs[11128]);
    assign layer2_outputs[4385] = layer1_outputs[8198];
    assign layer2_outputs[4386] = ~(layer1_outputs[3830]) | (layer1_outputs[1563]);
    assign layer2_outputs[4387] = (layer1_outputs[6066]) | (layer1_outputs[8280]);
    assign layer2_outputs[4388] = ~(layer1_outputs[10204]);
    assign layer2_outputs[4389] = layer1_outputs[7674];
    assign layer2_outputs[4390] = ~(layer1_outputs[1134]);
    assign layer2_outputs[4391] = layer1_outputs[539];
    assign layer2_outputs[4392] = (layer1_outputs[926]) & ~(layer1_outputs[7067]);
    assign layer2_outputs[4393] = ~(layer1_outputs[3257]) | (layer1_outputs[7024]);
    assign layer2_outputs[4394] = layer1_outputs[6106];
    assign layer2_outputs[4395] = ~((layer1_outputs[12472]) | (layer1_outputs[4555]));
    assign layer2_outputs[4396] = (layer1_outputs[576]) & ~(layer1_outputs[11306]);
    assign layer2_outputs[4397] = ~(layer1_outputs[9865]);
    assign layer2_outputs[4398] = ~(layer1_outputs[325]);
    assign layer2_outputs[4399] = layer1_outputs[7389];
    assign layer2_outputs[4400] = ~(layer1_outputs[6766]);
    assign layer2_outputs[4401] = layer1_outputs[5213];
    assign layer2_outputs[4402] = ~(layer1_outputs[1916]) | (layer1_outputs[5326]);
    assign layer2_outputs[4403] = ~(layer1_outputs[10987]);
    assign layer2_outputs[4404] = 1'b1;
    assign layer2_outputs[4405] = layer1_outputs[6092];
    assign layer2_outputs[4406] = ~(layer1_outputs[8914]) | (layer1_outputs[10072]);
    assign layer2_outputs[4407] = ~(layer1_outputs[9781]);
    assign layer2_outputs[4408] = (layer1_outputs[12719]) & ~(layer1_outputs[1642]);
    assign layer2_outputs[4409] = (layer1_outputs[12236]) ^ (layer1_outputs[6128]);
    assign layer2_outputs[4410] = ~(layer1_outputs[1263]);
    assign layer2_outputs[4411] = layer1_outputs[6095];
    assign layer2_outputs[4412] = layer1_outputs[6136];
    assign layer2_outputs[4413] = 1'b1;
    assign layer2_outputs[4414] = 1'b1;
    assign layer2_outputs[4415] = ~(layer1_outputs[5923]) | (layer1_outputs[12771]);
    assign layer2_outputs[4416] = (layer1_outputs[3435]) & ~(layer1_outputs[7117]);
    assign layer2_outputs[4417] = layer1_outputs[10380];
    assign layer2_outputs[4418] = layer1_outputs[5281];
    assign layer2_outputs[4419] = (layer1_outputs[2150]) ^ (layer1_outputs[216]);
    assign layer2_outputs[4420] = layer1_outputs[2872];
    assign layer2_outputs[4421] = ~(layer1_outputs[1429]);
    assign layer2_outputs[4422] = ~(layer1_outputs[2676]);
    assign layer2_outputs[4423] = (layer1_outputs[10911]) ^ (layer1_outputs[3744]);
    assign layer2_outputs[4424] = (layer1_outputs[1441]) & ~(layer1_outputs[5222]);
    assign layer2_outputs[4425] = ~(layer1_outputs[11329]);
    assign layer2_outputs[4426] = ~(layer1_outputs[10640]) | (layer1_outputs[55]);
    assign layer2_outputs[4427] = layer1_outputs[5213];
    assign layer2_outputs[4428] = layer1_outputs[547];
    assign layer2_outputs[4429] = ~(layer1_outputs[3809]);
    assign layer2_outputs[4430] = (layer1_outputs[8866]) & (layer1_outputs[4346]);
    assign layer2_outputs[4431] = ~((layer1_outputs[9864]) ^ (layer1_outputs[12072]));
    assign layer2_outputs[4432] = layer1_outputs[2288];
    assign layer2_outputs[4433] = (layer1_outputs[4469]) & ~(layer1_outputs[1107]);
    assign layer2_outputs[4434] = ~((layer1_outputs[5533]) ^ (layer1_outputs[12153]));
    assign layer2_outputs[4435] = (layer1_outputs[10838]) ^ (layer1_outputs[690]);
    assign layer2_outputs[4436] = layer1_outputs[2608];
    assign layer2_outputs[4437] = (layer1_outputs[10393]) & ~(layer1_outputs[12436]);
    assign layer2_outputs[4438] = (layer1_outputs[1499]) & (layer1_outputs[3756]);
    assign layer2_outputs[4439] = layer1_outputs[516];
    assign layer2_outputs[4440] = ~(layer1_outputs[12266]);
    assign layer2_outputs[4441] = layer1_outputs[6511];
    assign layer2_outputs[4442] = ~(layer1_outputs[5818]) | (layer1_outputs[4034]);
    assign layer2_outputs[4443] = ~((layer1_outputs[2905]) ^ (layer1_outputs[2580]));
    assign layer2_outputs[4444] = ~(layer1_outputs[6390]);
    assign layer2_outputs[4445] = (layer1_outputs[1969]) | (layer1_outputs[6559]);
    assign layer2_outputs[4446] = layer1_outputs[9361];
    assign layer2_outputs[4447] = 1'b0;
    assign layer2_outputs[4448] = (layer1_outputs[1589]) ^ (layer1_outputs[5131]);
    assign layer2_outputs[4449] = layer1_outputs[1621];
    assign layer2_outputs[4450] = ~(layer1_outputs[2908]) | (layer1_outputs[10244]);
    assign layer2_outputs[4451] = ~((layer1_outputs[6979]) & (layer1_outputs[8411]));
    assign layer2_outputs[4452] = (layer1_outputs[10024]) ^ (layer1_outputs[11628]);
    assign layer2_outputs[4453] = layer1_outputs[8373];
    assign layer2_outputs[4454] = (layer1_outputs[12288]) & ~(layer1_outputs[8608]);
    assign layer2_outputs[4455] = (layer1_outputs[1691]) ^ (layer1_outputs[9862]);
    assign layer2_outputs[4456] = ~(layer1_outputs[8263]);
    assign layer2_outputs[4457] = layer1_outputs[552];
    assign layer2_outputs[4458] = layer1_outputs[631];
    assign layer2_outputs[4459] = ~(layer1_outputs[9340]);
    assign layer2_outputs[4460] = layer1_outputs[5527];
    assign layer2_outputs[4461] = layer1_outputs[3324];
    assign layer2_outputs[4462] = ~((layer1_outputs[9446]) & (layer1_outputs[3397]));
    assign layer2_outputs[4463] = (layer1_outputs[8386]) & ~(layer1_outputs[6326]);
    assign layer2_outputs[4464] = ~((layer1_outputs[2831]) ^ (layer1_outputs[2947]));
    assign layer2_outputs[4465] = ~((layer1_outputs[1143]) ^ (layer1_outputs[2564]));
    assign layer2_outputs[4466] = (layer1_outputs[6576]) ^ (layer1_outputs[9444]);
    assign layer2_outputs[4467] = layer1_outputs[10068];
    assign layer2_outputs[4468] = ~(layer1_outputs[7949]);
    assign layer2_outputs[4469] = ~(layer1_outputs[5383]);
    assign layer2_outputs[4470] = ~(layer1_outputs[11161]);
    assign layer2_outputs[4471] = (layer1_outputs[2879]) ^ (layer1_outputs[308]);
    assign layer2_outputs[4472] = layer1_outputs[7931];
    assign layer2_outputs[4473] = layer1_outputs[386];
    assign layer2_outputs[4474] = (layer1_outputs[12277]) ^ (layer1_outputs[8206]);
    assign layer2_outputs[4475] = (layer1_outputs[2276]) & ~(layer1_outputs[2024]);
    assign layer2_outputs[4476] = layer1_outputs[6602];
    assign layer2_outputs[4477] = layer1_outputs[2219];
    assign layer2_outputs[4478] = ~((layer1_outputs[8902]) ^ (layer1_outputs[12709]));
    assign layer2_outputs[4479] = layer1_outputs[8712];
    assign layer2_outputs[4480] = ~(layer1_outputs[5371]);
    assign layer2_outputs[4481] = ~((layer1_outputs[2359]) ^ (layer1_outputs[565]));
    assign layer2_outputs[4482] = ~(layer1_outputs[12640]) | (layer1_outputs[9734]);
    assign layer2_outputs[4483] = (layer1_outputs[11110]) & ~(layer1_outputs[7061]);
    assign layer2_outputs[4484] = ~((layer1_outputs[8996]) ^ (layer1_outputs[4522]));
    assign layer2_outputs[4485] = ~(layer1_outputs[2661]) | (layer1_outputs[1580]);
    assign layer2_outputs[4486] = ~(layer1_outputs[8136]);
    assign layer2_outputs[4487] = ~(layer1_outputs[4032]);
    assign layer2_outputs[4488] = ~((layer1_outputs[9148]) ^ (layer1_outputs[10788]));
    assign layer2_outputs[4489] = (layer1_outputs[567]) & ~(layer1_outputs[3968]);
    assign layer2_outputs[4490] = ~(layer1_outputs[4917]);
    assign layer2_outputs[4491] = (layer1_outputs[919]) | (layer1_outputs[7565]);
    assign layer2_outputs[4492] = ~((layer1_outputs[4329]) & (layer1_outputs[12004]));
    assign layer2_outputs[4493] = (layer1_outputs[3860]) | (layer1_outputs[10255]);
    assign layer2_outputs[4494] = ~((layer1_outputs[4257]) | (layer1_outputs[6]));
    assign layer2_outputs[4495] = layer1_outputs[9277];
    assign layer2_outputs[4496] = ~(layer1_outputs[5382]);
    assign layer2_outputs[4497] = ~(layer1_outputs[9472]) | (layer1_outputs[4743]);
    assign layer2_outputs[4498] = ~((layer1_outputs[6404]) ^ (layer1_outputs[12781]));
    assign layer2_outputs[4499] = ~(layer1_outputs[12060]);
    assign layer2_outputs[4500] = ~((layer1_outputs[197]) | (layer1_outputs[2535]));
    assign layer2_outputs[4501] = (layer1_outputs[8026]) | (layer1_outputs[1012]);
    assign layer2_outputs[4502] = (layer1_outputs[4104]) | (layer1_outputs[10672]);
    assign layer2_outputs[4503] = (layer1_outputs[7466]) & ~(layer1_outputs[2506]);
    assign layer2_outputs[4504] = ~((layer1_outputs[7139]) ^ (layer1_outputs[6724]));
    assign layer2_outputs[4505] = layer1_outputs[3462];
    assign layer2_outputs[4506] = (layer1_outputs[3232]) & (layer1_outputs[6864]);
    assign layer2_outputs[4507] = (layer1_outputs[502]) ^ (layer1_outputs[1777]);
    assign layer2_outputs[4508] = ~(layer1_outputs[6498]);
    assign layer2_outputs[4509] = ~(layer1_outputs[4293]);
    assign layer2_outputs[4510] = layer1_outputs[4199];
    assign layer2_outputs[4511] = layer1_outputs[2088];
    assign layer2_outputs[4512] = ~(layer1_outputs[10211]) | (layer1_outputs[904]);
    assign layer2_outputs[4513] = layer1_outputs[5748];
    assign layer2_outputs[4514] = layer1_outputs[9210];
    assign layer2_outputs[4515] = ~(layer1_outputs[10723]);
    assign layer2_outputs[4516] = ~(layer1_outputs[8880]);
    assign layer2_outputs[4517] = layer1_outputs[3552];
    assign layer2_outputs[4518] = ~(layer1_outputs[9862]) | (layer1_outputs[2511]);
    assign layer2_outputs[4519] = ~((layer1_outputs[7437]) | (layer1_outputs[8084]));
    assign layer2_outputs[4520] = layer1_outputs[7755];
    assign layer2_outputs[4521] = (layer1_outputs[1279]) & (layer1_outputs[6189]);
    assign layer2_outputs[4522] = ~((layer1_outputs[4381]) ^ (layer1_outputs[1716]));
    assign layer2_outputs[4523] = layer1_outputs[8589];
    assign layer2_outputs[4524] = (layer1_outputs[7644]) & ~(layer1_outputs[2620]);
    assign layer2_outputs[4525] = layer1_outputs[12487];
    assign layer2_outputs[4526] = (layer1_outputs[5590]) ^ (layer1_outputs[6646]);
    assign layer2_outputs[4527] = ~(layer1_outputs[11525]);
    assign layer2_outputs[4528] = ~((layer1_outputs[8304]) | (layer1_outputs[1634]));
    assign layer2_outputs[4529] = ~(layer1_outputs[513]);
    assign layer2_outputs[4530] = (layer1_outputs[3418]) & (layer1_outputs[8331]);
    assign layer2_outputs[4531] = (layer1_outputs[12599]) | (layer1_outputs[4302]);
    assign layer2_outputs[4532] = (layer1_outputs[1186]) | (layer1_outputs[4372]);
    assign layer2_outputs[4533] = ~(layer1_outputs[7079]);
    assign layer2_outputs[4534] = ~(layer1_outputs[2479]);
    assign layer2_outputs[4535] = ~(layer1_outputs[7841]);
    assign layer2_outputs[4536] = layer1_outputs[1674];
    assign layer2_outputs[4537] = layer1_outputs[2606];
    assign layer2_outputs[4538] = layer1_outputs[9218];
    assign layer2_outputs[4539] = ~((layer1_outputs[5730]) ^ (layer1_outputs[2142]));
    assign layer2_outputs[4540] = (layer1_outputs[3289]) & ~(layer1_outputs[3748]);
    assign layer2_outputs[4541] = ~((layer1_outputs[4347]) ^ (layer1_outputs[9534]));
    assign layer2_outputs[4542] = (layer1_outputs[10685]) ^ (layer1_outputs[12344]);
    assign layer2_outputs[4543] = ~((layer1_outputs[4094]) ^ (layer1_outputs[3206]));
    assign layer2_outputs[4544] = ~((layer1_outputs[6499]) ^ (layer1_outputs[3071]));
    assign layer2_outputs[4545] = ~((layer1_outputs[10165]) | (layer1_outputs[3806]));
    assign layer2_outputs[4546] = layer1_outputs[4156];
    assign layer2_outputs[4547] = ~(layer1_outputs[11847]);
    assign layer2_outputs[4548] = ~(layer1_outputs[12074]);
    assign layer2_outputs[4549] = (layer1_outputs[1436]) ^ (layer1_outputs[8134]);
    assign layer2_outputs[4550] = ~(layer1_outputs[3220]) | (layer1_outputs[12435]);
    assign layer2_outputs[4551] = ~(layer1_outputs[2635]) | (layer1_outputs[2631]);
    assign layer2_outputs[4552] = ~(layer1_outputs[11381]);
    assign layer2_outputs[4553] = layer1_outputs[1622];
    assign layer2_outputs[4554] = (layer1_outputs[7214]) & (layer1_outputs[2549]);
    assign layer2_outputs[4555] = layer1_outputs[10157];
    assign layer2_outputs[4556] = ~(layer1_outputs[12708]);
    assign layer2_outputs[4557] = ~(layer1_outputs[3427]) | (layer1_outputs[11214]);
    assign layer2_outputs[4558] = ~(layer1_outputs[3384]) | (layer1_outputs[3262]);
    assign layer2_outputs[4559] = layer1_outputs[316];
    assign layer2_outputs[4560] = ~(layer1_outputs[2514]);
    assign layer2_outputs[4561] = (layer1_outputs[9573]) | (layer1_outputs[422]);
    assign layer2_outputs[4562] = (layer1_outputs[968]) & ~(layer1_outputs[1293]);
    assign layer2_outputs[4563] = (layer1_outputs[1846]) & ~(layer1_outputs[1728]);
    assign layer2_outputs[4564] = layer1_outputs[1939];
    assign layer2_outputs[4565] = ~(layer1_outputs[2060]);
    assign layer2_outputs[4566] = ~((layer1_outputs[10554]) & (layer1_outputs[750]));
    assign layer2_outputs[4567] = layer1_outputs[8293];
    assign layer2_outputs[4568] = layer1_outputs[2194];
    assign layer2_outputs[4569] = ~(layer1_outputs[4183]);
    assign layer2_outputs[4570] = ~((layer1_outputs[8135]) | (layer1_outputs[6764]));
    assign layer2_outputs[4571] = (layer1_outputs[11704]) & ~(layer1_outputs[5319]);
    assign layer2_outputs[4572] = ~(layer1_outputs[6815]);
    assign layer2_outputs[4573] = layer1_outputs[5109];
    assign layer2_outputs[4574] = ~(layer1_outputs[10498]);
    assign layer2_outputs[4575] = layer1_outputs[4008];
    assign layer2_outputs[4576] = ~((layer1_outputs[10173]) ^ (layer1_outputs[8786]));
    assign layer2_outputs[4577] = ~(layer1_outputs[7690]);
    assign layer2_outputs[4578] = ~(layer1_outputs[5825]) | (layer1_outputs[5777]);
    assign layer2_outputs[4579] = (layer1_outputs[3478]) ^ (layer1_outputs[4888]);
    assign layer2_outputs[4580] = layer1_outputs[10392];
    assign layer2_outputs[4581] = (layer1_outputs[5750]) ^ (layer1_outputs[1479]);
    assign layer2_outputs[4582] = ~(layer1_outputs[6706]);
    assign layer2_outputs[4583] = ~(layer1_outputs[10632]);
    assign layer2_outputs[4584] = layer1_outputs[7089];
    assign layer2_outputs[4585] = layer1_outputs[11615];
    assign layer2_outputs[4586] = ~(layer1_outputs[5302]);
    assign layer2_outputs[4587] = ~((layer1_outputs[6440]) ^ (layer1_outputs[10877]));
    assign layer2_outputs[4588] = (layer1_outputs[9668]) & ~(layer1_outputs[12304]);
    assign layer2_outputs[4589] = layer1_outputs[3407];
    assign layer2_outputs[4590] = ~((layer1_outputs[8837]) ^ (layer1_outputs[6470]));
    assign layer2_outputs[4591] = ~((layer1_outputs[5414]) ^ (layer1_outputs[12013]));
    assign layer2_outputs[4592] = ~(layer1_outputs[10986]);
    assign layer2_outputs[4593] = ~(layer1_outputs[4633]);
    assign layer2_outputs[4594] = ~(layer1_outputs[4266]);
    assign layer2_outputs[4595] = layer1_outputs[5053];
    assign layer2_outputs[4596] = ~(layer1_outputs[11266]) | (layer1_outputs[11315]);
    assign layer2_outputs[4597] = ~(layer1_outputs[7943]);
    assign layer2_outputs[4598] = layer1_outputs[7619];
    assign layer2_outputs[4599] = (layer1_outputs[8030]) & (layer1_outputs[11232]);
    assign layer2_outputs[4600] = ~(layer1_outputs[12105]);
    assign layer2_outputs[4601] = (layer1_outputs[5104]) & ~(layer1_outputs[791]);
    assign layer2_outputs[4602] = ~(layer1_outputs[1108]);
    assign layer2_outputs[4603] = ~(layer1_outputs[5521]);
    assign layer2_outputs[4604] = ~(layer1_outputs[2829]);
    assign layer2_outputs[4605] = (layer1_outputs[3227]) ^ (layer1_outputs[11023]);
    assign layer2_outputs[4606] = layer1_outputs[7926];
    assign layer2_outputs[4607] = (layer1_outputs[6758]) & (layer1_outputs[6306]);
    assign layer2_outputs[4608] = ~(layer1_outputs[276]);
    assign layer2_outputs[4609] = (layer1_outputs[4269]) & ~(layer1_outputs[2792]);
    assign layer2_outputs[4610] = (layer1_outputs[12775]) & ~(layer1_outputs[5234]);
    assign layer2_outputs[4611] = layer1_outputs[10702];
    assign layer2_outputs[4612] = ~(layer1_outputs[11630]);
    assign layer2_outputs[4613] = ~(layer1_outputs[5172]);
    assign layer2_outputs[4614] = layer1_outputs[127];
    assign layer2_outputs[4615] = (layer1_outputs[8932]) & ~(layer1_outputs[4446]);
    assign layer2_outputs[4616] = (layer1_outputs[10010]) & ~(layer1_outputs[335]);
    assign layer2_outputs[4617] = ~(layer1_outputs[1934]);
    assign layer2_outputs[4618] = (layer1_outputs[5239]) & ~(layer1_outputs[8248]);
    assign layer2_outputs[4619] = layer1_outputs[3075];
    assign layer2_outputs[4620] = ~((layer1_outputs[6175]) ^ (layer1_outputs[7473]));
    assign layer2_outputs[4621] = layer1_outputs[7339];
    assign layer2_outputs[4622] = ~((layer1_outputs[10819]) | (layer1_outputs[8984]));
    assign layer2_outputs[4623] = layer1_outputs[7313];
    assign layer2_outputs[4624] = layer1_outputs[2907];
    assign layer2_outputs[4625] = ~(layer1_outputs[409]) | (layer1_outputs[11892]);
    assign layer2_outputs[4626] = ~((layer1_outputs[1689]) ^ (layer1_outputs[222]));
    assign layer2_outputs[4627] = ~((layer1_outputs[8895]) & (layer1_outputs[2084]));
    assign layer2_outputs[4628] = layer1_outputs[7166];
    assign layer2_outputs[4629] = ~(layer1_outputs[5800]);
    assign layer2_outputs[4630] = ~(layer1_outputs[3498]);
    assign layer2_outputs[4631] = layer1_outputs[9641];
    assign layer2_outputs[4632] = ~(layer1_outputs[5791]);
    assign layer2_outputs[4633] = layer1_outputs[9326];
    assign layer2_outputs[4634] = layer1_outputs[8821];
    assign layer2_outputs[4635] = ~(layer1_outputs[3495]);
    assign layer2_outputs[4636] = (layer1_outputs[2422]) & ~(layer1_outputs[4081]);
    assign layer2_outputs[4637] = layer1_outputs[3124];
    assign layer2_outputs[4638] = layer1_outputs[6318];
    assign layer2_outputs[4639] = ~(layer1_outputs[6911]);
    assign layer2_outputs[4640] = ~((layer1_outputs[10319]) | (layer1_outputs[6552]));
    assign layer2_outputs[4641] = ~(layer1_outputs[353]);
    assign layer2_outputs[4642] = (layer1_outputs[10330]) & ~(layer1_outputs[3970]);
    assign layer2_outputs[4643] = ~(layer1_outputs[7196]);
    assign layer2_outputs[4644] = ~((layer1_outputs[4127]) & (layer1_outputs[1040]));
    assign layer2_outputs[4645] = (layer1_outputs[3292]) | (layer1_outputs[9452]);
    assign layer2_outputs[4646] = (layer1_outputs[549]) | (layer1_outputs[2293]);
    assign layer2_outputs[4647] = ~(layer1_outputs[264]);
    assign layer2_outputs[4648] = (layer1_outputs[9334]) | (layer1_outputs[4606]);
    assign layer2_outputs[4649] = layer1_outputs[9146];
    assign layer2_outputs[4650] = ~(layer1_outputs[6635]);
    assign layer2_outputs[4651] = layer1_outputs[11530];
    assign layer2_outputs[4652] = (layer1_outputs[12098]) ^ (layer1_outputs[12430]);
    assign layer2_outputs[4653] = (layer1_outputs[659]) & ~(layer1_outputs[9204]);
    assign layer2_outputs[4654] = layer1_outputs[243];
    assign layer2_outputs[4655] = ~(layer1_outputs[5342]) | (layer1_outputs[889]);
    assign layer2_outputs[4656] = (layer1_outputs[5028]) | (layer1_outputs[1798]);
    assign layer2_outputs[4657] = layer1_outputs[9081];
    assign layer2_outputs[4658] = (layer1_outputs[5956]) ^ (layer1_outputs[3651]);
    assign layer2_outputs[4659] = ~(layer1_outputs[11690]) | (layer1_outputs[9773]);
    assign layer2_outputs[4660] = ~(layer1_outputs[8703]);
    assign layer2_outputs[4661] = ~(layer1_outputs[4982]);
    assign layer2_outputs[4662] = layer1_outputs[9564];
    assign layer2_outputs[4663] = ~((layer1_outputs[2353]) | (layer1_outputs[5179]));
    assign layer2_outputs[4664] = layer1_outputs[131];
    assign layer2_outputs[4665] = ~(layer1_outputs[10704]) | (layer1_outputs[26]);
    assign layer2_outputs[4666] = ~(layer1_outputs[2650]);
    assign layer2_outputs[4667] = layer1_outputs[357];
    assign layer2_outputs[4668] = ~(layer1_outputs[4709]);
    assign layer2_outputs[4669] = ~(layer1_outputs[2526]);
    assign layer2_outputs[4670] = (layer1_outputs[9289]) & ~(layer1_outputs[10825]);
    assign layer2_outputs[4671] = (layer1_outputs[12484]) & ~(layer1_outputs[12029]);
    assign layer2_outputs[4672] = layer1_outputs[7893];
    assign layer2_outputs[4673] = ~(layer1_outputs[9827]);
    assign layer2_outputs[4674] = 1'b0;
    assign layer2_outputs[4675] = layer1_outputs[6506];
    assign layer2_outputs[4676] = (layer1_outputs[11603]) | (layer1_outputs[4141]);
    assign layer2_outputs[4677] = (layer1_outputs[7888]) & ~(layer1_outputs[4130]);
    assign layer2_outputs[4678] = ~(layer1_outputs[8776]);
    assign layer2_outputs[4679] = (layer1_outputs[9025]) ^ (layer1_outputs[1746]);
    assign layer2_outputs[4680] = ~(layer1_outputs[12182]);
    assign layer2_outputs[4681] = ~((layer1_outputs[10985]) | (layer1_outputs[9600]));
    assign layer2_outputs[4682] = (layer1_outputs[4218]) & ~(layer1_outputs[9765]);
    assign layer2_outputs[4683] = ~((layer1_outputs[3180]) ^ (layer1_outputs[12015]));
    assign layer2_outputs[4684] = ~(layer1_outputs[5134]);
    assign layer2_outputs[4685] = layer1_outputs[12794];
    assign layer2_outputs[4686] = layer1_outputs[854];
    assign layer2_outputs[4687] = (layer1_outputs[12490]) & (layer1_outputs[1147]);
    assign layer2_outputs[4688] = (layer1_outputs[7076]) ^ (layer1_outputs[3400]);
    assign layer2_outputs[4689] = (layer1_outputs[10448]) & (layer1_outputs[10827]);
    assign layer2_outputs[4690] = layer1_outputs[4374];
    assign layer2_outputs[4691] = ~(layer1_outputs[7766]);
    assign layer2_outputs[4692] = ~(layer1_outputs[602]);
    assign layer2_outputs[4693] = (layer1_outputs[1812]) & ~(layer1_outputs[1131]);
    assign layer2_outputs[4694] = layer1_outputs[7432];
    assign layer2_outputs[4695] = ~(layer1_outputs[2286]);
    assign layer2_outputs[4696] = ~((layer1_outputs[2812]) | (layer1_outputs[8325]));
    assign layer2_outputs[4697] = ~(layer1_outputs[3740]);
    assign layer2_outputs[4698] = ~(layer1_outputs[9317]);
    assign layer2_outputs[4699] = ~(layer1_outputs[12243]);
    assign layer2_outputs[4700] = (layer1_outputs[4122]) & (layer1_outputs[10565]);
    assign layer2_outputs[4701] = ~(layer1_outputs[11072]);
    assign layer2_outputs[4702] = ~(layer1_outputs[6987]);
    assign layer2_outputs[4703] = ~(layer1_outputs[10793]);
    assign layer2_outputs[4704] = ~((layer1_outputs[9132]) | (layer1_outputs[4074]));
    assign layer2_outputs[4705] = layer1_outputs[4745];
    assign layer2_outputs[4706] = ~(layer1_outputs[10017]);
    assign layer2_outputs[4707] = layer1_outputs[7589];
    assign layer2_outputs[4708] = ~((layer1_outputs[2417]) & (layer1_outputs[1678]));
    assign layer2_outputs[4709] = ~((layer1_outputs[2582]) ^ (layer1_outputs[9664]));
    assign layer2_outputs[4710] = layer1_outputs[2132];
    assign layer2_outputs[4711] = (layer1_outputs[594]) & (layer1_outputs[291]);
    assign layer2_outputs[4712] = (layer1_outputs[7152]) ^ (layer1_outputs[6640]);
    assign layer2_outputs[4713] = 1'b1;
    assign layer2_outputs[4714] = ~((layer1_outputs[3633]) ^ (layer1_outputs[3060]));
    assign layer2_outputs[4715] = ~((layer1_outputs[4815]) ^ (layer1_outputs[9050]));
    assign layer2_outputs[4716] = ~(layer1_outputs[4739]);
    assign layer2_outputs[4717] = ~(layer1_outputs[1543]);
    assign layer2_outputs[4718] = (layer1_outputs[12273]) & ~(layer1_outputs[7194]);
    assign layer2_outputs[4719] = ~(layer1_outputs[2427]);
    assign layer2_outputs[4720] = ~(layer1_outputs[12235]);
    assign layer2_outputs[4721] = (layer1_outputs[8778]) & ~(layer1_outputs[2300]);
    assign layer2_outputs[4722] = ~(layer1_outputs[10104]) | (layer1_outputs[10372]);
    assign layer2_outputs[4723] = layer1_outputs[8913];
    assign layer2_outputs[4724] = ~(layer1_outputs[7683]) | (layer1_outputs[8959]);
    assign layer2_outputs[4725] = ~((layer1_outputs[3945]) ^ (layer1_outputs[11656]));
    assign layer2_outputs[4726] = (layer1_outputs[12148]) & ~(layer1_outputs[3962]);
    assign layer2_outputs[4727] = ~(layer1_outputs[7841]) | (layer1_outputs[7444]);
    assign layer2_outputs[4728] = ~(layer1_outputs[6645]);
    assign layer2_outputs[4729] = ~(layer1_outputs[10650]);
    assign layer2_outputs[4730] = (layer1_outputs[9101]) ^ (layer1_outputs[3509]);
    assign layer2_outputs[4731] = layer1_outputs[5210];
    assign layer2_outputs[4732] = (layer1_outputs[12516]) & ~(layer1_outputs[7860]);
    assign layer2_outputs[4733] = (layer1_outputs[1338]) & (layer1_outputs[10086]);
    assign layer2_outputs[4734] = ~((layer1_outputs[3319]) ^ (layer1_outputs[11991]));
    assign layer2_outputs[4735] = ~((layer1_outputs[6684]) | (layer1_outputs[593]));
    assign layer2_outputs[4736] = ~((layer1_outputs[9721]) ^ (layer1_outputs[11386]));
    assign layer2_outputs[4737] = ~((layer1_outputs[10905]) ^ (layer1_outputs[3231]));
    assign layer2_outputs[4738] = ~(layer1_outputs[9987]);
    assign layer2_outputs[4739] = ~(layer1_outputs[11246]) | (layer1_outputs[11928]);
    assign layer2_outputs[4740] = layer1_outputs[4730];
    assign layer2_outputs[4741] = (layer1_outputs[4666]) & ~(layer1_outputs[3245]);
    assign layer2_outputs[4742] = ~(layer1_outputs[12111]);
    assign layer2_outputs[4743] = layer1_outputs[8502];
    assign layer2_outputs[4744] = ~(layer1_outputs[8100]) | (layer1_outputs[8165]);
    assign layer2_outputs[4745] = layer1_outputs[3842];
    assign layer2_outputs[4746] = (layer1_outputs[8142]) ^ (layer1_outputs[1461]);
    assign layer2_outputs[4747] = layer1_outputs[4299];
    assign layer2_outputs[4748] = ~(layer1_outputs[7931]);
    assign layer2_outputs[4749] = (layer1_outputs[5806]) | (layer1_outputs[11028]);
    assign layer2_outputs[4750] = (layer1_outputs[12559]) | (layer1_outputs[4143]);
    assign layer2_outputs[4751] = (layer1_outputs[5011]) & (layer1_outputs[5697]);
    assign layer2_outputs[4752] = ~(layer1_outputs[5789]);
    assign layer2_outputs[4753] = ~(layer1_outputs[589]);
    assign layer2_outputs[4754] = ~(layer1_outputs[9892]);
    assign layer2_outputs[4755] = (layer1_outputs[2782]) & ~(layer1_outputs[9825]);
    assign layer2_outputs[4756] = layer1_outputs[9752];
    assign layer2_outputs[4757] = ~(layer1_outputs[8553]) | (layer1_outputs[12037]);
    assign layer2_outputs[4758] = layer1_outputs[5710];
    assign layer2_outputs[4759] = ~((layer1_outputs[329]) ^ (layer1_outputs[8068]));
    assign layer2_outputs[4760] = layer1_outputs[953];
    assign layer2_outputs[4761] = ~(layer1_outputs[1967]) | (layer1_outputs[10939]);
    assign layer2_outputs[4762] = layer1_outputs[7829];
    assign layer2_outputs[4763] = ~((layer1_outputs[11206]) | (layer1_outputs[8210]));
    assign layer2_outputs[4764] = layer1_outputs[2684];
    assign layer2_outputs[4765] = layer1_outputs[1294];
    assign layer2_outputs[4766] = layer1_outputs[8086];
    assign layer2_outputs[4767] = (layer1_outputs[6641]) | (layer1_outputs[1894]);
    assign layer2_outputs[4768] = ~(layer1_outputs[8837]);
    assign layer2_outputs[4769] = (layer1_outputs[312]) & (layer1_outputs[4520]);
    assign layer2_outputs[4770] = layer1_outputs[10238];
    assign layer2_outputs[4771] = ~(layer1_outputs[11558]);
    assign layer2_outputs[4772] = ~(layer1_outputs[5688]);
    assign layer2_outputs[4773] = (layer1_outputs[3268]) ^ (layer1_outputs[6115]);
    assign layer2_outputs[4774] = (layer1_outputs[3748]) | (layer1_outputs[6626]);
    assign layer2_outputs[4775] = layer1_outputs[3103];
    assign layer2_outputs[4776] = ~((layer1_outputs[11210]) ^ (layer1_outputs[7542]));
    assign layer2_outputs[4777] = layer1_outputs[6021];
    assign layer2_outputs[4778] = ~(layer1_outputs[2602]);
    assign layer2_outputs[4779] = ~(layer1_outputs[3449]) | (layer1_outputs[1083]);
    assign layer2_outputs[4780] = ~(layer1_outputs[8817]);
    assign layer2_outputs[4781] = ~(layer1_outputs[10377]);
    assign layer2_outputs[4782] = ~(layer1_outputs[10423]);
    assign layer2_outputs[4783] = (layer1_outputs[12740]) & ~(layer1_outputs[2949]);
    assign layer2_outputs[4784] = ~(layer1_outputs[3893]);
    assign layer2_outputs[4785] = ~(layer1_outputs[8119]);
    assign layer2_outputs[4786] = ~(layer1_outputs[1865]);
    assign layer2_outputs[4787] = (layer1_outputs[6261]) & (layer1_outputs[6612]);
    assign layer2_outputs[4788] = layer1_outputs[10466];
    assign layer2_outputs[4789] = layer1_outputs[6100];
    assign layer2_outputs[4790] = layer1_outputs[11126];
    assign layer2_outputs[4791] = ~(layer1_outputs[1359]);
    assign layer2_outputs[4792] = ~((layer1_outputs[3834]) ^ (layer1_outputs[12135]));
    assign layer2_outputs[4793] = (layer1_outputs[648]) & (layer1_outputs[5368]);
    assign layer2_outputs[4794] = layer1_outputs[4490];
    assign layer2_outputs[4795] = (layer1_outputs[2590]) ^ (layer1_outputs[9289]);
    assign layer2_outputs[4796] = ~((layer1_outputs[175]) ^ (layer1_outputs[3030]));
    assign layer2_outputs[4797] = ~((layer1_outputs[9965]) | (layer1_outputs[163]));
    assign layer2_outputs[4798] = layer1_outputs[8699];
    assign layer2_outputs[4799] = ~(layer1_outputs[11549]);
    assign layer2_outputs[4800] = (layer1_outputs[6090]) & ~(layer1_outputs[7054]);
    assign layer2_outputs[4801] = ~((layer1_outputs[3135]) ^ (layer1_outputs[11748]));
    assign layer2_outputs[4802] = ~(layer1_outputs[9437]);
    assign layer2_outputs[4803] = ~(layer1_outputs[10265]);
    assign layer2_outputs[4804] = ~((layer1_outputs[6476]) | (layer1_outputs[11072]));
    assign layer2_outputs[4805] = ~(layer1_outputs[657]);
    assign layer2_outputs[4806] = ~(layer1_outputs[1578]);
    assign layer2_outputs[4807] = ~(layer1_outputs[10268]);
    assign layer2_outputs[4808] = layer1_outputs[168];
    assign layer2_outputs[4809] = layer1_outputs[6832];
    assign layer2_outputs[4810] = ~((layer1_outputs[7417]) & (layer1_outputs[11629]));
    assign layer2_outputs[4811] = (layer1_outputs[12614]) & ~(layer1_outputs[5084]);
    assign layer2_outputs[4812] = (layer1_outputs[7602]) | (layer1_outputs[10842]);
    assign layer2_outputs[4813] = ~((layer1_outputs[7940]) ^ (layer1_outputs[1273]));
    assign layer2_outputs[4814] = (layer1_outputs[6406]) & (layer1_outputs[2530]);
    assign layer2_outputs[4815] = (layer1_outputs[8828]) & ~(layer1_outputs[3601]);
    assign layer2_outputs[4816] = layer1_outputs[7242];
    assign layer2_outputs[4817] = layer1_outputs[7684];
    assign layer2_outputs[4818] = (layer1_outputs[9192]) ^ (layer1_outputs[5078]);
    assign layer2_outputs[4819] = ~((layer1_outputs[6834]) ^ (layer1_outputs[9513]));
    assign layer2_outputs[4820] = ~(layer1_outputs[6357]);
    assign layer2_outputs[4821] = layer1_outputs[12058];
    assign layer2_outputs[4822] = ~(layer1_outputs[7694]);
    assign layer2_outputs[4823] = (layer1_outputs[7867]) ^ (layer1_outputs[8907]);
    assign layer2_outputs[4824] = ~((layer1_outputs[4387]) ^ (layer1_outputs[8518]));
    assign layer2_outputs[4825] = layer1_outputs[6965];
    assign layer2_outputs[4826] = ~(layer1_outputs[1688]);
    assign layer2_outputs[4827] = ~(layer1_outputs[10951]) | (layer1_outputs[1113]);
    assign layer2_outputs[4828] = layer1_outputs[3814];
    assign layer2_outputs[4829] = ~(layer1_outputs[9872]) | (layer1_outputs[11546]);
    assign layer2_outputs[4830] = ~((layer1_outputs[1310]) ^ (layer1_outputs[9302]));
    assign layer2_outputs[4831] = (layer1_outputs[2569]) & ~(layer1_outputs[5471]);
    assign layer2_outputs[4832] = ~(layer1_outputs[7692]);
    assign layer2_outputs[4833] = layer1_outputs[10684];
    assign layer2_outputs[4834] = ~(layer1_outputs[4938]);
    assign layer2_outputs[4835] = (layer1_outputs[3979]) ^ (layer1_outputs[8448]);
    assign layer2_outputs[4836] = (layer1_outputs[1756]) | (layer1_outputs[1530]);
    assign layer2_outputs[4837] = layer1_outputs[4342];
    assign layer2_outputs[4838] = layer1_outputs[12103];
    assign layer2_outputs[4839] = (layer1_outputs[8510]) ^ (layer1_outputs[1303]);
    assign layer2_outputs[4840] = ~((layer1_outputs[343]) ^ (layer1_outputs[1454]));
    assign layer2_outputs[4841] = layer1_outputs[12520];
    assign layer2_outputs[4842] = ~(layer1_outputs[12270]);
    assign layer2_outputs[4843] = (layer1_outputs[7022]) | (layer1_outputs[12707]);
    assign layer2_outputs[4844] = (layer1_outputs[8469]) ^ (layer1_outputs[2246]);
    assign layer2_outputs[4845] = ~((layer1_outputs[12105]) ^ (layer1_outputs[441]));
    assign layer2_outputs[4846] = ~(layer1_outputs[561]);
    assign layer2_outputs[4847] = (layer1_outputs[5136]) & (layer1_outputs[9270]);
    assign layer2_outputs[4848] = ~((layer1_outputs[6145]) ^ (layer1_outputs[2190]));
    assign layer2_outputs[4849] = ~(layer1_outputs[10008]) | (layer1_outputs[12332]);
    assign layer2_outputs[4850] = ~((layer1_outputs[8197]) & (layer1_outputs[1392]));
    assign layer2_outputs[4851] = ~(layer1_outputs[8463]);
    assign layer2_outputs[4852] = ~(layer1_outputs[9684]);
    assign layer2_outputs[4853] = (layer1_outputs[3521]) & ~(layer1_outputs[7040]);
    assign layer2_outputs[4854] = layer1_outputs[7485];
    assign layer2_outputs[4855] = ~((layer1_outputs[3132]) & (layer1_outputs[4155]));
    assign layer2_outputs[4856] = layer1_outputs[1014];
    assign layer2_outputs[4857] = (layer1_outputs[3503]) & ~(layer1_outputs[10613]);
    assign layer2_outputs[4858] = layer1_outputs[2844];
    assign layer2_outputs[4859] = ~(layer1_outputs[7729]);
    assign layer2_outputs[4860] = ~((layer1_outputs[1463]) | (layer1_outputs[5612]));
    assign layer2_outputs[4861] = ~(layer1_outputs[4211]);
    assign layer2_outputs[4862] = (layer1_outputs[10359]) & ~(layer1_outputs[7236]);
    assign layer2_outputs[4863] = (layer1_outputs[9145]) ^ (layer1_outputs[11990]);
    assign layer2_outputs[4864] = ~((layer1_outputs[6254]) ^ (layer1_outputs[5378]));
    assign layer2_outputs[4865] = layer1_outputs[827];
    assign layer2_outputs[4866] = (layer1_outputs[12432]) ^ (layer1_outputs[318]);
    assign layer2_outputs[4867] = (layer1_outputs[3597]) & (layer1_outputs[10349]);
    assign layer2_outputs[4868] = layer1_outputs[3737];
    assign layer2_outputs[4869] = ~(layer1_outputs[542]);
    assign layer2_outputs[4870] = layer1_outputs[12260];
    assign layer2_outputs[4871] = (layer1_outputs[8434]) & (layer1_outputs[6715]);
    assign layer2_outputs[4872] = (layer1_outputs[7403]) & ~(layer1_outputs[7278]);
    assign layer2_outputs[4873] = ~(layer1_outputs[10920]);
    assign layer2_outputs[4874] = ~(layer1_outputs[9033]) | (layer1_outputs[5903]);
    assign layer2_outputs[4875] = (layer1_outputs[588]) ^ (layer1_outputs[10707]);
    assign layer2_outputs[4876] = ~(layer1_outputs[10134]) | (layer1_outputs[3608]);
    assign layer2_outputs[4877] = layer1_outputs[2241];
    assign layer2_outputs[4878] = layer1_outputs[8463];
    assign layer2_outputs[4879] = layer1_outputs[11410];
    assign layer2_outputs[4880] = ~((layer1_outputs[6366]) ^ (layer1_outputs[2646]));
    assign layer2_outputs[4881] = layer1_outputs[12766];
    assign layer2_outputs[4882] = ~(layer1_outputs[9375]);
    assign layer2_outputs[4883] = ~((layer1_outputs[5813]) | (layer1_outputs[946]));
    assign layer2_outputs[4884] = ~(layer1_outputs[8103]);
    assign layer2_outputs[4885] = layer1_outputs[9900];
    assign layer2_outputs[4886] = ~(layer1_outputs[581]);
    assign layer2_outputs[4887] = (layer1_outputs[4664]) & ~(layer1_outputs[7811]);
    assign layer2_outputs[4888] = ~(layer1_outputs[3364]);
    assign layer2_outputs[4889] = ~(layer1_outputs[9982]);
    assign layer2_outputs[4890] = (layer1_outputs[5079]) & ~(layer1_outputs[914]);
    assign layer2_outputs[4891] = layer1_outputs[2165];
    assign layer2_outputs[4892] = (layer1_outputs[3941]) & (layer1_outputs[12419]);
    assign layer2_outputs[4893] = (layer1_outputs[6396]) & ~(layer1_outputs[10754]);
    assign layer2_outputs[4894] = (layer1_outputs[1396]) ^ (layer1_outputs[8094]);
    assign layer2_outputs[4895] = ~((layer1_outputs[3180]) & (layer1_outputs[9591]));
    assign layer2_outputs[4896] = layer1_outputs[3528];
    assign layer2_outputs[4897] = ~((layer1_outputs[8429]) & (layer1_outputs[10465]));
    assign layer2_outputs[4898] = (layer1_outputs[6777]) ^ (layer1_outputs[11049]);
    assign layer2_outputs[4899] = ~(layer1_outputs[6053]) | (layer1_outputs[5363]);
    assign layer2_outputs[4900] = layer1_outputs[8857];
    assign layer2_outputs[4901] = layer1_outputs[9443];
    assign layer2_outputs[4902] = (layer1_outputs[7723]) & ~(layer1_outputs[12620]);
    assign layer2_outputs[4903] = ~(layer1_outputs[7659]);
    assign layer2_outputs[4904] = (layer1_outputs[5071]) | (layer1_outputs[1839]);
    assign layer2_outputs[4905] = (layer1_outputs[7094]) & ~(layer1_outputs[11505]);
    assign layer2_outputs[4906] = layer1_outputs[9704];
    assign layer2_outputs[4907] = layer1_outputs[10315];
    assign layer2_outputs[4908] = (layer1_outputs[9809]) ^ (layer1_outputs[1686]);
    assign layer2_outputs[4909] = (layer1_outputs[2331]) | (layer1_outputs[8057]);
    assign layer2_outputs[4910] = (layer1_outputs[3928]) & (layer1_outputs[3039]);
    assign layer2_outputs[4911] = layer1_outputs[1621];
    assign layer2_outputs[4912] = (layer1_outputs[9937]) ^ (layer1_outputs[2493]);
    assign layer2_outputs[4913] = ~(layer1_outputs[3483]);
    assign layer2_outputs[4914] = layer1_outputs[3831];
    assign layer2_outputs[4915] = ~((layer1_outputs[4404]) ^ (layer1_outputs[8410]));
    assign layer2_outputs[4916] = layer1_outputs[11750];
    assign layer2_outputs[4917] = ~(layer1_outputs[11642]);
    assign layer2_outputs[4918] = layer1_outputs[9074];
    assign layer2_outputs[4919] = ~(layer1_outputs[12102]);
    assign layer2_outputs[4920] = (layer1_outputs[11167]) & (layer1_outputs[5528]);
    assign layer2_outputs[4921] = ~((layer1_outputs[11556]) | (layer1_outputs[2780]));
    assign layer2_outputs[4922] = ~((layer1_outputs[5385]) ^ (layer1_outputs[1683]));
    assign layer2_outputs[4923] = ~(layer1_outputs[3647]);
    assign layer2_outputs[4924] = ~(layer1_outputs[4057]);
    assign layer2_outputs[4925] = layer1_outputs[2355];
    assign layer2_outputs[4926] = ~(layer1_outputs[4097]);
    assign layer2_outputs[4927] = ~((layer1_outputs[5636]) | (layer1_outputs[6486]));
    assign layer2_outputs[4928] = ~(layer1_outputs[1690]);
    assign layer2_outputs[4929] = ~(layer1_outputs[11948]);
    assign layer2_outputs[4930] = ~((layer1_outputs[1715]) ^ (layer1_outputs[6373]));
    assign layer2_outputs[4931] = ~(layer1_outputs[7445]);
    assign layer2_outputs[4932] = (layer1_outputs[2089]) & ~(layer1_outputs[6790]);
    assign layer2_outputs[4933] = ~(layer1_outputs[4956]) | (layer1_outputs[7648]);
    assign layer2_outputs[4934] = ~((layer1_outputs[3564]) ^ (layer1_outputs[5406]));
    assign layer2_outputs[4935] = layer1_outputs[9398];
    assign layer2_outputs[4936] = (layer1_outputs[1611]) & ~(layer1_outputs[894]);
    assign layer2_outputs[4937] = ~(layer1_outputs[5689]);
    assign layer2_outputs[4938] = layer1_outputs[7885];
    assign layer2_outputs[4939] = layer1_outputs[9072];
    assign layer2_outputs[4940] = ~(layer1_outputs[10595]);
    assign layer2_outputs[4941] = ~((layer1_outputs[5477]) ^ (layer1_outputs[1734]));
    assign layer2_outputs[4942] = (layer1_outputs[6871]) ^ (layer1_outputs[9820]);
    assign layer2_outputs[4943] = layer1_outputs[7235];
    assign layer2_outputs[4944] = (layer1_outputs[9750]) ^ (layer1_outputs[3049]);
    assign layer2_outputs[4945] = layer1_outputs[36];
    assign layer2_outputs[4946] = layer1_outputs[11462];
    assign layer2_outputs[4947] = (layer1_outputs[774]) | (layer1_outputs[5257]);
    assign layer2_outputs[4948] = ~(layer1_outputs[11882]);
    assign layer2_outputs[4949] = (layer1_outputs[4843]) | (layer1_outputs[10467]);
    assign layer2_outputs[4950] = ~(layer1_outputs[6273]);
    assign layer2_outputs[4951] = ~(layer1_outputs[6846]);
    assign layer2_outputs[4952] = layer1_outputs[5359];
    assign layer2_outputs[4953] = (layer1_outputs[5242]) ^ (layer1_outputs[2009]);
    assign layer2_outputs[4954] = (layer1_outputs[5270]) ^ (layer1_outputs[10833]);
    assign layer2_outputs[4955] = (layer1_outputs[5346]) & ~(layer1_outputs[2529]);
    assign layer2_outputs[4956] = layer1_outputs[2633];
    assign layer2_outputs[4957] = ~((layer1_outputs[2641]) | (layer1_outputs[10878]));
    assign layer2_outputs[4958] = (layer1_outputs[7631]) & (layer1_outputs[7537]);
    assign layer2_outputs[4959] = layer1_outputs[1258];
    assign layer2_outputs[4960] = (layer1_outputs[1720]) & ~(layer1_outputs[6071]);
    assign layer2_outputs[4961] = ~((layer1_outputs[11474]) | (layer1_outputs[2002]));
    assign layer2_outputs[4962] = layer1_outputs[11921];
    assign layer2_outputs[4963] = ~(layer1_outputs[2139]);
    assign layer2_outputs[4964] = (layer1_outputs[10092]) & ~(layer1_outputs[12644]);
    assign layer2_outputs[4965] = (layer1_outputs[2311]) & (layer1_outputs[3110]);
    assign layer2_outputs[4966] = ~(layer1_outputs[12565]);
    assign layer2_outputs[4967] = ~((layer1_outputs[5556]) | (layer1_outputs[4500]));
    assign layer2_outputs[4968] = ~(layer1_outputs[8574]) | (layer1_outputs[11412]);
    assign layer2_outputs[4969] = (layer1_outputs[5820]) | (layer1_outputs[7165]);
    assign layer2_outputs[4970] = layer1_outputs[10575];
    assign layer2_outputs[4971] = layer1_outputs[12513];
    assign layer2_outputs[4972] = ~(layer1_outputs[7948]) | (layer1_outputs[5327]);
    assign layer2_outputs[4973] = ~((layer1_outputs[11576]) ^ (layer1_outputs[9622]));
    assign layer2_outputs[4974] = ~(layer1_outputs[6034]);
    assign layer2_outputs[4975] = layer1_outputs[6801];
    assign layer2_outputs[4976] = ~(layer1_outputs[12324]);
    assign layer2_outputs[4977] = (layer1_outputs[3791]) & ~(layer1_outputs[7760]);
    assign layer2_outputs[4978] = ~(layer1_outputs[12797]);
    assign layer2_outputs[4979] = ~(layer1_outputs[6931]);
    assign layer2_outputs[4980] = ~(layer1_outputs[2701]);
    assign layer2_outputs[4981] = layer1_outputs[3219];
    assign layer2_outputs[4982] = (layer1_outputs[3359]) & ~(layer1_outputs[1233]);
    assign layer2_outputs[4983] = (layer1_outputs[5644]) & (layer1_outputs[11345]);
    assign layer2_outputs[4984] = ~(layer1_outputs[1501]) | (layer1_outputs[3486]);
    assign layer2_outputs[4985] = ~(layer1_outputs[11942]);
    assign layer2_outputs[4986] = ~((layer1_outputs[12208]) & (layer1_outputs[5250]));
    assign layer2_outputs[4987] = layer1_outputs[4478];
    assign layer2_outputs[4988] = ~(layer1_outputs[9787]);
    assign layer2_outputs[4989] = ~(layer1_outputs[11468]);
    assign layer2_outputs[4990] = layer1_outputs[12096];
    assign layer2_outputs[4991] = (layer1_outputs[12530]) | (layer1_outputs[11651]);
    assign layer2_outputs[4992] = (layer1_outputs[6783]) | (layer1_outputs[2630]);
    assign layer2_outputs[4993] = ~(layer1_outputs[12639]) | (layer1_outputs[7539]);
    assign layer2_outputs[4994] = ~(layer1_outputs[2399]) | (layer1_outputs[10101]);
    assign layer2_outputs[4995] = (layer1_outputs[636]) | (layer1_outputs[11160]);
    assign layer2_outputs[4996] = (layer1_outputs[3835]) & ~(layer1_outputs[7122]);
    assign layer2_outputs[4997] = layer1_outputs[5050];
    assign layer2_outputs[4998] = ~((layer1_outputs[5129]) & (layer1_outputs[7122]));
    assign layer2_outputs[4999] = layer1_outputs[5863];
    assign layer2_outputs[5000] = layer1_outputs[1015];
    assign layer2_outputs[5001] = (layer1_outputs[7373]) & ~(layer1_outputs[8131]);
    assign layer2_outputs[5002] = ~(layer1_outputs[2007]);
    assign layer2_outputs[5003] = ~(layer1_outputs[7410]);
    assign layer2_outputs[5004] = ~((layer1_outputs[6050]) & (layer1_outputs[12051]));
    assign layer2_outputs[5005] = ~(layer1_outputs[3369]) | (layer1_outputs[6508]);
    assign layer2_outputs[5006] = ~((layer1_outputs[11480]) & (layer1_outputs[2522]));
    assign layer2_outputs[5007] = layer1_outputs[5180];
    assign layer2_outputs[5008] = layer1_outputs[12038];
    assign layer2_outputs[5009] = ~(layer1_outputs[9102]);
    assign layer2_outputs[5010] = layer1_outputs[7123];
    assign layer2_outputs[5011] = ~(layer1_outputs[12181]);
    assign layer2_outputs[5012] = (layer1_outputs[8004]) ^ (layer1_outputs[912]);
    assign layer2_outputs[5013] = ~(layer1_outputs[2694]);
    assign layer2_outputs[5014] = ~(layer1_outputs[10808]);
    assign layer2_outputs[5015] = (layer1_outputs[11780]) & ~(layer1_outputs[12723]);
    assign layer2_outputs[5016] = (layer1_outputs[2585]) & ~(layer1_outputs[7225]);
    assign layer2_outputs[5017] = (layer1_outputs[11188]) & ~(layer1_outputs[4495]);
    assign layer2_outputs[5018] = ~(layer1_outputs[7119]);
    assign layer2_outputs[5019] = ~((layer1_outputs[406]) & (layer1_outputs[8578]));
    assign layer2_outputs[5020] = ~(layer1_outputs[11372]) | (layer1_outputs[10473]);
    assign layer2_outputs[5021] = layer1_outputs[3706];
    assign layer2_outputs[5022] = (layer1_outputs[12001]) & (layer1_outputs[2011]);
    assign layer2_outputs[5023] = layer1_outputs[11345];
    assign layer2_outputs[5024] = (layer1_outputs[11617]) ^ (layer1_outputs[4714]);
    assign layer2_outputs[5025] = ~((layer1_outputs[12080]) ^ (layer1_outputs[4188]));
    assign layer2_outputs[5026] = (layer1_outputs[9541]) ^ (layer1_outputs[7047]);
    assign layer2_outputs[5027] = ~((layer1_outputs[10950]) | (layer1_outputs[7704]));
    assign layer2_outputs[5028] = ~((layer1_outputs[10605]) | (layer1_outputs[8187]));
    assign layer2_outputs[5029] = ~(layer1_outputs[7359]);
    assign layer2_outputs[5030] = layer1_outputs[11312];
    assign layer2_outputs[5031] = ~((layer1_outputs[8595]) | (layer1_outputs[12287]));
    assign layer2_outputs[5032] = ~((layer1_outputs[3954]) & (layer1_outputs[10275]));
    assign layer2_outputs[5033] = layer1_outputs[7091];
    assign layer2_outputs[5034] = (layer1_outputs[7411]) ^ (layer1_outputs[500]);
    assign layer2_outputs[5035] = layer1_outputs[4197];
    assign layer2_outputs[5036] = (layer1_outputs[9164]) ^ (layer1_outputs[182]);
    assign layer2_outputs[5037] = ~(layer1_outputs[2541]);
    assign layer2_outputs[5038] = ~(layer1_outputs[3477]);
    assign layer2_outputs[5039] = layer1_outputs[8040];
    assign layer2_outputs[5040] = (layer1_outputs[8964]) ^ (layer1_outputs[11271]);
    assign layer2_outputs[5041] = layer1_outputs[12533];
    assign layer2_outputs[5042] = ~((layer1_outputs[9327]) | (layer1_outputs[704]));
    assign layer2_outputs[5043] = ~(layer1_outputs[4146]);
    assign layer2_outputs[5044] = layer1_outputs[10487];
    assign layer2_outputs[5045] = ~((layer1_outputs[403]) ^ (layer1_outputs[3958]));
    assign layer2_outputs[5046] = ~(layer1_outputs[3392]) | (layer1_outputs[7945]);
    assign layer2_outputs[5047] = ~(layer1_outputs[4602]);
    assign layer2_outputs[5048] = layer1_outputs[8313];
    assign layer2_outputs[5049] = (layer1_outputs[6697]) & (layer1_outputs[12749]);
    assign layer2_outputs[5050] = (layer1_outputs[456]) & ~(layer1_outputs[2582]);
    assign layer2_outputs[5051] = ~(layer1_outputs[2660]);
    assign layer2_outputs[5052] = ~(layer1_outputs[4656]);
    assign layer2_outputs[5053] = layer1_outputs[1599];
    assign layer2_outputs[5054] = layer1_outputs[12034];
    assign layer2_outputs[5055] = (layer1_outputs[379]) & ~(layer1_outputs[3015]);
    assign layer2_outputs[5056] = layer1_outputs[10140];
    assign layer2_outputs[5057] = ~(layer1_outputs[9305]);
    assign layer2_outputs[5058] = ~(layer1_outputs[12419]);
    assign layer2_outputs[5059] = ~(layer1_outputs[12445]);
    assign layer2_outputs[5060] = ~(layer1_outputs[6583]);
    assign layer2_outputs[5061] = ~(layer1_outputs[10562]);
    assign layer2_outputs[5062] = (layer1_outputs[1604]) & ~(layer1_outputs[10524]);
    assign layer2_outputs[5063] = (layer1_outputs[9692]) & (layer1_outputs[6079]);
    assign layer2_outputs[5064] = ~((layer1_outputs[11938]) | (layer1_outputs[798]));
    assign layer2_outputs[5065] = (layer1_outputs[4334]) & ~(layer1_outputs[12038]);
    assign layer2_outputs[5066] = ~(layer1_outputs[10675]);
    assign layer2_outputs[5067] = layer1_outputs[1440];
    assign layer2_outputs[5068] = ~((layer1_outputs[3465]) | (layer1_outputs[10656]));
    assign layer2_outputs[5069] = layer1_outputs[7932];
    assign layer2_outputs[5070] = ~((layer1_outputs[9489]) | (layer1_outputs[4269]));
    assign layer2_outputs[5071] = (layer1_outputs[3898]) & (layer1_outputs[4789]);
    assign layer2_outputs[5072] = layer1_outputs[6158];
    assign layer2_outputs[5073] = (layer1_outputs[9716]) & ~(layer1_outputs[11411]);
    assign layer2_outputs[5074] = 1'b0;
    assign layer2_outputs[5075] = (layer1_outputs[2272]) | (layer1_outputs[6806]);
    assign layer2_outputs[5076] = ~(layer1_outputs[3228]);
    assign layer2_outputs[5077] = ~(layer1_outputs[2451]);
    assign layer2_outputs[5078] = ~((layer1_outputs[6524]) & (layer1_outputs[6788]));
    assign layer2_outputs[5079] = ~(layer1_outputs[10862]) | (layer1_outputs[5255]);
    assign layer2_outputs[5080] = (layer1_outputs[4367]) ^ (layer1_outputs[10245]);
    assign layer2_outputs[5081] = layer1_outputs[3735];
    assign layer2_outputs[5082] = layer1_outputs[3984];
    assign layer2_outputs[5083] = ~(layer1_outputs[4825]);
    assign layer2_outputs[5084] = (layer1_outputs[10052]) ^ (layer1_outputs[8281]);
    assign layer2_outputs[5085] = ~(layer1_outputs[1552]);
    assign layer2_outputs[5086] = (layer1_outputs[4499]) & ~(layer1_outputs[9198]);
    assign layer2_outputs[5087] = ~(layer1_outputs[7503]);
    assign layer2_outputs[5088] = ~(layer1_outputs[3247]) | (layer1_outputs[6518]);
    assign layer2_outputs[5089] = layer1_outputs[2133];
    assign layer2_outputs[5090] = ~(layer1_outputs[1922]) | (layer1_outputs[4403]);
    assign layer2_outputs[5091] = layer1_outputs[2354];
    assign layer2_outputs[5092] = ~((layer1_outputs[8113]) ^ (layer1_outputs[12241]));
    assign layer2_outputs[5093] = (layer1_outputs[6532]) | (layer1_outputs[9895]);
    assign layer2_outputs[5094] = layer1_outputs[4434];
    assign layer2_outputs[5095] = layer1_outputs[9285];
    assign layer2_outputs[5096] = (layer1_outputs[9011]) ^ (layer1_outputs[10592]);
    assign layer2_outputs[5097] = (layer1_outputs[6380]) & ~(layer1_outputs[8337]);
    assign layer2_outputs[5098] = ~(layer1_outputs[333]) | (layer1_outputs[5171]);
    assign layer2_outputs[5099] = ~(layer1_outputs[6437]) | (layer1_outputs[7546]);
    assign layer2_outputs[5100] = layer1_outputs[11129];
    assign layer2_outputs[5101] = ~(layer1_outputs[7837]) | (layer1_outputs[7138]);
    assign layer2_outputs[5102] = (layer1_outputs[4352]) | (layer1_outputs[1174]);
    assign layer2_outputs[5103] = (layer1_outputs[3891]) & ~(layer1_outputs[10118]);
    assign layer2_outputs[5104] = layer1_outputs[4943];
    assign layer2_outputs[5105] = (layer1_outputs[5332]) ^ (layer1_outputs[2424]);
    assign layer2_outputs[5106] = ~(layer1_outputs[8825]) | (layer1_outputs[10199]);
    assign layer2_outputs[5107] = (layer1_outputs[2052]) ^ (layer1_outputs[8891]);
    assign layer2_outputs[5108] = layer1_outputs[8192];
    assign layer2_outputs[5109] = ~(layer1_outputs[11925]);
    assign layer2_outputs[5110] = ~((layer1_outputs[1262]) ^ (layer1_outputs[478]));
    assign layer2_outputs[5111] = layer1_outputs[6702];
    assign layer2_outputs[5112] = (layer1_outputs[10927]) & ~(layer1_outputs[9797]);
    assign layer2_outputs[5113] = ~(layer1_outputs[2759]);
    assign layer2_outputs[5114] = (layer1_outputs[8754]) ^ (layer1_outputs[7478]);
    assign layer2_outputs[5115] = (layer1_outputs[5683]) | (layer1_outputs[4762]);
    assign layer2_outputs[5116] = ~(layer1_outputs[9908]);
    assign layer2_outputs[5117] = ~(layer1_outputs[5673]);
    assign layer2_outputs[5118] = layer1_outputs[10070];
    assign layer2_outputs[5119] = ~(layer1_outputs[11665]);
    assign layer2_outputs[5120] = ~(layer1_outputs[10532]) | (layer1_outputs[9423]);
    assign layer2_outputs[5121] = (layer1_outputs[9155]) ^ (layer1_outputs[6848]);
    assign layer2_outputs[5122] = layer1_outputs[12228];
    assign layer2_outputs[5123] = ~((layer1_outputs[4663]) ^ (layer1_outputs[4353]));
    assign layer2_outputs[5124] = ~(layer1_outputs[10451]);
    assign layer2_outputs[5125] = ~(layer1_outputs[11841]) | (layer1_outputs[12219]);
    assign layer2_outputs[5126] = ~(layer1_outputs[7768]);
    assign layer2_outputs[5127] = (layer1_outputs[10347]) & ~(layer1_outputs[2211]);
    assign layer2_outputs[5128] = layer1_outputs[12410];
    assign layer2_outputs[5129] = ~(layer1_outputs[298]);
    assign layer2_outputs[5130] = 1'b0;
    assign layer2_outputs[5131] = layer1_outputs[5838];
    assign layer2_outputs[5132] = (layer1_outputs[6320]) ^ (layer1_outputs[11231]);
    assign layer2_outputs[5133] = layer1_outputs[12741];
    assign layer2_outputs[5134] = layer1_outputs[12760];
    assign layer2_outputs[5135] = layer1_outputs[11307];
    assign layer2_outputs[5136] = layer1_outputs[6718];
    assign layer2_outputs[5137] = layer1_outputs[2726];
    assign layer2_outputs[5138] = ~(layer1_outputs[10926]);
    assign layer2_outputs[5139] = ~(layer1_outputs[2220]);
    assign layer2_outputs[5140] = layer1_outputs[3211];
    assign layer2_outputs[5141] = (layer1_outputs[3289]) & ~(layer1_outputs[1911]);
    assign layer2_outputs[5142] = ~(layer1_outputs[3404]);
    assign layer2_outputs[5143] = (layer1_outputs[10303]) ^ (layer1_outputs[7703]);
    assign layer2_outputs[5144] = ~((layer1_outputs[2523]) ^ (layer1_outputs[1840]));
    assign layer2_outputs[5145] = ~(layer1_outputs[6688]) | (layer1_outputs[1377]);
    assign layer2_outputs[5146] = ~(layer1_outputs[7645]);
    assign layer2_outputs[5147] = ~((layer1_outputs[9956]) ^ (layer1_outputs[3390]));
    assign layer2_outputs[5148] = layer1_outputs[7003];
    assign layer2_outputs[5149] = (layer1_outputs[3015]) & ~(layer1_outputs[10489]);
    assign layer2_outputs[5150] = ~(layer1_outputs[5963]) | (layer1_outputs[12089]);
    assign layer2_outputs[5151] = layer1_outputs[4271];
    assign layer2_outputs[5152] = ~((layer1_outputs[2784]) ^ (layer1_outputs[5218]));
    assign layer2_outputs[5153] = layer1_outputs[11545];
    assign layer2_outputs[5154] = (layer1_outputs[10981]) ^ (layer1_outputs[7537]);
    assign layer2_outputs[5155] = ~((layer1_outputs[12600]) ^ (layer1_outputs[917]));
    assign layer2_outputs[5156] = ~(layer1_outputs[8634]);
    assign layer2_outputs[5157] = layer1_outputs[1198];
    assign layer2_outputs[5158] = ~(layer1_outputs[11806]);
    assign layer2_outputs[5159] = layer1_outputs[6704];
    assign layer2_outputs[5160] = (layer1_outputs[12337]) ^ (layer1_outputs[6482]);
    assign layer2_outputs[5161] = (layer1_outputs[9358]) ^ (layer1_outputs[5764]);
    assign layer2_outputs[5162] = (layer1_outputs[10331]) & (layer1_outputs[10484]);
    assign layer2_outputs[5163] = layer1_outputs[8327];
    assign layer2_outputs[5164] = ~((layer1_outputs[12647]) ^ (layer1_outputs[10916]));
    assign layer2_outputs[5165] = layer1_outputs[6483];
    assign layer2_outputs[5166] = ~(layer1_outputs[11074]) | (layer1_outputs[7345]);
    assign layer2_outputs[5167] = (layer1_outputs[2914]) ^ (layer1_outputs[447]);
    assign layer2_outputs[5168] = ~((layer1_outputs[7754]) & (layer1_outputs[8094]));
    assign layer2_outputs[5169] = layer1_outputs[1655];
    assign layer2_outputs[5170] = ~(layer1_outputs[4330]);
    assign layer2_outputs[5171] = ~(layer1_outputs[7572]);
    assign layer2_outputs[5172] = layer1_outputs[6932];
    assign layer2_outputs[5173] = layer1_outputs[4593];
    assign layer2_outputs[5174] = ~((layer1_outputs[382]) ^ (layer1_outputs[11794]));
    assign layer2_outputs[5175] = ~(layer1_outputs[5722]);
    assign layer2_outputs[5176] = layer1_outputs[326];
    assign layer2_outputs[5177] = ~((layer1_outputs[9393]) | (layer1_outputs[5596]));
    assign layer2_outputs[5178] = ~(layer1_outputs[2900]) | (layer1_outputs[11380]);
    assign layer2_outputs[5179] = layer1_outputs[1180];
    assign layer2_outputs[5180] = ~(layer1_outputs[301]);
    assign layer2_outputs[5181] = ~(layer1_outputs[8254]) | (layer1_outputs[3528]);
    assign layer2_outputs[5182] = (layer1_outputs[336]) ^ (layer1_outputs[10843]);
    assign layer2_outputs[5183] = (layer1_outputs[2113]) ^ (layer1_outputs[9029]);
    assign layer2_outputs[5184] = ~(layer1_outputs[5496]);
    assign layer2_outputs[5185] = layer1_outputs[12788];
    assign layer2_outputs[5186] = ~(layer1_outputs[931]) | (layer1_outputs[10536]);
    assign layer2_outputs[5187] = ~((layer1_outputs[7685]) | (layer1_outputs[3551]));
    assign layer2_outputs[5188] = (layer1_outputs[5021]) ^ (layer1_outputs[3364]);
    assign layer2_outputs[5189] = ~(layer1_outputs[4927]) | (layer1_outputs[4815]);
    assign layer2_outputs[5190] = ~((layer1_outputs[3673]) ^ (layer1_outputs[4216]));
    assign layer2_outputs[5191] = layer1_outputs[8145];
    assign layer2_outputs[5192] = ~(layer1_outputs[6082]);
    assign layer2_outputs[5193] = layer1_outputs[5892];
    assign layer2_outputs[5194] = ~(layer1_outputs[2126]) | (layer1_outputs[10761]);
    assign layer2_outputs[5195] = ~(layer1_outputs[11600]);
    assign layer2_outputs[5196] = (layer1_outputs[11943]) ^ (layer1_outputs[72]);
    assign layer2_outputs[5197] = ~((layer1_outputs[395]) ^ (layer1_outputs[5174]));
    assign layer2_outputs[5198] = (layer1_outputs[2028]) & (layer1_outputs[367]);
    assign layer2_outputs[5199] = ~(layer1_outputs[12677]);
    assign layer2_outputs[5200] = layer1_outputs[10123];
    assign layer2_outputs[5201] = layer1_outputs[5311];
    assign layer2_outputs[5202] = ~(layer1_outputs[3178]) | (layer1_outputs[7232]);
    assign layer2_outputs[5203] = ~(layer1_outputs[8705]);
    assign layer2_outputs[5204] = ~(layer1_outputs[10568]) | (layer1_outputs[7084]);
    assign layer2_outputs[5205] = ~(layer1_outputs[6279]);
    assign layer2_outputs[5206] = layer1_outputs[10713];
    assign layer2_outputs[5207] = ~(layer1_outputs[1058]);
    assign layer2_outputs[5208] = ~(layer1_outputs[1882]);
    assign layer2_outputs[5209] = ~((layer1_outputs[11461]) & (layer1_outputs[5006]));
    assign layer2_outputs[5210] = ~((layer1_outputs[267]) & (layer1_outputs[3119]));
    assign layer2_outputs[5211] = layer1_outputs[5794];
    assign layer2_outputs[5212] = (layer1_outputs[8554]) ^ (layer1_outputs[3724]);
    assign layer2_outputs[5213] = (layer1_outputs[11107]) & (layer1_outputs[8560]);
    assign layer2_outputs[5214] = ~(layer1_outputs[3034]);
    assign layer2_outputs[5215] = layer1_outputs[7189];
    assign layer2_outputs[5216] = ~((layer1_outputs[2976]) | (layer1_outputs[1414]));
    assign layer2_outputs[5217] = layer1_outputs[210];
    assign layer2_outputs[5218] = (layer1_outputs[7793]) & ~(layer1_outputs[8410]);
    assign layer2_outputs[5219] = (layer1_outputs[10053]) & ~(layer1_outputs[9040]);
    assign layer2_outputs[5220] = ~(layer1_outputs[3026]);
    assign layer2_outputs[5221] = (layer1_outputs[7682]) ^ (layer1_outputs[9078]);
    assign layer2_outputs[5222] = ~(layer1_outputs[5475]) | (layer1_outputs[6682]);
    assign layer2_outputs[5223] = ~(layer1_outputs[7456]) | (layer1_outputs[6420]);
    assign layer2_outputs[5224] = layer1_outputs[311];
    assign layer2_outputs[5225] = (layer1_outputs[6591]) | (layer1_outputs[8156]);
    assign layer2_outputs[5226] = ~(layer1_outputs[2701]);
    assign layer2_outputs[5227] = ~(layer1_outputs[4117]);
    assign layer2_outputs[5228] = layer1_outputs[12525];
    assign layer2_outputs[5229] = ~(layer1_outputs[1872]);
    assign layer2_outputs[5230] = ~((layer1_outputs[7504]) & (layer1_outputs[11463]));
    assign layer2_outputs[5231] = ~((layer1_outputs[12014]) & (layer1_outputs[5904]));
    assign layer2_outputs[5232] = (layer1_outputs[1772]) & (layer1_outputs[7209]);
    assign layer2_outputs[5233] = ~(layer1_outputs[12635]);
    assign layer2_outputs[5234] = layer1_outputs[6124];
    assign layer2_outputs[5235] = (layer1_outputs[12009]) | (layer1_outputs[6997]);
    assign layer2_outputs[5236] = ~((layer1_outputs[9717]) | (layer1_outputs[3359]));
    assign layer2_outputs[5237] = layer1_outputs[682];
    assign layer2_outputs[5238] = (layer1_outputs[11206]) | (layer1_outputs[2690]);
    assign layer2_outputs[5239] = ~(layer1_outputs[12292]) | (layer1_outputs[1383]);
    assign layer2_outputs[5240] = layer1_outputs[387];
    assign layer2_outputs[5241] = (layer1_outputs[12662]) | (layer1_outputs[5636]);
    assign layer2_outputs[5242] = ~(layer1_outputs[7933]);
    assign layer2_outputs[5243] = ~((layer1_outputs[10411]) | (layer1_outputs[12066]));
    assign layer2_outputs[5244] = ~(layer1_outputs[9496]) | (layer1_outputs[5744]);
    assign layer2_outputs[5245] = ~(layer1_outputs[11264]);
    assign layer2_outputs[5246] = layer1_outputs[11144];
    assign layer2_outputs[5247] = ~((layer1_outputs[321]) | (layer1_outputs[10113]));
    assign layer2_outputs[5248] = ~(layer1_outputs[10244]);
    assign layer2_outputs[5249] = layer1_outputs[172];
    assign layer2_outputs[5250] = ~((layer1_outputs[10680]) ^ (layer1_outputs[5287]));
    assign layer2_outputs[5251] = layer1_outputs[12124];
    assign layer2_outputs[5252] = ~(layer1_outputs[12707]) | (layer1_outputs[4620]);
    assign layer2_outputs[5253] = layer1_outputs[5684];
    assign layer2_outputs[5254] = ~(layer1_outputs[7154]);
    assign layer2_outputs[5255] = (layer1_outputs[1704]) & ~(layer1_outputs[3942]);
    assign layer2_outputs[5256] = ~(layer1_outputs[531]);
    assign layer2_outputs[5257] = layer1_outputs[3781];
    assign layer2_outputs[5258] = (layer1_outputs[4512]) & ~(layer1_outputs[3031]);
    assign layer2_outputs[5259] = (layer1_outputs[8379]) | (layer1_outputs[3041]);
    assign layer2_outputs[5260] = ~(layer1_outputs[12592]);
    assign layer2_outputs[5261] = ~((layer1_outputs[12450]) ^ (layer1_outputs[5219]));
    assign layer2_outputs[5262] = ~((layer1_outputs[8409]) & (layer1_outputs[12783]));
    assign layer2_outputs[5263] = (layer1_outputs[8878]) & ~(layer1_outputs[12067]);
    assign layer2_outputs[5264] = ~(layer1_outputs[11589]);
    assign layer2_outputs[5265] = ~(layer1_outputs[9486]);
    assign layer2_outputs[5266] = ~((layer1_outputs[10530]) & (layer1_outputs[10189]));
    assign layer2_outputs[5267] = ~((layer1_outputs[8806]) | (layer1_outputs[8772]));
    assign layer2_outputs[5268] = 1'b0;
    assign layer2_outputs[5269] = layer1_outputs[4224];
    assign layer2_outputs[5270] = ~(layer1_outputs[8797]);
    assign layer2_outputs[5271] = ~(layer1_outputs[2436]);
    assign layer2_outputs[5272] = ~(layer1_outputs[9517]);
    assign layer2_outputs[5273] = layer1_outputs[9279];
    assign layer2_outputs[5274] = ~(layer1_outputs[4629]) | (layer1_outputs[11331]);
    assign layer2_outputs[5275] = ~((layer1_outputs[10556]) & (layer1_outputs[5919]));
    assign layer2_outputs[5276] = (layer1_outputs[7901]) ^ (layer1_outputs[1596]);
    assign layer2_outputs[5277] = layer1_outputs[7998];
    assign layer2_outputs[5278] = ~(layer1_outputs[20]);
    assign layer2_outputs[5279] = (layer1_outputs[4899]) & ~(layer1_outputs[8663]);
    assign layer2_outputs[5280] = ~((layer1_outputs[12329]) & (layer1_outputs[417]));
    assign layer2_outputs[5281] = layer1_outputs[965];
    assign layer2_outputs[5282] = ~(layer1_outputs[833]);
    assign layer2_outputs[5283] = (layer1_outputs[10529]) & ~(layer1_outputs[4151]);
    assign layer2_outputs[5284] = layer1_outputs[12141];
    assign layer2_outputs[5285] = ~((layer1_outputs[6780]) & (layer1_outputs[1784]));
    assign layer2_outputs[5286] = (layer1_outputs[3324]) & ~(layer1_outputs[6424]);
    assign layer2_outputs[5287] = layer1_outputs[1230];
    assign layer2_outputs[5288] = ~(layer1_outputs[6700]);
    assign layer2_outputs[5289] = ~(layer1_outputs[6721]);
    assign layer2_outputs[5290] = ~(layer1_outputs[10622]);
    assign layer2_outputs[5291] = ~(layer1_outputs[12229]) | (layer1_outputs[5261]);
    assign layer2_outputs[5292] = ~(layer1_outputs[5997]);
    assign layer2_outputs[5293] = layer1_outputs[6043];
    assign layer2_outputs[5294] = ~(layer1_outputs[11363]);
    assign layer2_outputs[5295] = ~(layer1_outputs[9212]) | (layer1_outputs[3965]);
    assign layer2_outputs[5296] = layer1_outputs[1730];
    assign layer2_outputs[5297] = layer1_outputs[7199];
    assign layer2_outputs[5298] = (layer1_outputs[11804]) & ~(layer1_outputs[8500]);
    assign layer2_outputs[5299] = ~((layer1_outputs[1061]) & (layer1_outputs[3414]));
    assign layer2_outputs[5300] = ~((layer1_outputs[10410]) ^ (layer1_outputs[8726]));
    assign layer2_outputs[5301] = layer1_outputs[1444];
    assign layer2_outputs[5302] = layer1_outputs[5177];
    assign layer2_outputs[5303] = layer1_outputs[7300];
    assign layer2_outputs[5304] = ~((layer1_outputs[7017]) & (layer1_outputs[3322]));
    assign layer2_outputs[5305] = ~(layer1_outputs[5446]) | (layer1_outputs[9059]);
    assign layer2_outputs[5306] = ~(layer1_outputs[8820]);
    assign layer2_outputs[5307] = layer1_outputs[1353];
    assign layer2_outputs[5308] = ~((layer1_outputs[9791]) ^ (layer1_outputs[9363]));
    assign layer2_outputs[5309] = layer1_outputs[7469];
    assign layer2_outputs[5310] = (layer1_outputs[6293]) & (layer1_outputs[3204]);
    assign layer2_outputs[5311] = ~(layer1_outputs[10779]);
    assign layer2_outputs[5312] = (layer1_outputs[1035]) & (layer1_outputs[1993]);
    assign layer2_outputs[5313] = ~(layer1_outputs[11762]);
    assign layer2_outputs[5314] = (layer1_outputs[2250]) ^ (layer1_outputs[8902]);
    assign layer2_outputs[5315] = ~((layer1_outputs[11065]) & (layer1_outputs[10358]));
    assign layer2_outputs[5316] = layer1_outputs[219];
    assign layer2_outputs[5317] = ~(layer1_outputs[12732]);
    assign layer2_outputs[5318] = (layer1_outputs[10643]) ^ (layer1_outputs[902]);
    assign layer2_outputs[5319] = layer1_outputs[6190];
    assign layer2_outputs[5320] = (layer1_outputs[4470]) ^ (layer1_outputs[1156]);
    assign layer2_outputs[5321] = layer1_outputs[5874];
    assign layer2_outputs[5322] = ~(layer1_outputs[1453]);
    assign layer2_outputs[5323] = (layer1_outputs[9546]) ^ (layer1_outputs[412]);
    assign layer2_outputs[5324] = (layer1_outputs[1424]) | (layer1_outputs[4757]);
    assign layer2_outputs[5325] = ~(layer1_outputs[10550]);
    assign layer2_outputs[5326] = ~((layer1_outputs[8842]) ^ (layer1_outputs[12440]));
    assign layer2_outputs[5327] = ~(layer1_outputs[8354]);
    assign layer2_outputs[5328] = (layer1_outputs[38]) & (layer1_outputs[3263]);
    assign layer2_outputs[5329] = (layer1_outputs[11927]) ^ (layer1_outputs[7326]);
    assign layer2_outputs[5330] = ~(layer1_outputs[7072]);
    assign layer2_outputs[5331] = (layer1_outputs[4024]) & (layer1_outputs[1425]);
    assign layer2_outputs[5332] = layer1_outputs[4655];
    assign layer2_outputs[5333] = ~(layer1_outputs[8146]) | (layer1_outputs[6739]);
    assign layer2_outputs[5334] = ~((layer1_outputs[1792]) & (layer1_outputs[11108]));
    assign layer2_outputs[5335] = ~(layer1_outputs[5229]);
    assign layer2_outputs[5336] = ~(layer1_outputs[8531]) | (layer1_outputs[11816]);
    assign layer2_outputs[5337] = (layer1_outputs[2933]) & ~(layer1_outputs[12278]);
    assign layer2_outputs[5338] = ~(layer1_outputs[1803]) | (layer1_outputs[736]);
    assign layer2_outputs[5339] = ~(layer1_outputs[11163]);
    assign layer2_outputs[5340] = (layer1_outputs[8673]) & (layer1_outputs[61]);
    assign layer2_outputs[5341] = ~((layer1_outputs[9447]) ^ (layer1_outputs[1494]));
    assign layer2_outputs[5342] = ~(layer1_outputs[7728]);
    assign layer2_outputs[5343] = ~(layer1_outputs[6811]);
    assign layer2_outputs[5344] = ~(layer1_outputs[8036]);
    assign layer2_outputs[5345] = (layer1_outputs[11797]) ^ (layer1_outputs[4551]);
    assign layer2_outputs[5346] = ~(layer1_outputs[1656]);
    assign layer2_outputs[5347] = ~(layer1_outputs[5170]);
    assign layer2_outputs[5348] = (layer1_outputs[5774]) & (layer1_outputs[8513]);
    assign layer2_outputs[5349] = ~((layer1_outputs[9910]) & (layer1_outputs[1360]));
    assign layer2_outputs[5350] = (layer1_outputs[2296]) ^ (layer1_outputs[2768]);
    assign layer2_outputs[5351] = (layer1_outputs[5007]) & ~(layer1_outputs[11434]);
    assign layer2_outputs[5352] = layer1_outputs[6382];
    assign layer2_outputs[5353] = (layer1_outputs[3395]) | (layer1_outputs[2337]);
    assign layer2_outputs[5354] = (layer1_outputs[3143]) ^ (layer1_outputs[12075]);
    assign layer2_outputs[5355] = layer1_outputs[10170];
    assign layer2_outputs[5356] = layer1_outputs[2199];
    assign layer2_outputs[5357] = layer1_outputs[12680];
    assign layer2_outputs[5358] = (layer1_outputs[2136]) & ~(layer1_outputs[12770]);
    assign layer2_outputs[5359] = (layer1_outputs[998]) & ~(layer1_outputs[3627]);
    assign layer2_outputs[5360] = layer1_outputs[4227];
    assign layer2_outputs[5361] = (layer1_outputs[12524]) & ~(layer1_outputs[11547]);
    assign layer2_outputs[5362] = ~(layer1_outputs[11735]);
    assign layer2_outputs[5363] = ~(layer1_outputs[9201]);
    assign layer2_outputs[5364] = ~(layer1_outputs[4174]);
    assign layer2_outputs[5365] = (layer1_outputs[3442]) & (layer1_outputs[9121]);
    assign layer2_outputs[5366] = ~(layer1_outputs[7934]);
    assign layer2_outputs[5367] = (layer1_outputs[2545]) | (layer1_outputs[6447]);
    assign layer2_outputs[5368] = layer1_outputs[8808];
    assign layer2_outputs[5369] = ~(layer1_outputs[10915]);
    assign layer2_outputs[5370] = ~((layer1_outputs[9174]) ^ (layer1_outputs[9317]));
    assign layer2_outputs[5371] = (layer1_outputs[4385]) & ~(layer1_outputs[2681]);
    assign layer2_outputs[5372] = (layer1_outputs[1150]) & ~(layer1_outputs[2343]);
    assign layer2_outputs[5373] = (layer1_outputs[8111]) | (layer1_outputs[134]);
    assign layer2_outputs[5374] = ~((layer1_outputs[5119]) | (layer1_outputs[4425]));
    assign layer2_outputs[5375] = ~(layer1_outputs[3429]);
    assign layer2_outputs[5376] = layer1_outputs[11776];
    assign layer2_outputs[5377] = layer1_outputs[2];
    assign layer2_outputs[5378] = layer1_outputs[11714];
    assign layer2_outputs[5379] = ~((layer1_outputs[1116]) & (layer1_outputs[5929]));
    assign layer2_outputs[5380] = layer1_outputs[10326];
    assign layer2_outputs[5381] = ~(layer1_outputs[1767]) | (layer1_outputs[1407]);
    assign layer2_outputs[5382] = (layer1_outputs[7769]) ^ (layer1_outputs[6631]);
    assign layer2_outputs[5383] = ~(layer1_outputs[7897]);
    assign layer2_outputs[5384] = layer1_outputs[5152];
    assign layer2_outputs[5385] = (layer1_outputs[6307]) ^ (layer1_outputs[401]);
    assign layer2_outputs[5386] = (layer1_outputs[4846]) | (layer1_outputs[10312]);
    assign layer2_outputs[5387] = layer1_outputs[10262];
    assign layer2_outputs[5388] = layer1_outputs[5514];
    assign layer2_outputs[5389] = ~(layer1_outputs[9886]);
    assign layer2_outputs[5390] = ~(layer1_outputs[12463]);
    assign layer2_outputs[5391] = ~(layer1_outputs[1628]);
    assign layer2_outputs[5392] = (layer1_outputs[1788]) & (layer1_outputs[11902]);
    assign layer2_outputs[5393] = ~(layer1_outputs[2148]);
    assign layer2_outputs[5394] = layer1_outputs[5841];
    assign layer2_outputs[5395] = ~(layer1_outputs[12585]);
    assign layer2_outputs[5396] = layer1_outputs[2198];
    assign layer2_outputs[5397] = (layer1_outputs[6716]) | (layer1_outputs[3501]);
    assign layer2_outputs[5398] = ~((layer1_outputs[7256]) & (layer1_outputs[2478]));
    assign layer2_outputs[5399] = (layer1_outputs[5943]) ^ (layer1_outputs[7248]);
    assign layer2_outputs[5400] = ~(layer1_outputs[7922]);
    assign layer2_outputs[5401] = (layer1_outputs[5689]) | (layer1_outputs[444]);
    assign layer2_outputs[5402] = ~(layer1_outputs[5199]);
    assign layer2_outputs[5403] = ~(layer1_outputs[5632]);
    assign layer2_outputs[5404] = (layer1_outputs[10937]) & ~(layer1_outputs[4028]);
    assign layer2_outputs[5405] = ~((layer1_outputs[10609]) & (layer1_outputs[3010]));
    assign layer2_outputs[5406] = ~((layer1_outputs[8250]) & (layer1_outputs[8]));
    assign layer2_outputs[5407] = ~(layer1_outputs[4445]) | (layer1_outputs[78]);
    assign layer2_outputs[5408] = (layer1_outputs[9972]) ^ (layer1_outputs[10634]);
    assign layer2_outputs[5409] = layer1_outputs[9990];
    assign layer2_outputs[5410] = layer1_outputs[19];
    assign layer2_outputs[5411] = ~(layer1_outputs[12373]) | (layer1_outputs[3167]);
    assign layer2_outputs[5412] = ~(layer1_outputs[1319]) | (layer1_outputs[9131]);
    assign layer2_outputs[5413] = layer1_outputs[8022];
    assign layer2_outputs[5414] = layer1_outputs[2159];
    assign layer2_outputs[5415] = ~(layer1_outputs[6726]);
    assign layer2_outputs[5416] = ~((layer1_outputs[6475]) & (layer1_outputs[7040]));
    assign layer2_outputs[5417] = layer1_outputs[11472];
    assign layer2_outputs[5418] = ~(layer1_outputs[10917]);
    assign layer2_outputs[5419] = ~(layer1_outputs[6001]);
    assign layer2_outputs[5420] = (layer1_outputs[7231]) | (layer1_outputs[12217]);
    assign layer2_outputs[5421] = (layer1_outputs[12482]) & ~(layer1_outputs[11267]);
    assign layer2_outputs[5422] = layer1_outputs[9949];
    assign layer2_outputs[5423] = layer1_outputs[504];
    assign layer2_outputs[5424] = ~(layer1_outputs[1669]);
    assign layer2_outputs[5425] = layer1_outputs[3045];
    assign layer2_outputs[5426] = ~((layer1_outputs[1565]) | (layer1_outputs[3095]));
    assign layer2_outputs[5427] = layer1_outputs[2380];
    assign layer2_outputs[5428] = layer1_outputs[1019];
    assign layer2_outputs[5429] = (layer1_outputs[10062]) & ~(layer1_outputs[3169]);
    assign layer2_outputs[5430] = ~(layer1_outputs[2563]);
    assign layer2_outputs[5431] = layer1_outputs[10286];
    assign layer2_outputs[5432] = layer1_outputs[4186];
    assign layer2_outputs[5433] = ~(layer1_outputs[9904]);
    assign layer2_outputs[5434] = ~(layer1_outputs[2305]);
    assign layer2_outputs[5435] = ~(layer1_outputs[6167]);
    assign layer2_outputs[5436] = ~(layer1_outputs[6873]) | (layer1_outputs[1962]);
    assign layer2_outputs[5437] = ~(layer1_outputs[3667]);
    assign layer2_outputs[5438] = (layer1_outputs[6049]) & ~(layer1_outputs[6101]);
    assign layer2_outputs[5439] = (layer1_outputs[5123]) & ~(layer1_outputs[12102]);
    assign layer2_outputs[5440] = ~((layer1_outputs[806]) ^ (layer1_outputs[2465]));
    assign layer2_outputs[5441] = layer1_outputs[10710];
    assign layer2_outputs[5442] = ~((layer1_outputs[287]) | (layer1_outputs[4948]));
    assign layer2_outputs[5443] = layer1_outputs[7180];
    assign layer2_outputs[5444] = layer1_outputs[5183];
    assign layer2_outputs[5445] = ~(layer1_outputs[6473]);
    assign layer2_outputs[5446] = (layer1_outputs[12133]) & ~(layer1_outputs[1944]);
    assign layer2_outputs[5447] = ~(layer1_outputs[2099]) | (layer1_outputs[8335]);
    assign layer2_outputs[5448] = ~(layer1_outputs[8600]);
    assign layer2_outputs[5449] = (layer1_outputs[5158]) & ~(layer1_outputs[7659]);
    assign layer2_outputs[5450] = layer1_outputs[9084];
    assign layer2_outputs[5451] = (layer1_outputs[153]) & ~(layer1_outputs[3942]);
    assign layer2_outputs[5452] = ~(layer1_outputs[4482]);
    assign layer2_outputs[5453] = layer1_outputs[2852];
    assign layer2_outputs[5454] = ~(layer1_outputs[7745]);
    assign layer2_outputs[5455] = layer1_outputs[4895];
    assign layer2_outputs[5456] = ~(layer1_outputs[4010]) | (layer1_outputs[5945]);
    assign layer2_outputs[5457] = (layer1_outputs[8620]) | (layer1_outputs[11437]);
    assign layer2_outputs[5458] = layer1_outputs[285];
    assign layer2_outputs[5459] = ~(layer1_outputs[1873]);
    assign layer2_outputs[5460] = layer1_outputs[6922];
    assign layer2_outputs[5461] = ~(layer1_outputs[5651]) | (layer1_outputs[11101]);
    assign layer2_outputs[5462] = ~(layer1_outputs[12248]);
    assign layer2_outputs[5463] = ~(layer1_outputs[1207]);
    assign layer2_outputs[5464] = (layer1_outputs[5159]) & (layer1_outputs[6245]);
    assign layer2_outputs[5465] = layer1_outputs[6865];
    assign layer2_outputs[5466] = layer1_outputs[11504];
    assign layer2_outputs[5467] = ~(layer1_outputs[11921]) | (layer1_outputs[12296]);
    assign layer2_outputs[5468] = ~((layer1_outputs[1244]) | (layer1_outputs[9718]));
    assign layer2_outputs[5469] = ~(layer1_outputs[9343]);
    assign layer2_outputs[5470] = layer1_outputs[4702];
    assign layer2_outputs[5471] = (layer1_outputs[2654]) ^ (layer1_outputs[8685]);
    assign layer2_outputs[5472] = layer1_outputs[4427];
    assign layer2_outputs[5473] = 1'b0;
    assign layer2_outputs[5474] = (layer1_outputs[12689]) & ~(layer1_outputs[11498]);
    assign layer2_outputs[5475] = ~(layer1_outputs[1769]);
    assign layer2_outputs[5476] = layer1_outputs[1119];
    assign layer2_outputs[5477] = layer1_outputs[9997];
    assign layer2_outputs[5478] = layer1_outputs[6492];
    assign layer2_outputs[5479] = ~((layer1_outputs[9629]) ^ (layer1_outputs[962]));
    assign layer2_outputs[5480] = ~(layer1_outputs[11700]) | (layer1_outputs[7752]);
    assign layer2_outputs[5481] = (layer1_outputs[5965]) | (layer1_outputs[5551]);
    assign layer2_outputs[5482] = layer1_outputs[11834];
    assign layer2_outputs[5483] = ~((layer1_outputs[8918]) & (layer1_outputs[12381]));
    assign layer2_outputs[5484] = ~(layer1_outputs[4710]) | (layer1_outputs[482]);
    assign layer2_outputs[5485] = (layer1_outputs[11249]) | (layer1_outputs[10918]);
    assign layer2_outputs[5486] = ~(layer1_outputs[10974]);
    assign layer2_outputs[5487] = ~(layer1_outputs[12285]) | (layer1_outputs[3608]);
    assign layer2_outputs[5488] = ~(layer1_outputs[8757]) | (layer1_outputs[6064]);
    assign layer2_outputs[5489] = ~((layer1_outputs[6185]) ^ (layer1_outputs[12793]));
    assign layer2_outputs[5490] = layer1_outputs[9421];
    assign layer2_outputs[5491] = (layer1_outputs[11505]) ^ (layer1_outputs[8271]);
    assign layer2_outputs[5492] = (layer1_outputs[1472]) & ~(layer1_outputs[7112]);
    assign layer2_outputs[5493] = ~(layer1_outputs[11791]);
    assign layer2_outputs[5494] = layer1_outputs[2999];
    assign layer2_outputs[5495] = layer1_outputs[11276];
    assign layer2_outputs[5496] = (layer1_outputs[4409]) ^ (layer1_outputs[5457]);
    assign layer2_outputs[5497] = layer1_outputs[2499];
    assign layer2_outputs[5498] = layer1_outputs[11081];
    assign layer2_outputs[5499] = (layer1_outputs[3023]) | (layer1_outputs[2700]);
    assign layer2_outputs[5500] = layer1_outputs[1056];
    assign layer2_outputs[5501] = ~(layer1_outputs[11575]);
    assign layer2_outputs[5502] = (layer1_outputs[2781]) | (layer1_outputs[633]);
    assign layer2_outputs[5503] = layer1_outputs[4823];
    assign layer2_outputs[5504] = (layer1_outputs[11086]) & ~(layer1_outputs[2621]);
    assign layer2_outputs[5505] = ~((layer1_outputs[8824]) ^ (layer1_outputs[4575]));
    assign layer2_outputs[5506] = ~((layer1_outputs[3254]) & (layer1_outputs[869]));
    assign layer2_outputs[5507] = (layer1_outputs[4449]) & (layer1_outputs[828]);
    assign layer2_outputs[5508] = (layer1_outputs[10525]) & (layer1_outputs[5535]);
    assign layer2_outputs[5509] = ~(layer1_outputs[9936]) | (layer1_outputs[5087]);
    assign layer2_outputs[5510] = ~((layer1_outputs[8921]) ^ (layer1_outputs[8629]));
    assign layer2_outputs[5511] = (layer1_outputs[6478]) & (layer1_outputs[6282]);
    assign layer2_outputs[5512] = (layer1_outputs[7797]) & ~(layer1_outputs[4176]);
    assign layer2_outputs[5513] = (layer1_outputs[8731]) ^ (layer1_outputs[10091]);
    assign layer2_outputs[5514] = (layer1_outputs[12604]) ^ (layer1_outputs[10972]);
    assign layer2_outputs[5515] = layer1_outputs[8823];
    assign layer2_outputs[5516] = ~(layer1_outputs[5459]);
    assign layer2_outputs[5517] = ~(layer1_outputs[1458]);
    assign layer2_outputs[5518] = layer1_outputs[5126];
    assign layer2_outputs[5519] = ~((layer1_outputs[9695]) | (layer1_outputs[11272]));
    assign layer2_outputs[5520] = layer1_outputs[9491];
    assign layer2_outputs[5521] = (layer1_outputs[11275]) ^ (layer1_outputs[1696]);
    assign layer2_outputs[5522] = ~((layer1_outputs[6193]) ^ (layer1_outputs[12362]));
    assign layer2_outputs[5523] = ~((layer1_outputs[12573]) | (layer1_outputs[12319]));
    assign layer2_outputs[5524] = ~((layer1_outputs[2600]) ^ (layer1_outputs[4222]));
    assign layer2_outputs[5525] = ~((layer1_outputs[5146]) ^ (layer1_outputs[10713]));
    assign layer2_outputs[5526] = (layer1_outputs[4688]) & (layer1_outputs[7556]);
    assign layer2_outputs[5527] = ~(layer1_outputs[311]);
    assign layer2_outputs[5528] = ~(layer1_outputs[6845]);
    assign layer2_outputs[5529] = layer1_outputs[10982];
    assign layer2_outputs[5530] = ~(layer1_outputs[4453]);
    assign layer2_outputs[5531] = ~((layer1_outputs[634]) & (layer1_outputs[11042]));
    assign layer2_outputs[5532] = layer1_outputs[785];
    assign layer2_outputs[5533] = (layer1_outputs[5624]) | (layer1_outputs[8477]);
    assign layer2_outputs[5534] = ~(layer1_outputs[9467]);
    assign layer2_outputs[5535] = (layer1_outputs[6827]) | (layer1_outputs[180]);
    assign layer2_outputs[5536] = layer1_outputs[9486];
    assign layer2_outputs[5537] = ~((layer1_outputs[207]) | (layer1_outputs[7383]));
    assign layer2_outputs[5538] = ~((layer1_outputs[10044]) | (layer1_outputs[10061]));
    assign layer2_outputs[5539] = layer1_outputs[10456];
    assign layer2_outputs[5540] = ~(layer1_outputs[11928]);
    assign layer2_outputs[5541] = (layer1_outputs[3279]) & ~(layer1_outputs[5905]);
    assign layer2_outputs[5542] = (layer1_outputs[9783]) & ~(layer1_outputs[3114]);
    assign layer2_outputs[5543] = (layer1_outputs[5695]) | (layer1_outputs[3385]);
    assign layer2_outputs[5544] = ~(layer1_outputs[9364]);
    assign layer2_outputs[5545] = ~(layer1_outputs[9960]);
    assign layer2_outputs[5546] = ~(layer1_outputs[5599]);
    assign layer2_outputs[5547] = ~(layer1_outputs[10901]);
    assign layer2_outputs[5548] = ~((layer1_outputs[2956]) ^ (layer1_outputs[4855]));
    assign layer2_outputs[5549] = ~((layer1_outputs[8785]) | (layer1_outputs[11717]));
    assign layer2_outputs[5550] = ~((layer1_outputs[9593]) & (layer1_outputs[8135]));
    assign layer2_outputs[5551] = ~(layer1_outputs[6268]);
    assign layer2_outputs[5552] = layer1_outputs[8319];
    assign layer2_outputs[5553] = (layer1_outputs[2326]) ^ (layer1_outputs[12208]);
    assign layer2_outputs[5554] = ~(layer1_outputs[9855]);
    assign layer2_outputs[5555] = ~(layer1_outputs[2167]);
    assign layer2_outputs[5556] = layer1_outputs[5460];
    assign layer2_outputs[5557] = ~(layer1_outputs[7075]);
    assign layer2_outputs[5558] = layer1_outputs[6562];
    assign layer2_outputs[5559] = ~((layer1_outputs[6657]) ^ (layer1_outputs[4354]));
    assign layer2_outputs[5560] = (layer1_outputs[6158]) & (layer1_outputs[4698]);
    assign layer2_outputs[5561] = (layer1_outputs[192]) | (layer1_outputs[3229]);
    assign layer2_outputs[5562] = layer1_outputs[10675];
    assign layer2_outputs[5563] = layer1_outputs[292];
    assign layer2_outputs[5564] = layer1_outputs[11953];
    assign layer2_outputs[5565] = layer1_outputs[11640];
    assign layer2_outputs[5566] = (layer1_outputs[1649]) ^ (layer1_outputs[10668]);
    assign layer2_outputs[5567] = (layer1_outputs[12786]) & ~(layer1_outputs[12755]);
    assign layer2_outputs[5568] = ~(layer1_outputs[4848]);
    assign layer2_outputs[5569] = ~(layer1_outputs[10092]);
    assign layer2_outputs[5570] = ~(layer1_outputs[6168]);
    assign layer2_outputs[5571] = layer1_outputs[1256];
    assign layer2_outputs[5572] = (layer1_outputs[3369]) ^ (layer1_outputs[1345]);
    assign layer2_outputs[5573] = layer1_outputs[8879];
    assign layer2_outputs[5574] = layer1_outputs[12203];
    assign layer2_outputs[5575] = layer1_outputs[1208];
    assign layer2_outputs[5576] = ~(layer1_outputs[5570]);
    assign layer2_outputs[5577] = layer1_outputs[5884];
    assign layer2_outputs[5578] = ~(layer1_outputs[3963]);
    assign layer2_outputs[5579] = ~(layer1_outputs[3923]) | (layer1_outputs[8290]);
    assign layer2_outputs[5580] = ~((layer1_outputs[6687]) & (layer1_outputs[1849]));
    assign layer2_outputs[5581] = layer1_outputs[5540];
    assign layer2_outputs[5582] = layer1_outputs[3712];
    assign layer2_outputs[5583] = layer1_outputs[7685];
    assign layer2_outputs[5584] = (layer1_outputs[11093]) ^ (layer1_outputs[3246]);
    assign layer2_outputs[5585] = ~(layer1_outputs[11569]);
    assign layer2_outputs[5586] = layer1_outputs[263];
    assign layer2_outputs[5587] = ~((layer1_outputs[3194]) ^ (layer1_outputs[7675]));
    assign layer2_outputs[5588] = (layer1_outputs[10845]) ^ (layer1_outputs[515]);
    assign layer2_outputs[5589] = ~(layer1_outputs[10791]);
    assign layer2_outputs[5590] = (layer1_outputs[10168]) & ~(layer1_outputs[11009]);
    assign layer2_outputs[5591] = (layer1_outputs[10886]) ^ (layer1_outputs[1730]);
    assign layer2_outputs[5592] = ~((layer1_outputs[1751]) ^ (layer1_outputs[9503]));
    assign layer2_outputs[5593] = ~(layer1_outputs[717]);
    assign layer2_outputs[5594] = ~((layer1_outputs[5020]) & (layer1_outputs[5833]));
    assign layer2_outputs[5595] = (layer1_outputs[10305]) | (layer1_outputs[6782]);
    assign layer2_outputs[5596] = ~(layer1_outputs[2843]);
    assign layer2_outputs[5597] = ~(layer1_outputs[11241]);
    assign layer2_outputs[5598] = ~(layer1_outputs[6790]) | (layer1_outputs[31]);
    assign layer2_outputs[5599] = ~(layer1_outputs[4614]);
    assign layer2_outputs[5600] = layer1_outputs[9258];
    assign layer2_outputs[5601] = ~(layer1_outputs[1207]);
    assign layer2_outputs[5602] = layer1_outputs[12667];
    assign layer2_outputs[5603] = ~(layer1_outputs[533]);
    assign layer2_outputs[5604] = layer1_outputs[12757];
    assign layer2_outputs[5605] = ~(layer1_outputs[6840]);
    assign layer2_outputs[5606] = ~(layer1_outputs[8089]);
    assign layer2_outputs[5607] = (layer1_outputs[103]) & ~(layer1_outputs[5988]);
    assign layer2_outputs[5608] = layer1_outputs[9160];
    assign layer2_outputs[5609] = (layer1_outputs[5866]) ^ (layer1_outputs[7755]);
    assign layer2_outputs[5610] = layer1_outputs[2938];
    assign layer2_outputs[5611] = (layer1_outputs[8290]) & ~(layer1_outputs[228]);
    assign layer2_outputs[5612] = ~(layer1_outputs[2841]);
    assign layer2_outputs[5613] = ~(layer1_outputs[4000]);
    assign layer2_outputs[5614] = layer1_outputs[12041];
    assign layer2_outputs[5615] = (layer1_outputs[5822]) | (layer1_outputs[2153]);
    assign layer2_outputs[5616] = ~((layer1_outputs[12242]) ^ (layer1_outputs[10773]));
    assign layer2_outputs[5617] = ~(layer1_outputs[11269]);
    assign layer2_outputs[5618] = ~(layer1_outputs[8618]);
    assign layer2_outputs[5619] = (layer1_outputs[11446]) & ~(layer1_outputs[8967]);
    assign layer2_outputs[5620] = ~((layer1_outputs[3498]) | (layer1_outputs[5033]));
    assign layer2_outputs[5621] = ~(layer1_outputs[2756]);
    assign layer2_outputs[5622] = ~(layer1_outputs[5119]);
    assign layer2_outputs[5623] = ~((layer1_outputs[4013]) & (layer1_outputs[6992]));
    assign layer2_outputs[5624] = layer1_outputs[11805];
    assign layer2_outputs[5625] = ~(layer1_outputs[10782]);
    assign layer2_outputs[5626] = ~(layer1_outputs[11800]);
    assign layer2_outputs[5627] = (layer1_outputs[6019]) & ~(layer1_outputs[1183]);
    assign layer2_outputs[5628] = ~(layer1_outputs[866]);
    assign layer2_outputs[5629] = ~(layer1_outputs[9825]) | (layer1_outputs[4171]);
    assign layer2_outputs[5630] = (layer1_outputs[10143]) & ~(layer1_outputs[2249]);
    assign layer2_outputs[5631] = ~(layer1_outputs[10023]);
    assign layer2_outputs[5632] = layer1_outputs[10732];
    assign layer2_outputs[5633] = layer1_outputs[8676];
    assign layer2_outputs[5634] = (layer1_outputs[7980]) & ~(layer1_outputs[12194]);
    assign layer2_outputs[5635] = ~((layer1_outputs[6925]) & (layer1_outputs[319]));
    assign layer2_outputs[5636] = layer1_outputs[8903];
    assign layer2_outputs[5637] = (layer1_outputs[4478]) | (layer1_outputs[8384]);
    assign layer2_outputs[5638] = ~(layer1_outputs[10393]);
    assign layer2_outputs[5639] = ~(layer1_outputs[3233]);
    assign layer2_outputs[5640] = ~(layer1_outputs[7896]);
    assign layer2_outputs[5641] = ~(layer1_outputs[5487]);
    assign layer2_outputs[5642] = ~(layer1_outputs[1759]);
    assign layer2_outputs[5643] = ~(layer1_outputs[8352]);
    assign layer2_outputs[5644] = (layer1_outputs[7364]) ^ (layer1_outputs[7826]);
    assign layer2_outputs[5645] = ~(layer1_outputs[9225]);
    assign layer2_outputs[5646] = ~(layer1_outputs[5678]);
    assign layer2_outputs[5647] = ~(layer1_outputs[2067]);
    assign layer2_outputs[5648] = ~(layer1_outputs[2939]);
    assign layer2_outputs[5649] = layer1_outputs[11904];
    assign layer2_outputs[5650] = ~((layer1_outputs[5282]) & (layer1_outputs[8342]));
    assign layer2_outputs[5651] = ~((layer1_outputs[10241]) | (layer1_outputs[3801]));
    assign layer2_outputs[5652] = ~(layer1_outputs[7646]);
    assign layer2_outputs[5653] = (layer1_outputs[6876]) | (layer1_outputs[11416]);
    assign layer2_outputs[5654] = (layer1_outputs[3945]) ^ (layer1_outputs[8932]);
    assign layer2_outputs[5655] = layer1_outputs[3008];
    assign layer2_outputs[5656] = ~((layer1_outputs[7253]) ^ (layer1_outputs[8416]));
    assign layer2_outputs[5657] = (layer1_outputs[9647]) ^ (layer1_outputs[3397]);
    assign layer2_outputs[5658] = ~(layer1_outputs[1497]);
    assign layer2_outputs[5659] = layer1_outputs[10046];
    assign layer2_outputs[5660] = ~(layer1_outputs[3630]);
    assign layer2_outputs[5661] = (layer1_outputs[2425]) & (layer1_outputs[3240]);
    assign layer2_outputs[5662] = ~((layer1_outputs[1676]) | (layer1_outputs[284]));
    assign layer2_outputs[5663] = ~(layer1_outputs[6795]);
    assign layer2_outputs[5664] = ~((layer1_outputs[9632]) & (layer1_outputs[4447]));
    assign layer2_outputs[5665] = layer1_outputs[4378];
    assign layer2_outputs[5666] = ~(layer1_outputs[3170]);
    assign layer2_outputs[5667] = (layer1_outputs[1271]) & (layer1_outputs[3774]);
    assign layer2_outputs[5668] = layer1_outputs[3988];
    assign layer2_outputs[5669] = (layer1_outputs[5417]) & ~(layer1_outputs[3813]);
    assign layer2_outputs[5670] = layer1_outputs[7729];
    assign layer2_outputs[5671] = ~(layer1_outputs[7716]);
    assign layer2_outputs[5672] = ~((layer1_outputs[11801]) ^ (layer1_outputs[899]));
    assign layer2_outputs[5673] = (layer1_outputs[8805]) & ~(layer1_outputs[1020]);
    assign layer2_outputs[5674] = layer1_outputs[11864];
    assign layer2_outputs[5675] = ~((layer1_outputs[1585]) ^ (layer1_outputs[2004]));
    assign layer2_outputs[5676] = ~(layer1_outputs[39]) | (layer1_outputs[4080]);
    assign layer2_outputs[5677] = (layer1_outputs[4230]) | (layer1_outputs[1631]);
    assign layer2_outputs[5678] = layer1_outputs[8080];
    assign layer2_outputs[5679] = ~(layer1_outputs[12179]);
    assign layer2_outputs[5680] = layer1_outputs[4868];
    assign layer2_outputs[5681] = layer1_outputs[8142];
    assign layer2_outputs[5682] = ~((layer1_outputs[7358]) ^ (layer1_outputs[8091]));
    assign layer2_outputs[5683] = ~((layer1_outputs[10227]) ^ (layer1_outputs[350]));
    assign layer2_outputs[5684] = ~(layer1_outputs[5757]);
    assign layer2_outputs[5685] = ~(layer1_outputs[12431]) | (layer1_outputs[7889]);
    assign layer2_outputs[5686] = ~(layer1_outputs[7618]);
    assign layer2_outputs[5687] = ~((layer1_outputs[862]) & (layer1_outputs[7201]));
    assign layer2_outputs[5688] = (layer1_outputs[9530]) & ~(layer1_outputs[8282]);
    assign layer2_outputs[5689] = (layer1_outputs[7954]) & ~(layer1_outputs[12622]);
    assign layer2_outputs[5690] = ~(layer1_outputs[10327]);
    assign layer2_outputs[5691] = layer1_outputs[11346];
    assign layer2_outputs[5692] = ~(layer1_outputs[3972]);
    assign layer2_outputs[5693] = (layer1_outputs[9311]) ^ (layer1_outputs[8083]);
    assign layer2_outputs[5694] = layer1_outputs[11667];
    assign layer2_outputs[5695] = ~(layer1_outputs[8259]);
    assign layer2_outputs[5696] = ~(layer1_outputs[4585]);
    assign layer2_outputs[5697] = (layer1_outputs[9922]) | (layer1_outputs[3632]);
    assign layer2_outputs[5698] = (layer1_outputs[11379]) | (layer1_outputs[8994]);
    assign layer2_outputs[5699] = ~(layer1_outputs[6690]);
    assign layer2_outputs[5700] = ~((layer1_outputs[8487]) | (layer1_outputs[7015]));
    assign layer2_outputs[5701] = ~(layer1_outputs[8378]);
    assign layer2_outputs[5702] = (layer1_outputs[12046]) & ~(layer1_outputs[1636]);
    assign layer2_outputs[5703] = ~(layer1_outputs[9027]);
    assign layer2_outputs[5704] = ~(layer1_outputs[9814]);
    assign layer2_outputs[5705] = ~((layer1_outputs[8585]) ^ (layer1_outputs[9364]));
    assign layer2_outputs[5706] = layer1_outputs[358];
    assign layer2_outputs[5707] = ~((layer1_outputs[486]) & (layer1_outputs[3091]));
    assign layer2_outputs[5708] = ~(layer1_outputs[9197]);
    assign layer2_outputs[5709] = layer1_outputs[7681];
    assign layer2_outputs[5710] = (layer1_outputs[700]) ^ (layer1_outputs[9408]);
    assign layer2_outputs[5711] = (layer1_outputs[12262]) & (layer1_outputs[12281]);
    assign layer2_outputs[5712] = layer1_outputs[183];
    assign layer2_outputs[5713] = (layer1_outputs[8440]) & (layer1_outputs[8468]);
    assign layer2_outputs[5714] = (layer1_outputs[2414]) & ~(layer1_outputs[8207]);
    assign layer2_outputs[5715] = (layer1_outputs[3371]) ^ (layer1_outputs[7796]);
    assign layer2_outputs[5716] = (layer1_outputs[9055]) & ~(layer1_outputs[6850]);
    assign layer2_outputs[5717] = ~(layer1_outputs[1545]) | (layer1_outputs[4686]);
    assign layer2_outputs[5718] = ~(layer1_outputs[2140]);
    assign layer2_outputs[5719] = layer1_outputs[8030];
    assign layer2_outputs[5720] = ~(layer1_outputs[2091]);
    assign layer2_outputs[5721] = (layer1_outputs[8456]) & ~(layer1_outputs[1151]);
    assign layer2_outputs[5722] = ~(layer1_outputs[4179]);
    assign layer2_outputs[5723] = ~((layer1_outputs[4176]) & (layer1_outputs[3809]));
    assign layer2_outputs[5724] = layer1_outputs[11833];
    assign layer2_outputs[5725] = ~((layer1_outputs[8233]) & (layer1_outputs[6784]));
    assign layer2_outputs[5726] = ~((layer1_outputs[7240]) & (layer1_outputs[3007]));
    assign layer2_outputs[5727] = ~((layer1_outputs[3382]) ^ (layer1_outputs[6720]));
    assign layer2_outputs[5728] = layer1_outputs[6819];
    assign layer2_outputs[5729] = (layer1_outputs[5532]) | (layer1_outputs[8140]);
    assign layer2_outputs[5730] = layer1_outputs[2811];
    assign layer2_outputs[5731] = (layer1_outputs[6109]) ^ (layer1_outputs[9898]);
    assign layer2_outputs[5732] = ~(layer1_outputs[10841]);
    assign layer2_outputs[5733] = (layer1_outputs[164]) | (layer1_outputs[11187]);
    assign layer2_outputs[5734] = ~((layer1_outputs[7159]) | (layer1_outputs[7201]));
    assign layer2_outputs[5735] = layer1_outputs[7971];
    assign layer2_outputs[5736] = ~(layer1_outputs[7288]);
    assign layer2_outputs[5737] = ~(layer1_outputs[8483]) | (layer1_outputs[2020]);
    assign layer2_outputs[5738] = layer1_outputs[6942];
    assign layer2_outputs[5739] = ~(layer1_outputs[3440]);
    assign layer2_outputs[5740] = ~(layer1_outputs[10677]) | (layer1_outputs[1909]);
    assign layer2_outputs[5741] = ~(layer1_outputs[6803]);
    assign layer2_outputs[5742] = ~(layer1_outputs[1105]);
    assign layer2_outputs[5743] = ~(layer1_outputs[11095]) | (layer1_outputs[7531]);
    assign layer2_outputs[5744] = layer1_outputs[9853];
    assign layer2_outputs[5745] = ~(layer1_outputs[3122]);
    assign layer2_outputs[5746] = ~(layer1_outputs[8662]);
    assign layer2_outputs[5747] = ~((layer1_outputs[4216]) & (layer1_outputs[329]));
    assign layer2_outputs[5748] = ~(layer1_outputs[10716]) | (layer1_outputs[12257]);
    assign layer2_outputs[5749] = ~((layer1_outputs[10156]) | (layer1_outputs[7703]));
    assign layer2_outputs[5750] = (layer1_outputs[3298]) & (layer1_outputs[5770]);
    assign layer2_outputs[5751] = layer1_outputs[3304];
    assign layer2_outputs[5752] = ~((layer1_outputs[2736]) & (layer1_outputs[2149]));
    assign layer2_outputs[5753] = layer1_outputs[11624];
    assign layer2_outputs[5754] = layer1_outputs[4809];
    assign layer2_outputs[5755] = ~(layer1_outputs[1951]) | (layer1_outputs[10670]);
    assign layer2_outputs[5756] = layer1_outputs[5122];
    assign layer2_outputs[5757] = layer1_outputs[10236];
    assign layer2_outputs[5758] = ~(layer1_outputs[3017]);
    assign layer2_outputs[5759] = layer1_outputs[4464];
    assign layer2_outputs[5760] = ~((layer1_outputs[8123]) | (layer1_outputs[9384]));
    assign layer2_outputs[5761] = (layer1_outputs[9491]) ^ (layer1_outputs[10334]);
    assign layer2_outputs[5762] = layer1_outputs[8323];
    assign layer2_outputs[5763] = (layer1_outputs[6624]) & ~(layer1_outputs[6281]);
    assign layer2_outputs[5764] = ~(layer1_outputs[541]);
    assign layer2_outputs[5765] = ~(layer1_outputs[4335]);
    assign layer2_outputs[5766] = (layer1_outputs[4215]) ^ (layer1_outputs[2507]);
    assign layer2_outputs[5767] = layer1_outputs[239];
    assign layer2_outputs[5768] = ~((layer1_outputs[6534]) ^ (layer1_outputs[10144]));
    assign layer2_outputs[5769] = (layer1_outputs[7912]) ^ (layer1_outputs[5977]);
    assign layer2_outputs[5770] = (layer1_outputs[2549]) & ~(layer1_outputs[11020]);
    assign layer2_outputs[5771] = ~(layer1_outputs[3328]);
    assign layer2_outputs[5772] = ~(layer1_outputs[7614]);
    assign layer2_outputs[5773] = layer1_outputs[11403];
    assign layer2_outputs[5774] = (layer1_outputs[7605]) | (layer1_outputs[2276]);
    assign layer2_outputs[5775] = ~(layer1_outputs[20]);
    assign layer2_outputs[5776] = ~(layer1_outputs[9397]);
    assign layer2_outputs[5777] = layer1_outputs[4708];
    assign layer2_outputs[5778] = ~(layer1_outputs[2578]);
    assign layer2_outputs[5779] = ~(layer1_outputs[9776]);
    assign layer2_outputs[5780] = ~((layer1_outputs[1022]) & (layer1_outputs[5782]));
    assign layer2_outputs[5781] = layer1_outputs[8830];
    assign layer2_outputs[5782] = ~((layer1_outputs[4194]) ^ (layer1_outputs[1130]));
    assign layer2_outputs[5783] = ~(layer1_outputs[8790]);
    assign layer2_outputs[5784] = ~(layer1_outputs[4796]);
    assign layer2_outputs[5785] = layer1_outputs[8774];
    assign layer2_outputs[5786] = 1'b0;
    assign layer2_outputs[5787] = ~((layer1_outputs[4030]) ^ (layer1_outputs[1057]));
    assign layer2_outputs[5788] = (layer1_outputs[679]) & (layer1_outputs[8816]);
    assign layer2_outputs[5789] = (layer1_outputs[613]) & (layer1_outputs[9385]);
    assign layer2_outputs[5790] = ~(layer1_outputs[3582]);
    assign layer2_outputs[5791] = layer1_outputs[8601];
    assign layer2_outputs[5792] = (layer1_outputs[2662]) & (layer1_outputs[11989]);
    assign layer2_outputs[5793] = (layer1_outputs[6980]) & (layer1_outputs[975]);
    assign layer2_outputs[5794] = (layer1_outputs[9159]) ^ (layer1_outputs[1633]);
    assign layer2_outputs[5795] = ~((layer1_outputs[11568]) ^ (layer1_outputs[11158]));
    assign layer2_outputs[5796] = layer1_outputs[12410];
    assign layer2_outputs[5797] = ~((layer1_outputs[11344]) & (layer1_outputs[11352]));
    assign layer2_outputs[5798] = layer1_outputs[2982];
    assign layer2_outputs[5799] = ~(layer1_outputs[10983]) | (layer1_outputs[6300]);
    assign layer2_outputs[5800] = (layer1_outputs[3276]) & ~(layer1_outputs[8350]);
    assign layer2_outputs[5801] = ~(layer1_outputs[5534]);
    assign layer2_outputs[5802] = layer1_outputs[12564];
    assign layer2_outputs[5803] = ~(layer1_outputs[10124]) | (layer1_outputs[10320]);
    assign layer2_outputs[5804] = ~(layer1_outputs[4819]);
    assign layer2_outputs[5805] = ~((layer1_outputs[7356]) ^ (layer1_outputs[4379]));
    assign layer2_outputs[5806] = ~(layer1_outputs[2139]);
    assign layer2_outputs[5807] = ~(layer1_outputs[4340]);
    assign layer2_outputs[5808] = layer1_outputs[7448];
    assign layer2_outputs[5809] = ~(layer1_outputs[9655]);
    assign layer2_outputs[5810] = ~(layer1_outputs[5542]);
    assign layer2_outputs[5811] = (layer1_outputs[5971]) ^ (layer1_outputs[6744]);
    assign layer2_outputs[5812] = ~((layer1_outputs[7412]) & (layer1_outputs[8098]));
    assign layer2_outputs[5813] = ~(layer1_outputs[10473]) | (layer1_outputs[3795]);
    assign layer2_outputs[5814] = ~(layer1_outputs[2137]);
    assign layer2_outputs[5815] = layer1_outputs[4315];
    assign layer2_outputs[5816] = ~(layer1_outputs[1641]);
    assign layer2_outputs[5817] = (layer1_outputs[12528]) ^ (layer1_outputs[4131]);
    assign layer2_outputs[5818] = (layer1_outputs[2513]) & (layer1_outputs[1384]);
    assign layer2_outputs[5819] = (layer1_outputs[7406]) ^ (layer1_outputs[11353]);
    assign layer2_outputs[5820] = ~(layer1_outputs[11097]) | (layer1_outputs[10343]);
    assign layer2_outputs[5821] = (layer1_outputs[2187]) & ~(layer1_outputs[1120]);
    assign layer2_outputs[5822] = (layer1_outputs[4557]) | (layer1_outputs[11538]);
    assign layer2_outputs[5823] = (layer1_outputs[5868]) & ~(layer1_outputs[3841]);
    assign layer2_outputs[5824] = ~((layer1_outputs[11920]) | (layer1_outputs[2932]));
    assign layer2_outputs[5825] = layer1_outputs[5468];
    assign layer2_outputs[5826] = ~(layer1_outputs[11767]) | (layer1_outputs[6559]);
    assign layer2_outputs[5827] = ~(layer1_outputs[3794]) | (layer1_outputs[4654]);
    assign layer2_outputs[5828] = ~(layer1_outputs[7304]) | (layer1_outputs[9451]);
    assign layer2_outputs[5829] = layer1_outputs[10982];
    assign layer2_outputs[5830] = (layer1_outputs[7990]) & ~(layer1_outputs[5273]);
    assign layer2_outputs[5831] = (layer1_outputs[12224]) ^ (layer1_outputs[5645]);
    assign layer2_outputs[5832] = (layer1_outputs[1108]) ^ (layer1_outputs[7471]);
    assign layer2_outputs[5833] = layer1_outputs[12722];
    assign layer2_outputs[5834] = ~(layer1_outputs[7617]);
    assign layer2_outputs[5835] = layer1_outputs[12321];
    assign layer2_outputs[5836] = ~(layer1_outputs[4837]);
    assign layer2_outputs[5837] = (layer1_outputs[5593]) & ~(layer1_outputs[3202]);
    assign layer2_outputs[5838] = ~(layer1_outputs[4567]);
    assign layer2_outputs[5839] = ~(layer1_outputs[11557]);
    assign layer2_outputs[5840] = ~(layer1_outputs[8046]);
    assign layer2_outputs[5841] = (layer1_outputs[8371]) ^ (layer1_outputs[3536]);
    assign layer2_outputs[5842] = (layer1_outputs[2063]) & ~(layer1_outputs[8504]);
    assign layer2_outputs[5843] = ~(layer1_outputs[12538]);
    assign layer2_outputs[5844] = layer1_outputs[6427];
    assign layer2_outputs[5845] = layer1_outputs[480];
    assign layer2_outputs[5846] = ~((layer1_outputs[5184]) & (layer1_outputs[10890]));
    assign layer2_outputs[5847] = ~(layer1_outputs[2367]);
    assign layer2_outputs[5848] = layer1_outputs[3207];
    assign layer2_outputs[5849] = ~(layer1_outputs[10795]);
    assign layer2_outputs[5850] = layer1_outputs[10443];
    assign layer2_outputs[5851] = ~((layer1_outputs[11983]) ^ (layer1_outputs[1200]));
    assign layer2_outputs[5852] = layer1_outputs[1291];
    assign layer2_outputs[5853] = layer1_outputs[7208];
    assign layer2_outputs[5854] = (layer1_outputs[7376]) & (layer1_outputs[1547]);
    assign layer2_outputs[5855] = ~(layer1_outputs[6809]) | (layer1_outputs[4107]);
    assign layer2_outputs[5856] = (layer1_outputs[1950]) & ~(layer1_outputs[921]);
    assign layer2_outputs[5857] = ~((layer1_outputs[10674]) & (layer1_outputs[12157]));
    assign layer2_outputs[5858] = (layer1_outputs[7071]) & ~(layer1_outputs[7311]);
    assign layer2_outputs[5859] = (layer1_outputs[10749]) ^ (layer1_outputs[4013]);
    assign layer2_outputs[5860] = ~(layer1_outputs[5682]) | (layer1_outputs[3216]);
    assign layer2_outputs[5861] = (layer1_outputs[2738]) | (layer1_outputs[5574]);
    assign layer2_outputs[5862] = ~((layer1_outputs[3434]) ^ (layer1_outputs[4906]));
    assign layer2_outputs[5863] = layer1_outputs[2059];
    assign layer2_outputs[5864] = layer1_outputs[2648];
    assign layer2_outputs[5865] = (layer1_outputs[1091]) | (layer1_outputs[2166]);
    assign layer2_outputs[5866] = ~((layer1_outputs[12684]) ^ (layer1_outputs[2573]));
    assign layer2_outputs[5867] = ~(layer1_outputs[12739]) | (layer1_outputs[4307]);
    assign layer2_outputs[5868] = ~((layer1_outputs[1767]) | (layer1_outputs[4623]));
    assign layer2_outputs[5869] = ~((layer1_outputs[4595]) ^ (layer1_outputs[12452]));
    assign layer2_outputs[5870] = layer1_outputs[3157];
    assign layer2_outputs[5871] = ~(layer1_outputs[5380]);
    assign layer2_outputs[5872] = ~((layer1_outputs[10517]) & (layer1_outputs[12003]));
    assign layer2_outputs[5873] = ~(layer1_outputs[5350]);
    assign layer2_outputs[5874] = ~(layer1_outputs[9245]);
    assign layer2_outputs[5875] = ~(layer1_outputs[4583]);
    assign layer2_outputs[5876] = ~(layer1_outputs[7098]);
    assign layer2_outputs[5877] = ~(layer1_outputs[9166]) | (layer1_outputs[1884]);
    assign layer2_outputs[5878] = ~(layer1_outputs[11011]);
    assign layer2_outputs[5879] = ~((layer1_outputs[6925]) | (layer1_outputs[6474]));
    assign layer2_outputs[5880] = layer1_outputs[8973];
    assign layer2_outputs[5881] = layer1_outputs[1076];
    assign layer2_outputs[5882] = ~(layer1_outputs[3402]);
    assign layer2_outputs[5883] = layer1_outputs[2383];
    assign layer2_outputs[5884] = layer1_outputs[1727];
    assign layer2_outputs[5885] = ~((layer1_outputs[10345]) ^ (layer1_outputs[6824]));
    assign layer2_outputs[5886] = layer1_outputs[12551];
    assign layer2_outputs[5887] = (layer1_outputs[8307]) & ~(layer1_outputs[1837]);
    assign layer2_outputs[5888] = (layer1_outputs[5324]) ^ (layer1_outputs[68]);
    assign layer2_outputs[5889] = layer1_outputs[8464];
    assign layer2_outputs[5890] = ~((layer1_outputs[7109]) ^ (layer1_outputs[4058]));
    assign layer2_outputs[5891] = (layer1_outputs[10105]) | (layer1_outputs[3047]);
    assign layer2_outputs[5892] = ~(layer1_outputs[8792]);
    assign layer2_outputs[5893] = layer1_outputs[354];
    assign layer2_outputs[5894] = ~(layer1_outputs[7738]) | (layer1_outputs[11700]);
    assign layer2_outputs[5895] = layer1_outputs[2356];
    assign layer2_outputs[5896] = ~((layer1_outputs[3981]) ^ (layer1_outputs[3929]));
    assign layer2_outputs[5897] = (layer1_outputs[10589]) ^ (layer1_outputs[6537]);
    assign layer2_outputs[5898] = layer1_outputs[6858];
    assign layer2_outputs[5899] = (layer1_outputs[338]) ^ (layer1_outputs[3930]);
    assign layer2_outputs[5900] = ~(layer1_outputs[7680]);
    assign layer2_outputs[5901] = layer1_outputs[4140];
    assign layer2_outputs[5902] = ~(layer1_outputs[1856]);
    assign layer2_outputs[5903] = layer1_outputs[11233];
    assign layer2_outputs[5904] = layer1_outputs[11027];
    assign layer2_outputs[5905] = ~(layer1_outputs[5231]);
    assign layer2_outputs[5906] = 1'b1;
    assign layer2_outputs[5907] = layer1_outputs[11478];
    assign layer2_outputs[5908] = ~(layer1_outputs[4251]);
    assign layer2_outputs[5909] = ~((layer1_outputs[1386]) ^ (layer1_outputs[5387]));
    assign layer2_outputs[5910] = ~(layer1_outputs[987]) | (layer1_outputs[5152]);
    assign layer2_outputs[5911] = layer1_outputs[8496];
    assign layer2_outputs[5912] = layer1_outputs[6806];
    assign layer2_outputs[5913] = ~(layer1_outputs[4469]);
    assign layer2_outputs[5914] = ~(layer1_outputs[9484]);
    assign layer2_outputs[5915] = (layer1_outputs[4859]) & (layer1_outputs[11086]);
    assign layer2_outputs[5916] = ~(layer1_outputs[1322]) | (layer1_outputs[7613]);
    assign layer2_outputs[5917] = ~((layer1_outputs[522]) & (layer1_outputs[2033]));
    assign layer2_outputs[5918] = layer1_outputs[9497];
    assign layer2_outputs[5919] = layer1_outputs[11214];
    assign layer2_outputs[5920] = (layer1_outputs[7147]) | (layer1_outputs[9297]);
    assign layer2_outputs[5921] = ~(layer1_outputs[9051]);
    assign layer2_outputs[5922] = ~(layer1_outputs[7069]);
    assign layer2_outputs[5923] = (layer1_outputs[10273]) ^ (layer1_outputs[12438]);
    assign layer2_outputs[5924] = (layer1_outputs[952]) ^ (layer1_outputs[7875]);
    assign layer2_outputs[5925] = layer1_outputs[11807];
    assign layer2_outputs[5926] = ~(layer1_outputs[1438]);
    assign layer2_outputs[5927] = layer1_outputs[6195];
    assign layer2_outputs[5928] = ~(layer1_outputs[228]);
    assign layer2_outputs[5929] = ~((layer1_outputs[8862]) ^ (layer1_outputs[2220]));
    assign layer2_outputs[5930] = layer1_outputs[11816];
    assign layer2_outputs[5931] = ~((layer1_outputs[7421]) ^ (layer1_outputs[2711]));
    assign layer2_outputs[5932] = layer1_outputs[2789];
    assign layer2_outputs[5933] = ~((layer1_outputs[4045]) ^ (layer1_outputs[10147]));
    assign layer2_outputs[5934] = layer1_outputs[485];
    assign layer2_outputs[5935] = layer1_outputs[12719];
    assign layer2_outputs[5936] = ~((layer1_outputs[7671]) ^ (layer1_outputs[9821]));
    assign layer2_outputs[5937] = ~((layer1_outputs[11773]) | (layer1_outputs[120]));
    assign layer2_outputs[5938] = (layer1_outputs[11398]) & ~(layer1_outputs[8549]);
    assign layer2_outputs[5939] = layer1_outputs[11882];
    assign layer2_outputs[5940] = ~(layer1_outputs[11827]) | (layer1_outputs[2088]);
    assign layer2_outputs[5941] = ~(layer1_outputs[11317]);
    assign layer2_outputs[5942] = (layer1_outputs[6166]) ^ (layer1_outputs[3626]);
    assign layer2_outputs[5943] = layer1_outputs[6659];
    assign layer2_outputs[5944] = ~(layer1_outputs[4312]);
    assign layer2_outputs[5945] = layer1_outputs[885];
    assign layer2_outputs[5946] = layer1_outputs[825];
    assign layer2_outputs[5947] = ~((layer1_outputs[12729]) ^ (layer1_outputs[1636]));
    assign layer2_outputs[5948] = ~((layer1_outputs[695]) | (layer1_outputs[8488]));
    assign layer2_outputs[5949] = layer1_outputs[3686];
    assign layer2_outputs[5950] = ~((layer1_outputs[1534]) | (layer1_outputs[11584]));
    assign layer2_outputs[5951] = layer1_outputs[3342];
    assign layer2_outputs[5952] = (layer1_outputs[11895]) & (layer1_outputs[9666]);
    assign layer2_outputs[5953] = ~(layer1_outputs[12239]);
    assign layer2_outputs[5954] = (layer1_outputs[427]) & ~(layer1_outputs[7318]);
    assign layer2_outputs[5955] = ~(layer1_outputs[3341]);
    assign layer2_outputs[5956] = ~(layer1_outputs[3683]) | (layer1_outputs[12731]);
    assign layer2_outputs[5957] = ~(layer1_outputs[9238]) | (layer1_outputs[3140]);
    assign layer2_outputs[5958] = layer1_outputs[38];
    assign layer2_outputs[5959] = layer1_outputs[2604];
    assign layer2_outputs[5960] = ~(layer1_outputs[8292]);
    assign layer2_outputs[5961] = ~(layer1_outputs[12405]);
    assign layer2_outputs[5962] = ~(layer1_outputs[3301]) | (layer1_outputs[4133]);
    assign layer2_outputs[5963] = ~(layer1_outputs[9100]);
    assign layer2_outputs[5964] = ~(layer1_outputs[6172]) | (layer1_outputs[8152]);
    assign layer2_outputs[5965] = ~((layer1_outputs[3141]) ^ (layer1_outputs[628]));
    assign layer2_outputs[5966] = ~(layer1_outputs[12023]) | (layer1_outputs[8217]);
    assign layer2_outputs[5967] = layer1_outputs[7769];
    assign layer2_outputs[5968] = (layer1_outputs[7156]) & ~(layer1_outputs[10806]);
    assign layer2_outputs[5969] = (layer1_outputs[11669]) & (layer1_outputs[2990]);
    assign layer2_outputs[5970] = ~(layer1_outputs[11696]);
    assign layer2_outputs[5971] = layer1_outputs[2190];
    assign layer2_outputs[5972] = ~(layer1_outputs[1505]);
    assign layer2_outputs[5973] = layer1_outputs[1770];
    assign layer2_outputs[5974] = layer1_outputs[9754];
    assign layer2_outputs[5975] = (layer1_outputs[6105]) & (layer1_outputs[12673]);
    assign layer2_outputs[5976] = ~(layer1_outputs[8974]);
    assign layer2_outputs[5977] = ~(layer1_outputs[3824]);
    assign layer2_outputs[5978] = ~(layer1_outputs[9798]);
    assign layer2_outputs[5979] = ~(layer1_outputs[11713]) | (layer1_outputs[11895]);
    assign layer2_outputs[5980] = ~((layer1_outputs[3525]) & (layer1_outputs[10810]));
    assign layer2_outputs[5981] = (layer1_outputs[3765]) & ~(layer1_outputs[5221]);
    assign layer2_outputs[5982] = ~(layer1_outputs[799]);
    assign layer2_outputs[5983] = ~((layer1_outputs[11169]) | (layer1_outputs[607]));
    assign layer2_outputs[5984] = ~(layer1_outputs[9091]);
    assign layer2_outputs[5985] = (layer1_outputs[2881]) & (layer1_outputs[2736]);
    assign layer2_outputs[5986] = (layer1_outputs[2362]) & ~(layer1_outputs[7071]);
    assign layer2_outputs[5987] = layer1_outputs[4221];
    assign layer2_outputs[5988] = ~(layer1_outputs[6679]);
    assign layer2_outputs[5989] = ~((layer1_outputs[11779]) ^ (layer1_outputs[10602]));
    assign layer2_outputs[5990] = ~(layer1_outputs[4684]);
    assign layer2_outputs[5991] = ~(layer1_outputs[11968]);
    assign layer2_outputs[5992] = ~(layer1_outputs[9411]);
    assign layer2_outputs[5993] = (layer1_outputs[3887]) & (layer1_outputs[5587]);
    assign layer2_outputs[5994] = (layer1_outputs[7518]) & (layer1_outputs[12521]);
    assign layer2_outputs[5995] = ~(layer1_outputs[11653]) | (layer1_outputs[11580]);
    assign layer2_outputs[5996] = ~(layer1_outputs[7213]);
    assign layer2_outputs[5997] = ~((layer1_outputs[3242]) | (layer1_outputs[24]));
    assign layer2_outputs[5998] = ~(layer1_outputs[11659]);
    assign layer2_outputs[5999] = ~(layer1_outputs[7599]);
    assign layer2_outputs[6000] = layer1_outputs[10552];
    assign layer2_outputs[6001] = ~(layer1_outputs[8510]) | (layer1_outputs[1268]);
    assign layer2_outputs[6002] = (layer1_outputs[12601]) ^ (layer1_outputs[10562]);
    assign layer2_outputs[6003] = ~(layer1_outputs[4428]);
    assign layer2_outputs[6004] = (layer1_outputs[2470]) & ~(layer1_outputs[6751]);
    assign layer2_outputs[6005] = layer1_outputs[6374];
    assign layer2_outputs[6006] = ~(layer1_outputs[9357]);
    assign layer2_outputs[6007] = layer1_outputs[8628];
    assign layer2_outputs[6008] = layer1_outputs[7647];
    assign layer2_outputs[6009] = (layer1_outputs[12717]) & (layer1_outputs[7264]);
    assign layer2_outputs[6010] = layer1_outputs[5772];
    assign layer2_outputs[6011] = layer1_outputs[10456];
    assign layer2_outputs[6012] = layer1_outputs[7442];
    assign layer2_outputs[6013] = ~(layer1_outputs[7817]);
    assign layer2_outputs[6014] = ~(layer1_outputs[8079]);
    assign layer2_outputs[6015] = ~(layer1_outputs[2685]);
    assign layer2_outputs[6016] = (layer1_outputs[10381]) & ~(layer1_outputs[6007]);
    assign layer2_outputs[6017] = ~(layer1_outputs[527]) | (layer1_outputs[3290]);
    assign layer2_outputs[6018] = ~(layer1_outputs[725]) | (layer1_outputs[6617]);
    assign layer2_outputs[6019] = ~(layer1_outputs[8883]);
    assign layer2_outputs[6020] = ~(layer1_outputs[10887]);
    assign layer2_outputs[6021] = ~((layer1_outputs[4167]) | (layer1_outputs[11104]));
    assign layer2_outputs[6022] = ~(layer1_outputs[10317]);
    assign layer2_outputs[6023] = (layer1_outputs[1355]) ^ (layer1_outputs[1341]);
    assign layer2_outputs[6024] = ~((layer1_outputs[2238]) | (layer1_outputs[6729]));
    assign layer2_outputs[6025] = ~(layer1_outputs[1157]);
    assign layer2_outputs[6026] = ~((layer1_outputs[6228]) & (layer1_outputs[8080]));
    assign layer2_outputs[6027] = layer1_outputs[2682];
    assign layer2_outputs[6028] = ~((layer1_outputs[3213]) ^ (layer1_outputs[5740]));
    assign layer2_outputs[6029] = ~(layer1_outputs[5720]);
    assign layer2_outputs[6030] = (layer1_outputs[6989]) & (layer1_outputs[11427]);
    assign layer2_outputs[6031] = ~(layer1_outputs[10719]) | (layer1_outputs[8146]);
    assign layer2_outputs[6032] = layer1_outputs[9374];
    assign layer2_outputs[6033] = layer1_outputs[11405];
    assign layer2_outputs[6034] = ~(layer1_outputs[8900]);
    assign layer2_outputs[6035] = (layer1_outputs[10186]) & ~(layer1_outputs[8106]);
    assign layer2_outputs[6036] = (layer1_outputs[11295]) ^ (layer1_outputs[9557]);
    assign layer2_outputs[6037] = layer1_outputs[3458];
    assign layer2_outputs[6038] = ~(layer1_outputs[12564]);
    assign layer2_outputs[6039] = ~(layer1_outputs[12145]) | (layer1_outputs[9917]);
    assign layer2_outputs[6040] = layer1_outputs[3954];
    assign layer2_outputs[6041] = (layer1_outputs[11727]) & ~(layer1_outputs[310]);
    assign layer2_outputs[6042] = layer1_outputs[12536];
    assign layer2_outputs[6043] = ~(layer1_outputs[4973]);
    assign layer2_outputs[6044] = layer1_outputs[2057];
    assign layer2_outputs[6045] = (layer1_outputs[5655]) & ~(layer1_outputs[5906]);
    assign layer2_outputs[6046] = ~(layer1_outputs[8940]);
    assign layer2_outputs[6047] = ~(layer1_outputs[11414]) | (layer1_outputs[2019]);
    assign layer2_outputs[6048] = ~(layer1_outputs[1139]) | (layer1_outputs[6812]);
    assign layer2_outputs[6049] = layer1_outputs[10913];
    assign layer2_outputs[6050] = (layer1_outputs[9915]) & ~(layer1_outputs[1168]);
    assign layer2_outputs[6051] = (layer1_outputs[810]) & (layer1_outputs[4636]);
    assign layer2_outputs[6052] = ~(layer1_outputs[9520]);
    assign layer2_outputs[6053] = ~(layer1_outputs[1970]) | (layer1_outputs[12168]);
    assign layer2_outputs[6054] = ~((layer1_outputs[3759]) & (layer1_outputs[10361]));
    assign layer2_outputs[6055] = ~((layer1_outputs[3585]) & (layer1_outputs[187]));
    assign layer2_outputs[6056] = ~(layer1_outputs[8509]);
    assign layer2_outputs[6057] = ~(layer1_outputs[3309]);
    assign layer2_outputs[6058] = layer1_outputs[10543];
    assign layer2_outputs[6059] = ~(layer1_outputs[11205]);
    assign layer2_outputs[6060] = layer1_outputs[6842];
    assign layer2_outputs[6061] = ~((layer1_outputs[7505]) ^ (layer1_outputs[9110]));
    assign layer2_outputs[6062] = 1'b1;
    assign layer2_outputs[6063] = ~(layer1_outputs[9743]);
    assign layer2_outputs[6064] = layer1_outputs[9896];
    assign layer2_outputs[6065] = (layer1_outputs[6123]) & (layer1_outputs[3099]);
    assign layer2_outputs[6066] = ~(layer1_outputs[9316]);
    assign layer2_outputs[6067] = (layer1_outputs[10402]) & ~(layer1_outputs[728]);
    assign layer2_outputs[6068] = layer1_outputs[9744];
    assign layer2_outputs[6069] = ~(layer1_outputs[275]) | (layer1_outputs[11813]);
    assign layer2_outputs[6070] = ~(layer1_outputs[1387]);
    assign layer2_outputs[6071] = ~(layer1_outputs[6279]) | (layer1_outputs[1276]);
    assign layer2_outputs[6072] = (layer1_outputs[2439]) & (layer1_outputs[775]);
    assign layer2_outputs[6073] = ~(layer1_outputs[4258]) | (layer1_outputs[5939]);
    assign layer2_outputs[6074] = ~(layer1_outputs[119]);
    assign layer2_outputs[6075] = (layer1_outputs[8592]) & ~(layer1_outputs[11728]);
    assign layer2_outputs[6076] = (layer1_outputs[5396]) ^ (layer1_outputs[9871]);
    assign layer2_outputs[6077] = (layer1_outputs[1773]) ^ (layer1_outputs[3414]);
    assign layer2_outputs[6078] = (layer1_outputs[7250]) & ~(layer1_outputs[2319]);
    assign layer2_outputs[6079] = ~(layer1_outputs[8390]) | (layer1_outputs[8906]);
    assign layer2_outputs[6080] = layer1_outputs[3254];
    assign layer2_outputs[6081] = layer1_outputs[3341];
    assign layer2_outputs[6082] = (layer1_outputs[8651]) & ~(layer1_outputs[11892]);
    assign layer2_outputs[6083] = ~(layer1_outputs[10618]) | (layer1_outputs[11495]);
    assign layer2_outputs[6084] = ~((layer1_outputs[11924]) | (layer1_outputs[9987]));
    assign layer2_outputs[6085] = layer1_outputs[5469];
    assign layer2_outputs[6086] = layer1_outputs[8560];
    assign layer2_outputs[6087] = ~((layer1_outputs[1187]) ^ (layer1_outputs[12488]));
    assign layer2_outputs[6088] = (layer1_outputs[2602]) & ~(layer1_outputs[4414]);
    assign layer2_outputs[6089] = ~((layer1_outputs[7418]) ^ (layer1_outputs[8163]));
    assign layer2_outputs[6090] = (layer1_outputs[8763]) | (layer1_outputs[7413]);
    assign layer2_outputs[6091] = layer1_outputs[8481];
    assign layer2_outputs[6092] = layer1_outputs[6061];
    assign layer2_outputs[6093] = ~(layer1_outputs[8108]) | (layer1_outputs[12524]);
    assign layer2_outputs[6094] = (layer1_outputs[9818]) ^ (layer1_outputs[8317]);
    assign layer2_outputs[6095] = ~((layer1_outputs[1453]) | (layer1_outputs[7317]));
    assign layer2_outputs[6096] = (layer1_outputs[9703]) & ~(layer1_outputs[1963]);
    assign layer2_outputs[6097] = ~((layer1_outputs[8561]) & (layer1_outputs[4762]));
    assign layer2_outputs[6098] = layer1_outputs[5462];
    assign layer2_outputs[6099] = layer1_outputs[7033];
    assign layer2_outputs[6100] = ~(layer1_outputs[3510]);
    assign layer2_outputs[6101] = layer1_outputs[8909];
    assign layer2_outputs[6102] = layer1_outputs[2777];
    assign layer2_outputs[6103] = layer1_outputs[87];
    assign layer2_outputs[6104] = ~((layer1_outputs[10186]) ^ (layer1_outputs[2158]));
    assign layer2_outputs[6105] = (layer1_outputs[7963]) & ~(layer1_outputs[12486]);
    assign layer2_outputs[6106] = (layer1_outputs[2217]) & (layer1_outputs[425]);
    assign layer2_outputs[6107] = layer1_outputs[12325];
    assign layer2_outputs[6108] = layer1_outputs[9980];
    assign layer2_outputs[6109] = (layer1_outputs[11186]) ^ (layer1_outputs[3980]);
    assign layer2_outputs[6110] = ~((layer1_outputs[5937]) & (layer1_outputs[11329]));
    assign layer2_outputs[6111] = ~((layer1_outputs[1327]) ^ (layer1_outputs[8922]));
    assign layer2_outputs[6112] = ~((layer1_outputs[6124]) | (layer1_outputs[5785]));
    assign layer2_outputs[6113] = ~((layer1_outputs[8332]) & (layer1_outputs[8264]));
    assign layer2_outputs[6114] = (layer1_outputs[9940]) ^ (layer1_outputs[2550]);
    assign layer2_outputs[6115] = ~((layer1_outputs[9887]) & (layer1_outputs[6897]));
    assign layer2_outputs[6116] = layer1_outputs[5650];
    assign layer2_outputs[6117] = (layer1_outputs[10184]) & ~(layer1_outputs[7764]);
    assign layer2_outputs[6118] = (layer1_outputs[4202]) & ~(layer1_outputs[10990]);
    assign layer2_outputs[6119] = ~(layer1_outputs[1474]);
    assign layer2_outputs[6120] = ~(layer1_outputs[10323]);
    assign layer2_outputs[6121] = ~((layer1_outputs[4854]) & (layer1_outputs[3381]));
    assign layer2_outputs[6122] = (layer1_outputs[8954]) ^ (layer1_outputs[6343]);
    assign layer2_outputs[6123] = ~(layer1_outputs[12662]);
    assign layer2_outputs[6124] = (layer1_outputs[10197]) & ~(layer1_outputs[3176]);
    assign layer2_outputs[6125] = ~(layer1_outputs[5663]) | (layer1_outputs[9321]);
    assign layer2_outputs[6126] = (layer1_outputs[6605]) & ~(layer1_outputs[9443]);
    assign layer2_outputs[6127] = layer1_outputs[3133];
    assign layer2_outputs[6128] = ~((layer1_outputs[938]) & (layer1_outputs[12354]));
    assign layer2_outputs[6129] = ~(layer1_outputs[2679]);
    assign layer2_outputs[6130] = layer1_outputs[1603];
    assign layer2_outputs[6131] = layer1_outputs[10924];
    assign layer2_outputs[6132] = ~(layer1_outputs[4888]);
    assign layer2_outputs[6133] = layer1_outputs[12760];
    assign layer2_outputs[6134] = ~(layer1_outputs[5163]) | (layer1_outputs[2020]);
    assign layer2_outputs[6135] = ~(layer1_outputs[12720]);
    assign layer2_outputs[6136] = ~((layer1_outputs[134]) | (layer1_outputs[9948]));
    assign layer2_outputs[6137] = layer1_outputs[2554];
    assign layer2_outputs[6138] = ~(layer1_outputs[3513]) | (layer1_outputs[5189]);
    assign layer2_outputs[6139] = (layer1_outputs[1259]) & ~(layer1_outputs[9460]);
    assign layer2_outputs[6140] = layer1_outputs[9003];
    assign layer2_outputs[6141] = ~(layer1_outputs[9255]) | (layer1_outputs[4764]);
    assign layer2_outputs[6142] = ~(layer1_outputs[4237]);
    assign layer2_outputs[6143] = ~(layer1_outputs[8852]) | (layer1_outputs[4727]);
    assign layer2_outputs[6144] = layer1_outputs[880];
    assign layer2_outputs[6145] = ~(layer1_outputs[4462]);
    assign layer2_outputs[6146] = ~((layer1_outputs[8122]) ^ (layer1_outputs[8236]));
    assign layer2_outputs[6147] = layer1_outputs[5056];
    assign layer2_outputs[6148] = (layer1_outputs[194]) ^ (layer1_outputs[4095]);
    assign layer2_outputs[6149] = (layer1_outputs[691]) & (layer1_outputs[12752]);
    assign layer2_outputs[6150] = (layer1_outputs[1149]) | (layer1_outputs[12459]);
    assign layer2_outputs[6151] = ~(layer1_outputs[8302]);
    assign layer2_outputs[6152] = layer1_outputs[3629];
    assign layer2_outputs[6153] = layer1_outputs[4937];
    assign layer2_outputs[6154] = ~(layer1_outputs[7886]);
    assign layer2_outputs[6155] = layer1_outputs[7988];
    assign layer2_outputs[6156] = ~((layer1_outputs[2951]) & (layer1_outputs[7832]));
    assign layer2_outputs[6157] = ~((layer1_outputs[8358]) & (layer1_outputs[6062]));
    assign layer2_outputs[6158] = layer1_outputs[5083];
    assign layer2_outputs[6159] = ~(layer1_outputs[6515]) | (layer1_outputs[8337]);
    assign layer2_outputs[6160] = ~((layer1_outputs[9016]) | (layer1_outputs[2253]));
    assign layer2_outputs[6161] = layer1_outputs[6604];
    assign layer2_outputs[6162] = ~(layer1_outputs[8960]);
    assign layer2_outputs[6163] = ~(layer1_outputs[9226]);
    assign layer2_outputs[6164] = ~(layer1_outputs[10457]);
    assign layer2_outputs[6165] = ~(layer1_outputs[1680]) | (layer1_outputs[9295]);
    assign layer2_outputs[6166] = ~(layer1_outputs[3618]);
    assign layer2_outputs[6167] = ~(layer1_outputs[10817]);
    assign layer2_outputs[6168] = ~(layer1_outputs[5381]);
    assign layer2_outputs[6169] = ~(layer1_outputs[5941]);
    assign layer2_outputs[6170] = layer1_outputs[3421];
    assign layer2_outputs[6171] = layer1_outputs[11364];
    assign layer2_outputs[6172] = (layer1_outputs[9754]) ^ (layer1_outputs[1154]);
    assign layer2_outputs[6173] = ~(layer1_outputs[3468]);
    assign layer2_outputs[6174] = layer1_outputs[1467];
    assign layer2_outputs[6175] = layer1_outputs[7547];
    assign layer2_outputs[6176] = 1'b1;
    assign layer2_outputs[6177] = (layer1_outputs[5122]) | (layer1_outputs[10630]);
    assign layer2_outputs[6178] = ~(layer1_outputs[3283]);
    assign layer2_outputs[6179] = layer1_outputs[10311];
    assign layer2_outputs[6180] = (layer1_outputs[5306]) & ~(layer1_outputs[6134]);
    assign layer2_outputs[6181] = 1'b1;
    assign layer2_outputs[6182] = layer1_outputs[2051];
    assign layer2_outputs[6183] = ~((layer1_outputs[844]) | (layer1_outputs[12629]));
    assign layer2_outputs[6184] = 1'b1;
    assign layer2_outputs[6185] = (layer1_outputs[1511]) | (layer1_outputs[8503]);
    assign layer2_outputs[6186] = (layer1_outputs[5130]) | (layer1_outputs[2262]);
    assign layer2_outputs[6187] = ~(layer1_outputs[9181]);
    assign layer2_outputs[6188] = ~(layer1_outputs[11782]) | (layer1_outputs[4900]);
    assign layer2_outputs[6189] = (layer1_outputs[2035]) ^ (layer1_outputs[12725]);
    assign layer2_outputs[6190] = ~(layer1_outputs[4354]);
    assign layer2_outputs[6191] = ~(layer1_outputs[8110]);
    assign layer2_outputs[6192] = (layer1_outputs[10651]) ^ (layer1_outputs[12698]);
    assign layer2_outputs[6193] = ~(layer1_outputs[10744]);
    assign layer2_outputs[6194] = ~(layer1_outputs[8817]);
    assign layer2_outputs[6195] = layer1_outputs[7559];
    assign layer2_outputs[6196] = layer1_outputs[1829];
    assign layer2_outputs[6197] = (layer1_outputs[11246]) & ~(layer1_outputs[7447]);
    assign layer2_outputs[6198] = ~((layer1_outputs[11535]) & (layer1_outputs[10784]));
    assign layer2_outputs[6199] = (layer1_outputs[2519]) ^ (layer1_outputs[52]);
    assign layer2_outputs[6200] = ~(layer1_outputs[8485]) | (layer1_outputs[8353]);
    assign layer2_outputs[6201] = ~((layer1_outputs[1774]) & (layer1_outputs[9841]));
    assign layer2_outputs[6202] = 1'b0;
    assign layer2_outputs[6203] = ~((layer1_outputs[12682]) & (layer1_outputs[7970]));
    assign layer2_outputs[6204] = ~(layer1_outputs[9043]);
    assign layer2_outputs[6205] = ~(layer1_outputs[237]) | (layer1_outputs[4248]);
    assign layer2_outputs[6206] = layer1_outputs[11893];
    assign layer2_outputs[6207] = (layer1_outputs[2005]) & ~(layer1_outputs[1038]);
    assign layer2_outputs[6208] = ~(layer1_outputs[3611]) | (layer1_outputs[11450]);
    assign layer2_outputs[6209] = ~(layer1_outputs[9743]);
    assign layer2_outputs[6210] = ~(layer1_outputs[11670]);
    assign layer2_outputs[6211] = ~(layer1_outputs[8804]);
    assign layer2_outputs[6212] = ~((layer1_outputs[338]) ^ (layer1_outputs[7712]));
    assign layer2_outputs[6213] = (layer1_outputs[7469]) & ~(layer1_outputs[681]);
    assign layer2_outputs[6214] = layer1_outputs[10156];
    assign layer2_outputs[6215] = ~(layer1_outputs[614]);
    assign layer2_outputs[6216] = ~(layer1_outputs[2115]);
    assign layer2_outputs[6217] = (layer1_outputs[2435]) & (layer1_outputs[8565]);
    assign layer2_outputs[6218] = ~(layer1_outputs[1071]);
    assign layer2_outputs[6219] = ~(layer1_outputs[2315]) | (layer1_outputs[10288]);
    assign layer2_outputs[6220] = ~(layer1_outputs[4787]);
    assign layer2_outputs[6221] = (layer1_outputs[9521]) ^ (layer1_outputs[9116]);
    assign layer2_outputs[6222] = ~(layer1_outputs[11369]);
    assign layer2_outputs[6223] = ~(layer1_outputs[5600]);
    assign layer2_outputs[6224] = ~(layer1_outputs[6207]);
    assign layer2_outputs[6225] = (layer1_outputs[4115]) & ~(layer1_outputs[5062]);
    assign layer2_outputs[6226] = ~((layer1_outputs[11588]) ^ (layer1_outputs[665]));
    assign layer2_outputs[6227] = (layer1_outputs[6891]) ^ (layer1_outputs[12572]);
    assign layer2_outputs[6228] = (layer1_outputs[9050]) | (layer1_outputs[8881]);
    assign layer2_outputs[6229] = (layer1_outputs[4817]) ^ (layer1_outputs[12378]);
    assign layer2_outputs[6230] = ~((layer1_outputs[7844]) & (layer1_outputs[7434]));
    assign layer2_outputs[6231] = layer1_outputs[8319];
    assign layer2_outputs[6232] = ~((layer1_outputs[2285]) ^ (layer1_outputs[4324]));
    assign layer2_outputs[6233] = ~(layer1_outputs[7858]);
    assign layer2_outputs[6234] = (layer1_outputs[1884]) ^ (layer1_outputs[8208]);
    assign layer2_outputs[6235] = ~(layer1_outputs[3832]) | (layer1_outputs[4676]);
    assign layer2_outputs[6236] = layer1_outputs[6250];
    assign layer2_outputs[6237] = (layer1_outputs[12210]) & ~(layer1_outputs[11213]);
    assign layer2_outputs[6238] = ~(layer1_outputs[2335]) | (layer1_outputs[7229]);
    assign layer2_outputs[6239] = (layer1_outputs[5115]) & (layer1_outputs[12003]);
    assign layer2_outputs[6240] = layer1_outputs[2314];
    assign layer2_outputs[6241] = layer1_outputs[432];
    assign layer2_outputs[6242] = (layer1_outputs[10481]) | (layer1_outputs[3088]);
    assign layer2_outputs[6243] = layer1_outputs[8976];
    assign layer2_outputs[6244] = layer1_outputs[712];
    assign layer2_outputs[6245] = ~(layer1_outputs[3825]) | (layer1_outputs[7830]);
    assign layer2_outputs[6246] = ~(layer1_outputs[12559]);
    assign layer2_outputs[6247] = layer1_outputs[709];
    assign layer2_outputs[6248] = ~(layer1_outputs[8322]);
    assign layer2_outputs[6249] = ~(layer1_outputs[429]);
    assign layer2_outputs[6250] = ~(layer1_outputs[5870]) | (layer1_outputs[11829]);
    assign layer2_outputs[6251] = (layer1_outputs[2034]) | (layer1_outputs[11303]);
    assign layer2_outputs[6252] = layer1_outputs[10700];
    assign layer2_outputs[6253] = ~(layer1_outputs[8035]);
    assign layer2_outputs[6254] = ~(layer1_outputs[2466]);
    assign layer2_outputs[6255] = layer1_outputs[12359];
    assign layer2_outputs[6256] = (layer1_outputs[2858]) & ~(layer1_outputs[8491]);
    assign layer2_outputs[6257] = layer1_outputs[4603];
    assign layer2_outputs[6258] = layer1_outputs[1381];
    assign layer2_outputs[6259] = ~(layer1_outputs[12661]);
    assign layer2_outputs[6260] = (layer1_outputs[1088]) ^ (layer1_outputs[9968]);
    assign layer2_outputs[6261] = ~(layer1_outputs[8472]);
    assign layer2_outputs[6262] = (layer1_outputs[5285]) | (layer1_outputs[1728]);
    assign layer2_outputs[6263] = ~(layer1_outputs[2870]) | (layer1_outputs[9550]);
    assign layer2_outputs[6264] = layer1_outputs[4208];
    assign layer2_outputs[6265] = ~(layer1_outputs[5815]);
    assign layer2_outputs[6266] = (layer1_outputs[9010]) & ~(layer1_outputs[9201]);
    assign layer2_outputs[6267] = (layer1_outputs[11916]) & ~(layer1_outputs[6644]);
    assign layer2_outputs[6268] = (layer1_outputs[9729]) | (layer1_outputs[7198]);
    assign layer2_outputs[6269] = ~(layer1_outputs[4839]);
    assign layer2_outputs[6270] = ~(layer1_outputs[7488]);
    assign layer2_outputs[6271] = layer1_outputs[81];
    assign layer2_outputs[6272] = layer1_outputs[12136];
    assign layer2_outputs[6273] = ~((layer1_outputs[10756]) & (layer1_outputs[963]));
    assign layer2_outputs[6274] = (layer1_outputs[3061]) ^ (layer1_outputs[8739]);
    assign layer2_outputs[6275] = (layer1_outputs[9206]) | (layer1_outputs[1903]);
    assign layer2_outputs[6276] = ~(layer1_outputs[9911]);
    assign layer2_outputs[6277] = ~((layer1_outputs[7132]) ^ (layer1_outputs[126]));
    assign layer2_outputs[6278] = ~(layer1_outputs[7816]);
    assign layer2_outputs[6279] = ~(layer1_outputs[12611]);
    assign layer2_outputs[6280] = ~(layer1_outputs[8598]);
    assign layer2_outputs[6281] = ~(layer1_outputs[6133]);
    assign layer2_outputs[6282] = layer1_outputs[4644];
    assign layer2_outputs[6283] = ~(layer1_outputs[3513]);
    assign layer2_outputs[6284] = layer1_outputs[536];
    assign layer2_outputs[6285] = ~((layer1_outputs[3795]) | (layer1_outputs[439]));
    assign layer2_outputs[6286] = layer1_outputs[3394];
    assign layer2_outputs[6287] = layer1_outputs[4566];
    assign layer2_outputs[6288] = layer1_outputs[4932];
    assign layer2_outputs[6289] = (layer1_outputs[2280]) & ~(layer1_outputs[7990]);
    assign layer2_outputs[6290] = (layer1_outputs[416]) & (layer1_outputs[11858]);
    assign layer2_outputs[6291] = ~(layer1_outputs[2179]);
    assign layer2_outputs[6292] = 1'b1;
    assign layer2_outputs[6293] = ~(layer1_outputs[1736]);
    assign layer2_outputs[6294] = ~(layer1_outputs[3463]);
    assign layer2_outputs[6295] = (layer1_outputs[11038]) & ~(layer1_outputs[744]);
    assign layer2_outputs[6296] = (layer1_outputs[1450]) & (layer1_outputs[5147]);
    assign layer2_outputs[6297] = layer1_outputs[8867];
    assign layer2_outputs[6298] = ~(layer1_outputs[9390]);
    assign layer2_outputs[6299] = ~((layer1_outputs[2317]) ^ (layer1_outputs[10747]));
    assign layer2_outputs[6300] = ~((layer1_outputs[3346]) ^ (layer1_outputs[5181]));
    assign layer2_outputs[6301] = layer1_outputs[317];
    assign layer2_outputs[6302] = (layer1_outputs[10258]) ^ (layer1_outputs[12494]);
    assign layer2_outputs[6303] = ~(layer1_outputs[8013]);
    assign layer2_outputs[6304] = ~(layer1_outputs[9065]);
    assign layer2_outputs[6305] = ~((layer1_outputs[11943]) ^ (layer1_outputs[10493]));
    assign layer2_outputs[6306] = ~(layer1_outputs[11109]);
    assign layer2_outputs[6307] = ~(layer1_outputs[1750]);
    assign layer2_outputs[6308] = ~((layer1_outputs[3046]) | (layer1_outputs[6976]));
    assign layer2_outputs[6309] = ~(layer1_outputs[6581]);
    assign layer2_outputs[6310] = ~(layer1_outputs[10118]);
    assign layer2_outputs[6311] = ~(layer1_outputs[5572]);
    assign layer2_outputs[6312] = ~(layer1_outputs[9301]);
    assign layer2_outputs[6313] = ~((layer1_outputs[8706]) | (layer1_outputs[9010]));
    assign layer2_outputs[6314] = (layer1_outputs[5484]) & ~(layer1_outputs[3081]);
    assign layer2_outputs[6315] = layer1_outputs[6169];
    assign layer2_outputs[6316] = ~(layer1_outputs[1916]);
    assign layer2_outputs[6317] = (layer1_outputs[1755]) | (layer1_outputs[12421]);
    assign layer2_outputs[6318] = ~((layer1_outputs[4935]) & (layer1_outputs[869]));
    assign layer2_outputs[6319] = layer1_outputs[8611];
    assign layer2_outputs[6320] = ~((layer1_outputs[2974]) | (layer1_outputs[10770]));
    assign layer2_outputs[6321] = layer1_outputs[10358];
    assign layer2_outputs[6322] = layer1_outputs[414];
    assign layer2_outputs[6323] = ~((layer1_outputs[1799]) & (layer1_outputs[501]));
    assign layer2_outputs[6324] = layer1_outputs[8285];
    assign layer2_outputs[6325] = ~(layer1_outputs[1360]);
    assign layer2_outputs[6326] = ~(layer1_outputs[7188]);
    assign layer2_outputs[6327] = ~(layer1_outputs[9021]);
    assign layer2_outputs[6328] = (layer1_outputs[5701]) & (layer1_outputs[4304]);
    assign layer2_outputs[6329] = ~(layer1_outputs[8522]);
    assign layer2_outputs[6330] = ~(layer1_outputs[5218]);
    assign layer2_outputs[6331] = layer1_outputs[6610];
    assign layer2_outputs[6332] = ~((layer1_outputs[8935]) & (layer1_outputs[8252]));
    assign layer2_outputs[6333] = (layer1_outputs[1697]) & ~(layer1_outputs[6152]);
    assign layer2_outputs[6334] = layer1_outputs[8289];
    assign layer2_outputs[6335] = ~((layer1_outputs[2261]) ^ (layer1_outputs[3958]));
    assign layer2_outputs[6336] = ~(layer1_outputs[160]) | (layer1_outputs[5989]);
    assign layer2_outputs[6337] = layer1_outputs[10695];
    assign layer2_outputs[6338] = ~(layer1_outputs[4296]);
    assign layer2_outputs[6339] = layer1_outputs[6851];
    assign layer2_outputs[6340] = layer1_outputs[10233];
    assign layer2_outputs[6341] = ~(layer1_outputs[9463]);
    assign layer2_outputs[6342] = ~((layer1_outputs[8184]) | (layer1_outputs[7210]));
    assign layer2_outputs[6343] = (layer1_outputs[3783]) ^ (layer1_outputs[12272]);
    assign layer2_outputs[6344] = (layer1_outputs[10871]) & ~(layer1_outputs[12560]);
    assign layer2_outputs[6345] = (layer1_outputs[3197]) & (layer1_outputs[877]);
    assign layer2_outputs[6346] = ~(layer1_outputs[3530]);
    assign layer2_outputs[6347] = (layer1_outputs[4552]) ^ (layer1_outputs[11733]);
    assign layer2_outputs[6348] = (layer1_outputs[7874]) & (layer1_outputs[10596]);
    assign layer2_outputs[6349] = ~(layer1_outputs[10870]) | (layer1_outputs[2722]);
    assign layer2_outputs[6350] = ~(layer1_outputs[9020]);
    assign layer2_outputs[6351] = ~((layer1_outputs[9828]) ^ (layer1_outputs[1608]));
    assign layer2_outputs[6352] = ~(layer1_outputs[2177]) | (layer1_outputs[2344]);
    assign layer2_outputs[6353] = ~((layer1_outputs[205]) ^ (layer1_outputs[6549]));
    assign layer2_outputs[6354] = layer1_outputs[359];
    assign layer2_outputs[6355] = layer1_outputs[5110];
    assign layer2_outputs[6356] = (layer1_outputs[11215]) ^ (layer1_outputs[2615]);
    assign layer2_outputs[6357] = layer1_outputs[76];
    assign layer2_outputs[6358] = ~((layer1_outputs[4340]) & (layer1_outputs[8314]));
    assign layer2_outputs[6359] = ~((layer1_outputs[5657]) & (layer1_outputs[7546]));
    assign layer2_outputs[6360] = (layer1_outputs[6733]) | (layer1_outputs[11175]);
    assign layer2_outputs[6361] = (layer1_outputs[6882]) & ~(layer1_outputs[7405]);
    assign layer2_outputs[6362] = (layer1_outputs[8557]) | (layer1_outputs[11674]);
    assign layer2_outputs[6363] = (layer1_outputs[5724]) ^ (layer1_outputs[2928]);
    assign layer2_outputs[6364] = ~(layer1_outputs[12776]) | (layer1_outputs[11498]);
    assign layer2_outputs[6365] = ~(layer1_outputs[6159]);
    assign layer2_outputs[6366] = ~((layer1_outputs[9829]) ^ (layer1_outputs[4825]));
    assign layer2_outputs[6367] = layer1_outputs[820];
    assign layer2_outputs[6368] = (layer1_outputs[854]) & (layer1_outputs[11497]);
    assign layer2_outputs[6369] = layer1_outputs[6108];
    assign layer2_outputs[6370] = (layer1_outputs[7528]) | (layer1_outputs[12002]);
    assign layer2_outputs[6371] = ~(layer1_outputs[10587]);
    assign layer2_outputs[6372] = ~(layer1_outputs[1257]);
    assign layer2_outputs[6373] = ~(layer1_outputs[5171]);
    assign layer2_outputs[6374] = ~(layer1_outputs[1163]);
    assign layer2_outputs[6375] = ~(layer1_outputs[12309]);
    assign layer2_outputs[6376] = ~(layer1_outputs[4210]);
    assign layer2_outputs[6377] = layer1_outputs[7842];
    assign layer2_outputs[6378] = (layer1_outputs[6275]) & ~(layer1_outputs[2659]);
    assign layer2_outputs[6379] = ~(layer1_outputs[363]) | (layer1_outputs[11170]);
    assign layer2_outputs[6380] = ~((layer1_outputs[2753]) ^ (layer1_outputs[9394]));
    assign layer2_outputs[6381] = (layer1_outputs[5787]) ^ (layer1_outputs[3975]);
    assign layer2_outputs[6382] = ~((layer1_outputs[6193]) ^ (layer1_outputs[6004]));
    assign layer2_outputs[6383] = ~(layer1_outputs[9749]);
    assign layer2_outputs[6384] = ~(layer1_outputs[4125]);
    assign layer2_outputs[6385] = layer1_outputs[3215];
    assign layer2_outputs[6386] = ~(layer1_outputs[10271]);
    assign layer2_outputs[6387] = ~(layer1_outputs[6728]);
    assign layer2_outputs[6388] = (layer1_outputs[965]) & ~(layer1_outputs[7513]);
    assign layer2_outputs[6389] = layer1_outputs[7090];
    assign layer2_outputs[6390] = (layer1_outputs[1812]) & ~(layer1_outputs[9698]);
    assign layer2_outputs[6391] = ~(layer1_outputs[983]) | (layer1_outputs[12342]);
    assign layer2_outputs[6392] = ~((layer1_outputs[12019]) ^ (layer1_outputs[1190]));
    assign layer2_outputs[6393] = (layer1_outputs[6435]) & (layer1_outputs[4037]);
    assign layer2_outputs[6394] = ~(layer1_outputs[4511]) | (layer1_outputs[10505]);
    assign layer2_outputs[6395] = (layer1_outputs[4748]) ^ (layer1_outputs[865]);
    assign layer2_outputs[6396] = layer1_outputs[7891];
    assign layer2_outputs[6397] = ~(layer1_outputs[5019]) | (layer1_outputs[2237]);
    assign layer2_outputs[6398] = ~(layer1_outputs[11645]) | (layer1_outputs[2090]);
    assign layer2_outputs[6399] = ~(layer1_outputs[4048]);
    assign layer2_outputs[6400] = ~(layer1_outputs[3994]) | (layer1_outputs[2511]);
    assign layer2_outputs[6401] = (layer1_outputs[9122]) & (layer1_outputs[12395]);
    assign layer2_outputs[6402] = ~(layer1_outputs[5850]);
    assign layer2_outputs[6403] = ~(layer1_outputs[7222]) | (layer1_outputs[8562]);
    assign layer2_outputs[6404] = ~(layer1_outputs[5117]);
    assign layer2_outputs[6405] = ~(layer1_outputs[927]);
    assign layer2_outputs[6406] = (layer1_outputs[2764]) & ~(layer1_outputs[7623]);
    assign layer2_outputs[6407] = (layer1_outputs[9512]) ^ (layer1_outputs[4840]);
    assign layer2_outputs[6408] = (layer1_outputs[11304]) & (layer1_outputs[2156]);
    assign layer2_outputs[6409] = layer1_outputs[3299];
    assign layer2_outputs[6410] = ~(layer1_outputs[2564]);
    assign layer2_outputs[6411] = (layer1_outputs[6804]) ^ (layer1_outputs[11357]);
    assign layer2_outputs[6412] = layer1_outputs[4502];
    assign layer2_outputs[6413] = (layer1_outputs[9502]) | (layer1_outputs[7711]);
    assign layer2_outputs[6414] = ~((layer1_outputs[1852]) | (layer1_outputs[3937]));
    assign layer2_outputs[6415] = layer1_outputs[7932];
    assign layer2_outputs[6416] = ~((layer1_outputs[1943]) | (layer1_outputs[5251]));
    assign layer2_outputs[6417] = (layer1_outputs[6960]) ^ (layer1_outputs[12518]);
    assign layer2_outputs[6418] = layer1_outputs[9548];
    assign layer2_outputs[6419] = ~(layer1_outputs[2309]);
    assign layer2_outputs[6420] = (layer1_outputs[4977]) | (layer1_outputs[5259]);
    assign layer2_outputs[6421] = ~(layer1_outputs[755]);
    assign layer2_outputs[6422] = ~(layer1_outputs[2351]);
    assign layer2_outputs[6423] = (layer1_outputs[5266]) & ~(layer1_outputs[10773]);
    assign layer2_outputs[6424] = (layer1_outputs[11840]) ^ (layer1_outputs[6515]);
    assign layer2_outputs[6425] = (layer1_outputs[6500]) | (layer1_outputs[9147]);
    assign layer2_outputs[6426] = ~(layer1_outputs[11199]);
    assign layer2_outputs[6427] = layer1_outputs[11926];
    assign layer2_outputs[6428] = (layer1_outputs[12214]) | (layer1_outputs[8361]);
    assign layer2_outputs[6429] = layer1_outputs[6075];
    assign layer2_outputs[6430] = ~(layer1_outputs[1231]);
    assign layer2_outputs[6431] = ~(layer1_outputs[11841]);
    assign layer2_outputs[6432] = layer1_outputs[2542];
    assign layer2_outputs[6433] = ~(layer1_outputs[7400]);
    assign layer2_outputs[6434] = (layer1_outputs[2041]) & (layer1_outputs[2533]);
    assign layer2_outputs[6435] = ~(layer1_outputs[41]) | (layer1_outputs[1974]);
    assign layer2_outputs[6436] = ~(layer1_outputs[10275]);
    assign layer2_outputs[6437] = layer1_outputs[8490];
    assign layer2_outputs[6438] = layer1_outputs[1333];
    assign layer2_outputs[6439] = ~((layer1_outputs[12068]) ^ (layer1_outputs[5895]));
    assign layer2_outputs[6440] = ~((layer1_outputs[1393]) | (layer1_outputs[5000]));
    assign layer2_outputs[6441] = ~(layer1_outputs[1717]) | (layer1_outputs[7945]);
    assign layer2_outputs[6442] = ~(layer1_outputs[3075]) | (layer1_outputs[10231]);
    assign layer2_outputs[6443] = (layer1_outputs[9655]) | (layer1_outputs[12251]);
    assign layer2_outputs[6444] = ~(layer1_outputs[4988]);
    assign layer2_outputs[6445] = ~((layer1_outputs[3444]) & (layer1_outputs[3233]));
    assign layer2_outputs[6446] = ~(layer1_outputs[6845]);
    assign layer2_outputs[6447] = ~((layer1_outputs[1996]) & (layer1_outputs[6802]));
    assign layer2_outputs[6448] = (layer1_outputs[10837]) & (layer1_outputs[1672]);
    assign layer2_outputs[6449] = layer1_outputs[6668];
    assign layer2_outputs[6450] = ~(layer1_outputs[2418]);
    assign layer2_outputs[6451] = ~(layer1_outputs[9053]);
    assign layer2_outputs[6452] = ~(layer1_outputs[1226]) | (layer1_outputs[11667]);
    assign layer2_outputs[6453] = ~(layer1_outputs[9371]);
    assign layer2_outputs[6454] = ~((layer1_outputs[5725]) | (layer1_outputs[3820]));
    assign layer2_outputs[6455] = layer1_outputs[5621];
    assign layer2_outputs[6456] = ~(layer1_outputs[1507]);
    assign layer2_outputs[6457] = ~((layer1_outputs[3459]) & (layer1_outputs[7104]));
    assign layer2_outputs[6458] = (layer1_outputs[11101]) & (layer1_outputs[1503]);
    assign layer2_outputs[6459] = layer1_outputs[2824];
    assign layer2_outputs[6460] = (layer1_outputs[5085]) & (layer1_outputs[6640]);
    assign layer2_outputs[6461] = layer1_outputs[11785];
    assign layer2_outputs[6462] = ~(layer1_outputs[9519]);
    assign layer2_outputs[6463] = (layer1_outputs[8002]) ^ (layer1_outputs[9977]);
    assign layer2_outputs[6464] = (layer1_outputs[11577]) | (layer1_outputs[440]);
    assign layer2_outputs[6465] = layer1_outputs[9836];
    assign layer2_outputs[6466] = ~((layer1_outputs[5859]) ^ (layer1_outputs[546]));
    assign layer2_outputs[6467] = ~((layer1_outputs[9409]) & (layer1_outputs[5392]));
    assign layer2_outputs[6468] = ~(layer1_outputs[2377]);
    assign layer2_outputs[6469] = layer1_outputs[2884];
    assign layer2_outputs[6470] = layer1_outputs[8454];
    assign layer2_outputs[6471] = ~((layer1_outputs[4161]) | (layer1_outputs[8159]));
    assign layer2_outputs[6472] = layer1_outputs[11407];
    assign layer2_outputs[6473] = (layer1_outputs[9334]) | (layer1_outputs[7393]);
    assign layer2_outputs[6474] = ~((layer1_outputs[7279]) ^ (layer1_outputs[7045]));
    assign layer2_outputs[6475] = ~(layer1_outputs[5947]);
    assign layer2_outputs[6476] = ~(layer1_outputs[10059]);
    assign layer2_outputs[6477] = (layer1_outputs[2410]) & ~(layer1_outputs[1123]);
    assign layer2_outputs[6478] = ~(layer1_outputs[2869]);
    assign layer2_outputs[6479] = ~(layer1_outputs[1320]);
    assign layer2_outputs[6480] = ~(layer1_outputs[1264]) | (layer1_outputs[10074]);
    assign layer2_outputs[6481] = (layer1_outputs[2474]) & ~(layer1_outputs[898]);
    assign layer2_outputs[6482] = (layer1_outputs[7459]) & ~(layer1_outputs[6058]);
    assign layer2_outputs[6483] = layer1_outputs[10324];
    assign layer2_outputs[6484] = ~(layer1_outputs[4154]) | (layer1_outputs[7737]);
    assign layer2_outputs[6485] = layer1_outputs[10041];
    assign layer2_outputs[6486] = ~(layer1_outputs[11480]);
    assign layer2_outputs[6487] = layer1_outputs[9202];
    assign layer2_outputs[6488] = ~(layer1_outputs[8722]);
    assign layer2_outputs[6489] = ~(layer1_outputs[9946]);
    assign layer2_outputs[6490] = ~(layer1_outputs[5164]);
    assign layer2_outputs[6491] = layer1_outputs[2566];
    assign layer2_outputs[6492] = layer1_outputs[11946];
    assign layer2_outputs[6493] = layer1_outputs[3365];
    assign layer2_outputs[6494] = ~(layer1_outputs[12074]) | (layer1_outputs[5247]);
    assign layer2_outputs[6495] = ~(layer1_outputs[5616]) | (layer1_outputs[1325]);
    assign layer2_outputs[6496] = layer1_outputs[807];
    assign layer2_outputs[6497] = 1'b1;
    assign layer2_outputs[6498] = layer1_outputs[1192];
    assign layer2_outputs[6499] = layer1_outputs[8887];
    assign layer2_outputs[6500] = ~((layer1_outputs[2235]) & (layer1_outputs[5604]));
    assign layer2_outputs[6501] = (layer1_outputs[8983]) & (layer1_outputs[776]);
    assign layer2_outputs[6502] = ~((layer1_outputs[999]) ^ (layer1_outputs[3820]));
    assign layer2_outputs[6503] = layer1_outputs[2479];
    assign layer2_outputs[6504] = ~(layer1_outputs[8576]);
    assign layer2_outputs[6505] = layer1_outputs[11489];
    assign layer2_outputs[6506] = (layer1_outputs[11258]) ^ (layer1_outputs[6555]);
    assign layer2_outputs[6507] = layer1_outputs[9764];
    assign layer2_outputs[6508] = layer1_outputs[796];
    assign layer2_outputs[6509] = (layer1_outputs[9387]) | (layer1_outputs[11828]);
    assign layer2_outputs[6510] = layer1_outputs[5133];
    assign layer2_outputs[6511] = (layer1_outputs[7355]) | (layer1_outputs[10616]);
    assign layer2_outputs[6512] = layer1_outputs[10563];
    assign layer2_outputs[6513] = ~(layer1_outputs[1097]);
    assign layer2_outputs[6514] = layer1_outputs[9504];
    assign layer2_outputs[6515] = ~((layer1_outputs[10869]) ^ (layer1_outputs[3195]));
    assign layer2_outputs[6516] = layer1_outputs[4285];
    assign layer2_outputs[6517] = ~(layer1_outputs[10469]);
    assign layer2_outputs[6518] = ~(layer1_outputs[9328]);
    assign layer2_outputs[6519] = ~((layer1_outputs[8188]) ^ (layer1_outputs[695]));
    assign layer2_outputs[6520] = ~(layer1_outputs[7317]);
    assign layer2_outputs[6521] = layer1_outputs[2444];
    assign layer2_outputs[6522] = ~((layer1_outputs[4983]) & (layer1_outputs[118]));
    assign layer2_outputs[6523] = ~(layer1_outputs[296]);
    assign layer2_outputs[6524] = ~(layer1_outputs[23]);
    assign layer2_outputs[6525] = (layer1_outputs[5022]) ^ (layer1_outputs[10078]);
    assign layer2_outputs[6526] = layer1_outputs[11869];
    assign layer2_outputs[6527] = layer1_outputs[4317];
    assign layer2_outputs[6528] = ~(layer1_outputs[7960]);
    assign layer2_outputs[6529] = 1'b0;
    assign layer2_outputs[6530] = layer1_outputs[6753];
    assign layer2_outputs[6531] = ~(layer1_outputs[11867]);
    assign layer2_outputs[6532] = 1'b1;
    assign layer2_outputs[6533] = ~(layer1_outputs[7310]);
    assign layer2_outputs[6534] = layer1_outputs[4313];
    assign layer2_outputs[6535] = (layer1_outputs[5630]) & ~(layer1_outputs[4437]);
    assign layer2_outputs[6536] = (layer1_outputs[6209]) ^ (layer1_outputs[9821]);
    assign layer2_outputs[6537] = ~(layer1_outputs[2722]);
    assign layer2_outputs[6538] = ~(layer1_outputs[76]);
    assign layer2_outputs[6539] = ~(layer1_outputs[9208]);
    assign layer2_outputs[6540] = ~((layer1_outputs[4235]) | (layer1_outputs[1868]));
    assign layer2_outputs[6541] = ~(layer1_outputs[4014]);
    assign layer2_outputs[6542] = ~(layer1_outputs[10299]);
    assign layer2_outputs[6543] = (layer1_outputs[860]) ^ (layer1_outputs[12586]);
    assign layer2_outputs[6544] = (layer1_outputs[4484]) ^ (layer1_outputs[6433]);
    assign layer2_outputs[6545] = ~(layer1_outputs[4097]);
    assign layer2_outputs[6546] = ~((layer1_outputs[11650]) ^ (layer1_outputs[12765]));
    assign layer2_outputs[6547] = (layer1_outputs[2174]) | (layer1_outputs[6968]);
    assign layer2_outputs[6548] = ~(layer1_outputs[11456]);
    assign layer2_outputs[6549] = ~((layer1_outputs[2438]) & (layer1_outputs[9322]));
    assign layer2_outputs[6550] = ~(layer1_outputs[7825]) | (layer1_outputs[3264]);
    assign layer2_outputs[6551] = (layer1_outputs[7581]) & (layer1_outputs[6095]);
    assign layer2_outputs[6552] = (layer1_outputs[11874]) & ~(layer1_outputs[1344]);
    assign layer2_outputs[6553] = ~(layer1_outputs[9487]);
    assign layer2_outputs[6554] = ~(layer1_outputs[3595]) | (layer1_outputs[5843]);
    assign layer2_outputs[6555] = ~(layer1_outputs[11010]);
    assign layer2_outputs[6556] = ~((layer1_outputs[1644]) ^ (layer1_outputs[4533]));
    assign layer2_outputs[6557] = ~((layer1_outputs[4435]) | (layer1_outputs[4963]));
    assign layer2_outputs[6558] = ~(layer1_outputs[5369]);
    assign layer2_outputs[6559] = layer1_outputs[4814];
    assign layer2_outputs[6560] = (layer1_outputs[10360]) & ~(layer1_outputs[604]);
    assign layer2_outputs[6561] = layer1_outputs[7161];
    assign layer2_outputs[6562] = (layer1_outputs[1204]) & (layer1_outputs[5669]);
    assign layer2_outputs[6563] = ~((layer1_outputs[5316]) & (layer1_outputs[1801]));
    assign layer2_outputs[6564] = ~(layer1_outputs[293]) | (layer1_outputs[1180]);
    assign layer2_outputs[6565] = ~(layer1_outputs[2904]);
    assign layer2_outputs[6566] = ~((layer1_outputs[11729]) | (layer1_outputs[557]));
    assign layer2_outputs[6567] = (layer1_outputs[8899]) & ~(layer1_outputs[537]);
    assign layer2_outputs[6568] = ~((layer1_outputs[5578]) & (layer1_outputs[8674]));
    assign layer2_outputs[6569] = ~((layer1_outputs[8215]) & (layer1_outputs[2780]));
    assign layer2_outputs[6570] = (layer1_outputs[890]) & ~(layer1_outputs[12425]);
    assign layer2_outputs[6571] = layer1_outputs[991];
    assign layer2_outputs[6572] = ~(layer1_outputs[9436]);
    assign layer2_outputs[6573] = layer1_outputs[4273];
    assign layer2_outputs[6574] = ~(layer1_outputs[10992]);
    assign layer2_outputs[6575] = ~(layer1_outputs[10511]) | (layer1_outputs[6838]);
    assign layer2_outputs[6576] = ~(layer1_outputs[7090]);
    assign layer2_outputs[6577] = ~((layer1_outputs[2389]) ^ (layer1_outputs[1717]));
    assign layer2_outputs[6578] = layer1_outputs[9371];
    assign layer2_outputs[6579] = layer1_outputs[10849];
    assign layer2_outputs[6580] = (layer1_outputs[7603]) ^ (layer1_outputs[3482]);
    assign layer2_outputs[6581] = ~(layer1_outputs[1863]);
    assign layer2_outputs[6582] = layer1_outputs[719];
    assign layer2_outputs[6583] = (layer1_outputs[12091]) & ~(layer1_outputs[1215]);
    assign layer2_outputs[6584] = ~(layer1_outputs[10514]);
    assign layer2_outputs[6585] = (layer1_outputs[2581]) & ~(layer1_outputs[7425]);
    assign layer2_outputs[6586] = ~(layer1_outputs[8888]) | (layer1_outputs[10914]);
    assign layer2_outputs[6587] = layer1_outputs[10866];
    assign layer2_outputs[6588] = ~(layer1_outputs[8196]);
    assign layer2_outputs[6589] = ~((layer1_outputs[11936]) ^ (layer1_outputs[6182]));
    assign layer2_outputs[6590] = 1'b1;
    assign layer2_outputs[6591] = ~(layer1_outputs[9116]);
    assign layer2_outputs[6592] = layer1_outputs[5070];
    assign layer2_outputs[6593] = layer1_outputs[2861];
    assign layer2_outputs[6594] = (layer1_outputs[9428]) & ~(layer1_outputs[9470]);
    assign layer2_outputs[6595] = ~(layer1_outputs[8606]);
    assign layer2_outputs[6596] = layer1_outputs[6730];
    assign layer2_outputs[6597] = ~(layer1_outputs[3455]);
    assign layer2_outputs[6598] = (layer1_outputs[9466]) & (layer1_outputs[426]);
    assign layer2_outputs[6599] = layer1_outputs[9823];
    assign layer2_outputs[6600] = ~((layer1_outputs[2168]) ^ (layer1_outputs[9895]));
    assign layer2_outputs[6601] = (layer1_outputs[5606]) & ~(layer1_outputs[6907]);
    assign layer2_outputs[6602] = (layer1_outputs[11674]) ^ (layer1_outputs[7722]);
    assign layer2_outputs[6603] = layer1_outputs[22];
    assign layer2_outputs[6604] = (layer1_outputs[8034]) | (layer1_outputs[10499]);
    assign layer2_outputs[6605] = (layer1_outputs[6823]) | (layer1_outputs[10783]);
    assign layer2_outputs[6606] = layer1_outputs[11137];
    assign layer2_outputs[6607] = (layer1_outputs[9095]) & ~(layer1_outputs[7792]);
    assign layer2_outputs[6608] = ~((layer1_outputs[3808]) ^ (layer1_outputs[10718]));
    assign layer2_outputs[6609] = layer1_outputs[12293];
    assign layer2_outputs[6610] = ~((layer1_outputs[8622]) ^ (layer1_outputs[2823]));
    assign layer2_outputs[6611] = ~((layer1_outputs[5308]) & (layer1_outputs[2172]));
    assign layer2_outputs[6612] = (layer1_outputs[11393]) ^ (layer1_outputs[9757]);
    assign layer2_outputs[6613] = ~((layer1_outputs[7952]) | (layer1_outputs[11387]));
    assign layer2_outputs[6614] = layer1_outputs[6210];
    assign layer2_outputs[6615] = ~(layer1_outputs[1357]);
    assign layer2_outputs[6616] = ~(layer1_outputs[3792]);
    assign layer2_outputs[6617] = layer1_outputs[4033];
    assign layer2_outputs[6618] = (layer1_outputs[1113]) & (layer1_outputs[7773]);
    assign layer2_outputs[6619] = layer1_outputs[7180];
    assign layer2_outputs[6620] = (layer1_outputs[10064]) & ~(layer1_outputs[8238]);
    assign layer2_outputs[6621] = (layer1_outputs[10580]) ^ (layer1_outputs[7670]);
    assign layer2_outputs[6622] = (layer1_outputs[4100]) & (layer1_outputs[7973]);
    assign layer2_outputs[6623] = ~(layer1_outputs[8764]);
    assign layer2_outputs[6624] = layer1_outputs[11000];
    assign layer2_outputs[6625] = ~(layer1_outputs[142]);
    assign layer2_outputs[6626] = layer1_outputs[6866];
    assign layer2_outputs[6627] = (layer1_outputs[4209]) ^ (layer1_outputs[5799]);
    assign layer2_outputs[6628] = ~(layer1_outputs[994]);
    assign layer2_outputs[6629] = ~((layer1_outputs[5562]) ^ (layer1_outputs[139]));
    assign layer2_outputs[6630] = layer1_outputs[8765];
    assign layer2_outputs[6631] = layer1_outputs[3642];
    assign layer2_outputs[6632] = ~(layer1_outputs[2460]);
    assign layer2_outputs[6633] = (layer1_outputs[11908]) | (layer1_outputs[10193]);
    assign layer2_outputs[6634] = layer1_outputs[8967];
    assign layer2_outputs[6635] = layer1_outputs[77];
    assign layer2_outputs[6636] = layer1_outputs[2243];
    assign layer2_outputs[6637] = layer1_outputs[5966];
    assign layer2_outputs[6638] = ~(layer1_outputs[6910]);
    assign layer2_outputs[6639] = ~((layer1_outputs[2476]) & (layer1_outputs[9450]));
    assign layer2_outputs[6640] = ~(layer1_outputs[8939]);
    assign layer2_outputs[6641] = (layer1_outputs[6560]) ^ (layer1_outputs[12519]);
    assign layer2_outputs[6642] = (layer1_outputs[1919]) & ~(layer1_outputs[8454]);
    assign layer2_outputs[6643] = layer1_outputs[9237];
    assign layer2_outputs[6644] = (layer1_outputs[3752]) & ~(layer1_outputs[7073]);
    assign layer2_outputs[6645] = layer1_outputs[11837];
    assign layer2_outputs[6646] = ~(layer1_outputs[4744]);
    assign layer2_outputs[6647] = ~(layer1_outputs[8989]) | (layer1_outputs[1223]);
    assign layer2_outputs[6648] = (layer1_outputs[6140]) | (layer1_outputs[9905]);
    assign layer2_outputs[6649] = ~((layer1_outputs[6227]) | (layer1_outputs[11988]));
    assign layer2_outputs[6650] = layer1_outputs[3022];
    assign layer2_outputs[6651] = layer1_outputs[4120];
    assign layer2_outputs[6652] = (layer1_outputs[6668]) | (layer1_outputs[6975]);
    assign layer2_outputs[6653] = (layer1_outputs[6574]) & (layer1_outputs[9982]);
    assign layer2_outputs[6654] = ~((layer1_outputs[643]) ^ (layer1_outputs[10612]));
    assign layer2_outputs[6655] = (layer1_outputs[10178]) & ~(layer1_outputs[8390]);
    assign layer2_outputs[6656] = ~(layer1_outputs[11973]);
    assign layer2_outputs[6657] = layer1_outputs[1942];
    assign layer2_outputs[6658] = layer1_outputs[8407];
    assign layer2_outputs[6659] = ~(layer1_outputs[4358]);
    assign layer2_outputs[6660] = ~((layer1_outputs[6807]) ^ (layer1_outputs[1251]));
    assign layer2_outputs[6661] = layer1_outputs[12211];
    assign layer2_outputs[6662] = ~(layer1_outputs[9628]);
    assign layer2_outputs[6663] = (layer1_outputs[11312]) & ~(layer1_outputs[9238]);
    assign layer2_outputs[6664] = ~(layer1_outputs[8037]);
    assign layer2_outputs[6665] = layer1_outputs[4864];
    assign layer2_outputs[6666] = (layer1_outputs[6953]) ^ (layer1_outputs[4901]);
    assign layer2_outputs[6667] = layer1_outputs[6019];
    assign layer2_outputs[6668] = ~(layer1_outputs[773]);
    assign layer2_outputs[6669] = (layer1_outputs[10471]) | (layer1_outputs[429]);
    assign layer2_outputs[6670] = ~(layer1_outputs[12704]);
    assign layer2_outputs[6671] = ~((layer1_outputs[10097]) | (layer1_outputs[9558]));
    assign layer2_outputs[6672] = layer1_outputs[2765];
    assign layer2_outputs[6673] = ~(layer1_outputs[4703]);
    assign layer2_outputs[6674] = (layer1_outputs[8081]) & ~(layer1_outputs[6448]);
    assign layer2_outputs[6675] = ~(layer1_outputs[3159]) | (layer1_outputs[4347]);
    assign layer2_outputs[6676] = layer1_outputs[3849];
    assign layer2_outputs[6677] = ~((layer1_outputs[5286]) ^ (layer1_outputs[2086]));
    assign layer2_outputs[6678] = layer1_outputs[4368];
    assign layer2_outputs[6679] = ~((layer1_outputs[2568]) ^ (layer1_outputs[8971]));
    assign layer2_outputs[6680] = ~(layer1_outputs[11531]) | (layer1_outputs[7843]);
    assign layer2_outputs[6681] = layer1_outputs[2406];
    assign layer2_outputs[6682] = ~(layer1_outputs[2157]);
    assign layer2_outputs[6683] = ~(layer1_outputs[5711]);
    assign layer2_outputs[6684] = ~(layer1_outputs[10856]);
    assign layer2_outputs[6685] = layer1_outputs[7983];
    assign layer2_outputs[6686] = layer1_outputs[419];
    assign layer2_outputs[6687] = ~(layer1_outputs[6798]);
    assign layer2_outputs[6688] = ~(layer1_outputs[12471]);
    assign layer2_outputs[6689] = layer1_outputs[11626];
    assign layer2_outputs[6690] = layer1_outputs[4454];
    assign layer2_outputs[6691] = layer1_outputs[1322];
    assign layer2_outputs[6692] = ~(layer1_outputs[8461]) | (layer1_outputs[11992]);
    assign layer2_outputs[6693] = ~((layer1_outputs[5005]) | (layer1_outputs[1823]));
    assign layer2_outputs[6694] = ~(layer1_outputs[8388]) | (layer1_outputs[7964]);
    assign layer2_outputs[6695] = (layer1_outputs[5108]) ^ (layer1_outputs[12618]);
    assign layer2_outputs[6696] = ~((layer1_outputs[4071]) & (layer1_outputs[6863]));
    assign layer2_outputs[6697] = ~((layer1_outputs[12026]) ^ (layer1_outputs[10434]));
    assign layer2_outputs[6698] = ~(layer1_outputs[12050]);
    assign layer2_outputs[6699] = ~(layer1_outputs[6154]);
    assign layer2_outputs[6700] = ~(layer1_outputs[12495]);
    assign layer2_outputs[6701] = 1'b1;
    assign layer2_outputs[6702] = layer1_outputs[345];
    assign layer2_outputs[6703] = ~((layer1_outputs[6461]) | (layer1_outputs[2871]));
    assign layer2_outputs[6704] = ~(layer1_outputs[4511]);
    assign layer2_outputs[6705] = (layer1_outputs[601]) & ~(layer1_outputs[11220]);
    assign layer2_outputs[6706] = layer1_outputs[1409];
    assign layer2_outputs[6707] = 1'b0;
    assign layer2_outputs[6708] = layer1_outputs[8245];
    assign layer2_outputs[6709] = (layer1_outputs[8636]) & (layer1_outputs[10714]);
    assign layer2_outputs[6710] = ~(layer1_outputs[2585]) | (layer1_outputs[12728]);
    assign layer2_outputs[6711] = layer1_outputs[11325];
    assign layer2_outputs[6712] = (layer1_outputs[3187]) & (layer1_outputs[2811]);
    assign layer2_outputs[6713] = layer1_outputs[3058];
    assign layer2_outputs[6714] = ~(layer1_outputs[1955]);
    assign layer2_outputs[6715] = ~(layer1_outputs[11608]);
    assign layer2_outputs[6716] = ~((layer1_outputs[5753]) ^ (layer1_outputs[166]));
    assign layer2_outputs[6717] = layer1_outputs[7847];
    assign layer2_outputs[6718] = ~((layer1_outputs[3050]) & (layer1_outputs[9036]));
    assign layer2_outputs[6719] = ~(layer1_outputs[2298]);
    assign layer2_outputs[6720] = ~((layer1_outputs[6597]) ^ (layer1_outputs[8995]));
    assign layer2_outputs[6721] = 1'b0;
    assign layer2_outputs[6722] = layer1_outputs[9318];
    assign layer2_outputs[6723] = layer1_outputs[5361];
    assign layer2_outputs[6724] = ~(layer1_outputs[1223]);
    assign layer2_outputs[6725] = layer1_outputs[8611];
    assign layer2_outputs[6726] = layer1_outputs[250];
    assign layer2_outputs[6727] = 1'b1;
    assign layer2_outputs[6728] = ~(layer1_outputs[9768]);
    assign layer2_outputs[6729] = (layer1_outputs[8632]) & ~(layer1_outputs[5320]);
    assign layer2_outputs[6730] = (layer1_outputs[7262]) ^ (layer1_outputs[11564]);
    assign layer2_outputs[6731] = layer1_outputs[1677];
    assign layer2_outputs[6732] = ~(layer1_outputs[8232]);
    assign layer2_outputs[6733] = ~(layer1_outputs[6792]);
    assign layer2_outputs[6734] = layer1_outputs[991];
    assign layer2_outputs[6735] = layer1_outputs[12533];
    assign layer2_outputs[6736] = layer1_outputs[10836];
    assign layer2_outputs[6737] = ~((layer1_outputs[2011]) | (layer1_outputs[11513]));
    assign layer2_outputs[6738] = ~((layer1_outputs[9418]) ^ (layer1_outputs[6617]));
    assign layer2_outputs[6739] = (layer1_outputs[2321]) & ~(layer1_outputs[6056]);
    assign layer2_outputs[6740] = ~((layer1_outputs[11740]) & (layer1_outputs[525]));
    assign layer2_outputs[6741] = ~((layer1_outputs[8710]) & (layer1_outputs[5646]));
    assign layer2_outputs[6742] = layer1_outputs[8159];
    assign layer2_outputs[6743] = ~((layer1_outputs[10671]) & (layer1_outputs[12706]));
    assign layer2_outputs[6744] = layer1_outputs[9712];
    assign layer2_outputs[6745] = ~((layer1_outputs[12730]) ^ (layer1_outputs[2452]));
    assign layer2_outputs[6746] = (layer1_outputs[4476]) | (layer1_outputs[9611]);
    assign layer2_outputs[6747] = layer1_outputs[12571];
    assign layer2_outputs[6748] = ~((layer1_outputs[10131]) ^ (layer1_outputs[4102]));
    assign layer2_outputs[6749] = ~(layer1_outputs[5436]) | (layer1_outputs[6216]);
    assign layer2_outputs[6750] = ~(layer1_outputs[5967]);
    assign layer2_outputs[6751] = layer1_outputs[10217];
    assign layer2_outputs[6752] = ~(layer1_outputs[220]);
    assign layer2_outputs[6753] = ~(layer1_outputs[9081]);
    assign layer2_outputs[6754] = ~(layer1_outputs[851]) | (layer1_outputs[3669]);
    assign layer2_outputs[6755] = ~((layer1_outputs[8219]) | (layer1_outputs[12423]));
    assign layer2_outputs[6756] = (layer1_outputs[8598]) & ~(layer1_outputs[6302]);
    assign layer2_outputs[6757] = (layer1_outputs[12002]) | (layer1_outputs[276]);
    assign layer2_outputs[6758] = layer1_outputs[6536];
    assign layer2_outputs[6759] = (layer1_outputs[5759]) ^ (layer1_outputs[9848]);
    assign layer2_outputs[6760] = layer1_outputs[3275];
    assign layer2_outputs[6761] = ~((layer1_outputs[9412]) ^ (layer1_outputs[5512]));
    assign layer2_outputs[6762] = layer1_outputs[10128];
    assign layer2_outputs[6763] = ~(layer1_outputs[752]);
    assign layer2_outputs[6764] = layer1_outputs[7021];
    assign layer2_outputs[6765] = ~(layer1_outputs[4005]);
    assign layer2_outputs[6766] = ~(layer1_outputs[791]);
    assign layer2_outputs[6767] = ~((layer1_outputs[1948]) & (layer1_outputs[2868]));
    assign layer2_outputs[6768] = layer1_outputs[9472];
    assign layer2_outputs[6769] = (layer1_outputs[7855]) & (layer1_outputs[5446]);
    assign layer2_outputs[6770] = ~((layer1_outputs[3196]) ^ (layer1_outputs[4901]));
    assign layer2_outputs[6771] = (layer1_outputs[484]) ^ (layer1_outputs[6336]);
    assign layer2_outputs[6772] = layer1_outputs[11873];
    assign layer2_outputs[6773] = ~((layer1_outputs[10648]) ^ (layer1_outputs[1342]));
    assign layer2_outputs[6774] = ~(layer1_outputs[1762]);
    assign layer2_outputs[6775] = (layer1_outputs[6748]) & (layer1_outputs[12774]);
    assign layer2_outputs[6776] = ~(layer1_outputs[722]);
    assign layer2_outputs[6777] = (layer1_outputs[5696]) & (layer1_outputs[10791]);
    assign layer2_outputs[6778] = layer1_outputs[12556];
    assign layer2_outputs[6779] = layer1_outputs[4978];
    assign layer2_outputs[6780] = (layer1_outputs[8328]) & (layer1_outputs[9228]);
    assign layer2_outputs[6781] = ~(layer1_outputs[111]);
    assign layer2_outputs[6782] = ~(layer1_outputs[11330]);
    assign layer2_outputs[6783] = ~((layer1_outputs[10636]) ^ (layer1_outputs[7266]));
    assign layer2_outputs[6784] = ~(layer1_outputs[7392]);
    assign layer2_outputs[6785] = layer1_outputs[10405];
    assign layer2_outputs[6786] = ~(layer1_outputs[7440]);
    assign layer2_outputs[6787] = ~((layer1_outputs[11076]) | (layer1_outputs[10310]));
    assign layer2_outputs[6788] = (layer1_outputs[6619]) & ~(layer1_outputs[10117]);
    assign layer2_outputs[6789] = ~(layer1_outputs[5253]) | (layer1_outputs[5252]);
    assign layer2_outputs[6790] = layer1_outputs[10736];
    assign layer2_outputs[6791] = layer1_outputs[8566];
    assign layer2_outputs[6792] = (layer1_outputs[5485]) | (layer1_outputs[3073]);
    assign layer2_outputs[6793] = (layer1_outputs[398]) & (layer1_outputs[2991]);
    assign layer2_outputs[6794] = ~(layer1_outputs[986]);
    assign layer2_outputs[6795] = (layer1_outputs[3096]) & ~(layer1_outputs[5245]);
    assign layer2_outputs[6796] = layer1_outputs[1982];
    assign layer2_outputs[6797] = layer1_outputs[7975];
    assign layer2_outputs[6798] = ~((layer1_outputs[1731]) & (layer1_outputs[12730]));
    assign layer2_outputs[6799] = (layer1_outputs[2512]) | (layer1_outputs[1489]);
    assign layer2_outputs[6800] = ~(layer1_outputs[3162]) | (layer1_outputs[9974]);
    assign layer2_outputs[6801] = (layer1_outputs[12569]) | (layer1_outputs[11819]);
    assign layer2_outputs[6802] = ~(layer1_outputs[8892]) | (layer1_outputs[9780]);
    assign layer2_outputs[6803] = layer1_outputs[7640];
    assign layer2_outputs[6804] = ~(layer1_outputs[10482]);
    assign layer2_outputs[6805] = (layer1_outputs[4089]) ^ (layer1_outputs[8488]);
    assign layer2_outputs[6806] = layer1_outputs[1481];
    assign layer2_outputs[6807] = layer1_outputs[5835];
    assign layer2_outputs[6808] = ~(layer1_outputs[6340]);
    assign layer2_outputs[6809] = ~(layer1_outputs[6231]);
    assign layer2_outputs[6810] = ~((layer1_outputs[4542]) ^ (layer1_outputs[6348]));
    assign layer2_outputs[6811] = ~(layer1_outputs[2409]);
    assign layer2_outputs[6812] = ~(layer1_outputs[12644]);
    assign layer2_outputs[6813] = ~(layer1_outputs[83]);
    assign layer2_outputs[6814] = ~((layer1_outputs[8901]) ^ (layer1_outputs[5874]));
    assign layer2_outputs[6815] = ~((layer1_outputs[12493]) | (layer1_outputs[2156]));
    assign layer2_outputs[6816] = (layer1_outputs[118]) & ~(layer1_outputs[3239]);
    assign layer2_outputs[6817] = (layer1_outputs[765]) ^ (layer1_outputs[7993]);
    assign layer2_outputs[6818] = layer1_outputs[6539];
    assign layer2_outputs[6819] = ~(layer1_outputs[9381]);
    assign layer2_outputs[6820] = layer1_outputs[271];
    assign layer2_outputs[6821] = ~((layer1_outputs[5668]) ^ (layer1_outputs[7446]));
    assign layer2_outputs[6822] = ~(layer1_outputs[7696]);
    assign layer2_outputs[6823] = ~((layer1_outputs[9396]) & (layer1_outputs[10934]));
    assign layer2_outputs[6824] = ~(layer1_outputs[10703]);
    assign layer2_outputs[6825] = ~((layer1_outputs[5595]) | (layer1_outputs[8045]));
    assign layer2_outputs[6826] = layer1_outputs[8068];
    assign layer2_outputs[6827] = (layer1_outputs[683]) ^ (layer1_outputs[9024]);
    assign layer2_outputs[6828] = layer1_outputs[11402];
    assign layer2_outputs[6829] = ~(layer1_outputs[6650]);
    assign layer2_outputs[6830] = (layer1_outputs[2446]) & (layer1_outputs[455]);
    assign layer2_outputs[6831] = ~((layer1_outputs[4050]) & (layer1_outputs[8311]));
    assign layer2_outputs[6832] = ~(layer1_outputs[11625]);
    assign layer2_outputs[6833] = ~((layer1_outputs[4844]) ^ (layer1_outputs[12303]));
    assign layer2_outputs[6834] = ~(layer1_outputs[4505]);
    assign layer2_outputs[6835] = layer1_outputs[5472];
    assign layer2_outputs[6836] = ~((layer1_outputs[9571]) ^ (layer1_outputs[8206]));
    assign layer2_outputs[6837] = ~(layer1_outputs[1118]);
    assign layer2_outputs[6838] = ~(layer1_outputs[10807]);
    assign layer2_outputs[6839] = ~(layer1_outputs[5051]);
    assign layer2_outputs[6840] = ~(layer1_outputs[8755]);
    assign layer2_outputs[6841] = (layer1_outputs[4021]) ^ (layer1_outputs[6595]);
    assign layer2_outputs[6842] = (layer1_outputs[9375]) | (layer1_outputs[6347]);
    assign layer2_outputs[6843] = layer1_outputs[9925];
    assign layer2_outputs[6844] = ~((layer1_outputs[1628]) & (layer1_outputs[7681]));
    assign layer2_outputs[6845] = ~(layer1_outputs[9137]);
    assign layer2_outputs[6846] = ~((layer1_outputs[1926]) & (layer1_outputs[9800]));
    assign layer2_outputs[6847] = layer1_outputs[7673];
    assign layer2_outputs[6848] = layer1_outputs[9442];
    assign layer2_outputs[6849] = ~(layer1_outputs[5075]);
    assign layer2_outputs[6850] = (layer1_outputs[9483]) ^ (layer1_outputs[11286]);
    assign layer2_outputs[6851] = layer1_outputs[9715];
    assign layer2_outputs[6852] = (layer1_outputs[5464]) & (layer1_outputs[9391]);
    assign layer2_outputs[6853] = ~(layer1_outputs[4472]) | (layer1_outputs[8840]);
    assign layer2_outputs[6854] = ~(layer1_outputs[3851]);
    assign layer2_outputs[6855] = layer1_outputs[11451];
    assign layer2_outputs[6856] = (layer1_outputs[7522]) | (layer1_outputs[3177]);
    assign layer2_outputs[6857] = layer1_outputs[5734];
    assign layer2_outputs[6858] = ~(layer1_outputs[618]);
    assign layer2_outputs[6859] = ~(layer1_outputs[5443]);
    assign layer2_outputs[6860] = ~(layer1_outputs[4515]);
    assign layer2_outputs[6861] = ~((layer1_outputs[9094]) & (layer1_outputs[12471]));
    assign layer2_outputs[6862] = layer1_outputs[6148];
    assign layer2_outputs[6863] = layer1_outputs[1445];
    assign layer2_outputs[6864] = ~(layer1_outputs[12521]);
    assign layer2_outputs[6865] = (layer1_outputs[8092]) | (layer1_outputs[458]);
    assign layer2_outputs[6866] = ~(layer1_outputs[184]);
    assign layer2_outputs[6867] = (layer1_outputs[8610]) & ~(layer1_outputs[4942]);
    assign layer2_outputs[6868] = (layer1_outputs[7296]) & ~(layer1_outputs[4312]);
    assign layer2_outputs[6869] = (layer1_outputs[12111]) | (layer1_outputs[8894]);
    assign layer2_outputs[6870] = ~(layer1_outputs[2328]) | (layer1_outputs[5914]);
    assign layer2_outputs[6871] = layer1_outputs[10783];
    assign layer2_outputs[6872] = ~(layer1_outputs[10699]) | (layer1_outputs[6653]);
    assign layer2_outputs[6873] = ~(layer1_outputs[5850]);
    assign layer2_outputs[6874] = ~((layer1_outputs[5958]) & (layer1_outputs[1396]));
    assign layer2_outputs[6875] = ~(layer1_outputs[11786]) | (layer1_outputs[6504]);
    assign layer2_outputs[6876] = layer1_outputs[11819];
    assign layer2_outputs[6877] = ~(layer1_outputs[1163]) | (layer1_outputs[1871]);
    assign layer2_outputs[6878] = (layer1_outputs[4253]) & (layer1_outputs[12322]);
    assign layer2_outputs[6879] = ~(layer1_outputs[9488]);
    assign layer2_outputs[6880] = ~(layer1_outputs[5935]);
    assign layer2_outputs[6881] = layer1_outputs[2787];
    assign layer2_outputs[6882] = ~(layer1_outputs[8515]);
    assign layer2_outputs[6883] = ~(layer1_outputs[6240]) | (layer1_outputs[11348]);
    assign layer2_outputs[6884] = ~(layer1_outputs[8015]) | (layer1_outputs[12073]);
    assign layer2_outputs[6885] = ~(layer1_outputs[2126]) | (layer1_outputs[3192]);
    assign layer2_outputs[6886] = layer1_outputs[10815];
    assign layer2_outputs[6887] = ~(layer1_outputs[10786]);
    assign layer2_outputs[6888] = ~(layer1_outputs[5659]) | (layer1_outputs[3399]);
    assign layer2_outputs[6889] = ~((layer1_outputs[5042]) & (layer1_outputs[7700]));
    assign layer2_outputs[6890] = ~((layer1_outputs[5356]) ^ (layer1_outputs[553]));
    assign layer2_outputs[6891] = ~(layer1_outputs[1093]);
    assign layer2_outputs[6892] = (layer1_outputs[6952]) ^ (layer1_outputs[4583]);
    assign layer2_outputs[6893] = (layer1_outputs[692]) | (layer1_outputs[8961]);
    assign layer2_outputs[6894] = ~(layer1_outputs[6959]);
    assign layer2_outputs[6895] = layer1_outputs[2748];
    assign layer2_outputs[6896] = (layer1_outputs[7886]) ^ (layer1_outputs[8934]);
    assign layer2_outputs[6897] = (layer1_outputs[12125]) & ~(layer1_outputs[3698]);
    assign layer2_outputs[6898] = layer1_outputs[6002];
    assign layer2_outputs[6899] = ~(layer1_outputs[10464]);
    assign layer2_outputs[6900] = (layer1_outputs[6398]) & ~(layer1_outputs[3918]);
    assign layer2_outputs[6901] = layer1_outputs[9941];
    assign layer2_outputs[6902] = ~((layer1_outputs[6899]) & (layer1_outputs[9109]));
    assign layer2_outputs[6903] = layer1_outputs[4230];
    assign layer2_outputs[6904] = ~((layer1_outputs[5590]) ^ (layer1_outputs[7426]));
    assign layer2_outputs[6905] = ~(layer1_outputs[4153]);
    assign layer2_outputs[6906] = (layer1_outputs[10499]) & ~(layer1_outputs[7843]);
    assign layer2_outputs[6907] = layer1_outputs[3238];
    assign layer2_outputs[6908] = (layer1_outputs[3739]) | (layer1_outputs[9777]);
    assign layer2_outputs[6909] = ~(layer1_outputs[7223]);
    assign layer2_outputs[6910] = layer1_outputs[2948];
    assign layer2_outputs[6911] = ~(layer1_outputs[6660]);
    assign layer2_outputs[6912] = ~((layer1_outputs[7846]) ^ (layer1_outputs[4249]));
    assign layer2_outputs[6913] = ~((layer1_outputs[11234]) & (layer1_outputs[1705]));
    assign layer2_outputs[6914] = layer1_outputs[1439];
    assign layer2_outputs[6915] = layer1_outputs[3195];
    assign layer2_outputs[6916] = ~(layer1_outputs[5483]);
    assign layer2_outputs[6917] = ~(layer1_outputs[5267]);
    assign layer2_outputs[6918] = layer1_outputs[7544];
    assign layer2_outputs[6919] = layer1_outputs[751];
    assign layer2_outputs[6920] = ~(layer1_outputs[6189]);
    assign layer2_outputs[6921] = ~(layer1_outputs[6103]) | (layer1_outputs[12308]);
    assign layer2_outputs[6922] = ~(layer1_outputs[7166]) | (layer1_outputs[1561]);
    assign layer2_outputs[6923] = (layer1_outputs[3348]) | (layer1_outputs[4143]);
    assign layer2_outputs[6924] = layer1_outputs[9999];
    assign layer2_outputs[6925] = layer1_outputs[4221];
    assign layer2_outputs[6926] = layer1_outputs[12221];
    assign layer2_outputs[6927] = ~(layer1_outputs[8006]);
    assign layer2_outputs[6928] = ~(layer1_outputs[2888]);
    assign layer2_outputs[6929] = (layer1_outputs[6839]) & (layer1_outputs[4025]);
    assign layer2_outputs[6930] = ~(layer1_outputs[12531]);
    assign layer2_outputs[6931] = (layer1_outputs[11297]) | (layer1_outputs[9599]);
    assign layer2_outputs[6932] = (layer1_outputs[10917]) & ~(layer1_outputs[8535]);
    assign layer2_outputs[6933] = ~(layer1_outputs[9008]);
    assign layer2_outputs[6934] = (layer1_outputs[7293]) & (layer1_outputs[70]);
    assign layer2_outputs[6935] = ~(layer1_outputs[11886]);
    assign layer2_outputs[6936] = ~((layer1_outputs[2611]) & (layer1_outputs[2480]));
    assign layer2_outputs[6937] = ~(layer1_outputs[7543]) | (layer1_outputs[11186]);
    assign layer2_outputs[6938] = ~(layer1_outputs[2894]);
    assign layer2_outputs[6939] = ~((layer1_outputs[8580]) | (layer1_outputs[6330]));
    assign layer2_outputs[6940] = layer1_outputs[3682];
    assign layer2_outputs[6941] = layer1_outputs[9641];
    assign layer2_outputs[6942] = layer1_outputs[7399];
    assign layer2_outputs[6943] = (layer1_outputs[7741]) & ~(layer1_outputs[9978]);
    assign layer2_outputs[6944] = ~((layer1_outputs[7743]) | (layer1_outputs[4626]));
    assign layer2_outputs[6945] = ~(layer1_outputs[11711]) | (layer1_outputs[10197]);
    assign layer2_outputs[6946] = ~(layer1_outputs[11408]);
    assign layer2_outputs[6947] = (layer1_outputs[9212]) & (layer1_outputs[11180]);
    assign layer2_outputs[6948] = layer1_outputs[9918];
    assign layer2_outputs[6949] = layer1_outputs[12413];
    assign layer2_outputs[6950] = (layer1_outputs[11162]) | (layer1_outputs[11956]);
    assign layer2_outputs[6951] = ~(layer1_outputs[9088]);
    assign layer2_outputs[6952] = ~(layer1_outputs[9591]);
    assign layer2_outputs[6953] = ~((layer1_outputs[6755]) | (layer1_outputs[5813]));
    assign layer2_outputs[6954] = ~(layer1_outputs[555]);
    assign layer2_outputs[6955] = ~(layer1_outputs[4295]);
    assign layer2_outputs[6956] = (layer1_outputs[7297]) & ~(layer1_outputs[5648]);
    assign layer2_outputs[6957] = ~(layer1_outputs[7393]) | (layer1_outputs[7467]);
    assign layer2_outputs[6958] = ~(layer1_outputs[7881]) | (layer1_outputs[11930]);
    assign layer2_outputs[6959] = ~(layer1_outputs[7612]);
    assign layer2_outputs[6960] = layer1_outputs[1880];
    assign layer2_outputs[6961] = ~(layer1_outputs[8033]);
    assign layer2_outputs[6962] = ~(layer1_outputs[9202]);
    assign layer2_outputs[6963] = (layer1_outputs[1712]) & ~(layer1_outputs[11481]);
    assign layer2_outputs[6964] = ~(layer1_outputs[2048]);
    assign layer2_outputs[6965] = layer1_outputs[1084];
    assign layer2_outputs[6966] = ~((layer1_outputs[2138]) & (layer1_outputs[10408]));
    assign layer2_outputs[6967] = ~(layer1_outputs[8127]);
    assign layer2_outputs[6968] = (layer1_outputs[11623]) & (layer1_outputs[11022]);
    assign layer2_outputs[6969] = ~(layer1_outputs[10551]) | (layer1_outputs[12777]);
    assign layer2_outputs[6970] = ~(layer1_outputs[10743]) | (layer1_outputs[1650]);
    assign layer2_outputs[6971] = layer1_outputs[1838];
    assign layer2_outputs[6972] = (layer1_outputs[4976]) & ~(layer1_outputs[7241]);
    assign layer2_outputs[6973] = ~(layer1_outputs[11071]) | (layer1_outputs[3546]);
    assign layer2_outputs[6974] = ~(layer1_outputs[9523]);
    assign layer2_outputs[6975] = (layer1_outputs[3186]) | (layer1_outputs[8875]);
    assign layer2_outputs[6976] = layer1_outputs[10648];
    assign layer2_outputs[6977] = layer1_outputs[4277];
    assign layer2_outputs[6978] = (layer1_outputs[7839]) ^ (layer1_outputs[3468]);
    assign layer2_outputs[6979] = ~(layer1_outputs[1269]);
    assign layer2_outputs[6980] = ~((layer1_outputs[8369]) ^ (layer1_outputs[2713]));
    assign layer2_outputs[6981] = (layer1_outputs[10009]) & (layer1_outputs[1277]);
    assign layer2_outputs[6982] = ~((layer1_outputs[12434]) | (layer1_outputs[5960]));
    assign layer2_outputs[6983] = (layer1_outputs[4451]) & (layer1_outputs[2448]);
    assign layer2_outputs[6984] = (layer1_outputs[452]) & ~(layer1_outputs[9624]);
    assign layer2_outputs[6985] = ~((layer1_outputs[8815]) & (layer1_outputs[4584]));
    assign layer2_outputs[6986] = layer1_outputs[1054];
    assign layer2_outputs[6987] = ~(layer1_outputs[10789]);
    assign layer2_outputs[6988] = ~((layer1_outputs[8038]) & (layer1_outputs[632]));
    assign layer2_outputs[6989] = layer1_outputs[2916];
    assign layer2_outputs[6990] = ~(layer1_outputs[8399]);
    assign layer2_outputs[6991] = (layer1_outputs[3875]) & (layer1_outputs[6035]);
    assign layer2_outputs[6992] = layer1_outputs[3775];
    assign layer2_outputs[6993] = layer1_outputs[11032];
    assign layer2_outputs[6994] = layer1_outputs[6881];
    assign layer2_outputs[6995] = ~(layer1_outputs[3432]);
    assign layer2_outputs[6996] = (layer1_outputs[1692]) & (layer1_outputs[3922]);
    assign layer2_outputs[6997] = layer1_outputs[2725];
    assign layer2_outputs[6998] = layer1_outputs[4236];
    assign layer2_outputs[6999] = ~(layer1_outputs[10378]);
    assign layer2_outputs[7000] = ~(layer1_outputs[3792]);
    assign layer2_outputs[7001] = (layer1_outputs[7513]) & (layer1_outputs[1493]);
    assign layer2_outputs[7002] = layer1_outputs[950];
    assign layer2_outputs[7003] = (layer1_outputs[963]) ^ (layer1_outputs[8740]);
    assign layer2_outputs[7004] = (layer1_outputs[1529]) & ~(layer1_outputs[12080]);
    assign layer2_outputs[7005] = layer1_outputs[9191];
    assign layer2_outputs[7006] = layer1_outputs[8115];
    assign layer2_outputs[7007] = (layer1_outputs[11590]) | (layer1_outputs[12333]);
    assign layer2_outputs[7008] = ~(layer1_outputs[815]);
    assign layer2_outputs[7009] = layer1_outputs[12258];
    assign layer2_outputs[7010] = (layer1_outputs[5801]) & ~(layer1_outputs[4563]);
    assign layer2_outputs[7011] = (layer1_outputs[6332]) & (layer1_outputs[8208]);
    assign layer2_outputs[7012] = (layer1_outputs[12301]) & (layer1_outputs[4877]);
    assign layer2_outputs[7013] = (layer1_outputs[995]) & ~(layer1_outputs[4077]);
    assign layer2_outputs[7014] = layer1_outputs[10334];
    assign layer2_outputs[7015] = (layer1_outputs[7254]) & ~(layer1_outputs[4152]);
    assign layer2_outputs[7016] = ~(layer1_outputs[6163]);
    assign layer2_outputs[7017] = (layer1_outputs[2693]) & (layer1_outputs[6629]);
    assign layer2_outputs[7018] = layer1_outputs[3663];
    assign layer2_outputs[7019] = ~(layer1_outputs[2561]);
    assign layer2_outputs[7020] = (layer1_outputs[5524]) & (layer1_outputs[7668]);
    assign layer2_outputs[7021] = ~((layer1_outputs[12420]) & (layer1_outputs[8397]));
    assign layer2_outputs[7022] = ~(layer1_outputs[6624]);
    assign layer2_outputs[7023] = ~(layer1_outputs[3221]) | (layer1_outputs[9688]);
    assign layer2_outputs[7024] = ~((layer1_outputs[5778]) ^ (layer1_outputs[2647]));
    assign layer2_outputs[7025] = layer1_outputs[9220];
    assign layer2_outputs[7026] = ~((layer1_outputs[11875]) & (layer1_outputs[9585]));
    assign layer2_outputs[7027] = (layer1_outputs[3174]) & ~(layer1_outputs[4]);
    assign layer2_outputs[7028] = layer1_outputs[1073];
    assign layer2_outputs[7029] = (layer1_outputs[11661]) & ~(layer1_outputs[12566]);
    assign layer2_outputs[7030] = layer1_outputs[9489];
    assign layer2_outputs[7031] = ~((layer1_outputs[8230]) ^ (layer1_outputs[12474]));
    assign layer2_outputs[7032] = layer1_outputs[8191];
    assign layer2_outputs[7033] = (layer1_outputs[8940]) & (layer1_outputs[2714]);
    assign layer2_outputs[7034] = (layer1_outputs[7538]) | (layer1_outputs[9293]);
    assign layer2_outputs[7035] = ~((layer1_outputs[7374]) | (layer1_outputs[5803]));
    assign layer2_outputs[7036] = ~(layer1_outputs[3989]) | (layer1_outputs[7848]);
    assign layer2_outputs[7037] = layer1_outputs[811];
    assign layer2_outputs[7038] = ~(layer1_outputs[6061]);
    assign layer2_outputs[7039] = ~(layer1_outputs[9669]);
    assign layer2_outputs[7040] = (layer1_outputs[7845]) ^ (layer1_outputs[12389]);
    assign layer2_outputs[7041] = ~((layer1_outputs[2726]) & (layer1_outputs[3722]));
    assign layer2_outputs[7042] = ~(layer1_outputs[4744]);
    assign layer2_outputs[7043] = (layer1_outputs[3896]) & (layer1_outputs[1687]);
    assign layer2_outputs[7044] = layer1_outputs[9735];
    assign layer2_outputs[7045] = layer1_outputs[9715];
    assign layer2_outputs[7046] = ~((layer1_outputs[961]) & (layer1_outputs[4985]));
    assign layer2_outputs[7047] = ~((layer1_outputs[1640]) & (layer1_outputs[11412]));
    assign layer2_outputs[7048] = 1'b0;
    assign layer2_outputs[7049] = ~((layer1_outputs[7979]) | (layer1_outputs[1670]));
    assign layer2_outputs[7050] = ~(layer1_outputs[3106]);
    assign layer2_outputs[7051] = layer1_outputs[10164];
    assign layer2_outputs[7052] = ~(layer1_outputs[7411]);
    assign layer2_outputs[7053] = (layer1_outputs[9703]) & ~(layer1_outputs[9673]);
    assign layer2_outputs[7054] = (layer1_outputs[4399]) | (layer1_outputs[3342]);
    assign layer2_outputs[7055] = (layer1_outputs[9724]) ^ (layer1_outputs[9810]);
    assign layer2_outputs[7056] = layer1_outputs[10546];
    assign layer2_outputs[7057] = ~(layer1_outputs[9898]);
    assign layer2_outputs[7058] = ~(layer1_outputs[1235]);
    assign layer2_outputs[7059] = ~((layer1_outputs[3308]) ^ (layer1_outputs[11709]));
    assign layer2_outputs[7060] = ~(layer1_outputs[2576]);
    assign layer2_outputs[7061] = layer1_outputs[11054];
    assign layer2_outputs[7062] = layer1_outputs[8423];
    assign layer2_outputs[7063] = ~((layer1_outputs[4322]) ^ (layer1_outputs[8527]));
    assign layer2_outputs[7064] = ~((layer1_outputs[10000]) ^ (layer1_outputs[2985]));
    assign layer2_outputs[7065] = layer1_outputs[4586];
    assign layer2_outputs[7066] = ~((layer1_outputs[622]) ^ (layer1_outputs[6033]));
    assign layer2_outputs[7067] = (layer1_outputs[9415]) & ~(layer1_outputs[6556]);
    assign layer2_outputs[7068] = layer1_outputs[10260];
    assign layer2_outputs[7069] = ~((layer1_outputs[12174]) & (layer1_outputs[402]));
    assign layer2_outputs[7070] = layer1_outputs[8145];
    assign layer2_outputs[7071] = ~(layer1_outputs[6285]);
    assign layer2_outputs[7072] = ~(layer1_outputs[453]);
    assign layer2_outputs[7073] = (layer1_outputs[5238]) | (layer1_outputs[9816]);
    assign layer2_outputs[7074] = layer1_outputs[2268];
    assign layer2_outputs[7075] = layer1_outputs[743];
    assign layer2_outputs[7076] = (layer1_outputs[8022]) | (layer1_outputs[5737]);
    assign layer2_outputs[7077] = ~((layer1_outputs[8855]) | (layer1_outputs[7333]));
    assign layer2_outputs[7078] = layer1_outputs[3810];
    assign layer2_outputs[7079] = ~(layer1_outputs[3160]);
    assign layer2_outputs[7080] = (layer1_outputs[6421]) & (layer1_outputs[7551]);
    assign layer2_outputs[7081] = layer1_outputs[7996];
    assign layer2_outputs[7082] = ~(layer1_outputs[9199]) | (layer1_outputs[6939]);
    assign layer2_outputs[7083] = layer1_outputs[9208];
    assign layer2_outputs[7084] = (layer1_outputs[11373]) & (layer1_outputs[387]);
    assign layer2_outputs[7085] = (layer1_outputs[5216]) ^ (layer1_outputs[12537]);
    assign layer2_outputs[7086] = (layer1_outputs[6232]) ^ (layer1_outputs[1759]);
    assign layer2_outputs[7087] = (layer1_outputs[11638]) ^ (layer1_outputs[8427]);
    assign layer2_outputs[7088] = ~((layer1_outputs[7674]) | (layer1_outputs[12796]));
    assign layer2_outputs[7089] = (layer1_outputs[2219]) & ~(layer1_outputs[4164]);
    assign layer2_outputs[7090] = ~((layer1_outputs[11783]) | (layer1_outputs[9856]));
    assign layer2_outputs[7091] = layer1_outputs[11447];
    assign layer2_outputs[7092] = layer1_outputs[3824];
    assign layer2_outputs[7093] = ~((layer1_outputs[9687]) & (layer1_outputs[7572]));
    assign layer2_outputs[7094] = ~(layer1_outputs[3389]);
    assign layer2_outputs[7095] = ~((layer1_outputs[4724]) ^ (layer1_outputs[950]));
    assign layer2_outputs[7096] = (layer1_outputs[2765]) & ~(layer1_outputs[3433]);
    assign layer2_outputs[7097] = ~(layer1_outputs[5770]) | (layer1_outputs[1044]);
    assign layer2_outputs[7098] = ~(layer1_outputs[7782]) | (layer1_outputs[5608]);
    assign layer2_outputs[7099] = (layer1_outputs[6596]) & ~(layer1_outputs[10801]);
    assign layer2_outputs[7100] = layer1_outputs[8591];
    assign layer2_outputs[7101] = (layer1_outputs[11832]) | (layer1_outputs[7573]);
    assign layer2_outputs[7102] = layer1_outputs[10084];
    assign layer2_outputs[7103] = ~(layer1_outputs[11293]);
    assign layer2_outputs[7104] = layer1_outputs[7285];
    assign layer2_outputs[7105] = layer1_outputs[4735];
    assign layer2_outputs[7106] = ~(layer1_outputs[7155]);
    assign layer2_outputs[7107] = ~((layer1_outputs[12294]) | (layer1_outputs[1904]));
    assign layer2_outputs[7108] = ~((layer1_outputs[10131]) & (layer1_outputs[7964]));
    assign layer2_outputs[7109] = ~(layer1_outputs[12104]);
    assign layer2_outputs[7110] = ~(layer1_outputs[2906]);
    assign layer2_outputs[7111] = ~((layer1_outputs[10436]) ^ (layer1_outputs[10627]));
    assign layer2_outputs[7112] = layer1_outputs[46];
    assign layer2_outputs[7113] = layer1_outputs[10908];
    assign layer2_outputs[7114] = layer1_outputs[2356];
    assign layer2_outputs[7115] = layer1_outputs[8928];
    assign layer2_outputs[7116] = layer1_outputs[7336];
    assign layer2_outputs[7117] = ~(layer1_outputs[3265]) | (layer1_outputs[3951]);
    assign layer2_outputs[7118] = layer1_outputs[4758];
    assign layer2_outputs[7119] = ~(layer1_outputs[1581]);
    assign layer2_outputs[7120] = ~(layer1_outputs[10325]);
    assign layer2_outputs[7121] = ~(layer1_outputs[9916]) | (layer1_outputs[10874]);
    assign layer2_outputs[7122] = layer1_outputs[4804];
    assign layer2_outputs[7123] = (layer1_outputs[2365]) & ~(layer1_outputs[4987]);
    assign layer2_outputs[7124] = ~((layer1_outputs[10407]) ^ (layer1_outputs[766]));
    assign layer2_outputs[7125] = layer1_outputs[6978];
    assign layer2_outputs[7126] = ~(layer1_outputs[4535]);
    assign layer2_outputs[7127] = ~((layer1_outputs[9076]) | (layer1_outputs[8223]));
    assign layer2_outputs[7128] = (layer1_outputs[2154]) & ~(layer1_outputs[6429]);
    assign layer2_outputs[7129] = ~((layer1_outputs[9005]) & (layer1_outputs[11467]));
    assign layer2_outputs[7130] = ~(layer1_outputs[12199]);
    assign layer2_outputs[7131] = (layer1_outputs[11019]) & ~(layer1_outputs[11765]);
    assign layer2_outputs[7132] = (layer1_outputs[5316]) & ~(layer1_outputs[12695]);
    assign layer2_outputs[7133] = layer1_outputs[9469];
    assign layer2_outputs[7134] = ~(layer1_outputs[10433]);
    assign layer2_outputs[7135] = layer1_outputs[7063];
    assign layer2_outputs[7136] = ~(layer1_outputs[6454]);
    assign layer2_outputs[7137] = ~((layer1_outputs[223]) | (layer1_outputs[5698]));
    assign layer2_outputs[7138] = (layer1_outputs[3173]) ^ (layer1_outputs[2304]);
    assign layer2_outputs[7139] = ~(layer1_outputs[667]);
    assign layer2_outputs[7140] = layer1_outputs[10893];
    assign layer2_outputs[7141] = ~((layer1_outputs[11950]) ^ (layer1_outputs[9913]));
    assign layer2_outputs[7142] = (layer1_outputs[650]) ^ (layer1_outputs[8258]);
    assign layer2_outputs[7143] = ~(layer1_outputs[2450]);
    assign layer2_outputs[7144] = ~((layer1_outputs[12466]) | (layer1_outputs[8010]));
    assign layer2_outputs[7145] = ~((layer1_outputs[1650]) ^ (layer1_outputs[11860]));
    assign layer2_outputs[7146] = layer1_outputs[12714];
    assign layer2_outputs[7147] = (layer1_outputs[9349]) & ~(layer1_outputs[5247]);
    assign layer2_outputs[7148] = layer1_outputs[7008];
    assign layer2_outputs[7149] = (layer1_outputs[6852]) & (layer1_outputs[7327]);
    assign layer2_outputs[7150] = layer1_outputs[2317];
    assign layer2_outputs[7151] = ~(layer1_outputs[852]);
    assign layer2_outputs[7152] = (layer1_outputs[5797]) | (layer1_outputs[11520]);
    assign layer2_outputs[7153] = layer1_outputs[1485];
    assign layer2_outputs[7154] = (layer1_outputs[8779]) & ~(layer1_outputs[1220]);
    assign layer2_outputs[7155] = ~(layer1_outputs[2497]);
    assign layer2_outputs[7156] = ~((layer1_outputs[1413]) | (layer1_outputs[7910]));
    assign layer2_outputs[7157] = ~(layer1_outputs[714]);
    assign layer2_outputs[7158] = ~(layer1_outputs[3406]);
    assign layer2_outputs[7159] = 1'b1;
    assign layer2_outputs[7160] = ~(layer1_outputs[11977]);
    assign layer2_outputs[7161] = ~(layer1_outputs[680]) | (layer1_outputs[7695]);
    assign layer2_outputs[7162] = ~(layer1_outputs[7930]);
    assign layer2_outputs[7163] = (layer1_outputs[10202]) | (layer1_outputs[5678]);
    assign layer2_outputs[7164] = (layer1_outputs[3437]) ^ (layer1_outputs[10291]);
    assign layer2_outputs[7165] = (layer1_outputs[5358]) ^ (layer1_outputs[1196]);
    assign layer2_outputs[7166] = ~((layer1_outputs[2889]) | (layer1_outputs[5994]));
    assign layer2_outputs[7167] = ~((layer1_outputs[915]) | (layer1_outputs[10952]));
    assign layer2_outputs[7168] = ~((layer1_outputs[11878]) ^ (layer1_outputs[10612]));
    assign layer2_outputs[7169] = ~(layer1_outputs[8306]) | (layer1_outputs[4821]);
    assign layer2_outputs[7170] = layer1_outputs[9382];
    assign layer2_outputs[7171] = (layer1_outputs[10943]) & ~(layer1_outputs[10745]);
    assign layer2_outputs[7172] = ~((layer1_outputs[8688]) | (layer1_outputs[1485]));
    assign layer2_outputs[7173] = layer1_outputs[6902];
    assign layer2_outputs[7174] = (layer1_outputs[10240]) ^ (layer1_outputs[12224]);
    assign layer2_outputs[7175] = layer1_outputs[5743];
    assign layer2_outputs[7176] = ~((layer1_outputs[3333]) ^ (layer1_outputs[730]));
    assign layer2_outputs[7177] = layer1_outputs[10399];
    assign layer2_outputs[7178] = ~((layer1_outputs[2434]) | (layer1_outputs[608]));
    assign layer2_outputs[7179] = 1'b1;
    assign layer2_outputs[7180] = layer1_outputs[746];
    assign layer2_outputs[7181] = ~(layer1_outputs[9082]);
    assign layer2_outputs[7182] = ~((layer1_outputs[5556]) | (layer1_outputs[9250]));
    assign layer2_outputs[7183] = layer1_outputs[837];
    assign layer2_outputs[7184] = ~(layer1_outputs[4823]);
    assign layer2_outputs[7185] = layer1_outputs[3118];
    assign layer2_outputs[7186] = ~((layer1_outputs[5747]) ^ (layer1_outputs[2799]));
    assign layer2_outputs[7187] = ~(layer1_outputs[8263]);
    assign layer2_outputs[7188] = ~(layer1_outputs[9897]);
    assign layer2_outputs[7189] = ~(layer1_outputs[10409]);
    assign layer2_outputs[7190] = layer1_outputs[316];
    assign layer2_outputs[7191] = ~(layer1_outputs[8358]);
    assign layer2_outputs[7192] = ~((layer1_outputs[1535]) & (layer1_outputs[10169]));
    assign layer2_outputs[7193] = (layer1_outputs[3638]) & (layer1_outputs[4279]);
    assign layer2_outputs[7194] = (layer1_outputs[9338]) & ~(layer1_outputs[1920]);
    assign layer2_outputs[7195] = layer1_outputs[10691];
    assign layer2_outputs[7196] = (layer1_outputs[11118]) & ~(layer1_outputs[11351]);
    assign layer2_outputs[7197] = ~(layer1_outputs[120]);
    assign layer2_outputs[7198] = ~(layer1_outputs[985]) | (layer1_outputs[2206]);
    assign layer2_outputs[7199] = ~(layer1_outputs[12304]);
    assign layer2_outputs[7200] = ~((layer1_outputs[2866]) ^ (layer1_outputs[9853]));
    assign layer2_outputs[7201] = layer1_outputs[586];
    assign layer2_outputs[7202] = ~(layer1_outputs[6317]);
    assign layer2_outputs[7203] = ~(layer1_outputs[3245]);
    assign layer2_outputs[7204] = ~(layer1_outputs[8962]);
    assign layer2_outputs[7205] = ~(layer1_outputs[4242]) | (layer1_outputs[1104]);
    assign layer2_outputs[7206] = ~((layer1_outputs[11829]) & (layer1_outputs[11793]));
    assign layer2_outputs[7207] = ~(layer1_outputs[12534]);
    assign layer2_outputs[7208] = ~((layer1_outputs[2471]) & (layer1_outputs[5327]));
    assign layer2_outputs[7209] = (layer1_outputs[10066]) & ~(layer1_outputs[878]);
    assign layer2_outputs[7210] = ~((layer1_outputs[3020]) | (layer1_outputs[12015]));
    assign layer2_outputs[7211] = layer1_outputs[7420];
    assign layer2_outputs[7212] = ~(layer1_outputs[2089]);
    assign layer2_outputs[7213] = ~((layer1_outputs[8955]) | (layer1_outputs[5505]));
    assign layer2_outputs[7214] = (layer1_outputs[10757]) & (layer1_outputs[8550]);
    assign layer2_outputs[7215] = layer1_outputs[5900];
    assign layer2_outputs[7216] = layer1_outputs[11311];
    assign layer2_outputs[7217] = ~(layer1_outputs[7758]) | (layer1_outputs[8106]);
    assign layer2_outputs[7218] = ~((layer1_outputs[8710]) ^ (layer1_outputs[4786]));
    assign layer2_outputs[7219] = ~((layer1_outputs[9917]) & (layer1_outputs[562]));
    assign layer2_outputs[7220] = ~(layer1_outputs[5097]);
    assign layer2_outputs[7221] = layer1_outputs[3208];
    assign layer2_outputs[7222] = ~(layer1_outputs[1457]);
    assign layer2_outputs[7223] = ~(layer1_outputs[9203]);
    assign layer2_outputs[7224] = 1'b1;
    assign layer2_outputs[7225] = (layer1_outputs[8559]) ^ (layer1_outputs[11884]);
    assign layer2_outputs[7226] = ~(layer1_outputs[11212]);
    assign layer2_outputs[7227] = ~((layer1_outputs[3701]) | (layer1_outputs[9725]));
    assign layer2_outputs[7228] = (layer1_outputs[12740]) & ~(layer1_outputs[2124]);
    assign layer2_outputs[7229] = ~(layer1_outputs[3141]) | (layer1_outputs[3935]);
    assign layer2_outputs[7230] = layer1_outputs[2121];
    assign layer2_outputs[7231] = layer1_outputs[5365];
    assign layer2_outputs[7232] = ~((layer1_outputs[1448]) ^ (layer1_outputs[255]));
    assign layer2_outputs[7233] = ~((layer1_outputs[5336]) ^ (layer1_outputs[1519]));
    assign layer2_outputs[7234] = ~(layer1_outputs[4835]);
    assign layer2_outputs[7235] = ~(layer1_outputs[4659]);
    assign layer2_outputs[7236] = ~(layer1_outputs[7407]) | (layer1_outputs[9362]);
    assign layer2_outputs[7237] = (layer1_outputs[2809]) ^ (layer1_outputs[9877]);
    assign layer2_outputs[7238] = ~((layer1_outputs[1238]) ^ (layer1_outputs[10548]));
    assign layer2_outputs[7239] = ~(layer1_outputs[4082]);
    assign layer2_outputs[7240] = ~(layer1_outputs[12437]);
    assign layer2_outputs[7241] = ~(layer1_outputs[8552]);
    assign layer2_outputs[7242] = layer1_outputs[7492];
    assign layer2_outputs[7243] = ~(layer1_outputs[2858]) | (layer1_outputs[6171]);
    assign layer2_outputs[7244] = ~(layer1_outputs[4772]) | (layer1_outputs[6180]);
    assign layer2_outputs[7245] = (layer1_outputs[5868]) & ~(layer1_outputs[10134]);
    assign layer2_outputs[7246] = ~(layer1_outputs[2480]);
    assign layer2_outputs[7247] = ~(layer1_outputs[8977]) | (layer1_outputs[7096]);
    assign layer2_outputs[7248] = (layer1_outputs[11718]) & (layer1_outputs[7200]);
    assign layer2_outputs[7249] = ~((layer1_outputs[8569]) | (layer1_outputs[5913]));
    assign layer2_outputs[7250] = (layer1_outputs[3269]) & ~(layer1_outputs[6955]);
    assign layer2_outputs[7251] = ~((layer1_outputs[5003]) ^ (layer1_outputs[417]));
    assign layer2_outputs[7252] = ~(layer1_outputs[11978]) | (layer1_outputs[12299]);
    assign layer2_outputs[7253] = ~(layer1_outputs[6338]);
    assign layer2_outputs[7254] = ~(layer1_outputs[1471]);
    assign layer2_outputs[7255] = layer1_outputs[7732];
    assign layer2_outputs[7256] = ~(layer1_outputs[1306]);
    assign layer2_outputs[7257] = ~((layer1_outputs[2759]) ^ (layer1_outputs[1477]));
    assign layer2_outputs[7258] = ~((layer1_outputs[2114]) & (layer1_outputs[9796]));
    assign layer2_outputs[7259] = layer1_outputs[7514];
    assign layer2_outputs[7260] = layer1_outputs[7244];
    assign layer2_outputs[7261] = ~(layer1_outputs[11134]);
    assign layer2_outputs[7262] = layer1_outputs[9468];
    assign layer2_outputs[7263] = layer1_outputs[9184];
    assign layer2_outputs[7264] = layer1_outputs[882];
    assign layer2_outputs[7265] = layer1_outputs[8236];
    assign layer2_outputs[7266] = ~((layer1_outputs[2379]) ^ (layer1_outputs[4683]));
    assign layer2_outputs[7267] = ~(layer1_outputs[4071]);
    assign layer2_outputs[7268] = (layer1_outputs[2398]) ^ (layer1_outputs[505]);
    assign layer2_outputs[7269] = (layer1_outputs[3200]) | (layer1_outputs[12615]);
    assign layer2_outputs[7270] = ~((layer1_outputs[2353]) ^ (layer1_outputs[2000]));
    assign layer2_outputs[7271] = (layer1_outputs[5723]) & (layer1_outputs[2577]);
    assign layer2_outputs[7272] = ~((layer1_outputs[1462]) ^ (layer1_outputs[5034]));
    assign layer2_outputs[7273] = layer1_outputs[245];
    assign layer2_outputs[7274] = layer1_outputs[8097];
    assign layer2_outputs[7275] = (layer1_outputs[832]) ^ (layer1_outputs[609]);
    assign layer2_outputs[7276] = ~(layer1_outputs[8964]) | (layer1_outputs[2708]);
    assign layer2_outputs[7277] = (layer1_outputs[3664]) & ~(layer1_outputs[2433]);
    assign layer2_outputs[7278] = layer1_outputs[7929];
    assign layer2_outputs[7279] = ~(layer1_outputs[3645]);
    assign layer2_outputs[7280] = layer1_outputs[6950];
    assign layer2_outputs[7281] = layer1_outputs[10555];
    assign layer2_outputs[7282] = ~(layer1_outputs[12767]);
    assign layer2_outputs[7283] = ~(layer1_outputs[6249]) | (layer1_outputs[7406]);
    assign layer2_outputs[7284] = (layer1_outputs[6349]) & ~(layer1_outputs[8810]);
    assign layer2_outputs[7285] = ~(layer1_outputs[3393]);
    assign layer2_outputs[7286] = ~(layer1_outputs[4715]);
    assign layer2_outputs[7287] = (layer1_outputs[2348]) ^ (layer1_outputs[12422]);
    assign layer2_outputs[7288] = ~((layer1_outputs[12265]) ^ (layer1_outputs[9387]));
    assign layer2_outputs[7289] = ~((layer1_outputs[11494]) | (layer1_outputs[6407]));
    assign layer2_outputs[7290] = (layer1_outputs[9044]) & ~(layer1_outputs[8773]);
    assign layer2_outputs[7291] = ~(layer1_outputs[7061]);
    assign layer2_outputs[7292] = ~((layer1_outputs[12071]) ^ (layer1_outputs[11231]));
    assign layer2_outputs[7293] = ~(layer1_outputs[1792]);
    assign layer2_outputs[7294] = ~(layer1_outputs[6791]);
    assign layer2_outputs[7295] = (layer1_outputs[3040]) & ~(layer1_outputs[8527]);
    assign layer2_outputs[7296] = layer1_outputs[861];
    assign layer2_outputs[7297] = ~(layer1_outputs[9988]);
    assign layer2_outputs[7298] = (layer1_outputs[11707]) & (layer1_outputs[11688]);
    assign layer2_outputs[7299] = (layer1_outputs[10396]) & ~(layer1_outputs[6579]);
    assign layer2_outputs[7300] = ~(layer1_outputs[3307]);
    assign layer2_outputs[7301] = ~(layer1_outputs[9459]);
    assign layer2_outputs[7302] = layer1_outputs[4100];
    assign layer2_outputs[7303] = (layer1_outputs[10685]) & ~(layer1_outputs[2006]);
    assign layer2_outputs[7304] = (layer1_outputs[7491]) | (layer1_outputs[4476]);
    assign layer2_outputs[7305] = layer1_outputs[4691];
    assign layer2_outputs[7306] = (layer1_outputs[6522]) ^ (layer1_outputs[11783]);
    assign layer2_outputs[7307] = layer1_outputs[6717];
    assign layer2_outputs[7308] = ~(layer1_outputs[3812]);
    assign layer2_outputs[7309] = ~(layer1_outputs[8615]);
    assign layer2_outputs[7310] = (layer1_outputs[4395]) | (layer1_outputs[11848]);
    assign layer2_outputs[7311] = 1'b0;
    assign layer2_outputs[7312] = 1'b0;
    assign layer2_outputs[7313] = ~(layer1_outputs[12759]);
    assign layer2_outputs[7314] = layer1_outputs[4999];
    assign layer2_outputs[7315] = (layer1_outputs[3871]) | (layer1_outputs[10191]);
    assign layer2_outputs[7316] = ~(layer1_outputs[9207]);
    assign layer2_outputs[7317] = layer1_outputs[4517];
    assign layer2_outputs[7318] = ~(layer1_outputs[11133]) | (layer1_outputs[9814]);
    assign layer2_outputs[7319] = layer1_outputs[12575];
    assign layer2_outputs[7320] = (layer1_outputs[2445]) & (layer1_outputs[11756]);
    assign layer2_outputs[7321] = (layer1_outputs[12638]) | (layer1_outputs[466]);
    assign layer2_outputs[7322] = 1'b0;
    assign layer2_outputs[7323] = ~(layer1_outputs[1976]);
    assign layer2_outputs[7324] = (layer1_outputs[12684]) ^ (layer1_outputs[11235]);
    assign layer2_outputs[7325] = ~(layer1_outputs[4291]);
    assign layer2_outputs[7326] = ~((layer1_outputs[5504]) | (layer1_outputs[10344]));
    assign layer2_outputs[7327] = (layer1_outputs[11802]) & ~(layer1_outputs[7649]);
    assign layer2_outputs[7328] = ~(layer1_outputs[2285]);
    assign layer2_outputs[7329] = ~(layer1_outputs[2741]);
    assign layer2_outputs[7330] = layer1_outputs[8972];
    assign layer2_outputs[7331] = ~(layer1_outputs[797]);
    assign layer2_outputs[7332] = 1'b0;
    assign layer2_outputs[7333] = ~(layer1_outputs[10725]);
    assign layer2_outputs[7334] = ~(layer1_outputs[9172]);
    assign layer2_outputs[7335] = ~(layer1_outputs[10719]);
    assign layer2_outputs[7336] = (layer1_outputs[5593]) & ~(layer1_outputs[11221]);
    assign layer2_outputs[7337] = ~((layer1_outputs[4042]) ^ (layer1_outputs[10282]));
    assign layer2_outputs[7338] = ~(layer1_outputs[11441]);
    assign layer2_outputs[7339] = ~(layer1_outputs[11473]);
    assign layer2_outputs[7340] = (layer1_outputs[7956]) ^ (layer1_outputs[7195]);
    assign layer2_outputs[7341] = ~(layer1_outputs[1329]);
    assign layer2_outputs[7342] = 1'b1;
    assign layer2_outputs[7343] = ~((layer1_outputs[8059]) ^ (layer1_outputs[12457]));
    assign layer2_outputs[7344] = ~(layer1_outputs[11360]);
    assign layer2_outputs[7345] = ~(layer1_outputs[6877]);
    assign layer2_outputs[7346] = ~(layer1_outputs[11773]);
    assign layer2_outputs[7347] = ~(layer1_outputs[12772]);
    assign layer2_outputs[7348] = (layer1_outputs[1522]) ^ (layer1_outputs[6623]);
    assign layer2_outputs[7349] = layer1_outputs[5220];
    assign layer2_outputs[7350] = ~(layer1_outputs[6044]);
    assign layer2_outputs[7351] = (layer1_outputs[8161]) ^ (layer1_outputs[8660]);
    assign layer2_outputs[7352] = ~((layer1_outputs[976]) & (layer1_outputs[2436]));
    assign layer2_outputs[7353] = ~(layer1_outputs[3492]);
    assign layer2_outputs[7354] = ~(layer1_outputs[760]) | (layer1_outputs[1957]);
    assign layer2_outputs[7355] = (layer1_outputs[10425]) & ~(layer1_outputs[2228]);
    assign layer2_outputs[7356] = ~(layer1_outputs[7534]);
    assign layer2_outputs[7357] = layer1_outputs[954];
    assign layer2_outputs[7358] = layer1_outputs[2771];
    assign layer2_outputs[7359] = ~(layer1_outputs[4649]);
    assign layer2_outputs[7360] = layer1_outputs[9094];
    assign layer2_outputs[7361] = (layer1_outputs[6628]) ^ (layer1_outputs[12089]);
    assign layer2_outputs[7362] = (layer1_outputs[4765]) ^ (layer1_outputs[11904]);
    assign layer2_outputs[7363] = layer1_outputs[9455];
    assign layer2_outputs[7364] = ~(layer1_outputs[1810]) | (layer1_outputs[5080]);
    assign layer2_outputs[7365] = ~(layer1_outputs[1134]);
    assign layer2_outputs[7366] = (layer1_outputs[11697]) | (layer1_outputs[9047]);
    assign layer2_outputs[7367] = ~(layer1_outputs[8888]);
    assign layer2_outputs[7368] = layer1_outputs[7811];
    assign layer2_outputs[7369] = ~(layer1_outputs[8625]);
    assign layer2_outputs[7370] = layer1_outputs[618];
    assign layer2_outputs[7371] = ~(layer1_outputs[8254]) | (layer1_outputs[7263]);
    assign layer2_outputs[7372] = ~(layer1_outputs[2926]);
    assign layer2_outputs[7373] = (layer1_outputs[2075]) ^ (layer1_outputs[5741]);
    assign layer2_outputs[7374] = ~(layer1_outputs[6419]);
    assign layer2_outputs[7375] = ~(layer1_outputs[8821]) | (layer1_outputs[2115]);
    assign layer2_outputs[7376] = layer1_outputs[4908];
    assign layer2_outputs[7377] = layer1_outputs[4553];
    assign layer2_outputs[7378] = (layer1_outputs[1368]) ^ (layer1_outputs[8715]);
    assign layer2_outputs[7379] = ~(layer1_outputs[2920]) | (layer1_outputs[6462]);
    assign layer2_outputs[7380] = layer1_outputs[7941];
    assign layer2_outputs[7381] = layer1_outputs[1888];
    assign layer2_outputs[7382] = layer1_outputs[7961];
    assign layer2_outputs[7383] = ~(layer1_outputs[5559]) | (layer1_outputs[6127]);
    assign layer2_outputs[7384] = (layer1_outputs[2870]) & (layer1_outputs[10784]);
    assign layer2_outputs[7385] = ~((layer1_outputs[9746]) | (layer1_outputs[12550]));
    assign layer2_outputs[7386] = ~((layer1_outputs[4358]) ^ (layer1_outputs[1885]));
    assign layer2_outputs[7387] = (layer1_outputs[1504]) & ~(layer1_outputs[5349]);
    assign layer2_outputs[7388] = ~((layer1_outputs[6694]) ^ (layer1_outputs[7898]));
    assign layer2_outputs[7389] = ~((layer1_outputs[5836]) | (layer1_outputs[1432]));
    assign layer2_outputs[7390] = ~(layer1_outputs[438]);
    assign layer2_outputs[7391] = (layer1_outputs[501]) & ~(layer1_outputs[1458]);
    assign layer2_outputs[7392] = ~((layer1_outputs[5876]) ^ (layer1_outputs[9103]));
    assign layer2_outputs[7393] = ~(layer1_outputs[8458]) | (layer1_outputs[739]);
    assign layer2_outputs[7394] = (layer1_outputs[3407]) | (layer1_outputs[2286]);
    assign layer2_outputs[7395] = (layer1_outputs[3563]) & ~(layer1_outputs[4641]);
    assign layer2_outputs[7396] = layer1_outputs[7860];
    assign layer2_outputs[7397] = ~((layer1_outputs[2807]) | (layer1_outputs[12457]));
    assign layer2_outputs[7398] = ~(layer1_outputs[6703]);
    assign layer2_outputs[7399] = ~((layer1_outputs[12563]) | (layer1_outputs[5945]));
    assign layer2_outputs[7400] = ~(layer1_outputs[12255]);
    assign layer2_outputs[7401] = ~((layer1_outputs[6642]) & (layer1_outputs[3529]));
    assign layer2_outputs[7402] = (layer1_outputs[10061]) ^ (layer1_outputs[2902]);
    assign layer2_outputs[7403] = (layer1_outputs[3081]) & ~(layer1_outputs[11328]);
    assign layer2_outputs[7404] = ~(layer1_outputs[6179]) | (layer1_outputs[10553]);
    assign layer2_outputs[7405] = layer1_outputs[9506];
    assign layer2_outputs[7406] = (layer1_outputs[4268]) ^ (layer1_outputs[150]);
    assign layer2_outputs[7407] = layer1_outputs[11043];
    assign layer2_outputs[7408] = layer1_outputs[12229];
    assign layer2_outputs[7409] = layer1_outputs[3646];
    assign layer2_outputs[7410] = ~(layer1_outputs[8492]);
    assign layer2_outputs[7411] = (layer1_outputs[11536]) ^ (layer1_outputs[7984]);
    assign layer2_outputs[7412] = ~((layer1_outputs[8272]) ^ (layer1_outputs[3301]));
    assign layer2_outputs[7413] = layer1_outputs[1649];
    assign layer2_outputs[7414] = ~(layer1_outputs[9745]);
    assign layer2_outputs[7415] = ~(layer1_outputs[9888]);
    assign layer2_outputs[7416] = ~(layer1_outputs[5528]);
    assign layer2_outputs[7417] = layer1_outputs[6771];
    assign layer2_outputs[7418] = ~((layer1_outputs[1447]) | (layer1_outputs[7424]));
    assign layer2_outputs[7419] = ~(layer1_outputs[5767]);
    assign layer2_outputs[7420] = ~(layer1_outputs[11722]) | (layer1_outputs[12162]);
    assign layer2_outputs[7421] = ~(layer1_outputs[4912]);
    assign layer2_outputs[7422] = layer1_outputs[2810];
    assign layer2_outputs[7423] = (layer1_outputs[2218]) & (layer1_outputs[6950]);
    assign layer2_outputs[7424] = ~((layer1_outputs[12426]) & (layer1_outputs[9617]));
    assign layer2_outputs[7425] = (layer1_outputs[10317]) & ~(layer1_outputs[2535]);
    assign layer2_outputs[7426] = layer1_outputs[11733];
    assign layer2_outputs[7427] = layer1_outputs[79];
    assign layer2_outputs[7428] = 1'b0;
    assign layer2_outputs[7429] = (layer1_outputs[5426]) | (layer1_outputs[10203]);
    assign layer2_outputs[7430] = ~(layer1_outputs[381]) | (layer1_outputs[8781]);
    assign layer2_outputs[7431] = ~(layer1_outputs[7776]);
    assign layer2_outputs[7432] = ~((layer1_outputs[10430]) ^ (layer1_outputs[9518]));
    assign layer2_outputs[7433] = ~((layer1_outputs[5700]) & (layer1_outputs[3559]));
    assign layer2_outputs[7434] = (layer1_outputs[5853]) & ~(layer1_outputs[8746]);
    assign layer2_outputs[7435] = layer1_outputs[421];
    assign layer2_outputs[7436] = ~((layer1_outputs[3768]) ^ (layer1_outputs[7262]));
    assign layer2_outputs[7437] = ~((layer1_outputs[7476]) ^ (layer1_outputs[3467]));
    assign layer2_outputs[7438] = ~(layer1_outputs[10372]);
    assign layer2_outputs[7439] = ~(layer1_outputs[10305]);
    assign layer2_outputs[7440] = layer1_outputs[12170];
    assign layer2_outputs[7441] = ~((layer1_outputs[3396]) ^ (layer1_outputs[2172]));
    assign layer2_outputs[7442] = ~(layer1_outputs[8623]);
    assign layer2_outputs[7443] = ~(layer1_outputs[12193]);
    assign layer2_outputs[7444] = (layer1_outputs[11838]) ^ (layer1_outputs[11039]);
    assign layer2_outputs[7445] = layer1_outputs[240];
    assign layer2_outputs[7446] = (layer1_outputs[7785]) ^ (layer1_outputs[5825]);
    assign layer2_outputs[7447] = (layer1_outputs[10216]) ^ (layer1_outputs[5175]);
    assign layer2_outputs[7448] = ~((layer1_outputs[7692]) ^ (layer1_outputs[7794]));
    assign layer2_outputs[7449] = ~(layer1_outputs[11230]) | (layer1_outputs[4237]);
    assign layer2_outputs[7450] = ~((layer1_outputs[9806]) ^ (layer1_outputs[7068]));
    assign layer2_outputs[7451] = ~(layer1_outputs[3793]);
    assign layer2_outputs[7452] = ~(layer1_outputs[8000]) | (layer1_outputs[1901]);
    assign layer2_outputs[7453] = layer1_outputs[7781];
    assign layer2_outputs[7454] = ~(layer1_outputs[9248]);
    assign layer2_outputs[7455] = ~(layer1_outputs[3429]);
    assign layer2_outputs[7456] = ~((layer1_outputs[8345]) & (layer1_outputs[4574]));
    assign layer2_outputs[7457] = (layer1_outputs[2071]) ^ (layer1_outputs[11727]);
    assign layer2_outputs[7458] = layer1_outputs[9136];
    assign layer2_outputs[7459] = ~(layer1_outputs[4657]);
    assign layer2_outputs[7460] = (layer1_outputs[4679]) | (layer1_outputs[6843]);
    assign layer2_outputs[7461] = ~((layer1_outputs[3618]) & (layer1_outputs[7016]));
    assign layer2_outputs[7462] = ~(layer1_outputs[5937]) | (layer1_outputs[5352]);
    assign layer2_outputs[7463] = ~(layer1_outputs[5362]) | (layer1_outputs[11976]);
    assign layer2_outputs[7464] = layer1_outputs[12164];
    assign layer2_outputs[7465] = (layer1_outputs[2023]) ^ (layer1_outputs[9167]);
    assign layer2_outputs[7466] = ~(layer1_outputs[2521]);
    assign layer2_outputs[7467] = layer1_outputs[572];
    assign layer2_outputs[7468] = (layer1_outputs[1612]) ^ (layer1_outputs[838]);
    assign layer2_outputs[7469] = ~(layer1_outputs[7489]) | (layer1_outputs[8812]);
    assign layer2_outputs[7470] = layer1_outputs[6452];
    assign layer2_outputs[7471] = (layer1_outputs[7719]) ^ (layer1_outputs[8199]);
    assign layer2_outputs[7472] = (layer1_outputs[12483]) ^ (layer1_outputs[8114]);
    assign layer2_outputs[7473] = layer1_outputs[5291];
    assign layer2_outputs[7474] = layer1_outputs[1428];
    assign layer2_outputs[7475] = ~(layer1_outputs[10318]);
    assign layer2_outputs[7476] = ~(layer1_outputs[2617]);
    assign layer2_outputs[7477] = 1'b0;
    assign layer2_outputs[7478] = ~(layer1_outputs[6908]);
    assign layer2_outputs[7479] = ~((layer1_outputs[4738]) ^ (layer1_outputs[8360]));
    assign layer2_outputs[7480] = layer1_outputs[3347];
    assign layer2_outputs[7481] = ~(layer1_outputs[8690]);
    assign layer2_outputs[7482] = (layer1_outputs[7276]) ^ (layer1_outputs[5883]);
    assign layer2_outputs[7483] = layer1_outputs[8393];
    assign layer2_outputs[7484] = (layer1_outputs[7042]) ^ (layer1_outputs[7028]);
    assign layer2_outputs[7485] = (layer1_outputs[7564]) & ~(layer1_outputs[4902]);
    assign layer2_outputs[7486] = ~(layer1_outputs[1124]);
    assign layer2_outputs[7487] = ~(layer1_outputs[2957]) | (layer1_outputs[11897]);
    assign layer2_outputs[7488] = 1'b0;
    assign layer2_outputs[7489] = (layer1_outputs[8633]) & (layer1_outputs[12039]);
    assign layer2_outputs[7490] = ~(layer1_outputs[3786]) | (layer1_outputs[7748]);
    assign layer2_outputs[7491] = ~(layer1_outputs[6643]);
    assign layer2_outputs[7492] = (layer1_outputs[7188]) & ~(layer1_outputs[4436]);
    assign layer2_outputs[7493] = ~((layer1_outputs[5334]) ^ (layer1_outputs[9221]));
    assign layer2_outputs[7494] = ~(layer1_outputs[9194]) | (layer1_outputs[11683]);
    assign layer2_outputs[7495] = (layer1_outputs[11070]) & ~(layer1_outputs[9432]);
    assign layer2_outputs[7496] = layer1_outputs[2732];
    assign layer2_outputs[7497] = ~(layer1_outputs[6025]);
    assign layer2_outputs[7498] = layer1_outputs[5187];
    assign layer2_outputs[7499] = layer1_outputs[4977];
    assign layer2_outputs[7500] = ~(layer1_outputs[160]);
    assign layer2_outputs[7501] = (layer1_outputs[12005]) & ~(layer1_outputs[3759]);
    assign layer2_outputs[7502] = layer1_outputs[434];
    assign layer2_outputs[7503] = ~(layer1_outputs[7254]);
    assign layer2_outputs[7504] = layer1_outputs[624];
    assign layer2_outputs[7505] = layer1_outputs[4341];
    assign layer2_outputs[7506] = ~(layer1_outputs[2263]) | (layer1_outputs[8124]);
    assign layer2_outputs[7507] = layer1_outputs[3240];
    assign layer2_outputs[7508] = ~(layer1_outputs[3426]);
    assign layer2_outputs[7509] = (layer1_outputs[5837]) ^ (layer1_outputs[1925]);
    assign layer2_outputs[7510] = ~((layer1_outputs[4952]) ^ (layer1_outputs[11817]));
    assign layer2_outputs[7511] = ~((layer1_outputs[10390]) ^ (layer1_outputs[6324]));
    assign layer2_outputs[7512] = (layer1_outputs[980]) ^ (layer1_outputs[5746]);
    assign layer2_outputs[7513] = ~(layer1_outputs[8496]) | (layer1_outputs[7954]);
    assign layer2_outputs[7514] = (layer1_outputs[9353]) & (layer1_outputs[10643]);
    assign layer2_outputs[7515] = ~(layer1_outputs[8773]);
    assign layer2_outputs[7516] = ~(layer1_outputs[7731]);
    assign layer2_outputs[7517] = (layer1_outputs[2284]) & (layer1_outputs[10370]);
    assign layer2_outputs[7518] = (layer1_outputs[7593]) & ~(layer1_outputs[2269]);
    assign layer2_outputs[7519] = ~(layer1_outputs[2558]);
    assign layer2_outputs[7520] = layer1_outputs[2301];
    assign layer2_outputs[7521] = (layer1_outputs[6707]) & (layer1_outputs[12671]);
    assign layer2_outputs[7522] = ~(layer1_outputs[868]);
    assign layer2_outputs[7523] = (layer1_outputs[5041]) & ~(layer1_outputs[2834]);
    assign layer2_outputs[7524] = ~(layer1_outputs[843]);
    assign layer2_outputs[7525] = layer1_outputs[6497];
    assign layer2_outputs[7526] = (layer1_outputs[492]) ^ (layer1_outputs[11196]);
    assign layer2_outputs[7527] = ~(layer1_outputs[1227]);
    assign layer2_outputs[7528] = (layer1_outputs[664]) & (layer1_outputs[755]);
    assign layer2_outputs[7529] = ~(layer1_outputs[6644]);
    assign layer2_outputs[7530] = layer1_outputs[12134];
    assign layer2_outputs[7531] = ~(layer1_outputs[9999]) | (layer1_outputs[9639]);
    assign layer2_outputs[7532] = (layer1_outputs[5057]) ^ (layer1_outputs[8362]);
    assign layer2_outputs[7533] = ~(layer1_outputs[12766]);
    assign layer2_outputs[7534] = layer1_outputs[12127];
    assign layer2_outputs[7535] = ~(layer1_outputs[7821]) | (layer1_outputs[11082]);
    assign layer2_outputs[7536] = (layer1_outputs[8200]) | (layer1_outputs[3317]);
    assign layer2_outputs[7537] = ~(layer1_outputs[1218]);
    assign layer2_outputs[7538] = layer1_outputs[1167];
    assign layer2_outputs[7539] = (layer1_outputs[3901]) & ~(layer1_outputs[10182]);
    assign layer2_outputs[7540] = (layer1_outputs[5771]) & (layer1_outputs[6183]);
    assign layer2_outputs[7541] = (layer1_outputs[404]) & ~(layer1_outputs[7520]);
    assign layer2_outputs[7542] = (layer1_outputs[9782]) | (layer1_outputs[10617]);
    assign layer2_outputs[7543] = ~(layer1_outputs[12485]);
    assign layer2_outputs[7544] = ~((layer1_outputs[1086]) ^ (layer1_outputs[8002]));
    assign layer2_outputs[7545] = (layer1_outputs[2751]) ^ (layer1_outputs[12006]);
    assign layer2_outputs[7546] = layer1_outputs[9437];
    assign layer2_outputs[7547] = layer1_outputs[2095];
    assign layer2_outputs[7548] = ~(layer1_outputs[12777]);
    assign layer2_outputs[7549] = layer1_outputs[2656];
    assign layer2_outputs[7550] = (layer1_outputs[3679]) & ~(layer1_outputs[6288]);
    assign layer2_outputs[7551] = ~(layer1_outputs[11630]);
    assign layer2_outputs[7552] = ~(layer1_outputs[1052]);
    assign layer2_outputs[7553] = ~(layer1_outputs[12451]);
    assign layer2_outputs[7554] = ~(layer1_outputs[11945]);
    assign layer2_outputs[7555] = (layer1_outputs[4423]) & ~(layer1_outputs[4907]);
    assign layer2_outputs[7556] = ~(layer1_outputs[7705]) | (layer1_outputs[12196]);
    assign layer2_outputs[7557] = layer1_outputs[7510];
    assign layer2_outputs[7558] = ~((layer1_outputs[6670]) | (layer1_outputs[5325]));
    assign layer2_outputs[7559] = ~((layer1_outputs[11411]) | (layer1_outputs[8403]));
    assign layer2_outputs[7560] = layer1_outputs[11013];
    assign layer2_outputs[7561] = layer1_outputs[10373];
    assign layer2_outputs[7562] = (layer1_outputs[8172]) & (layer1_outputs[5491]);
    assign layer2_outputs[7563] = layer1_outputs[4304];
    assign layer2_outputs[7564] = (layer1_outputs[1895]) & ~(layer1_outputs[8882]);
    assign layer2_outputs[7565] = ~(layer1_outputs[6009]);
    assign layer2_outputs[7566] = ~(layer1_outputs[10611]) | (layer1_outputs[3269]);
    assign layer2_outputs[7567] = (layer1_outputs[2213]) & ~(layer1_outputs[9490]);
    assign layer2_outputs[7568] = layer1_outputs[5745];
    assign layer2_outputs[7569] = ~(layer1_outputs[4522]) | (layer1_outputs[4110]);
    assign layer2_outputs[7570] = ~(layer1_outputs[8079]) | (layer1_outputs[850]);
    assign layer2_outputs[7571] = ~(layer1_outputs[5975]);
    assign layer2_outputs[7572] = ~(layer1_outputs[3749]) | (layer1_outputs[576]);
    assign layer2_outputs[7573] = ~((layer1_outputs[11818]) & (layer1_outputs[2941]));
    assign layer2_outputs[7574] = layer1_outputs[4709];
    assign layer2_outputs[7575] = layer1_outputs[2975];
    assign layer2_outputs[7576] = (layer1_outputs[5675]) | (layer1_outputs[7082]);
    assign layer2_outputs[7577] = (layer1_outputs[999]) & (layer1_outputs[8988]);
    assign layer2_outputs[7578] = (layer1_outputs[4487]) | (layer1_outputs[9865]);
    assign layer2_outputs[7579] = (layer1_outputs[1126]) | (layer1_outputs[2420]);
    assign layer2_outputs[7580] = layer1_outputs[12724];
    assign layer2_outputs[7581] = ~(layer1_outputs[11664]) | (layer1_outputs[4559]);
    assign layer2_outputs[7582] = layer1_outputs[10235];
    assign layer2_outputs[7583] = ~(layer1_outputs[3682]);
    assign layer2_outputs[7584] = ~(layer1_outputs[2777]);
    assign layer2_outputs[7585] = layer1_outputs[3852];
    assign layer2_outputs[7586] = ~((layer1_outputs[2524]) ^ (layer1_outputs[5641]));
    assign layer2_outputs[7587] = (layer1_outputs[7026]) & (layer1_outputs[6996]);
    assign layer2_outputs[7588] = (layer1_outputs[629]) & (layer1_outputs[2890]);
    assign layer2_outputs[7589] = ~(layer1_outputs[12776]) | (layer1_outputs[8633]);
    assign layer2_outputs[7590] = layer1_outputs[2852];
    assign layer2_outputs[7591] = 1'b0;
    assign layer2_outputs[7592] = ~(layer1_outputs[5536]) | (layer1_outputs[10980]);
    assign layer2_outputs[7593] = ~(layer1_outputs[3611]);
    assign layer2_outputs[7594] = ~((layer1_outputs[12050]) ^ (layer1_outputs[11527]));
    assign layer2_outputs[7595] = ~(layer1_outputs[4213]);
    assign layer2_outputs[7596] = ~((layer1_outputs[2019]) ^ (layer1_outputs[3430]));
    assign layer2_outputs[7597] = ~(layer1_outputs[2850]) | (layer1_outputs[4784]);
    assign layer2_outputs[7598] = layer1_outputs[7349];
    assign layer2_outputs[7599] = ~((layer1_outputs[7670]) ^ (layer1_outputs[5053]));
    assign layer2_outputs[7600] = layer1_outputs[6695];
    assign layer2_outputs[7601] = (layer1_outputs[3094]) & (layer1_outputs[4116]);
    assign layer2_outputs[7602] = ~(layer1_outputs[11668]);
    assign layer2_outputs[7603] = ~((layer1_outputs[12236]) | (layer1_outputs[11798]));
    assign layer2_outputs[7604] = layer1_outputs[9165];
    assign layer2_outputs[7605] = ~(layer1_outputs[10180]);
    assign layer2_outputs[7606] = layer1_outputs[698];
    assign layer2_outputs[7607] = ~(layer1_outputs[7730]) | (layer1_outputs[8348]);
    assign layer2_outputs[7608] = (layer1_outputs[8979]) & (layer1_outputs[4790]);
    assign layer2_outputs[7609] = ~((layer1_outputs[2140]) & (layer1_outputs[1371]));
    assign layer2_outputs[7610] = (layer1_outputs[2472]) | (layer1_outputs[99]);
    assign layer2_outputs[7611] = layer1_outputs[7812];
    assign layer2_outputs[7612] = (layer1_outputs[5950]) & ~(layer1_outputs[1620]);
    assign layer2_outputs[7613] = ~(layer1_outputs[5661]);
    assign layer2_outputs[7614] = ~(layer1_outputs[2965]);
    assign layer2_outputs[7615] = ~(layer1_outputs[5921]);
    assign layer2_outputs[7616] = ~((layer1_outputs[7002]) & (layer1_outputs[7613]));
    assign layer2_outputs[7617] = layer1_outputs[2676];
    assign layer2_outputs[7618] = ~((layer1_outputs[1696]) & (layer1_outputs[4309]));
    assign layer2_outputs[7619] = layer1_outputs[257];
    assign layer2_outputs[7620] = ~((layer1_outputs[12676]) ^ (layer1_outputs[491]));
    assign layer2_outputs[7621] = ~((layer1_outputs[11458]) | (layer1_outputs[7094]));
    assign layer2_outputs[7622] = ~((layer1_outputs[9388]) & (layer1_outputs[5956]));
    assign layer2_outputs[7623] = ~(layer1_outputs[3578]);
    assign layer2_outputs[7624] = ~(layer1_outputs[11127]);
    assign layer2_outputs[7625] = ~((layer1_outputs[7898]) | (layer1_outputs[6170]));
    assign layer2_outputs[7626] = ~((layer1_outputs[4617]) ^ (layer1_outputs[2318]));
    assign layer2_outputs[7627] = layer1_outputs[2897];
    assign layer2_outputs[7628] = layer1_outputs[9264];
    assign layer2_outputs[7629] = ~((layer1_outputs[6012]) & (layer1_outputs[7638]));
    assign layer2_outputs[7630] = ~((layer1_outputs[6585]) ^ (layer1_outputs[3587]));
    assign layer2_outputs[7631] = (layer1_outputs[9242]) ^ (layer1_outputs[7924]);
    assign layer2_outputs[7632] = (layer1_outputs[4262]) & ~(layer1_outputs[123]);
    assign layer2_outputs[7633] = ~(layer1_outputs[4283]) | (layer1_outputs[6821]);
    assign layer2_outputs[7634] = ~(layer1_outputs[3866]);
    assign layer2_outputs[7635] = ~(layer1_outputs[9685]);
    assign layer2_outputs[7636] = ~(layer1_outputs[9256]);
    assign layer2_outputs[7637] = ~(layer1_outputs[2690]) | (layer1_outputs[5573]);
    assign layer2_outputs[7638] = (layer1_outputs[3212]) ^ (layer1_outputs[2512]);
    assign layer2_outputs[7639] = ~(layer1_outputs[8723]);
    assign layer2_outputs[7640] = ~((layer1_outputs[2847]) & (layer1_outputs[7478]));
    assign layer2_outputs[7641] = layer1_outputs[5130];
    assign layer2_outputs[7642] = ~(layer1_outputs[922]);
    assign layer2_outputs[7643] = layer1_outputs[12424];
    assign layer2_outputs[7644] = ~((layer1_outputs[11860]) ^ (layer1_outputs[1910]));
    assign layer2_outputs[7645] = (layer1_outputs[10897]) & ~(layer1_outputs[8031]);
    assign layer2_outputs[7646] = ~(layer1_outputs[242]);
    assign layer2_outputs[7647] = (layer1_outputs[9941]) & (layer1_outputs[9518]);
    assign layer2_outputs[7648] = layer1_outputs[4751];
    assign layer2_outputs[7649] = ~((layer1_outputs[1191]) & (layer1_outputs[1704]));
    assign layer2_outputs[7650] = layer1_outputs[6613];
    assign layer2_outputs[7651] = ~((layer1_outputs[5706]) ^ (layer1_outputs[3128]));
    assign layer2_outputs[7652] = layer1_outputs[8422];
    assign layer2_outputs[7653] = (layer1_outputs[2204]) & ~(layer1_outputs[6628]);
    assign layer2_outputs[7654] = ~((layer1_outputs[5271]) ^ (layer1_outputs[2887]));
    assign layer2_outputs[7655] = ~((layer1_outputs[7925]) ^ (layer1_outputs[5628]));
    assign layer2_outputs[7656] = layer1_outputs[6415];
    assign layer2_outputs[7657] = ~((layer1_outputs[6681]) ^ (layer1_outputs[1869]));
    assign layer2_outputs[7658] = ~(layer1_outputs[7527]);
    assign layer2_outputs[7659] = ~(layer1_outputs[8415]);
    assign layer2_outputs[7660] = ~((layer1_outputs[7646]) | (layer1_outputs[6120]));
    assign layer2_outputs[7661] = layer1_outputs[2439];
    assign layer2_outputs[7662] = layer1_outputs[11070];
    assign layer2_outputs[7663] = ~(layer1_outputs[6370]);
    assign layer2_outputs[7664] = ~(layer1_outputs[6673]);
    assign layer2_outputs[7665] = (layer1_outputs[424]) ^ (layer1_outputs[3636]);
    assign layer2_outputs[7666] = (layer1_outputs[10400]) & ~(layer1_outputs[8766]);
    assign layer2_outputs[7667] = layer1_outputs[4909];
    assign layer2_outputs[7668] = ~(layer1_outputs[4168]);
    assign layer2_outputs[7669] = layer1_outputs[787];
    assign layer2_outputs[7670] = ~(layer1_outputs[1077]);
    assign layer2_outputs[7671] = (layer1_outputs[4662]) & ~(layer1_outputs[3948]);
    assign layer2_outputs[7672] = layer1_outputs[6137];
    assign layer2_outputs[7673] = ~((layer1_outputs[2953]) ^ (layer1_outputs[12584]));
    assign layer2_outputs[7674] = layer1_outputs[1700];
    assign layer2_outputs[7675] = ~(layer1_outputs[4641]);
    assign layer2_outputs[7676] = (layer1_outputs[3538]) & (layer1_outputs[6886]);
    assign layer2_outputs[7677] = layer1_outputs[2108];
    assign layer2_outputs[7678] = ~(layer1_outputs[3835]);
    assign layer2_outputs[7679] = 1'b1;
    assign layer2_outputs[7680] = ~((layer1_outputs[12175]) & (layer1_outputs[180]));
    assign layer2_outputs[7681] = layer1_outputs[9545];
    assign layer2_outputs[7682] = ~(layer1_outputs[11479]) | (layer1_outputs[8846]);
    assign layer2_outputs[7683] = ~(layer1_outputs[9805]);
    assign layer2_outputs[7684] = layer1_outputs[10717];
    assign layer2_outputs[7685] = (layer1_outputs[11622]) & (layer1_outputs[7797]);
    assign layer2_outputs[7686] = layer1_outputs[137];
    assign layer2_outputs[7687] = ~((layer1_outputs[6726]) ^ (layer1_outputs[2934]));
    assign layer2_outputs[7688] = (layer1_outputs[455]) & ~(layer1_outputs[7868]);
    assign layer2_outputs[7689] = ~((layer1_outputs[6053]) ^ (layer1_outputs[4869]));
    assign layer2_outputs[7690] = (layer1_outputs[7113]) | (layer1_outputs[5693]);
    assign layer2_outputs[7691] = ~((layer1_outputs[12552]) ^ (layer1_outputs[5118]));
    assign layer2_outputs[7692] = (layer1_outputs[2698]) ^ (layer1_outputs[11823]);
    assign layer2_outputs[7693] = ~(layer1_outputs[2384]);
    assign layer2_outputs[7694] = ~(layer1_outputs[4504]);
    assign layer2_outputs[7695] = layer1_outputs[9034];
    assign layer2_outputs[7696] = ~(layer1_outputs[3087]) | (layer1_outputs[4067]);
    assign layer2_outputs[7697] = (layer1_outputs[32]) | (layer1_outputs[196]);
    assign layer2_outputs[7698] = layer1_outputs[5897];
    assign layer2_outputs[7699] = (layer1_outputs[6738]) ^ (layer1_outputs[11103]);
    assign layer2_outputs[7700] = (layer1_outputs[4336]) & (layer1_outputs[10422]);
    assign layer2_outputs[7701] = ~(layer1_outputs[7975]) | (layer1_outputs[7441]);
    assign layer2_outputs[7702] = ~(layer1_outputs[5410]) | (layer1_outputs[10701]);
    assign layer2_outputs[7703] = (layer1_outputs[7496]) & ~(layer1_outputs[10451]);
    assign layer2_outputs[7704] = layer1_outputs[12798];
    assign layer2_outputs[7705] = ~((layer1_outputs[9636]) & (layer1_outputs[3234]));
    assign layer2_outputs[7706] = ~(layer1_outputs[787]);
    assign layer2_outputs[7707] = ~(layer1_outputs[7609]) | (layer1_outputs[2905]);
    assign layer2_outputs[7708] = (layer1_outputs[8775]) | (layer1_outputs[12348]);
    assign layer2_outputs[7709] = (layer1_outputs[8141]) & ~(layer1_outputs[5735]);
    assign layer2_outputs[7710] = (layer1_outputs[9890]) & ~(layer1_outputs[7584]);
    assign layer2_outputs[7711] = ~(layer1_outputs[10296]) | (layer1_outputs[1854]);
    assign layer2_outputs[7712] = (layer1_outputs[7869]) ^ (layer1_outputs[1133]);
    assign layer2_outputs[7713] = ~((layer1_outputs[3724]) ^ (layer1_outputs[4924]));
    assign layer2_outputs[7714] = ~(layer1_outputs[5506]) | (layer1_outputs[7495]);
    assign layer2_outputs[7715] = layer1_outputs[413];
    assign layer2_outputs[7716] = layer1_outputs[9279];
    assign layer2_outputs[7717] = ~(layer1_outputs[11767]);
    assign layer2_outputs[7718] = (layer1_outputs[6600]) & (layer1_outputs[1658]);
    assign layer2_outputs[7719] = layer1_outputs[2129];
    assign layer2_outputs[7720] = ~((layer1_outputs[10965]) | (layer1_outputs[5597]));
    assign layer2_outputs[7721] = ~((layer1_outputs[1476]) & (layer1_outputs[11470]));
    assign layer2_outputs[7722] = (layer1_outputs[256]) | (layer1_outputs[8368]);
    assign layer2_outputs[7723] = layer1_outputs[10391];
    assign layer2_outputs[7724] = layer1_outputs[6814];
    assign layer2_outputs[7725] = ~((layer1_outputs[10065]) | (layer1_outputs[829]));
    assign layer2_outputs[7726] = ~(layer1_outputs[4917]);
    assign layer2_outputs[7727] = layer1_outputs[12605];
    assign layer2_outputs[7728] = ~(layer1_outputs[5980]);
    assign layer2_outputs[7729] = ~(layer1_outputs[9243]) | (layer1_outputs[5855]);
    assign layer2_outputs[7730] = ~((layer1_outputs[10318]) & (layer1_outputs[12654]));
    assign layer2_outputs[7731] = ~((layer1_outputs[5067]) | (layer1_outputs[8815]));
    assign layer2_outputs[7732] = layer1_outputs[4903];
    assign layer2_outputs[7733] = ~(layer1_outputs[12609]);
    assign layer2_outputs[7734] = ~((layer1_outputs[7038]) ^ (layer1_outputs[4371]));
    assign layer2_outputs[7735] = (layer1_outputs[4996]) | (layer1_outputs[7810]);
    assign layer2_outputs[7736] = ~(layer1_outputs[11004]);
    assign layer2_outputs[7737] = (layer1_outputs[11724]) & ~(layer1_outputs[3696]);
    assign layer2_outputs[7738] = ~(layer1_outputs[2685]) | (layer1_outputs[1002]);
    assign layer2_outputs[7739] = layer1_outputs[5853];
    assign layer2_outputs[7740] = ~(layer1_outputs[801]);
    assign layer2_outputs[7741] = ~(layer1_outputs[1365]);
    assign layer2_outputs[7742] = ~(layer1_outputs[856]);
    assign layer2_outputs[7743] = ~(layer1_outputs[855]);
    assign layer2_outputs[7744] = ~(layer1_outputs[4877]);
    assign layer2_outputs[7745] = layer1_outputs[3062];
    assign layer2_outputs[7746] = (layer1_outputs[2054]) & (layer1_outputs[7129]);
    assign layer2_outputs[7747] = ~(layer1_outputs[9329]);
    assign layer2_outputs[7748] = (layer1_outputs[11443]) & ~(layer1_outputs[10825]);
    assign layer2_outputs[7749] = ~(layer1_outputs[6046]);
    assign layer2_outputs[7750] = ~(layer1_outputs[10720]) | (layer1_outputs[11564]);
    assign layer2_outputs[7751] = ~(layer1_outputs[7092]);
    assign layer2_outputs[7752] = (layer1_outputs[1336]) & ~(layer1_outputs[6916]);
    assign layer2_outputs[7753] = layer1_outputs[1773];
    assign layer2_outputs[7754] = layer1_outputs[1309];
    assign layer2_outputs[7755] = (layer1_outputs[6842]) & (layer1_outputs[9892]);
    assign layer2_outputs[7756] = layer1_outputs[5307];
    assign layer2_outputs[7757] = ~(layer1_outputs[9355]);
    assign layer2_outputs[7758] = ~((layer1_outputs[9592]) ^ (layer1_outputs[7062]));
    assign layer2_outputs[7759] = layer1_outputs[9930];
    assign layer2_outputs[7760] = ~(layer1_outputs[5150]);
    assign layer2_outputs[7761] = (layer1_outputs[6778]) & ~(layer1_outputs[807]);
    assign layer2_outputs[7762] = ~((layer1_outputs[4491]) | (layer1_outputs[12522]));
    assign layer2_outputs[7763] = ~((layer1_outputs[3236]) & (layer1_outputs[7191]));
    assign layer2_outputs[7764] = layer1_outputs[7444];
    assign layer2_outputs[7765] = (layer1_outputs[1021]) & ~(layer1_outputs[4677]);
    assign layer2_outputs[7766] = layer1_outputs[9009];
    assign layer2_outputs[7767] = ~((layer1_outputs[5116]) | (layer1_outputs[4661]));
    assign layer2_outputs[7768] = layer1_outputs[8357];
    assign layer2_outputs[7769] = layer1_outputs[4610];
    assign layer2_outputs[7770] = (layer1_outputs[7405]) & ~(layer1_outputs[5069]);
    assign layer2_outputs[7771] = ~(layer1_outputs[9077]);
    assign layer2_outputs[7772] = (layer1_outputs[3475]) & ~(layer1_outputs[10867]);
    assign layer2_outputs[7773] = (layer1_outputs[10206]) & (layer1_outputs[9601]);
    assign layer2_outputs[7774] = ~(layer1_outputs[6966]);
    assign layer2_outputs[7775] = (layer1_outputs[4774]) & (layer1_outputs[7396]);
    assign layer2_outputs[7776] = ~((layer1_outputs[8155]) ^ (layer1_outputs[8503]));
    assign layer2_outputs[7777] = (layer1_outputs[7836]) & ~(layer1_outputs[2015]);
    assign layer2_outputs[7778] = ~(layer1_outputs[7586]) | (layer1_outputs[6986]);
    assign layer2_outputs[7779] = (layer1_outputs[295]) | (layer1_outputs[9350]);
    assign layer2_outputs[7780] = ~(layer1_outputs[7799]) | (layer1_outputs[2633]);
    assign layer2_outputs[7781] = ~(layer1_outputs[4384]) | (layer1_outputs[894]);
    assign layer2_outputs[7782] = (layer1_outputs[8422]) & (layer1_outputs[346]);
    assign layer2_outputs[7783] = layer1_outputs[12370];
    assign layer2_outputs[7784] = ~((layer1_outputs[1558]) | (layer1_outputs[9236]));
    assign layer2_outputs[7785] = layer1_outputs[3693];
    assign layer2_outputs[7786] = (layer1_outputs[3086]) & ~(layer1_outputs[5887]);
    assign layer2_outputs[7787] = (layer1_outputs[3744]) | (layer1_outputs[10002]);
    assign layer2_outputs[7788] = ~(layer1_outputs[7554]) | (layer1_outputs[7432]);
    assign layer2_outputs[7789] = layer1_outputs[8037];
    assign layer2_outputs[7790] = ~(layer1_outputs[6915]);
    assign layer2_outputs[7791] = ~((layer1_outputs[4426]) | (layer1_outputs[3188]));
    assign layer2_outputs[7792] = ~(layer1_outputs[8167]);
    assign layer2_outputs[7793] = ~(layer1_outputs[10432]);
    assign layer2_outputs[7794] = ~((layer1_outputs[11566]) | (layer1_outputs[1176]));
    assign layer2_outputs[7795] = layer1_outputs[3440];
    assign layer2_outputs[7796] = ~((layer1_outputs[10263]) | (layer1_outputs[8609]));
    assign layer2_outputs[7797] = (layer1_outputs[8253]) & ~(layer1_outputs[1087]);
    assign layer2_outputs[7798] = (layer1_outputs[486]) & ~(layer1_outputs[2617]);
    assign layer2_outputs[7799] = ~((layer1_outputs[2053]) | (layer1_outputs[12169]));
    assign layer2_outputs[7800] = layer1_outputs[3635];
    assign layer2_outputs[7801] = ~(layer1_outputs[5568]) | (layer1_outputs[1178]);
    assign layer2_outputs[7802] = ~(layer1_outputs[10592]);
    assign layer2_outputs[7803] = layer1_outputs[7049];
    assign layer2_outputs[7804] = ~(layer1_outputs[626]);
    assign layer2_outputs[7805] = ~(layer1_outputs[4263]);
    assign layer2_outputs[7806] = ~(layer1_outputs[10020]);
    assign layer2_outputs[7807] = ~(layer1_outputs[7710]) | (layer1_outputs[8365]);
    assign layer2_outputs[7808] = ~((layer1_outputs[5508]) ^ (layer1_outputs[4235]));
    assign layer2_outputs[7809] = layer1_outputs[277];
    assign layer2_outputs[7810] = ~(layer1_outputs[1876]);
    assign layer2_outputs[7811] = (layer1_outputs[10731]) ^ (layer1_outputs[6373]);
    assign layer2_outputs[7812] = layer1_outputs[11390];
    assign layer2_outputs[7813] = ~(layer1_outputs[1205]);
    assign layer2_outputs[7814] = ~((layer1_outputs[5098]) ^ (layer1_outputs[841]));
    assign layer2_outputs[7815] = ~((layer1_outputs[1362]) | (layer1_outputs[8905]));
    assign layer2_outputs[7816] = (layer1_outputs[5760]) ^ (layer1_outputs[7625]);
    assign layer2_outputs[7817] = layer1_outputs[519];
    assign layer2_outputs[7818] = ~(layer1_outputs[1285]) | (layer1_outputs[7890]);
    assign layer2_outputs[7819] = ~((layer1_outputs[1447]) ^ (layer1_outputs[3976]));
    assign layer2_outputs[7820] = layer1_outputs[6809];
    assign layer2_outputs[7821] = (layer1_outputs[4534]) | (layer1_outputs[4934]);
    assign layer2_outputs[7822] = (layer1_outputs[3435]) | (layer1_outputs[8809]);
    assign layer2_outputs[7823] = layer1_outputs[3340];
    assign layer2_outputs[7824] = layer1_outputs[7803];
    assign layer2_outputs[7825] = ~(layer1_outputs[6267]);
    assign layer2_outputs[7826] = layer1_outputs[2306];
    assign layer2_outputs[7827] = layer1_outputs[8455];
    assign layer2_outputs[7828] = ~(layer1_outputs[7764]);
    assign layer2_outputs[7829] = (layer1_outputs[11391]) ^ (layer1_outputs[7020]);
    assign layer2_outputs[7830] = ~(layer1_outputs[1006]);
    assign layer2_outputs[7831] = (layer1_outputs[934]) & ~(layer1_outputs[3419]);
    assign layer2_outputs[7832] = (layer1_outputs[1708]) & ~(layer1_outputs[9014]);
    assign layer2_outputs[7833] = ~(layer1_outputs[874]);
    assign layer2_outputs[7834] = ~(layer1_outputs[4201]);
    assign layer2_outputs[7835] = ~((layer1_outputs[2339]) & (layer1_outputs[3719]));
    assign layer2_outputs[7836] = (layer1_outputs[12497]) | (layer1_outputs[5497]);
    assign layer2_outputs[7837] = (layer1_outputs[12512]) ^ (layer1_outputs[672]);
    assign layer2_outputs[7838] = ~(layer1_outputs[8708]);
    assign layer2_outputs[7839] = layer1_outputs[6358];
    assign layer2_outputs[7840] = ~((layer1_outputs[9792]) ^ (layer1_outputs[6578]));
    assign layer2_outputs[7841] = ~((layer1_outputs[8402]) & (layer1_outputs[5215]));
    assign layer2_outputs[7842] = (layer1_outputs[10122]) & ~(layer1_outputs[12385]);
    assign layer2_outputs[7843] = (layer1_outputs[10574]) ^ (layer1_outputs[8771]);
    assign layer2_outputs[7844] = ~((layer1_outputs[5591]) | (layer1_outputs[7689]));
    assign layer2_outputs[7845] = ~((layer1_outputs[1660]) & (layer1_outputs[8357]));
    assign layer2_outputs[7846] = (layer1_outputs[1370]) & ~(layer1_outputs[10936]);
    assign layer2_outputs[7847] = ~((layer1_outputs[7133]) ^ (layer1_outputs[411]));
    assign layer2_outputs[7848] = (layer1_outputs[37]) ^ (layer1_outputs[8653]);
    assign layer2_outputs[7849] = (layer1_outputs[4381]) & ~(layer1_outputs[12448]);
    assign layer2_outputs[7850] = ~(layer1_outputs[2373]);
    assign layer2_outputs[7851] = ~(layer1_outputs[11343]);
    assign layer2_outputs[7852] = layer1_outputs[3048];
    assign layer2_outputs[7853] = (layer1_outputs[2989]) & ~(layer1_outputs[10966]);
    assign layer2_outputs[7854] = layer1_outputs[7660];
    assign layer2_outputs[7855] = ~(layer1_outputs[6383]);
    assign layer2_outputs[7856] = layer1_outputs[4788];
    assign layer2_outputs[7857] = (layer1_outputs[7981]) | (layer1_outputs[9861]);
    assign layer2_outputs[7858] = ~((layer1_outputs[12244]) & (layer1_outputs[2508]));
    assign layer2_outputs[7859] = layer1_outputs[5080];
    assign layer2_outputs[7860] = ~(layer1_outputs[3612]);
    assign layer2_outputs[7861] = layer1_outputs[6384];
    assign layer2_outputs[7862] = ~(layer1_outputs[11944]);
    assign layer2_outputs[7863] = (layer1_outputs[7851]) & ~(layer1_outputs[1952]);
    assign layer2_outputs[7864] = ~((layer1_outputs[2377]) & (layer1_outputs[9111]));
    assign layer2_outputs[7865] = ~((layer1_outputs[5934]) | (layer1_outputs[10820]));
    assign layer2_outputs[7866] = layer1_outputs[533];
    assign layer2_outputs[7867] = (layer1_outputs[5461]) ^ (layer1_outputs[110]);
    assign layer2_outputs[7868] = ~(layer1_outputs[8619]);
    assign layer2_outputs[7869] = ~((layer1_outputs[8282]) & (layer1_outputs[8578]));
    assign layer2_outputs[7870] = (layer1_outputs[11544]) ^ (layer1_outputs[5961]);
    assign layer2_outputs[7871] = ~(layer1_outputs[12258]);
    assign layer2_outputs[7872] = ~(layer1_outputs[1059]);
    assign layer2_outputs[7873] = layer1_outputs[9409];
    assign layer2_outputs[7874] = layer1_outputs[11362];
    assign layer2_outputs[7875] = ~((layer1_outputs[10792]) | (layer1_outputs[6180]));
    assign layer2_outputs[7876] = ~(layer1_outputs[7021]);
    assign layer2_outputs[7877] = (layer1_outputs[315]) & (layer1_outputs[4343]);
    assign layer2_outputs[7878] = layer1_outputs[9195];
    assign layer2_outputs[7879] = (layer1_outputs[8844]) ^ (layer1_outputs[6789]);
    assign layer2_outputs[7880] = (layer1_outputs[6270]) & (layer1_outputs[12154]);
    assign layer2_outputs[7881] = layer1_outputs[3957];
    assign layer2_outputs[7882] = (layer1_outputs[10925]) & ~(layer1_outputs[11382]);
    assign layer2_outputs[7883] = layer1_outputs[2869];
    assign layer2_outputs[7884] = layer1_outputs[12473];
    assign layer2_outputs[7885] = ~((layer1_outputs[12139]) | (layer1_outputs[8204]));
    assign layer2_outputs[7886] = (layer1_outputs[777]) ^ (layer1_outputs[5775]);
    assign layer2_outputs[7887] = ~(layer1_outputs[1130]);
    assign layer2_outputs[7888] = ~(layer1_outputs[12031]) | (layer1_outputs[3267]);
    assign layer2_outputs[7889] = ~(layer1_outputs[7620]);
    assign layer2_outputs[7890] = ~(layer1_outputs[4925]);
    assign layer2_outputs[7891] = (layer1_outputs[4321]) | (layer1_outputs[3689]);
    assign layer2_outputs[7892] = (layer1_outputs[11154]) & ~(layer1_outputs[1188]);
    assign layer2_outputs[7893] = (layer1_outputs[3078]) & ~(layer1_outputs[10413]);
    assign layer2_outputs[7894] = layer1_outputs[12131];
    assign layer2_outputs[7895] = ~(layer1_outputs[3055]) | (layer1_outputs[5347]);
    assign layer2_outputs[7896] = ~(layer1_outputs[12233]);
    assign layer2_outputs[7897] = ~(layer1_outputs[4470]) | (layer1_outputs[3986]);
    assign layer2_outputs[7898] = (layer1_outputs[3778]) & ~(layer1_outputs[5337]);
    assign layer2_outputs[7899] = ~(layer1_outputs[3944]);
    assign layer2_outputs[7900] = layer1_outputs[3953];
    assign layer2_outputs[7901] = ~((layer1_outputs[8308]) | (layer1_outputs[2898]));
    assign layer2_outputs[7902] = layer1_outputs[7476];
    assign layer2_outputs[7903] = ~(layer1_outputs[1157]) | (layer1_outputs[10628]);
    assign layer2_outputs[7904] = ~(layer1_outputs[3330]);
    assign layer2_outputs[7905] = ~((layer1_outputs[11863]) | (layer1_outputs[5629]));
    assign layer2_outputs[7906] = layer1_outputs[10423];
    assign layer2_outputs[7907] = (layer1_outputs[6972]) ^ (layer1_outputs[3695]);
    assign layer2_outputs[7908] = ~((layer1_outputs[1348]) & (layer1_outputs[10018]));
    assign layer2_outputs[7909] = layer1_outputs[9648];
    assign layer2_outputs[7910] = layer1_outputs[1549];
    assign layer2_outputs[7911] = (layer1_outputs[8158]) | (layer1_outputs[2265]);
    assign layer2_outputs[7912] = ~((layer1_outputs[9837]) ^ (layer1_outputs[463]));
    assign layer2_outputs[7913] = layer1_outputs[10834];
    assign layer2_outputs[7914] = (layer1_outputs[1452]) & (layer1_outputs[9049]);
    assign layer2_outputs[7915] = ~(layer1_outputs[428]);
    assign layer2_outputs[7916] = ~(layer1_outputs[1827]);
    assign layer2_outputs[7917] = ~(layer1_outputs[3934]) | (layer1_outputs[12110]);
    assign layer2_outputs[7918] = ~((layer1_outputs[2103]) ^ (layer1_outputs[5246]));
    assign layer2_outputs[7919] = (layer1_outputs[5985]) & ~(layer1_outputs[10304]);
    assign layer2_outputs[7920] = ~(layer1_outputs[8937]);
    assign layer2_outputs[7921] = ~(layer1_outputs[8057]);
    assign layer2_outputs[7922] = (layer1_outputs[7360]) | (layer1_outputs[10266]);
    assign layer2_outputs[7923] = ~((layer1_outputs[5030]) & (layer1_outputs[8285]));
    assign layer2_outputs[7924] = (layer1_outputs[10298]) & ~(layer1_outputs[12636]);
    assign layer2_outputs[7925] = ~(layer1_outputs[3768]);
    assign layer2_outputs[7926] = (layer1_outputs[284]) | (layer1_outputs[5951]);
    assign layer2_outputs[7927] = ~((layer1_outputs[12394]) & (layer1_outputs[5666]));
    assign layer2_outputs[7928] = layer1_outputs[3906];
    assign layer2_outputs[7929] = layer1_outputs[1508];
    assign layer2_outputs[7930] = ~((layer1_outputs[2132]) ^ (layer1_outputs[2773]));
    assign layer2_outputs[7931] = layer1_outputs[6548];
    assign layer2_outputs[7932] = (layer1_outputs[10362]) & ~(layer1_outputs[1285]);
    assign layer2_outputs[7933] = layer1_outputs[12306];
    assign layer2_outputs[7934] = 1'b1;
    assign layer2_outputs[7935] = (layer1_outputs[5596]) & ~(layer1_outputs[5206]);
    assign layer2_outputs[7936] = (layer1_outputs[2609]) | (layer1_outputs[11922]);
    assign layer2_outputs[7937] = ~(layer1_outputs[2723]);
    assign layer2_outputs[7938] = (layer1_outputs[5121]) ^ (layer1_outputs[11474]);
    assign layer2_outputs[7939] = layer1_outputs[3612];
    assign layer2_outputs[7940] = layer1_outputs[5594];
    assign layer2_outputs[7941] = layer1_outputs[3199];
    assign layer2_outputs[7942] = ~(layer1_outputs[2872]);
    assign layer2_outputs[7943] = ~((layer1_outputs[830]) | (layer1_outputs[1456]));
    assign layer2_outputs[7944] = ~(layer1_outputs[8532]);
    assign layer2_outputs[7945] = layer1_outputs[11557];
    assign layer2_outputs[7946] = ~(layer1_outputs[6699]) | (layer1_outputs[10249]);
    assign layer2_outputs[7947] = layer1_outputs[7951];
    assign layer2_outputs[7948] = layer1_outputs[5002];
    assign layer2_outputs[7949] = ~(layer1_outputs[10729]);
    assign layer2_outputs[7950] = ~(layer1_outputs[815]);
    assign layer2_outputs[7951] = layer1_outputs[208];
    assign layer2_outputs[7952] = layer1_outputs[8457];
    assign layer2_outputs[7953] = ~((layer1_outputs[314]) | (layer1_outputs[689]));
    assign layer2_outputs[7954] = layer1_outputs[1473];
    assign layer2_outputs[7955] = (layer1_outputs[12219]) & (layer1_outputs[5404]);
    assign layer2_outputs[7956] = ~(layer1_outputs[554]);
    assign layer2_outputs[7957] = ~((layer1_outputs[12413]) ^ (layer1_outputs[2290]));
    assign layer2_outputs[7958] = ~((layer1_outputs[65]) ^ (layer1_outputs[11180]));
    assign layer2_outputs[7959] = ~(layer1_outputs[11602]);
    assign layer2_outputs[7960] = ~(layer1_outputs[6297]);
    assign layer2_outputs[7961] = ~(layer1_outputs[8088]) | (layer1_outputs[2915]);
    assign layer2_outputs[7962] = ~(layer1_outputs[11375]);
    assign layer2_outputs[7963] = ~(layer1_outputs[7368]);
    assign layer2_outputs[7964] = ~(layer1_outputs[10647]);
    assign layer2_outputs[7965] = ~(layer1_outputs[11658]);
    assign layer2_outputs[7966] = ~(layer1_outputs[9963]);
    assign layer2_outputs[7967] = ~((layer1_outputs[221]) | (layer1_outputs[1654]));
    assign layer2_outputs[7968] = (layer1_outputs[1480]) ^ (layer1_outputs[209]);
    assign layer2_outputs[7969] = layer1_outputs[8302];
    assign layer2_outputs[7970] = (layer1_outputs[11361]) & ~(layer1_outputs[1032]);
    assign layer2_outputs[7971] = ~(layer1_outputs[1774]);
    assign layer2_outputs[7972] = ~(layer1_outputs[12750]);
    assign layer2_outputs[7973] = 1'b0;
    assign layer2_outputs[7974] = (layer1_outputs[450]) & ~(layer1_outputs[7966]);
    assign layer2_outputs[7975] = ~(layer1_outputs[9758]);
    assign layer2_outputs[7976] = (layer1_outputs[1204]) ^ (layer1_outputs[6677]);
    assign layer2_outputs[7977] = ~((layer1_outputs[3055]) | (layer1_outputs[4545]));
    assign layer2_outputs[7978] = ~(layer1_outputs[9681]);
    assign layer2_outputs[7979] = (layer1_outputs[1500]) & ~(layer1_outputs[2652]);
    assign layer2_outputs[7980] = ~(layer1_outputs[5632]) | (layer1_outputs[6479]);
    assign layer2_outputs[7981] = layer1_outputs[11537];
    assign layer2_outputs[7982] = ~((layer1_outputs[9037]) ^ (layer1_outputs[6808]));
    assign layer2_outputs[7983] = ~(layer1_outputs[10690]) | (layer1_outputs[599]);
    assign layer2_outputs[7984] = ~((layer1_outputs[7263]) & (layer1_outputs[4604]));
    assign layer2_outputs[7985] = (layer1_outputs[12511]) | (layer1_outputs[3371]);
    assign layer2_outputs[7986] = layer1_outputs[3067];
    assign layer2_outputs[7987] = (layer1_outputs[689]) ^ (layer1_outputs[10155]);
    assign layer2_outputs[7988] = ~(layer1_outputs[1682]);
    assign layer2_outputs[7989] = ~((layer1_outputs[2854]) | (layer1_outputs[9933]));
    assign layer2_outputs[7990] = layer1_outputs[12165];
    assign layer2_outputs[7991] = layer1_outputs[750];
    assign layer2_outputs[7992] = ~((layer1_outputs[1580]) ^ (layer1_outputs[5341]));
    assign layer2_outputs[7993] = ~((layer1_outputs[5023]) ^ (layer1_outputs[6841]));
    assign layer2_outputs[7994] = ~(layer1_outputs[6838]);
    assign layer2_outputs[7995] = (layer1_outputs[11873]) & (layer1_outputs[1312]);
    assign layer2_outputs[7996] = layer1_outputs[7093];
    assign layer2_outputs[7997] = ~(layer1_outputs[183]);
    assign layer2_outputs[7998] = ~(layer1_outputs[3386]) | (layer1_outputs[856]);
    assign layer2_outputs[7999] = ~(layer1_outputs[11933]);
    assign layer2_outputs[8000] = layer1_outputs[7259];
    assign layer2_outputs[8001] = (layer1_outputs[1175]) & ~(layer1_outputs[2999]);
    assign layer2_outputs[8002] = ~(layer1_outputs[9204]);
    assign layer2_outputs[8003] = ~(layer1_outputs[10447]);
    assign layer2_outputs[8004] = ~(layer1_outputs[6735]);
    assign layer2_outputs[8005] = ~(layer1_outputs[9169]);
    assign layer2_outputs[8006] = ~(layer1_outputs[8639]) | (layer1_outputs[2761]);
    assign layer2_outputs[8007] = layer1_outputs[881];
    assign layer2_outputs[8008] = (layer1_outputs[11242]) & ~(layer1_outputs[12636]);
    assign layer2_outputs[8009] = ~(layer1_outputs[10258]) | (layer1_outputs[12187]);
    assign layer2_outputs[8010] = ~(layer1_outputs[8041]);
    assign layer2_outputs[8011] = ~(layer1_outputs[10207]);
    assign layer2_outputs[8012] = layer1_outputs[2311];
    assign layer2_outputs[8013] = ~((layer1_outputs[5804]) ^ (layer1_outputs[12787]));
    assign layer2_outputs[8014] = ~(layer1_outputs[10803]);
    assign layer2_outputs[8015] = (layer1_outputs[4697]) ^ (layer1_outputs[3134]);
    assign layer2_outputs[8016] = (layer1_outputs[7388]) & ~(layer1_outputs[4053]);
    assign layer2_outputs[8017] = ~(layer1_outputs[4667]);
    assign layer2_outputs[8018] = (layer1_outputs[1883]) & ~(layer1_outputs[1871]);
    assign layer2_outputs[8019] = 1'b0;
    assign layer2_outputs[8020] = layer1_outputs[9145];
    assign layer2_outputs[8021] = ~(layer1_outputs[11765]);
    assign layer2_outputs[8022] = ~(layer1_outputs[1915]);
    assign layer2_outputs[8023] = ~((layer1_outputs[12481]) ^ (layer1_outputs[5803]));
    assign layer2_outputs[8024] = layer1_outputs[1592];
    assign layer2_outputs[8025] = layer1_outputs[12393];
    assign layer2_outputs[8026] = ~(layer1_outputs[9061]) | (layer1_outputs[4637]);
    assign layer2_outputs[8027] = layer1_outputs[7075];
    assign layer2_outputs[8028] = ~(layer1_outputs[1817]);
    assign layer2_outputs[8029] = (layer1_outputs[6002]) | (layer1_outputs[6513]);
    assign layer2_outputs[8030] = ~(layer1_outputs[6692]);
    assign layer2_outputs[8031] = ~((layer1_outputs[4371]) ^ (layer1_outputs[1079]));
    assign layer2_outputs[8032] = layer1_outputs[8694];
    assign layer2_outputs[8033] = ~(layer1_outputs[7060]);
    assign layer2_outputs[8034] = layer1_outputs[7565];
    assign layer2_outputs[8035] = ~((layer1_outputs[7497]) ^ (layer1_outputs[1830]));
    assign layer2_outputs[8036] = (layer1_outputs[7292]) | (layer1_outputs[11113]);
    assign layer2_outputs[8037] = (layer1_outputs[12369]) ^ (layer1_outputs[11649]);
    assign layer2_outputs[8038] = layer1_outputs[7930];
    assign layer2_outputs[8039] = ~(layer1_outputs[6240]);
    assign layer2_outputs[8040] = (layer1_outputs[6928]) & ~(layer1_outputs[9966]);
    assign layer2_outputs[8041] = layer1_outputs[11462];
    assign layer2_outputs[8042] = ~(layer1_outputs[2359]) | (layer1_outputs[6523]);
    assign layer2_outputs[8043] = ~(layer1_outputs[3790]);
    assign layer2_outputs[8044] = ~((layer1_outputs[3016]) ^ (layer1_outputs[11323]));
    assign layer2_outputs[8045] = layer1_outputs[8064];
    assign layer2_outputs[8046] = (layer1_outputs[2538]) ^ (layer1_outputs[9900]);
    assign layer2_outputs[8047] = layer1_outputs[7633];
    assign layer2_outputs[8048] = ~(layer1_outputs[218]);
    assign layer2_outputs[8049] = (layer1_outputs[4887]) ^ (layer1_outputs[6947]);
    assign layer2_outputs[8050] = ~(layer1_outputs[4185]);
    assign layer2_outputs[8051] = layer1_outputs[2559];
    assign layer2_outputs[8052] = (layer1_outputs[1821]) & (layer1_outputs[11108]);
    assign layer2_outputs[8053] = (layer1_outputs[1278]) ^ (layer1_outputs[549]);
    assign layer2_outputs[8054] = ~(layer1_outputs[3747]);
    assign layer2_outputs[8055] = ~(layer1_outputs[1741]);
    assign layer2_outputs[8056] = ~(layer1_outputs[7150]);
    assign layer2_outputs[8057] = layer1_outputs[9185];
    assign layer2_outputs[8058] = ~(layer1_outputs[2962]) | (layer1_outputs[6535]);
    assign layer2_outputs[8059] = (layer1_outputs[9386]) | (layer1_outputs[11188]);
    assign layer2_outputs[8060] = (layer1_outputs[11063]) & ~(layer1_outputs[4833]);
    assign layer2_outputs[8061] = ~(layer1_outputs[12616]) | (layer1_outputs[5241]);
    assign layer2_outputs[8062] = ~(layer1_outputs[12095]) | (layer1_outputs[803]);
    assign layer2_outputs[8063] = layer1_outputs[9540];
    assign layer2_outputs[8064] = layer1_outputs[6814];
    assign layer2_outputs[8065] = ~(layer1_outputs[5797]) | (layer1_outputs[514]);
    assign layer2_outputs[8066] = (layer1_outputs[11120]) & (layer1_outputs[5733]);
    assign layer2_outputs[8067] = ~(layer1_outputs[6238]) | (layer1_outputs[5658]);
    assign layer2_outputs[8068] = layer1_outputs[6486];
    assign layer2_outputs[8069] = layer1_outputs[4687];
    assign layer2_outputs[8070] = (layer1_outputs[3025]) | (layer1_outputs[12100]);
    assign layer2_outputs[8071] = layer1_outputs[8528];
    assign layer2_outputs[8072] = ~((layer1_outputs[1265]) & (layer1_outputs[9700]));
    assign layer2_outputs[8073] = (layer1_outputs[3515]) | (layer1_outputs[11560]);
    assign layer2_outputs[8074] = ~((layer1_outputs[1301]) | (layer1_outputs[7691]));
    assign layer2_outputs[8075] = (layer1_outputs[10168]) & (layer1_outputs[8965]);
    assign layer2_outputs[8076] = 1'b0;
    assign layer2_outputs[8077] = (layer1_outputs[4333]) | (layer1_outputs[28]);
    assign layer2_outputs[8078] = ~(layer1_outputs[906]) | (layer1_outputs[6100]);
    assign layer2_outputs[8079] = layer1_outputs[6392];
    assign layer2_outputs[8080] = ~(layer1_outputs[5196]) | (layer1_outputs[5972]);
    assign layer2_outputs[8081] = ~((layer1_outputs[12697]) | (layer1_outputs[6519]));
    assign layer2_outputs[8082] = layer1_outputs[4573];
    assign layer2_outputs[8083] = ~(layer1_outputs[4214]);
    assign layer2_outputs[8084] = layer1_outputs[1870];
    assign layer2_outputs[8085] = ~(layer1_outputs[1095]) | (layer1_outputs[6076]);
    assign layer2_outputs[8086] = ~(layer1_outputs[7096]);
    assign layer2_outputs[8087] = layer1_outputs[8696];
    assign layer2_outputs[8088] = (layer1_outputs[7967]) ^ (layer1_outputs[10577]);
    assign layer2_outputs[8089] = ~(layer1_outputs[9385]);
    assign layer2_outputs[8090] = ~(layer1_outputs[10117]) | (layer1_outputs[8381]);
    assign layer2_outputs[8091] = ~(layer1_outputs[2246]);
    assign layer2_outputs[8092] = (layer1_outputs[1978]) & ~(layer1_outputs[5594]);
    assign layer2_outputs[8093] = layer1_outputs[2995];
    assign layer2_outputs[8094] = ~((layer1_outputs[2428]) ^ (layer1_outputs[6967]));
    assign layer2_outputs[8095] = layer1_outputs[1443];
    assign layer2_outputs[8096] = ~((layer1_outputs[11988]) ^ (layer1_outputs[7382]));
    assign layer2_outputs[8097] = ~((layer1_outputs[11431]) ^ (layer1_outputs[2877]));
    assign layer2_outputs[8098] = (layer1_outputs[5200]) & ~(layer1_outputs[7362]);
    assign layer2_outputs[8099] = ~(layer1_outputs[3313]);
    assign layer2_outputs[8100] = ~(layer1_outputs[6092]);
    assign layer2_outputs[8101] = ~((layer1_outputs[11485]) & (layer1_outputs[6793]));
    assign layer2_outputs[8102] = ~(layer1_outputs[4308]) | (layer1_outputs[12439]);
    assign layer2_outputs[8103] = (layer1_outputs[11016]) | (layer1_outputs[245]);
    assign layer2_outputs[8104] = layer1_outputs[8753];
    assign layer2_outputs[8105] = (layer1_outputs[11203]) ^ (layer1_outputs[7559]);
    assign layer2_outputs[8106] = (layer1_outputs[704]) ^ (layer1_outputs[1516]);
    assign layer2_outputs[8107] = (layer1_outputs[3404]) & ~(layer1_outputs[6590]);
    assign layer2_outputs[8108] = (layer1_outputs[260]) | (layer1_outputs[10137]);
    assign layer2_outputs[8109] = ~(layer1_outputs[10015]) | (layer1_outputs[3375]);
    assign layer2_outputs[8110] = ~(layer1_outputs[4087]) | (layer1_outputs[5566]);
    assign layer2_outputs[8111] = layer1_outputs[6278];
    assign layer2_outputs[8112] = ~(layer1_outputs[3279]);
    assign layer2_outputs[8113] = ~(layer1_outputs[1305]) | (layer1_outputs[11526]);
    assign layer2_outputs[8114] = ~(layer1_outputs[12118]);
    assign layer2_outputs[8115] = layer1_outputs[819];
    assign layer2_outputs[8116] = ~(layer1_outputs[673]);
    assign layer2_outputs[8117] = layer1_outputs[5245];
    assign layer2_outputs[8118] = ~(layer1_outputs[6874]);
    assign layer2_outputs[8119] = layer1_outputs[1406];
    assign layer2_outputs[8120] = layer1_outputs[7661];
    assign layer2_outputs[8121] = ~(layer1_outputs[9744]);
    assign layer2_outputs[8122] = ~((layer1_outputs[7158]) | (layer1_outputs[7261]));
    assign layer2_outputs[8123] = ~(layer1_outputs[10111]);
    assign layer2_outputs[8124] = (layer1_outputs[1985]) ^ (layer1_outputs[587]);
    assign layer2_outputs[8125] = layer1_outputs[1131];
    assign layer2_outputs[8126] = ~(layer1_outputs[4286]) | (layer1_outputs[641]);
    assign layer2_outputs[8127] = (layer1_outputs[10964]) & (layer1_outputs[5895]);
    assign layer2_outputs[8128] = layer1_outputs[3653];
    assign layer2_outputs[8129] = (layer1_outputs[10716]) | (layer1_outputs[4022]);
    assign layer2_outputs[8130] = ~(layer1_outputs[6509]);
    assign layer2_outputs[8131] = layer1_outputs[1268];
    assign layer2_outputs[8132] = ~((layer1_outputs[8978]) ^ (layer1_outputs[7147]));
    assign layer2_outputs[8133] = layer1_outputs[5679];
    assign layer2_outputs[8134] = ~((layer1_outputs[1761]) ^ (layer1_outputs[2002]));
    assign layer2_outputs[8135] = (layer1_outputs[9541]) ^ (layer1_outputs[1574]);
    assign layer2_outputs[8136] = layer1_outputs[4200];
    assign layer2_outputs[8137] = layer1_outputs[1579];
    assign layer2_outputs[8138] = ~((layer1_outputs[11291]) | (layer1_outputs[11507]));
    assign layer2_outputs[8139] = ~(layer1_outputs[942]) | (layer1_outputs[12594]);
    assign layer2_outputs[8140] = ~((layer1_outputs[11094]) & (layer1_outputs[366]));
    assign layer2_outputs[8141] = ~(layer1_outputs[634]);
    assign layer2_outputs[8142] = ~((layer1_outputs[3112]) | (layer1_outputs[4376]));
    assign layer2_outputs[8143] = ~((layer1_outputs[7714]) & (layer1_outputs[12230]));
    assign layer2_outputs[8144] = (layer1_outputs[2130]) & ~(layer1_outputs[7865]);
    assign layer2_outputs[8145] = layer1_outputs[9355];
    assign layer2_outputs[8146] = layer1_outputs[12582];
    assign layer2_outputs[8147] = layer1_outputs[3229];
    assign layer2_outputs[8148] = layer1_outputs[11707];
    assign layer2_outputs[8149] = ~(layer1_outputs[1335]);
    assign layer2_outputs[8150] = layer1_outputs[6805];
    assign layer2_outputs[8151] = ~(layer1_outputs[10636]);
    assign layer2_outputs[8152] = ~(layer1_outputs[11001]) | (layer1_outputs[2256]);
    assign layer2_outputs[8153] = layer1_outputs[1370];
    assign layer2_outputs[8154] = ~(layer1_outputs[6093]) | (layer1_outputs[5860]);
    assign layer2_outputs[8155] = (layer1_outputs[9041]) | (layer1_outputs[6945]);
    assign layer2_outputs[8156] = ~(layer1_outputs[12663]) | (layer1_outputs[8168]);
    assign layer2_outputs[8157] = ~(layer1_outputs[199]);
    assign layer2_outputs[8158] = (layer1_outputs[5858]) ^ (layer1_outputs[12425]);
    assign layer2_outputs[8159] = (layer1_outputs[3710]) | (layer1_outputs[8117]);
    assign layer2_outputs[8160] = layer1_outputs[4769];
    assign layer2_outputs[8161] = ~((layer1_outputs[952]) ^ (layer1_outputs[978]));
    assign layer2_outputs[8162] = ~((layer1_outputs[6327]) ^ (layer1_outputs[9940]));
    assign layer2_outputs[8163] = layer1_outputs[4524];
    assign layer2_outputs[8164] = ~((layer1_outputs[7862]) & (layer1_outputs[10379]));
    assign layer2_outputs[8165] = ~((layer1_outputs[2322]) & (layer1_outputs[3091]));
    assign layer2_outputs[8166] = ~(layer1_outputs[2348]) | (layer1_outputs[3755]);
    assign layer2_outputs[8167] = ~(layer1_outputs[1590]);
    assign layer2_outputs[8168] = (layer1_outputs[11912]) | (layer1_outputs[1785]);
    assign layer2_outputs[8169] = ~(layer1_outputs[12633]);
    assign layer2_outputs[8170] = ~(layer1_outputs[2396]);
    assign layer2_outputs[8171] = (layer1_outputs[3202]) | (layer1_outputs[11173]);
    assign layer2_outputs[8172] = ~(layer1_outputs[5927]);
    assign layer2_outputs[8173] = ~(layer1_outputs[9561]) | (layer1_outputs[30]);
    assign layer2_outputs[8174] = ~((layer1_outputs[9657]) & (layer1_outputs[4916]));
    assign layer2_outputs[8175] = layer1_outputs[12108];
    assign layer2_outputs[8176] = ~((layer1_outputs[10132]) & (layer1_outputs[3192]));
    assign layer2_outputs[8177] = layer1_outputs[11631];
    assign layer2_outputs[8178] = ~(layer1_outputs[4408]);
    assign layer2_outputs[8179] = ~(layer1_outputs[12741]) | (layer1_outputs[8050]);
    assign layer2_outputs[8180] = layer1_outputs[895];
    assign layer2_outputs[8181] = layer1_outputs[11953];
    assign layer2_outputs[8182] = ~(layer1_outputs[2528]) | (layer1_outputs[12649]);
    assign layer2_outputs[8183] = (layer1_outputs[7486]) | (layer1_outputs[11815]);
    assign layer2_outputs[8184] = ~(layer1_outputs[7725]);
    assign layer2_outputs[8185] = ~(layer1_outputs[12169]);
    assign layer2_outputs[8186] = (layer1_outputs[11251]) & ~(layer1_outputs[1442]);
    assign layer2_outputs[8187] = ~((layer1_outputs[2430]) | (layer1_outputs[2489]));
    assign layer2_outputs[8188] = ~(layer1_outputs[1196]) | (layer1_outputs[6120]);
    assign layer2_outputs[8189] = layer1_outputs[949];
    assign layer2_outputs[8190] = layer1_outputs[6675];
    assign layer2_outputs[8191] = ~((layer1_outputs[4093]) & (layer1_outputs[975]));
    assign layer2_outputs[8192] = ~(layer1_outputs[2197]);
    assign layer2_outputs[8193] = ~((layer1_outputs[6503]) ^ (layer1_outputs[949]));
    assign layer2_outputs[8194] = ~(layer1_outputs[5725]);
    assign layer2_outputs[8195] = ~((layer1_outputs[11644]) ^ (layer1_outputs[1316]));
    assign layer2_outputs[8196] = layer1_outputs[11539];
    assign layer2_outputs[8197] = ~(layer1_outputs[44]);
    assign layer2_outputs[8198] = layer1_outputs[8631];
    assign layer2_outputs[8199] = layer1_outputs[12069];
    assign layer2_outputs[8200] = ~(layer1_outputs[7239]);
    assign layer2_outputs[8201] = ~((layer1_outputs[10028]) ^ (layer1_outputs[4406]));
    assign layer2_outputs[8202] = (layer1_outputs[6424]) ^ (layer1_outputs[12400]);
    assign layer2_outputs[8203] = (layer1_outputs[12061]) | (layer1_outputs[2066]);
    assign layer2_outputs[8204] = ~(layer1_outputs[2505]) | (layer1_outputs[10340]);
    assign layer2_outputs[8205] = (layer1_outputs[2143]) ^ (layer1_outputs[1989]);
    assign layer2_outputs[8206] = ~((layer1_outputs[11573]) ^ (layer1_outputs[6525]));
    assign layer2_outputs[8207] = ~(layer1_outputs[9254]);
    assign layer2_outputs[8208] = ~(layer1_outputs[8060]) | (layer1_outputs[709]);
    assign layer2_outputs[8209] = (layer1_outputs[7732]) & ~(layer1_outputs[4250]);
    assign layer2_outputs[8210] = layer1_outputs[4205];
    assign layer2_outputs[8211] = ~(layer1_outputs[11606]) | (layer1_outputs[10968]);
    assign layer2_outputs[8212] = (layer1_outputs[10157]) | (layer1_outputs[6573]);
    assign layer2_outputs[8213] = (layer1_outputs[7482]) | (layer1_outputs[8676]);
    assign layer2_outputs[8214] = (layer1_outputs[11445]) & ~(layer1_outputs[4242]);
    assign layer2_outputs[8215] = ~(layer1_outputs[2505]) | (layer1_outputs[2782]);
    assign layer2_outputs[8216] = (layer1_outputs[7908]) ^ (layer1_outputs[9318]);
    assign layer2_outputs[8217] = ~(layer1_outputs[6114]) | (layer1_outputs[8083]);
    assign layer2_outputs[8218] = (layer1_outputs[711]) | (layer1_outputs[10066]);
    assign layer2_outputs[8219] = layer1_outputs[11387];
    assign layer2_outputs[8220] = (layer1_outputs[9292]) | (layer1_outputs[2055]);
    assign layer2_outputs[8221] = ~((layer1_outputs[3722]) ^ (layer1_outputs[6601]));
    assign layer2_outputs[8222] = ~(layer1_outputs[7067]) | (layer1_outputs[11336]);
    assign layer2_outputs[8223] = layer1_outputs[2260];
    assign layer2_outputs[8224] = layer1_outputs[7783];
    assign layer2_outputs[8225] = ~((layer1_outputs[11738]) ^ (layer1_outputs[11750]));
    assign layer2_outputs[8226] = ~(layer1_outputs[12351]);
    assign layer2_outputs[8227] = ~(layer1_outputs[8042]);
    assign layer2_outputs[8228] = ~(layer1_outputs[2423]);
    assign layer2_outputs[8229] = (layer1_outputs[4474]) & ~(layer1_outputs[7587]);
    assign layer2_outputs[8230] = ~((layer1_outputs[10303]) ^ (layer1_outputs[5894]));
    assign layer2_outputs[8231] = layer1_outputs[11367];
    assign layer2_outputs[8232] = layer1_outputs[4290];
    assign layer2_outputs[8233] = layer1_outputs[12451];
    assign layer2_outputs[8234] = ~(layer1_outputs[4845]);
    assign layer2_outputs[8235] = layer1_outputs[474];
    assign layer2_outputs[8236] = ~(layer1_outputs[423]);
    assign layer2_outputs[8237] = layer1_outputs[421];
    assign layer2_outputs[8238] = ~(layer1_outputs[5191]) | (layer1_outputs[3162]);
    assign layer2_outputs[8239] = ~((layer1_outputs[8203]) & (layer1_outputs[5086]));
    assign layer2_outputs[8240] = layer1_outputs[2724];
    assign layer2_outputs[8241] = ~(layer1_outputs[3593]);
    assign layer2_outputs[8242] = (layer1_outputs[3085]) & ~(layer1_outputs[11283]);
    assign layer2_outputs[8243] = ~(layer1_outputs[10683]);
    assign layer2_outputs[8244] = ~((layer1_outputs[4945]) | (layer1_outputs[11151]));
    assign layer2_outputs[8245] = ~((layer1_outputs[12407]) & (layer1_outputs[3971]));
    assign layer2_outputs[8246] = layer1_outputs[8593];
    assign layer2_outputs[8247] = ~((layer1_outputs[507]) & (layer1_outputs[11567]));
    assign layer2_outputs[8248] = layer1_outputs[805];
    assign layer2_outputs[8249] = layer1_outputs[481];
    assign layer2_outputs[8250] = ~(layer1_outputs[9762]);
    assign layer2_outputs[8251] = (layer1_outputs[6033]) & ~(layer1_outputs[6816]);
    assign layer2_outputs[8252] = (layer1_outputs[5567]) ^ (layer1_outputs[3687]);
    assign layer2_outputs[8253] = ~(layer1_outputs[126]);
    assign layer2_outputs[8254] = 1'b1;
    assign layer2_outputs[8255] = layer1_outputs[5882];
    assign layer2_outputs[8256] = ~(layer1_outputs[12373]) | (layer1_outputs[9931]);
    assign layer2_outputs[8257] = (layer1_outputs[334]) & ~(layer1_outputs[12768]);
    assign layer2_outputs[8258] = ~(layer1_outputs[9833]);
    assign layer2_outputs[8259] = ~(layer1_outputs[12580]) | (layer1_outputs[4839]);
    assign layer2_outputs[8260] = ~((layer1_outputs[10752]) | (layer1_outputs[8882]));
    assign layer2_outputs[8261] = ~(layer1_outputs[661]);
    assign layer2_outputs[8262] = ~(layer1_outputs[12138]);
    assign layer2_outputs[8263] = ~((layer1_outputs[8155]) | (layer1_outputs[12670]));
    assign layer2_outputs[8264] = layer1_outputs[1486];
    assign layer2_outputs[8265] = (layer1_outputs[5738]) & (layer1_outputs[8574]);
    assign layer2_outputs[8266] = ~(layer1_outputs[5642]);
    assign layer2_outputs[8267] = ~(layer1_outputs[6458]) | (layer1_outputs[313]);
    assign layer2_outputs[8268] = ~(layer1_outputs[2252]);
    assign layer2_outputs[8269] = (layer1_outputs[3932]) & (layer1_outputs[12201]);
    assign layer2_outputs[8270] = layer1_outputs[5838];
    assign layer2_outputs[8271] = layer1_outputs[5104];
    assign layer2_outputs[8272] = layer1_outputs[7408];
    assign layer2_outputs[8273] = ~((layer1_outputs[135]) & (layer1_outputs[8477]));
    assign layer2_outputs[8274] = ~(layer1_outputs[9778]);
    assign layer2_outputs[8275] = (layer1_outputs[1623]) | (layer1_outputs[4534]);
    assign layer2_outputs[8276] = layer1_outputs[7521];
    assign layer2_outputs[8277] = (layer1_outputs[10578]) | (layer1_outputs[5063]);
    assign layer2_outputs[8278] = layer1_outputs[11593];
    assign layer2_outputs[8279] = ~(layer1_outputs[12667]) | (layer1_outputs[11389]);
    assign layer2_outputs[8280] = ~((layer1_outputs[4991]) ^ (layer1_outputs[10086]));
    assign layer2_outputs[8281] = layer1_outputs[7009];
    assign layer2_outputs[8282] = (layer1_outputs[7024]) & ~(layer1_outputs[8216]);
    assign layer2_outputs[8283] = ~(layer1_outputs[6230]);
    assign layer2_outputs[8284] = (layer1_outputs[12231]) | (layer1_outputs[9231]);
    assign layer2_outputs[8285] = ~(layer1_outputs[8457]);
    assign layer2_outputs[8286] = (layer1_outputs[4670]) ^ (layer1_outputs[6021]);
    assign layer2_outputs[8287] = layer1_outputs[7839];
    assign layer2_outputs[8288] = ~((layer1_outputs[8788]) & (layer1_outputs[4953]));
    assign layer2_outputs[8289] = ~((layer1_outputs[4166]) & (layer1_outputs[770]));
    assign layer2_outputs[8290] = ~(layer1_outputs[7620]);
    assign layer2_outputs[8291] = ~(layer1_outputs[8748]) | (layer1_outputs[9714]);
    assign layer2_outputs[8292] = layer1_outputs[5921];
    assign layer2_outputs[8293] = ~(layer1_outputs[2508]);
    assign layer2_outputs[8294] = layer1_outputs[7977];
    assign layer2_outputs[8295] = (layer1_outputs[12030]) ^ (layer1_outputs[2429]);
    assign layer2_outputs[8296] = ~(layer1_outputs[7127]) | (layer1_outputs[12350]);
    assign layer2_outputs[8297] = ~(layer1_outputs[11639]) | (layer1_outputs[67]);
    assign layer2_outputs[8298] = layer1_outputs[7239];
    assign layer2_outputs[8299] = layer1_outputs[12310];
    assign layer2_outputs[8300] = (layer1_outputs[7298]) & ~(layer1_outputs[1148]);
    assign layer2_outputs[8301] = (layer1_outputs[9458]) & (layer1_outputs[3961]);
    assign layer2_outputs[8302] = layer1_outputs[5640];
    assign layer2_outputs[8303] = ~(layer1_outputs[786]);
    assign layer2_outputs[8304] = layer1_outputs[5348];
    assign layer2_outputs[8305] = layer1_outputs[12052];
    assign layer2_outputs[8306] = layer1_outputs[3452];
    assign layer2_outputs[8307] = ~(layer1_outputs[2646]) | (layer1_outputs[9040]);
    assign layer2_outputs[8308] = ~(layer1_outputs[8525]);
    assign layer2_outputs[8309] = (layer1_outputs[3852]) & (layer1_outputs[10660]);
    assign layer2_outputs[8310] = ~(layer1_outputs[4554]);
    assign layer2_outputs[8311] = layer1_outputs[1902];
    assign layer2_outputs[8312] = (layer1_outputs[11881]) & ~(layer1_outputs[9064]);
    assign layer2_outputs[8313] = ~(layer1_outputs[11026]);
    assign layer2_outputs[8314] = layer1_outputs[471];
    assign layer2_outputs[8315] = layer1_outputs[6047];
    assign layer2_outputs[8316] = ~((layer1_outputs[10922]) | (layer1_outputs[1368]));
    assign layer2_outputs[8317] = (layer1_outputs[9998]) & ~(layer1_outputs[1980]);
    assign layer2_outputs[8318] = (layer1_outputs[9740]) & (layer1_outputs[12394]);
    assign layer2_outputs[8319] = layer1_outputs[11240];
    assign layer2_outputs[8320] = ~((layer1_outputs[4989]) & (layer1_outputs[1288]));
    assign layer2_outputs[8321] = ~(layer1_outputs[7278]);
    assign layer2_outputs[8322] = layer1_outputs[12682];
    assign layer2_outputs[8323] = ~(layer1_outputs[6538]) | (layer1_outputs[5674]);
    assign layer2_outputs[8324] = (layer1_outputs[8742]) & (layer1_outputs[6712]);
    assign layer2_outputs[8325] = ~((layer1_outputs[9179]) ^ (layer1_outputs[8076]));
    assign layer2_outputs[8326] = layer1_outputs[248];
    assign layer2_outputs[8327] = layer1_outputs[11136];
    assign layer2_outputs[8328] = ~(layer1_outputs[10596]);
    assign layer2_outputs[8329] = ~(layer1_outputs[7179]);
    assign layer2_outputs[8330] = (layer1_outputs[10565]) & (layer1_outputs[4785]);
    assign layer2_outputs[8331] = layer1_outputs[462];
    assign layer2_outputs[8332] = ~(layer1_outputs[5015]);
    assign layer2_outputs[8333] = ~(layer1_outputs[12437]) | (layer1_outputs[7383]);
    assign layer2_outputs[8334] = layer1_outputs[11355];
    assign layer2_outputs[8335] = ~(layer1_outputs[3952]);
    assign layer2_outputs[8336] = layer1_outputs[9085];
    assign layer2_outputs[8337] = layer1_outputs[8524];
    assign layer2_outputs[8338] = ~(layer1_outputs[8778]);
    assign layer2_outputs[8339] = (layer1_outputs[1117]) & (layer1_outputs[865]);
    assign layer2_outputs[8340] = (layer1_outputs[8501]) | (layer1_outputs[8665]);
    assign layer2_outputs[8341] = layer1_outputs[418];
    assign layer2_outputs[8342] = layer1_outputs[887];
    assign layer2_outputs[8343] = ~((layer1_outputs[7010]) | (layer1_outputs[9333]));
    assign layer2_outputs[8344] = layer1_outputs[12660];
    assign layer2_outputs[8345] = ~(layer1_outputs[8521]);
    assign layer2_outputs[8346] = ~(layer1_outputs[4502]) | (layer1_outputs[8231]);
    assign layer2_outputs[8347] = layer1_outputs[2672];
    assign layer2_outputs[8348] = ~(layer1_outputs[3214]);
    assign layer2_outputs[8349] = ~((layer1_outputs[1562]) & (layer1_outputs[1605]));
    assign layer2_outputs[8350] = ~(layer1_outputs[1122]);
    assign layer2_outputs[8351] = ~(layer1_outputs[11492]);
    assign layer2_outputs[8352] = (layer1_outputs[4036]) & ~(layer1_outputs[1842]);
    assign layer2_outputs[8353] = ~(layer1_outputs[11281]) | (layer1_outputs[12117]);
    assign layer2_outputs[8354] = ~(layer1_outputs[3862]);
    assign layer2_outputs[8355] = (layer1_outputs[10037]) & (layer1_outputs[3944]);
    assign layer2_outputs[8356] = ~((layer1_outputs[9933]) & (layer1_outputs[5470]));
    assign layer2_outputs[8357] = ~((layer1_outputs[4059]) & (layer1_outputs[10359]));
    assign layer2_outputs[8358] = layer1_outputs[9265];
    assign layer2_outputs[8359] = ~(layer1_outputs[12642]);
    assign layer2_outputs[8360] = ~(layer1_outputs[3096]) | (layer1_outputs[745]);
    assign layer2_outputs[8361] = ~((layer1_outputs[9926]) | (layer1_outputs[3581]));
    assign layer2_outputs[8362] = 1'b0;
    assign layer2_outputs[8363] = (layer1_outputs[12737]) & ~(layer1_outputs[10988]);
    assign layer2_outputs[8364] = layer1_outputs[10045];
    assign layer2_outputs[8365] = layer1_outputs[11410];
    assign layer2_outputs[8366] = ~(layer1_outputs[11404]);
    assign layer2_outputs[8367] = ~(layer1_outputs[4672]);
    assign layer2_outputs[8368] = ~((layer1_outputs[10352]) | (layer1_outputs[10100]));
    assign layer2_outputs[8369] = ~(layer1_outputs[3300]);
    assign layer2_outputs[8370] = ~(layer1_outputs[4598]);
    assign layer2_outputs[8371] = ~((layer1_outputs[4692]) | (layer1_outputs[4980]));
    assign layer2_outputs[8372] = ~((layer1_outputs[4045]) | (layer1_outputs[2153]));
    assign layer2_outputs[8373] = ~((layer1_outputs[9504]) ^ (layer1_outputs[11747]));
    assign layer2_outputs[8374] = layer1_outputs[855];
    assign layer2_outputs[8375] = (layer1_outputs[651]) | (layer1_outputs[9016]);
    assign layer2_outputs[8376] = ~((layer1_outputs[9843]) ^ (layer1_outputs[10208]));
    assign layer2_outputs[8377] = ~((layer1_outputs[652]) ^ (layer1_outputs[5328]));
    assign layer2_outputs[8378] = ~((layer1_outputs[299]) & (layer1_outputs[6936]));
    assign layer2_outputs[8379] = (layer1_outputs[6226]) & ~(layer1_outputs[5805]);
    assign layer2_outputs[8380] = ~(layer1_outputs[3928]);
    assign layer2_outputs[8381] = layer1_outputs[1055];
    assign layer2_outputs[8382] = ~(layer1_outputs[1897]);
    assign layer2_outputs[8383] = layer1_outputs[7715];
    assign layer2_outputs[8384] = layer1_outputs[7267];
    assign layer2_outputs[8385] = layer1_outputs[1955];
    assign layer2_outputs[8386] = (layer1_outputs[11104]) | (layer1_outputs[5500]);
    assign layer2_outputs[8387] = ~(layer1_outputs[10050]) | (layer1_outputs[11077]);
    assign layer2_outputs[8388] = layer1_outputs[12090];
    assign layer2_outputs[8389] = (layer1_outputs[2352]) ^ (layer1_outputs[702]);
    assign layer2_outputs[8390] = ~(layer1_outputs[10953]);
    assign layer2_outputs[8391] = ~(layer1_outputs[10930]) | (layer1_outputs[9741]);
    assign layer2_outputs[8392] = ~(layer1_outputs[996]);
    assign layer2_outputs[8393] = ~((layer1_outputs[3466]) | (layer1_outputs[9765]));
    assign layer2_outputs[8394] = (layer1_outputs[2329]) & ~(layer1_outputs[11447]);
    assign layer2_outputs[8395] = ~(layer1_outputs[6200]);
    assign layer2_outputs[8396] = ~(layer1_outputs[1325]) | (layer1_outputs[6750]);
    assign layer2_outputs[8397] = ~(layer1_outputs[10192]) | (layer1_outputs[4093]);
    assign layer2_outputs[8398] = (layer1_outputs[4467]) ^ (layer1_outputs[5174]);
    assign layer2_outputs[8399] = ~(layer1_outputs[3314]);
    assign layer2_outputs[8400] = (layer1_outputs[4829]) ^ (layer1_outputs[11995]);
    assign layer2_outputs[8401] = ~(layer1_outputs[2562]);
    assign layer2_outputs[8402] = ~(layer1_outputs[7344]);
    assign layer2_outputs[8403] = (layer1_outputs[133]) ^ (layer1_outputs[4249]);
    assign layer2_outputs[8404] = ~(layer1_outputs[8401]);
    assign layer2_outputs[8405] = layer1_outputs[628];
    assign layer2_outputs[8406] = ~(layer1_outputs[2315]) | (layer1_outputs[6224]);
    assign layer2_outputs[8407] = layer1_outputs[2345];
    assign layer2_outputs[8408] = ~((layer1_outputs[2605]) | (layer1_outputs[12166]));
    assign layer2_outputs[8409] = layer1_outputs[11056];
    assign layer2_outputs[8410] = (layer1_outputs[3249]) | (layer1_outputs[5612]);
    assign layer2_outputs[8411] = layer1_outputs[7903];
    assign layer2_outputs[8412] = (layer1_outputs[12290]) ^ (layer1_outputs[11779]);
    assign layer2_outputs[8413] = ~(layer1_outputs[11901]);
    assign layer2_outputs[8414] = layer1_outputs[1555];
    assign layer2_outputs[8415] = (layer1_outputs[4288]) & ~(layer1_outputs[9683]);
    assign layer2_outputs[8416] = layer1_outputs[10346];
    assign layer2_outputs[8417] = ~((layer1_outputs[5138]) | (layer1_outputs[4507]));
    assign layer2_outputs[8418] = ~((layer1_outputs[5566]) | (layer1_outputs[8939]));
    assign layer2_outputs[8419] = ~((layer1_outputs[8363]) & (layer1_outputs[6836]));
    assign layer2_outputs[8420] = (layer1_outputs[11252]) ^ (layer1_outputs[1942]);
    assign layer2_outputs[8421] = layer1_outputs[699];
    assign layer2_outputs[8422] = (layer1_outputs[11010]) ^ (layer1_outputs[11834]);
    assign layer2_outputs[8423] = ~(layer1_outputs[7416]) | (layer1_outputs[9557]);
    assign layer2_outputs[8424] = ~(layer1_outputs[6072]) | (layer1_outputs[130]);
    assign layer2_outputs[8425] = ~(layer1_outputs[3641]);
    assign layer2_outputs[8426] = layer1_outputs[10575];
    assign layer2_outputs[8427] = (layer1_outputs[4265]) & ~(layer1_outputs[5588]);
    assign layer2_outputs[8428] = ~((layer1_outputs[8329]) & (layer1_outputs[6976]));
    assign layer2_outputs[8429] = (layer1_outputs[6994]) & ~(layer1_outputs[7242]);
    assign layer2_outputs[8430] = (layer1_outputs[5673]) & ~(layer1_outputs[1052]);
    assign layer2_outputs[8431] = ~(layer1_outputs[4126]);
    assign layer2_outputs[8432] = ~((layer1_outputs[11491]) | (layer1_outputs[11787]));
    assign layer2_outputs[8433] = ~(layer1_outputs[5551]) | (layer1_outputs[6202]);
    assign layer2_outputs[8434] = layer1_outputs[5101];
    assign layer2_outputs[8435] = layer1_outputs[1009];
    assign layer2_outputs[8436] = 1'b0;
    assign layer2_outputs[8437] = layer1_outputs[4090];
    assign layer2_outputs[8438] = ~(layer1_outputs[1300]);
    assign layer2_outputs[8439] = ~(layer1_outputs[11043]);
    assign layer2_outputs[8440] = ~((layer1_outputs[6801]) | (layer1_outputs[8175]));
    assign layer2_outputs[8441] = layer1_outputs[10215];
    assign layer2_outputs[8442] = layer1_outputs[12057];
    assign layer2_outputs[8443] = ~(layer1_outputs[9131]);
    assign layer2_outputs[8444] = ~(layer1_outputs[1470]) | (layer1_outputs[3246]);
    assign layer2_outputs[8445] = ~(layer1_outputs[10321]);
    assign layer2_outputs[8446] = layer1_outputs[1000];
    assign layer2_outputs[8447] = ~(layer1_outputs[9154]) | (layer1_outputs[5301]);
    assign layer2_outputs[8448] = ~(layer1_outputs[2829]);
    assign layer2_outputs[8449] = layer1_outputs[4326];
    assign layer2_outputs[8450] = ~(layer1_outputs[10938]) | (layer1_outputs[7759]);
    assign layer2_outputs[8451] = layer1_outputs[11316];
    assign layer2_outputs[8452] = (layer1_outputs[12602]) & ~(layer1_outputs[6088]);
    assign layer2_outputs[8453] = ~((layer1_outputs[11195]) | (layer1_outputs[10673]));
    assign layer2_outputs[8454] = (layer1_outputs[2715]) ^ (layer1_outputs[4361]);
    assign layer2_outputs[8455] = 1'b0;
    assign layer2_outputs[8456] = layer1_outputs[2223];
    assign layer2_outputs[8457] = (layer1_outputs[1616]) | (layer1_outputs[9971]);
    assign layer2_outputs[8458] = (layer1_outputs[1937]) & ~(layer1_outputs[4716]);
    assign layer2_outputs[8459] = (layer1_outputs[1610]) ^ (layer1_outputs[12542]);
    assign layer2_outputs[8460] = ~(layer1_outputs[4783]);
    assign layer2_outputs[8461] = ~(layer1_outputs[6075]);
    assign layer2_outputs[8462] = ~(layer1_outputs[2370]);
    assign layer2_outputs[8463] = layer1_outputs[156];
    assign layer2_outputs[8464] = layer1_outputs[2795];
    assign layer2_outputs[8465] = layer1_outputs[523];
    assign layer2_outputs[8466] = layer1_outputs[11321];
    assign layer2_outputs[8467] = ~(layer1_outputs[1560]) | (layer1_outputs[6430]);
    assign layer2_outputs[8468] = (layer1_outputs[7636]) & (layer1_outputs[7933]);
    assign layer2_outputs[8469] = ~(layer1_outputs[12476]);
    assign layer2_outputs[8470] = layer1_outputs[6686];
    assign layer2_outputs[8471] = (layer1_outputs[7041]) & (layer1_outputs[3120]);
    assign layer2_outputs[8472] = ~((layer1_outputs[3497]) ^ (layer1_outputs[8548]));
    assign layer2_outputs[8473] = layer1_outputs[3449];
    assign layer2_outputs[8474] = ~(layer1_outputs[7730]) | (layer1_outputs[2520]);
    assign layer2_outputs[8475] = (layer1_outputs[10392]) | (layer1_outputs[3153]);
    assign layer2_outputs[8476] = layer1_outputs[530];
    assign layer2_outputs[8477] = ~(layer1_outputs[5190]) | (layer1_outputs[12225]);
    assign layer2_outputs[8478] = (layer1_outputs[6937]) & ~(layer1_outputs[11208]);
    assign layer2_outputs[8479] = ~((layer1_outputs[6199]) ^ (layer1_outputs[11709]));
    assign layer2_outputs[8480] = (layer1_outputs[512]) & ~(layer1_outputs[2893]);
    assign layer2_outputs[8481] = ~(layer1_outputs[2070]);
    assign layer2_outputs[8482] = (layer1_outputs[5759]) & (layer1_outputs[3897]);
    assign layer2_outputs[8483] = (layer1_outputs[1732]) & (layer1_outputs[149]);
    assign layer2_outputs[8484] = ~((layer1_outputs[6442]) ^ (layer1_outputs[7823]));
    assign layer2_outputs[8485] = (layer1_outputs[7795]) ^ (layer1_outputs[3995]);
    assign layer2_outputs[8486] = (layer1_outputs[6621]) & ~(layer1_outputs[5269]);
    assign layer2_outputs[8487] = ~((layer1_outputs[9525]) | (layer1_outputs[35]));
    assign layer2_outputs[8488] = layer1_outputs[9295];
    assign layer2_outputs[8489] = ~((layer1_outputs[11413]) | (layer1_outputs[7206]));
    assign layer2_outputs[8490] = (layer1_outputs[3319]) & ~(layer1_outputs[10148]);
    assign layer2_outputs[8491] = ~(layer1_outputs[2042]);
    assign layer2_outputs[8492] = ~(layer1_outputs[4903]);
    assign layer2_outputs[8493] = layer1_outputs[8467];
    assign layer2_outputs[8494] = (layer1_outputs[9096]) & ~(layer1_outputs[9985]);
    assign layer2_outputs[8495] = layer1_outputs[10354];
    assign layer2_outputs[8496] = ~(layer1_outputs[7085]);
    assign layer2_outputs[8497] = ~(layer1_outputs[762]);
    assign layer2_outputs[8498] = ~(layer1_outputs[5740]) | (layer1_outputs[1336]);
    assign layer2_outputs[8499] = (layer1_outputs[7611]) & (layer1_outputs[1158]);
    assign layer2_outputs[8500] = (layer1_outputs[1265]) | (layer1_outputs[5672]);
    assign layer2_outputs[8501] = layer1_outputs[8707];
    assign layer2_outputs[8502] = layer1_outputs[9445];
    assign layer2_outputs[8503] = ~((layer1_outputs[588]) ^ (layer1_outputs[3090]));
    assign layer2_outputs[8504] = (layer1_outputs[12621]) | (layer1_outputs[12396]);
    assign layer2_outputs[8505] = (layer1_outputs[10414]) ^ (layer1_outputs[2817]);
    assign layer2_outputs[8506] = (layer1_outputs[3845]) ^ (layer1_outputs[11111]);
    assign layer2_outputs[8507] = ~(layer1_outputs[9830]) | (layer1_outputs[3158]);
    assign layer2_outputs[8508] = layer1_outputs[11804];
    assign layer2_outputs[8509] = (layer1_outputs[4558]) ^ (layer1_outputs[11920]);
    assign layer2_outputs[8510] = ~(layer1_outputs[4963]);
    assign layer2_outputs[8511] = ~(layer1_outputs[2049]) | (layer1_outputs[9122]);
    assign layer2_outputs[8512] = (layer1_outputs[2790]) & ~(layer1_outputs[4455]);
    assign layer2_outputs[8513] = (layer1_outputs[1185]) & (layer1_outputs[6797]);
    assign layer2_outputs[8514] = (layer1_outputs[863]) ^ (layer1_outputs[7689]);
    assign layer2_outputs[8515] = layer1_outputs[10903];
    assign layer2_outputs[8516] = ~(layer1_outputs[6112]);
    assign layer2_outputs[8517] = ~(layer1_outputs[4927]) | (layer1_outputs[11811]);
    assign layer2_outputs[8518] = ~(layer1_outputs[12618]);
    assign layer2_outputs[8519] = ~(layer1_outputs[9497]);
    assign layer2_outputs[8520] = ~((layer1_outputs[6758]) & (layer1_outputs[6919]));
    assign layer2_outputs[8521] = layer1_outputs[6091];
    assign layer2_outputs[8522] = layer1_outputs[1444];
    assign layer2_outputs[8523] = (layer1_outputs[8203]) & (layer1_outputs[415]);
    assign layer2_outputs[8524] = 1'b0;
    assign layer2_outputs[8525] = ~(layer1_outputs[6587]) | (layer1_outputs[4325]);
    assign layer2_outputs[8526] = (layer1_outputs[389]) | (layer1_outputs[5060]);
    assign layer2_outputs[8527] = (layer1_outputs[4932]) & ~(layer1_outputs[3615]);
    assign layer2_outputs[8528] = layer1_outputs[10526];
    assign layer2_outputs[8529] = (layer1_outputs[1928]) & ~(layer1_outputs[57]);
    assign layer2_outputs[8530] = ~((layer1_outputs[8975]) ^ (layer1_outputs[3966]));
    assign layer2_outputs[8531] = (layer1_outputs[6836]) & ~(layer1_outputs[1822]);
    assign layer2_outputs[8532] = ~(layer1_outputs[10932]);
    assign layer2_outputs[8533] = ~(layer1_outputs[2912]) | (layer1_outputs[2075]);
    assign layer2_outputs[8534] = layer1_outputs[8868];
    assign layer2_outputs[8535] = ~(layer1_outputs[4669]);
    assign layer2_outputs[8536] = ~(layer1_outputs[4424]);
    assign layer2_outputs[8537] = layer1_outputs[5664];
    assign layer2_outputs[8538] = (layer1_outputs[635]) | (layer1_outputs[12440]);
    assign layer2_outputs[8539] = layer1_outputs[12347];
    assign layer2_outputs[8540] = layer1_outputs[7905];
    assign layer2_outputs[8541] = ~(layer1_outputs[1915]);
    assign layer2_outputs[8542] = layer1_outputs[1737];
    assign layer2_outputs[8543] = ~(layer1_outputs[710]);
    assign layer2_outputs[8544] = (layer1_outputs[5580]) | (layer1_outputs[7232]);
    assign layer2_outputs[8545] = ~((layer1_outputs[5686]) | (layer1_outputs[4255]));
    assign layer2_outputs[8546] = layer1_outputs[6335];
    assign layer2_outputs[8547] = (layer1_outputs[7514]) ^ (layer1_outputs[6652]);
    assign layer2_outputs[8548] = ~(layer1_outputs[3278]) | (layer1_outputs[9162]);
    assign layer2_outputs[8549] = ~(layer1_outputs[1635]);
    assign layer2_outputs[8550] = layer1_outputs[663];
    assign layer2_outputs[8551] = (layer1_outputs[12547]) & ~(layer1_outputs[3750]);
    assign layer2_outputs[8552] = ~(layer1_outputs[726]);
    assign layer2_outputs[8553] = (layer1_outputs[782]) ^ (layer1_outputs[5494]);
    assign layer2_outputs[8554] = ~(layer1_outputs[8313]);
    assign layer2_outputs[8555] = (layer1_outputs[9322]) & ~(layer1_outputs[7941]);
    assign layer2_outputs[8556] = ~(layer1_outputs[1496]);
    assign layer2_outputs[8557] = layer1_outputs[4415];
    assign layer2_outputs[8558] = layer1_outputs[8114];
    assign layer2_outputs[8559] = (layer1_outputs[7183]) & ~(layer1_outputs[3568]);
    assign layer2_outputs[8560] = (layer1_outputs[5118]) | (layer1_outputs[9549]);
    assign layer2_outputs[8561] = ~(layer1_outputs[9290]);
    assign layer2_outputs[8562] = ~(layer1_outputs[11437]);
    assign layer2_outputs[8563] = ~(layer1_outputs[5768]);
    assign layer2_outputs[8564] = (layer1_outputs[3573]) & ~(layer1_outputs[7533]);
    assign layer2_outputs[8565] = ~((layer1_outputs[1715]) & (layer1_outputs[6484]));
    assign layer2_outputs[8566] = layer1_outputs[2699];
    assign layer2_outputs[8567] = (layer1_outputs[8712]) ^ (layer1_outputs[621]);
    assign layer2_outputs[8568] = (layer1_outputs[113]) & (layer1_outputs[5763]);
    assign layer2_outputs[8569] = ~(layer1_outputs[4719]) | (layer1_outputs[9783]);
    assign layer2_outputs[8570] = ~((layer1_outputs[8517]) ^ (layer1_outputs[9675]));
    assign layer2_outputs[8571] = (layer1_outputs[654]) ^ (layer1_outputs[5794]);
    assign layer2_outputs[8572] = (layer1_outputs[4510]) ^ (layer1_outputs[4350]);
    assign layer2_outputs[8573] = ~(layer1_outputs[4245]);
    assign layer2_outputs[8574] = ~((layer1_outputs[1399]) ^ (layer1_outputs[9902]));
    assign layer2_outputs[8575] = ~(layer1_outputs[11760]);
    assign layer2_outputs[8576] = (layer1_outputs[7658]) & (layer1_outputs[749]);
    assign layer2_outputs[8577] = ~((layer1_outputs[1141]) & (layer1_outputs[9890]));
    assign layer2_outputs[8578] = layer1_outputs[4043];
    assign layer2_outputs[8579] = (layer1_outputs[5510]) & ~(layer1_outputs[6139]);
    assign layer2_outputs[8580] = layer1_outputs[7734];
    assign layer2_outputs[8581] = ~(layer1_outputs[11219]);
    assign layer2_outputs[8582] = layer1_outputs[10772];
    assign layer2_outputs[8583] = (layer1_outputs[11384]) | (layer1_outputs[8073]);
    assign layer2_outputs[8584] = ~((layer1_outputs[683]) ^ (layer1_outputs[7835]));
    assign layer2_outputs[8585] = ~(layer1_outputs[6303]);
    assign layer2_outputs[8586] = layer1_outputs[756];
    assign layer2_outputs[8587] = (layer1_outputs[10129]) & (layer1_outputs[1748]);
    assign layer2_outputs[8588] = (layer1_outputs[12197]) & ~(layer1_outputs[6843]);
    assign layer2_outputs[8589] = (layer1_outputs[2697]) & ~(layer1_outputs[7244]);
    assign layer2_outputs[8590] = ~(layer1_outputs[2808]);
    assign layer2_outputs[8591] = ~(layer1_outputs[1001]);
    assign layer2_outputs[8592] = (layer1_outputs[1643]) & ~(layer1_outputs[9608]);
    assign layer2_outputs[8593] = (layer1_outputs[6982]) & ~(layer1_outputs[6803]);
    assign layer2_outputs[8594] = layer1_outputs[6069];
    assign layer2_outputs[8595] = layer1_outputs[6017];
    assign layer2_outputs[8596] = ~(layer1_outputs[1921]);
    assign layer2_outputs[8597] = (layer1_outputs[12202]) ^ (layer1_outputs[2342]);
    assign layer2_outputs[8598] = ~((layer1_outputs[11432]) & (layer1_outputs[9584]));
    assign layer2_outputs[8599] = ~(layer1_outputs[11140]) | (layer1_outputs[3674]);
    assign layer2_outputs[8600] = (layer1_outputs[2931]) & (layer1_outputs[7351]);
    assign layer2_outputs[8601] = layer1_outputs[4466];
    assign layer2_outputs[8602] = ~((layer1_outputs[5718]) | (layer1_outputs[5284]));
    assign layer2_outputs[8603] = ~(layer1_outputs[6554]) | (layer1_outputs[212]);
    assign layer2_outputs[8604] = ~(layer1_outputs[4345]);
    assign layer2_outputs[8605] = ~(layer1_outputs[10039]);
    assign layer2_outputs[8606] = ~((layer1_outputs[10844]) | (layer1_outputs[1111]));
    assign layer2_outputs[8607] = ~(layer1_outputs[11680]);
    assign layer2_outputs[8608] = (layer1_outputs[11142]) & ~(layer1_outputs[5460]);
    assign layer2_outputs[8609] = layer1_outputs[373];
    assign layer2_outputs[8610] = ~((layer1_outputs[3976]) | (layer1_outputs[6639]));
    assign layer2_outputs[8611] = ~(layer1_outputs[314]);
    assign layer2_outputs[8612] = ~(layer1_outputs[4000]);
    assign layer2_outputs[8613] = ~(layer1_outputs[1171]);
    assign layer2_outputs[8614] = (layer1_outputs[7614]) | (layer1_outputs[11341]);
    assign layer2_outputs[8615] = layer1_outputs[8082];
    assign layer2_outputs[8616] = layer1_outputs[10822];
    assign layer2_outputs[8617] = (layer1_outputs[11912]) | (layer1_outputs[9763]);
    assign layer2_outputs[8618] = (layer1_outputs[11720]) & (layer1_outputs[3564]);
    assign layer2_outputs[8619] = ~((layer1_outputs[10214]) & (layer1_outputs[4914]));
    assign layer2_outputs[8620] = ~(layer1_outputs[1816]);
    assign layer2_outputs[8621] = (layer1_outputs[4252]) & (layer1_outputs[11894]);
    assign layer2_outputs[8622] = ~(layer1_outputs[4962]);
    assign layer2_outputs[8623] = (layer1_outputs[4865]) & (layer1_outputs[6401]);
    assign layer2_outputs[8624] = ~(layer1_outputs[9138]) | (layer1_outputs[3814]);
    assign layer2_outputs[8625] = ~((layer1_outputs[7366]) ^ (layer1_outputs[4587]));
    assign layer2_outputs[8626] = layer1_outputs[2450];
    assign layer2_outputs[8627] = ~(layer1_outputs[1229]);
    assign layer2_outputs[8628] = (layer1_outputs[4929]) & ~(layer1_outputs[3888]);
    assign layer2_outputs[8629] = 1'b0;
    assign layer2_outputs[8630] = layer1_outputs[3108];
    assign layer2_outputs[8631] = (layer1_outputs[984]) | (layer1_outputs[3547]);
    assign layer2_outputs[8632] = ~(layer1_outputs[591]);
    assign layer2_outputs[8633] = layer1_outputs[8067];
    assign layer2_outputs[8634] = ~(layer1_outputs[9665]);
    assign layer2_outputs[8635] = (layer1_outputs[1851]) & (layer1_outputs[3713]);
    assign layer2_outputs[8636] = layer1_outputs[7501];
    assign layer2_outputs[8637] = layer1_outputs[10931];
    assign layer2_outputs[8638] = (layer1_outputs[4721]) | (layer1_outputs[1983]);
    assign layer2_outputs[8639] = layer1_outputs[7949];
    assign layer2_outputs[8640] = ~(layer1_outputs[913]) | (layer1_outputs[8132]);
    assign layer2_outputs[8641] = (layer1_outputs[1960]) | (layer1_outputs[2667]);
    assign layer2_outputs[8642] = layer1_outputs[6394];
    assign layer2_outputs[8643] = (layer1_outputs[12318]) & ~(layer1_outputs[7459]);
    assign layer2_outputs[8644] = (layer1_outputs[1398]) & ~(layer1_outputs[3894]);
    assign layer2_outputs[8645] = layer1_outputs[5969];
    assign layer2_outputs[8646] = layer1_outputs[2946];
    assign layer2_outputs[8647] = (layer1_outputs[5772]) ^ (layer1_outputs[7014]);
    assign layer2_outputs[8648] = (layer1_outputs[448]) & ~(layer1_outputs[178]);
    assign layer2_outputs[8649] = layer1_outputs[2638];
    assign layer2_outputs[8650] = ~(layer1_outputs[4928]);
    assign layer2_outputs[8651] = ~((layer1_outputs[2210]) & (layer1_outputs[6943]));
    assign layer2_outputs[8652] = ~((layer1_outputs[3636]) & (layer1_outputs[5692]));
    assign layer2_outputs[8653] = (layer1_outputs[3306]) & (layer1_outputs[7250]);
    assign layer2_outputs[8654] = layer1_outputs[6108];
    assign layer2_outputs[8655] = ~((layer1_outputs[5954]) ^ (layer1_outputs[8389]));
    assign layer2_outputs[8656] = (layer1_outputs[12040]) & ~(layer1_outputs[9697]);
    assign layer2_outputs[8657] = ~((layer1_outputs[8835]) ^ (layer1_outputs[3271]));
    assign layer2_outputs[8658] = layer1_outputs[10581];
    assign layer2_outputs[8659] = 1'b1;
    assign layer2_outputs[8660] = ~((layer1_outputs[5335]) & (layer1_outputs[6141]));
    assign layer2_outputs[8661] = ~(layer1_outputs[11662]);
    assign layer2_outputs[8662] = (layer1_outputs[4412]) & ~(layer1_outputs[4771]);
    assign layer2_outputs[8663] = 1'b0;
    assign layer2_outputs[8664] = ~(layer1_outputs[3719]);
    assign layer2_outputs[8665] = layer1_outputs[12619];
    assign layer2_outputs[8666] = ~(layer1_outputs[8381]) | (layer1_outputs[7271]);
    assign layer2_outputs[8667] = layer1_outputs[5237];
    assign layer2_outputs[8668] = ~(layer1_outputs[11372]) | (layer1_outputs[9801]);
    assign layer2_outputs[8669] = ~((layer1_outputs[6443]) ^ (layer1_outputs[10818]));
    assign layer2_outputs[8670] = ~((layer1_outputs[8195]) ^ (layer1_outputs[577]));
    assign layer2_outputs[8671] = ~(layer1_outputs[9108]) | (layer1_outputs[3648]);
    assign layer2_outputs[8672] = layer1_outputs[12370];
    assign layer2_outputs[8673] = (layer1_outputs[12726]) & ~(layer1_outputs[2840]);
    assign layer2_outputs[8674] = ~((layer1_outputs[677]) | (layer1_outputs[6365]));
    assign layer2_outputs[8675] = ~(layer1_outputs[4749]) | (layer1_outputs[2567]);
    assign layer2_outputs[8676] = (layer1_outputs[10264]) ^ (layer1_outputs[8100]);
    assign layer2_outputs[8677] = ~((layer1_outputs[9171]) | (layer1_outputs[3769]));
    assign layer2_outputs[8678] = ~((layer1_outputs[3642]) ^ (layer1_outputs[879]));
    assign layer2_outputs[8679] = ~(layer1_outputs[12386]);
    assign layer2_outputs[8680] = layer1_outputs[7419];
    assign layer2_outputs[8681] = ~(layer1_outputs[11929]);
    assign layer2_outputs[8682] = (layer1_outputs[4261]) & ~(layer1_outputs[2952]);
    assign layer2_outputs[8683] = (layer1_outputs[3802]) ^ (layer1_outputs[1468]);
    assign layer2_outputs[8684] = layer1_outputs[5292];
    assign layer2_outputs[8685] = layer1_outputs[12412];
    assign layer2_outputs[8686] = layer1_outputs[1342];
    assign layer2_outputs[8687] = (layer1_outputs[11986]) | (layer1_outputs[11429]);
    assign layer2_outputs[8688] = ~(layer1_outputs[5189]);
    assign layer2_outputs[8689] = ~((layer1_outputs[10876]) | (layer1_outputs[65]));
    assign layer2_outputs[8690] = ~(layer1_outputs[2099]);
    assign layer2_outputs[8691] = ~(layer1_outputs[8336]) | (layer1_outputs[9470]);
    assign layer2_outputs[8692] = layer1_outputs[7789];
    assign layer2_outputs[8693] = ~(layer1_outputs[6948]);
    assign layer2_outputs[8694] = ~(layer1_outputs[1240]);
    assign layer2_outputs[8695] = (layer1_outputs[1179]) ^ (layer1_outputs[4418]);
    assign layer2_outputs[8696] = (layer1_outputs[2290]) & (layer1_outputs[7152]);
    assign layer2_outputs[8697] = layer1_outputs[6291];
    assign layer2_outputs[8698] = ~((layer1_outputs[9481]) & (layer1_outputs[11375]));
    assign layer2_outputs[8699] = (layer1_outputs[9400]) & ~(layer1_outputs[8990]);
    assign layer2_outputs[8700] = (layer1_outputs[9564]) ^ (layer1_outputs[3072]);
    assign layer2_outputs[8701] = (layer1_outputs[272]) ^ (layer1_outputs[9473]);
    assign layer2_outputs[8702] = 1'b1;
    assign layer2_outputs[8703] = (layer1_outputs[5970]) | (layer1_outputs[10516]);
    assign layer2_outputs[8704] = ~(layer1_outputs[10195]) | (layer1_outputs[8522]);
    assign layer2_outputs[8705] = ~(layer1_outputs[6329]) | (layer1_outputs[9226]);
    assign layer2_outputs[8706] = ~((layer1_outputs[10606]) ^ (layer1_outputs[4605]));
    assign layer2_outputs[8707] = (layer1_outputs[4895]) & (layer1_outputs[9113]);
    assign layer2_outputs[8708] = layer1_outputs[6910];
    assign layer2_outputs[8709] = (layer1_outputs[5161]) | (layer1_outputs[2025]);
    assign layer2_outputs[8710] = ~(layer1_outputs[6788]);
    assign layer2_outputs[8711] = layer1_outputs[864];
    assign layer2_outputs[8712] = (layer1_outputs[3295]) | (layer1_outputs[11068]);
    assign layer2_outputs[8713] = (layer1_outputs[2940]) & ~(layer1_outputs[568]);
    assign layer2_outputs[8714] = layer1_outputs[2781];
    assign layer2_outputs[8715] = 1'b1;
    assign layer2_outputs[8716] = (layer1_outputs[6037]) | (layer1_outputs[4905]);
    assign layer2_outputs[8717] = ~(layer1_outputs[4015]);
    assign layer2_outputs[8718] = ~(layer1_outputs[17]);
    assign layer2_outputs[8719] = (layer1_outputs[9690]) & ~(layer1_outputs[10279]);
    assign layer2_outputs[8720] = layer1_outputs[1685];
    assign layer2_outputs[8721] = ~((layer1_outputs[8421]) & (layer1_outputs[8123]));
    assign layer2_outputs[8722] = ~(layer1_outputs[559]) | (layer1_outputs[10294]);
    assign layer2_outputs[8723] = ~(layer1_outputs[7872]);
    assign layer2_outputs[8724] = layer1_outputs[6128];
    assign layer2_outputs[8725] = ~((layer1_outputs[9561]) | (layer1_outputs[509]));
    assign layer2_outputs[8726] = ~(layer1_outputs[5345]) | (layer1_outputs[9083]);
    assign layer2_outputs[8727] = ~(layer1_outputs[5217]);
    assign layer2_outputs[8728] = ~((layer1_outputs[3614]) | (layer1_outputs[10268]));
    assign layer2_outputs[8729] = (layer1_outputs[1714]) ^ (layer1_outputs[4061]);
    assign layer2_outputs[8730] = ~(layer1_outputs[3859]) | (layer1_outputs[5962]);
    assign layer2_outputs[8731] = layer1_outputs[1255];
    assign layer2_outputs[8732] = ~((layer1_outputs[11445]) ^ (layer1_outputs[12614]));
    assign layer2_outputs[8733] = layer1_outputs[4992];
    assign layer2_outputs[8734] = ~(layer1_outputs[2702]);
    assign layer2_outputs[8735] = (layer1_outputs[4591]) & ~(layer1_outputs[5320]);
    assign layer2_outputs[8736] = ~((layer1_outputs[5571]) | (layer1_outputs[11970]));
    assign layer2_outputs[8737] = (layer1_outputs[5775]) & ~(layer1_outputs[3505]);
    assign layer2_outputs[8738] = (layer1_outputs[436]) ^ (layer1_outputs[10891]);
    assign layer2_outputs[8739] = ~(layer1_outputs[4413]);
    assign layer2_outputs[8740] = (layer1_outputs[3907]) & ~(layer1_outputs[8424]);
    assign layer2_outputs[8741] = ~((layer1_outputs[1840]) ^ (layer1_outputs[10924]));
    assign layer2_outputs[8742] = ~(layer1_outputs[6334]);
    assign layer2_outputs[8743] = (layer1_outputs[8962]) & (layer1_outputs[8845]);
    assign layer2_outputs[8744] = ~((layer1_outputs[6098]) & (layer1_outputs[3481]));
    assign layer2_outputs[8745] = layer1_outputs[4017];
    assign layer2_outputs[8746] = layer1_outputs[3069];
    assign layer2_outputs[8747] = layer1_outputs[3708];
    assign layer2_outputs[8748] = ~(layer1_outputs[7759]);
    assign layer2_outputs[8749] = (layer1_outputs[584]) & ~(layer1_outputs[9924]);
    assign layer2_outputs[8750] = (layer1_outputs[4975]) | (layer1_outputs[5182]);
    assign layer2_outputs[8751] = (layer1_outputs[1744]) & ~(layer1_outputs[1995]);
    assign layer2_outputs[8752] = ~(layer1_outputs[2421]);
    assign layer2_outputs[8753] = ~(layer1_outputs[6360]) | (layer1_outputs[6754]);
    assign layer2_outputs[8754] = (layer1_outputs[4725]) & (layer1_outputs[1987]);
    assign layer2_outputs[8755] = ~(layer1_outputs[7027]) | (layer1_outputs[1244]);
    assign layer2_outputs[8756] = ~(layer1_outputs[781]);
    assign layer2_outputs[8757] = ~((layer1_outputs[5428]) | (layer1_outputs[2806]));
    assign layer2_outputs[8758] = layer1_outputs[936];
    assign layer2_outputs[8759] = ~(layer1_outputs[1637]);
    assign layer2_outputs[8760] = (layer1_outputs[11971]) & ~(layer1_outputs[3448]);
    assign layer2_outputs[8761] = 1'b1;
    assign layer2_outputs[8762] = (layer1_outputs[5681]) ^ (layer1_outputs[1361]);
    assign layer2_outputs[8763] = (layer1_outputs[10016]) & (layer1_outputs[10200]);
    assign layer2_outputs[8764] = layer1_outputs[12107];
    assign layer2_outputs[8765] = (layer1_outputs[7347]) & ~(layer1_outputs[10149]);
    assign layer2_outputs[8766] = layer1_outputs[5336];
    assign layer2_outputs[8767] = layer1_outputs[10833];
    assign layer2_outputs[8768] = ~(layer1_outputs[1269]) | (layer1_outputs[9599]);
    assign layer2_outputs[8769] = ~((layer1_outputs[7243]) & (layer1_outputs[5524]));
    assign layer2_outputs[8770] = layer1_outputs[7582];
    assign layer2_outputs[8771] = (layer1_outputs[2846]) & (layer1_outputs[4867]);
    assign layer2_outputs[8772] = ~((layer1_outputs[6765]) ^ (layer1_outputs[11741]));
    assign layer2_outputs[8773] = layer1_outputs[11077];
    assign layer2_outputs[8774] = ~(layer1_outputs[2296]);
    assign layer2_outputs[8775] = (layer1_outputs[7029]) & ~(layer1_outputs[5931]);
    assign layer2_outputs[8776] = (layer1_outputs[4178]) & (layer1_outputs[735]);
    assign layer2_outputs[8777] = ~(layer1_outputs[12773]) | (layer1_outputs[779]);
    assign layer2_outputs[8778] = (layer1_outputs[6536]) | (layer1_outputs[7237]);
    assign layer2_outputs[8779] = ~(layer1_outputs[12400]) | (layer1_outputs[4147]);
    assign layer2_outputs[8780] = (layer1_outputs[7929]) | (layer1_outputs[4967]);
    assign layer2_outputs[8781] = (layer1_outputs[2496]) & ~(layer1_outputs[6956]);
    assign layer2_outputs[8782] = ~((layer1_outputs[2947]) | (layer1_outputs[10026]));
    assign layer2_outputs[8783] = (layer1_outputs[8287]) & ~(layer1_outputs[6818]);
    assign layer2_outputs[8784] = (layer1_outputs[6526]) & (layer1_outputs[4327]);
    assign layer2_outputs[8785] = layer1_outputs[3652];
    assign layer2_outputs[8786] = layer1_outputs[12099];
    assign layer2_outputs[8787] = ~(layer1_outputs[1202]);
    assign layer2_outputs[8788] = layer1_outputs[9303];
    assign layer2_outputs[8789] = ~(layer1_outputs[5597]);
    assign layer2_outputs[8790] = ~(layer1_outputs[8228]) | (layer1_outputs[9770]);
    assign layer2_outputs[8791] = ~(layer1_outputs[2407]);
    assign layer2_outputs[8792] = ~(layer1_outputs[9]);
    assign layer2_outputs[8793] = ~((layer1_outputs[2503]) & (layer1_outputs[2122]));
    assign layer2_outputs[8794] = layer1_outputs[1779];
    assign layer2_outputs[8795] = (layer1_outputs[1394]) | (layer1_outputs[3675]);
    assign layer2_outputs[8796] = layer1_outputs[1819];
    assign layer2_outputs[8797] = ~(layer1_outputs[5488]);
    assign layer2_outputs[8798] = ~((layer1_outputs[11579]) & (layer1_outputs[3197]));
    assign layer2_outputs[8799] = ~(layer1_outputs[10112]) | (layer1_outputs[4266]);
    assign layer2_outputs[8800] = (layer1_outputs[7160]) ^ (layer1_outputs[4882]);
    assign layer2_outputs[8801] = ~(layer1_outputs[460]);
    assign layer2_outputs[8802] = (layer1_outputs[8870]) ^ (layer1_outputs[6658]);
    assign layer2_outputs[8803] = (layer1_outputs[5421]) & ~(layer1_outputs[2264]);
    assign layer2_outputs[8804] = layer1_outputs[2128];
    assign layer2_outputs[8805] = (layer1_outputs[10960]) ^ (layer1_outputs[11582]);
    assign layer2_outputs[8806] = layer1_outputs[7726];
    assign layer2_outputs[8807] = layer1_outputs[12248];
    assign layer2_outputs[8808] = ~(layer1_outputs[3514]);
    assign layer2_outputs[8809] = (layer1_outputs[11055]) ^ (layer1_outputs[9979]);
    assign layer2_outputs[8810] = (layer1_outputs[7959]) ^ (layer1_outputs[9736]);
    assign layer2_outputs[8811] = (layer1_outputs[5758]) | (layer1_outputs[12116]);
    assign layer2_outputs[8812] = ~((layer1_outputs[10512]) ^ (layer1_outputs[10637]));
    assign layer2_outputs[8813] = ~((layer1_outputs[737]) ^ (layer1_outputs[10662]));
    assign layer2_outputs[8814] = (layer1_outputs[7048]) | (layer1_outputs[1890]);
    assign layer2_outputs[8815] = ~((layer1_outputs[6720]) ^ (layer1_outputs[12271]));
    assign layer2_outputs[8816] = ~(layer1_outputs[10093]) | (layer1_outputs[6472]);
    assign layer2_outputs[8817] = layer1_outputs[5603];
    assign layer2_outputs[8818] = ~((layer1_outputs[10395]) ^ (layer1_outputs[3873]));
    assign layer2_outputs[8819] = ~(layer1_outputs[3241]);
    assign layer2_outputs[8820] = layer1_outputs[11655];
    assign layer2_outputs[8821] = ~(layer1_outputs[739]) | (layer1_outputs[9180]);
    assign layer2_outputs[8822] = layer1_outputs[8504];
    assign layer2_outputs[8823] = ~(layer1_outputs[163]);
    assign layer2_outputs[8824] = ~((layer1_outputs[12353]) | (layer1_outputs[11041]));
    assign layer2_outputs[8825] = (layer1_outputs[4232]) & (layer1_outputs[2940]);
    assign layer2_outputs[8826] = ~((layer1_outputs[6087]) ^ (layer1_outputs[2921]));
    assign layer2_outputs[8827] = ~(layer1_outputs[1144]);
    assign layer2_outputs[8828] = ~((layer1_outputs[8547]) ^ (layer1_outputs[9652]));
    assign layer2_outputs[8829] = (layer1_outputs[11511]) & (layer1_outputs[859]);
    assign layer2_outputs[8830] = ~((layer1_outputs[8230]) & (layer1_outputs[4379]));
    assign layer2_outputs[8831] = ~(layer1_outputs[5333]);
    assign layer2_outputs[8832] = layer1_outputs[11705];
    assign layer2_outputs[8833] = layer1_outputs[3142];
    assign layer2_outputs[8834] = layer1_outputs[9365];
    assign layer2_outputs[8835] = ~(layer1_outputs[6068]);
    assign layer2_outputs[8836] = ~((layer1_outputs[4785]) & (layer1_outputs[9745]));
    assign layer2_outputs[8837] = ~(layer1_outputs[660]);
    assign layer2_outputs[8838] = layer1_outputs[112];
    assign layer2_outputs[8839] = ~(layer1_outputs[11005]);
    assign layer2_outputs[8840] = ~(layer1_outputs[2645]) | (layer1_outputs[3574]);
    assign layer2_outputs[8841] = ~(layer1_outputs[11459]);
    assign layer2_outputs[8842] = (layer1_outputs[2186]) & ~(layer1_outputs[897]);
    assign layer2_outputs[8843] = layer1_outputs[325];
    assign layer2_outputs[8844] = (layer1_outputs[9258]) & (layer1_outputs[7439]);
    assign layer2_outputs[8845] = ~(layer1_outputs[6039]);
    assign layer2_outputs[8846] = (layer1_outputs[9670]) & (layer1_outputs[7409]);
    assign layer2_outputs[8847] = ~(layer1_outputs[6042]) | (layer1_outputs[1321]);
    assign layer2_outputs[8848] = ~(layer1_outputs[7217]);
    assign layer2_outputs[8849] = ~(layer1_outputs[6904]);
    assign layer2_outputs[8850] = ~(layer1_outputs[1546]);
    assign layer2_outputs[8851] = (layer1_outputs[6603]) ^ (layer1_outputs[4973]);
    assign layer2_outputs[8852] = layer1_outputs[3118];
    assign layer2_outputs[8853] = layer1_outputs[2492];
    assign layer2_outputs[8854] = (layer1_outputs[7748]) | (layer1_outputs[562]);
    assign layer2_outputs[8855] = ~((layer1_outputs[12358]) ^ (layer1_outputs[1274]));
    assign layer2_outputs[8856] = ~(layer1_outputs[5193]) | (layer1_outputs[6676]);
    assign layer2_outputs[8857] = layer1_outputs[1847];
    assign layer2_outputs[8858] = ~(layer1_outputs[5370]);
    assign layer2_outputs[8859] = layer1_outputs[6465];
    assign layer2_outputs[8860] = ~((layer1_outputs[3179]) ^ (layer1_outputs[12630]));
    assign layer2_outputs[8861] = 1'b1;
    assign layer2_outputs[8862] = ~((layer1_outputs[11431]) & (layer1_outputs[11201]));
    assign layer2_outputs[8863] = layer1_outputs[8244];
    assign layer2_outputs[8864] = ~(layer1_outputs[3375]);
    assign layer2_outputs[8865] = layer1_outputs[4990];
    assign layer2_outputs[8866] = ~((layer1_outputs[2908]) | (layer1_outputs[10290]));
    assign layer2_outputs[8867] = ~((layer1_outputs[10301]) & (layer1_outputs[4642]));
    assign layer2_outputs[8868] = (layer1_outputs[2747]) ^ (layer1_outputs[11560]);
    assign layer2_outputs[8869] = (layer1_outputs[12415]) ^ (layer1_outputs[8734]);
    assign layer2_outputs[8870] = ~(layer1_outputs[6626]) | (layer1_outputs[1406]);
    assign layer2_outputs[8871] = layer1_outputs[8709];
    assign layer2_outputs[8872] = (layer1_outputs[5499]) & (layer1_outputs[12446]);
    assign layer2_outputs[8873] = ~((layer1_outputs[12392]) ^ (layer1_outputs[1397]));
    assign layer2_outputs[8874] = (layer1_outputs[193]) ^ (layer1_outputs[5208]);
    assign layer2_outputs[8875] = layer1_outputs[503];
    assign layer2_outputs[8876] = (layer1_outputs[2682]) | (layer1_outputs[8382]);
    assign layer2_outputs[8877] = (layer1_outputs[4543]) & ~(layer1_outputs[11435]);
    assign layer2_outputs[8878] = ~(layer1_outputs[7955]);
    assign layer2_outputs[8879] = (layer1_outputs[9389]) & (layer1_outputs[229]);
    assign layer2_outputs[8880] = layer1_outputs[2291];
    assign layer2_outputs[8881] = ~(layer1_outputs[11520]);
    assign layer2_outputs[8882] = layer1_outputs[6208];
    assign layer2_outputs[8883] = ~(layer1_outputs[5561]);
    assign layer2_outputs[8884] = layer1_outputs[9842];
    assign layer2_outputs[8885] = ~(layer1_outputs[11635]);
    assign layer2_outputs[8886] = ~(layer1_outputs[1988]);
    assign layer2_outputs[8887] = (layer1_outputs[1166]) & (layer1_outputs[9393]);
    assign layer2_outputs[8888] = (layer1_outputs[1675]) & ~(layer1_outputs[2767]);
    assign layer2_outputs[8889] = ~(layer1_outputs[246]);
    assign layer2_outputs[8890] = 1'b1;
    assign layer2_outputs[8891] = 1'b1;
    assign layer2_outputs[8892] = ~((layer1_outputs[8031]) & (layer1_outputs[9181]));
    assign layer2_outputs[8893] = ~(layer1_outputs[4259]);
    assign layer2_outputs[8894] = (layer1_outputs[9779]) | (layer1_outputs[7091]);
    assign layer2_outputs[8895] = (layer1_outputs[973]) ^ (layer1_outputs[727]);
    assign layer2_outputs[8896] = (layer1_outputs[688]) | (layer1_outputs[8151]);
    assign layer2_outputs[8897] = ~(layer1_outputs[2751]);
    assign layer2_outputs[8898] = ~(layer1_outputs[648]) | (layer1_outputs[11642]);
    assign layer2_outputs[8899] = (layer1_outputs[9290]) & ~(layer1_outputs[8680]);
    assign layer2_outputs[8900] = ~((layer1_outputs[2826]) ^ (layer1_outputs[9586]));
    assign layer2_outputs[8901] = (layer1_outputs[5858]) ^ (layer1_outputs[3624]);
    assign layer2_outputs[8902] = (layer1_outputs[5235]) ^ (layer1_outputs[6722]);
    assign layer2_outputs[8903] = ~(layer1_outputs[7415]);
    assign layer2_outputs[8904] = ~((layer1_outputs[4939]) ^ (layer1_outputs[12585]));
    assign layer2_outputs[8905] = ~(layer1_outputs[4461]);
    assign layer2_outputs[8906] = (layer1_outputs[4864]) | (layer1_outputs[4194]);
    assign layer2_outputs[8907] = layer1_outputs[9771];
    assign layer2_outputs[8908] = layer1_outputs[3129];
    assign layer2_outputs[8909] = layer1_outputs[4282];
    assign layer2_outputs[8910] = ~(layer1_outputs[3247]) | (layer1_outputs[5360]);
    assign layer2_outputs[8911] = layer1_outputs[1281];
    assign layer2_outputs[8912] = ~((layer1_outputs[12352]) ^ (layer1_outputs[3594]));
    assign layer2_outputs[8913] = layer1_outputs[11370];
    assign layer2_outputs[8914] = (layer1_outputs[73]) & (layer1_outputs[3165]);
    assign layer2_outputs[8915] = layer1_outputs[6034];
    assign layer2_outputs[8916] = (layer1_outputs[3990]) & ~(layer1_outputs[10849]);
    assign layer2_outputs[8917] = ~(layer1_outputs[6835]);
    assign layer2_outputs[8918] = ~((layer1_outputs[11053]) & (layer1_outputs[30]));
    assign layer2_outputs[8919] = ~((layer1_outputs[9440]) & (layer1_outputs[9017]));
    assign layer2_outputs[8920] = (layer1_outputs[8573]) ^ (layer1_outputs[8720]);
    assign layer2_outputs[8921] = (layer1_outputs[5204]) ^ (layer1_outputs[5236]);
    assign layer2_outputs[8922] = ~(layer1_outputs[8244]);
    assign layer2_outputs[8923] = ~((layer1_outputs[5646]) ^ (layer1_outputs[834]));
    assign layer2_outputs[8924] = layer1_outputs[6259];
    assign layer2_outputs[8925] = layer1_outputs[2684];
    assign layer2_outputs[8926] = ~((layer1_outputs[3706]) | (layer1_outputs[10918]));
    assign layer2_outputs[8927] = ~(layer1_outputs[8818]);
    assign layer2_outputs[8928] = (layer1_outputs[7202]) & ~(layer1_outputs[1478]);
    assign layer2_outputs[8929] = ~(layer1_outputs[1668]);
    assign layer2_outputs[8930] = (layer1_outputs[12104]) & (layer1_outputs[7178]);
    assign layer2_outputs[8931] = ~((layer1_outputs[12123]) ^ (layer1_outputs[509]));
    assign layer2_outputs[8932] = (layer1_outputs[3738]) ^ (layer1_outputs[840]);
    assign layer2_outputs[8933] = ~(layer1_outputs[6011]) | (layer1_outputs[2563]);
    assign layer2_outputs[8934] = ~(layer1_outputs[135]) | (layer1_outputs[2653]);
    assign layer2_outputs[8935] = ~(layer1_outputs[1424]);
    assign layer2_outputs[8936] = ~(layer1_outputs[12540]);
    assign layer2_outputs[8937] = layer1_outputs[12528];
    assign layer2_outputs[8938] = layer1_outputs[11872];
    assign layer2_outputs[8939] = ~(layer1_outputs[10617]);
    assign layer2_outputs[8940] = ~(layer1_outputs[10853]);
    assign layer2_outputs[8941] = (layer1_outputs[1374]) ^ (layer1_outputs[6204]);
    assign layer2_outputs[8942] = ~(layer1_outputs[6823]);
    assign layer2_outputs[8943] = layer1_outputs[3074];
    assign layer2_outputs[8944] = ~(layer1_outputs[2816]);
    assign layer2_outputs[8945] = (layer1_outputs[7087]) | (layer1_outputs[10764]);
    assign layer2_outputs[8946] = layer1_outputs[4960];
    assign layer2_outputs[8947] = (layer1_outputs[7870]) | (layer1_outputs[10806]);
    assign layer2_outputs[8948] = ~(layer1_outputs[2545]) | (layer1_outputs[1309]);
    assign layer2_outputs[8949] = ~(layer1_outputs[7942]);
    assign layer2_outputs[8950] = ~(layer1_outputs[9742]);
    assign layer2_outputs[8951] = layer1_outputs[3294];
    assign layer2_outputs[8952] = 1'b1;
    assign layer2_outputs[8953] = ~(layer1_outputs[11548]);
    assign layer2_outputs[8954] = (layer1_outputs[4529]) & ~(layer1_outputs[4525]);
    assign layer2_outputs[8955] = (layer1_outputs[4529]) ^ (layer1_outputs[8554]);
    assign layer2_outputs[8956] = ~(layer1_outputs[6355]);
    assign layer2_outputs[8957] = ~(layer1_outputs[7216]) | (layer1_outputs[6887]);
    assign layer2_outputs[8958] = ~((layer1_outputs[5442]) | (layer1_outputs[5501]));
    assign layer2_outputs[8959] = ~((layer1_outputs[9691]) | (layer1_outputs[6111]));
    assign layer2_outputs[8960] = ~(layer1_outputs[4060]);
    assign layer2_outputs[8961] = ~(layer1_outputs[4624]);
    assign layer2_outputs[8962] = ~((layer1_outputs[1122]) | (layer1_outputs[6117]));
    assign layer2_outputs[8963] = layer1_outputs[1272];
    assign layer2_outputs[8964] = ~(layer1_outputs[2558]);
    assign layer2_outputs[8965] = ~(layer1_outputs[5332]) | (layer1_outputs[12790]);
    assign layer2_outputs[8966] = ~((layer1_outputs[11940]) | (layer1_outputs[8514]));
    assign layer2_outputs[8967] = ~((layer1_outputs[2636]) ^ (layer1_outputs[1179]));
    assign layer2_outputs[8968] = 1'b1;
    assign layer2_outputs[8969] = ~(layer1_outputs[11995]);
    assign layer2_outputs[8970] = (layer1_outputs[12786]) & (layer1_outputs[2709]);
    assign layer2_outputs[8971] = ~(layer1_outputs[9667]);
    assign layer2_outputs[8972] = ~(layer1_outputs[6580]);
    assign layer2_outputs[8973] = layer1_outputs[4088];
    assign layer2_outputs[8974] = (layer1_outputs[7058]) ^ (layer1_outputs[9186]);
    assign layer2_outputs[8975] = layer1_outputs[7924];
    assign layer2_outputs[8976] = layer1_outputs[7323];
    assign layer2_outputs[8977] = ~(layer1_outputs[3779]) | (layer1_outputs[4270]);
    assign layer2_outputs[8978] = (layer1_outputs[11116]) ^ (layer1_outputs[12580]);
    assign layer2_outputs[8979] = (layer1_outputs[8856]) & ~(layer1_outputs[911]);
    assign layer2_outputs[8980] = ~((layer1_outputs[9805]) | (layer1_outputs[2668]));
    assign layer2_outputs[8981] = ~(layer1_outputs[2983]);
    assign layer2_outputs[8982] = (layer1_outputs[3856]) & (layer1_outputs[5997]);
    assign layer2_outputs[8983] = ~((layer1_outputs[10620]) | (layer1_outputs[3454]));
    assign layer2_outputs[8984] = ~(layer1_outputs[3499]);
    assign layer2_outputs[8985] = ~((layer1_outputs[7549]) ^ (layer1_outputs[213]));
    assign layer2_outputs[8986] = (layer1_outputs[10852]) ^ (layer1_outputs[2973]);
    assign layer2_outputs[8987] = ~(layer1_outputs[8192]);
    assign layer2_outputs[8988] = ~(layer1_outputs[3476]);
    assign layer2_outputs[8989] = ~(layer1_outputs[10210]) | (layer1_outputs[4253]);
    assign layer2_outputs[8990] = ~(layer1_outputs[7969]);
    assign layer2_outputs[8991] = layer1_outputs[972];
    assign layer2_outputs[8992] = ~((layer1_outputs[7702]) ^ (layer1_outputs[7640]));
    assign layer2_outputs[8993] = (layer1_outputs[4400]) & (layer1_outputs[4468]);
    assign layer2_outputs[8994] = layer1_outputs[6397];
    assign layer2_outputs[8995] = (layer1_outputs[5670]) ^ (layer1_outputs[9728]);
    assign layer2_outputs[8996] = ~(layer1_outputs[4245]);
    assign layer2_outputs[8997] = (layer1_outputs[9239]) | (layer1_outputs[2459]);
    assign layer2_outputs[8998] = layer1_outputs[6388];
    assign layer2_outputs[8999] = ~(layer1_outputs[2877]);
    assign layer2_outputs[9000] = ~(layer1_outputs[4447]) | (layer1_outputs[2816]);
    assign layer2_outputs[9001] = (layer1_outputs[3982]) & ~(layer1_outputs[8927]);
    assign layer2_outputs[9002] = ~(layer1_outputs[11351]) | (layer1_outputs[6235]);
    assign layer2_outputs[9003] = layer1_outputs[9912];
    assign layer2_outputs[9004] = ~((layer1_outputs[11592]) ^ (layer1_outputs[10909]));
    assign layer2_outputs[9005] = layer1_outputs[10169];
    assign layer2_outputs[9006] = ~(layer1_outputs[6674]) | (layer1_outputs[7003]);
    assign layer2_outputs[9007] = ~((layer1_outputs[4309]) ^ (layer1_outputs[9894]));
    assign layer2_outputs[9008] = layer1_outputs[7148];
    assign layer2_outputs[9009] = (layer1_outputs[10705]) & ~(layer1_outputs[5692]);
    assign layer2_outputs[9010] = ~(layer1_outputs[1626]);
    assign layer2_outputs[9011] = ~(layer1_outputs[2763]);
    assign layer2_outputs[9012] = ~((layer1_outputs[5337]) ^ (layer1_outputs[10552]));
    assign layer2_outputs[9013] = layer1_outputs[10022];
    assign layer2_outputs[9014] = (layer1_outputs[11117]) & (layer1_outputs[859]);
    assign layer2_outputs[9015] = ~((layer1_outputs[12000]) | (layer1_outputs[5934]));
    assign layer2_outputs[9016] = ~(layer1_outputs[5226]);
    assign layer2_outputs[9017] = (layer1_outputs[6017]) & (layer1_outputs[24]);
    assign layer2_outputs[9018] = (layer1_outputs[6796]) | (layer1_outputs[1112]);
    assign layer2_outputs[9019] = (layer1_outputs[5881]) & (layer1_outputs[9174]);
    assign layer2_outputs[9020] = ~((layer1_outputs[9771]) & (layer1_outputs[10816]));
    assign layer2_outputs[9021] = layer1_outputs[10544];
    assign layer2_outputs[9022] = ~(layer1_outputs[1815]) | (layer1_outputs[6336]);
    assign layer2_outputs[9023] = (layer1_outputs[4181]) & ~(layer1_outputs[6711]);
    assign layer2_outputs[9024] = layer1_outputs[4590];
    assign layer2_outputs[9025] = layer1_outputs[11692];
    assign layer2_outputs[9026] = (layer1_outputs[9796]) | (layer1_outputs[4612]);
    assign layer2_outputs[9027] = ~(layer1_outputs[7339]);
    assign layer2_outputs[9028] = ~(layer1_outputs[8991]);
    assign layer2_outputs[9029] = (layer1_outputs[1041]) | (layer1_outputs[8270]);
    assign layer2_outputs[9030] = ~((layer1_outputs[6961]) & (layer1_outputs[12567]));
    assign layer2_outputs[9031] = layer1_outputs[9374];
    assign layer2_outputs[9032] = layer1_outputs[12071];
    assign layer2_outputs[9033] = layer1_outputs[9618];
    assign layer2_outputs[9034] = ~(layer1_outputs[1768]);
    assign layer2_outputs[9035] = ~(layer1_outputs[5274]);
    assign layer2_outputs[9036] = ~((layer1_outputs[4787]) & (layer1_outputs[3267]));
    assign layer2_outputs[9037] = layer1_outputs[2700];
    assign layer2_outputs[9038] = ~((layer1_outputs[1249]) ^ (layer1_outputs[3109]));
    assign layer2_outputs[9039] = ~((layer1_outputs[3565]) ^ (layer1_outputs[10475]));
    assign layer2_outputs[9040] = ~(layer1_outputs[1178]);
    assign layer2_outputs[9041] = (layer1_outputs[6411]) ^ (layer1_outputs[9671]);
    assign layer2_outputs[9042] = (layer1_outputs[4555]) & ~(layer1_outputs[3881]);
    assign layer2_outputs[9043] = layer1_outputs[10224];
    assign layer2_outputs[9044] = (layer1_outputs[4679]) & ~(layer1_outputs[12637]);
    assign layer2_outputs[9045] = layer1_outputs[935];
    assign layer2_outputs[9046] = ~(layer1_outputs[4816]);
    assign layer2_outputs[9047] = (layer1_outputs[3881]) | (layer1_outputs[11081]);
    assign layer2_outputs[9048] = (layer1_outputs[4092]) | (layer1_outputs[4403]);
    assign layer2_outputs[9049] = layer1_outputs[7596];
    assign layer2_outputs[9050] = ~(layer1_outputs[3083]);
    assign layer2_outputs[9051] = (layer1_outputs[5400]) & (layer1_outputs[9876]);
    assign layer2_outputs[9052] = layer1_outputs[12489];
    assign layer2_outputs[9053] = ~(layer1_outputs[10737]);
    assign layer2_outputs[9054] = ~(layer1_outputs[904]);
    assign layer2_outputs[9055] = ~(layer1_outputs[12626]);
    assign layer2_outputs[9056] = ~((layer1_outputs[3258]) | (layer1_outputs[6817]));
    assign layer2_outputs[9057] = ~(layer1_outputs[2813]);
    assign layer2_outputs[9058] = layer1_outputs[1945];
    assign layer2_outputs[9059] = layer1_outputs[6765];
    assign layer2_outputs[9060] = ~(layer1_outputs[4837]);
    assign layer2_outputs[9061] = (layer1_outputs[10711]) & ~(layer1_outputs[9708]);
    assign layer2_outputs[9062] = ~((layer1_outputs[4123]) & (layer1_outputs[6898]));
    assign layer2_outputs[9063] = ~(layer1_outputs[7042]);
    assign layer2_outputs[9064] = ~(layer1_outputs[1587]);
    assign layer2_outputs[9065] = (layer1_outputs[3539]) & (layer1_outputs[10051]);
    assign layer2_outputs[9066] = ~(layer1_outputs[5222]);
    assign layer2_outputs[9067] = (layer1_outputs[11778]) ^ (layer1_outputs[2105]);
    assign layer2_outputs[9068] = ~((layer1_outputs[2107]) & (layer1_outputs[2103]));
    assign layer2_outputs[9069] = ~(layer1_outputs[8475]) | (layer1_outputs[3059]);
    assign layer2_outputs[9070] = ~((layer1_outputs[1250]) & (layer1_outputs[6745]));
    assign layer2_outputs[9071] = ~(layer1_outputs[10874]) | (layer1_outputs[9002]);
    assign layer2_outputs[9072] = (layer1_outputs[9546]) & ~(layer1_outputs[1956]);
    assign layer2_outputs[9073] = layer1_outputs[11209];
    assign layer2_outputs[9074] = (layer1_outputs[3389]) ^ (layer1_outputs[8670]);
    assign layer2_outputs[9075] = ~(layer1_outputs[8922]);
    assign layer2_outputs[9076] = (layer1_outputs[7139]) ^ (layer1_outputs[2043]);
    assign layer2_outputs[9077] = (layer1_outputs[8599]) ^ (layer1_outputs[6408]);
    assign layer2_outputs[9078] = (layer1_outputs[12642]) & ~(layer1_outputs[5269]);
    assign layer2_outputs[9079] = ~(layer1_outputs[3403]);
    assign layer2_outputs[9080] = layer1_outputs[51];
    assign layer2_outputs[9081] = (layer1_outputs[5224]) & ~(layer1_outputs[6136]);
    assign layer2_outputs[9082] = ~(layer1_outputs[6988]);
    assign layer2_outputs[9083] = ~(layer1_outputs[6188]);
    assign layer2_outputs[9084] = ~((layer1_outputs[1088]) | (layer1_outputs[4370]));
    assign layer2_outputs[9085] = ~((layer1_outputs[9133]) & (layer1_outputs[1350]));
    assign layer2_outputs[9086] = (layer1_outputs[2026]) | (layer1_outputs[7268]);
    assign layer2_outputs[9087] = ~(layer1_outputs[3378]) | (layer1_outputs[4805]);
    assign layer2_outputs[9088] = ~((layer1_outputs[8342]) ^ (layer1_outputs[8077]));
    assign layer2_outputs[9089] = (layer1_outputs[1267]) & (layer1_outputs[5781]);
    assign layer2_outputs[9090] = (layer1_outputs[3912]) & (layer1_outputs[12502]);
    assign layer2_outputs[9091] = layer1_outputs[10026];
    assign layer2_outputs[9092] = layer1_outputs[4284];
    assign layer2_outputs[9093] = layer1_outputs[7806];
    assign layer2_outputs[9094] = (layer1_outputs[5014]) & ~(layer1_outputs[5238]);
    assign layer2_outputs[9095] = (layer1_outputs[10183]) ^ (layer1_outputs[5716]);
    assign layer2_outputs[9096] = ~(layer1_outputs[11178]);
    assign layer2_outputs[9097] = layer1_outputs[2200];
    assign layer2_outputs[9098] = (layer1_outputs[623]) & ~(layer1_outputs[7997]);
    assign layer2_outputs[9099] = (layer1_outputs[1110]) & ~(layer1_outputs[6054]);
    assign layer2_outputs[9100] = (layer1_outputs[7252]) | (layer1_outputs[12429]);
    assign layer2_outputs[9101] = ~(layer1_outputs[445]);
    assign layer2_outputs[9102] = layer1_outputs[10007];
    assign layer2_outputs[9103] = layer1_outputs[11005];
    assign layer2_outputs[9104] = ~(layer1_outputs[1997]);
    assign layer2_outputs[9105] = layer1_outputs[1235];
    assign layer2_outputs[9106] = ~(layer1_outputs[12551]);
    assign layer2_outputs[9107] = (layer1_outputs[2160]) & ~(layer1_outputs[8664]);
    assign layer2_outputs[9108] = ~(layer1_outputs[8341]);
    assign layer2_outputs[9109] = (layer1_outputs[7283]) & ~(layer1_outputs[9702]);
    assign layer2_outputs[9110] = layer1_outputs[6299];
    assign layer2_outputs[9111] = layer1_outputs[1005];
    assign layer2_outputs[9112] = layer1_outputs[6927];
    assign layer2_outputs[9113] = (layer1_outputs[8570]) & ~(layer1_outputs[11004]);
    assign layer2_outputs[9114] = ~(layer1_outputs[3268]);
    assign layer2_outputs[9115] = ~((layer1_outputs[11125]) & (layer1_outputs[4205]));
    assign layer2_outputs[9116] = (layer1_outputs[845]) & ~(layer1_outputs[12629]);
    assign layer2_outputs[9117] = layer1_outputs[7087];
    assign layer2_outputs[9118] = ~((layer1_outputs[12331]) | (layer1_outputs[6755]));
    assign layer2_outputs[9119] = ~(layer1_outputs[2713]);
    assign layer2_outputs[9120] = ~(layer1_outputs[5262]) | (layer1_outputs[4892]);
    assign layer2_outputs[9121] = ~(layer1_outputs[4258]) | (layer1_outputs[4808]);
    assign layer2_outputs[9122] = layer1_outputs[3941];
    assign layer2_outputs[9123] = layer1_outputs[6052];
    assign layer2_outputs[9124] = ~(layer1_outputs[8138]);
    assign layer2_outputs[9125] = ~(layer1_outputs[4890]);
    assign layer2_outputs[9126] = ~((layer1_outputs[6928]) & (layer1_outputs[10027]));
    assign layer2_outputs[9127] = (layer1_outputs[9521]) ^ (layer1_outputs[7264]);
    assign layer2_outputs[9128] = ~((layer1_outputs[7511]) ^ (layer1_outputs[2119]));
    assign layer2_outputs[9129] = layer1_outputs[4324];
    assign layer2_outputs[9130] = ~(layer1_outputs[6078]);
    assign layer2_outputs[9131] = layer1_outputs[9167];
    assign layer2_outputs[9132] = ~(layer1_outputs[326]);
    assign layer2_outputs[9133] = layer1_outputs[11947];
    assign layer2_outputs[9134] = (layer1_outputs[8530]) ^ (layer1_outputs[9396]);
    assign layer2_outputs[9135] = (layer1_outputs[4616]) & (layer1_outputs[3265]);
    assign layer2_outputs[9136] = (layer1_outputs[10651]) | (layer1_outputs[11612]);
    assign layer2_outputs[9137] = ~(layer1_outputs[11286]) | (layer1_outputs[10025]);
    assign layer2_outputs[9138] = ~(layer1_outputs[12011]) | (layer1_outputs[2720]);
    assign layer2_outputs[9139] = ~(layer1_outputs[4027]);
    assign layer2_outputs[9140] = (layer1_outputs[2860]) ^ (layer1_outputs[9811]);
    assign layer2_outputs[9141] = ~((layer1_outputs[2326]) & (layer1_outputs[8802]));
    assign layer2_outputs[9142] = (layer1_outputs[11463]) & ~(layer1_outputs[6052]);
    assign layer2_outputs[9143] = (layer1_outputs[12331]) & ~(layer1_outputs[6275]);
    assign layer2_outputs[9144] = ~(layer1_outputs[11038]);
    assign layer2_outputs[9145] = layer1_outputs[5403];
    assign layer2_outputs[9146] = ~(layer1_outputs[10174]);
    assign layer2_outputs[9147] = (layer1_outputs[12689]) & (layer1_outputs[749]);
    assign layer2_outputs[9148] = ~((layer1_outputs[3691]) ^ (layer1_outputs[3014]));
    assign layer2_outputs[9149] = layer1_outputs[1435];
    assign layer2_outputs[9150] = layer1_outputs[6432];
    assign layer2_outputs[9151] = layer1_outputs[1253];
    assign layer2_outputs[9152] = ~((layer1_outputs[1624]) ^ (layer1_outputs[9269]));
    assign layer2_outputs[9153] = layer1_outputs[6103];
    assign layer2_outputs[9154] = ~((layer1_outputs[1354]) ^ (layer1_outputs[714]));
    assign layer2_outputs[9155] = ~(layer1_outputs[4287]) | (layer1_outputs[9701]);
    assign layer2_outputs[9156] = ~((layer1_outputs[2597]) ^ (layer1_outputs[1968]));
    assign layer2_outputs[9157] = layer1_outputs[1004];
    assign layer2_outputs[9158] = (layer1_outputs[2110]) & ~(layer1_outputs[3046]);
    assign layer2_outputs[9159] = (layer1_outputs[8695]) & ~(layer1_outputs[12365]);
    assign layer2_outputs[9160] = layer1_outputs[10119];
    assign layer2_outputs[9161] = (layer1_outputs[11048]) & (layer1_outputs[9824]);
    assign layer2_outputs[9162] = (layer1_outputs[3161]) & ~(layer1_outputs[109]);
    assign layer2_outputs[9163] = layer1_outputs[3741];
    assign layer2_outputs[9164] = ~(layer1_outputs[1145]);
    assign layer2_outputs[9165] = ~(layer1_outputs[6347]);
    assign layer2_outputs[9166] = ~(layer1_outputs[9257]);
    assign layer2_outputs[9167] = layer1_outputs[544];
    assign layer2_outputs[9168] = (layer1_outputs[9981]) ^ (layer1_outputs[7774]);
    assign layer2_outputs[9169] = (layer1_outputs[597]) & ~(layer1_outputs[2370]);
    assign layer2_outputs[9170] = ~(layer1_outputs[8760]);
    assign layer2_outputs[9171] = layer1_outputs[1327];
    assign layer2_outputs[9172] = ~((layer1_outputs[7028]) ^ (layer1_outputs[9660]));
    assign layer2_outputs[9173] = (layer1_outputs[80]) & ~(layer1_outputs[5034]);
    assign layer2_outputs[9174] = layer1_outputs[9077];
    assign layer2_outputs[9175] = ~(layer1_outputs[2975]);
    assign layer2_outputs[9176] = layer1_outputs[6083];
    assign layer2_outputs[9177] = layer1_outputs[8467];
    assign layer2_outputs[9178] = (layer1_outputs[5718]) ^ (layer1_outputs[10171]);
    assign layer2_outputs[9179] = ~(layer1_outputs[1363]);
    assign layer2_outputs[9180] = ~(layer1_outputs[7706]);
    assign layer2_outputs[9181] = (layer1_outputs[2081]) & (layer1_outputs[5097]);
    assign layer2_outputs[9182] = ~((layer1_outputs[9178]) ^ (layer1_outputs[7973]));
    assign layer2_outputs[9183] = (layer1_outputs[9880]) | (layer1_outputs[4466]);
    assign layer2_outputs[9184] = ~(layer1_outputs[7335]);
    assign layer2_outputs[9185] = ~(layer1_outputs[6768]);
    assign layer2_outputs[9186] = layer1_outputs[4673];
    assign layer2_outputs[9187] = ~((layer1_outputs[7197]) & (layer1_outputs[3846]));
    assign layer2_outputs[9188] = (layer1_outputs[10695]) & ~(layer1_outputs[3351]);
    assign layer2_outputs[9189] = layer1_outputs[9069];
    assign layer2_outputs[9190] = ~(layer1_outputs[7055]);
    assign layer2_outputs[9191] = layer1_outputs[3472];
    assign layer2_outputs[9192] = ~((layer1_outputs[2097]) ^ (layer1_outputs[3357]));
    assign layer2_outputs[9193] = layer1_outputs[12701];
    assign layer2_outputs[9194] = (layer1_outputs[3730]) & (layer1_outputs[3415]);
    assign layer2_outputs[9195] = ~((layer1_outputs[11530]) ^ (layer1_outputs[12534]));
    assign layer2_outputs[9196] = 1'b1;
    assign layer2_outputs[9197] = layer1_outputs[5705];
    assign layer2_outputs[9198] = ~(layer1_outputs[3309]);
    assign layer2_outputs[9199] = (layer1_outputs[12747]) | (layer1_outputs[9944]);
    assign layer2_outputs[9200] = ~(layer1_outputs[6194]);
    assign layer2_outputs[9201] = layer1_outputs[4807];
    assign layer2_outputs[9202] = ~(layer1_outputs[1824]);
    assign layer2_outputs[9203] = ~(layer1_outputs[2312]);
    assign layer2_outputs[9204] = ~(layer1_outputs[10295]);
    assign layer2_outputs[9205] = ~(layer1_outputs[1378]);
    assign layer2_outputs[9206] = ~(layer1_outputs[6521]);
    assign layer2_outputs[9207] = ~((layer1_outputs[12048]) & (layer1_outputs[11583]));
    assign layer2_outputs[9208] = ~(layer1_outputs[9503]) | (layer1_outputs[6827]);
    assign layer2_outputs[9209] = (layer1_outputs[4969]) & (layer1_outputs[3151]);
    assign layer2_outputs[9210] = ~(layer1_outputs[12209]);
    assign layer2_outputs[9211] = ~((layer1_outputs[4034]) & (layer1_outputs[2730]));
    assign layer2_outputs[9212] = layer1_outputs[543];
    assign layer2_outputs[9213] = ~((layer1_outputs[4109]) | (layer1_outputs[538]));
    assign layer2_outputs[9214] = layer1_outputs[11676];
    assign layer2_outputs[9215] = ~(layer1_outputs[3511]) | (layer1_outputs[8004]);
    assign layer2_outputs[9216] = ~(layer1_outputs[5676]) | (layer1_outputs[2838]);
    assign layer2_outputs[9217] = ~(layer1_outputs[2688]);
    assign layer2_outputs[9218] = ~(layer1_outputs[7049]) | (layer1_outputs[3908]);
    assign layer2_outputs[9219] = layer1_outputs[5248];
    assign layer2_outputs[9220] = ~((layer1_outputs[10572]) | (layer1_outputs[6223]));
    assign layer2_outputs[9221] = (layer1_outputs[12087]) & (layer1_outputs[10109]);
    assign layer2_outputs[9222] = layer1_outputs[6917];
    assign layer2_outputs[9223] = ~(layer1_outputs[8804]) | (layer1_outputs[9438]);
    assign layer2_outputs[9224] = ~(layer1_outputs[9866]) | (layer1_outputs[8174]);
    assign layer2_outputs[9225] = ~((layer1_outputs[8793]) ^ (layer1_outputs[1976]));
    assign layer2_outputs[9226] = (layer1_outputs[7245]) ^ (layer1_outputs[5014]);
    assign layer2_outputs[9227] = (layer1_outputs[4811]) & (layer1_outputs[66]);
    assign layer2_outputs[9228] = ~(layer1_outputs[12240]);
    assign layer2_outputs[9229] = (layer1_outputs[9957]) & ~(layer1_outputs[2734]);
    assign layer2_outputs[9230] = layer1_outputs[12030];
    assign layer2_outputs[9231] = ~((layer1_outputs[3315]) & (layer1_outputs[2275]));
    assign layer2_outputs[9232] = layer1_outputs[11095];
    assign layer2_outputs[9233] = ~(layer1_outputs[4700]);
    assign layer2_outputs[9234] = ~((layer1_outputs[10644]) | (layer1_outputs[2623]));
    assign layer2_outputs[9235] = ~((layer1_outputs[12412]) | (layer1_outputs[2969]));
    assign layer2_outputs[9236] = 1'b0;
    assign layer2_outputs[9237] = ~((layer1_outputs[6614]) ^ (layer1_outputs[4923]));
    assign layer2_outputs[9238] = (layer1_outputs[660]) & ~(layer1_outputs[6870]);
    assign layer2_outputs[9239] = (layer1_outputs[12638]) | (layer1_outputs[5620]);
    assign layer2_outputs[9240] = (layer1_outputs[554]) & (layer1_outputs[2647]);
    assign layer2_outputs[9241] = layer1_outputs[2518];
    assign layer2_outputs[9242] = ~((layer1_outputs[8715]) ^ (layer1_outputs[915]));
    assign layer2_outputs[9243] = ~(layer1_outputs[4523]);
    assign layer2_outputs[9244] = ~((layer1_outputs[3242]) ^ (layer1_outputs[7450]));
    assign layer2_outputs[9245] = (layer1_outputs[9183]) ^ (layer1_outputs[7151]);
    assign layer2_outputs[9246] = ~(layer1_outputs[5028]);
    assign layer2_outputs[9247] = ~(layer1_outputs[2620]);
    assign layer2_outputs[9248] = layer1_outputs[4736];
    assign layer2_outputs[9249] = layer1_outputs[4252];
    assign layer2_outputs[9250] = ~(layer1_outputs[11428]) | (layer1_outputs[9563]);
    assign layer2_outputs[9251] = ~((layer1_outputs[4821]) | (layer1_outputs[6028]));
    assign layer2_outputs[9252] = (layer1_outputs[7808]) | (layer1_outputs[9485]);
    assign layer2_outputs[9253] = ~(layer1_outputs[3002]);
    assign layer2_outputs[9254] = ~(layer1_outputs[9335]);
    assign layer2_outputs[9255] = ~(layer1_outputs[543]);
    assign layer2_outputs[9256] = layer1_outputs[8993];
    assign layer2_outputs[9257] = (layer1_outputs[4496]) & ~(layer1_outputs[5134]);
    assign layer2_outputs[9258] = layer1_outputs[210];
    assign layer2_outputs[9259] = ~(layer1_outputs[12167]);
    assign layer2_outputs[9260] = ~(layer1_outputs[10778]);
    assign layer2_outputs[9261] = layer1_outputs[7582];
    assign layer2_outputs[9262] = ~((layer1_outputs[8984]) & (layer1_outputs[11712]));
    assign layer2_outputs[9263] = (layer1_outputs[11607]) & (layer1_outputs[12368]);
    assign layer2_outputs[9264] = (layer1_outputs[7555]) | (layer1_outputs[4067]);
    assign layer2_outputs[9265] = ~(layer1_outputs[4166]);
    assign layer2_outputs[9266] = layer1_outputs[3451];
    assign layer2_outputs[9267] = ~((layer1_outputs[12001]) | (layer1_outputs[12384]));
    assign layer2_outputs[9268] = ~(layer1_outputs[9445]);
    assign layer2_outputs[9269] = ~(layer1_outputs[10055]);
    assign layer2_outputs[9270] = ~((layer1_outputs[12261]) & (layer1_outputs[5328]));
    assign layer2_outputs[9271] = (layer1_outputs[11415]) ^ (layer1_outputs[7691]);
    assign layer2_outputs[9272] = ~(layer1_outputs[12769]);
    assign layer2_outputs[9273] = (layer1_outputs[12056]) & ~(layer1_outputs[11073]);
    assign layer2_outputs[9274] = ~((layer1_outputs[1553]) ^ (layer1_outputs[6966]));
    assign layer2_outputs[9275] = (layer1_outputs[7422]) & ~(layer1_outputs[1941]);
    assign layer2_outputs[9276] = layer1_outputs[3400];
    assign layer2_outputs[9277] = (layer1_outputs[7927]) & ~(layer1_outputs[8518]);
    assign layer2_outputs[9278] = layer1_outputs[12500];
    assign layer2_outputs[9279] = (layer1_outputs[9804]) & ~(layer1_outputs[4736]);
    assign layer2_outputs[9280] = ~((layer1_outputs[3914]) & (layer1_outputs[2850]));
    assign layer2_outputs[9281] = (layer1_outputs[12489]) & (layer1_outputs[7529]);
    assign layer2_outputs[9282] = layer1_outputs[8802];
    assign layer2_outputs[9283] = ~((layer1_outputs[442]) & (layer1_outputs[11047]));
    assign layer2_outputs[9284] = (layer1_outputs[9924]) ^ (layer1_outputs[2263]);
    assign layer2_outputs[9285] = (layer1_outputs[7884]) | (layer1_outputs[5486]);
    assign layer2_outputs[9286] = layer1_outputs[6829];
    assign layer2_outputs[9287] = layer1_outputs[4297];
    assign layer2_outputs[9288] = ~(layer1_outputs[8253]) | (layer1_outputs[370]);
    assign layer2_outputs[9289] = ~(layer1_outputs[610]);
    assign layer2_outputs[9290] = ~((layer1_outputs[3917]) | (layer1_outputs[12494]));
    assign layer2_outputs[9291] = layer1_outputs[8609];
    assign layer2_outputs[9292] = layer1_outputs[5931];
    assign layer2_outputs[9293] = ~(layer1_outputs[10586]);
    assign layer2_outputs[9294] = ~(layer1_outputs[10394]) | (layer1_outputs[7508]);
    assign layer2_outputs[9295] = (layer1_outputs[7701]) ^ (layer1_outputs[1680]);
    assign layer2_outputs[9296] = (layer1_outputs[5416]) & ~(layer1_outputs[9728]);
    assign layer2_outputs[9297] = (layer1_outputs[8231]) | (layer1_outputs[1586]);
    assign layer2_outputs[9298] = ~(layer1_outputs[2432]) | (layer1_outputs[5407]);
    assign layer2_outputs[9299] = layer1_outputs[1874];
    assign layer2_outputs[9300] = layer1_outputs[9358];
    assign layer2_outputs[9301] = ~((layer1_outputs[6927]) ^ (layer1_outputs[11121]));
    assign layer2_outputs[9302] = (layer1_outputs[3134]) | (layer1_outputs[1090]);
    assign layer2_outputs[9303] = layer1_outputs[10488];
    assign layer2_outputs[9304] = layer1_outputs[4439];
    assign layer2_outputs[9305] = ~(layer1_outputs[9688]);
    assign layer2_outputs[9306] = layer1_outputs[277];
    assign layer2_outputs[9307] = (layer1_outputs[7325]) & ~(layer1_outputs[5666]);
    assign layer2_outputs[9308] = 1'b1;
    assign layer2_outputs[9309] = layer1_outputs[7131];
    assign layer2_outputs[9310] = ~(layer1_outputs[7220]);
    assign layer2_outputs[9311] = ~(layer1_outputs[5220]);
    assign layer2_outputs[9312] = (layer1_outputs[615]) ^ (layer1_outputs[11119]);
    assign layer2_outputs[9313] = ~((layer1_outputs[2334]) ^ (layer1_outputs[11284]));
    assign layer2_outputs[9314] = (layer1_outputs[3607]) | (layer1_outputs[1290]);
    assign layer2_outputs[9315] = layer1_outputs[10948];
    assign layer2_outputs[9316] = (layer1_outputs[9928]) ^ (layer1_outputs[3308]);
    assign layer2_outputs[9317] = layer1_outputs[12677];
    assign layer2_outputs[9318] = ~(layer1_outputs[8234]) | (layer1_outputs[2254]);
    assign layer2_outputs[9319] = layer1_outputs[6359];
    assign layer2_outputs[9320] = ~(layer1_outputs[4314]);
    assign layer2_outputs[9321] = ~((layer1_outputs[10362]) ^ (layer1_outputs[9927]));
    assign layer2_outputs[9322] = layer1_outputs[3960];
    assign layer2_outputs[9323] = layer1_outputs[11865];
    assign layer2_outputs[9324] = (layer1_outputs[2638]) | (layer1_outputs[2138]);
    assign layer2_outputs[9325] = ~((layer1_outputs[11903]) ^ (layer1_outputs[8356]));
    assign layer2_outputs[9326] = (layer1_outputs[430]) & ~(layer1_outputs[2016]);
    assign layer2_outputs[9327] = (layer1_outputs[3889]) & ~(layer1_outputs[3405]);
    assign layer2_outputs[9328] = layer1_outputs[2621];
    assign layer2_outputs[9329] = ~(layer1_outputs[12748]);
    assign layer2_outputs[9330] = (layer1_outputs[6265]) & ~(layer1_outputs[8433]);
    assign layer2_outputs[9331] = ~((layer1_outputs[10517]) | (layer1_outputs[3567]));
    assign layer2_outputs[9332] = ~(layer1_outputs[459]);
    assign layer2_outputs[9333] = ~(layer1_outputs[12452]);
    assign layer2_outputs[9334] = ~((layer1_outputs[10922]) & (layer1_outputs[11732]));
    assign layer2_outputs[9335] = layer1_outputs[2513];
    assign layer2_outputs[9336] = ~(layer1_outputs[10507]);
    assign layer2_outputs[9337] = (layer1_outputs[2798]) & (layer1_outputs[12342]);
    assign layer2_outputs[9338] = ~((layer1_outputs[7438]) ^ (layer1_outputs[9128]));
    assign layer2_outputs[9339] = ~(layer1_outputs[1194]);
    assign layer2_outputs[9340] = ~(layer1_outputs[2859]);
    assign layer2_outputs[9341] = layer1_outputs[10454];
    assign layer2_outputs[9342] = layer1_outputs[1968];
    assign layer2_outputs[9343] = (layer1_outputs[3235]) & ~(layer1_outputs[9120]);
    assign layer2_outputs[9344] = (layer1_outputs[4645]) & (layer1_outputs[4595]);
    assign layer2_outputs[9345] = ~(layer1_outputs[8468]) | (layer1_outputs[4280]);
    assign layer2_outputs[9346] = ~((layer1_outputs[6364]) & (layer1_outputs[8055]));
    assign layer2_outputs[9347] = layer1_outputs[9960];
    assign layer2_outputs[9348] = ~(layer1_outputs[3936]);
    assign layer2_outputs[9349] = ~(layer1_outputs[10747]);
    assign layer2_outputs[9350] = ~(layer1_outputs[1625]);
    assign layer2_outputs[9351] = layer1_outputs[6544];
    assign layer2_outputs[9352] = layer1_outputs[3883];
    assign layer2_outputs[9353] = (layer1_outputs[789]) & (layer1_outputs[4231]);
    assign layer2_outputs[9354] = ~((layer1_outputs[5459]) & (layer1_outputs[1245]));
    assign layer2_outputs[9355] = ~(layer1_outputs[2609]);
    assign layer2_outputs[9356] = (layer1_outputs[7069]) & ~(layer1_outputs[3217]);
    assign layer2_outputs[9357] = ~((layer1_outputs[10557]) ^ (layer1_outputs[3933]));
    assign layer2_outputs[9358] = layer1_outputs[5993];
    assign layer2_outputs[9359] = ~(layer1_outputs[10958]);
    assign layer2_outputs[9360] = layer1_outputs[7451];
    assign layer2_outputs[9361] = ~(layer1_outputs[11821]);
    assign layer2_outputs[9362] = (layer1_outputs[10353]) & ~(layer1_outputs[6813]);
    assign layer2_outputs[9363] = ~(layer1_outputs[7775]);
    assign layer2_outputs[9364] = 1'b1;
    assign layer2_outputs[9365] = ~((layer1_outputs[12593]) & (layer1_outputs[6968]));
    assign layer2_outputs[9366] = layer1_outputs[10626];
    assign layer2_outputs[9367] = ~(layer1_outputs[1212]);
    assign layer2_outputs[9368] = ~((layer1_outputs[1508]) ^ (layer1_outputs[2029]));
    assign layer2_outputs[9369] = layer1_outputs[11528];
    assign layer2_outputs[9370] = (layer1_outputs[8363]) | (layer1_outputs[7676]);
    assign layer2_outputs[9371] = ~(layer1_outputs[2418]) | (layer1_outputs[2127]);
    assign layer2_outputs[9372] = layer1_outputs[225];
    assign layer2_outputs[9373] = ~(layer1_outputs[10037]);
    assign layer2_outputs[9374] = ~((layer1_outputs[359]) ^ (layer1_outputs[5235]));
    assign layer2_outputs[9375] = (layer1_outputs[279]) ^ (layer1_outputs[11035]);
    assign layer2_outputs[9376] = (layer1_outputs[8588]) | (layer1_outputs[19]);
    assign layer2_outputs[9377] = ~(layer1_outputs[11572]);
    assign layer2_outputs[9378] = ~(layer1_outputs[8650]);
    assign layer2_outputs[9379] = layer1_outputs[6045];
    assign layer2_outputs[9380] = ~((layer1_outputs[1087]) ^ (layer1_outputs[3933]));
    assign layer2_outputs[9381] = (layer1_outputs[12657]) & (layer1_outputs[9447]);
    assign layer2_outputs[9382] = ~((layer1_outputs[4422]) ^ (layer1_outputs[11418]));
    assign layer2_outputs[9383] = layer1_outputs[4780];
    assign layer2_outputs[9384] = 1'b1;
    assign layer2_outputs[9385] = ~(layer1_outputs[12653]);
    assign layer2_outputs[9386] = ~((layer1_outputs[6104]) & (layer1_outputs[3326]));
    assign layer2_outputs[9387] = ~((layer1_outputs[11216]) ^ (layer1_outputs[12315]));
    assign layer2_outputs[9388] = 1'b0;
    assign layer2_outputs[9389] = (layer1_outputs[7741]) & ~(layer1_outputs[8963]);
    assign layer2_outputs[9390] = layer1_outputs[9863];
    assign layer2_outputs[9391] = layer1_outputs[8209];
    assign layer2_outputs[9392] = layer1_outputs[12517];
    assign layer2_outputs[9393] = ~(layer1_outputs[1785]);
    assign layer2_outputs[9394] = layer1_outputs[5482];
    assign layer2_outputs[9395] = layer1_outputs[9535];
    assign layer2_outputs[9396] = layer1_outputs[9742];
    assign layer2_outputs[9397] = ~(layer1_outputs[3469]);
    assign layer2_outputs[9398] = (layer1_outputs[5876]) ^ (layer1_outputs[7140]);
    assign layer2_outputs[9399] = (layer1_outputs[11029]) & ~(layer1_outputs[12711]);
    assign layer2_outputs[9400] = layer1_outputs[4782];
    assign layer2_outputs[9401] = (layer1_outputs[10895]) ^ (layer1_outputs[4667]);
    assign layer2_outputs[9402] = ~((layer1_outputs[4952]) ^ (layer1_outputs[3864]));
    assign layer2_outputs[9403] = (layer1_outputs[6804]) & ~(layer1_outputs[3720]);
    assign layer2_outputs[9404] = (layer1_outputs[220]) ^ (layer1_outputs[2778]);
    assign layer2_outputs[9405] = ~(layer1_outputs[778]);
    assign layer2_outputs[9406] = layer1_outputs[12792];
    assign layer2_outputs[9407] = ~((layer1_outputs[9115]) | (layer1_outputs[11239]));
    assign layer2_outputs[9408] = (layer1_outputs[516]) | (layer1_outputs[12020]);
    assign layer2_outputs[9409] = ~((layer1_outputs[12447]) ^ (layer1_outputs[5663]));
    assign layer2_outputs[9410] = ~(layer1_outputs[4857]);
    assign layer2_outputs[9411] = (layer1_outputs[10659]) & ~(layer1_outputs[5873]);
    assign layer2_outputs[9412] = (layer1_outputs[6086]) & ~(layer1_outputs[669]);
    assign layer2_outputs[9413] = layer1_outputs[7718];
    assign layer2_outputs[9414] = (layer1_outputs[11302]) & ~(layer1_outputs[5832]);
    assign layer2_outputs[9415] = layer1_outputs[2199];
    assign layer2_outputs[9416] = ~((layer1_outputs[5038]) ^ (layer1_outputs[2618]));
    assign layer2_outputs[9417] = layer1_outputs[3464];
    assign layer2_outputs[9418] = ~(layer1_outputs[10371]);
    assign layer2_outputs[9419] = (layer1_outputs[8814]) & ~(layer1_outputs[4651]);
    assign layer2_outputs[9420] = (layer1_outputs[11146]) & ~(layer1_outputs[461]);
    assign layer2_outputs[9421] = ~((layer1_outputs[2151]) ^ (layer1_outputs[8909]));
    assign layer2_outputs[9422] = (layer1_outputs[17]) & ~(layer1_outputs[11150]);
    assign layer2_outputs[9423] = (layer1_outputs[12791]) ^ (layer1_outputs[2961]);
    assign layer2_outputs[9424] = ~((layer1_outputs[1618]) & (layer1_outputs[7149]));
    assign layer2_outputs[9425] = (layer1_outputs[10075]) ^ (layer1_outputs[3087]);
    assign layer2_outputs[9426] = ~(layer1_outputs[6170]) | (layer1_outputs[10429]);
    assign layer2_outputs[9427] = ~(layer1_outputs[11742]);
    assign layer2_outputs[9428] = ~((layer1_outputs[5377]) & (layer1_outputs[8702]));
    assign layer2_outputs[9429] = (layer1_outputs[2297]) & ~(layer1_outputs[8727]);
    assign layer2_outputs[9430] = (layer1_outputs[1556]) & ~(layer1_outputs[770]);
    assign layer2_outputs[9431] = ~((layer1_outputs[7484]) ^ (layer1_outputs[8583]));
    assign layer2_outputs[9432] = layer1_outputs[6262];
    assign layer2_outputs[9433] = (layer1_outputs[8278]) ^ (layer1_outputs[1417]);
    assign layer2_outputs[9434] = ~(layer1_outputs[10559]);
    assign layer2_outputs[9435] = ~(layer1_outputs[11610]);
    assign layer2_outputs[9436] = (layer1_outputs[5754]) & (layer1_outputs[11621]);
    assign layer2_outputs[9437] = 1'b0;
    assign layer2_outputs[9438] = (layer1_outputs[11218]) & ~(layer1_outputs[1323]);
    assign layer2_outputs[9439] = ~(layer1_outputs[12613]);
    assign layer2_outputs[9440] = 1'b1;
    assign layer2_outputs[9441] = ~(layer1_outputs[9542]);
    assign layer2_outputs[9442] = (layer1_outputs[6210]) & (layer1_outputs[2442]);
    assign layer2_outputs[9443] = layer1_outputs[7992];
    assign layer2_outputs[9444] = (layer1_outputs[10969]) ^ (layer1_outputs[3484]);
    assign layer2_outputs[9445] = layer1_outputs[5375];
    assign layer2_outputs[9446] = (layer1_outputs[6466]) & (layer1_outputs[7838]);
    assign layer2_outputs[9447] = (layer1_outputs[1121]) ^ (layer1_outputs[11096]);
    assign layer2_outputs[9448] = ~(layer1_outputs[10039]);
    assign layer2_outputs[9449] = (layer1_outputs[1057]) | (layer1_outputs[9992]);
    assign layer2_outputs[9450] = layer1_outputs[8059];
    assign layer2_outputs[9451] = ~(layer1_outputs[12546]);
    assign layer2_outputs[9452] = layer1_outputs[3819];
    assign layer2_outputs[9453] = ~((layer1_outputs[9810]) | (layer1_outputs[9835]));
    assign layer2_outputs[9454] = ~(layer1_outputs[11789]);
    assign layer2_outputs[9455] = (layer1_outputs[10798]) ^ (layer1_outputs[10068]);
    assign layer2_outputs[9456] = ~(layer1_outputs[4756]);
    assign layer2_outputs[9457] = ~((layer1_outputs[11318]) & (layer1_outputs[7943]));
    assign layer2_outputs[9458] = ~(layer1_outputs[10956]) | (layer1_outputs[4940]);
    assign layer2_outputs[9459] = layer1_outputs[10415];
    assign layer2_outputs[9460] = layer1_outputs[7137];
    assign layer2_outputs[9461] = ~((layer1_outputs[2635]) & (layer1_outputs[11787]));
    assign layer2_outputs[9462] = ~((layer1_outputs[335]) ^ (layer1_outputs[11076]));
    assign layer2_outputs[9463] = (layer1_outputs[6648]) & ~(layer1_outputs[6083]);
    assign layer2_outputs[9464] = (layer1_outputs[1751]) & (layer1_outputs[2643]);
    assign layer2_outputs[9465] = (layer1_outputs[10863]) ^ (layer1_outputs[8175]);
    assign layer2_outputs[9466] = ~(layer1_outputs[3471]);
    assign layer2_outputs[9467] = (layer1_outputs[236]) ^ (layer1_outputs[4630]);
    assign layer2_outputs[9468] = (layer1_outputs[617]) ^ (layer1_outputs[7423]);
    assign layer2_outputs[9469] = layer1_outputs[5157];
    assign layer2_outputs[9470] = ~((layer1_outputs[7593]) & (layer1_outputs[6477]));
    assign layer2_outputs[9471] = layer1_outputs[6251];
    assign layer2_outputs[9472] = layer1_outputs[3296];
    assign layer2_outputs[9473] = ~(layer1_outputs[7006]);
    assign layer2_outputs[9474] = (layer1_outputs[737]) ^ (layer1_outputs[6026]);
    assign layer2_outputs[9475] = ~(layer1_outputs[10104]);
    assign layer2_outputs[9476] = ~(layer1_outputs[2187]);
    assign layer2_outputs[9477] = (layer1_outputs[9367]) & (layer1_outputs[11871]);
    assign layer2_outputs[9478] = (layer1_outputs[8679]) | (layer1_outputs[6436]);
    assign layer2_outputs[9479] = ~((layer1_outputs[4489]) & (layer1_outputs[9256]));
    assign layer2_outputs[9480] = (layer1_outputs[6991]) ^ (layer1_outputs[924]);
    assign layer2_outputs[9481] = ~(layer1_outputs[1573]);
    assign layer2_outputs[9482] = layer1_outputs[4];
    assign layer2_outputs[9483] = ~(layer1_outputs[10072]);
    assign layer2_outputs[9484] = ~(layer1_outputs[2277]);
    assign layer2_outputs[9485] = ~(layer1_outputs[2105]) | (layer1_outputs[9803]);
    assign layer2_outputs[9486] = layer1_outputs[6165];
    assign layer2_outputs[9487] = ~(layer1_outputs[2052]);
    assign layer2_outputs[9488] = layer1_outputs[2444];
    assign layer2_outputs[9489] = ~(layer1_outputs[6894]);
    assign layer2_outputs[9490] = ~(layer1_outputs[11124]) | (layer1_outputs[2643]);
    assign layer2_outputs[9491] = (layer1_outputs[6245]) ^ (layer1_outputs[2752]);
    assign layer2_outputs[9492] = layer1_outputs[5693];
    assign layer2_outputs[9493] = (layer1_outputs[2207]) | (layer1_outputs[2529]);
    assign layer2_outputs[9494] = ~((layer1_outputs[6641]) & (layer1_outputs[10377]));
    assign layer2_outputs[9495] = (layer1_outputs[8197]) ^ (layer1_outputs[892]);
    assign layer2_outputs[9496] = layer1_outputs[6282];
    assign layer2_outputs[9497] = (layer1_outputs[9671]) & ~(layer1_outputs[9287]);
    assign layer2_outputs[9498] = ~(layer1_outputs[885]) | (layer1_outputs[3310]);
    assign layer2_outputs[9499] = layer1_outputs[7299];
    assign layer2_outputs[9500] = (layer1_outputs[5089]) & (layer1_outputs[9881]);
    assign layer2_outputs[9501] = (layer1_outputs[8966]) & (layer1_outputs[3776]);
    assign layer2_outputs[9502] = layer1_outputs[2804];
    assign layer2_outputs[9503] = ~(layer1_outputs[4771]);
    assign layer2_outputs[9504] = ~((layer1_outputs[8655]) | (layer1_outputs[5162]));
    assign layer2_outputs[9505] = ~(layer1_outputs[1140]) | (layer1_outputs[7030]);
    assign layer2_outputs[9506] = layer1_outputs[7834];
    assign layer2_outputs[9507] = (layer1_outputs[11845]) & ~(layer1_outputs[11339]);
    assign layer2_outputs[9508] = ~((layer1_outputs[8812]) & (layer1_outputs[1272]));
    assign layer2_outputs[9509] = ~((layer1_outputs[9761]) | (layer1_outputs[1624]));
    assign layer2_outputs[9510] = layer1_outputs[10411];
    assign layer2_outputs[9511] = layer1_outputs[1945];
    assign layer2_outputs[9512] = ~((layer1_outputs[3890]) & (layer1_outputs[12752]));
    assign layer2_outputs[9513] = layer1_outputs[5445];
    assign layer2_outputs[9514] = ~(layer1_outputs[11637]);
    assign layer2_outputs[9515] = (layer1_outputs[8916]) & (layer1_outputs[6453]);
    assign layer2_outputs[9516] = (layer1_outputs[10352]) ^ (layer1_outputs[7679]);
    assign layer2_outputs[9517] = ~(layer1_outputs[9649]) | (layer1_outputs[9215]);
    assign layer2_outputs[9518] = layer1_outputs[4453];
    assign layer2_outputs[9519] = ~(layer1_outputs[10237]);
    assign layer2_outputs[9520] = layer1_outputs[1010];
    assign layer2_outputs[9521] = layer1_outputs[11956];
    assign layer2_outputs[9522] = layer1_outputs[5492];
    assign layer2_outputs[9523] = (layer1_outputs[3817]) & (layer1_outputs[5864]);
    assign layer2_outputs[9524] = ~((layer1_outputs[8534]) & (layer1_outputs[2979]));
    assign layer2_outputs[9525] = ~(layer1_outputs[9178]);
    assign layer2_outputs[9526] = ~(layer1_outputs[3657]);
    assign layer2_outputs[9527] = layer1_outputs[6497];
    assign layer2_outputs[9528] = ~(layer1_outputs[6963]) | (layer1_outputs[3148]);
    assign layer2_outputs[9529] = ~(layer1_outputs[1914]);
    assign layer2_outputs[9530] = (layer1_outputs[2211]) ^ (layer1_outputs[12793]);
    assign layer2_outputs[9531] = ~(layer1_outputs[11877]);
    assign layer2_outputs[9532] = ~(layer1_outputs[5167]) | (layer1_outputs[4768]);
    assign layer2_outputs[9533] = (layer1_outputs[12388]) & ~(layer1_outputs[8249]);
    assign layer2_outputs[9534] = ~(layer1_outputs[5824]);
    assign layer2_outputs[9535] = ~(layer1_outputs[8184]);
    assign layer2_outputs[9536] = layer1_outputs[12720];
    assign layer2_outputs[9537] = ~(layer1_outputs[4822]);
    assign layer2_outputs[9538] = (layer1_outputs[2176]) ^ (layer1_outputs[5025]);
    assign layer2_outputs[9539] = layer1_outputs[12664];
    assign layer2_outputs[9540] = ~(layer1_outputs[5948]);
    assign layer2_outputs[9541] = ~(layer1_outputs[8911]) | (layer1_outputs[4441]);
    assign layer2_outputs[9542] = ~((layer1_outputs[7341]) | (layer1_outputs[9190]));
    assign layer2_outputs[9543] = layer1_outputs[12087];
    assign layer2_outputs[9544] = (layer1_outputs[11981]) | (layer1_outputs[12348]);
    assign layer2_outputs[9545] = ~((layer1_outputs[5103]) | (layer1_outputs[10843]));
    assign layer2_outputs[9546] = (layer1_outputs[7211]) ^ (layer1_outputs[12366]);
    assign layer2_outputs[9547] = layer1_outputs[2413];
    assign layer2_outputs[9548] = (layer1_outputs[2226]) ^ (layer1_outputs[4592]);
    assign layer2_outputs[9549] = ~(layer1_outputs[3777]);
    assign layer2_outputs[9550] = (layer1_outputs[10067]) & ~(layer1_outputs[10005]);
    assign layer2_outputs[9551] = (layer1_outputs[7486]) ^ (layer1_outputs[2964]);
    assign layer2_outputs[9552] = layer1_outputs[7982];
    assign layer2_outputs[9553] = layer1_outputs[9243];
    assign layer2_outputs[9554] = ~(layer1_outputs[9991]);
    assign layer2_outputs[9555] = layer1_outputs[3761];
    assign layer2_outputs[9556] = (layer1_outputs[6237]) & ~(layer1_outputs[11872]);
    assign layer2_outputs[9557] = (layer1_outputs[11476]) ^ (layer1_outputs[8449]);
    assign layer2_outputs[9558] = ~(layer1_outputs[2785]);
    assign layer2_outputs[9559] = layer1_outputs[3033];
    assign layer2_outputs[9560] = ~(layer1_outputs[5147]);
    assign layer2_outputs[9561] = layer1_outputs[11218];
    assign layer2_outputs[9562] = ~((layer1_outputs[6219]) & (layer1_outputs[12648]));
    assign layer2_outputs[9563] = (layer1_outputs[11523]) ^ (layer1_outputs[12623]);
    assign layer2_outputs[9564] = ~(layer1_outputs[12279]);
    assign layer2_outputs[9565] = ~(layer1_outputs[2475]);
    assign layer2_outputs[9566] = (layer1_outputs[12213]) & ~(layer1_outputs[8983]);
    assign layer2_outputs[9567] = ~((layer1_outputs[11718]) | (layer1_outputs[6513]));
    assign layer2_outputs[9568] = layer1_outputs[4506];
    assign layer2_outputs[9569] = layer1_outputs[3695];
    assign layer2_outputs[9570] = ~(layer1_outputs[2610]) | (layer1_outputs[5188]);
    assign layer2_outputs[9571] = ~(layer1_outputs[7604]) | (layer1_outputs[2773]);
    assign layer2_outputs[9572] = ~(layer1_outputs[10219]);
    assign layer2_outputs[9573] = ~(layer1_outputs[1938]) | (layer1_outputs[4127]);
    assign layer2_outputs[9574] = ~(layer1_outputs[6620]);
    assign layer2_outputs[9575] = ~(layer1_outputs[3653]);
    assign layer2_outputs[9576] = ~(layer1_outputs[457]);
    assign layer2_outputs[9577] = layer1_outputs[11282];
    assign layer2_outputs[9578] = (layer1_outputs[12780]) & ~(layer1_outputs[4333]);
    assign layer2_outputs[9579] = ~(layer1_outputs[9013]);
    assign layer2_outputs[9580] = ~((layer1_outputs[3823]) & (layer1_outputs[629]));
    assign layer2_outputs[9581] = (layer1_outputs[11939]) ^ (layer1_outputs[8508]);
    assign layer2_outputs[9582] = (layer1_outputs[10945]) & ~(layer1_outputs[10201]);
    assign layer2_outputs[9583] = ~((layer1_outputs[10779]) & (layer1_outputs[8291]));
    assign layer2_outputs[9584] = (layer1_outputs[330]) & ~(layer1_outputs[11347]);
    assign layer2_outputs[9585] = 1'b1;
    assign layer2_outputs[9586] = layer1_outputs[2428];
    assign layer2_outputs[9587] = ~(layer1_outputs[4462]);
    assign layer2_outputs[9588] = layer1_outputs[9705];
    assign layer2_outputs[9589] = ~(layer1_outputs[4114]);
    assign layer2_outputs[9590] = ~(layer1_outputs[11708]);
    assign layer2_outputs[9591] = ~(layer1_outputs[6914]);
    assign layer2_outputs[9592] = (layer1_outputs[1020]) & ~(layer1_outputs[4611]);
    assign layer2_outputs[9593] = layer1_outputs[2796];
    assign layer2_outputs[9594] = ~(layer1_outputs[5338]) | (layer1_outputs[6787]);
    assign layer2_outputs[9595] = (layer1_outputs[7664]) & (layer1_outputs[10162]);
    assign layer2_outputs[9596] = layer1_outputs[7895];
    assign layer2_outputs[9597] = layer1_outputs[7887];
    assign layer2_outputs[9598] = ~(layer1_outputs[2424]);
    assign layer2_outputs[9599] = 1'b1;
    assign layer2_outputs[9600] = ~((layer1_outputs[6613]) ^ (layer1_outputs[9642]));
    assign layer2_outputs[9601] = ~(layer1_outputs[3632]);
    assign layer2_outputs[9602] = ~(layer1_outputs[4711]);
    assign layer2_outputs[9603] = (layer1_outputs[3872]) | (layer1_outputs[5660]);
    assign layer2_outputs[9604] = ~(layer1_outputs[11439]);
    assign layer2_outputs[9605] = ~(layer1_outputs[10708]);
    assign layer2_outputs[9606] = (layer1_outputs[1791]) ^ (layer1_outputs[10941]);
    assign layer2_outputs[9607] = (layer1_outputs[4338]) ^ (layer1_outputs[7450]);
    assign layer2_outputs[9608] = ~((layer1_outputs[6592]) ^ (layer1_outputs[7849]));
    assign layer2_outputs[9609] = ~(layer1_outputs[5144]) | (layer1_outputs[12422]);
    assign layer2_outputs[9610] = layer1_outputs[6141];
    assign layer2_outputs[9611] = ~(layer1_outputs[125]) | (layer1_outputs[2358]);
    assign layer2_outputs[9612] = ~((layer1_outputs[5462]) ^ (layer1_outputs[11793]));
    assign layer2_outputs[9613] = ~((layer1_outputs[526]) ^ (layer1_outputs[11506]));
    assign layer2_outputs[9614] = ~((layer1_outputs[9467]) & (layer1_outputs[9747]));
    assign layer2_outputs[9615] = layer1_outputs[2415];
    assign layer2_outputs[9616] = ~(layer1_outputs[703]);
    assign layer2_outputs[9617] = layer1_outputs[7311];
    assign layer2_outputs[9618] = layer1_outputs[10049];
    assign layer2_outputs[9619] = ~((layer1_outputs[11127]) | (layer1_outputs[620]));
    assign layer2_outputs[9620] = layer1_outputs[9537];
    assign layer2_outputs[9621] = (layer1_outputs[170]) & ~(layer1_outputs[6581]);
    assign layer2_outputs[9622] = ~(layer1_outputs[7001]);
    assign layer2_outputs[9623] = (layer1_outputs[10447]) & ~(layer1_outputs[3163]);
    assign layer2_outputs[9624] = (layer1_outputs[3551]) & (layer1_outputs[6233]);
    assign layer2_outputs[9625] = (layer1_outputs[11171]) ^ (layer1_outputs[11164]);
    assign layer2_outputs[9626] = layer1_outputs[10116];
    assign layer2_outputs[9627] = ~((layer1_outputs[3641]) ^ (layer1_outputs[10989]));
    assign layer2_outputs[9628] = (layer1_outputs[7618]) ^ (layer1_outputs[2524]);
    assign layer2_outputs[9629] = (layer1_outputs[10335]) & ~(layer1_outputs[12654]);
    assign layer2_outputs[9630] = (layer1_outputs[9244]) | (layer1_outputs[11602]);
    assign layer2_outputs[9631] = layer1_outputs[10591];
    assign layer2_outputs[9632] = (layer1_outputs[3084]) | (layer1_outputs[4581]);
    assign layer2_outputs[9633] = ~((layer1_outputs[5253]) ^ (layer1_outputs[79]));
    assign layer2_outputs[9634] = ~(layer1_outputs[6420]);
    assign layer2_outputs[9635] = (layer1_outputs[11503]) & ~(layer1_outputs[5834]);
    assign layer2_outputs[9636] = ~(layer1_outputs[12228]);
    assign layer2_outputs[9637] = (layer1_outputs[95]) ^ (layer1_outputs[758]);
    assign layer2_outputs[9638] = layer1_outputs[3272];
    assign layer2_outputs[9639] = ~((layer1_outputs[6377]) | (layer1_outputs[10508]));
    assign layer2_outputs[9640] = ~(layer1_outputs[10175]);
    assign layer2_outputs[9641] = (layer1_outputs[5557]) & ~(layer1_outputs[12378]);
    assign layer2_outputs[9642] = (layer1_outputs[6456]) & ~(layer1_outputs[9323]);
    assign layer2_outputs[9643] = (layer1_outputs[9662]) & ~(layer1_outputs[472]);
    assign layer2_outputs[9644] = (layer1_outputs[7763]) ^ (layer1_outputs[6199]);
    assign layer2_outputs[9645] = ~((layer1_outputs[7698]) ^ (layer1_outputs[391]));
    assign layer2_outputs[9646] = ~(layer1_outputs[2443]);
    assign layer2_outputs[9647] = (layer1_outputs[3250]) ^ (layer1_outputs[7634]);
    assign layer2_outputs[9648] = layer1_outputs[4118];
    assign layer2_outputs[9649] = ~(layer1_outputs[6344]);
    assign layer2_outputs[9650] = ~((layer1_outputs[1013]) & (layer1_outputs[5532]));
    assign layer2_outputs[9651] = ~(layer1_outputs[5912]);
    assign layer2_outputs[9652] = ~(layer1_outputs[4435]);
    assign layer2_outputs[9653] = ~((layer1_outputs[5755]) ^ (layer1_outputs[3861]));
    assign layer2_outputs[9654] = ~(layer1_outputs[12067]) | (layer1_outputs[4170]);
    assign layer2_outputs[9655] = ~((layer1_outputs[11310]) ^ (layer1_outputs[11504]));
    assign layer2_outputs[9656] = ~((layer1_outputs[872]) ^ (layer1_outputs[11166]));
    assign layer2_outputs[9657] = ~(layer1_outputs[2955]);
    assign layer2_outputs[9658] = ~(layer1_outputs[407]) | (layer1_outputs[4028]);
    assign layer2_outputs[9659] = layer1_outputs[9421];
    assign layer2_outputs[9660] = ~((layer1_outputs[9923]) ^ (layer1_outputs[8223]));
    assign layer2_outputs[9661] = ~(layer1_outputs[6174]);
    assign layer2_outputs[9662] = layer1_outputs[11770];
    assign layer2_outputs[9663] = ~(layer1_outputs[6805]) | (layer1_outputs[7506]);
    assign layer2_outputs[9664] = ~(layer1_outputs[2871]) | (layer1_outputs[4708]);
    assign layer2_outputs[9665] = ~(layer1_outputs[10031]) | (layer1_outputs[3413]);
    assign layer2_outputs[9666] = (layer1_outputs[11485]) | (layer1_outputs[9552]);
    assign layer2_outputs[9667] = layer1_outputs[7645];
    assign layer2_outputs[9668] = layer1_outputs[1677];
    assign layer2_outputs[9669] = ~((layer1_outputs[12298]) | (layer1_outputs[11148]));
    assign layer2_outputs[9670] = layer1_outputs[5990];
    assign layer2_outputs[9671] = (layer1_outputs[460]) & ~(layer1_outputs[12527]);
    assign layer2_outputs[9672] = 1'b0;
    assign layer2_outputs[9673] = ~(layer1_outputs[7367]);
    assign layer2_outputs[9674] = ~(layer1_outputs[5343]);
    assign layer2_outputs[9675] = layer1_outputs[12607];
    assign layer2_outputs[9676] = layer1_outputs[7218];
    assign layer2_outputs[9677] = layer1_outputs[6800];
    assign layer2_outputs[9678] = layer1_outputs[11729];
    assign layer2_outputs[9679] = ~(layer1_outputs[7865]);
    assign layer2_outputs[9680] = (layer1_outputs[4226]) & (layer1_outputs[5628]);
    assign layer2_outputs[9681] = layer1_outputs[8173];
    assign layer2_outputs[9682] = ~(layer1_outputs[6042]) | (layer1_outputs[7321]);
    assign layer2_outputs[9683] = layer1_outputs[11803];
    assign layer2_outputs[9684] = layer1_outputs[4049];
    assign layer2_outputs[9685] = (layer1_outputs[4190]) | (layer1_outputs[1518]);
    assign layer2_outputs[9686] = ~(layer1_outputs[2214]) | (layer1_outputs[251]);
    assign layer2_outputs[9687] = (layer1_outputs[2291]) | (layer1_outputs[9506]);
    assign layer2_outputs[9688] = ~(layer1_outputs[4179]) | (layer1_outputs[8493]);
    assign layer2_outputs[9689] = layer1_outputs[8617];
    assign layer2_outputs[9690] = ~(layer1_outputs[5454]) | (layer1_outputs[12674]);
    assign layer2_outputs[9691] = (layer1_outputs[1600]) & (layer1_outputs[5139]);
    assign layer2_outputs[9692] = ~(layer1_outputs[3662]);
    assign layer2_outputs[9693] = layer1_outputs[40];
    assign layer2_outputs[9694] = layer1_outputs[6410];
    assign layer2_outputs[9695] = ~((layer1_outputs[12150]) | (layer1_outputs[8240]));
    assign layer2_outputs[9696] = layer1_outputs[9061];
    assign layer2_outputs[9697] = ~(layer1_outputs[11113]);
    assign layer2_outputs[9698] = ~((layer1_outputs[7600]) & (layer1_outputs[2268]));
    assign layer2_outputs[9699] = layer1_outputs[8631];
    assign layer2_outputs[9700] = ~(layer1_outputs[7552]) | (layer1_outputs[11307]);
    assign layer2_outputs[9701] = ~(layer1_outputs[10172]);
    assign layer2_outputs[9702] = layer1_outputs[5653];
    assign layer2_outputs[9703] = ~(layer1_outputs[4872]) | (layer1_outputs[11554]);
    assign layer2_outputs[9704] = ~(layer1_outputs[8739]);
    assign layer2_outputs[9705] = ~(layer1_outputs[11282]) | (layer1_outputs[4559]);
    assign layer2_outputs[9706] = (layer1_outputs[7378]) & (layer1_outputs[9291]);
    assign layer2_outputs[9707] = ~(layer1_outputs[10232]);
    assign layer2_outputs[9708] = (layer1_outputs[9846]) & ~(layer1_outputs[1629]);
    assign layer2_outputs[9709] = (layer1_outputs[2727]) & ~(layer1_outputs[5722]);
    assign layer2_outputs[9710] = ~(layer1_outputs[977]);
    assign layer2_outputs[9711] = layer1_outputs[8119];
    assign layer2_outputs[9712] = ~(layer1_outputs[5910]);
    assign layer2_outputs[9713] = (layer1_outputs[4050]) & (layer1_outputs[5766]);
    assign layer2_outputs[9714] = ~((layer1_outputs[1936]) | (layer1_outputs[3991]));
    assign layer2_outputs[9715] = ~(layer1_outputs[11252]);
    assign layer2_outputs[9716] = layer1_outputs[738];
    assign layer2_outputs[9717] = (layer1_outputs[713]) | (layer1_outputs[9453]);
    assign layer2_outputs[9718] = ~(layer1_outputs[4492]) | (layer1_outputs[6074]);
    assign layer2_outputs[9719] = layer1_outputs[1848];
    assign layer2_outputs[9720] = (layer1_outputs[9989]) & ~(layer1_outputs[8024]);
    assign layer2_outputs[9721] = ~((layer1_outputs[11274]) ^ (layer1_outputs[5928]));
    assign layer2_outputs[9722] = ~((layer1_outputs[3220]) ^ (layer1_outputs[8459]));
    assign layer2_outputs[9723] = ~(layer1_outputs[5650]);
    assign layer2_outputs[9724] = (layer1_outputs[8486]) ^ (layer1_outputs[12176]);
    assign layer2_outputs[9725] = ~(layer1_outputs[4571]);
    assign layer2_outputs[9726] = (layer1_outputs[7190]) | (layer1_outputs[1537]);
    assign layer2_outputs[9727] = ~((layer1_outputs[12581]) ^ (layer1_outputs[9555]));
    assign layer2_outputs[9728] = layer1_outputs[6399];
    assign layer2_outputs[9729] = (layer1_outputs[1542]) & ~(layer1_outputs[7667]);
    assign layer2_outputs[9730] = 1'b0;
    assign layer2_outputs[9731] = (layer1_outputs[3916]) ^ (layer1_outputs[1411]);
    assign layer2_outputs[9732] = layer1_outputs[8708];
    assign layer2_outputs[9733] = ~(layer1_outputs[8048]);
    assign layer2_outputs[9734] = ~(layer1_outputs[2146]);
    assign layer2_outputs[9735] = ~(layer1_outputs[8372]);
    assign layer2_outputs[9736] = ~(layer1_outputs[1413]);
    assign layer2_outputs[9737] = layer1_outputs[2260];
    assign layer2_outputs[9738] = ~(layer1_outputs[8738]);
    assign layer2_outputs[9739] = ~(layer1_outputs[514]);
    assign layer2_outputs[9740] = ~(layer1_outputs[5940]);
    assign layer2_outputs[9741] = ~(layer1_outputs[11857]);
    assign layer2_outputs[9742] = ~((layer1_outputs[1544]) & (layer1_outputs[5709]));
    assign layer2_outputs[9743] = ~((layer1_outputs[12747]) | (layer1_outputs[4142]));
    assign layer2_outputs[9744] = ~(layer1_outputs[7827]);
    assign layer2_outputs[9745] = ~((layer1_outputs[3857]) ^ (layer1_outputs[3490]));
    assign layer2_outputs[9746] = ~((layer1_outputs[3175]) ^ (layer1_outputs[10478]));
    assign layer2_outputs[9747] = ~(layer1_outputs[12142]);
    assign layer2_outputs[9748] = ~((layer1_outputs[625]) ^ (layer1_outputs[2818]));
    assign layer2_outputs[9749] = ~(layer1_outputs[3286]);
    assign layer2_outputs[9750] = ~(layer1_outputs[3621]);
    assign layer2_outputs[9751] = layer1_outputs[6923];
    assign layer2_outputs[9752] = layer1_outputs[8063];
    assign layer2_outputs[9753] = ~(layer1_outputs[8339]);
    assign layer2_outputs[9754] = ~((layer1_outputs[11224]) | (layer1_outputs[3550]));
    assign layer2_outputs[9755] = (layer1_outputs[1479]) ^ (layer1_outputs[1664]);
    assign layer2_outputs[9756] = ~(layer1_outputs[12242]);
    assign layer2_outputs[9757] = ~(layer1_outputs[4288]);
    assign layer2_outputs[9758] = ~(layer1_outputs[3185]) | (layer1_outputs[2702]);
    assign layer2_outputs[9759] = layer1_outputs[6036];
    assign layer2_outputs[9760] = ~(layer1_outputs[7365]);
    assign layer2_outputs[9761] = layer1_outputs[10809];
    assign layer2_outputs[9762] = layer1_outputs[212];
    assign layer2_outputs[9763] = (layer1_outputs[12188]) & (layer1_outputs[6361]);
    assign layer2_outputs[9764] = layer1_outputs[761];
    assign layer2_outputs[9765] = ~(layer1_outputs[3790]);
    assign layer2_outputs[9766] = layer1_outputs[1994];
    assign layer2_outputs[9767] = layer1_outputs[4195];
    assign layer2_outputs[9768] = (layer1_outputs[12546]) ^ (layer1_outputs[2655]);
    assign layer2_outputs[9769] = ~(layer1_outputs[10229]);
    assign layer2_outputs[9770] = layer1_outputs[4599];
    assign layer2_outputs[9771] = (layer1_outputs[5633]) & (layer1_outputs[631]);
    assign layer2_outputs[9772] = ~(layer1_outputs[6532]);
    assign layer2_outputs[9773] = ~(layer1_outputs[10553]);
    assign layer2_outputs[9774] = layer1_outputs[8526];
    assign layer2_outputs[9775] = ~(layer1_outputs[5737]);
    assign layer2_outputs[9776] = ~((layer1_outputs[3376]) | (layer1_outputs[9207]));
    assign layer2_outputs[9777] = ~((layer1_outputs[4452]) ^ (layer1_outputs[12726]));
    assign layer2_outputs[9778] = layer1_outputs[8674];
    assign layer2_outputs[9779] = layer1_outputs[3800];
    assign layer2_outputs[9780] = ~(layer1_outputs[6636]) | (layer1_outputs[362]);
    assign layer2_outputs[9781] = ~((layer1_outputs[8762]) ^ (layer1_outputs[520]));
    assign layer2_outputs[9782] = layer1_outputs[1416];
    assign layer2_outputs[9783] = (layer1_outputs[8586]) ^ (layer1_outputs[10739]);
    assign layer2_outputs[9784] = (layer1_outputs[4286]) & ~(layer1_outputs[11089]);
    assign layer2_outputs[9785] = (layer1_outputs[9309]) & ~(layer1_outputs[11937]);
    assign layer2_outputs[9786] = ~(layer1_outputs[4668]);
    assign layer2_outputs[9787] = layer1_outputs[9308];
    assign layer2_outputs[9788] = (layer1_outputs[1804]) & ~(layer1_outputs[6089]);
    assign layer2_outputs[9789] = (layer1_outputs[2118]) & ~(layer1_outputs[11045]);
    assign layer2_outputs[9790] = (layer1_outputs[3909]) & (layer1_outputs[5401]);
    assign layer2_outputs[9791] = (layer1_outputs[9031]) & ~(layer1_outputs[8025]);
    assign layer2_outputs[9792] = (layer1_outputs[4038]) ^ (layer1_outputs[6223]);
    assign layer2_outputs[9793] = (layer1_outputs[4341]) & (layer1_outputs[10595]);
    assign layer2_outputs[9794] = (layer1_outputs[8214]) & ~(layer1_outputs[9264]);
    assign layer2_outputs[9795] = ~((layer1_outputs[733]) | (layer1_outputs[12484]));
    assign layer2_outputs[9796] = ~(layer1_outputs[3464]) | (layer1_outputs[6883]);
    assign layer2_outputs[9797] = (layer1_outputs[7630]) & ~(layer1_outputs[10537]);
    assign layer2_outputs[9798] = ~(layer1_outputs[3690]);
    assign layer2_outputs[9799] = (layer1_outputs[8404]) & ~(layer1_outputs[1123]);
    assign layer2_outputs[9800] = (layer1_outputs[8831]) & (layer1_outputs[5935]);
    assign layer2_outputs[9801] = ~((layer1_outputs[5529]) ^ (layer1_outputs[2674]));
    assign layer2_outputs[9802] = ~(layer1_outputs[11197]);
    assign layer2_outputs[9803] = ~(layer1_outputs[7436]);
    assign layer2_outputs[9804] = ~(layer1_outputs[2362]) | (layer1_outputs[569]);
    assign layer2_outputs[9805] = ~(layer1_outputs[11901]) | (layer1_outputs[12446]);
    assign layer2_outputs[9806] = layer1_outputs[2009];
    assign layer2_outputs[9807] = ~(layer1_outputs[11715]);
    assign layer2_outputs[9808] = ~(layer1_outputs[6187]) | (layer1_outputs[3980]);
    assign layer2_outputs[9809] = (layer1_outputs[5149]) ^ (layer1_outputs[4752]);
    assign layer2_outputs[9810] = ~((layer1_outputs[2071]) | (layer1_outputs[10890]));
    assign layer2_outputs[9811] = (layer1_outputs[2053]) & ~(layer1_outputs[4437]);
    assign layer2_outputs[9812] = ~(layer1_outputs[640]);
    assign layer2_outputs[9813] = ~((layer1_outputs[7580]) | (layer1_outputs[5631]));
    assign layer2_outputs[9814] = layer1_outputs[8284];
    assign layer2_outputs[9815] = ~(layer1_outputs[12008]);
    assign layer2_outputs[9816] = (layer1_outputs[8406]) & ~(layer1_outputs[8512]);
    assign layer2_outputs[9817] = (layer1_outputs[2804]) & ~(layer1_outputs[8199]);
    assign layer2_outputs[9818] = (layer1_outputs[8698]) & (layer1_outputs[7006]);
    assign layer2_outputs[9819] = layer1_outputs[4460];
    assign layer2_outputs[9820] = ~(layer1_outputs[5217]);
    assign layer2_outputs[9821] = ~((layer1_outputs[11130]) ^ (layer1_outputs[5977]));
    assign layer2_outputs[9822] = ~((layer1_outputs[6008]) | (layer1_outputs[7465]));
    assign layer2_outputs[9823] = (layer1_outputs[558]) | (layer1_outputs[1146]);
    assign layer2_outputs[9824] = ~(layer1_outputs[1828]) | (layer1_outputs[5671]);
    assign layer2_outputs[9825] = (layer1_outputs[11244]) & ~(layer1_outputs[5448]);
    assign layer2_outputs[9826] = ~(layer1_outputs[11386]);
    assign layer2_outputs[9827] = ~((layer1_outputs[7336]) ^ (layer1_outputs[6466]));
    assign layer2_outputs[9828] = ~(layer1_outputs[8169]) | (layer1_outputs[5736]);
    assign layer2_outputs[9829] = layer1_outputs[6186];
    assign layer2_outputs[9830] = layer1_outputs[6426];
    assign layer2_outputs[9831] = ~(layer1_outputs[4239]) | (layer1_outputs[11621]);
    assign layer2_outputs[9832] = layer1_outputs[12397];
    assign layer2_outputs[9833] = (layer1_outputs[10642]) & ~(layer1_outputs[3739]);
    assign layer2_outputs[9834] = ~((layer1_outputs[8176]) | (layer1_outputs[5619]));
    assign layer2_outputs[9835] = (layer1_outputs[9032]) & (layer1_outputs[12745]);
    assign layer2_outputs[9836] = 1'b0;
    assign layer2_outputs[9837] = ~(layer1_outputs[12199]);
    assign layer2_outputs[9838] = ~(layer1_outputs[2100]);
    assign layer2_outputs[9839] = layer1_outputs[7120];
    assign layer2_outputs[9840] = ~(layer1_outputs[8672]) | (layer1_outputs[670]);
    assign layer2_outputs[9841] = ~(layer1_outputs[1957]);
    assign layer2_outputs[9842] = (layer1_outputs[1384]) & (layer1_outputs[6362]);
    assign layer2_outputs[9843] = (layer1_outputs[9124]) ^ (layer1_outputs[3169]);
    assign layer2_outputs[9844] = (layer1_outputs[10835]) ^ (layer1_outputs[2366]);
    assign layer2_outputs[9845] = layer1_outputs[565];
    assign layer2_outputs[9846] = ~(layer1_outputs[10106]);
    assign layer2_outputs[9847] = (layer1_outputs[10677]) ^ (layer1_outputs[5389]);
    assign layer2_outputs[9848] = 1'b1;
    assign layer2_outputs[9849] = ~(layer1_outputs[7204]) | (layer1_outputs[5387]);
    assign layer2_outputs[9850] = layer1_outputs[6157];
    assign layer2_outputs[9851] = (layer1_outputs[10272]) & (layer1_outputs[3771]);
    assign layer2_outputs[9852] = ~(layer1_outputs[3822]);
    assign layer2_outputs[9853] = (layer1_outputs[10698]) ^ (layer1_outputs[87]);
    assign layer2_outputs[9854] = ~(layer1_outputs[1866]) | (layer1_outputs[3977]);
    assign layer2_outputs[9855] = (layer1_outputs[3545]) & ~(layer1_outputs[5939]);
    assign layer2_outputs[9856] = ~((layer1_outputs[6663]) ^ (layer1_outputs[2299]));
    assign layer2_outputs[9857] = (layer1_outputs[8168]) ^ (layer1_outputs[12186]);
    assign layer2_outputs[9858] = ~(layer1_outputs[7300]);
    assign layer2_outputs[9859] = (layer1_outputs[11175]) ^ (layer1_outputs[10488]);
    assign layer2_outputs[9860] = (layer1_outputs[5920]) & ~(layer1_outputs[5800]);
    assign layer2_outputs[9861] = (layer1_outputs[5607]) ^ (layer1_outputs[4568]);
    assign layer2_outputs[9862] = ~((layer1_outputs[89]) ^ (layer1_outputs[3590]));
    assign layer2_outputs[9863] = layer1_outputs[11870];
    assign layer2_outputs[9864] = ~(layer1_outputs[11570]) | (layer1_outputs[5401]);
    assign layer2_outputs[9865] = ~(layer1_outputs[12712]);
    assign layer2_outputs[9866] = ~((layer1_outputs[5281]) ^ (layer1_outputs[11247]));
    assign layer2_outputs[9867] = ~(layer1_outputs[575]);
    assign layer2_outputs[9868] = layer1_outputs[3175];
    assign layer2_outputs[9869] = layer1_outputs[8077];
    assign layer2_outputs[9870] = (layer1_outputs[9197]) & (layer1_outputs[12597]);
    assign layer2_outputs[9871] = (layer1_outputs[10699]) & ~(layer1_outputs[5323]);
    assign layer2_outputs[9872] = (layer1_outputs[12185]) | (layer1_outputs[143]);
    assign layer2_outputs[9873] = ~(layer1_outputs[6709]);
    assign layer2_outputs[9874] = ~(layer1_outputs[793]);
    assign layer2_outputs[9875] = ~((layer1_outputs[9475]) | (layer1_outputs[5996]));
    assign layer2_outputs[9876] = ~(layer1_outputs[8841]) | (layer1_outputs[58]);
    assign layer2_outputs[9877] = ~(layer1_outputs[132]);
    assign layer2_outputs[9878] = ~((layer1_outputs[10945]) & (layer1_outputs[1980]));
    assign layer2_outputs[9879] = ~((layer1_outputs[7612]) ^ (layer1_outputs[1474]));
    assign layer2_outputs[9880] = (layer1_outputs[4530]) & (layer1_outputs[9632]);
    assign layer2_outputs[9881] = (layer1_outputs[42]) & ~(layer1_outputs[7012]);
    assign layer2_outputs[9882] = ~(layer1_outputs[5423]);
    assign layer2_outputs[9883] = ~((layer1_outputs[7009]) ^ (layer1_outputs[10722]));
    assign layer2_outputs[9884] = ~(layer1_outputs[3089]);
    assign layer2_outputs[9885] = ~((layer1_outputs[8924]) & (layer1_outputs[78]));
    assign layer2_outputs[9886] = (layer1_outputs[1402]) | (layer1_outputs[4578]);
    assign layer2_outputs[9887] = ~(layer1_outputs[3546]);
    assign layer2_outputs[9888] = ~(layer1_outputs[6616]);
    assign layer2_outputs[9889] = (layer1_outputs[1337]) & ~(layer1_outputs[7413]);
    assign layer2_outputs[9890] = ~(layer1_outputs[3913]) | (layer1_outputs[11339]);
    assign layer2_outputs[9891] = ~(layer1_outputs[5600]);
    assign layer2_outputs[9892] = ~(layer1_outputs[12383]);
    assign layer2_outputs[9893] = layer1_outputs[8328];
    assign layer2_outputs[9894] = ~((layer1_outputs[88]) | (layer1_outputs[252]));
    assign layer2_outputs[9895] = ~(layer1_outputs[5434]);
    assign layer2_outputs[9896] = (layer1_outputs[9266]) | (layer1_outputs[11030]);
    assign layer2_outputs[9897] = ~(layer1_outputs[3874]);
    assign layer2_outputs[9898] = (layer1_outputs[10354]) ^ (layer1_outputs[2666]);
    assign layer2_outputs[9899] = ~((layer1_outputs[10919]) ^ (layer1_outputs[8418]));
    assign layer2_outputs[9900] = ~(layer1_outputs[8066]);
    assign layer2_outputs[9901] = ~(layer1_outputs[2598]);
    assign layer2_outputs[9902] = ~(layer1_outputs[4356]);
    assign layer2_outputs[9903] = ~(layer1_outputs[446]);
    assign layer2_outputs[9904] = layer1_outputs[8138];
    assign layer2_outputs[9905] = ~(layer1_outputs[5924]);
    assign layer2_outputs[9906] = (layer1_outputs[7833]) & ~(layer1_outputs[1612]);
    assign layer2_outputs[9907] = (layer1_outputs[3949]) & (layer1_outputs[7837]);
    assign layer2_outputs[9908] = (layer1_outputs[12587]) & ~(layer1_outputs[8761]);
    assign layer2_outputs[9909] = layer1_outputs[4201];
    assign layer2_outputs[9910] = layer1_outputs[1579];
    assign layer2_outputs[9911] = layer1_outputs[11857];
    assign layer2_outputs[9912] = ~(layer1_outputs[10332]);
    assign layer2_outputs[9913] = layer1_outputs[5896];
    assign layer2_outputs[9914] = ~(layer1_outputs[10482]);
    assign layer2_outputs[9915] = (layer1_outputs[6737]) & ~(layer1_outputs[7351]);
    assign layer2_outputs[9916] = (layer1_outputs[5783]) | (layer1_outputs[7337]);
    assign layer2_outputs[9917] = ~(layer1_outputs[1003]);
    assign layer2_outputs[9918] = ~(layer1_outputs[12055]) | (layer1_outputs[6351]);
    assign layer2_outputs[9919] = (layer1_outputs[1234]) | (layer1_outputs[6208]);
    assign layer2_outputs[9920] = ~(layer1_outputs[3415]);
    assign layer2_outputs[9921] = 1'b1;
    assign layer2_outputs[9922] = ~(layer1_outputs[3805]) | (layer1_outputs[295]);
    assign layer2_outputs[9923] = ~((layer1_outputs[11962]) & (layer1_outputs[2980]));
    assign layer2_outputs[9924] = ~(layer1_outputs[8129]) | (layer1_outputs[6987]);
    assign layer2_outputs[9925] = ~((layer1_outputs[12167]) | (layer1_outputs[11279]));
    assign layer2_outputs[9926] = (layer1_outputs[9214]) & (layer1_outputs[12323]);
    assign layer2_outputs[9927] = ~(layer1_outputs[5465]) | (layer1_outputs[10813]);
    assign layer2_outputs[9928] = layer1_outputs[5667];
    assign layer2_outputs[9929] = (layer1_outputs[9570]) ^ (layer1_outputs[9023]);
    assign layer2_outputs[9930] = layer1_outputs[11259];
    assign layer2_outputs[9931] = ~(layer1_outputs[8816]);
    assign layer2_outputs[9932] = ~(layer1_outputs[2830]);
    assign layer2_outputs[9933] = (layer1_outputs[12624]) & ~(layer1_outputs[7666]);
    assign layer2_outputs[9934] = ~(layer1_outputs[2948]);
    assign layer2_outputs[9935] = (layer1_outputs[4351]) ^ (layer1_outputs[1478]);
    assign layer2_outputs[9936] = (layer1_outputs[5397]) & ~(layer1_outputs[10496]);
    assign layer2_outputs[9937] = ~(layer1_outputs[6892]);
    assign layer2_outputs[9938] = layer1_outputs[10014];
    assign layer2_outputs[9939] = (layer1_outputs[3152]) ^ (layer1_outputs[12509]);
    assign layer2_outputs[9940] = (layer1_outputs[3189]) & ~(layer1_outputs[7635]);
    assign layer2_outputs[9941] = layer1_outputs[8929];
    assign layer2_outputs[9942] = ~(layer1_outputs[4801]);
    assign layer2_outputs[9943] = (layer1_outputs[1787]) | (layer1_outputs[10465]);
    assign layer2_outputs[9944] = ~(layer1_outputs[10879]);
    assign layer2_outputs[9945] = (layer1_outputs[5668]) & (layer1_outputs[6722]);
    assign layer2_outputs[9946] = (layer1_outputs[10099]) ^ (layer1_outputs[12550]);
    assign layer2_outputs[9947] = layer1_outputs[4503];
    assign layer2_outputs[9948] = (layer1_outputs[278]) & (layer1_outputs[3358]);
    assign layer2_outputs[9949] = ~(layer1_outputs[3817]);
    assign layer2_outputs[9950] = (layer1_outputs[12233]) & (layer1_outputs[11488]);
    assign layer2_outputs[9951] = layer1_outputs[1039];
    assign layer2_outputs[9952] = (layer1_outputs[12286]) & (layer1_outputs[2982]);
    assign layer2_outputs[9953] = ~(layer1_outputs[7817]) | (layer1_outputs[7385]);
    assign layer2_outputs[9954] = ~((layer1_outputs[2464]) ^ (layer1_outputs[3486]));
    assign layer2_outputs[9955] = ~((layer1_outputs[6566]) & (layer1_outputs[140]));
    assign layer2_outputs[9956] = ~(layer1_outputs[5538]);
    assign layer2_outputs[9957] = ~(layer1_outputs[9041]);
    assign layer2_outputs[9958] = (layer1_outputs[896]) ^ (layer1_outputs[860]);
    assign layer2_outputs[9959] = ~((layer1_outputs[5752]) ^ (layer1_outputs[1742]));
    assign layer2_outputs[9960] = layer1_outputs[9986];
    assign layer2_outputs[9961] = ~(layer1_outputs[2376]);
    assign layer2_outputs[9962] = (layer1_outputs[6584]) & ~(layer1_outputs[3164]);
    assign layer2_outputs[9963] = ~(layer1_outputs[7923]);
    assign layer2_outputs[9964] = (layer1_outputs[4106]) & ~(layer1_outputs[2837]);
    assign layer2_outputs[9965] = (layer1_outputs[9086]) ^ (layer1_outputs[7739]);
    assign layer2_outputs[9966] = layer1_outputs[5437];
    assign layer2_outputs[9967] = ~(layer1_outputs[1219]) | (layer1_outputs[4464]);
    assign layer2_outputs[9968] = layer1_outputs[2125];
    assign layer2_outputs[9969] = layer1_outputs[10861];
    assign layer2_outputs[9970] = layer1_outputs[234];
    assign layer2_outputs[9971] = (layer1_outputs[3640]) & ~(layer1_outputs[11068]);
    assign layer2_outputs[9972] = ~((layer1_outputs[3039]) ^ (layer1_outputs[1186]));
    assign layer2_outputs[9973] = layer1_outputs[8782];
    assign layer2_outputs[9974] = layer1_outputs[3270];
    assign layer2_outputs[9975] = layer1_outputs[206];
    assign layer2_outputs[9976] = ~((layer1_outputs[7697]) | (layer1_outputs[11963]));
    assign layer2_outputs[9977] = ~(layer1_outputs[5578]) | (layer1_outputs[6353]);
    assign layer2_outputs[9978] = layer1_outputs[3703];
    assign layer2_outputs[9979] = ~((layer1_outputs[11973]) ^ (layer1_outputs[4497]));
    assign layer2_outputs[9980] = ~(layer1_outputs[10860]);
    assign layer2_outputs[9981] = (layer1_outputs[12115]) | (layer1_outputs[5037]);
    assign layer2_outputs[9982] = (layer1_outputs[2666]) ^ (layer1_outputs[7871]);
    assign layer2_outputs[9983] = ~(layer1_outputs[432]) | (layer1_outputs[2163]);
    assign layer2_outputs[9984] = ~((layer1_outputs[11285]) & (layer1_outputs[888]));
    assign layer2_outputs[9985] = (layer1_outputs[8954]) & (layer1_outputs[6885]);
    assign layer2_outputs[9986] = layer1_outputs[11481];
    assign layer2_outputs[9987] = layer1_outputs[340];
    assign layer2_outputs[9988] = layer1_outputs[10755];
    assign layer2_outputs[9989] = ~((layer1_outputs[2453]) ^ (layer1_outputs[6402]));
    assign layer2_outputs[9990] = ~(layer1_outputs[7184]);
    assign layer2_outputs[9991] = (layer1_outputs[3035]) & ~(layer1_outputs[1355]);
    assign layer2_outputs[9992] = layer1_outputs[6934];
    assign layer2_outputs[9993] = ~(layer1_outputs[676]) | (layer1_outputs[11253]);
    assign layer2_outputs[9994] = ~(layer1_outputs[6931]);
    assign layer2_outputs[9995] = layer1_outputs[1539];
    assign layer2_outputs[9996] = layer1_outputs[4192];
    assign layer2_outputs[9997] = ~((layer1_outputs[5410]) ^ (layer1_outputs[7804]));
    assign layer2_outputs[9998] = ~((layer1_outputs[468]) & (layer1_outputs[1423]));
    assign layer2_outputs[9999] = (layer1_outputs[8261]) & ~(layer1_outputs[7402]);
    assign layer2_outputs[10000] = ~(layer1_outputs[8959]);
    assign layer2_outputs[10001] = (layer1_outputs[7506]) & (layer1_outputs[1397]);
    assign layer2_outputs[10002] = ~(layer1_outputs[9786]);
    assign layer2_outputs[10003] = (layer1_outputs[1005]) & ~(layer1_outputs[11130]);
    assign layer2_outputs[10004] = layer1_outputs[9969];
    assign layer2_outputs[10005] = layer1_outputs[3721];
    assign layer2_outputs[10006] = ~(layer1_outputs[2215]) | (layer1_outputs[7199]);
    assign layer2_outputs[10007] = ~(layer1_outputs[10387]) | (layer1_outputs[6293]);
    assign layer2_outputs[10008] = (layer1_outputs[9075]) | (layer1_outputs[173]);
    assign layer2_outputs[10009] = (layer1_outputs[341]) & (layer1_outputs[2404]);
    assign layer2_outputs[10010] = ~(layer1_outputs[12679]);
    assign layer2_outputs[10011] = layer1_outputs[7828];
    assign layer2_outputs[10012] = (layer1_outputs[1053]) & (layer1_outputs[1852]);
    assign layer2_outputs[10013] = (layer1_outputs[3147]) & ~(layer1_outputs[4850]);
    assign layer2_outputs[10014] = ~(layer1_outputs[1093]);
    assign layer2_outputs[10015] = layer1_outputs[10573];
    assign layer2_outputs[10016] = layer1_outputs[3418];
    assign layer2_outputs[10017] = (layer1_outputs[9220]) & ~(layer1_outputs[5216]);
    assign layer2_outputs[10018] = ~(layer1_outputs[6917]);
    assign layer2_outputs[10019] = (layer1_outputs[5986]) & ~(layer1_outputs[4701]);
    assign layer2_outputs[10020] = (layer1_outputs[4366]) & ~(layer1_outputs[4018]);
    assign layer2_outputs[10021] = (layer1_outputs[7320]) & ~(layer1_outputs[1863]);
    assign layer2_outputs[10022] = layer1_outputs[1476];
    assign layer2_outputs[10023] = ~((layer1_outputs[3354]) ^ (layer1_outputs[2366]));
    assign layer2_outputs[10024] = layer1_outputs[5616];
    assign layer2_outputs[10025] = ~(layer1_outputs[8768]);
    assign layer2_outputs[10026] = (layer1_outputs[1892]) | (layer1_outputs[198]);
    assign layer2_outputs[10027] = ~((layer1_outputs[4383]) | (layer1_outputs[10875]));
    assign layer2_outputs[10028] = layer1_outputs[6627];
    assign layer2_outputs[10029] = ~(layer1_outputs[1975]) | (layer1_outputs[9333]);
    assign layer2_outputs[10030] = ~((layer1_outputs[7144]) ^ (layer1_outputs[1635]));
    assign layer2_outputs[10031] = (layer1_outputs[513]) ^ (layer1_outputs[6142]);
    assign layer2_outputs[10032] = (layer1_outputs[9241]) | (layer1_outputs[3417]);
    assign layer2_outputs[10033] = layer1_outputs[3787];
    assign layer2_outputs[10034] = ~((layer1_outputs[5270]) ^ (layer1_outputs[2375]));
    assign layer2_outputs[10035] = ~(layer1_outputs[4966]);
    assign layer2_outputs[10036] = ~((layer1_outputs[1420]) & (layer1_outputs[8355]));
    assign layer2_outputs[10037] = ~(layer1_outputs[449]) | (layer1_outputs[3126]);
    assign layer2_outputs[10038] = layer1_outputs[6934];
    assign layer2_outputs[10039] = ~(layer1_outputs[6677]) | (layer1_outputs[5526]);
    assign layer2_outputs[10040] = (layer1_outputs[2421]) & ~(layer1_outputs[10943]);
    assign layer2_outputs[10041] = (layer1_outputs[8557]) | (layer1_outputs[12123]);
    assign layer2_outputs[10042] = layer1_outputs[10603];
    assign layer2_outputs[10043] = ~(layer1_outputs[8318]);
    assign layer2_outputs[10044] = ~(layer1_outputs[1260]);
    assign layer2_outputs[10045] = ~(layer1_outputs[3650]) | (layer1_outputs[11929]);
    assign layer2_outputs[10046] = (layer1_outputs[6343]) | (layer1_outputs[4027]);
    assign layer2_outputs[10047] = ~((layer1_outputs[1718]) | (layer1_outputs[2215]));
    assign layer2_outputs[10048] = ~((layer1_outputs[4965]) & (layer1_outputs[2392]));
    assign layer2_outputs[10049] = ~(layer1_outputs[2970]);
    assign layer2_outputs[10050] = layer1_outputs[1694];
    assign layer2_outputs[10051] = ~(layer1_outputs[12535]);
    assign layer2_outputs[10052] = ~(layer1_outputs[1692]);
    assign layer2_outputs[10053] = ~(layer1_outputs[3794]);
    assign layer2_outputs[10054] = layer1_outputs[9994];
    assign layer2_outputs[10055] = (layer1_outputs[12212]) & ~(layer1_outputs[8677]);
    assign layer2_outputs[10056] = ~(layer1_outputs[2769]);
    assign layer2_outputs[10057] = layer1_outputs[5481];
    assign layer2_outputs[10058] = (layer1_outputs[7010]) & (layer1_outputs[3333]);
    assign layer2_outputs[10059] = (layer1_outputs[11054]) ^ (layer1_outputs[4577]);
    assign layer2_outputs[10060] = layer1_outputs[8264];
    assign layer2_outputs[10061] = ~(layer1_outputs[12178]);
    assign layer2_outputs[10062] = ~(layer1_outputs[7225]);
    assign layer2_outputs[10063] = layer1_outputs[10133];
    assign layer2_outputs[10064] = (layer1_outputs[5455]) ^ (layer1_outputs[10615]);
    assign layer2_outputs[10065] = layer1_outputs[11555];
    assign layer2_outputs[10066] = ~(layer1_outputs[152]);
    assign layer2_outputs[10067] = (layer1_outputs[2239]) ^ (layer1_outputs[2232]);
    assign layer2_outputs[10068] = (layer1_outputs[7876]) & ~(layer1_outputs[90]);
    assign layer2_outputs[10069] = (layer1_outputs[6671]) & ~(layer1_outputs[339]);
    assign layer2_outputs[10070] = ~(layer1_outputs[10458]);
    assign layer2_outputs[10071] = layer1_outputs[5609];
    assign layer2_outputs[10072] = (layer1_outputs[6242]) & ~(layer1_outputs[3576]);
    assign layer2_outputs[10073] = ~((layer1_outputs[3902]) | (layer1_outputs[1460]));
    assign layer2_outputs[10074] = layer1_outputs[7631];
    assign layer2_outputs[10075] = ~(layer1_outputs[6463]);
    assign layer2_outputs[10076] = (layer1_outputs[9731]) | (layer1_outputs[11471]);
    assign layer2_outputs[10077] = (layer1_outputs[3124]) & ~(layer1_outputs[12141]);
    assign layer2_outputs[10078] = ~((layer1_outputs[367]) | (layer1_outputs[5439]));
    assign layer2_outputs[10079] = ~(layer1_outputs[9348]);
    assign layer2_outputs[10080] = layer1_outputs[8777];
    assign layer2_outputs[10081] = layer1_outputs[12146];
    assign layer2_outputs[10082] = (layer1_outputs[592]) & ~(layer1_outputs[3125]);
    assign layer2_outputs[10083] = (layer1_outputs[790]) ^ (layer1_outputs[4065]);
    assign layer2_outputs[10084] = (layer1_outputs[1084]) & ~(layer1_outputs[4509]);
    assign layer2_outputs[10085] = (layer1_outputs[5485]) & ~(layer1_outputs[8042]);
    assign layer2_outputs[10086] = ~(layer1_outputs[4300]);
    assign layer2_outputs[10087] = ~((layer1_outputs[101]) ^ (layer1_outputs[8584]));
    assign layer2_outputs[10088] = (layer1_outputs[4444]) | (layer1_outputs[9694]);
    assign layer2_outputs[10089] = ~((layer1_outputs[3920]) ^ (layer1_outputs[9529]));
    assign layer2_outputs[10090] = (layer1_outputs[4099]) ^ (layer1_outputs[10347]);
    assign layer2_outputs[10091] = ~((layer1_outputs[11891]) & (layer1_outputs[5755]));
    assign layer2_outputs[10092] = ~(layer1_outputs[2750]);
    assign layer2_outputs[10093] = ~(layer1_outputs[1597]);
    assign layer2_outputs[10094] = ~(layer1_outputs[1895]) | (layer1_outputs[10775]);
    assign layer2_outputs[10095] = ~(layer1_outputs[235]);
    assign layer2_outputs[10096] = ~((layer1_outputs[5729]) & (layer1_outputs[3690]));
    assign layer2_outputs[10097] = (layer1_outputs[8506]) ^ (layer1_outputs[11986]);
    assign layer2_outputs[10098] = layer1_outputs[9404];
    assign layer2_outputs[10099] = ~(layer1_outputs[1997]) | (layer1_outputs[11202]);
    assign layer2_outputs[10100] = ~(layer1_outputs[8855]) | (layer1_outputs[10160]);
    assign layer2_outputs[10101] = layer1_outputs[2757];
    assign layer2_outputs[10102] = layer1_outputs[10668];
    assign layer2_outputs[10103] = layer1_outputs[11998];
    assign layer2_outputs[10104] = (layer1_outputs[7363]) & (layer1_outputs[4988]);
    assign layer2_outputs[10105] = 1'b1;
    assign layer2_outputs[10106] = layer1_outputs[12159];
    assign layer2_outputs[10107] = (layer1_outputs[9340]) | (layer1_outputs[782]);
    assign layer2_outputs[10108] = layer1_outputs[1509];
    assign layer2_outputs[10109] = layer1_outputs[1641];
    assign layer2_outputs[10110] = ~(layer1_outputs[2030]);
    assign layer2_outputs[10111] = (layer1_outputs[2815]) | (layer1_outputs[10252]);
    assign layer2_outputs[10112] = (layer1_outputs[7830]) & (layer1_outputs[9832]);
    assign layer2_outputs[10113] = ~((layer1_outputs[1768]) & (layer1_outputs[3598]));
    assign layer2_outputs[10114] = ~(layer1_outputs[156]);
    assign layer2_outputs[10115] = ~(layer1_outputs[1949]) | (layer1_outputs[11633]);
    assign layer2_outputs[10116] = ~(layer1_outputs[6909]) | (layer1_outputs[7019]);
    assign layer2_outputs[10117] = (layer1_outputs[6144]) & (layer1_outputs[5346]);
    assign layer2_outputs[10118] = layer1_outputs[3378];
    assign layer2_outputs[10119] = layer1_outputs[1825];
    assign layer2_outputs[10120] = ~((layer1_outputs[7733]) ^ (layer1_outputs[8649]));
    assign layer2_outputs[10121] = (layer1_outputs[5898]) ^ (layer1_outputs[5588]);
    assign layer2_outputs[10122] = (layer1_outputs[8475]) ^ (layer1_outputs[11585]);
    assign layer2_outputs[10123] = ~((layer1_outputs[4794]) ^ (layer1_outputs[11295]));
    assign layer2_outputs[10124] = (layer1_outputs[1745]) & (layer1_outputs[8143]);
    assign layer2_outputs[10125] = layer1_outputs[11666];
    assign layer2_outputs[10126] = (layer1_outputs[3989]) ^ (layer1_outputs[8065]);
    assign layer2_outputs[10127] = 1'b0;
    assign layer2_outputs[10128] = layer1_outputs[12407];
    assign layer2_outputs[10129] = (layer1_outputs[5976]) ^ (layer1_outputs[6852]);
    assign layer2_outputs[10130] = ~(layer1_outputs[4627]);
    assign layer2_outputs[10131] = ~(layer1_outputs[4084]);
    assign layer2_outputs[10132] = ~(layer1_outputs[3038]);
    assign layer2_outputs[10133] = layer1_outputs[10418];
    assign layer2_outputs[10134] = layer1_outputs[11325];
    assign layer2_outputs[10135] = layer1_outputs[3499];
    assign layer2_outputs[10136] = ~(layer1_outputs[12734]);
    assign layer2_outputs[10137] = (layer1_outputs[7915]) & ~(layer1_outputs[12264]);
    assign layer2_outputs[10138] = 1'b0;
    assign layer2_outputs[10139] = (layer1_outputs[5452]) & ~(layer1_outputs[1260]);
    assign layer2_outputs[10140] = (layer1_outputs[7431]) ^ (layer1_outputs[9140]);
    assign layer2_outputs[10141] = ~((layer1_outputs[12110]) ^ (layer1_outputs[11417]));
    assign layer2_outputs[10142] = layer1_outputs[940];
    assign layer2_outputs[10143] = (layer1_outputs[11515]) ^ (layer1_outputs[8523]);
    assign layer2_outputs[10144] = ~(layer1_outputs[5517]);
    assign layer2_outputs[10145] = ~((layer1_outputs[5135]) ^ (layer1_outputs[1197]));
    assign layer2_outputs[10146] = layer1_outputs[7541];
    assign layer2_outputs[10147] = layer1_outputs[9839];
    assign layer2_outputs[10148] = ~(layer1_outputs[3905]) | (layer1_outputs[9623]);
    assign layer2_outputs[10149] = ~(layer1_outputs[6346]) | (layer1_outputs[11304]);
    assign layer2_outputs[10150] = ~(layer1_outputs[3784]);
    assign layer2_outputs[10151] = layer1_outputs[10503];
    assign layer2_outputs[10152] = ~(layer1_outputs[4203]);
    assign layer2_outputs[10153] = layer1_outputs[1465];
    assign layer2_outputs[10154] = ~(layer1_outputs[910]);
    assign layer2_outputs[10155] = layer1_outputs[372];
    assign layer2_outputs[10156] = ~((layer1_outputs[9172]) & (layer1_outputs[4662]));
    assign layer2_outputs[10157] = ~(layer1_outputs[8229]);
    assign layer2_outputs[10158] = ~(layer1_outputs[62]) | (layer1_outputs[4955]);
    assign layer2_outputs[10159] = ~(layer1_outputs[162]);
    assign layer2_outputs[10160] = (layer1_outputs[2458]) ^ (layer1_outputs[1714]);
    assign layer2_outputs[10161] = (layer1_outputs[9528]) | (layer1_outputs[9831]);
    assign layer2_outputs[10162] = ~(layer1_outputs[10652]);
    assign layer2_outputs[10163] = ~(layer1_outputs[9026]);
    assign layer2_outputs[10164] = ~((layer1_outputs[5643]) & (layer1_outputs[3560]));
    assign layer2_outputs[10165] = ~(layer1_outputs[6879]);
    assign layer2_outputs[10166] = layer1_outputs[10837];
    assign layer2_outputs[10167] = layer1_outputs[11287];
    assign layer2_outputs[10168] = layer1_outputs[12652];
    assign layer2_outputs[10169] = (layer1_outputs[8341]) & ~(layer1_outputs[11392]);
    assign layer2_outputs[10170] = ~((layer1_outputs[3553]) | (layer1_outputs[6678]));
    assign layer2_outputs[10171] = ~(layer1_outputs[12205]);
    assign layer2_outputs[10172] = layer1_outputs[7985];
    assign layer2_outputs[10173] = (layer1_outputs[8320]) ^ (layer1_outputs[2168]);
    assign layer2_outputs[10174] = (layer1_outputs[897]) & ~(layer1_outputs[4348]);
    assign layer2_outputs[10175] = ~(layer1_outputs[5742]) | (layer1_outputs[6101]);
    assign layer2_outputs[10176] = ~(layer1_outputs[7141]);
    assign layer2_outputs[10177] = layer1_outputs[1843];
    assign layer2_outputs[10178] = ~(layer1_outputs[6494]);
    assign layer2_outputs[10179] = (layer1_outputs[10052]) | (layer1_outputs[10353]);
    assign layer2_outputs[10180] = ~(layer1_outputs[6970]) | (layer1_outputs[8333]);
    assign layer2_outputs[10181] = (layer1_outputs[1256]) & ~(layer1_outputs[7286]);
    assign layer2_outputs[10182] = ~(layer1_outputs[12316]) | (layer1_outputs[8297]);
    assign layer2_outputs[10183] = (layer1_outputs[5186]) & (layer1_outputs[3344]);
    assign layer2_outputs[10184] = layer1_outputs[465];
    assign layer2_outputs[10185] = (layer1_outputs[7211]) ^ (layer1_outputs[3327]);
    assign layer2_outputs[10186] = ~(layer1_outputs[9454]);
    assign layer2_outputs[10187] = layer1_outputs[6480];
    assign layer2_outputs[10188] = ~(layer1_outputs[11395]);
    assign layer2_outputs[10189] = (layer1_outputs[7495]) & ~(layer1_outputs[4867]);
    assign layer2_outputs[10190] = layer1_outputs[636];
    assign layer2_outputs[10191] = (layer1_outputs[9480]) & ~(layer1_outputs[10292]);
    assign layer2_outputs[10192] = ~(layer1_outputs[2728]);
    assign layer2_outputs[10193] = (layer1_outputs[12610]) | (layer1_outputs[12748]);
    assign layer2_outputs[10194] = ~(layer1_outputs[5425]);
    assign layer2_outputs[10195] = layer1_outputs[1096];
    assign layer2_outputs[10196] = (layer1_outputs[8324]) ^ (layer1_outputs[4452]);
    assign layer2_outputs[10197] = layer1_outputs[9570];
    assign layer2_outputs[10198] = (layer1_outputs[1517]) | (layer1_outputs[200]);
    assign layer2_outputs[10199] = layer1_outputs[10311];
    assign layer2_outputs[10200] = ~((layer1_outputs[7384]) ^ (layer1_outputs[10307]));
    assign layer2_outputs[10201] = ~(layer1_outputs[4085]);
    assign layer2_outputs[10202] = layer1_outputs[5509];
    assign layer2_outputs[10203] = layer1_outputs[8714];
    assign layer2_outputs[10204] = (layer1_outputs[12163]) & ~(layer1_outputs[5771]);
    assign layer2_outputs[10205] = ~((layer1_outputs[10084]) | (layer1_outputs[11746]));
    assign layer2_outputs[10206] = ~(layer1_outputs[7000]);
    assign layer2_outputs[10207] = (layer1_outputs[5966]) ^ (layer1_outputs[12151]);
    assign layer2_outputs[10208] = ~(layer1_outputs[1707]) | (layer1_outputs[5513]);
    assign layer2_outputs[10209] = ~(layer1_outputs[7578]) | (layer1_outputs[10501]);
    assign layer2_outputs[10210] = ~(layer1_outputs[5252]);
    assign layer2_outputs[10211] = ~((layer1_outputs[8758]) ^ (layer1_outputs[9526]));
    assign layer2_outputs[10212] = layer1_outputs[10923];
    assign layer2_outputs[10213] = ~(layer1_outputs[121]);
    assign layer2_outputs[10214] = layer1_outputs[4467];
    assign layer2_outputs[10215] = ~(layer1_outputs[8898]) | (layer1_outputs[4892]);
    assign layer2_outputs[10216] = ~(layer1_outputs[3155]);
    assign layer2_outputs[10217] = (layer1_outputs[8151]) | (layer1_outputs[3190]);
    assign layer2_outputs[10218] = ~(layer1_outputs[10208]) | (layer1_outputs[9087]);
    assign layer2_outputs[10219] = ~(layer1_outputs[2937]);
    assign layer2_outputs[10220] = ~(layer1_outputs[7989]);
    assign layer2_outputs[10221] = (layer1_outputs[10232]) ^ (layer1_outputs[1395]);
    assign layer2_outputs[10222] = layer1_outputs[8269];
    assign layer2_outputs[10223] = (layer1_outputs[7259]) & (layer1_outputs[2494]);
    assign layer2_outputs[10224] = ~(layer1_outputs[9335]);
    assign layer2_outputs[10225] = (layer1_outputs[2441]) & ~(layer1_outputs[2161]);
    assign layer2_outputs[10226] = ~((layer1_outputs[567]) & (layer1_outputs[6474]));
    assign layer2_outputs[10227] = ~(layer1_outputs[1899]);
    assign layer2_outputs[10228] = layer1_outputs[7529];
    assign layer2_outputs[10229] = ~(layer1_outputs[2391]);
    assign layer2_outputs[10230] = ~((layer1_outputs[6837]) & (layer1_outputs[411]));
    assign layer2_outputs[10231] = layer1_outputs[9114];
    assign layer2_outputs[10232] = ~(layer1_outputs[10150]) | (layer1_outputs[7335]);
    assign layer2_outputs[10233] = ~(layer1_outputs[12597]);
    assign layer2_outputs[10234] = layer1_outputs[8626];
    assign layer2_outputs[10235] = layer1_outputs[4124];
    assign layer2_outputs[10236] = ~((layer1_outputs[6873]) ^ (layer1_outputs[2173]));
    assign layer2_outputs[10237] = ~(layer1_outputs[4875]) | (layer1_outputs[8719]);
    assign layer2_outputs[10238] = (layer1_outputs[12268]) & (layer1_outputs[510]);
    assign layer2_outputs[10239] = (layer1_outputs[9450]) & ~(layer1_outputs[7498]);
    assign layer2_outputs[10240] = ~((layer1_outputs[5857]) & (layer1_outputs[6140]));
    assign layer2_outputs[10241] = ~(layer1_outputs[10203]);
    assign layer2_outputs[10242] = layer1_outputs[12449];
    assign layer2_outputs[10243] = layer1_outputs[6328];
    assign layer2_outputs[10244] = (layer1_outputs[12149]) ^ (layer1_outputs[7013]);
    assign layer2_outputs[10245] = ~(layer1_outputs[6656]) | (layer1_outputs[8836]);
    assign layer2_outputs[10246] = ~((layer1_outputs[12380]) ^ (layer1_outputs[7074]));
    assign layer2_outputs[10247] = ~(layer1_outputs[3261]);
    assign layer2_outputs[10248] = (layer1_outputs[12309]) & ~(layer1_outputs[10873]);
    assign layer2_outputs[10249] = (layer1_outputs[3167]) & (layer1_outputs[2477]);
    assign layer2_outputs[10250] = ~(layer1_outputs[2028]) | (layer1_outputs[12109]);
    assign layer2_outputs[10251] = layer1_outputs[11439];
    assign layer2_outputs[10252] = (layer1_outputs[9388]) & ~(layer1_outputs[11977]);
    assign layer2_outputs[10253] = ~((layer1_outputs[1213]) & (layer1_outputs[9171]));
    assign layer2_outputs[10254] = ~((layer1_outputs[12337]) | (layer1_outputs[10800]));
    assign layer2_outputs[10255] = layer1_outputs[9269];
    assign layer2_outputs[10256] = ~(layer1_outputs[2644]);
    assign layer2_outputs[10257] = layer1_outputs[9030];
    assign layer2_outputs[10258] = layer1_outputs[4995];
    assign layer2_outputs[10259] = (layer1_outputs[9410]) & ~(layer1_outputs[4869]);
    assign layer2_outputs[10260] = ~((layer1_outputs[2090]) & (layer1_outputs[7636]));
    assign layer2_outputs[10261] = ~((layer1_outputs[8636]) ^ (layer1_outputs[7380]));
    assign layer2_outputs[10262] = ~((layer1_outputs[7840]) | (layer1_outputs[5493]));
    assign layer2_outputs[10263] = ~((layer1_outputs[12408]) | (layer1_outputs[227]));
    assign layer2_outputs[10264] = (layer1_outputs[10452]) ^ (layer1_outputs[6227]);
    assign layer2_outputs[10265] = ~(layer1_outputs[3097]) | (layer1_outputs[3797]);
    assign layer2_outputs[10266] = ~(layer1_outputs[8692]) | (layer1_outputs[10259]);
    assign layer2_outputs[10267] = ~((layer1_outputs[10501]) | (layer1_outputs[5368]));
    assign layer2_outputs[10268] = ~((layer1_outputs[10125]) & (layer1_outputs[9399]));
    assign layer2_outputs[10269] = (layer1_outputs[7662]) | (layer1_outputs[7316]);
    assign layer2_outputs[10270] = layer1_outputs[10226];
    assign layer2_outputs[10271] = layer1_outputs[6567];
    assign layer2_outputs[10272] = layer1_outputs[10470];
    assign layer2_outputs[10273] = (layer1_outputs[8961]) | (layer1_outputs[7879]);
    assign layer2_outputs[10274] = (layer1_outputs[3829]) & (layer1_outputs[3839]);
    assign layer2_outputs[10275] = layer1_outputs[11931];
    assign layer2_outputs[10276] = (layer1_outputs[3482]) | (layer1_outputs[9137]);
    assign layer2_outputs[10277] = ~(layer1_outputs[3939]);
    assign layer2_outputs[10278] = ~(layer1_outputs[3596]) | (layer1_outputs[11654]);
    assign layer2_outputs[10279] = (layer1_outputs[3133]) & (layer1_outputs[10206]);
    assign layer2_outputs[10280] = layer1_outputs[2591];
    assign layer2_outputs[10281] = ~(layer1_outputs[1416]);
    assign layer2_outputs[10282] = layer1_outputs[7548];
    assign layer2_outputs[10283] = layer1_outputs[2412];
    assign layer2_outputs[10284] = ~((layer1_outputs[268]) ^ (layer1_outputs[6800]));
    assign layer2_outputs[10285] = ~((layer1_outputs[7519]) | (layer1_outputs[1450]));
    assign layer2_outputs[10286] = layer1_outputs[11125];
    assign layer2_outputs[10287] = (layer1_outputs[11571]) & (layer1_outputs[8020]);
    assign layer2_outputs[10288] = ~((layer1_outputs[8897]) ^ (layer1_outputs[2693]));
    assign layer2_outputs[10289] = ~(layer1_outputs[5811]);
    assign layer2_outputs[10290] = ~(layer1_outputs[8965]);
    assign layer2_outputs[10291] = ~(layer1_outputs[11476]);
    assign layer2_outputs[10292] = layer1_outputs[4285];
    assign layer2_outputs[10293] = ~(layer1_outputs[2904]);
    assign layer2_outputs[10294] = ~(layer1_outputs[9712]);
    assign layer2_outputs[10295] = (layer1_outputs[1347]) & (layer1_outputs[12]);
    assign layer2_outputs[10296] = (layer1_outputs[256]) | (layer1_outputs[6338]);
    assign layer2_outputs[10297] = (layer1_outputs[5584]) | (layer1_outputs[3974]);
    assign layer2_outputs[10298] = ~(layer1_outputs[2595]);
    assign layer2_outputs[10299] = (layer1_outputs[2151]) ^ (layer1_outputs[6350]);
    assign layer2_outputs[10300] = ~((layer1_outputs[9619]) ^ (layer1_outputs[8466]));
    assign layer2_outputs[10301] = layer1_outputs[11556];
    assign layer2_outputs[10302] = ~(layer1_outputs[579]);
    assign layer2_outputs[10303] = layer1_outputs[6429];
    assign layer2_outputs[10304] = (layer1_outputs[8750]) & (layer1_outputs[2588]);
    assign layer2_outputs[10305] = ~(layer1_outputs[499]) | (layer1_outputs[3156]);
    assign layer2_outputs[10306] = layer1_outputs[6280];
    assign layer2_outputs[10307] = (layer1_outputs[6680]) & (layer1_outputs[6011]);
    assign layer2_outputs[10308] = (layer1_outputs[9676]) ^ (layer1_outputs[5394]);
    assign layer2_outputs[10309] = (layer1_outputs[5502]) | (layer1_outputs[262]);
    assign layer2_outputs[10310] = (layer1_outputs[11034]) & (layer1_outputs[3362]);
    assign layer2_outputs[10311] = ~(layer1_outputs[6155]) | (layer1_outputs[5821]);
    assign layer2_outputs[10312] = ~(layer1_outputs[11049]);
    assign layer2_outputs[10313] = (layer1_outputs[7129]) & ~(layer1_outputs[3651]);
    assign layer2_outputs[10314] = ~(layer1_outputs[2104]);
    assign layer2_outputs[10315] = ~(layer1_outputs[5386]) | (layer1_outputs[4523]);
    assign layer2_outputs[10316] = (layer1_outputs[11334]) & ~(layer1_outputs[4967]);
    assign layer2_outputs[10317] = layer1_outputs[511];
    assign layer2_outputs[10318] = ~((layer1_outputs[11131]) | (layer1_outputs[8835]));
    assign layer2_outputs[10319] = layer1_outputs[2109];
    assign layer2_outputs[10320] = layer1_outputs[6578];
    assign layer2_outputs[10321] = ~(layer1_outputs[11563]);
    assign layer2_outputs[10322] = layer1_outputs[4741];
    assign layer2_outputs[10323] = layer1_outputs[9634];
    assign layer2_outputs[10324] = ~(layer1_outputs[1156]);
    assign layer2_outputs[10325] = (layer1_outputs[8414]) & (layer1_outputs[7713]);
    assign layer2_outputs[10326] = layer1_outputs[2085];
    assign layer2_outputs[10327] = layer1_outputs[10583];
    assign layer2_outputs[10328] = ~((layer1_outputs[6292]) & (layer1_outputs[11871]));
    assign layer2_outputs[10329] = ~(layer1_outputs[1827]) | (layer1_outputs[1808]);
    assign layer2_outputs[10330] = layer1_outputs[10977];
    assign layer2_outputs[10331] = ~(layer1_outputs[6960]);
    assign layer2_outputs[10332] = layer1_outputs[5004];
    assign layer2_outputs[10333] = ~(layer1_outputs[5125]);
    assign layer2_outputs[10334] = ~((layer1_outputs[6982]) & (layer1_outputs[3259]));
    assign layer2_outputs[10335] = ~(layer1_outputs[7391]);
    assign layer2_outputs[10336] = ~(layer1_outputs[9571]);
    assign layer2_outputs[10337] = (layer1_outputs[10720]) & (layer1_outputs[8513]);
    assign layer2_outputs[10338] = ~(layer1_outputs[9740]);
    assign layer2_outputs[10339] = (layer1_outputs[5938]) & ~(layer1_outputs[1407]);
    assign layer2_outputs[10340] = ~(layer1_outputs[10862]);
    assign layer2_outputs[10341] = layer1_outputs[10054];
    assign layer2_outputs[10342] = ~(layer1_outputs[6304]) | (layer1_outputs[12091]);
    assign layer2_outputs[10343] = ~(layer1_outputs[1083]) | (layer1_outputs[9461]);
    assign layer2_outputs[10344] = ~((layer1_outputs[3411]) | (layer1_outputs[6163]));
    assign layer2_outputs[10345] = layer1_outputs[3526];
    assign layer2_outputs[10346] = ~(layer1_outputs[6787]);
    assign layer2_outputs[10347] = ~((layer1_outputs[3426]) | (layer1_outputs[540]));
    assign layer2_outputs[10348] = ~((layer1_outputs[11678]) & (layer1_outputs[8797]));
    assign layer2_outputs[10349] = ~(layer1_outputs[4607]) | (layer1_outputs[8951]);
    assign layer2_outputs[10350] = (layer1_outputs[2897]) & ~(layer1_outputs[5138]);
    assign layer2_outputs[10351] = (layer1_outputs[2278]) ^ (layer1_outputs[5613]);
    assign layer2_outputs[10352] = ~(layer1_outputs[6005]);
    assign layer2_outputs[10353] = layer1_outputs[10599];
    assign layer2_outputs[10354] = ~(layer1_outputs[11685]) | (layer1_outputs[1240]);
    assign layer2_outputs[10355] = layer1_outputs[10056];
    assign layer2_outputs[10356] = layer1_outputs[11845];
    assign layer2_outputs[10357] = ~(layer1_outputs[7370]);
    assign layer2_outputs[10358] = layer1_outputs[9046];
    assign layer2_outputs[10359] = ~(layer1_outputs[9307]);
    assign layer2_outputs[10360] = ~(layer1_outputs[8545]);
    assign layer2_outputs[10361] = layer1_outputs[8563];
    assign layer2_outputs[10362] = ~((layer1_outputs[3108]) ^ (layer1_outputs[12780]));
    assign layer2_outputs[10363] = ~(layer1_outputs[3516]) | (layer1_outputs[7292]);
    assign layer2_outputs[10364] = ~(layer1_outputs[2224]);
    assign layer2_outputs[10365] = ~(layer1_outputs[10966]);
    assign layer2_outputs[10366] = layer1_outputs[11242];
    assign layer2_outputs[10367] = layer1_outputs[3424];
    assign layer2_outputs[10368] = ~(layer1_outputs[11166]);
    assign layer2_outputs[10369] = ~((layer1_outputs[1556]) ^ (layer1_outputs[10888]));
    assign layer2_outputs[10370] = (layer1_outputs[9473]) ^ (layer1_outputs[10972]);
    assign layer2_outputs[10371] = (layer1_outputs[11502]) & ~(layer1_outputs[5079]);
    assign layer2_outputs[10372] = layer1_outputs[10417];
    assign layer2_outputs[10373] = ~(layer1_outputs[8953]);
    assign layer2_outputs[10374] = (layer1_outputs[4546]) & ~(layer1_outputs[1775]);
    assign layer2_outputs[10375] = ~((layer1_outputs[11183]) & (layer1_outputs[1779]));
    assign layer2_outputs[10376] = (layer1_outputs[11211]) & ~(layer1_outputs[9313]);
    assign layer2_outputs[10377] = (layer1_outputs[6598]) & ~(layer1_outputs[5571]);
    assign layer2_outputs[10378] = (layer1_outputs[1504]) & ~(layer1_outputs[12332]);
    assign layer2_outputs[10379] = layer1_outputs[3244];
    assign layer2_outputs[10380] = layer1_outputs[9275];
    assign layer2_outputs[10381] = (layer1_outputs[3328]) ^ (layer1_outputs[2475]);
    assign layer2_outputs[10382] = layer1_outputs[1547];
    assign layer2_outputs[10383] = ~(layer1_outputs[7571]);
    assign layer2_outputs[10384] = ~(layer1_outputs[12701]);
    assign layer2_outputs[10385] = 1'b0;
    assign layer2_outputs[10386] = ~((layer1_outputs[4200]) ^ (layer1_outputs[6090]));
    assign layer2_outputs[10387] = ~((layer1_outputs[3116]) & (layer1_outputs[3424]));
    assign layer2_outputs[10388] = layer1_outputs[9816];
    assign layer2_outputs[10389] = (layer1_outputs[4350]) & ~(layer1_outputs[5120]);
    assign layer2_outputs[10390] = ~(layer1_outputs[9616]);
    assign layer2_outputs[10391] = ~((layer1_outputs[1132]) | (layer1_outputs[1047]));
    assign layer2_outputs[10392] = ~(layer1_outputs[2032]);
    assign layer2_outputs[10393] = ~(layer1_outputs[443]);
    assign layer2_outputs[10394] = ~((layer1_outputs[5020]) & (layer1_outputs[11671]));
    assign layer2_outputs[10395] = layer1_outputs[10226];
    assign layer2_outputs[10396] = (layer1_outputs[6565]) | (layer1_outputs[1711]);
    assign layer2_outputs[10397] = ~(layer1_outputs[5815]);
    assign layer2_outputs[10398] = layer1_outputs[12402];
    assign layer2_outputs[10399] = ~(layer1_outputs[1278]);
    assign layer2_outputs[10400] = ~(layer1_outputs[2539]);
    assign layer2_outputs[10401] = ~(layer1_outputs[6993]);
    assign layer2_outputs[10402] = ~(layer1_outputs[2896]);
    assign layer2_outputs[10403] = (layer1_outputs[8879]) & ~(layer1_outputs[6146]);
    assign layer2_outputs[10404] = (layer1_outputs[6779]) & ~(layer1_outputs[11401]);
    assign layer2_outputs[10405] = ~(layer1_outputs[1046]);
    assign layer2_outputs[10406] = ~(layer1_outputs[1887]);
    assign layer2_outputs[10407] = ~(layer1_outputs[6822]) | (layer1_outputs[11734]);
    assign layer2_outputs[10408] = ~(layer1_outputs[12223]);
    assign layer2_outputs[10409] = ~(layer1_outputs[5508]);
    assign layer2_outputs[10410] = ~((layer1_outputs[254]) & (layer1_outputs[1099]));
    assign layer2_outputs[10411] = (layer1_outputs[12545]) & (layer1_outputs[4729]);
    assign layer2_outputs[10412] = ~((layer1_outputs[521]) & (layer1_outputs[6318]));
    assign layer2_outputs[10413] = ~(layer1_outputs[5955]);
    assign layer2_outputs[10414] = layer1_outputs[4168];
    assign layer2_outputs[10415] = ~((layer1_outputs[7574]) ^ (layer1_outputs[1129]));
    assign layer2_outputs[10416] = ~(layer1_outputs[9812]);
    assign layer2_outputs[10417] = ~((layer1_outputs[10585]) ^ (layer1_outputs[5550]));
    assign layer2_outputs[10418] = ~(layer1_outputs[446]);
    assign layer2_outputs[10419] = (layer1_outputs[2942]) ^ (layer1_outputs[11450]);
    assign layer2_outputs[10420] = layer1_outputs[5734];
    assign layer2_outputs[10421] = layer1_outputs[2325];
    assign layer2_outputs[10422] = (layer1_outputs[10355]) & ~(layer1_outputs[12234]);
    assign layer2_outputs[10423] = ~(layer1_outputs[2431]) | (layer1_outputs[3677]);
    assign layer2_outputs[10424] = ~(layer1_outputs[2895]);
    assign layer2_outputs[10425] = layer1_outputs[4849];
    assign layer2_outputs[10426] = (layer1_outputs[1861]) & ~(layer1_outputs[4656]);
    assign layer2_outputs[10427] = (layer1_outputs[11310]) ^ (layer1_outputs[9850]);
    assign layer2_outputs[10428] = ~(layer1_outputs[12362]);
    assign layer2_outputs[10429] = layer1_outputs[10485];
    assign layer2_outputs[10430] = layer1_outputs[8811];
    assign layer2_outputs[10431] = (layer1_outputs[11898]) | (layer1_outputs[5195]);
    assign layer2_outputs[10432] = ~((layer1_outputs[9903]) & (layer1_outputs[430]));
    assign layer2_outputs[10433] = ~((layer1_outputs[6328]) | (layer1_outputs[6844]));
    assign layer2_outputs[10434] = (layer1_outputs[7408]) & (layer1_outputs[7920]);
    assign layer2_outputs[10435] = layer1_outputs[3149];
    assign layer2_outputs[10436] = (layer1_outputs[5922]) | (layer1_outputs[10752]);
    assign layer2_outputs[10437] = (layer1_outputs[12605]) | (layer1_outputs[11381]);
    assign layer2_outputs[10438] = (layer1_outputs[5928]) & ~(layer1_outputs[8529]);
    assign layer2_outputs[10439] = (layer1_outputs[7720]) & (layer1_outputs[4921]);
    assign layer2_outputs[10440] = (layer1_outputs[7626]) & ~(layer1_outputs[12189]);
    assign layer2_outputs[10441] = layer1_outputs[1102];
    assign layer2_outputs[10442] = layer1_outputs[11644];
    assign layer2_outputs[10443] = (layer1_outputs[1844]) ^ (layer1_outputs[9653]);
    assign layer2_outputs[10444] = layer1_outputs[8719];
    assign layer2_outputs[10445] = layer1_outputs[6572];
    assign layer2_outputs[10446] = ~((layer1_outputs[10737]) | (layer1_outputs[1763]));
    assign layer2_outputs[10447] = layer1_outputs[857];
    assign layer2_outputs[10448] = layer1_outputs[12554];
    assign layer2_outputs[10449] = ~((layer1_outputs[4594]) | (layer1_outputs[8392]));
    assign layer2_outputs[10450] = ~((layer1_outputs[2360]) | (layer1_outputs[10681]));
    assign layer2_outputs[10451] = ~(layer1_outputs[11689]) | (layer1_outputs[11899]);
    assign layer2_outputs[10452] = layer1_outputs[9074];
    assign layer2_outputs[10453] = ~(layer1_outputs[3401]);
    assign layer2_outputs[10454] = layer1_outputs[12404];
    assign layer2_outputs[10455] = (layer1_outputs[12183]) | (layer1_outputs[10625]);
    assign layer2_outputs[10456] = ~(layer1_outputs[2864]);
    assign layer2_outputs[10457] = ~(layer1_outputs[2120]);
    assign layer2_outputs[10458] = ~(layer1_outputs[3572]);
    assign layer2_outputs[10459] = ~(layer1_outputs[1719]);
    assign layer2_outputs[10460] = ~((layer1_outputs[9923]) | (layer1_outputs[5243]));
    assign layer2_outputs[10461] = ~((layer1_outputs[1222]) | (layer1_outputs[6073]));
    assign layer2_outputs[10462] = layer1_outputs[7443];
    assign layer2_outputs[10463] = ~((layer1_outputs[4111]) | (layer1_outputs[1906]));
    assign layer2_outputs[10464] = layer1_outputs[10690];
    assign layer2_outputs[10465] = layer1_outputs[1068];
    assign layer2_outputs[10466] = ~(layer1_outputs[3421]);
    assign layer2_outputs[10467] = layer1_outputs[3616];
    assign layer2_outputs[10468] = ~(layer1_outputs[9766]);
    assign layer2_outputs[10469] = ~(layer1_outputs[5547]);
    assign layer2_outputs[10470] = 1'b0;
    assign layer2_outputs[10471] = (layer1_outputs[10420]) & ~(layer1_outputs[7762]);
    assign layer2_outputs[10472] = ~((layer1_outputs[9235]) | (layer1_outputs[811]));
    assign layer2_outputs[10473] = ~((layer1_outputs[9589]) | (layer1_outputs[4138]));
    assign layer2_outputs[10474] = (layer1_outputs[7452]) | (layer1_outputs[664]);
    assign layer2_outputs[10475] = ~((layer1_outputs[11858]) | (layer1_outputs[9602]));
    assign layer2_outputs[10476] = ~(layer1_outputs[233]);
    assign layer2_outputs[10477] = layer1_outputs[4956];
    assign layer2_outputs[10478] = ~((layer1_outputs[1877]) ^ (layer1_outputs[3753]));
    assign layer2_outputs[10479] = layer1_outputs[4044];
    assign layer2_outputs[10480] = ~(layer1_outputs[12659]) | (layer1_outputs[6762]);
    assign layer2_outputs[10481] = ~(layer1_outputs[1877]);
    assign layer2_outputs[10482] = (layer1_outputs[10011]) & ~(layer1_outputs[5081]);
    assign layer2_outputs[10483] = layer1_outputs[1434];
    assign layer2_outputs[10484] = ~((layer1_outputs[5778]) & (layer1_outputs[10983]));
    assign layer2_outputs[10485] = ~(layer1_outputs[741]);
    assign layer2_outputs[10486] = ~(layer1_outputs[9710]) | (layer1_outputs[928]);
    assign layer2_outputs[10487] = layer1_outputs[7914];
    assign layer2_outputs[10488] = layer1_outputs[11191];
    assign layer2_outputs[10489] = layer1_outputs[8937];
    assign layer2_outputs[10490] = ~((layer1_outputs[4029]) | (layer1_outputs[6718]));
    assign layer2_outputs[10491] = (layer1_outputs[1926]) & ~(layer1_outputs[6590]);
    assign layer2_outputs[10492] = ~(layer1_outputs[1666]);
    assign layer2_outputs[10493] = layer1_outputs[12608];
    assign layer2_outputs[10494] = ~(layer1_outputs[1615]);
    assign layer2_outputs[10495] = (layer1_outputs[9325]) ^ (layer1_outputs[8010]);
    assign layer2_outputs[10496] = layer1_outputs[4092];
    assign layer2_outputs[10497] = (layer1_outputs[12360]) ^ (layer1_outputs[2392]);
    assign layer2_outputs[10498] = layer1_outputs[4210];
    assign layer2_outputs[10499] = layer1_outputs[769];
    assign layer2_outputs[10500] = ~((layer1_outputs[1100]) ^ (layer1_outputs[3964]));
    assign layer2_outputs[10501] = layer1_outputs[4761];
    assign layer2_outputs[10502] = 1'b1;
    assign layer2_outputs[10503] = ~(layer1_outputs[11023]) | (layer1_outputs[10135]);
    assign layer2_outputs[10504] = ~((layer1_outputs[677]) & (layer1_outputs[7996]));
    assign layer2_outputs[10505] = layer1_outputs[12308];
    assign layer2_outputs[10506] = layer1_outputs[11695];
    assign layer2_outputs[10507] = (layer1_outputs[3383]) ^ (layer1_outputs[10485]);
    assign layer2_outputs[10508] = (layer1_outputs[6280]) | (layer1_outputs[5507]);
    assign layer2_outputs[10509] = layer1_outputs[10046];
    assign layer2_outputs[10510] = (layer1_outputs[3940]) & ~(layer1_outputs[11378]);
    assign layer2_outputs[10511] = ~(layer1_outputs[8958]);
    assign layer2_outputs[10512] = (layer1_outputs[71]) | (layer1_outputs[7920]);
    assign layer2_outputs[10513] = layer1_outputs[9249];
    assign layer2_outputs[10514] = ~(layer1_outputs[948]);
    assign layer2_outputs[10515] = layer1_outputs[11183];
    assign layer2_outputs[10516] = (layer1_outputs[9097]) ^ (layer1_outputs[3474]);
    assign layer2_outputs[10517] = layer1_outputs[4946];
    assign layer2_outputs[10518] = ~(layer1_outputs[63]);
    assign layer2_outputs[10519] = (layer1_outputs[11910]) & ~(layer1_outputs[10913]);
    assign layer2_outputs[10520] = ~((layer1_outputs[12798]) & (layer1_outputs[1850]));
    assign layer2_outputs[10521] = ~(layer1_outputs[203]);
    assign layer2_outputs[10522] = ~(layer1_outputs[11952]);
    assign layer2_outputs[10523] = layer1_outputs[7374];
    assign layer2_outputs[10524] = layer1_outputs[8900];
    assign layer2_outputs[10525] = ~((layer1_outputs[2145]) ^ (layer1_outputs[9304]));
    assign layer2_outputs[10526] = layer1_outputs[5537];
    assign layer2_outputs[10527] = ~((layer1_outputs[1171]) | (layer1_outputs[8370]));
    assign layer2_outputs[10528] = ~((layer1_outputs[8294]) ^ (layer1_outputs[974]));
    assign layer2_outputs[10529] = ~(layer1_outputs[7672]);
    assign layer2_outputs[10530] = ~(layer1_outputs[6649]);
    assign layer2_outputs[10531] = layer1_outputs[9500];
    assign layer2_outputs[10532] = ~((layer1_outputs[4625]) & (layer1_outputs[7911]));
    assign layer2_outputs[10533] = (layer1_outputs[5065]) | (layer1_outputs[4587]);
    assign layer2_outputs[10534] = ~(layer1_outputs[5848]);
    assign layer2_outputs[10535] = ~(layer1_outputs[8638]) | (layer1_outputs[12195]);
    assign layer2_outputs[10536] = layer1_outputs[5817];
    assign layer2_outputs[10537] = ~(layer1_outputs[7283]) | (layer1_outputs[2622]);
    assign layer2_outputs[10538] = (layer1_outputs[9120]) & ~(layer1_outputs[3714]);
    assign layer2_outputs[10539] = (layer1_outputs[5114]) & ~(layer1_outputs[5521]);
    assign layer2_outputs[10540] = layer1_outputs[11801];
    assign layer2_outputs[10541] = ~(layer1_outputs[7881]);
    assign layer2_outputs[10542] = (layer1_outputs[6434]) | (layer1_outputs[10409]);
    assign layer2_outputs[10543] = (layer1_outputs[10115]) & (layer1_outputs[3507]);
    assign layer2_outputs[10544] = ~(layer1_outputs[11171]);
    assign layer2_outputs[10545] = layer1_outputs[11292];
    assign layer2_outputs[10546] = (layer1_outputs[4263]) & ~(layer1_outputs[5308]);
    assign layer2_outputs[10547] = (layer1_outputs[10013]) & (layer1_outputs[4046]);
    assign layer2_outputs[10548] = ~((layer1_outputs[1550]) ^ (layer1_outputs[11255]));
    assign layer2_outputs[10549] = ~((layer1_outputs[4119]) ^ (layer1_outputs[7394]));
    assign layer2_outputs[10550] = (layer1_outputs[11899]) ^ (layer1_outputs[406]);
    assign layer2_outputs[10551] = layer1_outputs[1237];
    assign layer2_outputs[10552] = ~(layer1_outputs[3128]);
    assign layer2_outputs[10553] = ~(layer1_outputs[10778]);
    assign layer2_outputs[10554] = layer1_outputs[560];
    assign layer2_outputs[10555] = ~((layer1_outputs[7963]) ^ (layer1_outputs[6030]));
    assign layer2_outputs[10556] = layer1_outputs[12353];
    assign layer2_outputs[10557] = layer1_outputs[5207];
    assign layer2_outputs[10558] = ~((layer1_outputs[4732]) | (layer1_outputs[12059]));
    assign layer2_outputs[10559] = ~(layer1_outputs[3663]);
    assign layer2_outputs[10560] = ~(layer1_outputs[10120]);
    assign layer2_outputs[10561] = ~(layer1_outputs[7778]);
    assign layer2_outputs[10562] = (layer1_outputs[2121]) & ~(layer1_outputs[10183]);
    assign layer2_outputs[10563] = (layer1_outputs[5767]) & ~(layer1_outputs[238]);
    assign layer2_outputs[10564] = layer1_outputs[2288];
    assign layer2_outputs[10565] = ~(layer1_outputs[2906]);
    assign layer2_outputs[10566] = ~(layer1_outputs[1328]);
    assign layer2_outputs[10567] = layer1_outputs[2022];
    assign layer2_outputs[10568] = ~(layer1_outputs[590]);
    assign layer2_outputs[10569] = layer1_outputs[563];
    assign layer2_outputs[10570] = ~((layer1_outputs[10421]) | (layer1_outputs[9874]));
    assign layer2_outputs[10571] = ~((layer1_outputs[6050]) & (layer1_outputs[2243]));
    assign layer2_outputs[10572] = ~((layer1_outputs[6540]) ^ (layer1_outputs[12453]));
    assign layer2_outputs[10573] = ~((layer1_outputs[3346]) | (layer1_outputs[4463]));
    assign layer2_outputs[10574] = ~(layer1_outputs[1917]);
    assign layer2_outputs[10575] = (layer1_outputs[5100]) | (layer1_outputs[6700]);
    assign layer2_outputs[10576] = layer1_outputs[1896];
    assign layer2_outputs[10577] = (layer1_outputs[3373]) & ~(layer1_outputs[5185]);
    assign layer2_outputs[10578] = (layer1_outputs[8854]) & ~(layer1_outputs[7341]);
    assign layer2_outputs[10579] = ~(layer1_outputs[9180]);
    assign layer2_outputs[10580] = (layer1_outputs[3035]) | (layer1_outputs[1414]);
    assign layer2_outputs[10581] = ~(layer1_outputs[5483]);
    assign layer2_outputs[10582] = (layer1_outputs[4876]) | (layer1_outputs[3660]);
    assign layer2_outputs[10583] = 1'b0;
    assign layer2_outputs[10584] = (layer1_outputs[2339]) & (layer1_outputs[11279]);
    assign layer2_outputs[10585] = ~((layer1_outputs[6080]) | (layer1_outputs[9224]));
    assign layer2_outputs[10586] = ~((layer1_outputs[4722]) & (layer1_outputs[7275]));
    assign layer2_outputs[10587] = (layer1_outputs[5330]) & (layer1_outputs[1726]);
    assign layer2_outputs[10588] = (layer1_outputs[1008]) ^ (layer1_outputs[2727]);
    assign layer2_outputs[10589] = layer1_outputs[12499];
    assign layer2_outputs[10590] = layer1_outputs[1614];
    assign layer2_outputs[10591] = ~(layer1_outputs[12694]) | (layer1_outputs[5946]);
    assign layer2_outputs[10592] = layer1_outputs[2517];
    assign layer2_outputs[10593] = layer1_outputs[7709];
    assign layer2_outputs[10594] = layer1_outputs[10967];
    assign layer2_outputs[10595] = ~((layer1_outputs[7962]) ^ (layer1_outputs[12756]));
    assign layer2_outputs[10596] = ~(layer1_outputs[12606]);
    assign layer2_outputs[10597] = (layer1_outputs[6492]) & (layer1_outputs[475]);
    assign layer2_outputs[10598] = ~(layer1_outputs[7516]);
    assign layer2_outputs[10599] = layer1_outputs[6575];
    assign layer2_outputs[10600] = layer1_outputs[8309];
    assign layer2_outputs[10601] = layer1_outputs[6364];
    assign layer2_outputs[10602] = (layer1_outputs[3312]) & ~(layer1_outputs[4779]);
    assign layer2_outputs[10603] = ~(layer1_outputs[2364]);
    assign layer2_outputs[10604] = (layer1_outputs[808]) & ~(layer1_outputs[2639]);
    assign layer2_outputs[10605] = (layer1_outputs[10249]) | (layer1_outputs[5505]);
    assign layer2_outputs[10606] = layer1_outputs[1820];
    assign layer2_outputs[10607] = ~(layer1_outputs[8644]);
    assign layer2_outputs[10608] = (layer1_outputs[1891]) & ~(layer1_outputs[12577]);
    assign layer2_outputs[10609] = ~(layer1_outputs[746]);
    assign layer2_outputs[10610] = (layer1_outputs[12769]) & ~(layer1_outputs[6266]);
    assign layer2_outputs[10611] = layer1_outputs[2965];
    assign layer2_outputs[10612] = layer1_outputs[9644];
    assign layer2_outputs[10613] = ~((layer1_outputs[7662]) & (layer1_outputs[6334]));
    assign layer2_outputs[10614] = layer1_outputs[5239];
    assign layer2_outputs[10615] = (layer1_outputs[7666]) ^ (layer1_outputs[12751]);
    assign layer2_outputs[10616] = ~(layer1_outputs[10847]) | (layer1_outputs[5016]);
    assign layer2_outputs[10617] = ~(layer1_outputs[2760]);
    assign layer2_outputs[10618] = ~((layer1_outputs[3150]) ^ (layer1_outputs[302]));
    assign layer2_outputs[10619] = (layer1_outputs[4274]) & ~(layer1_outputs[3927]);
    assign layer2_outputs[10620] = ~(layer1_outputs[12283]);
    assign layer2_outputs[10621] = ~(layer1_outputs[11660]);
    assign layer2_outputs[10622] = (layer1_outputs[5437]) & ~(layer1_outputs[11624]);
    assign layer2_outputs[10623] = layer1_outputs[1702];
    assign layer2_outputs[10624] = ~(layer1_outputs[11425]);
    assign layer2_outputs[10625] = layer1_outputs[4454];
    assign layer2_outputs[10626] = ~(layer1_outputs[676]);
    assign layer2_outputs[10627] = ~(layer1_outputs[600]);
    assign layer2_outputs[10628] = layer1_outputs[4797];
    assign layer2_outputs[10629] = ~(layer1_outputs[1115]);
    assign layer2_outputs[10630] = layer1_outputs[415];
    assign layer2_outputs[10631] = (layer1_outputs[8404]) & ~(layer1_outputs[9380]);
    assign layer2_outputs[10632] = (layer1_outputs[3693]) & (layer1_outputs[2721]);
    assign layer2_outputs[10633] = (layer1_outputs[8595]) ^ (layer1_outputs[3436]);
    assign layer2_outputs[10634] = (layer1_outputs[7394]) ^ (layer1_outputs[7683]);
    assign layer2_outputs[10635] = ~(layer1_outputs[10080]);
    assign layer2_outputs[10636] = (layer1_outputs[7725]) ^ (layer1_outputs[454]);
    assign layer2_outputs[10637] = ~((layer1_outputs[11152]) | (layer1_outputs[11065]));
    assign layer2_outputs[10638] = (layer1_outputs[9683]) | (layer1_outputs[1811]);
    assign layer2_outputs[10639] = layer1_outputs[12584];
    assign layer2_outputs[10640] = (layer1_outputs[9087]) & (layer1_outputs[6091]);
    assign layer2_outputs[10641] = (layer1_outputs[8637]) ^ (layer1_outputs[3969]);
    assign layer2_outputs[10642] = ~((layer1_outputs[6063]) ^ (layer1_outputs[8700]));
    assign layer2_outputs[10643] = ~(layer1_outputs[6731]);
    assign layer2_outputs[10644] = (layer1_outputs[6822]) ^ (layer1_outputs[3892]);
    assign layer2_outputs[10645] = (layer1_outputs[7063]) ^ (layer1_outputs[6897]);
    assign layer2_outputs[10646] = ~(layer1_outputs[4041]);
    assign layer2_outputs[10647] = layer1_outputs[12737];
    assign layer2_outputs[10648] = ~(layer1_outputs[3402]);
    assign layer2_outputs[10649] = ~(layer1_outputs[2728]);
    assign layer2_outputs[10650] = ~(layer1_outputs[8183]) | (layer1_outputs[138]);
    assign layer2_outputs[10651] = ~(layer1_outputs[6557]);
    assign layer2_outputs[10652] = (layer1_outputs[10149]) ^ (layer1_outputs[2859]);
    assign layer2_outputs[10653] = (layer1_outputs[5557]) ^ (layer1_outputs[8951]);
    assign layer2_outputs[10654] = (layer1_outputs[5798]) ^ (layer1_outputs[8612]);
    assign layer2_outputs[10655] = (layer1_outputs[12358]) ^ (layer1_outputs[1080]);
    assign layer2_outputs[10656] = ~(layer1_outputs[6342]) | (layer1_outputs[944]);
    assign layer2_outputs[10657] = layer1_outputs[12316];
    assign layer2_outputs[10658] = ~((layer1_outputs[574]) ^ (layer1_outputs[9568]));
    assign layer2_outputs[10659] = ~((layer1_outputs[6361]) & (layer1_outputs[5893]));
    assign layer2_outputs[10660] = layer1_outputs[10368];
    assign layer2_outputs[10661] = ~(layer1_outputs[4164]);
    assign layer2_outputs[10662] = (layer1_outputs[4513]) & ~(layer1_outputs[8541]);
    assign layer2_outputs[10663] = (layer1_outputs[2014]) & (layer1_outputs[4047]);
    assign layer2_outputs[10664] = (layer1_outputs[2225]) | (layer1_outputs[9646]);
    assign layer2_outputs[10665] = (layer1_outputs[11603]) ^ (layer1_outputs[12608]);
    assign layer2_outputs[10666] = (layer1_outputs[11653]) ^ (layer1_outputs[8170]);
    assign layer2_outputs[10667] = layer1_outputs[2608];
    assign layer2_outputs[10668] = (layer1_outputs[10583]) ^ (layer1_outputs[8102]);
    assign layer2_outputs[10669] = (layer1_outputs[10898]) & ~(layer1_outputs[3592]);
    assign layer2_outputs[10670] = ~(layer1_outputs[6454]);
    assign layer2_outputs[10671] = (layer1_outputs[10977]) & ~(layer1_outputs[4524]);
    assign layer2_outputs[10672] = (layer1_outputs[10999]) & ~(layer1_outputs[9140]);
    assign layer2_outputs[10673] = ~(layer1_outputs[986]);
    assign layer2_outputs[10674] = layer1_outputs[3591];
    assign layer2_outputs[10675] = ~(layer1_outputs[1288]);
    assign layer2_outputs[10676] = ~(layer1_outputs[7780]);
    assign layer2_outputs[10677] = ~((layer1_outputs[11636]) & (layer1_outputs[3970]));
    assign layer2_outputs[10678] = (layer1_outputs[5315]) | (layer1_outputs[4863]);
    assign layer2_outputs[10679] = (layer1_outputs[4737]) & (layer1_outputs[11607]);
    assign layer2_outputs[10680] = ~((layer1_outputs[4540]) ^ (layer1_outputs[7052]));
    assign layer2_outputs[10681] = ~((layer1_outputs[11961]) ^ (layer1_outputs[11236]));
    assign layer2_outputs[10682] = ~((layer1_outputs[1034]) | (layer1_outputs[4856]));
    assign layer2_outputs[10683] = ~(layer1_outputs[3600]);
    assign layer2_outputs[10684] = ~(layer1_outputs[1064]);
    assign layer2_outputs[10685] = ~(layer1_outputs[6495]);
    assign layer2_outputs[10686] = ~((layer1_outputs[9707]) & (layer1_outputs[10751]));
    assign layer2_outputs[10687] = ~((layer1_outputs[6499]) | (layer1_outputs[10139]));
    assign layer2_outputs[10688] = ~(layer1_outputs[6337]);
    assign layer2_outputs[10689] = layer1_outputs[9716];
    assign layer2_outputs[10690] = ~(layer1_outputs[9863]);
    assign layer2_outputs[10691] = (layer1_outputs[99]) & ~(layer1_outputs[7400]);
    assign layer2_outputs[10692] = ~((layer1_outputs[5276]) ^ (layer1_outputs[11123]));
    assign layer2_outputs[10693] = ~(layer1_outputs[6953]) | (layer1_outputs[2735]);
    assign layer2_outputs[10694] = layer1_outputs[5691];
    assign layer2_outputs[10695] = ~(layer1_outputs[4725]);
    assign layer2_outputs[10696] = ~(layer1_outputs[5687]) | (layer1_outputs[2507]);
    assign layer2_outputs[10697] = ~((layer1_outputs[11866]) & (layer1_outputs[2284]));
    assign layer2_outputs[10698] = ~(layer1_outputs[9276]) | (layer1_outputs[10098]);
    assign layer2_outputs[10699] = ~(layer1_outputs[2839]);
    assign layer2_outputs[10700] = ~((layer1_outputs[5729]) ^ (layer1_outputs[6225]));
    assign layer2_outputs[10701] = ~(layer1_outputs[12416]);
    assign layer2_outputs[10702] = layer1_outputs[8538];
    assign layer2_outputs[10703] = layer1_outputs[6381];
    assign layer2_outputs[10704] = ~((layer1_outputs[4789]) | (layer1_outputs[8277]));
    assign layer2_outputs[10705] = layer1_outputs[306];
    assign layer2_outputs[10706] = ~(layer1_outputs[10815]);
    assign layer2_outputs[10707] = (layer1_outputs[8618]) | (layer1_outputs[6213]);
    assign layer2_outputs[10708] = ~((layer1_outputs[1574]) & (layer1_outputs[4777]));
    assign layer2_outputs[10709] = ~(layer1_outputs[5302]);
    assign layer2_outputs[10710] = ~((layer1_outputs[1217]) & (layer1_outputs[2237]));
    assign layer2_outputs[10711] = layer1_outputs[6856];
    assign layer2_outputs[10712] = ~((layer1_outputs[5845]) & (layer1_outputs[10676]));
    assign layer2_outputs[10713] = layer1_outputs[12025];
    assign layer2_outputs[10714] = (layer1_outputs[9337]) ^ (layer1_outputs[9218]);
    assign layer2_outputs[10715] = ~(layer1_outputs[705]);
    assign layer2_outputs[10716] = (layer1_outputs[7563]) | (layer1_outputs[5151]);
    assign layer2_outputs[10717] = layer1_outputs[8439];
    assign layer2_outputs[10718] = ~((layer1_outputs[7742]) ^ (layer1_outputs[5555]));
    assign layer2_outputs[10719] = 1'b0;
    assign layer2_outputs[10720] = ~(layer1_outputs[5657]);
    assign layer2_outputs[10721] = layer1_outputs[6368];
    assign layer2_outputs[10722] = ~((layer1_outputs[3408]) ^ (layer1_outputs[2189]));
    assign layer2_outputs[10723] = ~((layer1_outputs[11945]) | (layer1_outputs[401]));
    assign layer2_outputs[10724] = ~((layer1_outputs[500]) & (layer1_outputs[2562]));
    assign layer2_outputs[10725] = ~((layer1_outputs[3221]) ^ (layer1_outputs[1711]));
    assign layer2_outputs[10726] = (layer1_outputs[688]) & ~(layer1_outputs[12710]);
    assign layer2_outputs[10727] = (layer1_outputs[4975]) & (layer1_outputs[5809]);
    assign layer2_outputs[10728] = layer1_outputs[2640];
    assign layer2_outputs[10729] = ~(layer1_outputs[10629]);
    assign layer2_outputs[10730] = ~(layer1_outputs[4136]) | (layer1_outputs[12665]);
    assign layer2_outputs[10731] = ~(layer1_outputs[286]);
    assign layer2_outputs[10732] = ~(layer1_outputs[2509]) | (layer1_outputs[11359]);
    assign layer2_outputs[10733] = layer1_outputs[6606];
    assign layer2_outputs[10734] = (layer1_outputs[5670]) ^ (layer1_outputs[11863]);
    assign layer2_outputs[10735] = ~(layer1_outputs[10071]);
    assign layer2_outputs[10736] = ~((layer1_outputs[6102]) ^ (layer1_outputs[9268]));
    assign layer2_outputs[10737] = ~(layer1_outputs[9057]);
    assign layer2_outputs[10738] = (layer1_outputs[1073]) & ~(layer1_outputs[5395]);
    assign layer2_outputs[10739] = ~((layer1_outputs[11224]) ^ (layer1_outputs[4108]));
    assign layer2_outputs[10740] = layer1_outputs[8646];
    assign layer2_outputs[10741] = layer1_outputs[1568];
    assign layer2_outputs[10742] = (layer1_outputs[5703]) ^ (layer1_outputs[3416]);
    assign layer2_outputs[10743] = (layer1_outputs[1602]) & ~(layer1_outputs[2973]);
    assign layer2_outputs[10744] = ~((layer1_outputs[4375]) & (layer1_outputs[780]));
    assign layer2_outputs[10745] = (layer1_outputs[9605]) ^ (layer1_outputs[3962]);
    assign layer2_outputs[10746] = layer1_outputs[4048];
    assign layer2_outputs[10747] = (layer1_outputs[8908]) & (layer1_outputs[1441]);
    assign layer2_outputs[10748] = layer1_outputs[12555];
    assign layer2_outputs[10749] = layer1_outputs[6764];
    assign layer2_outputs[10750] = ~(layer1_outputs[12439]);
    assign layer2_outputs[10751] = ~(layer1_outputs[8101]);
    assign layer2_outputs[10752] = layer1_outputs[5857];
    assign layer2_outputs[10753] = ~((layer1_outputs[9031]) & (layer1_outputs[7786]));
    assign layer2_outputs[10754] = layer1_outputs[6851];
    assign layer2_outputs[10755] = ~(layer1_outputs[2630]) | (layer1_outputs[3379]);
    assign layer2_outputs[10756] = ~(layer1_outputs[4418]);
    assign layer2_outputs[10757] = layer1_outputs[6496];
    assign layer2_outputs[10758] = (layer1_outputs[1051]) & (layer1_outputs[8072]);
    assign layer2_outputs[10759] = layer1_outputs[4276];
    assign layer2_outputs[10760] = ~(layer1_outputs[8055]);
    assign layer2_outputs[10761] = ~((layer1_outputs[11426]) & (layer1_outputs[9606]));
    assign layer2_outputs[10762] = ~(layer1_outputs[9299]) | (layer1_outputs[3631]);
    assign layer2_outputs[10763] = layer1_outputs[2894];
    assign layer2_outputs[10764] = ~(layer1_outputs[6003]);
    assign layer2_outputs[10765] = ~(layer1_outputs[3849]);
    assign layer2_outputs[10766] = ~(layer1_outputs[1789]);
    assign layer2_outputs[10767] = (layer1_outputs[1096]) & ~(layer1_outputs[4031]);
    assign layer2_outputs[10768] = layer1_outputs[3931];
    assign layer2_outputs[10769] = ~(layer1_outputs[7078]);
    assign layer2_outputs[10770] = ~(layer1_outputs[9592]);
    assign layer2_outputs[10771] = (layer1_outputs[9919]) & ~(layer1_outputs[8185]);
    assign layer2_outputs[10772] = (layer1_outputs[6354]) | (layer1_outputs[9665]);
    assign layer2_outputs[10773] = ~((layer1_outputs[7568]) ^ (layer1_outputs[2114]));
    assign layer2_outputs[10774] = ~(layer1_outputs[5168]);
    assign layer2_outputs[10775] = (layer1_outputs[6030]) & (layer1_outputs[150]);
    assign layer2_outputs[10776] = layer1_outputs[1776];
    assign layer2_outputs[10777] = layer1_outputs[5710];
    assign layer2_outputs[10778] = layer1_outputs[9286];
    assign layer2_outputs[10779] = layer1_outputs[2394];
    assign layer2_outputs[10780] = ~((layer1_outputs[7836]) & (layer1_outputs[9858]));
    assign layer2_outputs[10781] = ~(layer1_outputs[9687]);
    assign layer2_outputs[10782] = (layer1_outputs[10365]) | (layer1_outputs[1164]);
    assign layer2_outputs[10783] = ~((layer1_outputs[924]) | (layer1_outputs[10272]));
    assign layer2_outputs[10784] = layer1_outputs[3527];
    assign layer2_outputs[10785] = ~(layer1_outputs[506]) | (layer1_outputs[10534]);
    assign layer2_outputs[10786] = (layer1_outputs[9377]) & (layer1_outputs[9059]);
    assign layer2_outputs[10787] = (layer1_outputs[11510]) & ~(layer1_outputs[8683]);
    assign layer2_outputs[10788] = ~((layer1_outputs[12344]) ^ (layer1_outputs[6685]));
    assign layer2_outputs[10789] = layer1_outputs[1452];
    assign layer2_outputs[10790] = layer1_outputs[8847];
    assign layer2_outputs[10791] = ~(layer1_outputs[7707]) | (layer1_outputs[5072]);
    assign layer2_outputs[10792] = layer1_outputs[785];
    assign layer2_outputs[10793] = (layer1_outputs[9079]) & (layer1_outputs[9869]);
    assign layer2_outputs[10794] = (layer1_outputs[122]) | (layer1_outputs[12787]);
    assign layer2_outputs[10795] = ~(layer1_outputs[4270]) | (layer1_outputs[5285]);
    assign layer2_outputs[10796] = ~(layer1_outputs[1200]);
    assign layer2_outputs[10797] = ~(layer1_outputs[12736]) | (layer1_outputs[12723]);
    assign layer2_outputs[10798] = ~(layer1_outputs[3456]);
    assign layer2_outputs[10799] = ~(layer1_outputs[3225]);
    assign layer2_outputs[10800] = ~((layer1_outputs[10656]) ^ (layer1_outputs[8729]));
    assign layer2_outputs[10801] = ~((layer1_outputs[3479]) | (layer1_outputs[2454]));
    assign layer2_outputs[10802] = ~((layer1_outputs[8672]) ^ (layer1_outputs[966]));
    assign layer2_outputs[10803] = (layer1_outputs[8678]) ^ (layer1_outputs[7316]);
    assign layer2_outputs[10804] = ~((layer1_outputs[2186]) & (layer1_outputs[4106]));
    assign layer2_outputs[10805] = (layer1_outputs[3370]) ^ (layer1_outputs[3251]);
    assign layer2_outputs[10806] = ~(layer1_outputs[3253]);
    assign layer2_outputs[10807] = (layer1_outputs[7277]) ^ (layer1_outputs[6451]);
    assign layer2_outputs[10808] = ~(layer1_outputs[10003]);
    assign layer2_outputs[10809] = ~(layer1_outputs[5031]);
    assign layer2_outputs[10810] = ~((layer1_outputs[10194]) ^ (layer1_outputs[12624]));
    assign layer2_outputs[10811] = ~(layer1_outputs[4638]);
    assign layer2_outputs[10812] = ~((layer1_outputs[2887]) ^ (layer1_outputs[3090]));
    assign layer2_outputs[10813] = (layer1_outputs[3765]) & (layer1_outputs[7511]);
    assign layer2_outputs[10814] = layer1_outputs[5077];
    assign layer2_outputs[10815] = ~(layer1_outputs[3393]);
    assign layer2_outputs[10816] = ~(layer1_outputs[5116]) | (layer1_outputs[1936]);
    assign layer2_outputs[10817] = ~(layer1_outputs[2664]);
    assign layer2_outputs[10818] = ~(layer1_outputs[11759]);
    assign layer2_outputs[10819] = ~(layer1_outputs[8753]);
    assign layer2_outputs[10820] = ~((layer1_outputs[1669]) & (layer1_outputs[11856]));
    assign layer2_outputs[10821] = ~(layer1_outputs[6932]);
    assign layer2_outputs[10822] = (layer1_outputs[4712]) & ~(layer1_outputs[7669]);
    assign layer2_outputs[10823] = ~(layer1_outputs[900]);
    assign layer2_outputs[10824] = ~(layer1_outputs[11247]) | (layer1_outputs[5822]);
    assign layer2_outputs[10825] = ~(layer1_outputs[9808]);
    assign layer2_outputs[10826] = 1'b0;
    assign layer2_outputs[10827] = layer1_outputs[980];
    assign layer2_outputs[10828] = ~(layer1_outputs[4712]);
    assign layer2_outputs[10829] = ~(layer1_outputs[7877]) | (layer1_outputs[249]);
    assign layer2_outputs[10830] = ~(layer1_outputs[9963]) | (layer1_outputs[5607]);
    assign layer2_outputs[10831] = (layer1_outputs[11852]) & (layer1_outputs[9829]);
    assign layer2_outputs[10832] = ~((layer1_outputs[10023]) | (layer1_outputs[128]));
    assign layer2_outputs[10833] = ~((layer1_outputs[9417]) | (layer1_outputs[2264]));
    assign layer2_outputs[10834] = layer1_outputs[3819];
    assign layer2_outputs[10835] = (layer1_outputs[9556]) ^ (layer1_outputs[8701]);
    assign layer2_outputs[10836] = layer1_outputs[74];
    assign layer2_outputs[10837] = ~(layer1_outputs[4674]);
    assign layer2_outputs[10838] = layer1_outputs[278];
    assign layer2_outputs[10839] = ~(layer1_outputs[12463]);
    assign layer2_outputs[10840] = layer1_outputs[879];
    assign layer2_outputs[10841] = ~(layer1_outputs[2914]) | (layer1_outputs[379]);
    assign layer2_outputs[10842] = ~(layer1_outputs[12052]);
    assign layer2_outputs[10843] = ~(layer1_outputs[9459]);
    assign layer2_outputs[10844] = ~((layer1_outputs[2526]) ^ (layer1_outputs[1961]));
    assign layer2_outputs[10845] = ~(layer1_outputs[4535]);
    assign layer2_outputs[10846] = layer1_outputs[2578];
    assign layer2_outputs[10847] = ~(layer1_outputs[10611]);
    assign layer2_outputs[10848] = ~(layer1_outputs[4802]);
    assign layer2_outputs[10849] = ~((layer1_outputs[6178]) ^ (layer1_outputs[1879]));
    assign layer2_outputs[10850] = ~(layer1_outputs[11768]);
    assign layer2_outputs[10851] = ~(layer1_outputs[3757]);
    assign layer2_outputs[10852] = layer1_outputs[2112];
    assign layer2_outputs[10853] = (layer1_outputs[2920]) ^ (layer1_outputs[11150]);
    assign layer2_outputs[10854] = (layer1_outputs[11996]) | (layer1_outputs[9948]);
    assign layer2_outputs[10855] = layer1_outputs[6295];
    assign layer2_outputs[10856] = ~((layer1_outputs[8432]) | (layer1_outputs[9802]));
    assign layer2_outputs[10857] = layer1_outputs[4178];
    assign layer2_outputs[10858] = ~((layer1_outputs[12763]) | (layer1_outputs[237]));
    assign layer2_outputs[10859] = ~((layer1_outputs[4181]) ^ (layer1_outputs[11419]));
    assign layer2_outputs[10860] = layer1_outputs[2181];
    assign layer2_outputs[10861] = (layer1_outputs[9559]) ^ (layer1_outputs[4544]);
    assign layer2_outputs[10862] = ~((layer1_outputs[8845]) ^ (layer1_outputs[1671]));
    assign layer2_outputs[10863] = layer1_outputs[2472];
    assign layer2_outputs[10864] = ~((layer1_outputs[7099]) & (layer1_outputs[1725]));
    assign layer2_outputs[10865] = ~(layer1_outputs[2882]);
    assign layer2_outputs[10866] = ~(layer1_outputs[976]);
    assign layer2_outputs[10867] = ~((layer1_outputs[12438]) | (layer1_outputs[2469]));
    assign layer2_outputs[10868] = ~(layer1_outputs[1420]) | (layer1_outputs[11509]);
    assign layer2_outputs[10869] = ~((layer1_outputs[8179]) ^ (layer1_outputs[8039]));
    assign layer2_outputs[10870] = layer1_outputs[4707];
    assign layer2_outputs[10871] = (layer1_outputs[621]) & (layer1_outputs[2441]);
    assign layer2_outputs[10872] = ~(layer1_outputs[6354]);
    assign layer2_outputs[10873] = ~((layer1_outputs[2696]) ^ (layer1_outputs[3517]));
    assign layer2_outputs[10874] = ~(layer1_outputs[124]);
    assign layer2_outputs[10875] = layer1_outputs[3845];
    assign layer2_outputs[10876] = ~(layer1_outputs[8105]);
    assign layer2_outputs[10877] = layer1_outputs[11698];
    assign layer2_outputs[10878] = ~((layer1_outputs[11234]) & (layer1_outputs[98]));
    assign layer2_outputs[10879] = (layer1_outputs[2718]) | (layer1_outputs[108]);
    assign layer2_outputs[10880] = ~((layer1_outputs[11629]) & (layer1_outputs[6295]));
    assign layer2_outputs[10881] = ~(layer1_outputs[4498]);
    assign layer2_outputs[10882] = (layer1_outputs[10748]) & ~(layer1_outputs[7715]);
    assign layer2_outputs[10883] = (layer1_outputs[2051]) ^ (layer1_outputs[7358]);
    assign layer2_outputs[10884] = ~(layer1_outputs[6213]);
    assign layer2_outputs[10885] = (layer1_outputs[2347]) & (layer1_outputs[1492]);
    assign layer2_outputs[10886] = (layer1_outputs[4640]) & (layer1_outputs[4084]);
    assign layer2_outputs[10887] = ~((layer1_outputs[12387]) ^ (layer1_outputs[10138]));
    assign layer2_outputs[10888] = (layer1_outputs[5202]) & ~(layer1_outputs[2896]);
    assign layer2_outputs[10889] = layer1_outputs[2079];
    assign layer2_outputs[10890] = layer1_outputs[9343];
    assign layer2_outputs[10891] = layer1_outputs[11229];
    assign layer2_outputs[10892] = ~(layer1_outputs[11752]);
    assign layer2_outputs[10893] = layer1_outputs[4061];
    assign layer2_outputs[10894] = ~(layer1_outputs[3747]);
    assign layer2_outputs[10895] = ~(layer1_outputs[2012]) | (layer1_outputs[3264]);
    assign layer2_outputs[10896] = ~((layer1_outputs[5466]) ^ (layer1_outputs[929]));
    assign layer2_outputs[10897] = (layer1_outputs[9407]) ^ (layer1_outputs[11964]);
    assign layer2_outputs[10898] = (layer1_outputs[7877]) ^ (layer1_outputs[5639]);
    assign layer2_outputs[10899] = layer1_outputs[6658];
    assign layer2_outputs[10900] = ~(layer1_outputs[3550]);
    assign layer2_outputs[10901] = layer1_outputs[10545];
    assign layer2_outputs[10902] = ~((layer1_outputs[4749]) | (layer1_outputs[10645]));
    assign layer2_outputs[10903] = ~(layer1_outputs[5960]);
    assign layer2_outputs[10904] = ~(layer1_outputs[10712]);
    assign layer2_outputs[10905] = ~(layer1_outputs[12427]);
    assign layer2_outputs[10906] = ~(layer1_outputs[11189]);
    assign layer2_outputs[10907] = ~(layer1_outputs[1079]);
    assign layer2_outputs[10908] = ~(layer1_outputs[7798]);
    assign layer2_outputs[10909] = (layer1_outputs[11915]) & ~(layer1_outputs[4912]);
    assign layer2_outputs[10910] = ~(layer1_outputs[7103]);
    assign layer2_outputs[10911] = ~((layer1_outputs[5066]) & (layer1_outputs[2983]));
    assign layer2_outputs[10912] = ~(layer1_outputs[2093]);
    assign layer2_outputs[10913] = layer1_outputs[10718];
    assign layer2_outputs[10914] = (layer1_outputs[10057]) & ~(layer1_outputs[9627]);
    assign layer2_outputs[10915] = ~(layer1_outputs[5349]);
    assign layer2_outputs[10916] = ~(layer1_outputs[10689]);
    assign layer2_outputs[10917] = ~(layer1_outputs[9868]) | (layer1_outputs[8989]);
    assign layer2_outputs[10918] = ~(layer1_outputs[10765]) | (layer1_outputs[10154]);
    assign layer2_outputs[10919] = layer1_outputs[5155];
    assign layer2_outputs[10920] = layer1_outputs[8085];
    assign layer2_outputs[10921] = ~(layer1_outputs[7758]);
    assign layer2_outputs[10922] = ~(layer1_outputs[4439]);
    assign layer2_outputs[10923] = ~((layer1_outputs[6879]) | (layer1_outputs[7289]));
    assign layer2_outputs[10924] = layer1_outputs[6853];
    assign layer2_outputs[10925] = ~((layer1_outputs[286]) ^ (layer1_outputs[1287]));
    assign layer2_outputs[10926] = (layer1_outputs[450]) ^ (layer1_outputs[4450]);
    assign layer2_outputs[10927] = (layer1_outputs[3639]) & (layer1_outputs[6994]);
    assign layer2_outputs[10928] = ~((layer1_outputs[6535]) | (layer1_outputs[6409]));
    assign layer2_outputs[10929] = (layer1_outputs[1904]) ^ (layer1_outputs[7906]);
    assign layer2_outputs[10930] = ~(layer1_outputs[8512]);
    assign layer2_outputs[10931] = layer1_outputs[12367];
    assign layer2_outputs[10932] = ~(layer1_outputs[4836]) | (layer1_outputs[4189]);
    assign layer2_outputs[10933] = layer1_outputs[10659];
    assign layer2_outputs[10934] = layer1_outputs[5918];
    assign layer2_outputs[10935] = ~((layer1_outputs[6713]) ^ (layer1_outputs[11923]));
    assign layer2_outputs[10936] = ~((layer1_outputs[3352]) | (layer1_outputs[4769]));
    assign layer2_outputs[10937] = layer1_outputs[2204];
    assign layer2_outputs[10938] = ~(layer1_outputs[5223]);
    assign layer2_outputs[10939] = (layer1_outputs[5334]) & (layer1_outputs[6858]);
    assign layer2_outputs[10940] = ~((layer1_outputs[7592]) ^ (layer1_outputs[8252]));
    assign layer2_outputs[10941] = ~(layer1_outputs[685]);
    assign layer2_outputs[10942] = layer1_outputs[9597];
    assign layer2_outputs[10943] = layer1_outputs[955];
    assign layer2_outputs[10944] = ~(layer1_outputs[8782]) | (layer1_outputs[307]);
    assign layer2_outputs[10945] = layer1_outputs[6750];
    assign layer2_outputs[10946] = layer1_outputs[4003];
    assign layer2_outputs[10947] = ~((layer1_outputs[2016]) ^ (layer1_outputs[8447]));
    assign layer2_outputs[10948] = ~(layer1_outputs[5075]);
    assign layer2_outputs[10949] = ~(layer1_outputs[1870]);
    assign layer2_outputs[10950] = ~(layer1_outputs[10185]) | (layer1_outputs[10620]);
    assign layer2_outputs[10951] = ~(layer1_outputs[8220]);
    assign layer2_outputs[10952] = ~(layer1_outputs[2531]);
    assign layer2_outputs[10953] = layer1_outputs[8641];
    assign layer2_outputs[10954] = ~(layer1_outputs[12220]);
    assign layer2_outputs[10955] = layer1_outputs[10813];
    assign layer2_outputs[10956] = ~((layer1_outputs[6520]) ^ (layer1_outputs[12100]));
    assign layer2_outputs[10957] = (layer1_outputs[2248]) & ~(layer1_outputs[11979]);
    assign layer2_outputs[10958] = layer1_outputs[6064];
    assign layer2_outputs[10959] = ~(layer1_outputs[11619]);
    assign layer2_outputs[10960] = (layer1_outputs[11896]) ^ (layer1_outputs[11854]);
    assign layer2_outputs[10961] = ~(layer1_outputs[4883]);
    assign layer2_outputs[10962] = (layer1_outputs[4413]) ^ (layer1_outputs[5836]);
    assign layer2_outputs[10963] = ~((layer1_outputs[4829]) ^ (layer1_outputs[6939]));
    assign layer2_outputs[10964] = ~(layer1_outputs[2572]);
    assign layer2_outputs[10965] = (layer1_outputs[12441]) & ~(layer1_outputs[11448]);
    assign layer2_outputs[10966] = ~(layer1_outputs[4582]) | (layer1_outputs[1932]);
    assign layer2_outputs[10967] = (layer1_outputs[9433]) | (layer1_outputs[2415]);
    assign layer2_outputs[10968] = ~((layer1_outputs[6680]) ^ (layer1_outputs[959]));
    assign layer2_outputs[10969] = ~((layer1_outputs[1757]) ^ (layer1_outputs[4074]));
    assign layer2_outputs[10970] = (layer1_outputs[4561]) & ~(layer1_outputs[6238]);
    assign layer2_outputs[10971] = layer1_outputs[9723];
    assign layer2_outputs[10972] = layer1_outputs[8811];
    assign layer2_outputs[10973] = (layer1_outputs[9705]) | (layer1_outputs[12450]);
    assign layer2_outputs[10974] = (layer1_outputs[7756]) & ~(layer1_outputs[3700]);
    assign layer2_outputs[10975] = layer1_outputs[6367];
    assign layer2_outputs[10976] = layer1_outputs[10022];
    assign layer2_outputs[10977] = layer1_outputs[4577];
    assign layer2_outputs[10978] = (layer1_outputs[1954]) ^ (layer1_outputs[9828]);
    assign layer2_outputs[10979] = layer1_outputs[2087];
    assign layer2_outputs[10980] = ~(layer1_outputs[12764]);
    assign layer2_outputs[10981] = (layer1_outputs[1710]) & ~(layer1_outputs[979]);
    assign layer2_outputs[10982] = layer1_outputs[1532];
    assign layer2_outputs[10983] = layer1_outputs[7330];
    assign layer2_outputs[10984] = ~(layer1_outputs[2911]) | (layer1_outputs[12650]);
    assign layer2_outputs[10985] = layer1_outputs[10907];
    assign layer2_outputs[10986] = ~(layer1_outputs[4985]);
    assign layer2_outputs[10987] = layer1_outputs[718];
    assign layer2_outputs[10988] = layer1_outputs[7041];
    assign layer2_outputs[10989] = ~(layer1_outputs[10665]);
    assign layer2_outputs[10990] = layer1_outputs[12699];
    assign layer2_outputs[10991] = ~((layer1_outputs[7240]) ^ (layer1_outputs[3178]));
    assign layer2_outputs[10992] = layer1_outputs[6723];
    assign layer2_outputs[10993] = layer1_outputs[6018];
    assign layer2_outputs[10994] = (layer1_outputs[6168]) & ~(layer1_outputs[167]);
    assign layer2_outputs[10995] = ~(layer1_outputs[8033]);
    assign layer2_outputs[10996] = (layer1_outputs[11861]) & (layer1_outputs[5792]);
    assign layer2_outputs[10997] = (layer1_outputs[4693]) | (layer1_outputs[3924]);
    assign layer2_outputs[10998] = ~((layer1_outputs[2010]) ^ (layer1_outputs[7995]));
    assign layer2_outputs[10999] = ~((layer1_outputs[9236]) ^ (layer1_outputs[6552]));
    assign layer2_outputs[11000] = layer1_outputs[10725];
    assign layer2_outputs[11001] = ~(layer1_outputs[12417]);
    assign layer2_outputs[11002] = (layer1_outputs[2078]) & ~(layer1_outputs[7787]);
    assign layer2_outputs[11003] = ~(layer1_outputs[4631]);
    assign layer2_outputs[11004] = (layer1_outputs[1098]) | (layer1_outputs[4830]);
    assign layer2_outputs[11005] = layer1_outputs[4752];
    assign layer2_outputs[11006] = ~(layer1_outputs[8567]);
    assign layer2_outputs[11007] = layer1_outputs[11373];
    assign layer2_outputs[11008] = ~((layer1_outputs[8942]) & (layer1_outputs[10379]));
    assign layer2_outputs[11009] = ~(layer1_outputs[11198]) | (layer1_outputs[2177]);
    assign layer2_outputs[11010] = ~(layer1_outputs[1017]);
    assign layer2_outputs[11011] = ~(layer1_outputs[4654]) | (layer1_outputs[11935]);
    assign layer2_outputs[11012] = (layer1_outputs[2924]) & (layer1_outputs[9427]);
    assign layer2_outputs[11013] = (layer1_outputs[216]) & ~(layer1_outputs[5407]);
    assign layer2_outputs[11014] = ~((layer1_outputs[2073]) & (layer1_outputs[591]));
    assign layer2_outputs[11015] = (layer1_outputs[2141]) & (layer1_outputs[4722]);
    assign layer2_outputs[11016] = (layer1_outputs[3730]) & ~(layer1_outputs[2209]);
    assign layer2_outputs[11017] = ~((layer1_outputs[3720]) & (layer1_outputs[4069]));
    assign layer2_outputs[11018] = ~((layer1_outputs[11277]) & (layer1_outputs[7950]));
    assign layer2_outputs[11019] = (layer1_outputs[3288]) | (layer1_outputs[12153]);
    assign layer2_outputs[11020] = (layer1_outputs[10827]) & ~(layer1_outputs[1037]);
    assign layer2_outputs[11021] = ~(layer1_outputs[11732]);
    assign layer2_outputs[11022] = layer1_outputs[2550];
    assign layer2_outputs[11023] = ~(layer1_outputs[11353]);
    assign layer2_outputs[11024] = (layer1_outputs[4272]) & ~(layer1_outputs[7054]);
    assign layer2_outputs[11025] = ~((layer1_outputs[465]) ^ (layer1_outputs[2938]));
    assign layer2_outputs[11026] = ~(layer1_outputs[5933]) | (layer1_outputs[696]);
    assign layer2_outputs[11027] = ~((layer1_outputs[12218]) & (layer1_outputs[7823]));
    assign layer2_outputs[11028] = layer1_outputs[8661];
    assign layer2_outputs[11029] = layer1_outputs[3394];
    assign layer2_outputs[11030] = (layer1_outputs[6390]) ^ (layer1_outputs[8005]);
    assign layer2_outputs[11031] = 1'b0;
    assign layer2_outputs[11032] = ~(layer1_outputs[5457]);
    assign layer2_outputs[11033] = (layer1_outputs[1655]) ^ (layer1_outputs[3076]);
    assign layer2_outputs[11034] = ~((layer1_outputs[5867]) | (layer1_outputs[1507]));
    assign layer2_outputs[11035] = ~((layer1_outputs[5884]) | (layer1_outputs[12582]));
    assign layer2_outputs[11036] = ~(layer1_outputs[7735]);
    assign layer2_outputs[11037] = ~((layer1_outputs[3380]) ^ (layer1_outputs[11676]));
    assign layer2_outputs[11038] = ~(layer1_outputs[11177]);
    assign layer2_outputs[11039] = ~(layer1_outputs[12078]);
    assign layer2_outputs[11040] = (layer1_outputs[1069]) ^ (layer1_outputs[498]);
    assign layer2_outputs[11041] = ~(layer1_outputs[8287]);
    assign layer2_outputs[11042] = ~(layer1_outputs[6585]);
    assign layer2_outputs[11043] = 1'b1;
    assign layer2_outputs[11044] = ~(layer1_outputs[4088]);
    assign layer2_outputs[11045] = (layer1_outputs[12288]) & ~(layer1_outputs[10560]);
    assign layer2_outputs[11046] = ~(layer1_outputs[8017]);
    assign layer2_outputs[11047] = (layer1_outputs[259]) & ~(layer1_outputs[70]);
    assign layer2_outputs[11048] = ~(layer1_outputs[9155]);
    assign layer2_outputs[11049] = layer1_outputs[11144];
    assign layer2_outputs[11050] = layer1_outputs[10912];
    assign layer2_outputs[11051] = layer1_outputs[6965];
    assign layer2_outputs[11052] = ~((layer1_outputs[6324]) & (layer1_outputs[9159]));
    assign layer2_outputs[11053] = ~(layer1_outputs[525]);
    assign layer2_outputs[11054] = ~((layer1_outputs[3955]) ^ (layer1_outputs[7329]));
    assign layer2_outputs[11055] = layer1_outputs[6760];
    assign layer2_outputs[11056] = ~(layer1_outputs[4792]) | (layer1_outputs[1885]);
    assign layer2_outputs[11057] = ~(layer1_outputs[10051]);
    assign layer2_outputs[11058] = layer1_outputs[977];
    assign layer2_outputs[11059] = layer1_outputs[5598];
    assign layer2_outputs[11060] = ~(layer1_outputs[2753]);
    assign layer2_outputs[11061] = (layer1_outputs[2797]) & ~(layer1_outputs[1594]);
    assign layer2_outputs[11062] = (layer1_outputs[5665]) ^ (layer1_outputs[8343]);
    assign layer2_outputs[11063] = (layer1_outputs[9389]) & (layer1_outputs[8013]);
    assign layer2_outputs[11064] = (layer1_outputs[10978]) & ~(layer1_outputs[9158]);
    assign layer2_outputs[11065] = (layer1_outputs[5298]) & ~(layer1_outputs[2062]);
    assign layer2_outputs[11066] = layer1_outputs[10077];
    assign layer2_outputs[11067] = ~(layer1_outputs[2117]);
    assign layer2_outputs[11068] = ~(layer1_outputs[1307]);
    assign layer2_outputs[11069] = layer1_outputs[3363];
    assign layer2_outputs[11070] = ~((layer1_outputs[97]) & (layer1_outputs[4134]));
    assign layer2_outputs[11071] = (layer1_outputs[11155]) ^ (layer1_outputs[6160]);
    assign layer2_outputs[11072] = ~(layer1_outputs[4680]);
    assign layer2_outputs[11073] = ~(layer1_outputs[9233]) | (layer1_outputs[2665]);
    assign layer2_outputs[11074] = (layer1_outputs[7788]) ^ (layer1_outputs[7095]);
    assign layer2_outputs[11075] = layer1_outputs[663];
    assign layer2_outputs[11076] = (layer1_outputs[9000]) | (layer1_outputs[1578]);
    assign layer2_outputs[11077] = ~((layer1_outputs[8759]) & (layer1_outputs[7824]));
    assign layer2_outputs[11078] = ~(layer1_outputs[2201]);
    assign layer2_outputs[11079] = ~(layer1_outputs[9432]);
    assign layer2_outputs[11080] = (layer1_outputs[7607]) & ~(layer1_outputs[2494]);
    assign layer2_outputs[11081] = ~(layer1_outputs[918]);
    assign layer2_outputs[11082] = layer1_outputs[6206];
    assign layer2_outputs[11083] = ~((layer1_outputs[5490]) ^ (layer1_outputs[3844]));
    assign layer2_outputs[11084] = layer1_outputs[10649];
    assign layer2_outputs[11085] = (layer1_outputs[4909]) | (layer1_outputs[6923]);
    assign layer2_outputs[11086] = ~(layer1_outputs[8717]) | (layer1_outputs[11165]);
    assign layer2_outputs[11087] = ~((layer1_outputs[3520]) | (layer1_outputs[9042]));
    assign layer2_outputs[11088] = ~(layer1_outputs[11374]) | (layer1_outputs[3299]);
    assign layer2_outputs[11089] = layer1_outputs[1335];
    assign layer2_outputs[11090] = ~(layer1_outputs[10805]);
    assign layer2_outputs[11091] = ~((layer1_outputs[21]) & (layer1_outputs[7106]));
    assign layer2_outputs[11092] = ~(layer1_outputs[4532]);
    assign layer2_outputs[11093] = layer1_outputs[4530];
    assign layer2_outputs[11094] = (layer1_outputs[10798]) & ~(layer1_outputs[7965]);
    assign layer2_outputs[11095] = ~(layer1_outputs[5915]) | (layer1_outputs[10233]);
    assign layer2_outputs[11096] = (layer1_outputs[1729]) | (layer1_outputs[12738]);
    assign layer2_outputs[11097] = (layer1_outputs[9419]) & ~(layer1_outputs[7602]);
    assign layer2_outputs[11098] = layer1_outputs[6487];
    assign layer2_outputs[11099] = ~((layer1_outputs[1037]) ^ (layer1_outputs[2672]));
    assign layer2_outputs[11100] = ~(layer1_outputs[9763]);
    assign layer2_outputs[11101] = ~((layer1_outputs[7342]) | (layer1_outputs[11316]));
    assign layer2_outputs[11102] = layer1_outputs[1281];
    assign layer2_outputs[11103] = ~(layer1_outputs[4596]);
    assign layer2_outputs[11104] = ~(layer1_outputs[5357]);
    assign layer2_outputs[11105] = (layer1_outputs[10]) ^ (layer1_outputs[6557]);
    assign layer2_outputs[11106] = layer1_outputs[12444];
    assign layer2_outputs[11107] = ~(layer1_outputs[4987]);
    assign layer2_outputs[11108] = 1'b1;
    assign layer2_outputs[11109] = ~((layer1_outputs[11582]) | (layer1_outputs[3986]));
    assign layer2_outputs[11110] = layer1_outputs[6618];
    assign layer2_outputs[11111] = (layer1_outputs[1506]) ^ (layer1_outputs[11565]);
    assign layer2_outputs[11112] = (layer1_outputs[332]) & (layer1_outputs[6159]);
    assign layer2_outputs[11113] = ~(layer1_outputs[172]);
    assign layer2_outputs[11114] = (layer1_outputs[3236]) & ~(layer1_outputs[1911]);
    assign layer2_outputs[11115] = ~((layer1_outputs[8999]) & (layer1_outputs[8711]));
    assign layer2_outputs[11116] = (layer1_outputs[2802]) ^ (layer1_outputs[7319]);
    assign layer2_outputs[11117] = (layer1_outputs[2081]) & ~(layer1_outputs[9313]);
    assign layer2_outputs[11118] = ~((layer1_outputs[2232]) ^ (layer1_outputs[6073]));
    assign layer2_outputs[11119] = layer1_outputs[12596];
    assign layer2_outputs[11120] = ~((layer1_outputs[847]) ^ (layer1_outputs[1814]));
    assign layer2_outputs[11121] = layer1_outputs[9738];
    assign layer2_outputs[11122] = ~((layer1_outputs[6023]) ^ (layer1_outputs[2432]));
    assign layer2_outputs[11123] = ~(layer1_outputs[7480]) | (layer1_outputs[8757]);
    assign layer2_outputs[11124] = (layer1_outputs[11479]) ^ (layer1_outputs[10196]);
    assign layer2_outputs[11125] = (layer1_outputs[3922]) ^ (layer1_outputs[4423]);
    assign layer2_outputs[11126] = (layer1_outputs[11957]) & (layer1_outputs[1867]);
    assign layer2_outputs[11127] = ~((layer1_outputs[9434]) ^ (layer1_outputs[8247]));
    assign layer2_outputs[11128] = ~(layer1_outputs[2674]);
    assign layer2_outputs[11129] = layer1_outputs[6322];
    assign layer2_outputs[11130] = layer1_outputs[10019];
    assign layer2_outputs[11131] = (layer1_outputs[6935]) & ~(layer1_outputs[8997]);
    assign layer2_outputs[11132] = ~((layer1_outputs[11078]) ^ (layer1_outputs[5686]));
    assign layer2_outputs[11133] = layer1_outputs[6958];
    assign layer2_outputs[11134] = ~(layer1_outputs[12054]);
    assign layer2_outputs[11135] = layer1_outputs[5256];
    assign layer2_outputs[11136] = (layer1_outputs[10987]) ^ (layer1_outputs[9424]);
    assign layer2_outputs[11137] = ~(layer1_outputs[4012]);
    assign layer2_outputs[11138] = ~(layer1_outputs[9902]);
    assign layer2_outputs[11139] = layer1_outputs[1535];
    assign layer2_outputs[11140] = ~((layer1_outputs[6369]) | (layer1_outputs[3523]));
    assign layer2_outputs[11141] = ~(layer1_outputs[614]) | (layer1_outputs[1393]);
    assign layer2_outputs[11142] = layer1_outputs[1740];
    assign layer2_outputs[11143] = layer1_outputs[11094];
    assign layer2_outputs[11144] = (layer1_outputs[1289]) ^ (layer1_outputs[9945]);
    assign layer2_outputs[11145] = (layer1_outputs[9722]) & (layer1_outputs[3323]);
    assign layer2_outputs[11146] = ~(layer1_outputs[6059]) | (layer1_outputs[10958]);
    assign layer2_outputs[11147] = ~(layer1_outputs[10166]);
    assign layer2_outputs[11148] = ~((layer1_outputs[11605]) | (layer1_outputs[8499]));
    assign layer2_outputs[11149] = layer1_outputs[6273];
    assign layer2_outputs[11150] = layer1_outputs[1251];
    assign layer2_outputs[11151] = ~(layer1_outputs[377]);
    assign layer2_outputs[11152] = ~(layer1_outputs[7271]);
    assign layer2_outputs[11153] = layer1_outputs[12230];
    assign layer2_outputs[11154] = layer1_outputs[439];
    assign layer2_outputs[11155] = ~(layer1_outputs[5429]);
    assign layer2_outputs[11156] = ~(layer1_outputs[1241]);
    assign layer2_outputs[11157] = layer1_outputs[11919];
    assign layer2_outputs[11158] = (layer1_outputs[5608]) | (layer1_outputs[1445]);
    assign layer2_outputs[11159] = layer1_outputs[5433];
    assign layer2_outputs[11160] = ~(layer1_outputs[5871]) | (layer1_outputs[6088]);
    assign layer2_outputs[11161] = layer1_outputs[981];
    assign layer2_outputs[11162] = layer1_outputs[6040];
    assign layer2_outputs[11163] = (layer1_outputs[10610]) | (layer1_outputs[8678]);
    assign layer2_outputs[11164] = (layer1_outputs[7637]) ^ (layer1_outputs[7381]);
    assign layer2_outputs[11165] = layer1_outputs[4244];
    assign layer2_outputs[11166] = layer1_outputs[7601];
    assign layer2_outputs[11167] = layer1_outputs[9285];
    assign layer2_outputs[11168] = ~(layer1_outputs[31]);
    assign layer2_outputs[11169] = layer1_outputs[5131];
    assign layer2_outputs[11170] = layer1_outputs[12033];
    assign layer2_outputs[11171] = ~(layer1_outputs[12692]);
    assign layer2_outputs[11172] = (layer1_outputs[9858]) & ~(layer1_outputs[4605]);
    assign layer2_outputs[11173] = (layer1_outputs[5309]) ^ (layer1_outputs[84]);
    assign layer2_outputs[11174] = layer1_outputs[4689];
    assign layer2_outputs[11175] = (layer1_outputs[7257]) ^ (layer1_outputs[587]);
    assign layer2_outputs[11176] = layer1_outputs[9267];
    assign layer2_outputs[11177] = (layer1_outputs[6188]) | (layer1_outputs[6569]);
    assign layer2_outputs[11178] = layer1_outputs[6632];
    assign layer2_outputs[11179] = (layer1_outputs[5031]) & ~(layer1_outputs[4984]);
    assign layer2_outputs[11180] = ~((layer1_outputs[2094]) & (layer1_outputs[12691]));
    assign layer2_outputs[11181] = ~((layer1_outputs[9304]) ^ (layer1_outputs[7656]));
    assign layer2_outputs[11182] = ~(layer1_outputs[1981]);
    assign layer2_outputs[11183] = layer1_outputs[11832];
    assign layer2_outputs[11184] = ~(layer1_outputs[385]);
    assign layer2_outputs[11185] = ~((layer1_outputs[10445]) ^ (layer1_outputs[10631]));
    assign layer2_outputs[11186] = (layer1_outputs[5139]) & ~(layer1_outputs[11862]);
    assign layer2_outputs[11187] = ~(layer1_outputs[11521]) | (layer1_outputs[10520]);
    assign layer2_outputs[11188] = (layer1_outputs[10900]) & (layer1_outputs[3751]);
    assign layer2_outputs[11189] = layer1_outputs[4776];
    assign layer2_outputs[11190] = (layer1_outputs[7305]) & ~(layer1_outputs[920]);
    assign layer2_outputs[11191] = layer1_outputs[6231];
    assign layer2_outputs[11192] = (layer1_outputs[7831]) | (layer1_outputs[4241]);
    assign layer2_outputs[11193] = (layer1_outputs[767]) & ~(layer1_outputs[9397]);
    assign layer2_outputs[11194] = layer1_outputs[9663];
    assign layer2_outputs[11195] = 1'b1;
    assign layer2_outputs[11196] = (layer1_outputs[10521]) ^ (layer1_outputs[11955]);
    assign layer2_outputs[11197] = ~((layer1_outputs[11251]) ^ (layer1_outputs[8746]));
    assign layer2_outputs[11198] = (layer1_outputs[145]) ^ (layer1_outputs[3496]);
    assign layer2_outputs[11199] = (layer1_outputs[6711]) & (layer1_outputs[11492]);
    assign layer2_outputs[11200] = layer1_outputs[1499];
    assign layer2_outputs[11201] = ~((layer1_outputs[12536]) & (layer1_outputs[7866]));
    assign layer2_outputs[11202] = (layer1_outputs[11244]) & (layer1_outputs[8316]);
    assign layer2_outputs[11203] = (layer1_outputs[11822]) & ~(layer1_outputs[6849]);
    assign layer2_outputs[11204] = ~(layer1_outputs[5899]) | (layer1_outputs[2913]);
    assign layer2_outputs[11205] = ~((layer1_outputs[2144]) ^ (layer1_outputs[1905]));
    assign layer2_outputs[11206] = ~(layer1_outputs[47]);
    assign layer2_outputs[11207] = ~(layer1_outputs[6363]);
    assign layer2_outputs[11208] = ~(layer1_outputs[11909]);
    assign layer2_outputs[11209] = layer1_outputs[3256];
    assign layer2_outputs[11210] = ~(layer1_outputs[380]);
    assign layer2_outputs[11211] = layer1_outputs[8127];
    assign layer2_outputs[11212] = ~((layer1_outputs[9785]) | (layer1_outputs[12414]));
    assign layer2_outputs[11213] = ~((layer1_outputs[12133]) ^ (layer1_outputs[8659]));
    assign layer2_outputs[11214] = ~(layer1_outputs[9582]);
    assign layer2_outputs[11215] = ~(layer1_outputs[5096]) | (layer1_outputs[12289]);
    assign layer2_outputs[11216] = (layer1_outputs[2927]) & ~(layer1_outputs[2984]);
    assign layer2_outputs[11217] = ~((layer1_outputs[10669]) | (layer1_outputs[7183]));
    assign layer2_outputs[11218] = layer1_outputs[3037];
    assign layer2_outputs[11219] = (layer1_outputs[871]) & ~(layer1_outputs[4911]);
    assign layer2_outputs[11220] = (layer1_outputs[1706]) ^ (layer1_outputs[6012]);
    assign layer2_outputs[11221] = layer1_outputs[3704];
    assign layer2_outputs[11222] = ~(layer1_outputs[3901]);
    assign layer2_outputs[11223] = ~(layer1_outputs[10607]);
    assign layer2_outputs[11224] = (layer1_outputs[5035]) ^ (layer1_outputs[5044]);
    assign layer2_outputs[11225] = ~((layer1_outputs[1611]) | (layer1_outputs[12349]));
    assign layer2_outputs[11226] = layer1_outputs[560];
    assign layer2_outputs[11227] = ~((layer1_outputs[6482]) & (layer1_outputs[11059]));
    assign layer2_outputs[11228] = layer1_outputs[5887];
    assign layer2_outputs[11229] = layer1_outputs[5286];
    assign layer2_outputs[11230] = ~((layer1_outputs[177]) ^ (layer1_outputs[5058]));
    assign layer2_outputs[11231] = (layer1_outputs[11701]) & (layer1_outputs[12361]);
    assign layer2_outputs[11232] = ~((layer1_outputs[2328]) | (layer1_outputs[9912]));
    assign layer2_outputs[11233] = ~(layer1_outputs[4056]);
    assign layer2_outputs[11234] = ~(layer1_outputs[1068]);
    assign layer2_outputs[11235] = ~(layer1_outputs[4726]) | (layer1_outputs[10406]);
    assign layer2_outputs[11236] = (layer1_outputs[9658]) ^ (layer1_outputs[2160]);
    assign layer2_outputs[11237] = ~(layer1_outputs[11079]);
    assign layer2_outputs[11238] = layer1_outputs[12736];
    assign layer2_outputs[11239] = ~((layer1_outputs[10818]) & (layer1_outputs[3350]));
    assign layer2_outputs[11240] = layer1_outputs[11227];
    assign layer2_outputs[11241] = ~(layer1_outputs[7739]);
    assign layer2_outputs[11242] = (layer1_outputs[8087]) ^ (layer1_outputs[10673]);
    assign layer2_outputs[11243] = (layer1_outputs[3235]) & ~(layer1_outputs[106]);
    assign layer2_outputs[11244] = (layer1_outputs[1226]) & ~(layer1_outputs[3737]);
    assign layer2_outputs[11245] = (layer1_outputs[7193]) & ~(layer1_outputs[7625]);
    assign layer2_outputs[11246] = ~(layer1_outputs[7978]) | (layer1_outputs[988]);
    assign layer2_outputs[11247] = ~(layer1_outputs[613]) | (layer1_outputs[8567]);
    assign layer2_outputs[11248] = ~((layer1_outputs[5405]) ^ (layer1_outputs[9156]));
    assign layer2_outputs[11249] = layer1_outputs[11792];
    assign layer2_outputs[11250] = (layer1_outputs[3367]) | (layer1_outputs[7274]);
    assign layer2_outputs[11251] = layer1_outputs[2766];
    assign layer2_outputs[11252] = ~(layer1_outputs[8276]);
    assign layer2_outputs[11253] = ~(layer1_outputs[4580]);
    assign layer2_outputs[11254] = ~(layer1_outputs[2731]);
    assign layer2_outputs[11255] = (layer1_outputs[1626]) & (layer1_outputs[2692]);
    assign layer2_outputs[11256] = layer1_outputs[9339];
    assign layer2_outputs[11257] = layer1_outputs[3004];
    assign layer2_outputs[11258] = ~(layer1_outputs[8293]) | (layer1_outputs[6345]);
    assign layer2_outputs[11259] = (layer1_outputs[7301]) | (layer1_outputs[11364]);
    assign layer2_outputs[11260] = (layer1_outputs[9182]) | (layer1_outputs[11744]);
    assign layer2_outputs[11261] = (layer1_outputs[11535]) & (layer1_outputs[10455]);
    assign layer2_outputs[11262] = ~(layer1_outputs[1733]);
    assign layer2_outputs[11263] = ~((layer1_outputs[1034]) | (layer1_outputs[4016]));
    assign layer2_outputs[11264] = layer1_outputs[11522];
    assign layer2_outputs[11265] = layer1_outputs[3311];
    assign layer2_outputs[11266] = layer1_outputs[2402];
    assign layer2_outputs[11267] = ~(layer1_outputs[5132]);
    assign layer2_outputs[11268] = ~((layer1_outputs[8838]) | (layer1_outputs[1975]));
    assign layer2_outputs[11269] = ~(layer1_outputs[11990]) | (layer1_outputs[11301]);
    assign layer2_outputs[11270] = (layer1_outputs[9046]) & (layer1_outputs[12010]);
    assign layer2_outputs[11271] = layer1_outputs[8540];
    assign layer2_outputs[11272] = layer1_outputs[9878];
    assign layer2_outputs[11273] = 1'b0;
    assign layer2_outputs[11274] = layer1_outputs[12718];
    assign layer2_outputs[11275] = (layer1_outputs[2993]) | (layer1_outputs[9834]);
    assign layer2_outputs[11276] = ~((layer1_outputs[11272]) ^ (layer1_outputs[754]));
    assign layer2_outputs[11277] = ~((layer1_outputs[12254]) ^ (layer1_outputs[6921]));
    assign layer2_outputs[11278] = (layer1_outputs[9616]) & (layer1_outputs[6517]);
    assign layer2_outputs[11279] = layer1_outputs[6212];
    assign layer2_outputs[11280] = ~(layer1_outputs[9282]);
    assign layer2_outputs[11281] = layer1_outputs[5951];
    assign layer2_outputs[11282] = ~((layer1_outputs[10908]) ^ (layer1_outputs[3089]));
    assign layer2_outputs[11283] = (layer1_outputs[346]) & ~(layer1_outputs[9266]);
    assign layer2_outputs[11284] = ~((layer1_outputs[7848]) ^ (layer1_outputs[1317]));
    assign layer2_outputs[11285] = ~(layer1_outputs[5527]);
    assign layer2_outputs[11286] = ~((layer1_outputs[12354]) ^ (layer1_outputs[11008]));
    assign layer2_outputs[11287] = (layer1_outputs[9569]) | (layer1_outputs[10774]);
    assign layer2_outputs[11288] = ~((layer1_outputs[5111]) ^ (layer1_outputs[2111]));
    assign layer2_outputs[11289] = ~(layer1_outputs[2998]);
    assign layer2_outputs[11290] = ~(layer1_outputs[11349]);
    assign layer2_outputs[11291] = layer1_outputs[2007];
    assign layer2_outputs[11292] = (layer1_outputs[2072]) & ~(layer1_outputs[10329]);
    assign layer2_outputs[11293] = ~(layer1_outputs[7522]);
    assign layer2_outputs[11294] = ~(layer1_outputs[5943]);
    assign layer2_outputs[11295] = ~(layer1_outputs[6309]);
    assign layer2_outputs[11296] = (layer1_outputs[7946]) ^ (layer1_outputs[4156]);
    assign layer2_outputs[11297] = (layer1_outputs[12735]) & (layer1_outputs[11654]);
    assign layer2_outputs[11298] = ~(layer1_outputs[6551]);
    assign layer2_outputs[11299] = ~(layer1_outputs[12249]);
    assign layer2_outputs[11300] = layer1_outputs[3238];
    assign layer2_outputs[11301] = ~(layer1_outputs[6864]);
    assign layer2_outputs[11302] = ~(layer1_outputs[12479]);
    assign layer2_outputs[11303] = ~(layer1_outputs[6826]) | (layer1_outputs[10667]);
    assign layer2_outputs[11304] = ~((layer1_outputs[8433]) | (layer1_outputs[1672]));
    assign layer2_outputs[11305] = ~((layer1_outputs[8330]) | (layer1_outputs[12032]));
    assign layer2_outputs[11306] = (layer1_outputs[12454]) & (layer1_outputs[6337]);
    assign layer2_outputs[11307] = layer1_outputs[3879];
    assign layer2_outputs[11308] = ~((layer1_outputs[1361]) & (layer1_outputs[9543]));
    assign layer2_outputs[11309] = ~(layer1_outputs[11657]);
    assign layer2_outputs[11310] = layer1_outputs[6247];
    assign layer2_outputs[11311] = ~((layer1_outputs[5458]) ^ (layer1_outputs[11448]));
    assign layer2_outputs[11312] = ~(layer1_outputs[7044]);
    assign layer2_outputs[11313] = layer1_outputs[6743];
    assign layer2_outputs[11314] = (layer1_outputs[5531]) & ~(layer1_outputs[2294]);
    assign layer2_outputs[11315] = (layer1_outputs[7747]) ^ (layer1_outputs[12379]);
    assign layer2_outputs[11316] = (layer1_outputs[2310]) ^ (layer1_outputs[8580]);
    assign layer2_outputs[11317] = ~(layer1_outputs[11684]) | (layer1_outputs[4621]);
    assign layer2_outputs[11318] = (layer1_outputs[1897]) ^ (layer1_outputs[9793]);
    assign layer2_outputs[11319] = layer1_outputs[6049];
    assign layer2_outputs[11320] = 1'b1;
    assign layer2_outputs[11321] = layer1_outputs[5491];
    assign layer2_outputs[11322] = ~(layer1_outputs[5469]);
    assign layer2_outputs[11323] = (layer1_outputs[9768]) | (layer1_outputs[1]);
    assign layer2_outputs[11324] = ~(layer1_outputs[5992]);
    assign layer2_outputs[11325] = layer1_outputs[8509];
    assign layer2_outputs[11326] = (layer1_outputs[6619]) & ~(layer1_outputs[4367]);
    assign layer2_outputs[11327] = layer1_outputs[5310];
    assign layer2_outputs[11328] = ~(layer1_outputs[9429]);
    assign layer2_outputs[11329] = ~(layer1_outputs[4915]);
    assign layer2_outputs[11330] = (layer1_outputs[7749]) | (layer1_outputs[5000]);
    assign layer2_outputs[11331] = ~(layer1_outputs[6197]);
    assign layer2_outputs[11332] = ~(layer1_outputs[11724]);
    assign layer2_outputs[11333] = ~(layer1_outputs[6655]);
    assign layer2_outputs[11334] = layer1_outputs[3878];
    assign layer2_outputs[11335] = ~(layer1_outputs[12632]);
    assign layer2_outputs[11336] = (layer1_outputs[9555]) | (layer1_outputs[6903]);
    assign layer2_outputs[11337] = ~(layer1_outputs[147]);
    assign layer2_outputs[11338] = ~((layer1_outputs[1757]) ^ (layer1_outputs[6316]));
    assign layer2_outputs[11339] = layer1_outputs[12259];
    assign layer2_outputs[11340] = ~((layer1_outputs[5719]) ^ (layer1_outputs[6065]));
    assign layer2_outputs[11341] = ~(layer1_outputs[12129]);
    assign layer2_outputs[11342] = (layer1_outputs[3519]) ^ (layer1_outputs[5810]);
    assign layer2_outputs[11343] = layer1_outputs[12157];
    assign layer2_outputs[11344] = ~(layer1_outputs[4208]);
    assign layer2_outputs[11345] = ~(layer1_outputs[3960]) | (layer1_outputs[11906]);
    assign layer2_outputs[11346] = ~((layer1_outputs[4905]) ^ (layer1_outputs[3584]));
    assign layer2_outputs[11347] = ~(layer1_outputs[8179]);
    assign layer2_outputs[11348] = layer1_outputs[2882];
    assign layer2_outputs[11349] = ~(layer1_outputs[3496]);
    assign layer2_outputs[11350] = layer1_outputs[3679];
    assign layer2_outputs[11351] = ~((layer1_outputs[1378]) | (layer1_outputs[4223]));
    assign layer2_outputs[11352] = layer1_outputs[5451];
    assign layer2_outputs[11353] = ~((layer1_outputs[10814]) & (layer1_outputs[531]));
    assign layer2_outputs[11354] = layer1_outputs[10024];
    assign layer2_outputs[11355] = ~(layer1_outputs[4175]);
    assign layer2_outputs[11356] = (layer1_outputs[3199]) | (layer1_outputs[10557]);
    assign layer2_outputs[11357] = (layer1_outputs[1695]) & ~(layer1_outputs[9935]);
    assign layer2_outputs[11358] = ~(layer1_outputs[2546]);
    assign layer2_outputs[11359] = (layer1_outputs[1293]) | (layer1_outputs[2282]);
    assign layer2_outputs[11360] = layer1_outputs[12103];
    assign layer2_outputs[11361] = ~((layer1_outputs[11796]) | (layer1_outputs[2820]));
    assign layer2_outputs[11362] = ~(layer1_outputs[12355]) | (layer1_outputs[1851]);
    assign layer2_outputs[11363] = ~((layer1_outputs[2323]) ^ (layer1_outputs[11761]));
    assign layer2_outputs[11364] = ~(layer1_outputs[2017]);
    assign layer2_outputs[11365] = ~((layer1_outputs[4187]) | (layer1_outputs[5662]));
    assign layer2_outputs[11366] = layer1_outputs[8062];
    assign layer2_outputs[11367] = ~(layer1_outputs[1275]) | (layer1_outputs[11313]);
    assign layer2_outputs[11368] = layer1_outputs[9098];
    assign layer2_outputs[11369] = (layer1_outputs[12465]) & (layer1_outputs[9177]);
    assign layer2_outputs[11370] = ~(layer1_outputs[1598]);
    assign layer2_outputs[11371] = ~((layer1_outputs[2357]) & (layer1_outputs[6315]));
    assign layer2_outputs[11372] = (layer1_outputs[10472]) & ~(layer1_outputs[6531]);
    assign layer2_outputs[11373] = layer1_outputs[8917];
    assign layer2_outputs[11374] = ~(layer1_outputs[9230]);
    assign layer2_outputs[11375] = ~(layer1_outputs[3562]);
    assign layer2_outputs[11376] = ~(layer1_outputs[3201]);
    assign layer2_outputs[11377] = (layer1_outputs[10121]) & (layer1_outputs[10231]);
    assign layer2_outputs[11378] = ~(layer1_outputs[10536]);
    assign layer2_outputs[11379] = layer1_outputs[8076];
    assign layer2_outputs[11380] = (layer1_outputs[2543]) & ~(layer1_outputs[11349]);
    assign layer2_outputs[11381] = ~(layer1_outputs[5714]) | (layer1_outputs[4134]);
    assign layer2_outputs[11382] = (layer1_outputs[7131]) & (layer1_outputs[8669]);
    assign layer2_outputs[11383] = layer1_outputs[11019];
    assign layer2_outputs[11384] = (layer1_outputs[3029]) ^ (layer1_outputs[11438]);
    assign layer2_outputs[11385] = ~(layer1_outputs[1790]);
    assign layer2_outputs[11386] = ~(layer1_outputs[611]);
    assign layer2_outputs[11387] = layer1_outputs[3680];
    assign layer2_outputs[11388] = ~(layer1_outputs[11645]) | (layer1_outputs[9607]);
    assign layer2_outputs[11389] = layer1_outputs[6545];
    assign layer2_outputs[11390] = (layer1_outputs[7822]) & (layer1_outputs[3285]);
    assign layer2_outputs[11391] = (layer1_outputs[2809]) & ~(layer1_outputs[4553]);
    assign layer2_outputs[11392] = ~(layer1_outputs[6290]);
    assign layer2_outputs[11393] = (layer1_outputs[11467]) & ~(layer1_outputs[11714]);
    assign layer2_outputs[11394] = (layer1_outputs[2010]) & ~(layer1_outputs[5833]);
    assign layer2_outputs[11395] = (layer1_outputs[12768]) ^ (layer1_outputs[5094]);
    assign layer2_outputs[11396] = layer1_outputs[324];
    assign layer2_outputs[11397] = ~((layer1_outputs[10654]) & (layer1_outputs[12121]));
    assign layer2_outputs[11398] = layer1_outputs[9376];
    assign layer2_outputs[11399] = (layer1_outputs[8652]) ^ (layer1_outputs[11012]);
    assign layer2_outputs[11400] = ~((layer1_outputs[10952]) | (layer1_outputs[11090]));
    assign layer2_outputs[11401] = ~(layer1_outputs[8399]);
    assign layer2_outputs[11402] = layer1_outputs[6709];
    assign layer2_outputs[11403] = layer1_outputs[9723];
    assign layer2_outputs[11404] = ~(layer1_outputs[9704]);
    assign layer2_outputs[11405] = ~((layer1_outputs[12482]) | (layer1_outputs[8166]));
    assign layer2_outputs[11406] = ~(layer1_outputs[2729]);
    assign layer2_outputs[11407] = layer1_outputs[3102];
    assign layer2_outputs[11408] = ~((layer1_outputs[10121]) ^ (layer1_outputs[10346]));
    assign layer2_outputs[11409] = (layer1_outputs[10365]) | (layer1_outputs[11982]);
    assign layer2_outputs[11410] = ~(layer1_outputs[1321]);
    assign layer2_outputs[11411] = ~((layer1_outputs[990]) | (layer1_outputs[1109]));
    assign layer2_outputs[11412] = (layer1_outputs[1103]) & ~(layer1_outputs[375]);
    assign layer2_outputs[11413] = (layer1_outputs[12351]) & ~(layer1_outputs[12464]);
    assign layer2_outputs[11414] = (layer1_outputs[1104]) ^ (layer1_outputs[556]);
    assign layer2_outputs[11415] = ~((layer1_outputs[2501]) | (layer1_outputs[10590]));
    assign layer2_outputs[11416] = ~((layer1_outputs[8297]) | (layer1_outputs[7340]));
    assign layer2_outputs[11417] = ~(layer1_outputs[10351]);
    assign layer2_outputs[11418] = (layer1_outputs[3796]) ^ (layer1_outputs[2627]);
    assign layer2_outputs[11419] = 1'b1;
    assign layer2_outputs[11420] = (layer1_outputs[5342]) & (layer1_outputs[12117]);
    assign layer2_outputs[11421] = ~(layer1_outputs[9901]) | (layer1_outputs[2314]);
    assign layer2_outputs[11422] = ~(layer1_outputs[10429]);
    assign layer2_outputs[11423] = ~(layer1_outputs[678]);
    assign layer2_outputs[11424] = ~(layer1_outputs[7577]);
    assign layer2_outputs[11425] = ~(layer1_outputs[1522]) | (layer1_outputs[6774]);
    assign layer2_outputs[11426] = layer1_outputs[4481];
    assign layer2_outputs[11427] = (layer1_outputs[3406]) & ~(layer1_outputs[6774]);
    assign layer2_outputs[11428] = ~(layer1_outputs[12503]);
    assign layer2_outputs[11429] = ~((layer1_outputs[906]) | (layer1_outputs[360]));
    assign layer2_outputs[11430] = (layer1_outputs[8873]) & ~(layer1_outputs[6844]);
    assign layer2_outputs[11431] = (layer1_outputs[12765]) ^ (layer1_outputs[3076]);
    assign layer2_outputs[11432] = ~(layer1_outputs[10047]) | (layer1_outputs[8021]);
    assign layer2_outputs[11433] = ~(layer1_outputs[11134]);
    assign layer2_outputs[11434] = layer1_outputs[5344];
    assign layer2_outputs[11435] = ~(layer1_outputs[1593]);
    assign layer2_outputs[11436] = (layer1_outputs[10376]) & (layer1_outputs[11797]);
    assign layer2_outputs[11437] = (layer1_outputs[4484]) & ~(layer1_outputs[8310]);
    assign layer2_outputs[11438] = (layer1_outputs[5263]) ^ (layer1_outputs[7785]);
    assign layer2_outputs[11439] = 1'b0;
    assign layer2_outputs[11440] = (layer1_outputs[10295]) ^ (layer1_outputs[8926]);
    assign layer2_outputs[11441] = (layer1_outputs[12774]) | (layer1_outputs[10676]);
    assign layer2_outputs[11442] = ~(layer1_outputs[2568]);
    assign layer2_outputs[11443] = ~(layer1_outputs[1857]);
    assign layer2_outputs[11444] = ~(layer1_outputs[11289]);
    assign layer2_outputs[11445] = ~(layer1_outputs[6132]);
    assign layer2_outputs[11446] = ~((layer1_outputs[2320]) ^ (layer1_outputs[6312]));
    assign layer2_outputs[11447] = layer1_outputs[4537];
    assign layer2_outputs[11448] = layer1_outputs[5968];
    assign layer2_outputs[11449] = layer1_outputs[5249];
    assign layer2_outputs[11450] = ~((layer1_outputs[8147]) | (layer1_outputs[9519]));
    assign layer2_outputs[11451] = layer1_outputs[11176];
    assign layer2_outputs[11452] = layer1_outputs[3811];
    assign layer2_outputs[11453] = (layer1_outputs[310]) | (layer1_outputs[7712]);
    assign layer2_outputs[11454] = layer1_outputs[9995];
    assign layer2_outputs[11455] = ~((layer1_outputs[3776]) | (layer1_outputs[1284]));
    assign layer2_outputs[11456] = ~(layer1_outputs[7116]);
    assign layer2_outputs[11457] = layer1_outputs[832];
    assign layer2_outputs[11458] = ~(layer1_outputs[298]);
    assign layer2_outputs[11459] = ~(layer1_outputs[3732]);
    assign layer2_outputs[11460] = ~(layer1_outputs[12274]);
    assign layer2_outputs[11461] = ~(layer1_outputs[5577]);
    assign layer2_outputs[11462] = layer1_outputs[6575];
    assign layer2_outputs[11463] = layer1_outputs[8021];
    assign layer2_outputs[11464] = ~((layer1_outputs[128]) & (layer1_outputs[12632]));
    assign layer2_outputs[11465] = (layer1_outputs[848]) ^ (layer1_outputs[54]);
    assign layer2_outputs[11466] = ~(layer1_outputs[8279]);
    assign layer2_outputs[11467] = ~(layer1_outputs[518]) | (layer1_outputs[10533]);
    assign layer2_outputs[11468] = layer1_outputs[1305];
    assign layer2_outputs[11469] = ~(layer1_outputs[16]);
    assign layer2_outputs[11470] = (layer1_outputs[4493]) & ~(layer1_outputs[2361]);
    assign layer2_outputs[11471] = ~(layer1_outputs[3349]);
    assign layer2_outputs[11472] = ~((layer1_outputs[7523]) | (layer1_outputs[4311]));
    assign layer2_outputs[11473] = layer1_outputs[4627];
    assign layer2_outputs[11474] = ~(layer1_outputs[2041]);
    assign layer2_outputs[11475] = ~((layer1_outputs[10106]) | (layer1_outputs[3823]));
    assign layer2_outputs[11476] = ~(layer1_outputs[1992]);
    assign layer2_outputs[11477] = ~((layer1_outputs[6719]) | (layer1_outputs[5958]));
    assign layer2_outputs[11478] = ~(layer1_outputs[5074]);
    assign layer2_outputs[11479] = ~(layer1_outputs[6935]);
    assign layer2_outputs[11480] = ~(layer1_outputs[12255]);
    assign layer2_outputs[11481] = layer1_outputs[10614];
    assign layer2_outputs[11482] = ~(layer1_outputs[4891]);
    assign layer2_outputs[11483] = ~((layer1_outputs[6598]) | (layer1_outputs[5141]));
    assign layer2_outputs[11484] = layer1_outputs[10594];
    assign layer2_outputs[11485] = ~((layer1_outputs[5768]) & (layer1_outputs[8726]));
    assign layer2_outputs[11486] = layer1_outputs[7179];
    assign layer2_outputs[11487] = ~(layer1_outputs[5197]) | (layer1_outputs[11574]);
    assign layer2_outputs[11488] = ~(layer1_outputs[9251]);
    assign layer2_outputs[11489] = ~(layer1_outputs[12715]);
    assign layer2_outputs[11490] = ~(layer1_outputs[264]);
    assign layer2_outputs[11491] = (layer1_outputs[6483]) & ~(layer1_outputs[4007]);
    assign layer2_outputs[11492] = layer1_outputs[7864];
    assign layer2_outputs[11493] = (layer1_outputs[1107]) & ~(layer1_outputs[8947]);
    assign layer2_outputs[11494] = layer1_outputs[12278];
    assign layer2_outputs[11495] = (layer1_outputs[8303]) & ~(layer1_outputs[363]);
    assign layer2_outputs[11496] = ~(layer1_outputs[8647]);
    assign layer2_outputs[11497] = layer1_outputs[3057];
    assign layer2_outputs[11498] = ~(layer1_outputs[4363]);
    assign layer2_outputs[11499] = layer1_outputs[7461];
    assign layer2_outputs[11500] = layer1_outputs[858];
    assign layer2_outputs[11501] = ~(layer1_outputs[2544]);
    assign layer2_outputs[11502] = layer1_outputs[2363];
    assign layer2_outputs[11503] = ~((layer1_outputs[3281]) | (layer1_outputs[11354]));
    assign layer2_outputs[11504] = layer1_outputs[8144];
    assign layer2_outputs[11505] = layer1_outputs[11058];
    assign layer2_outputs[11506] = (layer1_outputs[10820]) | (layer1_outputs[7767]);
    assign layer2_outputs[11507] = (layer1_outputs[10243]) ^ (layer1_outputs[4630]);
    assign layer2_outputs[11508] = ~(layer1_outputs[7414]);
    assign layer2_outputs[11509] = ~((layer1_outputs[7377]) & (layer1_outputs[9686]));
    assign layer2_outputs[11510] = ~(layer1_outputs[6234]);
    assign layer2_outputs[11511] = layer1_outputs[2251];
    assign layer2_outputs[11512] = ~((layer1_outputs[7937]) & (layer1_outputs[7462]));
    assign layer2_outputs[11513] = (layer1_outputs[1033]) | (layer1_outputs[1408]);
    assign layer2_outputs[11514] = (layer1_outputs[700]) ^ (layer1_outputs[9193]);
    assign layer2_outputs[11515] = layer1_outputs[3446];
    assign layer2_outputs[11516] = (layer1_outputs[8014]) ^ (layer1_outputs[2242]);
    assign layer2_outputs[11517] = layer1_outputs[11114];
    assign layer2_outputs[11518] = (layer1_outputs[5173]) ^ (layer1_outputs[6385]);
    assign layer2_outputs[11519] = layer1_outputs[2909];
    assign layer2_outputs[11520] = ~(layer1_outputs[6403]);
    assign layer2_outputs[11521] = (layer1_outputs[7170]) & (layer1_outputs[7298]);
    assign layer2_outputs[11522] = ~((layer1_outputs[2242]) ^ (layer1_outputs[302]));
    assign layer2_outputs[11523] = layer1_outputs[5861];
    assign layer2_outputs[11524] = ~((layer1_outputs[8614]) & (layer1_outputs[8196]));
    assign layer2_outputs[11525] = ~((layer1_outputs[4443]) | (layer1_outputs[6037]));
    assign layer2_outputs[11526] = ~((layer1_outputs[9341]) ^ (layer1_outputs[12343]));
    assign layer2_outputs[11527] = layer1_outputs[4957];
    assign layer2_outputs[11528] = layer1_outputs[11859];
    assign layer2_outputs[11529] = layer1_outputs[1340];
    assign layer2_outputs[11530] = layer1_outputs[1389];
    assign layer2_outputs[11531] = ~(layer1_outputs[7050]) | (layer1_outputs[4893]);
    assign layer2_outputs[11532] = ~(layer1_outputs[6349]);
    assign layer2_outputs[11533] = ~(layer1_outputs[4223]);
    assign layer2_outputs[11534] = layer1_outputs[328];
    assign layer2_outputs[11535] = layer1_outputs[7876];
    assign layer2_outputs[11536] = (layer1_outputs[5242]) ^ (layer1_outputs[8535]);
    assign layer2_outputs[11537] = ~((layer1_outputs[1380]) & (layer1_outputs[7643]));
    assign layer2_outputs[11538] = (layer1_outputs[4976]) & ~(layer1_outputs[2425]);
    assign layer2_outputs[11539] = ~(layer1_outputs[269]) | (layer1_outputs[7155]);
    assign layer2_outputs[11540] = (layer1_outputs[10091]) | (layer1_outputs[11135]);
    assign layer2_outputs[11541] = ~(layer1_outputs[5066]);
    assign layer2_outputs[11542] = (layer1_outputs[7421]) ^ (layer1_outputs[2463]);
    assign layer2_outputs[11543] = ~(layer1_outputs[11080]);
    assign layer2_outputs[11544] = layer1_outputs[4233];
    assign layer2_outputs[11545] = ~((layer1_outputs[1572]) | (layer1_outputs[1023]));
    assign layer2_outputs[11546] = ~(layer1_outputs[12268]);
    assign layer2_outputs[11547] = layer1_outputs[3821];
    assign layer2_outputs[11548] = layer1_outputs[7363];
    assign layer2_outputs[11549] = (layer1_outputs[6779]) & ~(layer1_outputs[1174]);
    assign layer2_outputs[11550] = (layer1_outputs[8340]) ^ (layer1_outputs[5082]);
    assign layer2_outputs[11551] = layer1_outputs[2517];
    assign layer2_outputs[11552] = ~((layer1_outputs[4675]) ^ (layer1_outputs[11753]));
    assign layer2_outputs[11553] = (layer1_outputs[743]) & (layer1_outputs[1857]);
    assign layer2_outputs[11554] = (layer1_outputs[6374]) & ~(layer1_outputs[1161]);
    assign layer2_outputs[11555] = ~((layer1_outputs[10916]) & (layer1_outputs[3598]));
    assign layer2_outputs[11556] = ~(layer1_outputs[9959]);
    assign layer2_outputs[11557] = layer1_outputs[727];
    assign layer2_outputs[11558] = ~(layer1_outputs[4569]) | (layer1_outputs[285]);
    assign layer2_outputs[11559] = ~(layer1_outputs[528]) | (layer1_outputs[4961]);
    assign layer2_outputs[11560] = ~((layer1_outputs[6290]) | (layer1_outputs[10486]));
    assign layer2_outputs[11561] = (layer1_outputs[12302]) & (layer1_outputs[11059]);
    assign layer2_outputs[11562] = layer1_outputs[8081];
    assign layer2_outputs[11563] = ~((layer1_outputs[324]) & (layer1_outputs[9983]));
    assign layer2_outputs[11564] = ~((layer1_outputs[9533]) ^ (layer1_outputs[5477]));
    assign layer2_outputs[11565] = layer1_outputs[11088];
    assign layer2_outputs[11566] = ~(layer1_outputs[964]) | (layer1_outputs[10032]);
    assign layer2_outputs[11567] = (layer1_outputs[9349]) & ~(layer1_outputs[451]);
    assign layer2_outputs[11568] = ~((layer1_outputs[1063]) ^ (layer1_outputs[477]));
    assign layer2_outputs[11569] = ~(layer1_outputs[2878]);
    assign layer2_outputs[11570] = (layer1_outputs[3030]) & ~(layer1_outputs[7190]);
    assign layer2_outputs[11571] = (layer1_outputs[9330]) & ~(layer1_outputs[12566]);
    assign layer2_outputs[11572] = ~(layer1_outputs[8701]);
    assign layer2_outputs[11573] = (layer1_outputs[5975]) & (layer1_outputs[6962]);
    assign layer2_outputs[11574] = ~(layer1_outputs[10545]) | (layer1_outputs[5841]);
    assign layer2_outputs[11575] = ~(layer1_outputs[10749]);
    assign layer2_outputs[11576] = layer1_outputs[3396];
    assign layer2_outputs[11577] = (layer1_outputs[5323]) & (layer1_outputs[1577]);
    assign layer2_outputs[11578] = ~(layer1_outputs[1571]);
    assign layer2_outputs[11579] = (layer1_outputs[12347]) ^ (layer1_outputs[4344]);
    assign layer2_outputs[11580] = ~(layer1_outputs[8156]) | (layer1_outputs[7427]);
    assign layer2_outputs[11581] = (layer1_outputs[4538]) ^ (layer1_outputs[9707]);
    assign layer2_outputs[11582] = ~(layer1_outputs[1969]);
    assign layer2_outputs[11583] = ~(layer1_outputs[10090]);
    assign layer2_outputs[11584] = ~((layer1_outputs[10363]) | (layer1_outputs[1540]));
    assign layer2_outputs[11585] = layer1_outputs[5464];
    assign layer2_outputs[11586] = layer1_outputs[10902];
    assign layer2_outputs[11587] = ~(layer1_outputs[9601]);
    assign layer2_outputs[11588] = layer1_outputs[7251];
    assign layer2_outputs[11589] = ~(layer1_outputs[1412]);
    assign layer2_outputs[11590] = layer1_outputs[1078];
    assign layer2_outputs[11591] = (layer1_outputs[9943]) & ~(layer1_outputs[11270]);
    assign layer2_outputs[11592] = layer1_outputs[6488];
    assign layer2_outputs[11593] = (layer1_outputs[12059]) ^ (layer1_outputs[4389]);
    assign layer2_outputs[11594] = ~(layer1_outputs[2710]) | (layer1_outputs[747]);
    assign layer2_outputs[11595] = layer1_outputs[1576];
    assign layer2_outputs[11596] = layer1_outputs[9146];
    assign layer2_outputs[11597] = ~(layer1_outputs[10771]);
    assign layer2_outputs[11598] = layer1_outputs[1310];
    assign layer2_outputs[11599] = ~(layer1_outputs[3530]);
    assign layer2_outputs[11600] = (layer1_outputs[7607]) ^ (layer1_outputs[10036]);
    assign layer2_outputs[11601] = layer1_outputs[12500];
    assign layer2_outputs[11602] = ~(layer1_outputs[5944]);
    assign layer2_outputs[11603] = ~(layer1_outputs[3548]);
    assign layer2_outputs[11604] = layer1_outputs[9149];
    assign layer2_outputs[11605] = layer1_outputs[12511];
    assign layer2_outputs[11606] = ~(layer1_outputs[11979]);
    assign layer2_outputs[11607] = (layer1_outputs[6255]) & ~(layer1_outputs[8400]);
    assign layer2_outputs[11608] = layer1_outputs[10098];
    assign layer2_outputs[11609] = layer1_outputs[11482];
    assign layer2_outputs[11610] = layer1_outputs[6102];
    assign layer2_outputs[11611] = ~(layer1_outputs[9806]);
    assign layer2_outputs[11612] = ~(layer1_outputs[2943]) | (layer1_outputs[5829]);
    assign layer2_outputs[11613] = layer1_outputs[1937];
    assign layer2_outputs[11614] = ~(layer1_outputs[3231]);
    assign layer2_outputs[11615] = (layer1_outputs[11685]) & ~(layer1_outputs[4763]);
    assign layer2_outputs[11616] = layer1_outputs[11885];
    assign layer2_outputs[11617] = ~(layer1_outputs[10906]) | (layer1_outputs[7926]);
    assign layer2_outputs[11618] = (layer1_outputs[2607]) & ~(layer1_outputs[4852]);
    assign layer2_outputs[11619] = ~(layer1_outputs[3461]);
    assign layer2_outputs[11620] = (layer1_outputs[10174]) ^ (layer1_outputs[10283]);
    assign layer2_outputs[11621] = layer1_outputs[11932];
    assign layer2_outputs[11622] = ~((layer1_outputs[943]) ^ (layer1_outputs[3609]));
    assign layer2_outputs[11623] = layer1_outputs[3900];
    assign layer2_outputs[11624] = layer1_outputs[11280];
    assign layer2_outputs[11625] = (layer1_outputs[1017]) & (layer1_outputs[11725]);
    assign layer2_outputs[11626] = ~(layer1_outputs[2515]);
    assign layer2_outputs[11627] = (layer1_outputs[9568]) & (layer1_outputs[1563]);
    assign layer2_outputs[11628] = (layer1_outputs[3057]) ^ (layer1_outputs[2056]);
    assign layer2_outputs[11629] = ~((layer1_outputs[10883]) ^ (layer1_outputs[9370]));
    assign layer2_outputs[11630] = layer1_outputs[1211];
    assign layer2_outputs[11631] = layer1_outputs[9139];
    assign layer2_outputs[11632] = layer1_outputs[7611];
    assign layer2_outputs[11633] = ~(layer1_outputs[1772]);
    assign layer2_outputs[11634] = layer1_outputs[12594];
    assign layer2_outputs[11635] = (layer1_outputs[4281]) | (layer1_outputs[10887]);
    assign layer2_outputs[11636] = layer1_outputs[597];
    assign layer2_outputs[11637] = ~(layer1_outputs[11613]);
    assign layer2_outputs[11638] = (layer1_outputs[5488]) ^ (layer1_outputs[8181]);
    assign layer2_outputs[11639] = layer1_outputs[10384];
    assign layer2_outputs[11640] = (layer1_outputs[4485]) & ~(layer1_outputs[4499]);
    assign layer2_outputs[11641] = (layer1_outputs[344]) ^ (layer1_outputs[715]);
    assign layer2_outputs[11642] = layer1_outputs[12253];
    assign layer2_outputs[11643] = layer1_outputs[6973];
    assign layer2_outputs[11644] = layer1_outputs[5145];
    assign layer2_outputs[11645] = ~(layer1_outputs[7806]);
    assign layer2_outputs[11646] = layer1_outputs[1189];
    assign layer2_outputs[11647] = layer1_outputs[9070];
    assign layer2_outputs[11648] = ~(layer1_outputs[8626]);
    assign layer2_outputs[11649] = ~((layer1_outputs[3664]) ^ (layer1_outputs[1813]));
    assign layer2_outputs[11650] = ~(layer1_outputs[3646]);
    assign layer2_outputs[11651] = ~(layer1_outputs[8150]);
    assign layer2_outputs[11652] = layer1_outputs[6003];
    assign layer2_outputs[11653] = layer1_outputs[10302];
    assign layer2_outputs[11654] = ~((layer1_outputs[12286]) & (layer1_outputs[4954]));
    assign layer2_outputs[11655] = ~(layer1_outputs[11641]);
    assign layer2_outputs[11656] = ~((layer1_outputs[698]) & (layer1_outputs[10637]));
    assign layer2_outputs[11657] = ~(layer1_outputs[1512]);
    assign layer2_outputs[11658] = (layer1_outputs[7810]) & ~(layer1_outputs[6278]);
    assign layer2_outputs[11659] = ~(layer1_outputs[3746]);
    assign layer2_outputs[11660] = ~((layer1_outputs[11996]) ^ (layer1_outputs[10759]));
    assign layer2_outputs[11661] = ~(layer1_outputs[12473]);
    assign layer2_outputs[11662] = (layer1_outputs[12699]) & ~(layer1_outputs[12287]);
    assign layer2_outputs[11663] = ~((layer1_outputs[2560]) ^ (layer1_outputs[7812]));
    assign layer2_outputs[11664] = (layer1_outputs[1213]) & ~(layer1_outputs[1527]);
    assign layer2_outputs[11665] = layer1_outputs[4303];
    assign layer2_outputs[11666] = layer1_outputs[12144];
    assign layer2_outputs[11667] = layer1_outputs[4799];
    assign layer2_outputs[11668] = ~(layer1_outputs[10435]);
    assign layer2_outputs[11669] = ~(layer1_outputs[6014]);
    assign layer2_outputs[11670] = ~(layer1_outputs[12250]);
    assign layer2_outputs[11671] = (layer1_outputs[2414]) | (layer1_outputs[5949]);
    assign layer2_outputs[11672] = (layer1_outputs[8559]) & (layer1_outputs[2446]);
    assign layer2_outputs[11673] = ~(layer1_outputs[10310]);
    assign layer2_outputs[11674] = (layer1_outputs[5765]) ^ (layer1_outputs[9429]);
    assign layer2_outputs[11675] = ~((layer1_outputs[12499]) ^ (layer1_outputs[4487]));
    assign layer2_outputs[11676] = layer1_outputs[1237];
    assign layer2_outputs[11677] = ~(layer1_outputs[5869]);
    assign layer2_outputs[11678] = ~(layer1_outputs[1048]) | (layer1_outputs[11122]);
    assign layer2_outputs[11679] = (layer1_outputs[1510]) | (layer1_outputs[10522]);
    assign layer2_outputs[11680] = layer1_outputs[1914];
    assign layer2_outputs[11681] = ~((layer1_outputs[2766]) ^ (layer1_outputs[7059]));
    assign layer2_outputs[11682] = ~(layer1_outputs[5525]);
    assign layer2_outputs[11683] = layer1_outputs[6820];
    assign layer2_outputs[11684] = ~(layer1_outputs[867]);
    assign layer2_outputs[11685] = ~(layer1_outputs[10838]) | (layer1_outputs[9635]);
    assign layer2_outputs[11686] = (layer1_outputs[6875]) & ~(layer1_outputs[2373]);
    assign layer2_outputs[11687] = ~((layer1_outputs[5808]) & (layer1_outputs[9936]));
    assign layer2_outputs[11688] = (layer1_outputs[1498]) & ~(layer1_outputs[4330]);
    assign layer2_outputs[11689] = ~((layer1_outputs[2050]) | (layer1_outputs[8485]));
    assign layer2_outputs[11690] = ~(layer1_outputs[8953]);
    assign layer2_outputs[11691] = layer1_outputs[8144];
    assign layer2_outputs[11692] = (layer1_outputs[5908]) & ~(layer1_outputs[236]);
    assign layer2_outputs[11693] = ~((layer1_outputs[6869]) ^ (layer1_outputs[7824]));
    assign layer2_outputs[11694] = ~((layer1_outputs[7628]) | (layer1_outputs[7562]));
    assign layer2_outputs[11695] = layer1_outputs[1598];
    assign layer2_outputs[11696] = layer1_outputs[11547];
    assign layer2_outputs[11697] = ~((layer1_outputs[3593]) ^ (layer1_outputs[5806]));
    assign layer2_outputs[11698] = ~(layer1_outputs[11646]);
    assign layer2_outputs[11699] = layer1_outputs[11020];
    assign layer2_outputs[11700] = ~(layer1_outputs[8027]);
    assign layer2_outputs[11701] = ~((layer1_outputs[12270]) & (layer1_outputs[10663]));
    assign layer2_outputs[11702] = (layer1_outputs[479]) & ~(layer1_outputs[1459]);
    assign layer2_outputs[11703] = layer1_outputs[5008];
    assign layer2_outputs[11704] = (layer1_outputs[10508]) ^ (layer1_outputs[1199]);
    assign layer2_outputs[11705] = ~(layer1_outputs[5494]);
    assign layer2_outputs[11706] = ~(layer1_outputs[4411]);
    assign layer2_outputs[11707] = layer1_outputs[287];
    assign layer2_outputs[11708] = (layer1_outputs[423]) & (layer1_outputs[3194]);
    assign layer2_outputs[11709] = layer1_outputs[4978];
    assign layer2_outputs[11710] = ~(layer1_outputs[8327]);
    assign layer2_outputs[11711] = layer1_outputs[792];
    assign layer2_outputs[11712] = ~(layer1_outputs[3676]);
    assign layer2_outputs[11713] = ~(layer1_outputs[9143]);
    assign layer2_outputs[11714] = layer1_outputs[7256];
    assign layer2_outputs[11715] = ~(layer1_outputs[10151]);
    assign layer2_outputs[11716] = layer1_outputs[6710];
    assign layer2_outputs[11717] = layer1_outputs[10452];
    assign layer2_outputs[11718] = ~((layer1_outputs[1961]) ^ (layer1_outputs[3321]));
    assign layer2_outputs[11719] = layer1_outputs[5721];
    assign layer2_outputs[11720] = ~(layer1_outputs[8494]) | (layer1_outputs[6672]);
    assign layer2_outputs[11721] = ~(layer1_outputs[5440]);
    assign layer2_outputs[11722] = layer1_outputs[5635];
    assign layer2_outputs[11723] = ~(layer1_outputs[10444]);
    assign layer2_outputs[11724] = layer1_outputs[4009];
    assign layer2_outputs[11725] = ~((layer1_outputs[8295]) | (layer1_outputs[3855]));
    assign layer2_outputs[11726] = ~(layer1_outputs[11342]);
    assign layer2_outputs[11727] = layer1_outputs[545];
    assign layer2_outputs[11728] = (layer1_outputs[2059]) & (layer1_outputs[3973]);
    assign layer2_outputs[11729] = ~(layer1_outputs[12700]) | (layer1_outputs[231]);
    assign layer2_outputs[11730] = layer1_outputs[8270];
    assign layer2_outputs[11731] = layer1_outputs[11507];
    assign layer2_outputs[11732] = (layer1_outputs[4611]) & ~(layer1_outputs[8703]);
    assign layer2_outputs[11733] = ~((layer1_outputs[7776]) & (layer1_outputs[5694]));
    assign layer2_outputs[11734] = (layer1_outputs[4859]) ^ (layer1_outputs[3335]);
    assign layer2_outputs[11735] = ~(layer1_outputs[7777]);
    assign layer2_outputs[11736] = layer1_outputs[9659];
    assign layer2_outputs[11737] = layer1_outputs[5509];
    assign layer2_outputs[11738] = layer1_outputs[4974];
    assign layer2_outputs[11739] = ~(layer1_outputs[4563]) | (layer1_outputs[10797]);
    assign layer2_outputs[11740] = ~((layer1_outputs[10891]) | (layer1_outputs[8048]));
    assign layer2_outputs[11741] = ~(layer1_outputs[827]);
    assign layer2_outputs[11742] = ~(layer1_outputs[4986]);
    assign layer2_outputs[11743] = (layer1_outputs[6714]) ^ (layer1_outputs[11418]);
    assign layer2_outputs[11744] = ~(layer1_outputs[6913]);
    assign layer2_outputs[11745] = layer1_outputs[5630];
    assign layer2_outputs[11746] = ~((layer1_outputs[10556]) ^ (layer1_outputs[8658]));
    assign layer2_outputs[11747] = (layer1_outputs[203]) & ~(layer1_outputs[6004]);
    assign layer2_outputs[11748] = layer1_outputs[9274];
    assign layer2_outputs[11749] = layer1_outputs[7107];
    assign layer2_outputs[11750] = ~(layer1_outputs[10714]) | (layer1_outputs[4570]);
    assign layer2_outputs[11751] = ~(layer1_outputs[3772]);
    assign layer2_outputs[11752] = 1'b0;
    assign layer2_outputs[11753] = ~(layer1_outputs[10355]);
    assign layer2_outputs[11754] = layer1_outputs[6230];
    assign layer2_outputs[11755] = ~((layer1_outputs[765]) | (layer1_outputs[1538]));
    assign layer2_outputs[11756] = ~((layer1_outputs[10728]) ^ (layer1_outputs[9123]));
    assign layer2_outputs[11757] = ~(layer1_outputs[5268]);
    assign layer2_outputs[11758] = ~((layer1_outputs[8776]) & (layer1_outputs[10609]));
    assign layer2_outputs[11759] = ~(layer1_outputs[9915]) | (layer1_outputs[8450]);
    assign layer2_outputs[11760] = (layer1_outputs[1376]) & ~(layer1_outputs[834]);
    assign layer2_outputs[11761] = ~(layer1_outputs[908]);
    assign layer2_outputs[11762] = layer1_outputs[1491];
    assign layer2_outputs[11763] = layer1_outputs[3370];
    assign layer2_outputs[11764] = layer1_outputs[11377];
    assign layer2_outputs[11765] = ~(layer1_outputs[11165]) | (layer1_outputs[3587]);
    assign layer2_outputs[11766] = ~((layer1_outputs[1713]) ^ (layer1_outputs[185]));
    assign layer2_outputs[11767] = layer1_outputs[7629];
    assign layer2_outputs[11768] = layer1_outputs[1318];
    assign layer2_outputs[11769] = layer1_outputs[6020];
    assign layer2_outputs[11770] = ~((layer1_outputs[11731]) ^ (layer1_outputs[4997]));
    assign layer2_outputs[11771] = (layer1_outputs[9065]) ^ (layer1_outputs[10076]);
    assign layer2_outputs[11772] = ~(layer1_outputs[5749]);
    assign layer2_outputs[11773] = ~((layer1_outputs[3428]) ^ (layer1_outputs[7863]));
    assign layer2_outputs[11774] = ~(layer1_outputs[6639]);
    assign layer2_outputs[11775] = ~(layer1_outputs[1491]);
    assign layer2_outputs[11776] = layer1_outputs[8751];
    assign layer2_outputs[11777] = (layer1_outputs[6759]) & ~(layer1_outputs[4968]);
    assign layer2_outputs[11778] = layer1_outputs[8162];
    assign layer2_outputs[11779] = (layer1_outputs[8743]) & ~(layer1_outputs[2557]);
    assign layer2_outputs[11780] = ~(layer1_outputs[2398]);
    assign layer2_outputs[11781] = (layer1_outputs[2308]) ^ (layer1_outputs[12433]);
    assign layer2_outputs[11782] = (layer1_outputs[8890]) & ~(layer1_outputs[12513]);
    assign layer2_outputs[11783] = ~((layer1_outputs[4590]) & (layer1_outputs[11223]));
    assign layer2_outputs[11784] = ~((layer1_outputs[12231]) | (layer1_outputs[3086]));
    assign layer2_outputs[11785] = layer1_outputs[9866];
    assign layer2_outputs[11786] = ~((layer1_outputs[11332]) ^ (layer1_outputs[12356]));
    assign layer2_outputs[11787] = ~(layer1_outputs[11066]);
    assign layer2_outputs[11788] = ~(layer1_outputs[7599]);
    assign layer2_outputs[11789] = ~(layer1_outputs[12402]) | (layer1_outputs[11449]);
    assign layer2_outputs[11790] = (layer1_outputs[2014]) & ~(layer1_outputs[2916]);
    assign layer2_outputs[11791] = layer1_outputs[9471];
    assign layer2_outputs[11792] = layer1_outputs[8649];
    assign layer2_outputs[11793] = layer1_outputs[10198];
    assign layer2_outputs[11794] = ~(layer1_outputs[1998]);
    assign layer2_outputs[11795] = layer1_outputs[2026];
    assign layer2_outputs[11796] = ~(layer1_outputs[11496]);
    assign layer2_outputs[11797] = ~(layer1_outputs[5637]);
    assign layer2_outputs[11798] = (layer1_outputs[12024]) ^ (layer1_outputs[12427]);
    assign layer2_outputs[11799] = ~(layer1_outputs[3625]);
    assign layer2_outputs[11800] = ~(layer1_outputs[10689]);
    assign layer2_outputs[11801] = ~((layer1_outputs[4760]) & (layer1_outputs[10539]));
    assign layer2_outputs[11802] = (layer1_outputs[41]) & ~(layer1_outputs[5408]);
    assign layer2_outputs[11803] = ~((layer1_outputs[8704]) ^ (layer1_outputs[4827]));
    assign layer2_outputs[11804] = layer1_outputs[14];
    assign layer2_outputs[11805] = ~(layer1_outputs[8705]);
    assign layer2_outputs[11806] = ~(layer1_outputs[6776]);
    assign layer2_outputs[11807] = ~((layer1_outputs[11751]) & (layer1_outputs[3617]));
    assign layer2_outputs[11808] = (layer1_outputs[2086]) ^ (layer1_outputs[7410]);
    assign layer2_outputs[11809] = ~(layer1_outputs[11616]);
    assign layer2_outputs[11810] = (layer1_outputs[1028]) & ~(layer1_outputs[6661]);
    assign layer2_outputs[11811] = ~((layer1_outputs[11515]) | (layer1_outputs[11006]));
    assign layer2_outputs[11812] = layer1_outputs[9436];
    assign layer2_outputs[11813] = ~((layer1_outputs[2193]) ^ (layer1_outputs[10471]));
    assign layer2_outputs[11814] = layer1_outputs[12543];
    assign layer2_outputs[11815] = (layer1_outputs[3592]) & (layer1_outputs[1766]);
    assign layer2_outputs[11816] = ~(layer1_outputs[5354]) | (layer1_outputs[9235]);
    assign layer2_outputs[11817] = ~(layer1_outputs[12789]) | (layer1_outputs[4267]);
    assign layer2_outputs[11818] = ~(layer1_outputs[7987]);
    assign layer2_outputs[11819] = ~(layer1_outputs[12468]);
    assign layer2_outputs[11820] = ~(layer1_outputs[6690]) | (layer1_outputs[5304]);
    assign layer2_outputs[11821] = (layer1_outputs[2462]) & (layer1_outputs[1674]);
    assign layer2_outputs[11822] = (layer1_outputs[7309]) & (layer1_outputs[5651]);
    assign layer2_outputs[11823] = (layer1_outputs[814]) ^ (layer1_outputs[3917]);
    assign layer2_outputs[11824] = layer1_outputs[3210];
    assign layer2_outputs[11825] = ~(layer1_outputs[7686]);
    assign layer2_outputs[11826] = (layer1_outputs[7994]) | (layer1_outputs[8336]);
    assign layer2_outputs[11827] = ~(layer1_outputs[9067]);
    assign layer2_outputs[11828] = ~(layer1_outputs[11993]);
    assign layer2_outputs[11829] = ~(layer1_outputs[12650]);
    assign layer2_outputs[11830] = 1'b0;
    assign layer2_outputs[11831] = (layer1_outputs[1796]) ^ (layer1_outputs[8408]);
    assign layer2_outputs[11832] = (layer1_outputs[12673]) & (layer1_outputs[204]);
    assign layer2_outputs[11833] = (layer1_outputs[1838]) & ~(layer1_outputs[1990]);
    assign layer2_outputs[11834] = ~(layer1_outputs[4065]);
    assign layer2_outputs[11835] = layer1_outputs[9914];
    assign layer2_outputs[11836] = (layer1_outputs[4960]) | (layer1_outputs[12431]);
    assign layer2_outputs[11837] = ~(layer1_outputs[5321]);
    assign layer2_outputs[11838] = layer1_outputs[5723];
    assign layer2_outputs[11839] = ~(layer1_outputs[8261]);
    assign layer2_outputs[11840] = layer1_outputs[4236];
    assign layer2_outputs[11841] = layer1_outputs[8830];
    assign layer2_outputs[11842] = layer1_outputs[4874];
    assign layer2_outputs[11843] = ~(layer1_outputs[2111]);
    assign layer2_outputs[11844] = (layer1_outputs[5667]) & (layer1_outputs[3529]);
    assign layer2_outputs[11845] = ~(layer1_outputs[7112]) | (layer1_outputs[12788]);
    assign layer2_outputs[11846] = (layer1_outputs[2654]) ^ (layer1_outputs[2997]);
    assign layer2_outputs[11847] = (layer1_outputs[5897]) & (layer1_outputs[2029]);
    assign layer2_outputs[11848] = ~((layer1_outputs[443]) | (layer1_outputs[3053]));
    assign layer2_outputs[11849] = layer1_outputs[907];
    assign layer2_outputs[11850] = ~(layer1_outputs[5364]);
    assign layer2_outputs[11851] = ~(layer1_outputs[11968]);
    assign layer2_outputs[11852] = (layer1_outputs[2065]) & (layer1_outputs[171]);
    assign layer2_outputs[11853] = ~(layer1_outputs[9778]);
    assign layer2_outputs[11854] = (layer1_outputs[10470]) & ~(layer1_outputs[9379]);
    assign layer2_outputs[11855] = ~((layer1_outputs[7080]) ^ (layer1_outputs[10151]));
    assign layer2_outputs[11856] = layer1_outputs[4949];
    assign layer2_outputs[11857] = ~(layer1_outputs[4420]);
    assign layer2_outputs[11858] = layer1_outputs[9028];
    assign layer2_outputs[11859] = ~((layer1_outputs[4373]) ^ (layer1_outputs[6184]));
    assign layer2_outputs[11860] = layer1_outputs[5831];
    assign layer2_outputs[11861] = (layer1_outputs[12639]) | (layer1_outputs[12165]);
    assign layer2_outputs[11862] = layer1_outputs[5989];
    assign layer2_outputs[11863] = ~(layer1_outputs[757]);
    assign layer2_outputs[11864] = ~(layer1_outputs[8061]) | (layer1_outputs[7116]);
    assign layer2_outputs[11865] = (layer1_outputs[5819]) | (layer1_outputs[5902]);
    assign layer2_outputs[11866] = layer1_outputs[8288];
    assign layer2_outputs[11867] = ~(layer1_outputs[8364]);
    assign layer2_outputs[11868] = ~((layer1_outputs[1843]) | (layer1_outputs[606]));
    assign layer2_outputs[11869] = (layer1_outputs[3799]) | (layer1_outputs[2552]);
    assign layer2_outputs[11870] = ~((layer1_outputs[8495]) ^ (layer1_outputs[3391]));
    assign layer2_outputs[11871] = ~((layer1_outputs[708]) & (layer1_outputs[6698]));
    assign layer2_outputs[11872] = ~(layer1_outputs[12531]);
    assign layer2_outputs[11873] = ~(layer1_outputs[8760]);
    assign layer2_outputs[11874] = (layer1_outputs[1953]) & (layer1_outputs[11055]);
    assign layer2_outputs[11875] = ~(layer1_outputs[1421]);
    assign layer2_outputs[11876] = (layer1_outputs[9228]) & ~(layer1_outputs[8482]);
    assign layer2_outputs[11877] = ~(layer1_outputs[7796]);
    assign layer2_outputs[11878] = layer1_outputs[3065];
    assign layer2_outputs[11879] = ~(layer1_outputs[1875]) | (layer1_outputs[7282]);
    assign layer2_outputs[11880] = (layer1_outputs[12355]) & (layer1_outputs[8756]);
    assign layer2_outputs[11881] = (layer1_outputs[11917]) ^ (layer1_outputs[5516]);
    assign layer2_outputs[11882] = ~(layer1_outputs[10001]) | (layer1_outputs[4383]);
    assign layer2_outputs[11883] = ~(layer1_outputs[2047]) | (layer1_outputs[8438]);
    assign layer2_outputs[11884] = (layer1_outputs[5909]) | (layer1_outputs[9310]);
    assign layer2_outputs[11885] = layer1_outputs[365];
    assign layer2_outputs[11886] = (layer1_outputs[5372]) & ~(layer1_outputs[3833]);
    assign layer2_outputs[11887] = ~(layer1_outputs[5796]);
    assign layer2_outputs[11888] = ~((layer1_outputs[11914]) | (layer1_outputs[9813]));
    assign layer2_outputs[11889] = layer1_outputs[6957];
    assign layer2_outputs[11890] = ~((layer1_outputs[200]) | (layer1_outputs[9440]));
    assign layer2_outputs[11891] = ~(layer1_outputs[4241]);
    assign layer2_outputs[11892] = ~(layer1_outputs[11875]);
    assign layer2_outputs[11893] = ~((layer1_outputs[10056]) ^ (layer1_outputs[7257]));
    assign layer2_outputs[11894] = ~(layer1_outputs[11513]);
    assign layer2_outputs[11895] = (layer1_outputs[8793]) & ~(layer1_outputs[5431]);
    assign layer2_outputs[11896] = (layer1_outputs[9675]) | (layer1_outputs[5799]);
    assign layer2_outputs[11897] = ~(layer1_outputs[12011]);
    assign layer2_outputs[11898] = ~(layer1_outputs[1832]);
    assign layer2_outputs[11899] = (layer1_outputs[10854]) ^ (layer1_outputs[4212]);
    assign layer2_outputs[11900] = (layer1_outputs[11057]) & ~(layer1_outputs[3374]);
    assign layer2_outputs[11901] = ~(layer1_outputs[8684]) | (layer1_outputs[10840]);
    assign layer2_outputs[11902] = ~((layer1_outputs[7650]) & (layer1_outputs[817]));
    assign layer2_outputs[11903] = ~(layer1_outputs[9667]);
    assign layer2_outputs[11904] = (layer1_outputs[4376]) & ~(layer1_outputs[4386]);
    assign layer2_outputs[11905] = layer1_outputs[6204];
    assign layer2_outputs[11906] = layer1_outputs[10814];
    assign layer2_outputs[11907] = layer1_outputs[138];
    assign layer2_outputs[11908] = (layer1_outputs[8771]) ^ (layer1_outputs[5965]);
    assign layer2_outputs[11909] = ~(layer1_outputs[4410]) | (layer1_outputs[3921]);
    assign layer2_outputs[11910] = ~(layer1_outputs[8304]);
    assign layer2_outputs[11911] = layer1_outputs[11143];
    assign layer2_outputs[11912] = layer1_outputs[4584];
    assign layer2_outputs[11913] = (layer1_outputs[10140]) | (layer1_outputs[1901]);
    assign layer2_outputs[11914] = ~((layer1_outputs[4545]) | (layer1_outputs[5540]));
    assign layer2_outputs[11915] = ~(layer1_outputs[7236]);
    assign layer2_outputs[11916] = ~((layer1_outputs[12343]) ^ (layer1_outputs[2800]));
    assign layer2_outputs[11917] = ~(layer1_outputs[6666]) | (layer1_outputs[1358]);
    assign layer2_outputs[11918] = ~((layer1_outputs[11684]) | (layer1_outputs[6151]));
    assign layer2_outputs[11919] = (layer1_outputs[10161]) & (layer1_outputs[3479]);
    assign layer2_outputs[11920] = ~(layer1_outputs[11098]);
    assign layer2_outputs[11921] = layer1_outputs[5048];
    assign layer2_outputs[11922] = (layer1_outputs[3314]) | (layer1_outputs[8125]);
    assign layer2_outputs[11923] = layer1_outputs[11036];
    assign layer2_outputs[11924] = ~(layer1_outputs[8153]);
    assign layer2_outputs[11925] = ~(layer1_outputs[12529]);
    assign layer2_outputs[11926] = ~((layer1_outputs[3699]) | (layer1_outputs[5425]));
    assign layer2_outputs[11927] = ~((layer1_outputs[6032]) & (layer1_outputs[12092]));
    assign layer2_outputs[11928] = (layer1_outputs[5345]) ^ (layer1_outputs[9593]);
    assign layer2_outputs[11929] = layer1_outputs[4025];
    assign layer2_outputs[11930] = layer1_outputs[4622];
    assign layer2_outputs[11931] = layer1_outputs[5645];
    assign layer2_outputs[11932] = ~(layer1_outputs[10220]);
    assign layer2_outputs[11933] = ~(layer1_outputs[8516]) | (layer1_outputs[272]);
    assign layer2_outputs[11934] = ~(layer1_outputs[11672]) | (layer1_outputs[5629]);
    assign layer2_outputs[11935] = ~((layer1_outputs[12009]) ^ (layer1_outputs[6096]));
    assign layer2_outputs[11936] = ~((layer1_outputs[2061]) ^ (layer1_outputs[6395]));
    assign layer2_outputs[11937] = (layer1_outputs[4505]) | (layer1_outputs[4191]);
    assign layer2_outputs[11938] = ~(layer1_outputs[12277]);
    assign layer2_outputs[11939] = ~(layer1_outputs[590]);
    assign layer2_outputs[11940] = ~(layer1_outputs[2133]);
    assign layer2_outputs[11941] = ~((layer1_outputs[10804]) | (layer1_outputs[5310]));
    assign layer2_outputs[11942] = layer1_outputs[8437];
    assign layer2_outputs[11943] = (layer1_outputs[8029]) & (layer1_outputs[2553]);
    assign layer2_outputs[11944] = layer1_outputs[4868];
    assign layer2_outputs[11945] = (layer1_outputs[9005]) & ~(layer1_outputs[1910]);
    assign layer2_outputs[11946] = ~(layer1_outputs[8446]) | (layer1_outputs[10474]);
    assign layer2_outputs[11947] = ~((layer1_outputs[11342]) ^ (layer1_outputs[10768]));
    assign layer2_outputs[11948] = layer1_outputs[2221];
    assign layer2_outputs[11949] = ~(layer1_outputs[1364]);
    assign layer2_outputs[11950] = ~(layer1_outputs[6015]);
    assign layer2_outputs[11951] = ~((layer1_outputs[7535]) & (layer1_outputs[2181]));
    assign layer2_outputs[11952] = (layer1_outputs[6662]) ^ (layer1_outputs[9280]);
    assign layer2_outputs[11953] = layer1_outputs[7126];
    assign layer2_outputs[11954] = layer1_outputs[3910];
    assign layer2_outputs[11955] = layer1_outputs[11954];
    assign layer2_outputs[11956] = ~(layer1_outputs[1765]);
    assign layer2_outputs[11957] = ~(layer1_outputs[1520]) | (layer1_outputs[10146]);
    assign layer2_outputs[11958] = layer1_outputs[8442];
    assign layer2_outputs[11959] = ~(layer1_outputs[552]);
    assign layer2_outputs[11960] = (layer1_outputs[8053]) ^ (layer1_outputs[8883]);
    assign layer2_outputs[11961] = (layer1_outputs[6678]) & ~(layer1_outputs[12461]);
    assign layer2_outputs[11962] = ~(layer1_outputs[404]);
    assign layer2_outputs[11963] = (layer1_outputs[9425]) & (layer1_outputs[5576]);
    assign layer2_outputs[11964] = (layer1_outputs[12396]) & ~(layer1_outputs[1930]);
    assign layer2_outputs[11965] = ~(layer1_outputs[8800]);
    assign layer2_outputs[11966] = (layer1_outputs[1807]) ^ (layer1_outputs[12301]);
    assign layer2_outputs[11967] = ~(layer1_outputs[8300]);
    assign layer2_outputs[11968] = layer1_outputs[11652];
    assign layer2_outputs[11969] = ~(layer1_outputs[12161]);
    assign layer2_outputs[11970] = layer1_outputs[2745];
    assign layer2_outputs[11971] = ~((layer1_outputs[8180]) | (layer1_outputs[369]));
    assign layer2_outputs[11972] = (layer1_outputs[6485]) & ~(layer1_outputs[6257]);
    assign layer2_outputs[11973] = ~(layer1_outputs[7050]) | (layer1_outputs[1209]);
    assign layer2_outputs[11974] = ~(layer1_outputs[5779]) | (layer1_outputs[9309]);
    assign layer2_outputs[11975] = ~(layer1_outputs[8152]) | (layer1_outputs[1514]);
    assign layer2_outputs[11976] = ~(layer1_outputs[7461]) | (layer1_outputs[8408]);
    assign layer2_outputs[11977] = layer1_outputs[1297];
    assign layer2_outputs[11978] = layer1_outputs[4234];
    assign layer2_outputs[11979] = layer1_outputs[9604];
    assign layer2_outputs[11980] = layer1_outputs[1283];
    assign layer2_outputs[11981] = ~((layer1_outputs[3395]) ^ (layer1_outputs[9481]));
    assign layer2_outputs[11982] = layer1_outputs[11398];
    assign layer2_outputs[11983] = layer1_outputs[7609];
    assign layer2_outputs[11984] = layer1_outputs[833];
    assign layer2_outputs[11985] = (layer1_outputs[933]) & ~(layer1_outputs[5373]);
    assign layer2_outputs[11986] = ~(layer1_outputs[1984]);
    assign layer2_outputs[11987] = ~(layer1_outputs[6493]) | (layer1_outputs[4442]);
    assign layer2_outputs[11988] = layer1_outputs[12782];
    assign layer2_outputs[11989] = (layer1_outputs[1029]) & ~(layer1_outputs[9974]);
    assign layer2_outputs[11990] = (layer1_outputs[720]) & (layer1_outputs[5127]);
    assign layer2_outputs[11991] = ~(layer1_outputs[2554]);
    assign layer2_outputs[11992] = ~((layer1_outputs[2230]) | (layer1_outputs[4746]));
    assign layer2_outputs[11993] = layer1_outputs[8099];
    assign layer2_outputs[11994] = 1'b0;
    assign layer2_outputs[11995] = ~(layer1_outputs[2145]);
    assign layer2_outputs[11996] = ~(layer1_outputs[8766]);
    assign layer2_outputs[11997] = ~(layer1_outputs[2218]);
    assign layer2_outputs[11998] = ~(layer1_outputs[11754]);
    assign layer2_outputs[11999] = layer1_outputs[2767];
    assign layer2_outputs[12000] = ~((layer1_outputs[7475]) & (layer1_outputs[5679]));
    assign layer2_outputs[12001] = ~((layer1_outputs[3946]) | (layer1_outputs[935]));
    assign layer2_outputs[12002] = layer1_outputs[9229];
    assign layer2_outputs[12003] = layer1_outputs[6715];
    assign layer2_outputs[12004] = (layer1_outputs[4832]) ^ (layer1_outputs[7483]);
    assign layer2_outputs[12005] = ~(layer1_outputs[9133]);
    assign layer2_outputs[12006] = (layer1_outputs[12578]) ^ (layer1_outputs[9337]);
    assign layer2_outputs[12007] = ~(layer1_outputs[2239]) | (layer1_outputs[1027]);
    assign layer2_outputs[12008] = (layer1_outputs[12214]) ^ (layer1_outputs[10621]);
    assign layer2_outputs[12009] = (layer1_outputs[4805]) & ~(layer1_outputs[11152]);
    assign layer2_outputs[12010] = ~(layer1_outputs[6878]);
    assign layer2_outputs[12011] = ~(layer1_outputs[5503]);
    assign layer2_outputs[12012] = ~(layer1_outputs[6150]);
    assign layer2_outputs[12013] = ~(layer1_outputs[3868]);
    assign layer2_outputs[12014] = (layer1_outputs[5183]) & ~(layer1_outputs[7795]);
    assign layer2_outputs[12015] = layer1_outputs[11423];
    assign layer2_outputs[12016] = (layer1_outputs[8008]) | (layer1_outputs[6125]);
    assign layer2_outputs[12017] = layer1_outputs[5082];
    assign layer2_outputs[12018] = 1'b0;
    assign layer2_outputs[12019] = (layer1_outputs[11565]) & ~(layer1_outputs[763]);
    assign layer2_outputs[12020] = (layer1_outputs[7234]) ^ (layer1_outputs[8443]);
    assign layer2_outputs[12021] = ~(layer1_outputs[957]);
    assign layer2_outputs[12022] = 1'b1;
    assign layer2_outputs[12023] = layer1_outputs[5015];
    assign layer2_outputs[12024] = layer1_outputs[11762];
    assign layer2_outputs[12025] = ~(layer1_outputs[7526]);
    assign layer2_outputs[12026] = (layer1_outputs[7275]) | (layer1_outputs[8234]);
    assign layer2_outputs[12027] = (layer1_outputs[2039]) ^ (layer1_outputs[6186]);
    assign layer2_outputs[12028] = (layer1_outputs[11543]) & ~(layer1_outputs[11452]);
    assign layer2_outputs[12029] = ~(layer1_outputs[3645]);
    assign layer2_outputs[12030] = (layer1_outputs[4265]) | (layer1_outputs[10073]);
    assign layer2_outputs[12031] = layer1_outputs[12206];
    assign layer2_outputs[12032] = ~(layer1_outputs[2525]);
    assign layer2_outputs[12033] = ~(layer1_outputs[9111]);
    assign layer2_outputs[12034] = ~((layer1_outputs[4229]) | (layer1_outputs[10601]));
    assign layer2_outputs[12035] = (layer1_outputs[4157]) ^ (layer1_outputs[3213]);
    assign layer2_outputs[12036] = ~((layer1_outputs[1480]) ^ (layer1_outputs[3833]));
    assign layer2_outputs[12037] = ~((layer1_outputs[10946]) ^ (layer1_outputs[9947]));
    assign layer2_outputs[12038] = ~(layer1_outputs[6284]) | (layer1_outputs[11776]);
    assign layer2_outputs[12039] = layer1_outputs[10535];
    assign layer2_outputs[12040] = ~((layer1_outputs[849]) ^ (layer1_outputs[9772]));
    assign layer2_outputs[12041] = layer1_outputs[9774];
    assign layer2_outputs[12042] = ~(layer1_outputs[1428]) | (layer1_outputs[11854]);
    assign layer2_outputs[12043] = ~(layer1_outputs[8375]);
    assign layer2_outputs[12044] = layer1_outputs[10010];
    assign layer2_outputs[12045] = ~(layer1_outputs[3310]);
    assign layer2_outputs[12046] = layer1_outputs[5487];
    assign layer2_outputs[12047] = ~(layer1_outputs[5481]) | (layer1_outputs[4540]);
    assign layer2_outputs[12048] = ~(layer1_outputs[5991]);
    assign layer2_outputs[12049] = ~((layer1_outputs[10923]) | (layer1_outputs[8415]));
    assign layer2_outputs[12050] = layer1_outputs[7433];
    assign layer2_outputs[12051] = ~((layer1_outputs[3985]) | (layer1_outputs[9670]));
    assign layer2_outputs[12052] = ~(layer1_outputs[5471]);
    assign layer2_outputs[12053] = (layer1_outputs[7853]) | (layer1_outputs[12078]);
    assign layer2_outputs[12054] = ~(layer1_outputs[1330]) | (layer1_outputs[8078]);
    assign layer2_outputs[12055] = layer1_outputs[3082];
    assign layer2_outputs[12056] = layer1_outputs[10350];
    assign layer2_outputs[12057] = ~((layer1_outputs[7329]) & (layer1_outputs[12131]));
    assign layer2_outputs[12058] = layer1_outputs[11771];
    assign layer2_outputs[12059] = (layer1_outputs[8398]) & ~(layer1_outputs[4486]);
    assign layer2_outputs[12060] = ~(layer1_outputs[5515]) | (layer1_outputs[8255]);
    assign layer2_outputs[12061] = ~(layer1_outputs[9586]);
    assign layer2_outputs[12062] = ~(layer1_outputs[12401]);
    assign layer2_outputs[12063] = ~(layer1_outputs[7947]) | (layer1_outputs[4784]);
    assign layer2_outputs[12064] = layer1_outputs[9556];
    assign layer2_outputs[12065] = layer1_outputs[6381];
    assign layer2_outputs[12066] = ~(layer1_outputs[729]) | (layer1_outputs[4747]);
    assign layer2_outputs[12067] = ~(layer1_outputs[10341]) | (layer1_outputs[7983]);
    assign layer2_outputs[12068] = ~((layer1_outputs[8443]) & (layer1_outputs[2241]));
    assign layer2_outputs[12069] = ~((layer1_outputs[8247]) ^ (layer1_outputs[504]));
    assign layer2_outputs[12070] = ~((layer1_outputs[6272]) & (layer1_outputs[7958]));
    assign layer2_outputs[12071] = ~(layer1_outputs[6243]);
    assign layer2_outputs[12072] = ~((layer1_outputs[637]) ^ (layer1_outputs[8941]));
    assign layer2_outputs[12073] = ~(layer1_outputs[11011]);
    assign layer2_outputs[12074] = (layer1_outputs[4256]) | (layer1_outputs[10981]);
    assign layer2_outputs[12075] = (layer1_outputs[5756]) & ~(layer1_outputs[8207]);
    assign layer2_outputs[12076] = layer1_outputs[3884];
    assign layer2_outputs[12077] = layer1_outputs[10641];
    assign layer2_outputs[12078] = (layer1_outputs[25]) ^ (layer1_outputs[6326]);
    assign layer2_outputs[12079] = layer1_outputs[10895];
    assign layer2_outputs[12080] = layer1_outputs[1343];
    assign layer2_outputs[12081] = (layer1_outputs[1662]) ^ (layer1_outputs[9168]);
    assign layer2_outputs[12082] = ~(layer1_outputs[7746]);
    assign layer2_outputs[12083] = (layer1_outputs[6423]) ^ (layer1_outputs[4388]);
    assign layer2_outputs[12084] = layer1_outputs[253];
    assign layer2_outputs[12085] = (layer1_outputs[2604]) & ~(layer1_outputs[3422]);
    assign layer2_outputs[12086] = (layer1_outputs[10715]) & ~(layer1_outputs[2174]);
    assign layer2_outputs[12087] = ~(layer1_outputs[12340]);
    assign layer2_outputs[12088] = ~(layer1_outputs[3158]);
    assign layer2_outputs[12089] = ~((layer1_outputs[2776]) ^ (layer1_outputs[3526]));
    assign layer2_outputs[12090] = ~(layer1_outputs[12058]);
    assign layer2_outputs[12091] = (layer1_outputs[10382]) | (layer1_outputs[1225]);
    assign layer2_outputs[12092] = layer1_outputs[8556];
    assign layer2_outputs[12093] = layer1_outputs[681];
    assign layer2_outputs[12094] = ~((layer1_outputs[9035]) ^ (layer1_outputs[5109]));
    assign layer2_outputs[12095] = ~(layer1_outputs[12477]);
    assign layer2_outputs[12096] = ~(layer1_outputs[5341]) | (layer1_outputs[10341]);
    assign layer2_outputs[12097] = (layer1_outputs[86]) & ~(layer1_outputs[10163]);
    assign layer2_outputs[12098] = layer1_outputs[9614];
    assign layer2_outputs[12099] = layer1_outputs[2783];
    assign layer2_outputs[12100] = (layer1_outputs[9321]) | (layer1_outputs[10082]);
    assign layer2_outputs[12101] = layer1_outputs[2021];
    assign layer2_outputs[12102] = ~((layer1_outputs[847]) & (layer1_outputs[11790]));
    assign layer2_outputs[12103] = (layer1_outputs[3977]) ^ (layer1_outputs[796]);
    assign layer2_outputs[12104] = (layer1_outputs[2135]) & ~(layer1_outputs[2261]);
    assign layer2_outputs[12105] = (layer1_outputs[3443]) & (layer1_outputs[8908]);
    assign layer2_outputs[12106] = ~(layer1_outputs[5647]) | (layer1_outputs[2481]);
    assign layer2_outputs[12107] = layer1_outputs[7693];
    assign layer2_outputs[12108] = ~(layer1_outputs[3248]) | (layer1_outputs[7479]);
    assign layer2_outputs[12109] = ~((layer1_outputs[4713]) ^ (layer1_outputs[11380]));
    assign layer2_outputs[12110] = layer1_outputs[1927];
    assign layer2_outputs[12111] = (layer1_outputs[12145]) ^ (layer1_outputs[1164]);
    assign layer2_outputs[12112] = ~(layer1_outputs[122]) | (layer1_outputs[6746]);
    assign layer2_outputs[12113] = layer1_outputs[10468];
    assign layer2_outputs[12114] = layer1_outputs[740];
    assign layer2_outputs[12115] = ~((layer1_outputs[2388]) & (layer1_outputs[11544]));
    assign layer2_outputs[12116] = ~(layer1_outputs[2815]);
    assign layer2_outputs[12117] = layer1_outputs[10210];
    assign layer2_outputs[12118] = layer1_outputs[3349];
    assign layer2_outputs[12119] = ~(layer1_outputs[2064]);
    assign layer2_outputs[12120] = layer1_outputs[2866];
    assign layer2_outputs[12121] = ~(layer1_outputs[3474]) | (layer1_outputs[10242]);
    assign layer2_outputs[12122] = ~(layer1_outputs[9627]) | (layer1_outputs[3886]);
    assign layer2_outputs[12123] = (layer1_outputs[2551]) & ~(layer1_outputs[12164]);
    assign layer2_outputs[12124] = (layer1_outputs[8600]) ^ (layer1_outputs[11618]);
    assign layer2_outputs[12125] = layer1_outputs[9479];
    assign layer2_outputs[12126] = (layer1_outputs[3631]) & (layer1_outputs[6495]);
    assign layer2_outputs[12127] = ~((layer1_outputs[6870]) ^ (layer1_outputs[3733]));
    assign layer2_outputs[12128] = layer1_outputs[8137];
    assign layer2_outputs[12129] = ~((layer1_outputs[10746]) & (layer1_outputs[5203]));
    assign layer2_outputs[12130] = ~((layer1_outputs[4920]) ^ (layer1_outputs[7813]));
    assign layer2_outputs[12131] = ~((layer1_outputs[4801]) ^ (layer1_outputs[5732]));
    assign layer2_outputs[12132] = ~((layer1_outputs[1438]) | (layer1_outputs[578]));
    assign layer2_outputs[12133] = ~((layer1_outputs[9209]) & (layer1_outputs[8682]));
    assign layer2_outputs[12134] = ~(layer1_outputs[8335]);
    assign layer2_outputs[12135] = layer1_outputs[11815];
    assign layer2_outputs[12136] = layer1_outputs[9656];
    assign layer2_outputs[12137] = ~(layer1_outputs[9093]) | (layer1_outputs[1919]);
    assign layer2_outputs[12138] = layer1_outputs[2683];
    assign layer2_outputs[12139] = ~((layer1_outputs[3353]) | (layer1_outputs[7209]));
    assign layer2_outputs[12140] = (layer1_outputs[6458]) & ~(layer1_outputs[0]);
    assign layer2_outputs[12141] = ~(layer1_outputs[1697]) | (layer1_outputs[147]);
    assign layer2_outputs[12142] = layer1_outputs[3077];
    assign layer2_outputs[12143] = ~(layer1_outputs[1803]);
    assign layer2_outputs[12144] = layer1_outputs[2787];
    assign layer2_outputs[12145] = ~(layer1_outputs[4609]);
    assign layer2_outputs[12146] = ~(layer1_outputs[6562]);
    assign layer2_outputs[12147] = ~(layer1_outputs[6248]) | (layer1_outputs[1607]);
    assign layer2_outputs[12148] = ~((layer1_outputs[6862]) & (layer1_outputs[7401]));
    assign layer2_outputs[12149] = layer1_outputs[2144];
    assign layer2_outputs[12150] = layer1_outputs[6867];
    assign layer2_outputs[12151] = layer1_outputs[2742];
    assign layer2_outputs[12152] = ~(layer1_outputs[10639]);
    assign layer2_outputs[12153] = ~(layer1_outputs[11719]) | (layer1_outputs[4268]);
    assign layer2_outputs[12154] = layer1_outputs[11391];
    assign layer2_outputs[12155] = layer1_outputs[3638];
    assign layer2_outputs[12156] = (layer1_outputs[9731]) & (layer1_outputs[8905]);
    assign layer2_outputs[12157] = layer1_outputs[7034];
    assign layer2_outputs[12158] = ~((layer1_outputs[4105]) ^ (layer1_outputs[12581]));
    assign layer2_outputs[12159] = (layer1_outputs[5190]) & (layer1_outputs[8303]);
    assign layer2_outputs[12160] = ~((layer1_outputs[5598]) | (layer1_outputs[7756]));
    assign layer2_outputs[12161] = ~(layer1_outputs[211]) | (layer1_outputs[5312]);
    assign layer2_outputs[12162] = (layer1_outputs[6734]) ^ (layer1_outputs[10516]);
    assign layer2_outputs[12163] = (layer1_outputs[4483]) & (layer1_outputs[4931]);
    assign layer2_outputs[12164] = (layer1_outputs[358]) & ~(layer1_outputs[8424]);
    assign layer2_outputs[12165] = layer1_outputs[9794];
    assign layer2_outputs[12166] = (layer1_outputs[12062]) & ~(layer1_outputs[2868]);
    assign layer2_outputs[12167] = ~(layer1_outputs[5507]);
    assign layer2_outputs[12168] = ~(layer1_outputs[2236]) | (layer1_outputs[474]);
    assign layer2_outputs[12169] = (layer1_outputs[1631]) & ~(layer1_outputs[5165]);
    assign layer2_outputs[12170] = ~((layer1_outputs[2889]) ^ (layer1_outputs[6410]));
    assign layer2_outputs[12171] = ~(layer1_outputs[11191]);
    assign layer2_outputs[12172] = ~(layer1_outputs[11182]) | (layer1_outputs[7364]);
    assign layer2_outputs[12173] = layer1_outputs[851];
    assign layer2_outputs[12174] = layer1_outputs[2484];
    assign layer2_outputs[12175] = ~(layer1_outputs[5264]);
    assign layer2_outputs[12176] = ~(layer1_outputs[6319]);
    assign layer2_outputs[12177] = ~(layer1_outputs[1162]);
    assign layer2_outputs[12178] = ~(layer1_outputs[8370]);
    assign layer2_outputs[12179] = ~(layer1_outputs[9324]);
    assign layer2_outputs[12180] = ~((layer1_outputs[7246]) | (layer1_outputs[12601]));
    assign layer2_outputs[12181] = ~((layer1_outputs[7960]) | (layer1_outputs[9245]));
    assign layer2_outputs[12182] = (layer1_outputs[1616]) & (layer1_outputs[11542]);
    assign layer2_outputs[12183] = ~(layer1_outputs[9123]);
    assign layer2_outputs[12184] = (layer1_outputs[10942]) ^ (layer1_outputs[10883]);
    assign layer2_outputs[12185] = ~(layer1_outputs[4386]);
    assign layer2_outputs[12186] = layer1_outputs[7542];
    assign layer2_outputs[12187] = layer1_outputs[9369];
    assign layer2_outputs[12188] = ~(layer1_outputs[2278]);
    assign layer2_outputs[12189] = layer1_outputs[9468];
    assign layer2_outputs[12190] = layer1_outputs[694];
    assign layer2_outputs[12191] = layer1_outputs[8561];
    assign layer2_outputs[12192] = ~(layer1_outputs[6386]);
    assign layer2_outputs[12193] = ~(layer1_outputs[3428]) | (layer1_outputs[12161]);
    assign layer2_outputs[12194] = ~(layer1_outputs[247]);
    assign layer2_outputs[12195] = (layer1_outputs[8724]) ^ (layer1_outputs[7076]);
    assign layer2_outputs[12196] = layer1_outputs[8843];
    assign layer2_outputs[12197] = ~(layer1_outputs[8012]);
    assign layer2_outputs[12198] = layer1_outputs[10247];
    assign layer2_outputs[12199] = ~(layer1_outputs[10571]);
    assign layer2_outputs[12200] = (layer1_outputs[7187]) ^ (layer1_outputs[5572]);
    assign layer2_outputs[12201] = ~((layer1_outputs[4091]) & (layer1_outputs[10910]));
    assign layer2_outputs[12202] = ~((layer1_outputs[1137]) ^ (layer1_outputs[1562]));
    assign layer2_outputs[12203] = (layer1_outputs[7445]) ^ (layer1_outputs[6439]);
    assign layer2_outputs[12204] = ~((layer1_outputs[7948]) & (layer1_outputs[611]));
    assign layer2_outputs[12205] = ~((layer1_outputs[3899]) & (layer1_outputs[2929]));
    assign layer2_outputs[12206] = ~((layer1_outputs[2492]) | (layer1_outputs[9034]));
    assign layer2_outputs[12207] = (layer1_outputs[5205]) & ~(layer1_outputs[6171]);
    assign layer2_outputs[12208] = ~(layer1_outputs[5530]);
    assign layer2_outputs[12209] = ~(layer1_outputs[7862]);
    assign layer2_outputs[12210] = ~((layer1_outputs[8886]) ^ (layer1_outputs[11461]));
    assign layer2_outputs[12211] = layer1_outputs[2743];
    assign layer2_outputs[12212] = ~(layer1_outputs[7097]) | (layer1_outputs[1912]);
    assign layer2_outputs[12213] = ~(layer1_outputs[2330]) | (layer1_outputs[5448]);
    assign layer2_outputs[12214] = ~(layer1_outputs[11525]);
    assign layer2_outputs[12215] = layer1_outputs[3427];
    assign layer2_outputs[12216] = (layer1_outputs[11465]) ^ (layer1_outputs[6297]);
    assign layer2_outputs[12217] = layer1_outputs[2565];
    assign layer2_outputs[12218] = layer1_outputs[3893];
    assign layer2_outputs[12219] = layer1_outputs[10254];
    assign layer2_outputs[12220] = ~((layer1_outputs[12595]) & (layer1_outputs[12063]));
    assign layer2_outputs[12221] = ~((layer1_outputs[1661]) ^ (layer1_outputs[12693]));
    assign layer2_outputs[12222] = ~(layer1_outputs[11913]);
    assign layer2_outputs[12223] = ~(layer1_outputs[8402]);
    assign layer2_outputs[12224] = ~((layer1_outputs[6861]) & (layer1_outputs[11935]));
    assign layer2_outputs[12225] = (layer1_outputs[2544]) & (layer1_outputs[1575]);
    assign layer2_outputs[12226] = ~((layer1_outputs[10763]) | (layer1_outputs[6345]));
    assign layer2_outputs[12227] = (layer1_outputs[6409]) ^ (layer1_outputs[1833]);
    assign layer2_outputs[12228] = ~(layer1_outputs[10523]) | (layer1_outputs[6846]);
    assign layer2_outputs[12229] = ~(layer1_outputs[835]);
    assign layer2_outputs[12230] = ~(layer1_outputs[5273]);
    assign layer2_outputs[12231] = (layer1_outputs[12057]) & ~(layer1_outputs[3524]);
    assign layer2_outputs[12232] = ~(layer1_outputs[12694]) | (layer1_outputs[6202]);
    assign layer2_outputs[12233] = ~(layer1_outputs[12643]) | (layer1_outputs[6629]);
    assign layer2_outputs[12234] = ~(layer1_outputs[8116]);
    assign layer2_outputs[12235] = ~(layer1_outputs[3522]);
    assign layer2_outputs[12236] = ~((layer1_outputs[4854]) | (layer1_outputs[175]));
    assign layer2_outputs[12237] = layer1_outputs[6821];
    assign layer2_outputs[12238] = ~(layer1_outputs[96]);
    assign layer2_outputs[12239] = layer1_outputs[5713];
    assign layer2_outputs[12240] = layer1_outputs[11691];
    assign layer2_outputs[12241] = ~(layer1_outputs[271]);
    assign layer2_outputs[12242] = layer1_outputs[2203];
    assign layer2_outputs[12243] = ~((layer1_outputs[1043]) ^ (layer1_outputs[1435]));
    assign layer2_outputs[12244] = (layer1_outputs[7135]) & (layer1_outputs[3571]);
    assign layer2_outputs[12245] = ~((layer1_outputs[585]) & (layer1_outputs[6296]));
    assign layer2_outputs[12246] = (layer1_outputs[7125]) ^ (layer1_outputs[11844]);
    assign layer2_outputs[12247] = ~(layer1_outputs[2689]);
    assign layer2_outputs[12248] = ~(layer1_outputs[7146]) | (layer1_outputs[8436]);
    assign layer2_outputs[12249] = ~(layer1_outputs[11905]);
    assign layer2_outputs[12250] = ~(layer1_outputs[62]);
    assign layer2_outputs[12251] = (layer1_outputs[9607]) ^ (layer1_outputs[8668]);
    assign layer2_outputs[12252] = ~((layer1_outputs[10124]) ^ (layer1_outputs[8191]));
    assign layer2_outputs[12253] = ~((layer1_outputs[1749]) & (layer1_outputs[171]));
    assign layer2_outputs[12254] = (layer1_outputs[10439]) ^ (layer1_outputs[4225]);
    assign layer2_outputs[12255] = layer1_outputs[11099];
    assign layer2_outputs[12256] = ~((layer1_outputs[3897]) ^ (layer1_outputs[12557]));
    assign layer2_outputs[12257] = (layer1_outputs[639]) & (layer1_outputs[9899]);
    assign layer2_outputs[12258] = layer1_outputs[7974];
    assign layer2_outputs[12259] = ~((layer1_outputs[8699]) | (layer1_outputs[5420]));
    assign layer2_outputs[12260] = ~((layer1_outputs[1613]) | (layer1_outputs[6498]));
    assign layer2_outputs[12261] = (layer1_outputs[813]) & ~(layer1_outputs[12340]);
    assign layer2_outputs[12262] = (layer1_outputs[3497]) | (layer1_outputs[1198]);
    assign layer2_outputs[12263] = layer1_outputs[6165];
    assign layer2_outputs[12264] = ~(layer1_outputs[5279]);
    assign layer2_outputs[12265] = ~(layer1_outputs[2275]);
    assign layer2_outputs[12266] = ~(layer1_outputs[5995]);
    assign layer2_outputs[12267] = layer1_outputs[11190];
    assign layer2_outputs[12268] = ~(layer1_outputs[4295]);
    assign layer2_outputs[12269] = (layer1_outputs[1532]) ^ (layer1_outputs[7543]);
    assign layer2_outputs[12270] = ~(layer1_outputs[5495]);
    assign layer2_outputs[12271] = ~((layer1_outputs[11136]) & (layer1_outputs[3715]));
    assign layer2_outputs[12272] = (layer1_outputs[5489]) & (layer1_outputs[5583]);
    assign layer2_outputs[12273] = ~((layer1_outputs[11749]) | (layer1_outputs[5791]));
    assign layer2_outputs[12274] = (layer1_outputs[2976]) | (layer1_outputs[2981]);
    assign layer2_outputs[12275] = layer1_outputs[9038];
    assign layer2_outputs[12276] = ~(layer1_outputs[5911]);
    assign layer2_outputs[12277] = ~(layer1_outputs[5382]) | (layer1_outputs[9602]);
    assign layer2_outputs[12278] = ~(layer1_outputs[5441]) | (layer1_outputs[7846]);
    assign layer2_outputs[12279] = layer1_outputs[1080];
    assign layer2_outputs[12280] = ~((layer1_outputs[8661]) ^ (layer1_outputs[4790]));
    assign layer2_outputs[12281] = layer1_outputs[809];
    assign layer2_outputs[12282] = (layer1_outputs[11311]) ^ (layer1_outputs[8491]);
    assign layer2_outputs[12283] = ~(layer1_outputs[7477]) | (layer1_outputs[3297]);
    assign layer2_outputs[12284] = ~(layer1_outputs[8121]);
    assign layer2_outputs[12285] = ~((layer1_outputs[340]) ^ (layer1_outputs[3548]));
    assign layer2_outputs[12286] = (layer1_outputs[12035]) ^ (layer1_outputs[9861]);
    assign layer2_outputs[12287] = ~(layer1_outputs[5603]);
    assign layer2_outputs[12288] = layer1_outputs[9674];
    assign layer2_outputs[12289] = (layer1_outputs[6469]) & ~(layer1_outputs[5761]);
    assign layer2_outputs[12290] = layer1_outputs[11811];
    assign layer2_outputs[12291] = ~(layer1_outputs[3208]);
    assign layer2_outputs[12292] = ~(layer1_outputs[7671]);
    assign layer2_outputs[12293] = ~(layer1_outputs[93]);
    assign layer2_outputs[12294] = (layer1_outputs[2618]) ^ (layer1_outputs[4830]);
    assign layer2_outputs[12295] = layer1_outputs[9231];
    assign layer2_outputs[12296] = ~(layer1_outputs[12683]) | (layer1_outputs[3093]);
    assign layer2_outputs[12297] = ~((layer1_outputs[8643]) & (layer1_outputs[2170]));
    assign layer2_outputs[12298] = ~(layer1_outputs[8930]);
    assign layer2_outputs[12299] = (layer1_outputs[5453]) ^ (layer1_outputs[10388]);
    assign layer2_outputs[12300] = ~((layer1_outputs[9619]) ^ (layer1_outputs[5918]));
    assign layer2_outputs[12301] = ~(layer1_outputs[9531]);
    assign layer2_outputs[12302] = (layer1_outputs[9836]) | (layer1_outputs[4325]);
    assign layer2_outputs[12303] = ~(layer1_outputs[11268]);
    assign layer2_outputs[12304] = layer1_outputs[11430];
    assign layer2_outputs[12305] = (layer1_outputs[9110]) ^ (layer1_outputs[5277]);
    assign layer2_outputs[12306] = layer1_outputs[2785];
    assign layer2_outputs[12307] = layer1_outputs[3280];
    assign layer2_outputs[12308] = ~((layer1_outputs[4767]) ^ (layer1_outputs[2189]));
    assign layer2_outputs[12309] = layer1_outputs[3532];
    assign layer2_outputs[12310] = (layer1_outputs[4177]) ^ (layer1_outputs[11663]);
    assign layer2_outputs[12311] = ~(layer1_outputs[5952]) | (layer1_outputs[2851]);
    assign layer2_outputs[12312] = ~(layer1_outputs[6520]);
    assign layer2_outputs[12313] = layer1_outputs[1837];
    assign layer2_outputs[12314] = ~((layer1_outputs[4428]) ^ (layer1_outputs[2216]));
    assign layer2_outputs[12315] = layer1_outputs[11843];
    assign layer2_outputs[12316] = ~(layer1_outputs[7579]);
    assign layer2_outputs[12317] = ~(layer1_outputs[2378]);
    assign layer2_outputs[12318] = 1'b1;
    assign layer2_outputs[12319] = ~(layer1_outputs[10029]) | (layer1_outputs[1437]);
    assign layer2_outputs[12320] = ~((layer1_outputs[3902]) ^ (layer1_outputs[1629]));
    assign layer2_outputs[12321] = (layer1_outputs[11376]) ^ (layer1_outputs[5783]);
    assign layer2_outputs[12322] = layer1_outputs[3337];
    assign layer2_outputs[12323] = ~(layer1_outputs[12475]) | (layer1_outputs[206]);
    assign layer2_outputs[12324] = ~((layer1_outputs[6544]) | (layer1_outputs[5498]));
    assign layer2_outputs[12325] = (layer1_outputs[11193]) & (layer1_outputs[2293]);
    assign layer2_outputs[12326] = 1'b1;
    assign layer2_outputs[12327] = layer1_outputs[7936];
    assign layer2_outputs[12328] = ~((layer1_outputs[12492]) | (layer1_outputs[2463]));
    assign layer2_outputs[12329] = ~(layer1_outputs[9729]);
    assign layer2_outputs[12330] = ~(layer1_outputs[3812]);
    assign layer2_outputs[12331] = (layer1_outputs[1341]) ^ (layer1_outputs[12527]);
    assign layer2_outputs[12332] = layer1_outputs[10195];
    assign layer2_outputs[12333] = layer1_outputs[11694];
    assign layer2_outputs[12334] = (layer1_outputs[9225]) & ~(layer1_outputs[10479]);
    assign layer2_outputs[12335] = ~(layer1_outputs[8662]);
    assign layer2_outputs[12336] = layer1_outputs[5953];
    assign layer2_outputs[12337] = layer1_outputs[15];
    assign layer2_outputs[12338] = layer1_outputs[1795];
    assign layer2_outputs[12339] = (layer1_outputs[8019]) | (layer1_outputs[3868]);
    assign layer2_outputs[12340] = (layer1_outputs[300]) & (layer1_outputs[8235]);
    assign layer2_outputs[12341] = layer1_outputs[12523];
    assign layer2_outputs[12342] = ~((layer1_outputs[8689]) ^ (layer1_outputs[8202]));
    assign layer2_outputs[12343] = ~(layer1_outputs[6683]) | (layer1_outputs[3009]);
    assign layer2_outputs[12344] = layer1_outputs[1404];
    assign layer2_outputs[12345] = layer1_outputs[8];
    assign layer2_outputs[12346] = ~(layer1_outputs[12313]) | (layer1_outputs[2937]);
    assign layer2_outputs[12347] = ~(layer1_outputs[2837]);
    assign layer2_outputs[12348] = (layer1_outputs[11174]) ^ (layer1_outputs[4589]);
    assign layer2_outputs[12349] = layer1_outputs[1541];
    assign layer2_outputs[12350] = ~((layer1_outputs[6736]) | (layer1_outputs[1411]));
    assign layer2_outputs[12351] = layer1_outputs[6450];
    assign layer2_outputs[12352] = 1'b1;
    assign layer2_outputs[12353] = layer1_outputs[11384];
    assign layer2_outputs[12354] = layer1_outputs[4706];
    assign layer2_outputs[12355] = (layer1_outputs[7229]) ^ (layer1_outputs[11949]);
    assign layer2_outputs[12356] = (layer1_outputs[12645]) ^ (layer1_outputs[8624]);
    assign layer2_outputs[12357] = layer1_outputs[4696];
    assign layer2_outputs[12358] = (layer1_outputs[9484]) & ~(layer1_outputs[7218]);
    assign layer2_outputs[12359] = (layer1_outputs[1455]) & ~(layer1_outputs[279]);
    assign layer2_outputs[12360] = ~(layer1_outputs[6313]) | (layer1_outputs[3036]);
    assign layer2_outputs[12361] = ~(layer1_outputs[4970]) | (layer1_outputs[4984]);
    assign layer2_outputs[12362] = (layer1_outputs[9222]) & (layer1_outputs[11799]);
    assign layer2_outputs[12363] = ~(layer1_outputs[9247]) | (layer1_outputs[11340]);
    assign layer2_outputs[12364] = ~(layer1_outputs[2018]);
    assign layer2_outputs[12365] = layer1_outputs[11284];
    assign layer2_outputs[12366] = (layer1_outputs[3001]) ^ (layer1_outputs[10101]);
    assign layer2_outputs[12367] = layer1_outputs[11323];
    assign layer2_outputs[12368] = ~(layer1_outputs[5699]);
    assign layer2_outputs[12369] = ~((layer1_outputs[6001]) | (layer1_outputs[488]));
    assign layer2_outputs[12370] = ~(layer1_outputs[7207]) | (layer1_outputs[3672]);
    assign layer2_outputs[12371] = (layer1_outputs[752]) ^ (layer1_outputs[12181]);
    assign layer2_outputs[12372] = layer1_outputs[10200];
    assign layer2_outputs[12373] = ~(layer1_outputs[10281]);
    assign layer2_outputs[12374] = ~(layer1_outputs[12084]) | (layer1_outputs[7917]);
    assign layer2_outputs[12375] = ~((layer1_outputs[7078]) | (layer1_outputs[6331]));
    assign layer2_outputs[12376] = ~(layer1_outputs[3033]);
    assign layer2_outputs[12377] = ~(layer1_outputs[3282]);
    assign layer2_outputs[12378] = 1'b1;
    assign layer2_outputs[12379] = layer1_outputs[2898];
    assign layer2_outputs[12380] = ~((layer1_outputs[3116]) ^ (layer1_outputs[1495]));
    assign layer2_outputs[12381] = layer1_outputs[5648];
    assign layer2_outputs[12382] = ~(layer1_outputs[1282]);
    assign layer2_outputs[12383] = ~(layer1_outputs[11658]) | (layer1_outputs[7458]);
    assign layer2_outputs[12384] = (layer1_outputs[1273]) & ~(layer1_outputs[92]);
    assign layer2_outputs[12385] = (layer1_outputs[3109]) ^ (layer1_outputs[6785]);
    assign layer2_outputs[12386] = layer1_outputs[2486];
    assign layer2_outputs[12387] = (layer1_outputs[3261]) & ~(layer1_outputs[8227]);
    assign layer2_outputs[12388] = ~(layer1_outputs[2357]);
    assign layer2_outputs[12389] = ~(layer1_outputs[3979]) | (layer1_outputs[10238]);
    assign layer2_outputs[12390] = (layer1_outputs[5061]) & ~(layer1_outputs[2295]);
    assign layer2_outputs[12391] = layer1_outputs[3556];
    assign layer2_outputs[12392] = ~(layer1_outputs[10579]) | (layer1_outputs[4412]);
    assign layer2_outputs[12393] = (layer1_outputs[10523]) & ~(layer1_outputs[12545]);
    assign layer2_outputs[12394] = ~(layer1_outputs[4233]);
    assign layer2_outputs[12395] = ~(layer1_outputs[1893]);
    assign layer2_outputs[12396] = (layer1_outputs[8493]) ^ (layer1_outputs[816]);
    assign layer2_outputs[12397] = ~(layer1_outputs[1790]);
    assign layer2_outputs[12398] = (layer1_outputs[6118]) ^ (layer1_outputs[5124]);
    assign layer2_outputs[12399] = ~(layer1_outputs[8916]);
    assign layer2_outputs[12400] = ~(layer1_outputs[2992]);
    assign layer2_outputs[12401] = ~(layer1_outputs[3816]);
    assign layer2_outputs[12402] = ~(layer1_outputs[9365]);
    assign layer2_outputs[12403] = (layer1_outputs[4822]) & ~(layer1_outputs[4646]);
    assign layer2_outputs[12404] = ~((layer1_outputs[12764]) | (layer1_outputs[686]));
    assign layer2_outputs[12405] = ~((layer1_outputs[7999]) ^ (layer1_outputs[8832]));
    assign layer2_outputs[12406] = (layer1_outputs[7909]) | (layer1_outputs[8880]);
    assign layer2_outputs[12407] = ~(layer1_outputs[2886]);
    assign layer2_outputs[12408] = layer1_outputs[4135];
    assign layer2_outputs[12409] = (layer1_outputs[547]) | (layer1_outputs[8667]);
    assign layer2_outputs[12410] = ~(layer1_outputs[4819]) | (layer1_outputs[3381]);
    assign layer2_outputs[12411] = ~((layer1_outputs[7338]) | (layer1_outputs[11392]));
    assign layer2_outputs[12412] = (layer1_outputs[632]) & (layer1_outputs[7561]);
    assign layer2_outputs[12413] = layer1_outputs[10426];
    assign layer2_outputs[12414] = layer1_outputs[6606];
    assign layer2_outputs[12415] = layer1_outputs[908];
    assign layer2_outputs[12416] = ~(layer1_outputs[9021]) | (layer1_outputs[7765]);
    assign layer2_outputs[12417] = ~((layer1_outputs[3872]) ^ (layer1_outputs[2487]));
    assign layer2_outputs[12418] = (layer1_outputs[11862]) & ~(layer1_outputs[6393]);
    assign layer2_outputs[12419] = ~(layer1_outputs[7182]);
    assign layer2_outputs[12420] = ~((layer1_outputs[6263]) | (layer1_outputs[10732]));
    assign layer2_outputs[12421] = layer1_outputs[7740];
    assign layer2_outputs[12422] = layer1_outputs[11775];
    assign layer2_outputs[12423] = 1'b1;
    assign layer2_outputs[12424] = ~(layer1_outputs[1958]);
    assign layer2_outputs[12425] = layer1_outputs[7567];
    assign layer2_outputs[12426] = ~(layer1_outputs[12479]) | (layer1_outputs[1035]);
    assign layer2_outputs[12427] = (layer1_outputs[5096]) & ~(layer1_outputs[1363]);
    assign layer2_outputs[12428] = ~(layer1_outputs[6479]);
    assign layer2_outputs[12429] = ~(layer1_outputs[9693]) | (layer1_outputs[5904]);
    assign layer2_outputs[12430] = ~(layer1_outputs[3249]) | (layer1_outputs[7716]);
    assign layer2_outputs[12431] = ~((layer1_outputs[3535]) ^ (layer1_outputs[12666]));
    assign layer2_outputs[12432] = ~(layer1_outputs[139]) | (layer1_outputs[3998]);
    assign layer2_outputs[12433] = ~((layer1_outputs[8733]) ^ (layer1_outputs[10984]));
    assign layer2_outputs[12434] = layer1_outputs[1765];
    assign layer2_outputs[12435] = ~(layer1_outputs[2295]);
    assign layer2_outputs[12436] = ~((layer1_outputs[1066]) ^ (layer1_outputs[4745]));
    assign layer2_outputs[12437] = layer1_outputs[10642];
    assign layer2_outputs[12438] = ~(layer1_outputs[53]);
    assign layer2_outputs[12439] = ~((layer1_outputs[8545]) ^ (layer1_outputs[2202]));
    assign layer2_outputs[12440] = ~(layer1_outputs[880]) | (layer1_outputs[5558]);
    assign layer2_outputs[12441] = ~((layer1_outputs[2371]) | (layer1_outputs[2001]));
    assign layer2_outputs[12442] = (layer1_outputs[4023]) & ~(layer1_outputs[4594]);
    assign layer2_outputs[12443] = (layer1_outputs[6026]) & (layer1_outputs[8221]);
    assign layer2_outputs[12444] = layer1_outputs[7853];
    assign layer2_outputs[12445] = ~(layer1_outputs[11742]) | (layer1_outputs[8426]);
    assign layer2_outputs[12446] = layer1_outputs[1462];
    assign layer2_outputs[12447] = layer1_outputs[3079];
    assign layer2_outputs[12448] = (layer1_outputs[12267]) ^ (layer1_outputs[2600]);
    assign layer2_outputs[12449] = ~((layer1_outputs[7376]) & (layer1_outputs[4894]));
    assign layer2_outputs[12450] = (layer1_outputs[1648]) & ~(layer1_outputs[7556]);
    assign layer2_outputs[12451] = ~(layer1_outputs[7717]);
    assign layer2_outputs[12452] = (layer1_outputs[7575]) & (layer1_outputs[5249]);
    assign layer2_outputs[12453] = layer1_outputs[7431];
    assign layer2_outputs[12454] = ~((layer1_outputs[8981]) ^ (layer1_outputs[7569]));
    assign layer2_outputs[12455] = ~(layer1_outputs[12643]);
    assign layer2_outputs[12456] = ~(layer1_outputs[3493]) | (layer1_outputs[831]);
    assign layer2_outputs[12457] = (layer1_outputs[6798]) ^ (layer1_outputs[2803]);
    assign layer2_outputs[12458] = ~((layer1_outputs[5560]) ^ (layer1_outputs[11812]));
    assign layer2_outputs[12459] = layer1_outputs[10497];
    assign layer2_outputs[12460] = layer1_outputs[10324];
    assign layer2_outputs[12461] = (layer1_outputs[4139]) & ~(layer1_outputs[3895]);
    assign layer2_outputs[12462] = layer1_outputs[9777];
    assign layer2_outputs[12463] = (layer1_outputs[5114]) ^ (layer1_outputs[7181]);
    assign layer2_outputs[12464] = ~((layer1_outputs[3321]) ^ (layer1_outputs[3480]));
    assign layer2_outputs[12465] = 1'b0;
    assign layer2_outputs[12466] = ~(layer1_outputs[4481]);
    assign layer2_outputs[12467] = (layer1_outputs[7260]) & (layer1_outputs[7696]);
    assign layer2_outputs[12468] = (layer1_outputs[9415]) | (layer1_outputs[1928]);
    assign layer2_outputs[12469] = ~(layer1_outputs[1638]);
    assign layer2_outputs[12470] = ~((layer1_outputs[6256]) & (layer1_outputs[9760]));
    assign layer2_outputs[12471] = ~(layer1_outputs[2367]);
    assign layer2_outputs[12472] = layer1_outputs[7644];
    assign layer2_outputs[12473] = ~(layer1_outputs[2271]) | (layer1_outputs[10360]);
    assign layer2_outputs[12474] = layer1_outputs[10654];
    assign layer2_outputs[12475] = layer1_outputs[4882];
    assign layer2_outputs[12476] = ~(layer1_outputs[1138]);
    assign layer2_outputs[12477] = layer1_outputs[6768];
    assign layer2_outputs[12478] = ~(layer1_outputs[10461]) | (layer1_outputs[12101]);
    assign layer2_outputs[12479] = (layer1_outputs[6241]) & ~(layer1_outputs[7589]);
    assign layer2_outputs[12480] = ~(layer1_outputs[2642]) | (layer1_outputs[6181]);
    assign layer2_outputs[12481] = ~((layer1_outputs[5933]) ^ (layer1_outputs[11220]));
    assign layer2_outputs[12482] = (layer1_outputs[7326]) & ~(layer1_outputs[7916]);
    assign layer2_outputs[12483] = layer1_outputs[3136];
    assign layer2_outputs[12484] = ~(layer1_outputs[11910]);
    assign layer2_outputs[12485] = layer1_outputs[3431];
    assign layer2_outputs[12486] = layer1_outputs[5541];
    assign layer2_outputs[12487] = (layer1_outputs[3332]) & (layer1_outputs[3100]);
    assign layer2_outputs[12488] = ~(layer1_outputs[8054]) | (layer1_outputs[459]);
    assign layer2_outputs[12489] = ~((layer1_outputs[2306]) | (layer1_outputs[679]));
    assign layer2_outputs[12490] = layer1_outputs[7672];
    assign layer2_outputs[12491] = (layer1_outputs[5344]) & ~(layer1_outputs[8219]);
    assign layer2_outputs[12492] = (layer1_outputs[540]) & ~(layer1_outputs[5626]);
    assign layer2_outputs[12493] = layer1_outputs[1133];
    assign layer2_outputs[12494] = layer1_outputs[12746];
    assign layer2_outputs[12495] = ~(layer1_outputs[4982]);
    assign layer2_outputs[12496] = (layer1_outputs[384]) & ~(layer1_outputs[1868]);
    assign layer2_outputs[12497] = ~(layer1_outputs[11120]);
    assign layer2_outputs[12498] = (layer1_outputs[844]) | (layer1_outputs[9769]);
    assign layer2_outputs[12499] = ~((layer1_outputs[2333]) & (layer1_outputs[10357]));
    assign layer2_outputs[12500] = ~(layer1_outputs[1112]) | (layer1_outputs[11409]);
    assign layer2_outputs[12501] = (layer1_outputs[2977]) ^ (layer1_outputs[4062]);
    assign layer2_outputs[12502] = (layer1_outputs[11394]) & (layer1_outputs[10860]);
    assign layer2_outputs[12503] = (layer1_outputs[2369]) & ~(layer1_outputs[3323]);
    assign layer2_outputs[12504] = ~(layer1_outputs[10564]);
    assign layer2_outputs[12505] = layer1_outputs[1847];
    assign layer2_outputs[12506] = ~((layer1_outputs[2599]) & (layer1_outputs[1898]));
    assign layer2_outputs[12507] = ~(layer1_outputs[4391]);
    assign layer2_outputs[12508] = ~(layer1_outputs[7499]) | (layer1_outputs[2860]);
    assign layer2_outputs[12509] = layer1_outputs[8046];
    assign layer2_outputs[12510] = ~((layer1_outputs[7557]) & (layer1_outputs[4863]));
    assign layer2_outputs[12511] = ~((layer1_outputs[1028]) ^ (layer1_outputs[9444]));
    assign layer2_outputs[12512] = (layer1_outputs[1849]) & ~(layer1_outputs[11090]);
    assign layer2_outputs[12513] = ~(layer1_outputs[6933]) | (layer1_outputs[4344]);
    assign layer2_outputs[12514] = (layer1_outputs[12013]) ^ (layer1_outputs[11172]);
    assign layer2_outputs[12515] = layer1_outputs[1739];
    assign layer2_outputs[12516] = ~(layer1_outputs[3006]);
    assign layer2_outputs[12517] = ~((layer1_outputs[12094]) & (layer1_outputs[7615]));
    assign layer2_outputs[12518] = layer1_outputs[5108];
    assign layer2_outputs[12519] = layer1_outputs[11330];
    assign layer2_outputs[12520] = ~((layer1_outputs[3032]) & (layer1_outputs[4613]));
    assign layer2_outputs[12521] = (layer1_outputs[3821]) & ~(layer1_outputs[3836]);
    assign layer2_outputs[12522] = ~(layer1_outputs[7953]) | (layer1_outputs[5856]);
    assign layer2_outputs[12523] = ~(layer1_outputs[5812]);
    assign layer2_outputs[12524] = layer1_outputs[11189];
    assign layer2_outputs[12525] = layer1_outputs[2953];
    assign layer2_outputs[12526] = ~(layer1_outputs[9054]) | (layer1_outputs[396]);
    assign layer2_outputs[12527] = ~(layer1_outputs[8437]);
    assign layer2_outputs[12528] = ~(layer1_outputs[5586]) | (layer1_outputs[2387]);
    assign layer2_outputs[12529] = layer1_outputs[989];
    assign layer2_outputs[12530] = ~(layer1_outputs[8957]);
    assign layer2_outputs[12531] = (layer1_outputs[10799]) | (layer1_outputs[9126]);
    assign layer2_outputs[12532] = ~((layer1_outputs[6761]) | (layer1_outputs[8588]));
    assign layer2_outputs[12533] = (layer1_outputs[11669]) & (layer1_outputs[6485]);
    assign layer2_outputs[12534] = ~((layer1_outputs[2984]) & (layer1_outputs[9532]));
    assign layer2_outputs[12535] = (layer1_outputs[108]) ^ (layer1_outputs[8124]);
    assign layer2_outputs[12536] = (layer1_outputs[11951]) | (layer1_outputs[12179]);
    assign layer2_outputs[12537] = ~((layer1_outputs[2918]) | (layer1_outputs[6461]));
    assign layer2_outputs[12538] = layer1_outputs[12004];
    assign layer2_outputs[12539] = ~(layer1_outputs[10873]) | (layer1_outputs[5036]);
    assign layer2_outputs[12540] = (layer1_outputs[11876]) ^ (layer1_outputs[9253]);
    assign layer2_outputs[12541] = (layer1_outputs[11663]) | (layer1_outputs[3659]);
    assign layer2_outputs[12542] = ~(layer1_outputs[8268]);
    assign layer2_outputs[12543] = ~(layer1_outputs[5210]);
    assign layer2_outputs[12544] = ~(layer1_outputs[3943]);
    assign layer2_outputs[12545] = ~((layer1_outputs[12575]) | (layer1_outputs[3172]));
    assign layer2_outputs[12546] = (layer1_outputs[3148]) ^ (layer1_outputs[3856]);
    assign layer2_outputs[12547] = ~(layer1_outputs[6289]);
    assign layer2_outputs[12548] = (layer1_outputs[10973]) & ~(layer1_outputs[7968]);
    assign layer2_outputs[12549] = layer1_outputs[2495];
    assign layer2_outputs[12550] = ~(layer1_outputs[1981]) | (layer1_outputs[1426]);
    assign layer2_outputs[12551] = layer1_outputs[12390];
    assign layer2_outputs[12552] = ~(layer1_outputs[12005]);
    assign layer2_outputs[12553] = ~(layer1_outputs[12312]);
    assign layer2_outputs[12554] = ~(layer1_outputs[10758]) | (layer1_outputs[7829]);
    assign layer2_outputs[12555] = layer1_outputs[8478];
    assign layer2_outputs[12556] = ~(layer1_outputs[10228]);
    assign layer2_outputs[12557] = ~(layer1_outputs[8860]);
    assign layer2_outputs[12558] = (layer1_outputs[3959]) & ~(layer1_outputs[951]);
    assign layer2_outputs[12559] = ~((layer1_outputs[7303]) ^ (layer1_outputs[6908]));
    assign layer2_outputs[12560] = ~((layer1_outputs[3251]) & (layer1_outputs[878]));
    assign layer2_outputs[12561] = (layer1_outputs[11133]) & (layer1_outputs[12220]);
    assign layer2_outputs[12562] = (layer1_outputs[288]) | (layer1_outputs[9934]);
    assign layer2_outputs[12563] = layer1_outputs[10185];
    assign layer2_outputs[12564] = (layer1_outputs[6543]) ^ (layer1_outputs[232]);
    assign layer2_outputs[12565] = layer1_outputs[9604];
    assign layer2_outputs[12566] = ~(layer1_outputs[12634]);
    assign layer2_outputs[12567] = (layer1_outputs[10537]) & ~(layer1_outputs[11327]);
    assign layer2_outputs[12568] = layer1_outputs[469];
    assign layer2_outputs[12569] = (layer1_outputs[1062]) | (layer1_outputs[5406]);
    assign layer2_outputs[12570] = ~((layer1_outputs[2385]) ^ (layer1_outputs[9246]));
    assign layer2_outputs[12571] = layer1_outputs[735];
    assign layer2_outputs[12572] = ~(layer1_outputs[11917]);
    assign layer2_outputs[12573] = (layer1_outputs[872]) & ~(layer1_outputs[6977]);
    assign layer2_outputs[12574] = ~(layer1_outputs[11368]);
    assign layer2_outputs[12575] = ~(layer1_outputs[1085]);
    assign layer2_outputs[12576] = ~((layer1_outputs[383]) & (layer1_outputs[4436]));
    assign layer2_outputs[12577] = (layer1_outputs[3120]) & ~(layer1_outputs[1986]);
    assign layer2_outputs[12578] = layer1_outputs[3926];
    assign layer2_outputs[12579] = ~((layer1_outputs[9085]) & (layer1_outputs[12265]));
    assign layer2_outputs[12580] = ~((layer1_outputs[7942]) & (layer1_outputs[10188]));
    assign layer2_outputs[12581] = (layer1_outputs[11237]) ^ (layer1_outputs[1960]);
    assign layer2_outputs[12582] = ~(layer1_outputs[7652]);
    assign layer2_outputs[12583] = (layer1_outputs[10851]) ^ (layer1_outputs[2005]);
    assign layer2_outputs[12584] = layer1_outputs[10087];
    assign layer2_outputs[12585] = ~(layer1_outputs[6284]);
    assign layer2_outputs[12586] = ~((layer1_outputs[9457]) & (layer1_outputs[6250]));
    assign layer2_outputs[12587] = ~(layer1_outputs[9331]);
    assign layer2_outputs[12588] = ~(layer1_outputs[9737]);
    assign layer2_outputs[12589] = layer1_outputs[3542];
    assign layer2_outputs[12590] = (layer1_outputs[1086]) & ~(layer1_outputs[10995]);
    assign layer2_outputs[12591] = ~((layer1_outputs[4972]) ^ (layer1_outputs[9554]));
    assign layer2_outputs[12592] = ~(layer1_outputs[7890]);
    assign layer2_outputs[12593] = ~(layer1_outputs[8799]);
    assign layer2_outputs[12594] = ~(layer1_outputs[7814]);
    assign layer2_outputs[12595] = (layer1_outputs[463]) ^ (layer1_outputs[11715]);
    assign layer2_outputs[12596] = (layer1_outputs[11601]) & ~(layer1_outputs[9342]);
    assign layer2_outputs[12597] = ~(layer1_outputs[9764]);
    assign layer2_outputs[12598] = layer1_outputs[5586];
    assign layer2_outputs[12599] = ~((layer1_outputs[7982]) ^ (layer1_outputs[1106]));
    assign layer2_outputs[12600] = ~((layer1_outputs[3630]) & (layer1_outputs[8505]));
    assign layer2_outputs[12601] = (layer1_outputs[569]) & (layer1_outputs[2169]);
    assign layer2_outputs[12602] = (layer1_outputs[2532]) ^ (layer1_outputs[12113]);
    assign layer2_outputs[12603] = (layer1_outputs[647]) & ~(layer1_outputs[7788]);
    assign layer2_outputs[12604] = ~(layer1_outputs[11622]);
    assign layer2_outputs[12605] = layer1_outputs[4781];
    assign layer2_outputs[12606] = (layer1_outputs[6412]) ^ (layer1_outputs[2234]);
    assign layer2_outputs[12607] = (layer1_outputs[5170]) ^ (layer1_outputs[12247]);
    assign layer2_outputs[12608] = layer1_outputs[2184];
    assign layer2_outputs[12609] = ~((layer1_outputs[9993]) ^ (layer1_outputs[816]));
    assign layer2_outputs[12610] = ~(layer1_outputs[8594]);
    assign layer2_outputs[12611] = layer1_outputs[1082];
    assign layer2_outputs[12612] = layer1_outputs[1239];
    assign layer2_outputs[12613] = layer1_outputs[12727];
    assign layer2_outputs[12614] = layer1_outputs[5948];
    assign layer2_outputs[12615] = layer1_outputs[804];
    assign layer2_outputs[12616] = ~(layer1_outputs[4874]);
    assign layer2_outputs[12617] = ~(layer1_outputs[9183]);
    assign layer2_outputs[12618] = layer1_outputs[5379];
    assign layer2_outputs[12619] = ~(layer1_outputs[9942]) | (layer1_outputs[2679]);
    assign layer2_outputs[12620] = (layer1_outputs[2606]) & ~(layer1_outputs[48]);
    assign layer2_outputs[12621] = ~(layer1_outputs[10349]);
    assign layer2_outputs[12622] = layer1_outputs[11123];
    assign layer2_outputs[12623] = (layer1_outputs[4842]) ^ (layer1_outputs[11772]);
    assign layer2_outputs[12624] = layer1_outputs[1402];
    assign layer2_outputs[12625] = (layer1_outputs[1888]) ^ (layer1_outputs[12598]);
    assign layer2_outputs[12626] = (layer1_outputs[230]) & ~(layer1_outputs[3702]);
    assign layer2_outputs[12627] = ~((layer1_outputs[9160]) ^ (layer1_outputs[9751]));
    assign layer2_outputs[12628] = layer1_outputs[4335];
    assign layer2_outputs[12629] = layer1_outputs[11739];
    assign layer2_outputs[12630] = ~((layer1_outputs[10994]) ^ (layer1_outputs[12063]));
    assign layer2_outputs[12631] = ~(layer1_outputs[6674]) | (layer1_outputs[2571]);
    assign layer2_outputs[12632] = ~(layer1_outputs[5788]);
    assign layer2_outputs[12633] = ~((layer1_outputs[348]) ^ (layer1_outputs[4778]));
    assign layer2_outputs[12634] = layer1_outputs[9471];
    assign layer2_outputs[12635] = 1'b0;
    assign layer2_outputs[12636] = (layer1_outputs[4171]) & ~(layer1_outputs[2763]);
    assign layer2_outputs[12637] = ~(layer1_outputs[3044]);
    assign layer2_outputs[12638] = (layer1_outputs[9144]) & (layer1_outputs[4716]);
    assign layer2_outputs[12639] = ~(layer1_outputs[230]);
    assign layer2_outputs[12640] = ~(layer1_outputs[5049]) | (layer1_outputs[11959]);
    assign layer2_outputs[12641] = layer1_outputs[5739];
    assign layer2_outputs[12642] = 1'b1;
    assign layer2_outputs[12643] = ~(layer1_outputs[1455]) | (layer1_outputs[3789]);
    assign layer2_outputs[12644] = ~(layer1_outputs[11812]);
    assign layer2_outputs[12645] = ~((layer1_outputs[6094]) & (layer1_outputs[4678]));
    assign layer2_outputs[12646] = ~((layer1_outputs[11355]) & (layer1_outputs[6502]));
    assign layer2_outputs[12647] = (layer1_outputs[6139]) & (layer1_outputs[11528]);
    assign layer2_outputs[12648] = layer1_outputs[6503];
    assign layer2_outputs[12649] = ~(layer1_outputs[6154]);
    assign layer2_outputs[12650] = (layer1_outputs[12567]) & ~(layer1_outputs[475]);
    assign layer2_outputs[12651] = (layer1_outputs[10839]) ^ (layer1_outputs[4087]);
    assign layer2_outputs[12652] = (layer1_outputs[5303]) ^ (layer1_outputs[7207]);
    assign layer2_outputs[12653] = ~(layer1_outputs[2966]) | (layer1_outputs[10526]);
    assign layer2_outputs[12654] = (layer1_outputs[5851]) | (layer1_outputs[5231]);
    assign layer2_outputs[12655] = ~(layer1_outputs[478]) | (layer1_outputs[10107]);
    assign layer2_outputs[12656] = ~((layer1_outputs[1521]) ^ (layer1_outputs[10809]));
    assign layer2_outputs[12657] = (layer1_outputs[8376]) | (layer1_outputs[673]);
    assign layer2_outputs[12658] = layer1_outputs[6263];
    assign layer2_outputs[12659] = (layer1_outputs[9018]) & ~(layer1_outputs[9574]);
    assign layer2_outputs[12660] = ~(layer1_outputs[3911]) | (layer1_outputs[7368]);
    assign layer2_outputs[12661] = ~((layer1_outputs[1431]) | (layer1_outputs[5613]));
    assign layer2_outputs[12662] = ~(layer1_outputs[2240]);
    assign layer2_outputs[12663] = ~((layer1_outputs[5154]) | (layer1_outputs[11147]));
    assign layer2_outputs[12664] = (layer1_outputs[3571]) ^ (layer1_outputs[2208]);
    assign layer2_outputs[12665] = ~(layer1_outputs[8249]) | (layer1_outputs[8403]);
    assign layer2_outputs[12666] = ~((layer1_outputs[2891]) | (layer1_outputs[6602]));
    assign layer2_outputs[12667] = layer1_outputs[9312];
    assign layer2_outputs[12668] = layer1_outputs[4202];
    assign layer2_outputs[12669] = (layer1_outputs[2466]) & (layer1_outputs[2991]);
    assign layer2_outputs[12670] = ~(layer1_outputs[5035]);
    assign layer2_outputs[12671] = (layer1_outputs[9493]) ^ (layer1_outputs[10164]);
    assign layer2_outputs[12672] = (layer1_outputs[1654]) & ~(layer1_outputs[8575]);
    assign layer2_outputs[12673] = layer1_outputs[4670];
    assign layer2_outputs[12674] = layer1_outputs[685];
    assign layer2_outputs[12675] = (layer1_outputs[7186]) ^ (layer1_outputs[5576]);
    assign layer2_outputs[12676] = ~((layer1_outputs[3573]) | (layer1_outputs[2680]));
    assign layer2_outputs[12677] = layer1_outputs[433];
    assign layer2_outputs[12678] = layer1_outputs[12497];
    assign layer2_outputs[12679] = ~(layer1_outputs[2797]) | (layer1_outputs[11636]);
    assign layer2_outputs[12680] = (layer1_outputs[1823]) | (layer1_outputs[7343]);
    assign layer2_outputs[12681] = (layer1_outputs[10257]) & ~(layer1_outputs[11486]);
    assign layer2_outputs[12682] = (layer1_outputs[9079]) & (layer1_outputs[5099]);
    assign layer2_outputs[12683] = (layer1_outputs[3691]) | (layer1_outputs[10584]);
    assign layer2_outputs[12684] = (layer1_outputs[1875]) & ~(layer1_outputs[3580]);
    assign layer2_outputs[12685] = ~(layer1_outputs[12393]);
    assign layer2_outputs[12686] = ~(layer1_outputs[3591]) | (layer1_outputs[9560]);
    assign layer2_outputs[12687] = ~(layer1_outputs[10458]);
    assign layer2_outputs[12688] = (layer1_outputs[8240]) ^ (layer1_outputs[92]);
    assign layer2_outputs[12689] = ~(layer1_outputs[853]);
    assign layer2_outputs[12690] = layer1_outputs[10969];
    assign layer2_outputs[12691] = ~(layer1_outputs[7074]);
    assign layer2_outputs[12692] = ~(layer1_outputs[10340]);
    assign layer2_outputs[12693] = (layer1_outputs[6912]) | (layer1_outputs[8696]);
    assign layer2_outputs[12694] = layer1_outputs[12612];
    assign layer2_outputs[12695] = layer1_outputs[3334];
    assign layer2_outputs[12696] = ~((layer1_outputs[6464]) ^ (layer1_outputs[3453]));
    assign layer2_outputs[12697] = layer1_outputs[10000];
    assign layer2_outputs[12698] = layer1_outputs[7479];
    assign layer2_outputs[12699] = (layer1_outputs[759]) & (layer1_outputs[3017]);
    assign layer2_outputs[12700] = 1'b0;
    assign layer2_outputs[12701] = (layer1_outputs[11160]) & ~(layer1_outputs[6527]);
    assign layer2_outputs[12702] = ~(layer1_outputs[89]);
    assign layer2_outputs[12703] = (layer1_outputs[11126]) & ~(layer1_outputs[4755]);
    assign layer2_outputs[12704] = 1'b0;
    assign layer2_outputs[12705] = layer1_outputs[9867];
    assign layer2_outputs[12706] = (layer1_outputs[736]) & (layer1_outputs[4544]);
    assign layer2_outputs[12707] = (layer1_outputs[11888]) & ~(layer1_outputs[3036]);
    assign layer2_outputs[12708] = layer1_outputs[4776];
    assign layer2_outputs[12709] = layer1_outputs[905];
    assign layer2_outputs[12710] = layer1_outputs[11671];
    assign layer2_outputs[12711] = ~(layer1_outputs[11264]);
    assign layer2_outputs[12712] = (layer1_outputs[8239]) ^ (layer1_outputs[4596]);
    assign layer2_outputs[12713] = layer1_outputs[9889];
    assign layer2_outputs[12714] = layer1_outputs[10111];
    assign layer2_outputs[12715] = ~(layer1_outputs[2008]);
    assign layer2_outputs[12716] = ~(layer1_outputs[7596]) | (layer1_outputs[2981]);
    assign layer2_outputs[12717] = ~((layer1_outputs[227]) & (layer1_outputs[11457]));
    assign layer2_outputs[12718] = ~(layer1_outputs[7633]) | (layer1_outputs[7247]);
    assign layer2_outputs[12719] = ~((layer1_outputs[11679]) & (layer1_outputs[8599]));
    assign layer2_outputs[12720] = ~(layer1_outputs[11914]);
    assign layer2_outputs[12721] = ~(layer1_outputs[11073]);
    assign layer2_outputs[12722] = layer1_outputs[6916];
    assign layer2_outputs[12723] = ~(layer1_outputs[9142]);
    assign layer2_outputs[12724] = (layer1_outputs[8544]) & ~(layer1_outputs[9025]);
    assign layer2_outputs[12725] = layer1_outputs[11604];
    assign layer2_outputs[12726] = (layer1_outputs[7457]) ^ (layer1_outputs[12501]);
    assign layer2_outputs[12727] = layer1_outputs[6893];
    assign layer2_outputs[12728] = layer1_outputs[7150];
    assign layer2_outputs[12729] = ~(layer1_outputs[6529]);
    assign layer2_outputs[12730] = layer1_outputs[2206];
    assign layer2_outputs[12731] = (layer1_outputs[12192]) ^ (layer1_outputs[10633]);
    assign layer2_outputs[12732] = layer1_outputs[6607];
    assign layer2_outputs[12733] = ~((layer1_outputs[4108]) | (layer1_outputs[1879]));
    assign layer2_outputs[12734] = layer1_outputs[9092];
    assign layer2_outputs[12735] = ~(layer1_outputs[9496]);
    assign layer2_outputs[12736] = ~(layer1_outputs[1810]) | (layer1_outputs[2985]);
    assign layer2_outputs[12737] = (layer1_outputs[3008]) ^ (layer1_outputs[11465]);
    assign layer2_outputs[12738] = layer1_outputs[9720];
    assign layer2_outputs[12739] = ~(layer1_outputs[7956]) | (layer1_outputs[368]);
    assign layer2_outputs[12740] = (layer1_outputs[10708]) & ~(layer1_outputs[8583]);
    assign layer2_outputs[12741] = (layer1_outputs[1058]) ^ (layer1_outputs[5058]);
    assign layer2_outputs[12742] = (layer1_outputs[4117]) ^ (layer1_outputs[4302]);
    assign layer2_outputs[12743] = ~(layer1_outputs[11789]);
    assign layer2_outputs[12744] = layer1_outputs[9937];
    assign layer2_outputs[12745] = layer1_outputs[10247];
    assign layer2_outputs[12746] = (layer1_outputs[1540]) & (layer1_outputs[10491]);
    assign layer2_outputs[12747] = ~((layer1_outputs[7085]) ^ (layer1_outputs[4323]));
    assign layer2_outputs[12748] = ~(layer1_outputs[10463]) | (layer1_outputs[9799]);
    assign layer2_outputs[12749] = ~(layer1_outputs[7328]);
    assign layer2_outputs[12750] = layer1_outputs[1523];
    assign layer2_outputs[12751] = 1'b1;
    assign layer2_outputs[12752] = layer1_outputs[1473];
    assign layer2_outputs[12753] = (layer1_outputs[2046]) & ~(layer1_outputs[9091]);
    assign layer2_outputs[12754] = (layer1_outputs[5976]) ^ (layer1_outputs[1921]);
    assign layer2_outputs[12755] = (layer1_outputs[5662]) & ~(layer1_outputs[1304]);
    assign layer2_outputs[12756] = layer1_outputs[8418];
    assign layer2_outputs[12757] = 1'b1;
    assign layer2_outputs[12758] = ~(layer1_outputs[3105]) | (layer1_outputs[10657]);
    assign layer2_outputs[12759] = (layer1_outputs[3940]) & ~(layer1_outputs[10128]);
    assign layer2_outputs[12760] = (layer1_outputs[10154]) | (layer1_outputs[4800]);
    assign layer2_outputs[12761] = (layer1_outputs[9281]) ^ (layer1_outputs[903]);
    assign layer2_outputs[12762] = ~(layer1_outputs[1923]) | (layer1_outputs[6944]);
    assign layer2_outputs[12763] = layer1_outputs[10803];
    assign layer2_outputs[12764] = ~(layer1_outputs[992]);
    assign layer2_outputs[12765] = ~((layer1_outputs[12543]) | (layer1_outputs[5013]));
    assign layer2_outputs[12766] = ~(layer1_outputs[1326]);
    assign layer2_outputs[12767] = layer1_outputs[9060];
    assign layer2_outputs[12768] = ~((layer1_outputs[10973]) | (layer1_outputs[10812]));
    assign layer2_outputs[12769] = layer1_outputs[178];
    assign layer2_outputs[12770] = ~(layer1_outputs[5458]) | (layer1_outputs[1566]);
    assign layer2_outputs[12771] = ~((layer1_outputs[3628]) | (layer1_outputs[4639]));
    assign layer2_outputs[12772] = (layer1_outputs[11229]) ^ (layer1_outputs[9773]);
    assign layer2_outputs[12773] = (layer1_outputs[6620]) | (layer1_outputs[11919]);
    assign layer2_outputs[12774] = ~((layer1_outputs[674]) & (layer1_outputs[1318]));
    assign layer2_outputs[12775] = ~(layer1_outputs[7578]);
    assign layer2_outputs[12776] = layer1_outputs[11824];
    assign layer2_outputs[12777] = ~(layer1_outputs[8987]);
    assign layer2_outputs[12778] = (layer1_outputs[3043]) & ~(layer1_outputs[1036]);
    assign layer2_outputs[12779] = ~((layer1_outputs[12150]) ^ (layer1_outputs[3405]));
    assign layer2_outputs[12780] = (layer1_outputs[8045]) ^ (layer1_outputs[4422]);
    assign layer2_outputs[12781] = (layer1_outputs[7449]) ^ (layer1_outputs[6419]);
    assign layer2_outputs[12782] = (layer1_outputs[9594]) & (layer1_outputs[11141]);
    assign layer2_outputs[12783] = ~((layer1_outputs[11157]) | (layer1_outputs[1701]));
    assign layer2_outputs[12784] = layer1_outputs[11455];
    assign layer2_outputs[12785] = layer1_outputs[479];
    assign layer2_outputs[12786] = ~(layer1_outputs[5311]) | (layer1_outputs[11902]);
    assign layer2_outputs[12787] = (layer1_outputs[8628]) ^ (layer1_outputs[12245]);
    assign layer2_outputs[12788] = ~((layer1_outputs[4161]) ^ (layer1_outputs[5694]));
    assign layer2_outputs[12789] = ~(layer1_outputs[3244]);
    assign layer2_outputs[12790] = ~((layer1_outputs[7249]) & (layer1_outputs[9985]));
    assign layer2_outputs[12791] = ~(layer1_outputs[9527]);
    assign layer2_outputs[12792] = (layer1_outputs[8998]) & (layer1_outputs[11298]);
    assign layer2_outputs[12793] = ~(layer1_outputs[11509]);
    assign layer2_outputs[12794] = ~(layer1_outputs[5500]);
    assign layer2_outputs[12795] = layer1_outputs[2129];
    assign layer2_outputs[12796] = layer1_outputs[10281];
    assign layer2_outputs[12797] = ~((layer1_outputs[10693]) & (layer1_outputs[5774]));
    assign layer2_outputs[12798] = ~((layer1_outputs[8605]) ^ (layer1_outputs[10213]));
    assign layer2_outputs[12799] = (layer1_outputs[4616]) | (layer1_outputs[7352]);
    assign outputs[0] = (layer2_outputs[3241]) & ~(layer2_outputs[40]);
    assign outputs[1] = ~((layer2_outputs[11896]) ^ (layer2_outputs[5388]));
    assign outputs[2] = (layer2_outputs[12741]) ^ (layer2_outputs[4720]);
    assign outputs[3] = ~(layer2_outputs[9654]) | (layer2_outputs[787]);
    assign outputs[4] = (layer2_outputs[7134]) ^ (layer2_outputs[4556]);
    assign outputs[5] = layer2_outputs[1508];
    assign outputs[6] = ~(layer2_outputs[5909]);
    assign outputs[7] = layer2_outputs[12707];
    assign outputs[8] = layer2_outputs[192];
    assign outputs[9] = layer2_outputs[4244];
    assign outputs[10] = ~(layer2_outputs[8345]);
    assign outputs[11] = ~(layer2_outputs[12373]);
    assign outputs[12] = ~(layer2_outputs[5295]) | (layer2_outputs[3894]);
    assign outputs[13] = (layer2_outputs[11018]) ^ (layer2_outputs[3391]);
    assign outputs[14] = layer2_outputs[921];
    assign outputs[15] = (layer2_outputs[12528]) ^ (layer2_outputs[2984]);
    assign outputs[16] = ~(layer2_outputs[10802]);
    assign outputs[17] = layer2_outputs[7337];
    assign outputs[18] = layer2_outputs[8746];
    assign outputs[19] = ~((layer2_outputs[7257]) | (layer2_outputs[12123]));
    assign outputs[20] = ~(layer2_outputs[2053]);
    assign outputs[21] = (layer2_outputs[12135]) & ~(layer2_outputs[10556]);
    assign outputs[22] = (layer2_outputs[6674]) ^ (layer2_outputs[1633]);
    assign outputs[23] = (layer2_outputs[3684]) & (layer2_outputs[10142]);
    assign outputs[24] = (layer2_outputs[671]) | (layer2_outputs[3030]);
    assign outputs[25] = ~(layer2_outputs[11018]);
    assign outputs[26] = layer2_outputs[1171];
    assign outputs[27] = (layer2_outputs[12384]) ^ (layer2_outputs[6870]);
    assign outputs[28] = ~(layer2_outputs[11074]);
    assign outputs[29] = ~(layer2_outputs[4273]);
    assign outputs[30] = ~((layer2_outputs[7397]) ^ (layer2_outputs[10243]));
    assign outputs[31] = (layer2_outputs[6742]) & ~(layer2_outputs[10906]);
    assign outputs[32] = ~(layer2_outputs[11964]);
    assign outputs[33] = ~(layer2_outputs[10954]);
    assign outputs[34] = ~(layer2_outputs[12150]);
    assign outputs[35] = (layer2_outputs[9233]) & ~(layer2_outputs[9256]);
    assign outputs[36] = ~((layer2_outputs[6547]) ^ (layer2_outputs[3808]));
    assign outputs[37] = layer2_outputs[11473];
    assign outputs[38] = ~(layer2_outputs[9081]);
    assign outputs[39] = (layer2_outputs[7205]) & (layer2_outputs[8433]);
    assign outputs[40] = layer2_outputs[5770];
    assign outputs[41] = ~(layer2_outputs[7859]);
    assign outputs[42] = (layer2_outputs[2806]) | (layer2_outputs[7050]);
    assign outputs[43] = layer2_outputs[3237];
    assign outputs[44] = ~(layer2_outputs[12017]);
    assign outputs[45] = ~(layer2_outputs[10537]) | (layer2_outputs[10977]);
    assign outputs[46] = layer2_outputs[8009];
    assign outputs[47] = ~(layer2_outputs[3456]);
    assign outputs[48] = layer2_outputs[8932];
    assign outputs[49] = layer2_outputs[4272];
    assign outputs[50] = layer2_outputs[5572];
    assign outputs[51] = (layer2_outputs[1675]) & (layer2_outputs[9045]);
    assign outputs[52] = ~(layer2_outputs[116]);
    assign outputs[53] = ~(layer2_outputs[10048]);
    assign outputs[54] = (layer2_outputs[3937]) ^ (layer2_outputs[2994]);
    assign outputs[55] = ~((layer2_outputs[10065]) ^ (layer2_outputs[5155]));
    assign outputs[56] = layer2_outputs[6539];
    assign outputs[57] = ~(layer2_outputs[6900]);
    assign outputs[58] = layer2_outputs[2874];
    assign outputs[59] = (layer2_outputs[2786]) ^ (layer2_outputs[540]);
    assign outputs[60] = ~(layer2_outputs[9297]);
    assign outputs[61] = layer2_outputs[7414];
    assign outputs[62] = (layer2_outputs[8491]) & ~(layer2_outputs[7037]);
    assign outputs[63] = ~((layer2_outputs[507]) ^ (layer2_outputs[6996]));
    assign outputs[64] = ~((layer2_outputs[477]) | (layer2_outputs[11495]));
    assign outputs[65] = (layer2_outputs[4224]) & ~(layer2_outputs[4887]);
    assign outputs[66] = layer2_outputs[6769];
    assign outputs[67] = layer2_outputs[961];
    assign outputs[68] = ~((layer2_outputs[1616]) ^ (layer2_outputs[3505]));
    assign outputs[69] = ~(layer2_outputs[4935]);
    assign outputs[70] = ~(layer2_outputs[9874]);
    assign outputs[71] = (layer2_outputs[3463]) | (layer2_outputs[7498]);
    assign outputs[72] = ~((layer2_outputs[3770]) ^ (layer2_outputs[207]));
    assign outputs[73] = ~(layer2_outputs[2040]);
    assign outputs[74] = ~((layer2_outputs[10065]) ^ (layer2_outputs[2134]));
    assign outputs[75] = ~((layer2_outputs[3235]) & (layer2_outputs[11906]));
    assign outputs[76] = (layer2_outputs[6215]) & ~(layer2_outputs[11074]);
    assign outputs[77] = (layer2_outputs[10163]) & ~(layer2_outputs[1720]);
    assign outputs[78] = layer2_outputs[9944];
    assign outputs[79] = (layer2_outputs[8760]) ^ (layer2_outputs[6173]);
    assign outputs[80] = ~(layer2_outputs[30]);
    assign outputs[81] = ~((layer2_outputs[5958]) | (layer2_outputs[12347]));
    assign outputs[82] = layer2_outputs[8443];
    assign outputs[83] = ~((layer2_outputs[1785]) ^ (layer2_outputs[9919]));
    assign outputs[84] = layer2_outputs[10781];
    assign outputs[85] = ~(layer2_outputs[7501]);
    assign outputs[86] = layer2_outputs[708];
    assign outputs[87] = ~((layer2_outputs[5205]) & (layer2_outputs[7545]));
    assign outputs[88] = layer2_outputs[11570];
    assign outputs[89] = ~(layer2_outputs[9842]);
    assign outputs[90] = ~((layer2_outputs[4510]) ^ (layer2_outputs[5340]));
    assign outputs[91] = ~(layer2_outputs[5288]);
    assign outputs[92] = ~(layer2_outputs[9684]);
    assign outputs[93] = ~((layer2_outputs[7306]) ^ (layer2_outputs[9397]));
    assign outputs[94] = ~(layer2_outputs[5773]);
    assign outputs[95] = ~(layer2_outputs[4957]);
    assign outputs[96] = (layer2_outputs[5497]) ^ (layer2_outputs[3393]);
    assign outputs[97] = ~((layer2_outputs[9573]) ^ (layer2_outputs[10858]));
    assign outputs[98] = ~(layer2_outputs[11831]);
    assign outputs[99] = layer2_outputs[2088];
    assign outputs[100] = ~(layer2_outputs[11799]);
    assign outputs[101] = (layer2_outputs[2310]) & ~(layer2_outputs[11090]);
    assign outputs[102] = ~(layer2_outputs[2450]);
    assign outputs[103] = (layer2_outputs[12430]) ^ (layer2_outputs[6329]);
    assign outputs[104] = ~((layer2_outputs[5506]) ^ (layer2_outputs[7677]));
    assign outputs[105] = ~(layer2_outputs[5108]);
    assign outputs[106] = (layer2_outputs[11783]) ^ (layer2_outputs[5017]);
    assign outputs[107] = ~(layer2_outputs[11834]);
    assign outputs[108] = layer2_outputs[5756];
    assign outputs[109] = layer2_outputs[7062];
    assign outputs[110] = layer2_outputs[159];
    assign outputs[111] = ~(layer2_outputs[11712]) | (layer2_outputs[7851]);
    assign outputs[112] = (layer2_outputs[6409]) & ~(layer2_outputs[2006]);
    assign outputs[113] = layer2_outputs[7326];
    assign outputs[114] = (layer2_outputs[1131]) ^ (layer2_outputs[6265]);
    assign outputs[115] = ~(layer2_outputs[8369]);
    assign outputs[116] = ~(layer2_outputs[4957]);
    assign outputs[117] = ~(layer2_outputs[6237]);
    assign outputs[118] = ~(layer2_outputs[12303]);
    assign outputs[119] = layer2_outputs[3697];
    assign outputs[120] = ~((layer2_outputs[9319]) ^ (layer2_outputs[11654]));
    assign outputs[121] = layer2_outputs[11418];
    assign outputs[122] = ~(layer2_outputs[11179]) | (layer2_outputs[6907]);
    assign outputs[123] = layer2_outputs[7482];
    assign outputs[124] = ~((layer2_outputs[7736]) ^ (layer2_outputs[3181]));
    assign outputs[125] = layer2_outputs[9609];
    assign outputs[126] = ~((layer2_outputs[2313]) & (layer2_outputs[3056]));
    assign outputs[127] = ~(layer2_outputs[2081]);
    assign outputs[128] = layer2_outputs[11197];
    assign outputs[129] = ~(layer2_outputs[11391]);
    assign outputs[130] = layer2_outputs[1800];
    assign outputs[131] = ~(layer2_outputs[593]);
    assign outputs[132] = ~(layer2_outputs[2147]);
    assign outputs[133] = layer2_outputs[11214];
    assign outputs[134] = layer2_outputs[1913];
    assign outputs[135] = ~((layer2_outputs[6581]) & (layer2_outputs[11961]));
    assign outputs[136] = ~(layer2_outputs[9130]) | (layer2_outputs[327]);
    assign outputs[137] = ~(layer2_outputs[7935]);
    assign outputs[138] = layer2_outputs[6208];
    assign outputs[139] = ~((layer2_outputs[7488]) ^ (layer2_outputs[7116]));
    assign outputs[140] = (layer2_outputs[8941]) & ~(layer2_outputs[86]);
    assign outputs[141] = layer2_outputs[9858];
    assign outputs[142] = layer2_outputs[11197];
    assign outputs[143] = layer2_outputs[7839];
    assign outputs[144] = ~(layer2_outputs[4637]);
    assign outputs[145] = ~((layer2_outputs[11475]) ^ (layer2_outputs[7229]));
    assign outputs[146] = ~(layer2_outputs[5767]);
    assign outputs[147] = layer2_outputs[8801];
    assign outputs[148] = ~((layer2_outputs[11630]) ^ (layer2_outputs[6371]));
    assign outputs[149] = ~(layer2_outputs[6179]);
    assign outputs[150] = layer2_outputs[126];
    assign outputs[151] = layer2_outputs[3609];
    assign outputs[152] = ~((layer2_outputs[10254]) ^ (layer2_outputs[7070]));
    assign outputs[153] = ~(layer2_outputs[11190]);
    assign outputs[154] = (layer2_outputs[9111]) & ~(layer2_outputs[10023]);
    assign outputs[155] = ~(layer2_outputs[1720]) | (layer2_outputs[6313]);
    assign outputs[156] = ~(layer2_outputs[10229]);
    assign outputs[157] = ~(layer2_outputs[7076]);
    assign outputs[158] = layer2_outputs[3102];
    assign outputs[159] = ~(layer2_outputs[6760]);
    assign outputs[160] = ~(layer2_outputs[10307]);
    assign outputs[161] = layer2_outputs[3731];
    assign outputs[162] = layer2_outputs[3616];
    assign outputs[163] = layer2_outputs[6723];
    assign outputs[164] = layer2_outputs[7118];
    assign outputs[165] = ~(layer2_outputs[12480]);
    assign outputs[166] = layer2_outputs[10703];
    assign outputs[167] = (layer2_outputs[1040]) & ~(layer2_outputs[8059]);
    assign outputs[168] = ~(layer2_outputs[3849]);
    assign outputs[169] = layer2_outputs[11490];
    assign outputs[170] = (layer2_outputs[3552]) ^ (layer2_outputs[9264]);
    assign outputs[171] = layer2_outputs[6231];
    assign outputs[172] = ~(layer2_outputs[8822]);
    assign outputs[173] = ~((layer2_outputs[3492]) ^ (layer2_outputs[7744]));
    assign outputs[174] = (layer2_outputs[3423]) & (layer2_outputs[10267]);
    assign outputs[175] = (layer2_outputs[12422]) & (layer2_outputs[5648]);
    assign outputs[176] = (layer2_outputs[2922]) ^ (layer2_outputs[10695]);
    assign outputs[177] = layer2_outputs[4462];
    assign outputs[178] = ~(layer2_outputs[9727]);
    assign outputs[179] = layer2_outputs[11451];
    assign outputs[180] = layer2_outputs[10133];
    assign outputs[181] = ~((layer2_outputs[3244]) | (layer2_outputs[8678]));
    assign outputs[182] = layer2_outputs[12403];
    assign outputs[183] = (layer2_outputs[5870]) ^ (layer2_outputs[11549]);
    assign outputs[184] = ~(layer2_outputs[6125]);
    assign outputs[185] = layer2_outputs[4234];
    assign outputs[186] = ~(layer2_outputs[2640]);
    assign outputs[187] = ~(layer2_outputs[11276]);
    assign outputs[188] = ~((layer2_outputs[12766]) ^ (layer2_outputs[6022]));
    assign outputs[189] = ~(layer2_outputs[11947]);
    assign outputs[190] = ~(layer2_outputs[7666]);
    assign outputs[191] = ~(layer2_outputs[7173]);
    assign outputs[192] = ~((layer2_outputs[11345]) ^ (layer2_outputs[8537]));
    assign outputs[193] = ~(layer2_outputs[7167]) | (layer2_outputs[3540]);
    assign outputs[194] = layer2_outputs[12184];
    assign outputs[195] = (layer2_outputs[9942]) ^ (layer2_outputs[11176]);
    assign outputs[196] = ~((layer2_outputs[12153]) ^ (layer2_outputs[6354]));
    assign outputs[197] = layer2_outputs[122];
    assign outputs[198] = ~(layer2_outputs[10683]);
    assign outputs[199] = ~((layer2_outputs[5603]) ^ (layer2_outputs[4161]));
    assign outputs[200] = layer2_outputs[1550];
    assign outputs[201] = (layer2_outputs[11988]) | (layer2_outputs[11876]);
    assign outputs[202] = ~(layer2_outputs[4324]);
    assign outputs[203] = ~(layer2_outputs[3597]);
    assign outputs[204] = ~(layer2_outputs[1615]);
    assign outputs[205] = layer2_outputs[12161];
    assign outputs[206] = ~(layer2_outputs[5260]);
    assign outputs[207] = layer2_outputs[715];
    assign outputs[208] = ~(layer2_outputs[10810]);
    assign outputs[209] = ~(layer2_outputs[4993]);
    assign outputs[210] = (layer2_outputs[9688]) & (layer2_outputs[4373]);
    assign outputs[211] = (layer2_outputs[3214]) & ~(layer2_outputs[2739]);
    assign outputs[212] = (layer2_outputs[10916]) & ~(layer2_outputs[6137]);
    assign outputs[213] = (layer2_outputs[2296]) ^ (layer2_outputs[1932]);
    assign outputs[214] = ~(layer2_outputs[3156]);
    assign outputs[215] = ~((layer2_outputs[6922]) ^ (layer2_outputs[2729]));
    assign outputs[216] = ~((layer2_outputs[3862]) ^ (layer2_outputs[9933]));
    assign outputs[217] = (layer2_outputs[8733]) ^ (layer2_outputs[10465]);
    assign outputs[218] = layer2_outputs[10413];
    assign outputs[219] = ~((layer2_outputs[10589]) ^ (layer2_outputs[6698]));
    assign outputs[220] = (layer2_outputs[1746]) & ~(layer2_outputs[186]);
    assign outputs[221] = ~(layer2_outputs[12150]);
    assign outputs[222] = (layer2_outputs[6509]) & ~(layer2_outputs[4882]);
    assign outputs[223] = layer2_outputs[7816];
    assign outputs[224] = (layer2_outputs[8385]) & ~(layer2_outputs[9665]);
    assign outputs[225] = ~(layer2_outputs[11319]);
    assign outputs[226] = ~(layer2_outputs[9268]);
    assign outputs[227] = ~((layer2_outputs[12390]) ^ (layer2_outputs[6636]));
    assign outputs[228] = (layer2_outputs[3598]) ^ (layer2_outputs[8165]);
    assign outputs[229] = layer2_outputs[822];
    assign outputs[230] = ~((layer2_outputs[843]) & (layer2_outputs[1688]));
    assign outputs[231] = ~(layer2_outputs[9137]);
    assign outputs[232] = ~(layer2_outputs[5773]);
    assign outputs[233] = ~(layer2_outputs[2607]);
    assign outputs[234] = (layer2_outputs[8307]) & (layer2_outputs[5517]);
    assign outputs[235] = layer2_outputs[1620];
    assign outputs[236] = (layer2_outputs[7376]) & (layer2_outputs[8711]);
    assign outputs[237] = layer2_outputs[244];
    assign outputs[238] = ~(layer2_outputs[7813]);
    assign outputs[239] = (layer2_outputs[9439]) & (layer2_outputs[10345]);
    assign outputs[240] = layer2_outputs[6877];
    assign outputs[241] = ~(layer2_outputs[8376]);
    assign outputs[242] = (layer2_outputs[11807]) & (layer2_outputs[9488]);
    assign outputs[243] = (layer2_outputs[8067]) & ~(layer2_outputs[7020]);
    assign outputs[244] = layer2_outputs[8611];
    assign outputs[245] = layer2_outputs[10981];
    assign outputs[246] = layer2_outputs[3105];
    assign outputs[247] = layer2_outputs[10439];
    assign outputs[248] = layer2_outputs[11769];
    assign outputs[249] = ~(layer2_outputs[586]);
    assign outputs[250] = layer2_outputs[9922];
    assign outputs[251] = ~(layer2_outputs[2410]);
    assign outputs[252] = ~(layer2_outputs[9459]);
    assign outputs[253] = (layer2_outputs[7681]) ^ (layer2_outputs[6327]);
    assign outputs[254] = (layer2_outputs[2462]) & (layer2_outputs[10890]);
    assign outputs[255] = ~((layer2_outputs[10499]) & (layer2_outputs[3788]));
    assign outputs[256] = (layer2_outputs[5772]) & (layer2_outputs[131]);
    assign outputs[257] = layer2_outputs[5941];
    assign outputs[258] = ~((layer2_outputs[2500]) ^ (layer2_outputs[456]));
    assign outputs[259] = layer2_outputs[4475];
    assign outputs[260] = ~((layer2_outputs[8603]) ^ (layer2_outputs[10805]));
    assign outputs[261] = layer2_outputs[11285];
    assign outputs[262] = (layer2_outputs[9152]) & ~(layer2_outputs[1680]);
    assign outputs[263] = layer2_outputs[638];
    assign outputs[264] = ~((layer2_outputs[5709]) ^ (layer2_outputs[10341]));
    assign outputs[265] = layer2_outputs[10204];
    assign outputs[266] = layer2_outputs[3900];
    assign outputs[267] = ~(layer2_outputs[2747]);
    assign outputs[268] = layer2_outputs[10752];
    assign outputs[269] = ~((layer2_outputs[6672]) | (layer2_outputs[519]));
    assign outputs[270] = ~(layer2_outputs[19]);
    assign outputs[271] = layer2_outputs[10959];
    assign outputs[272] = layer2_outputs[8511];
    assign outputs[273] = layer2_outputs[4155];
    assign outputs[274] = ~((layer2_outputs[3807]) ^ (layer2_outputs[6775]));
    assign outputs[275] = ~(layer2_outputs[7462]);
    assign outputs[276] = (layer2_outputs[6700]) & (layer2_outputs[8360]);
    assign outputs[277] = ~((layer2_outputs[7374]) ^ (layer2_outputs[6459]));
    assign outputs[278] = ~(layer2_outputs[7855]) | (layer2_outputs[3441]);
    assign outputs[279] = ~((layer2_outputs[825]) ^ (layer2_outputs[829]));
    assign outputs[280] = ~(layer2_outputs[1150]);
    assign outputs[281] = ~(layer2_outputs[7565]);
    assign outputs[282] = ~(layer2_outputs[1283]);
    assign outputs[283] = ~(layer2_outputs[10946]);
    assign outputs[284] = ~(layer2_outputs[2634]);
    assign outputs[285] = layer2_outputs[2834];
    assign outputs[286] = ~(layer2_outputs[5672]);
    assign outputs[287] = ~(layer2_outputs[9950]);
    assign outputs[288] = layer2_outputs[10227];
    assign outputs[289] = ~(layer2_outputs[10430]);
    assign outputs[290] = (layer2_outputs[5964]) & (layer2_outputs[3025]);
    assign outputs[291] = layer2_outputs[4227];
    assign outputs[292] = layer2_outputs[3034];
    assign outputs[293] = layer2_outputs[907];
    assign outputs[294] = layer2_outputs[591];
    assign outputs[295] = ~(layer2_outputs[1373]);
    assign outputs[296] = (layer2_outputs[1454]) ^ (layer2_outputs[10551]);
    assign outputs[297] = ~((layer2_outputs[5297]) ^ (layer2_outputs[1019]));
    assign outputs[298] = ~((layer2_outputs[3381]) | (layer2_outputs[5807]));
    assign outputs[299] = ~((layer2_outputs[10383]) ^ (layer2_outputs[9540]));
    assign outputs[300] = layer2_outputs[439];
    assign outputs[301] = ~((layer2_outputs[3374]) ^ (layer2_outputs[8626]));
    assign outputs[302] = layer2_outputs[12259];
    assign outputs[303] = (layer2_outputs[7226]) & (layer2_outputs[8752]);
    assign outputs[304] = layer2_outputs[5196];
    assign outputs[305] = ~(layer2_outputs[6852]);
    assign outputs[306] = ~((layer2_outputs[7575]) ^ (layer2_outputs[12060]));
    assign outputs[307] = ~((layer2_outputs[11599]) ^ (layer2_outputs[10301]));
    assign outputs[308] = ~((layer2_outputs[5881]) & (layer2_outputs[3387]));
    assign outputs[309] = layer2_outputs[2048];
    assign outputs[310] = ~(layer2_outputs[12139]);
    assign outputs[311] = ~(layer2_outputs[5339]);
    assign outputs[312] = (layer2_outputs[10265]) & ~(layer2_outputs[2128]);
    assign outputs[313] = (layer2_outputs[9979]) & (layer2_outputs[2305]);
    assign outputs[314] = layer2_outputs[8502];
    assign outputs[315] = ~(layer2_outputs[7874]);
    assign outputs[316] = layer2_outputs[4082];
    assign outputs[317] = layer2_outputs[4960];
    assign outputs[318] = layer2_outputs[8731];
    assign outputs[319] = ~((layer2_outputs[269]) ^ (layer2_outputs[6218]));
    assign outputs[320] = ~(layer2_outputs[3582]);
    assign outputs[321] = layer2_outputs[7617];
    assign outputs[322] = ~((layer2_outputs[6832]) | (layer2_outputs[3531]));
    assign outputs[323] = layer2_outputs[910];
    assign outputs[324] = ~(layer2_outputs[5172]);
    assign outputs[325] = (layer2_outputs[5057]) ^ (layer2_outputs[9674]);
    assign outputs[326] = (layer2_outputs[3212]) & ~(layer2_outputs[1869]);
    assign outputs[327] = ~(layer2_outputs[8345]);
    assign outputs[328] = ~(layer2_outputs[3141]);
    assign outputs[329] = layer2_outputs[1915];
    assign outputs[330] = ~((layer2_outputs[12740]) ^ (layer2_outputs[9435]));
    assign outputs[331] = layer2_outputs[2188];
    assign outputs[332] = layer2_outputs[2026];
    assign outputs[333] = (layer2_outputs[4672]) ^ (layer2_outputs[6094]);
    assign outputs[334] = layer2_outputs[10481];
    assign outputs[335] = ~((layer2_outputs[2944]) ^ (layer2_outputs[11247]));
    assign outputs[336] = layer2_outputs[9240];
    assign outputs[337] = layer2_outputs[6174];
    assign outputs[338] = (layer2_outputs[4966]) ^ (layer2_outputs[10464]);
    assign outputs[339] = layer2_outputs[3559];
    assign outputs[340] = ~(layer2_outputs[1862]);
    assign outputs[341] = ~(layer2_outputs[11516]) | (layer2_outputs[784]);
    assign outputs[342] = ~((layer2_outputs[3148]) ^ (layer2_outputs[1425]));
    assign outputs[343] = ~(layer2_outputs[3930]);
    assign outputs[344] = (layer2_outputs[10733]) ^ (layer2_outputs[9918]);
    assign outputs[345] = ~(layer2_outputs[2921]) | (layer2_outputs[8806]);
    assign outputs[346] = layer2_outputs[467];
    assign outputs[347] = layer2_outputs[7287];
    assign outputs[348] = ~(layer2_outputs[1383]);
    assign outputs[349] = ~(layer2_outputs[725]);
    assign outputs[350] = ~((layer2_outputs[6807]) ^ (layer2_outputs[11702]));
    assign outputs[351] = ~((layer2_outputs[3837]) & (layer2_outputs[9741]));
    assign outputs[352] = ~((layer2_outputs[1979]) ^ (layer2_outputs[11129]));
    assign outputs[353] = ~(layer2_outputs[7291]);
    assign outputs[354] = ~(layer2_outputs[9906]);
    assign outputs[355] = ~(layer2_outputs[9245]);
    assign outputs[356] = ~((layer2_outputs[12090]) ^ (layer2_outputs[10768]));
    assign outputs[357] = ~(layer2_outputs[2677]);
    assign outputs[358] = layer2_outputs[652];
    assign outputs[359] = ~((layer2_outputs[12091]) ^ (layer2_outputs[11405]));
    assign outputs[360] = ~(layer2_outputs[5915]);
    assign outputs[361] = ~((layer2_outputs[3969]) ^ (layer2_outputs[5284]));
    assign outputs[362] = ~(layer2_outputs[1187]) | (layer2_outputs[6064]);
    assign outputs[363] = (layer2_outputs[7152]) & ~(layer2_outputs[8220]);
    assign outputs[364] = ~((layer2_outputs[10195]) ^ (layer2_outputs[5548]));
    assign outputs[365] = layer2_outputs[10866];
    assign outputs[366] = ~(layer2_outputs[6315]);
    assign outputs[367] = (layer2_outputs[183]) & ~(layer2_outputs[6371]);
    assign outputs[368] = ~((layer2_outputs[10587]) ^ (layer2_outputs[5989]));
    assign outputs[369] = ~(layer2_outputs[1346]);
    assign outputs[370] = layer2_outputs[4029];
    assign outputs[371] = layer2_outputs[9703];
    assign outputs[372] = ~((layer2_outputs[9080]) ^ (layer2_outputs[9777]));
    assign outputs[373] = ~(layer2_outputs[11647]);
    assign outputs[374] = ~(layer2_outputs[7636]);
    assign outputs[375] = ~(layer2_outputs[11598]);
    assign outputs[376] = ~(layer2_outputs[10363]);
    assign outputs[377] = layer2_outputs[5042];
    assign outputs[378] = 1'b0;
    assign outputs[379] = (layer2_outputs[10743]) & (layer2_outputs[4376]);
    assign outputs[380] = ~((layer2_outputs[5355]) | (layer2_outputs[8342]));
    assign outputs[381] = ~((layer2_outputs[8644]) | (layer2_outputs[8285]));
    assign outputs[382] = ~(layer2_outputs[8377]);
    assign outputs[383] = layer2_outputs[7212];
    assign outputs[384] = ~(layer2_outputs[5062]);
    assign outputs[385] = ~((layer2_outputs[1870]) | (layer2_outputs[9594]));
    assign outputs[386] = (layer2_outputs[6121]) & (layer2_outputs[11628]);
    assign outputs[387] = (layer2_outputs[7179]) ^ (layer2_outputs[12035]);
    assign outputs[388] = ~((layer2_outputs[4847]) ^ (layer2_outputs[4073]));
    assign outputs[389] = (layer2_outputs[6443]) & ~(layer2_outputs[10789]);
    assign outputs[390] = layer2_outputs[11196];
    assign outputs[391] = (layer2_outputs[21]) ^ (layer2_outputs[9482]);
    assign outputs[392] = ~(layer2_outputs[5146]);
    assign outputs[393] = (layer2_outputs[12543]) & (layer2_outputs[12579]);
    assign outputs[394] = (layer2_outputs[4843]) ^ (layer2_outputs[1051]);
    assign outputs[395] = layer2_outputs[6443];
    assign outputs[396] = ~((layer2_outputs[11514]) & (layer2_outputs[7838]));
    assign outputs[397] = layer2_outputs[2158];
    assign outputs[398] = layer2_outputs[1891];
    assign outputs[399] = layer2_outputs[9135];
    assign outputs[400] = ~(layer2_outputs[3344]);
    assign outputs[401] = ~((layer2_outputs[4720]) & (layer2_outputs[11345]));
    assign outputs[402] = ~(layer2_outputs[11610]);
    assign outputs[403] = ~(layer2_outputs[12787]);
    assign outputs[404] = ~((layer2_outputs[12162]) ^ (layer2_outputs[9708]));
    assign outputs[405] = (layer2_outputs[79]) ^ (layer2_outputs[10436]);
    assign outputs[406] = ~((layer2_outputs[12386]) ^ (layer2_outputs[5952]));
    assign outputs[407] = ~(layer2_outputs[1473]) | (layer2_outputs[8842]);
    assign outputs[408] = layer2_outputs[8698];
    assign outputs[409] = ~(layer2_outputs[2492]) | (layer2_outputs[10882]);
    assign outputs[410] = ~(layer2_outputs[1678]);
    assign outputs[411] = layer2_outputs[2539];
    assign outputs[412] = layer2_outputs[8947];
    assign outputs[413] = layer2_outputs[1368];
    assign outputs[414] = (layer2_outputs[9345]) & (layer2_outputs[6778]);
    assign outputs[415] = ~((layer2_outputs[12179]) ^ (layer2_outputs[4133]));
    assign outputs[416] = ~(layer2_outputs[8147]);
    assign outputs[417] = ~(layer2_outputs[5541]);
    assign outputs[418] = ~(layer2_outputs[3962]) | (layer2_outputs[701]);
    assign outputs[419] = ~(layer2_outputs[1553]);
    assign outputs[420] = layer2_outputs[5843];
    assign outputs[421] = layer2_outputs[9215];
    assign outputs[422] = ~((layer2_outputs[2334]) ^ (layer2_outputs[63]));
    assign outputs[423] = ~(layer2_outputs[10437]);
    assign outputs[424] = (layer2_outputs[1868]) & ~(layer2_outputs[6402]);
    assign outputs[425] = layer2_outputs[3904];
    assign outputs[426] = ~(layer2_outputs[10239]);
    assign outputs[427] = layer2_outputs[1506];
    assign outputs[428] = layer2_outputs[3102];
    assign outputs[429] = ~(layer2_outputs[212]);
    assign outputs[430] = (layer2_outputs[1317]) ^ (layer2_outputs[10102]);
    assign outputs[431] = ~(layer2_outputs[3155]);
    assign outputs[432] = ~(layer2_outputs[1192]);
    assign outputs[433] = layer2_outputs[2412];
    assign outputs[434] = layer2_outputs[8418];
    assign outputs[435] = ~(layer2_outputs[12251]);
    assign outputs[436] = ~((layer2_outputs[1086]) ^ (layer2_outputs[11918]));
    assign outputs[437] = ~((layer2_outputs[7829]) | (layer2_outputs[12066]));
    assign outputs[438] = ~(layer2_outputs[8262]);
    assign outputs[439] = (layer2_outputs[10403]) & ~(layer2_outputs[6117]);
    assign outputs[440] = (layer2_outputs[9334]) & (layer2_outputs[5018]);
    assign outputs[441] = layer2_outputs[5028];
    assign outputs[442] = layer2_outputs[726];
    assign outputs[443] = ~(layer2_outputs[554]);
    assign outputs[444] = (layer2_outputs[9614]) ^ (layer2_outputs[12063]);
    assign outputs[445] = ~(layer2_outputs[10295]);
    assign outputs[446] = ~((layer2_outputs[10992]) | (layer2_outputs[12357]));
    assign outputs[447] = ~((layer2_outputs[2963]) ^ (layer2_outputs[8038]));
    assign outputs[448] = layer2_outputs[8916];
    assign outputs[449] = ~(layer2_outputs[2156]);
    assign outputs[450] = layer2_outputs[5553];
    assign outputs[451] = layer2_outputs[3649];
    assign outputs[452] = ~((layer2_outputs[103]) ^ (layer2_outputs[9742]));
    assign outputs[453] = ~(layer2_outputs[12556]) | (layer2_outputs[1168]);
    assign outputs[454] = layer2_outputs[7626];
    assign outputs[455] = ~((layer2_outputs[270]) ^ (layer2_outputs[11581]));
    assign outputs[456] = (layer2_outputs[9905]) ^ (layer2_outputs[4732]);
    assign outputs[457] = ~(layer2_outputs[8757]);
    assign outputs[458] = ~((layer2_outputs[1409]) & (layer2_outputs[2303]));
    assign outputs[459] = ~(layer2_outputs[2049]);
    assign outputs[460] = ~((layer2_outputs[443]) ^ (layer2_outputs[4164]));
    assign outputs[461] = layer2_outputs[9413];
    assign outputs[462] = layer2_outputs[5140];
    assign outputs[463] = ~((layer2_outputs[622]) ^ (layer2_outputs[7720]));
    assign outputs[464] = ~(layer2_outputs[8215]);
    assign outputs[465] = layer2_outputs[6431];
    assign outputs[466] = (layer2_outputs[4931]) & ~(layer2_outputs[826]);
    assign outputs[467] = ~((layer2_outputs[8850]) ^ (layer2_outputs[9289]));
    assign outputs[468] = ~(layer2_outputs[9034]);
    assign outputs[469] = layer2_outputs[2705];
    assign outputs[470] = (layer2_outputs[1248]) | (layer2_outputs[74]);
    assign outputs[471] = (layer2_outputs[9438]) & ~(layer2_outputs[10284]);
    assign outputs[472] = ~(layer2_outputs[4039]);
    assign outputs[473] = layer2_outputs[4399];
    assign outputs[474] = layer2_outputs[1391];
    assign outputs[475] = ~(layer2_outputs[2888]);
    assign outputs[476] = layer2_outputs[7920];
    assign outputs[477] = ~((layer2_outputs[10186]) ^ (layer2_outputs[5739]));
    assign outputs[478] = ~(layer2_outputs[5060]);
    assign outputs[479] = layer2_outputs[10244];
    assign outputs[480] = (layer2_outputs[12694]) | (layer2_outputs[6407]);
    assign outputs[481] = (layer2_outputs[2882]) ^ (layer2_outputs[5659]);
    assign outputs[482] = layer2_outputs[1699];
    assign outputs[483] = layer2_outputs[806];
    assign outputs[484] = ~(layer2_outputs[12263]);
    assign outputs[485] = ~((layer2_outputs[12497]) ^ (layer2_outputs[10687]));
    assign outputs[486] = layer2_outputs[9872];
    assign outputs[487] = (layer2_outputs[5845]) ^ (layer2_outputs[11013]);
    assign outputs[488] = ~(layer2_outputs[9678]);
    assign outputs[489] = layer2_outputs[12223];
    assign outputs[490] = ~(layer2_outputs[9280]);
    assign outputs[491] = ~(layer2_outputs[9365]) | (layer2_outputs[9868]);
    assign outputs[492] = ~(layer2_outputs[12589]);
    assign outputs[493] = (layer2_outputs[3025]) & ~(layer2_outputs[1213]);
    assign outputs[494] = ~(layer2_outputs[6894]);
    assign outputs[495] = ~(layer2_outputs[11072]);
    assign outputs[496] = (layer2_outputs[9929]) ^ (layer2_outputs[2334]);
    assign outputs[497] = layer2_outputs[2406];
    assign outputs[498] = ~((layer2_outputs[73]) ^ (layer2_outputs[10345]));
    assign outputs[499] = layer2_outputs[3626];
    assign outputs[500] = (layer2_outputs[11530]) ^ (layer2_outputs[5925]);
    assign outputs[501] = layer2_outputs[4288];
    assign outputs[502] = ~(layer2_outputs[11686]);
    assign outputs[503] = (layer2_outputs[223]) | (layer2_outputs[9051]);
    assign outputs[504] = ~(layer2_outputs[12407]);
    assign outputs[505] = layer2_outputs[8726];
    assign outputs[506] = ~((layer2_outputs[3474]) ^ (layer2_outputs[8042]));
    assign outputs[507] = ~((layer2_outputs[8275]) ^ (layer2_outputs[1896]));
    assign outputs[508] = ~(layer2_outputs[4492]);
    assign outputs[509] = (layer2_outputs[3649]) & ~(layer2_outputs[5413]);
    assign outputs[510] = (layer2_outputs[12133]) ^ (layer2_outputs[9231]);
    assign outputs[511] = (layer2_outputs[5467]) & (layer2_outputs[163]);
    assign outputs[512] = ~(layer2_outputs[3631]);
    assign outputs[513] = (layer2_outputs[11889]) ^ (layer2_outputs[3355]);
    assign outputs[514] = ~((layer2_outputs[1977]) ^ (layer2_outputs[11760]));
    assign outputs[515] = ~(layer2_outputs[7310]);
    assign outputs[516] = (layer2_outputs[7877]) ^ (layer2_outputs[12448]);
    assign outputs[517] = layer2_outputs[8365];
    assign outputs[518] = layer2_outputs[11228];
    assign outputs[519] = ~((layer2_outputs[12064]) ^ (layer2_outputs[10396]));
    assign outputs[520] = layer2_outputs[4060];
    assign outputs[521] = ~(layer2_outputs[2747]);
    assign outputs[522] = ~(layer2_outputs[3349]);
    assign outputs[523] = (layer2_outputs[6272]) & (layer2_outputs[10273]);
    assign outputs[524] = ~(layer2_outputs[496]);
    assign outputs[525] = ~(layer2_outputs[10492]);
    assign outputs[526] = ~(layer2_outputs[7254]) | (layer2_outputs[4894]);
    assign outputs[527] = (layer2_outputs[5653]) & ~(layer2_outputs[9593]);
    assign outputs[528] = layer2_outputs[10961];
    assign outputs[529] = layer2_outputs[616];
    assign outputs[530] = layer2_outputs[10627];
    assign outputs[531] = ~((layer2_outputs[11249]) | (layer2_outputs[9943]));
    assign outputs[532] = (layer2_outputs[2257]) & ~(layer2_outputs[10233]);
    assign outputs[533] = (layer2_outputs[6166]) | (layer2_outputs[395]);
    assign outputs[534] = ~(layer2_outputs[3768]);
    assign outputs[535] = layer2_outputs[1388];
    assign outputs[536] = (layer2_outputs[12590]) ^ (layer2_outputs[11468]);
    assign outputs[537] = ~(layer2_outputs[8738]);
    assign outputs[538] = (layer2_outputs[125]) ^ (layer2_outputs[7734]);
    assign outputs[539] = layer2_outputs[7861];
    assign outputs[540] = (layer2_outputs[6966]) & (layer2_outputs[9909]);
    assign outputs[541] = ~((layer2_outputs[12011]) & (layer2_outputs[4760]));
    assign outputs[542] = ~(layer2_outputs[6455]);
    assign outputs[543] = ~(layer2_outputs[8086]);
    assign outputs[544] = ~(layer2_outputs[1396]) | (layer2_outputs[6436]);
    assign outputs[545] = ~(layer2_outputs[5835]) | (layer2_outputs[11379]);
    assign outputs[546] = ~(layer2_outputs[353]);
    assign outputs[547] = ~(layer2_outputs[3185]);
    assign outputs[548] = (layer2_outputs[31]) ^ (layer2_outputs[9336]);
    assign outputs[549] = layer2_outputs[1507];
    assign outputs[550] = layer2_outputs[258];
    assign outputs[551] = ~(layer2_outputs[4001]) | (layer2_outputs[2388]);
    assign outputs[552] = ~(layer2_outputs[10460]);
    assign outputs[553] = ~(layer2_outputs[5012]);
    assign outputs[554] = layer2_outputs[9765];
    assign outputs[555] = (layer2_outputs[10782]) | (layer2_outputs[5643]);
    assign outputs[556] = ~(layer2_outputs[3163]) | (layer2_outputs[4572]);
    assign outputs[557] = ~(layer2_outputs[837]);
    assign outputs[558] = ~(layer2_outputs[1613]);
    assign outputs[559] = layer2_outputs[6183];
    assign outputs[560] = ~(layer2_outputs[10620]);
    assign outputs[561] = ~(layer2_outputs[1534]);
    assign outputs[562] = layer2_outputs[465];
    assign outputs[563] = (layer2_outputs[6480]) & ~(layer2_outputs[562]);
    assign outputs[564] = layer2_outputs[4127];
    assign outputs[565] = (layer2_outputs[1599]) & ~(layer2_outputs[9864]);
    assign outputs[566] = ~(layer2_outputs[5742]) | (layer2_outputs[12316]);
    assign outputs[567] = ~((layer2_outputs[426]) ^ (layer2_outputs[11826]));
    assign outputs[568] = layer2_outputs[3010];
    assign outputs[569] = ~(layer2_outputs[1754]);
    assign outputs[570] = (layer2_outputs[4180]) ^ (layer2_outputs[2096]);
    assign outputs[571] = ~(layer2_outputs[1797]);
    assign outputs[572] = ~(layer2_outputs[8287]);
    assign outputs[573] = (layer2_outputs[10493]) & ~(layer2_outputs[4156]);
    assign outputs[574] = ~(layer2_outputs[3916]) | (layer2_outputs[9129]);
    assign outputs[575] = (layer2_outputs[5052]) ^ (layer2_outputs[2776]);
    assign outputs[576] = ~(layer2_outputs[6173]) | (layer2_outputs[8022]);
    assign outputs[577] = layer2_outputs[11196];
    assign outputs[578] = layer2_outputs[9832];
    assign outputs[579] = (layer2_outputs[10378]) ^ (layer2_outputs[10570]);
    assign outputs[580] = ~(layer2_outputs[10027]);
    assign outputs[581] = ~(layer2_outputs[6611]);
    assign outputs[582] = ~(layer2_outputs[11226]);
    assign outputs[583] = (layer2_outputs[3751]) ^ (layer2_outputs[4793]);
    assign outputs[584] = ~(layer2_outputs[10636]);
    assign outputs[585] = ~(layer2_outputs[6422]);
    assign outputs[586] = (layer2_outputs[7645]) | (layer2_outputs[10385]);
    assign outputs[587] = layer2_outputs[6282];
    assign outputs[588] = layer2_outputs[4833];
    assign outputs[589] = ~(layer2_outputs[4905]);
    assign outputs[590] = ~(layer2_outputs[11865]);
    assign outputs[591] = ~(layer2_outputs[3748]);
    assign outputs[592] = ~((layer2_outputs[7199]) & (layer2_outputs[10321]));
    assign outputs[593] = ~((layer2_outputs[2778]) ^ (layer2_outputs[8193]));
    assign outputs[594] = ~(layer2_outputs[3204]) | (layer2_outputs[6073]);
    assign outputs[595] = layer2_outputs[10273];
    assign outputs[596] = (layer2_outputs[3079]) | (layer2_outputs[5439]);
    assign outputs[597] = (layer2_outputs[11480]) & ~(layer2_outputs[3018]);
    assign outputs[598] = ~(layer2_outputs[5814]) | (layer2_outputs[3101]);
    assign outputs[599] = ~(layer2_outputs[5846]);
    assign outputs[600] = ~(layer2_outputs[7027]);
    assign outputs[601] = ~(layer2_outputs[1627]) | (layer2_outputs[5196]);
    assign outputs[602] = layer2_outputs[7683];
    assign outputs[603] = (layer2_outputs[6926]) ^ (layer2_outputs[3270]);
    assign outputs[604] = ~((layer2_outputs[7316]) ^ (layer2_outputs[3150]));
    assign outputs[605] = (layer2_outputs[9849]) & ~(layer2_outputs[6209]);
    assign outputs[606] = layer2_outputs[2478];
    assign outputs[607] = (layer2_outputs[667]) ^ (layer2_outputs[7629]);
    assign outputs[608] = ~(layer2_outputs[8970]);
    assign outputs[609] = layer2_outputs[11128];
    assign outputs[610] = layer2_outputs[12023];
    assign outputs[611] = layer2_outputs[8403];
    assign outputs[612] = (layer2_outputs[21]) & ~(layer2_outputs[1143]);
    assign outputs[613] = ~(layer2_outputs[1264]);
    assign outputs[614] = ~(layer2_outputs[11237]);
    assign outputs[615] = layer2_outputs[9170];
    assign outputs[616] = (layer2_outputs[6925]) & ~(layer2_outputs[9562]);
    assign outputs[617] = ~(layer2_outputs[5504]);
    assign outputs[618] = layer2_outputs[6415];
    assign outputs[619] = layer2_outputs[10488];
    assign outputs[620] = ~((layer2_outputs[4896]) ^ (layer2_outputs[5916]));
    assign outputs[621] = ~((layer2_outputs[2397]) ^ (layer2_outputs[2716]));
    assign outputs[622] = ~((layer2_outputs[5417]) ^ (layer2_outputs[9582]));
    assign outputs[623] = (layer2_outputs[6669]) ^ (layer2_outputs[5826]);
    assign outputs[624] = ~((layer2_outputs[4055]) ^ (layer2_outputs[4968]));
    assign outputs[625] = ~((layer2_outputs[5375]) ^ (layer2_outputs[11650]));
    assign outputs[626] = layer2_outputs[5988];
    assign outputs[627] = ~(layer2_outputs[12035]);
    assign outputs[628] = (layer2_outputs[10953]) ^ (layer2_outputs[495]);
    assign outputs[629] = ~(layer2_outputs[7502]);
    assign outputs[630] = layer2_outputs[10515];
    assign outputs[631] = ~(layer2_outputs[9706]);
    assign outputs[632] = layer2_outputs[8375];
    assign outputs[633] = ~(layer2_outputs[10389]);
    assign outputs[634] = ~((layer2_outputs[6400]) & (layer2_outputs[12125]));
    assign outputs[635] = ~(layer2_outputs[132]);
    assign outputs[636] = ~(layer2_outputs[1180]) | (layer2_outputs[93]);
    assign outputs[637] = layer2_outputs[1935];
    assign outputs[638] = layer2_outputs[3910];
    assign outputs[639] = ~(layer2_outputs[2948]);
    assign outputs[640] = (layer2_outputs[10525]) & ~(layer2_outputs[6146]);
    assign outputs[641] = ~((layer2_outputs[3785]) & (layer2_outputs[4573]));
    assign outputs[642] = ~(layer2_outputs[2246]);
    assign outputs[643] = layer2_outputs[9318];
    assign outputs[644] = ~(layer2_outputs[6011]);
    assign outputs[645] = layer2_outputs[11988];
    assign outputs[646] = layer2_outputs[2749];
    assign outputs[647] = layer2_outputs[3441];
    assign outputs[648] = ~(layer2_outputs[12738]) | (layer2_outputs[6466]);
    assign outputs[649] = ~(layer2_outputs[6558]);
    assign outputs[650] = ~(layer2_outputs[3062]);
    assign outputs[651] = layer2_outputs[7285];
    assign outputs[652] = layer2_outputs[10005];
    assign outputs[653] = ~(layer2_outputs[1680]);
    assign outputs[654] = (layer2_outputs[99]) & ~(layer2_outputs[12496]);
    assign outputs[655] = layer2_outputs[2874];
    assign outputs[656] = (layer2_outputs[9673]) | (layer2_outputs[5675]);
    assign outputs[657] = ~((layer2_outputs[10030]) ^ (layer2_outputs[3912]));
    assign outputs[658] = (layer2_outputs[2266]) & ~(layer2_outputs[5617]);
    assign outputs[659] = ~(layer2_outputs[6849]);
    assign outputs[660] = ~((layer2_outputs[6765]) ^ (layer2_outputs[10803]));
    assign outputs[661] = ~(layer2_outputs[6575]);
    assign outputs[662] = ~(layer2_outputs[5991]);
    assign outputs[663] = layer2_outputs[8316];
    assign outputs[664] = ~((layer2_outputs[8782]) | (layer2_outputs[935]));
    assign outputs[665] = ~(layer2_outputs[7828]);
    assign outputs[666] = layer2_outputs[3528];
    assign outputs[667] = ~((layer2_outputs[5286]) | (layer2_outputs[1095]));
    assign outputs[668] = ~(layer2_outputs[12763]);
    assign outputs[669] = ~(layer2_outputs[2292]);
    assign outputs[670] = ~((layer2_outputs[11437]) | (layer2_outputs[8018]));
    assign outputs[671] = ~((layer2_outputs[3882]) ^ (layer2_outputs[4667]));
    assign outputs[672] = layer2_outputs[3604];
    assign outputs[673] = (layer2_outputs[10520]) ^ (layer2_outputs[11259]);
    assign outputs[674] = ~(layer2_outputs[6612]);
    assign outputs[675] = layer2_outputs[5799];
    assign outputs[676] = layer2_outputs[8641];
    assign outputs[677] = ~(layer2_outputs[1956]);
    assign outputs[678] = layer2_outputs[3729];
    assign outputs[679] = (layer2_outputs[5660]) & ~(layer2_outputs[1053]);
    assign outputs[680] = ~((layer2_outputs[3211]) ^ (layer2_outputs[6985]));
    assign outputs[681] = layer2_outputs[6283];
    assign outputs[682] = ~((layer2_outputs[7786]) & (layer2_outputs[10387]));
    assign outputs[683] = ~(layer2_outputs[5963]);
    assign outputs[684] = (layer2_outputs[9497]) & ~(layer2_outputs[9741]);
    assign outputs[685] = (layer2_outputs[3674]) & ~(layer2_outputs[12696]);
    assign outputs[686] = (layer2_outputs[7771]) | (layer2_outputs[1558]);
    assign outputs[687] = (layer2_outputs[11729]) & (layer2_outputs[7247]);
    assign outputs[688] = ~(layer2_outputs[2147]);
    assign outputs[689] = layer2_outputs[2036];
    assign outputs[690] = layer2_outputs[8006];
    assign outputs[691] = layer2_outputs[12204];
    assign outputs[692] = ~((layer2_outputs[10553]) ^ (layer2_outputs[3308]));
    assign outputs[693] = ~(layer2_outputs[5406]);
    assign outputs[694] = ~(layer2_outputs[11552]);
    assign outputs[695] = ~(layer2_outputs[379]) | (layer2_outputs[3536]);
    assign outputs[696] = ~((layer2_outputs[3478]) | (layer2_outputs[8531]));
    assign outputs[697] = ~(layer2_outputs[927]);
    assign outputs[698] = ~(layer2_outputs[8911]);
    assign outputs[699] = ~(layer2_outputs[458]);
    assign outputs[700] = layer2_outputs[27];
    assign outputs[701] = ~((layer2_outputs[10209]) ^ (layer2_outputs[3005]));
    assign outputs[702] = layer2_outputs[4215];
    assign outputs[703] = layer2_outputs[8029];
    assign outputs[704] = ~(layer2_outputs[3314]);
    assign outputs[705] = ~(layer2_outputs[5188]);
    assign outputs[706] = ~((layer2_outputs[9265]) ^ (layer2_outputs[6379]));
    assign outputs[707] = ~(layer2_outputs[9231]);
    assign outputs[708] = ~(layer2_outputs[12605]);
    assign outputs[709] = (layer2_outputs[4824]) ^ (layer2_outputs[11559]);
    assign outputs[710] = ~(layer2_outputs[3732]);
    assign outputs[711] = ~((layer2_outputs[1581]) | (layer2_outputs[355]));
    assign outputs[712] = (layer2_outputs[2062]) ^ (layer2_outputs[4379]);
    assign outputs[713] = layer2_outputs[961];
    assign outputs[714] = layer2_outputs[656];
    assign outputs[715] = ~(layer2_outputs[1966]);
    assign outputs[716] = ~(layer2_outputs[12069]);
    assign outputs[717] = ~((layer2_outputs[8462]) ^ (layer2_outputs[6791]));
    assign outputs[718] = ~(layer2_outputs[7061]);
    assign outputs[719] = layer2_outputs[520];
    assign outputs[720] = ~((layer2_outputs[11218]) ^ (layer2_outputs[153]));
    assign outputs[721] = ~((layer2_outputs[2853]) ^ (layer2_outputs[3702]));
    assign outputs[722] = layer2_outputs[8706];
    assign outputs[723] = layer2_outputs[12213];
    assign outputs[724] = (layer2_outputs[5974]) ^ (layer2_outputs[4424]);
    assign outputs[725] = (layer2_outputs[10121]) & ~(layer2_outputs[9816]);
    assign outputs[726] = (layer2_outputs[10746]) ^ (layer2_outputs[4816]);
    assign outputs[727] = (layer2_outputs[5247]) ^ (layer2_outputs[710]);
    assign outputs[728] = layer2_outputs[7234];
    assign outputs[729] = layer2_outputs[11008];
    assign outputs[730] = ~(layer2_outputs[1277]);
    assign outputs[731] = ~(layer2_outputs[12268]);
    assign outputs[732] = (layer2_outputs[10783]) | (layer2_outputs[364]);
    assign outputs[733] = ~(layer2_outputs[3732]);
    assign outputs[734] = ~(layer2_outputs[12106]) | (layer2_outputs[7294]);
    assign outputs[735] = ~(layer2_outputs[3307]);
    assign outputs[736] = layer2_outputs[4695];
    assign outputs[737] = ~(layer2_outputs[2932]);
    assign outputs[738] = (layer2_outputs[6003]) | (layer2_outputs[7144]);
    assign outputs[739] = ~((layer2_outputs[5574]) ^ (layer2_outputs[3971]));
    assign outputs[740] = layer2_outputs[5137];
    assign outputs[741] = layer2_outputs[8929];
    assign outputs[742] = layer2_outputs[5920];
    assign outputs[743] = layer2_outputs[5704];
    assign outputs[744] = layer2_outputs[10651];
    assign outputs[745] = ~(layer2_outputs[1682]);
    assign outputs[746] = ~((layer2_outputs[8889]) ^ (layer2_outputs[9100]));
    assign outputs[747] = ~(layer2_outputs[3564]);
    assign outputs[748] = ~(layer2_outputs[2508]);
    assign outputs[749] = ~(layer2_outputs[10970]);
    assign outputs[750] = ~((layer2_outputs[8066]) & (layer2_outputs[4548]));
    assign outputs[751] = layer2_outputs[2585];
    assign outputs[752] = layer2_outputs[11465];
    assign outputs[753] = (layer2_outputs[5621]) | (layer2_outputs[570]);
    assign outputs[754] = ~((layer2_outputs[3255]) & (layer2_outputs[11993]));
    assign outputs[755] = (layer2_outputs[10814]) & (layer2_outputs[9374]);
    assign outputs[756] = layer2_outputs[5149];
    assign outputs[757] = layer2_outputs[9519];
    assign outputs[758] = layer2_outputs[2860];
    assign outputs[759] = (layer2_outputs[3709]) & ~(layer2_outputs[1166]);
    assign outputs[760] = ~(layer2_outputs[7850]);
    assign outputs[761] = layer2_outputs[4804];
    assign outputs[762] = layer2_outputs[2998];
    assign outputs[763] = (layer2_outputs[5477]) ^ (layer2_outputs[1893]);
    assign outputs[764] = ~((layer2_outputs[2010]) ^ (layer2_outputs[3341]));
    assign outputs[765] = (layer2_outputs[2460]) ^ (layer2_outputs[6224]);
    assign outputs[766] = ~(layer2_outputs[9201]);
    assign outputs[767] = layer2_outputs[8080];
    assign outputs[768] = ~(layer2_outputs[12607]);
    assign outputs[769] = (layer2_outputs[4026]) ^ (layer2_outputs[8020]);
    assign outputs[770] = ~((layer2_outputs[8735]) ^ (layer2_outputs[7335]));
    assign outputs[771] = (layer2_outputs[1850]) & ~(layer2_outputs[6686]);
    assign outputs[772] = ~((layer2_outputs[7180]) ^ (layer2_outputs[7710]));
    assign outputs[773] = layer2_outputs[9916];
    assign outputs[774] = ~(layer2_outputs[10976]);
    assign outputs[775] = (layer2_outputs[5682]) & ~(layer2_outputs[1425]);
    assign outputs[776] = layer2_outputs[11629];
    assign outputs[777] = layer2_outputs[9894];
    assign outputs[778] = ~(layer2_outputs[9355]);
    assign outputs[779] = ~((layer2_outputs[10039]) ^ (layer2_outputs[8888]));
    assign outputs[780] = (layer2_outputs[12330]) & ~(layer2_outputs[2943]);
    assign outputs[781] = (layer2_outputs[11867]) & (layer2_outputs[9863]);
    assign outputs[782] = ~((layer2_outputs[8107]) ^ (layer2_outputs[2047]));
    assign outputs[783] = ~((layer2_outputs[3952]) ^ (layer2_outputs[4215]));
    assign outputs[784] = ~((layer2_outputs[7789]) ^ (layer2_outputs[50]));
    assign outputs[785] = ~(layer2_outputs[205]);
    assign outputs[786] = ~(layer2_outputs[11009]) | (layer2_outputs[9908]);
    assign outputs[787] = layer2_outputs[9046];
    assign outputs[788] = ~((layer2_outputs[8628]) ^ (layer2_outputs[5002]));
    assign outputs[789] = ~(layer2_outputs[9587]);
    assign outputs[790] = ~(layer2_outputs[11069]) | (layer2_outputs[10084]);
    assign outputs[791] = ~(layer2_outputs[11189]) | (layer2_outputs[3638]);
    assign outputs[792] = (layer2_outputs[12307]) ^ (layer2_outputs[2303]);
    assign outputs[793] = layer2_outputs[2998];
    assign outputs[794] = (layer2_outputs[9272]) | (layer2_outputs[4860]);
    assign outputs[795] = (layer2_outputs[10703]) | (layer2_outputs[2243]);
    assign outputs[796] = ~((layer2_outputs[2383]) | (layer2_outputs[7016]));
    assign outputs[797] = ~((layer2_outputs[3428]) ^ (layer2_outputs[11846]));
    assign outputs[798] = ~(layer2_outputs[2503]) | (layer2_outputs[7528]);
    assign outputs[799] = (layer2_outputs[2624]) | (layer2_outputs[1285]);
    assign outputs[800] = layer2_outputs[1604];
    assign outputs[801] = (layer2_outputs[2437]) | (layer2_outputs[12329]);
    assign outputs[802] = (layer2_outputs[4240]) | (layer2_outputs[1610]);
    assign outputs[803] = ~(layer2_outputs[9992]);
    assign outputs[804] = layer2_outputs[11958];
    assign outputs[805] = layer2_outputs[198];
    assign outputs[806] = (layer2_outputs[6659]) ^ (layer2_outputs[10010]);
    assign outputs[807] = ~(layer2_outputs[12159]);
    assign outputs[808] = (layer2_outputs[6941]) ^ (layer2_outputs[5366]);
    assign outputs[809] = (layer2_outputs[4120]) & (layer2_outputs[924]);
    assign outputs[810] = (layer2_outputs[8300]) & ~(layer2_outputs[11254]);
    assign outputs[811] = ~((layer2_outputs[11375]) ^ (layer2_outputs[9569]));
    assign outputs[812] = ~(layer2_outputs[3711]);
    assign outputs[813] = (layer2_outputs[3285]) & ~(layer2_outputs[6750]);
    assign outputs[814] = ~((layer2_outputs[5364]) ^ (layer2_outputs[12369]));
    assign outputs[815] = (layer2_outputs[11777]) ^ (layer2_outputs[11691]);
    assign outputs[816] = ~((layer2_outputs[9131]) ^ (layer2_outputs[10322]));
    assign outputs[817] = layer2_outputs[8457];
    assign outputs[818] = ~(layer2_outputs[10373]);
    assign outputs[819] = (layer2_outputs[1559]) & ~(layer2_outputs[3677]);
    assign outputs[820] = ~(layer2_outputs[960]);
    assign outputs[821] = ~(layer2_outputs[12178]);
    assign outputs[822] = ~((layer2_outputs[2357]) ^ (layer2_outputs[6666]));
    assign outputs[823] = (layer2_outputs[9299]) ^ (layer2_outputs[10033]);
    assign outputs[824] = layer2_outputs[1221];
    assign outputs[825] = (layer2_outputs[3764]) ^ (layer2_outputs[9247]);
    assign outputs[826] = (layer2_outputs[7745]) ^ (layer2_outputs[3001]);
    assign outputs[827] = ~((layer2_outputs[5635]) | (layer2_outputs[276]));
    assign outputs[828] = (layer2_outputs[5402]) ^ (layer2_outputs[8304]);
    assign outputs[829] = ~(layer2_outputs[8207]);
    assign outputs[830] = ~(layer2_outputs[2089]);
    assign outputs[831] = ~(layer2_outputs[796]);
    assign outputs[832] = (layer2_outputs[8055]) ^ (layer2_outputs[637]);
    assign outputs[833] = (layer2_outputs[6883]) & ~(layer2_outputs[10565]);
    assign outputs[834] = (layer2_outputs[2449]) & ~(layer2_outputs[1050]);
    assign outputs[835] = layer2_outputs[9290];
    assign outputs[836] = ~((layer2_outputs[3051]) ^ (layer2_outputs[7481]));
    assign outputs[837] = layer2_outputs[5213];
    assign outputs[838] = ~(layer2_outputs[12367]);
    assign outputs[839] = layer2_outputs[12223];
    assign outputs[840] = layer2_outputs[12172];
    assign outputs[841] = (layer2_outputs[2435]) ^ (layer2_outputs[2058]);
    assign outputs[842] = layer2_outputs[7484];
    assign outputs[843] = layer2_outputs[11942];
    assign outputs[844] = ~((layer2_outputs[5879]) | (layer2_outputs[11650]));
    assign outputs[845] = layer2_outputs[1809];
    assign outputs[846] = ~(layer2_outputs[5688]);
    assign outputs[847] = (layer2_outputs[7645]) & ~(layer2_outputs[6658]);
    assign outputs[848] = ~(layer2_outputs[382]);
    assign outputs[849] = ~((layer2_outputs[1930]) & (layer2_outputs[3575]));
    assign outputs[850] = ~(layer2_outputs[11448]);
    assign outputs[851] = ~((layer2_outputs[2508]) ^ (layer2_outputs[11104]));
    assign outputs[852] = ~(layer2_outputs[2094]);
    assign outputs[853] = ~((layer2_outputs[2802]) ^ (layer2_outputs[8225]));
    assign outputs[854] = ~(layer2_outputs[9864]);
    assign outputs[855] = layer2_outputs[2827];
    assign outputs[856] = (layer2_outputs[9676]) & (layer2_outputs[8179]);
    assign outputs[857] = layer2_outputs[11388];
    assign outputs[858] = ~((layer2_outputs[10172]) ^ (layer2_outputs[10151]));
    assign outputs[859] = layer2_outputs[12204];
    assign outputs[860] = layer2_outputs[3644];
    assign outputs[861] = ~(layer2_outputs[2946]);
    assign outputs[862] = ~(layer2_outputs[3014]);
    assign outputs[863] = ~(layer2_outputs[67]);
    assign outputs[864] = ~(layer2_outputs[3228]);
    assign outputs[865] = ~(layer2_outputs[5358]);
    assign outputs[866] = layer2_outputs[3489];
    assign outputs[867] = ~(layer2_outputs[1141]);
    assign outputs[868] = layer2_outputs[9190];
    assign outputs[869] = (layer2_outputs[4519]) ^ (layer2_outputs[11534]);
    assign outputs[870] = (layer2_outputs[10639]) ^ (layer2_outputs[7247]);
    assign outputs[871] = ~(layer2_outputs[896]);
    assign outputs[872] = layer2_outputs[9127];
    assign outputs[873] = (layer2_outputs[4077]) ^ (layer2_outputs[8781]);
    assign outputs[874] = ~((layer2_outputs[1012]) ^ (layer2_outputs[6481]));
    assign outputs[875] = ~((layer2_outputs[11342]) ^ (layer2_outputs[2326]));
    assign outputs[876] = layer2_outputs[1599];
    assign outputs[877] = (layer2_outputs[234]) | (layer2_outputs[2767]);
    assign outputs[878] = layer2_outputs[3558];
    assign outputs[879] = layer2_outputs[2562];
    assign outputs[880] = ~((layer2_outputs[7004]) ^ (layer2_outputs[3685]));
    assign outputs[881] = layer2_outputs[5953];
    assign outputs[882] = ~(layer2_outputs[809]);
    assign outputs[883] = layer2_outputs[11990];
    assign outputs[884] = ~(layer2_outputs[8136]);
    assign outputs[885] = ~(layer2_outputs[11312]);
    assign outputs[886] = ~(layer2_outputs[11122]);
    assign outputs[887] = layer2_outputs[8448];
    assign outputs[888] = ~((layer2_outputs[5201]) | (layer2_outputs[11377]));
    assign outputs[889] = ~((layer2_outputs[7345]) ^ (layer2_outputs[1858]));
    assign outputs[890] = ~(layer2_outputs[3026]);
    assign outputs[891] = layer2_outputs[4294];
    assign outputs[892] = ~(layer2_outputs[8965]);
    assign outputs[893] = ~((layer2_outputs[2500]) ^ (layer2_outputs[8521]));
    assign outputs[894] = ~((layer2_outputs[12592]) ^ (layer2_outputs[1376]));
    assign outputs[895] = layer2_outputs[8241];
    assign outputs[896] = (layer2_outputs[7430]) & ~(layer2_outputs[4370]);
    assign outputs[897] = ~((layer2_outputs[7183]) ^ (layer2_outputs[9897]));
    assign outputs[898] = layer2_outputs[7790];
    assign outputs[899] = (layer2_outputs[6029]) ^ (layer2_outputs[4930]);
    assign outputs[900] = (layer2_outputs[4822]) ^ (layer2_outputs[1553]);
    assign outputs[901] = ~((layer2_outputs[10347]) | (layer2_outputs[10846]));
    assign outputs[902] = ~(layer2_outputs[1134]);
    assign outputs[903] = (layer2_outputs[976]) ^ (layer2_outputs[10098]);
    assign outputs[904] = layer2_outputs[6525];
    assign outputs[905] = (layer2_outputs[11171]) ^ (layer2_outputs[12123]);
    assign outputs[906] = layer2_outputs[137];
    assign outputs[907] = ~(layer2_outputs[291]) | (layer2_outputs[12274]);
    assign outputs[908] = ~(layer2_outputs[11213]);
    assign outputs[909] = layer2_outputs[1926];
    assign outputs[910] = layer2_outputs[3709];
    assign outputs[911] = (layer2_outputs[550]) & (layer2_outputs[8515]);
    assign outputs[912] = ~(layer2_outputs[7713]);
    assign outputs[913] = layer2_outputs[5140];
    assign outputs[914] = (layer2_outputs[6085]) & (layer2_outputs[12489]);
    assign outputs[915] = ~(layer2_outputs[5688]);
    assign outputs[916] = ~((layer2_outputs[8497]) ^ (layer2_outputs[7702]));
    assign outputs[917] = (layer2_outputs[945]) ^ (layer2_outputs[3579]);
    assign outputs[918] = layer2_outputs[8043];
    assign outputs[919] = (layer2_outputs[12408]) & ~(layer2_outputs[7914]);
    assign outputs[920] = ~((layer2_outputs[10289]) & (layer2_outputs[1047]));
    assign outputs[921] = ~((layer2_outputs[7935]) ^ (layer2_outputs[326]));
    assign outputs[922] = ~(layer2_outputs[8074]) | (layer2_outputs[10061]);
    assign outputs[923] = layer2_outputs[6710];
    assign outputs[924] = ~(layer2_outputs[9779]);
    assign outputs[925] = (layer2_outputs[3179]) & (layer2_outputs[9266]);
    assign outputs[926] = (layer2_outputs[8357]) & ~(layer2_outputs[186]);
    assign outputs[927] = ~(layer2_outputs[2049]);
    assign outputs[928] = (layer2_outputs[6139]) ^ (layer2_outputs[8526]);
    assign outputs[929] = ~(layer2_outputs[5647]);
    assign outputs[930] = layer2_outputs[4438];
    assign outputs[931] = ~(layer2_outputs[5539]);
    assign outputs[932] = ~(layer2_outputs[7451]) | (layer2_outputs[890]);
    assign outputs[933] = layer2_outputs[8347];
    assign outputs[934] = ~(layer2_outputs[2297]);
    assign outputs[935] = (layer2_outputs[2221]) & ~(layer2_outputs[3421]);
    assign outputs[936] = ~((layer2_outputs[3987]) ^ (layer2_outputs[9564]));
    assign outputs[937] = (layer2_outputs[4823]) ^ (layer2_outputs[5164]);
    assign outputs[938] = (layer2_outputs[1574]) ^ (layer2_outputs[5420]);
    assign outputs[939] = (layer2_outputs[7046]) & ~(layer2_outputs[10885]);
    assign outputs[940] = layer2_outputs[7217];
    assign outputs[941] = layer2_outputs[12600];
    assign outputs[942] = layer2_outputs[10670];
    assign outputs[943] = (layer2_outputs[7303]) & (layer2_outputs[5480]);
    assign outputs[944] = ~(layer2_outputs[1798]);
    assign outputs[945] = ~((layer2_outputs[12494]) ^ (layer2_outputs[11974]));
    assign outputs[946] = layer2_outputs[10739];
    assign outputs[947] = layer2_outputs[11637];
    assign outputs[948] = layer2_outputs[11892];
    assign outputs[949] = ~((layer2_outputs[5759]) ^ (layer2_outputs[11620]));
    assign outputs[950] = layer2_outputs[4682];
    assign outputs[951] = layer2_outputs[12056];
    assign outputs[952] = ~(layer2_outputs[3243]) | (layer2_outputs[1086]);
    assign outputs[953] = ~(layer2_outputs[1918]);
    assign outputs[954] = (layer2_outputs[2870]) | (layer2_outputs[683]);
    assign outputs[955] = layer2_outputs[8295];
    assign outputs[956] = (layer2_outputs[1584]) ^ (layer2_outputs[3287]);
    assign outputs[957] = ~(layer2_outputs[11102]);
    assign outputs[958] = ~((layer2_outputs[8191]) & (layer2_outputs[5191]));
    assign outputs[959] = ~(layer2_outputs[35]);
    assign outputs[960] = ~(layer2_outputs[7157]) | (layer2_outputs[7989]);
    assign outputs[961] = ~(layer2_outputs[11079]);
    assign outputs[962] = layer2_outputs[1486];
    assign outputs[963] = ~((layer2_outputs[3603]) & (layer2_outputs[7836]));
    assign outputs[964] = ~(layer2_outputs[11617]) | (layer2_outputs[6466]);
    assign outputs[965] = ~(layer2_outputs[1962]);
    assign outputs[966] = ~(layer2_outputs[6060]);
    assign outputs[967] = ~(layer2_outputs[11003]);
    assign outputs[968] = ~((layer2_outputs[11160]) & (layer2_outputs[11677]));
    assign outputs[969] = layer2_outputs[1637];
    assign outputs[970] = ~(layer2_outputs[8741]);
    assign outputs[971] = ~(layer2_outputs[11102]);
    assign outputs[972] = layer2_outputs[9260];
    assign outputs[973] = ~(layer2_outputs[6484]) | (layer2_outputs[5231]);
    assign outputs[974] = layer2_outputs[3843];
    assign outputs[975] = (layer2_outputs[7432]) ^ (layer2_outputs[1251]);
    assign outputs[976] = ~((layer2_outputs[5368]) ^ (layer2_outputs[6841]));
    assign outputs[977] = layer2_outputs[4209];
    assign outputs[978] = (layer2_outputs[9197]) | (layer2_outputs[1344]);
    assign outputs[979] = layer2_outputs[7038];
    assign outputs[980] = layer2_outputs[6380];
    assign outputs[981] = ~(layer2_outputs[7823]);
    assign outputs[982] = ~(layer2_outputs[3958]);
    assign outputs[983] = layer2_outputs[4595];
    assign outputs[984] = ~(layer2_outputs[6754]);
    assign outputs[985] = ~(layer2_outputs[6580]);
    assign outputs[986] = ~(layer2_outputs[12565]);
    assign outputs[987] = (layer2_outputs[9698]) & (layer2_outputs[6364]);
    assign outputs[988] = ~(layer2_outputs[1264]);
    assign outputs[989] = ~(layer2_outputs[7112]) | (layer2_outputs[2894]);
    assign outputs[990] = layer2_outputs[11870];
    assign outputs[991] = ~(layer2_outputs[7092]) | (layer2_outputs[530]);
    assign outputs[992] = layer2_outputs[3984];
    assign outputs[993] = (layer2_outputs[12021]) ^ (layer2_outputs[8388]);
    assign outputs[994] = layer2_outputs[9785];
    assign outputs[995] = layer2_outputs[9397];
    assign outputs[996] = ~((layer2_outputs[3555]) | (layer2_outputs[8045]));
    assign outputs[997] = (layer2_outputs[2337]) ^ (layer2_outputs[3968]);
    assign outputs[998] = (layer2_outputs[2010]) & (layer2_outputs[7122]);
    assign outputs[999] = layer2_outputs[11569];
    assign outputs[1000] = (layer2_outputs[3666]) & ~(layer2_outputs[3398]);
    assign outputs[1001] = layer2_outputs[4543];
    assign outputs[1002] = ~(layer2_outputs[352]);
    assign outputs[1003] = ~(layer2_outputs[7840]);
    assign outputs[1004] = ~(layer2_outputs[2350]);
    assign outputs[1005] = layer2_outputs[11154];
    assign outputs[1006] = ~(layer2_outputs[7562]);
    assign outputs[1007] = layer2_outputs[3569];
    assign outputs[1008] = ~(layer2_outputs[9876]);
    assign outputs[1009] = ~(layer2_outputs[10975]);
    assign outputs[1010] = ~((layer2_outputs[3370]) ^ (layer2_outputs[12248]));
    assign outputs[1011] = ~(layer2_outputs[10745]);
    assign outputs[1012] = (layer2_outputs[11219]) | (layer2_outputs[11843]);
    assign outputs[1013] = layer2_outputs[4067];
    assign outputs[1014] = layer2_outputs[1447];
    assign outputs[1015] = layer2_outputs[213];
    assign outputs[1016] = (layer2_outputs[7899]) & (layer2_outputs[10331]);
    assign outputs[1017] = ~(layer2_outputs[8901]);
    assign outputs[1018] = ~(layer2_outputs[5504]);
    assign outputs[1019] = ~(layer2_outputs[416]);
    assign outputs[1020] = ~(layer2_outputs[7740]);
    assign outputs[1021] = ~(layer2_outputs[3627]);
    assign outputs[1022] = (layer2_outputs[7670]) ^ (layer2_outputs[5090]);
    assign outputs[1023] = (layer2_outputs[3451]) | (layer2_outputs[9230]);
    assign outputs[1024] = ~(layer2_outputs[11158]);
    assign outputs[1025] = layer2_outputs[6898];
    assign outputs[1026] = ~(layer2_outputs[12678]);
    assign outputs[1027] = layer2_outputs[7373];
    assign outputs[1028] = ~(layer2_outputs[11094]);
    assign outputs[1029] = layer2_outputs[12127];
    assign outputs[1030] = (layer2_outputs[1333]) ^ (layer2_outputs[1858]);
    assign outputs[1031] = (layer2_outputs[9410]) & ~(layer2_outputs[7520]);
    assign outputs[1032] = ~((layer2_outputs[7400]) ^ (layer2_outputs[8245]));
    assign outputs[1033] = layer2_outputs[12624];
    assign outputs[1034] = ~(layer2_outputs[4620]);
    assign outputs[1035] = layer2_outputs[1250];
    assign outputs[1036] = layer2_outputs[1275];
    assign outputs[1037] = ~(layer2_outputs[12254]);
    assign outputs[1038] = ~((layer2_outputs[316]) | (layer2_outputs[7820]));
    assign outputs[1039] = (layer2_outputs[8972]) ^ (layer2_outputs[11951]);
    assign outputs[1040] = ~((layer2_outputs[5170]) | (layer2_outputs[3238]));
    assign outputs[1041] = (layer2_outputs[5721]) | (layer2_outputs[7644]);
    assign outputs[1042] = layer2_outputs[9532];
    assign outputs[1043] = (layer2_outputs[7291]) ^ (layer2_outputs[11518]);
    assign outputs[1044] = ~(layer2_outputs[11029]) | (layer2_outputs[10720]);
    assign outputs[1045] = ~(layer2_outputs[9960]);
    assign outputs[1046] = ~((layer2_outputs[4927]) ^ (layer2_outputs[7282]));
    assign outputs[1047] = ~((layer2_outputs[2320]) ^ (layer2_outputs[1975]));
    assign outputs[1048] = ~((layer2_outputs[3881]) ^ (layer2_outputs[8380]));
    assign outputs[1049] = layer2_outputs[8472];
    assign outputs[1050] = ~(layer2_outputs[124]);
    assign outputs[1051] = ~(layer2_outputs[4369]);
    assign outputs[1052] = ~(layer2_outputs[3121]);
    assign outputs[1053] = ~(layer2_outputs[5245]);
    assign outputs[1054] = (layer2_outputs[769]) & ~(layer2_outputs[12555]);
    assign outputs[1055] = ~(layer2_outputs[6624]);
    assign outputs[1056] = ~(layer2_outputs[9466]);
    assign outputs[1057] = (layer2_outputs[11882]) & ~(layer2_outputs[5674]);
    assign outputs[1058] = ~(layer2_outputs[7536]);
    assign outputs[1059] = ~(layer2_outputs[7165]);
    assign outputs[1060] = ~(layer2_outputs[10193]);
    assign outputs[1061] = ~(layer2_outputs[3267]);
    assign outputs[1062] = layer2_outputs[10662];
    assign outputs[1063] = (layer2_outputs[9136]) & ~(layer2_outputs[777]);
    assign outputs[1064] = ~(layer2_outputs[12719]);
    assign outputs[1065] = layer2_outputs[7527];
    assign outputs[1066] = layer2_outputs[5763];
    assign outputs[1067] = ~((layer2_outputs[3873]) ^ (layer2_outputs[12495]));
    assign outputs[1068] = ~((layer2_outputs[1524]) ^ (layer2_outputs[6491]));
    assign outputs[1069] = (layer2_outputs[9885]) ^ (layer2_outputs[9846]);
    assign outputs[1070] = ~(layer2_outputs[11403]);
    assign outputs[1071] = layer2_outputs[10336];
    assign outputs[1072] = (layer2_outputs[9901]) & (layer2_outputs[5725]);
    assign outputs[1073] = layer2_outputs[6185];
    assign outputs[1074] = ~(layer2_outputs[12671]);
    assign outputs[1075] = ~((layer2_outputs[11830]) ^ (layer2_outputs[6735]));
    assign outputs[1076] = ~(layer2_outputs[2493]);
    assign outputs[1077] = (layer2_outputs[8572]) & (layer2_outputs[7236]);
    assign outputs[1078] = ~((layer2_outputs[4415]) ^ (layer2_outputs[7898]));
    assign outputs[1079] = layer2_outputs[9762];
    assign outputs[1080] = ~((layer2_outputs[2762]) & (layer2_outputs[1304]));
    assign outputs[1081] = ~(layer2_outputs[7269]) | (layer2_outputs[11886]);
    assign outputs[1082] = layer2_outputs[12472];
    assign outputs[1083] = layer2_outputs[3790];
    assign outputs[1084] = layer2_outputs[5379];
    assign outputs[1085] = ~(layer2_outputs[1955]);
    assign outputs[1086] = ~(layer2_outputs[8324]) | (layer2_outputs[1030]);
    assign outputs[1087] = (layer2_outputs[7073]) & (layer2_outputs[9824]);
    assign outputs[1088] = layer2_outputs[2201];
    assign outputs[1089] = ~((layer2_outputs[4132]) | (layer2_outputs[3425]));
    assign outputs[1090] = layer2_outputs[12585];
    assign outputs[1091] = layer2_outputs[5333];
    assign outputs[1092] = (layer2_outputs[8922]) & ~(layer2_outputs[7588]);
    assign outputs[1093] = (layer2_outputs[1593]) & (layer2_outputs[8477]);
    assign outputs[1094] = layer2_outputs[9862];
    assign outputs[1095] = layer2_outputs[12301];
    assign outputs[1096] = layer2_outputs[10002];
    assign outputs[1097] = (layer2_outputs[5067]) & ~(layer2_outputs[2715]);
    assign outputs[1098] = (layer2_outputs[2800]) ^ (layer2_outputs[8391]);
    assign outputs[1099] = layer2_outputs[11829];
    assign outputs[1100] = layer2_outputs[11880];
    assign outputs[1101] = ~((layer2_outputs[269]) | (layer2_outputs[4103]));
    assign outputs[1102] = layer2_outputs[5251];
    assign outputs[1103] = (layer2_outputs[5389]) ^ (layer2_outputs[12052]);
    assign outputs[1104] = ~(layer2_outputs[10748]);
    assign outputs[1105] = (layer2_outputs[3943]) & ~(layer2_outputs[3089]);
    assign outputs[1106] = layer2_outputs[4251];
    assign outputs[1107] = ~(layer2_outputs[1857]) | (layer2_outputs[11411]);
    assign outputs[1108] = (layer2_outputs[6483]) & ~(layer2_outputs[9143]);
    assign outputs[1109] = layer2_outputs[1025];
    assign outputs[1110] = ~((layer2_outputs[3753]) & (layer2_outputs[6455]));
    assign outputs[1111] = (layer2_outputs[8185]) & ~(layer2_outputs[3591]);
    assign outputs[1112] = (layer2_outputs[10872]) | (layer2_outputs[5744]);
    assign outputs[1113] = layer2_outputs[2420];
    assign outputs[1114] = ~((layer2_outputs[7951]) | (layer2_outputs[5208]));
    assign outputs[1115] = layer2_outputs[4006];
    assign outputs[1116] = layer2_outputs[828];
    assign outputs[1117] = (layer2_outputs[5455]) & ~(layer2_outputs[10457]);
    assign outputs[1118] = layer2_outputs[10134];
    assign outputs[1119] = ~(layer2_outputs[1270]);
    assign outputs[1120] = ~((layer2_outputs[10904]) ^ (layer2_outputs[10521]));
    assign outputs[1121] = (layer2_outputs[2990]) ^ (layer2_outputs[12399]);
    assign outputs[1122] = ~((layer2_outputs[326]) ^ (layer2_outputs[7123]));
    assign outputs[1123] = ~(layer2_outputs[4700]);
    assign outputs[1124] = ~(layer2_outputs[10971]);
    assign outputs[1125] = ~((layer2_outputs[2891]) ^ (layer2_outputs[2687]));
    assign outputs[1126] = ~(layer2_outputs[12264]);
    assign outputs[1127] = ~(layer2_outputs[5984]);
    assign outputs[1128] = layer2_outputs[225];
    assign outputs[1129] = (layer2_outputs[4767]) & ~(layer2_outputs[12548]);
    assign outputs[1130] = layer2_outputs[3146];
    assign outputs[1131] = (layer2_outputs[3568]) & ~(layer2_outputs[1882]);
    assign outputs[1132] = ~(layer2_outputs[10924]) | (layer2_outputs[11228]);
    assign outputs[1133] = ~(layer2_outputs[5159]);
    assign outputs[1134] = layer2_outputs[9385];
    assign outputs[1135] = (layer2_outputs[6162]) & (layer2_outputs[5666]);
    assign outputs[1136] = layer2_outputs[12405];
    assign outputs[1137] = layer2_outputs[5869];
    assign outputs[1138] = layer2_outputs[8013];
    assign outputs[1139] = (layer2_outputs[87]) & (layer2_outputs[7466]);
    assign outputs[1140] = ~(layer2_outputs[4013]);
    assign outputs[1141] = (layer2_outputs[4120]) & ~(layer2_outputs[10865]);
    assign outputs[1142] = ~(layer2_outputs[1307]);
    assign outputs[1143] = ~((layer2_outputs[10895]) ^ (layer2_outputs[7949]));
    assign outputs[1144] = layer2_outputs[10503];
    assign outputs[1145] = ~(layer2_outputs[4678]) | (layer2_outputs[5599]);
    assign outputs[1146] = (layer2_outputs[12317]) & ~(layer2_outputs[951]);
    assign outputs[1147] = ~(layer2_outputs[3842]);
    assign outputs[1148] = ~((layer2_outputs[9738]) ^ (layer2_outputs[6748]));
    assign outputs[1149] = ~(layer2_outputs[10441]);
    assign outputs[1150] = ~(layer2_outputs[8182]);
    assign outputs[1151] = layer2_outputs[10278];
    assign outputs[1152] = ~(layer2_outputs[8423]);
    assign outputs[1153] = (layer2_outputs[5929]) & (layer2_outputs[11502]);
    assign outputs[1154] = layer2_outputs[9064];
    assign outputs[1155] = layer2_outputs[9127];
    assign outputs[1156] = ~((layer2_outputs[6310]) ^ (layer2_outputs[892]));
    assign outputs[1157] = layer2_outputs[2427];
    assign outputs[1158] = ~(layer2_outputs[3712]);
    assign outputs[1159] = ~(layer2_outputs[5182]);
    assign outputs[1160] = ~((layer2_outputs[4347]) ^ (layer2_outputs[11635]));
    assign outputs[1161] = layer2_outputs[7503];
    assign outputs[1162] = ~((layer2_outputs[11121]) ^ (layer2_outputs[915]));
    assign outputs[1163] = (layer2_outputs[8991]) & ~(layer2_outputs[10461]);
    assign outputs[1164] = ~(layer2_outputs[5531]) | (layer2_outputs[9570]);
    assign outputs[1165] = ~((layer2_outputs[11505]) ^ (layer2_outputs[4653]));
    assign outputs[1166] = layer2_outputs[4912];
    assign outputs[1167] = ~((layer2_outputs[6161]) ^ (layer2_outputs[4245]));
    assign outputs[1168] = layer2_outputs[9012];
    assign outputs[1169] = ~(layer2_outputs[4692]);
    assign outputs[1170] = ~((layer2_outputs[2236]) & (layer2_outputs[7325]));
    assign outputs[1171] = ~((layer2_outputs[5621]) ^ (layer2_outputs[9963]));
    assign outputs[1172] = layer2_outputs[10217];
    assign outputs[1173] = ~(layer2_outputs[4546]);
    assign outputs[1174] = ~((layer2_outputs[2567]) & (layer2_outputs[11944]));
    assign outputs[1175] = ~((layer2_outputs[5934]) ^ (layer2_outputs[6328]));
    assign outputs[1176] = ~(layer2_outputs[7682]) | (layer2_outputs[1098]);
    assign outputs[1177] = (layer2_outputs[6314]) ^ (layer2_outputs[374]);
    assign outputs[1178] = ~(layer2_outputs[11321]);
    assign outputs[1179] = layer2_outputs[4107];
    assign outputs[1180] = layer2_outputs[10102];
    assign outputs[1181] = layer2_outputs[1903];
    assign outputs[1182] = layer2_outputs[4138];
    assign outputs[1183] = ~(layer2_outputs[5580]);
    assign outputs[1184] = ~(layer2_outputs[3654]);
    assign outputs[1185] = (layer2_outputs[289]) | (layer2_outputs[12015]);
    assign outputs[1186] = ~(layer2_outputs[9210]);
    assign outputs[1187] = layer2_outputs[8687];
    assign outputs[1188] = ~(layer2_outputs[8412]) | (layer2_outputs[11876]);
    assign outputs[1189] = (layer2_outputs[611]) ^ (layer2_outputs[1722]);
    assign outputs[1190] = (layer2_outputs[6845]) ^ (layer2_outputs[3496]);
    assign outputs[1191] = ~(layer2_outputs[5876]);
    assign outputs[1192] = (layer2_outputs[1314]) ^ (layer2_outputs[3832]);
    assign outputs[1193] = layer2_outputs[8401];
    assign outputs[1194] = ~(layer2_outputs[6697]);
    assign outputs[1195] = layer2_outputs[9287];
    assign outputs[1196] = layer2_outputs[4756];
    assign outputs[1197] = ~(layer2_outputs[8878]);
    assign outputs[1198] = ~(layer2_outputs[7755]);
    assign outputs[1199] = (layer2_outputs[4329]) ^ (layer2_outputs[11438]);
    assign outputs[1200] = ~(layer2_outputs[12564]);
    assign outputs[1201] = ~((layer2_outputs[7496]) ^ (layer2_outputs[3848]));
    assign outputs[1202] = ~(layer2_outputs[7991]);
    assign outputs[1203] = ~((layer2_outputs[9757]) ^ (layer2_outputs[9829]));
    assign outputs[1204] = ~((layer2_outputs[1987]) & (layer2_outputs[8367]));
    assign outputs[1205] = (layer2_outputs[9097]) ^ (layer2_outputs[10202]);
    assign outputs[1206] = ~(layer2_outputs[10984]);
    assign outputs[1207] = (layer2_outputs[5787]) & ~(layer2_outputs[1696]);
    assign outputs[1208] = ~(layer2_outputs[731]);
    assign outputs[1209] = ~((layer2_outputs[8578]) ^ (layer2_outputs[8864]));
    assign outputs[1210] = layer2_outputs[12535];
    assign outputs[1211] = layer2_outputs[6262];
    assign outputs[1212] = layer2_outputs[4100];
    assign outputs[1213] = ~((layer2_outputs[2995]) ^ (layer2_outputs[7931]));
    assign outputs[1214] = ~(layer2_outputs[4635]);
    assign outputs[1215] = ~((layer2_outputs[7672]) | (layer2_outputs[1567]));
    assign outputs[1216] = (layer2_outputs[4753]) & (layer2_outputs[3099]);
    assign outputs[1217] = layer2_outputs[2482];
    assign outputs[1218] = layer2_outputs[1644];
    assign outputs[1219] = ~((layer2_outputs[3676]) ^ (layer2_outputs[3503]));
    assign outputs[1220] = (layer2_outputs[1839]) & (layer2_outputs[5475]);
    assign outputs[1221] = layer2_outputs[581];
    assign outputs[1222] = (layer2_outputs[6277]) ^ (layer2_outputs[9696]);
    assign outputs[1223] = layer2_outputs[6158];
    assign outputs[1224] = ~((layer2_outputs[2661]) ^ (layer2_outputs[5334]));
    assign outputs[1225] = ~(layer2_outputs[2782]);
    assign outputs[1226] = ~(layer2_outputs[5747]) | (layer2_outputs[4643]);
    assign outputs[1227] = layer2_outputs[3870];
    assign outputs[1228] = layer2_outputs[11088];
    assign outputs[1229] = ~((layer2_outputs[1930]) & (layer2_outputs[3444]));
    assign outputs[1230] = ~((layer2_outputs[10363]) & (layer2_outputs[1924]));
    assign outputs[1231] = ~(layer2_outputs[3176]) | (layer2_outputs[9778]);
    assign outputs[1232] = layer2_outputs[2363];
    assign outputs[1233] = ~(layer2_outputs[8389]) | (layer2_outputs[11148]);
    assign outputs[1234] = ~(layer2_outputs[6984]);
    assign outputs[1235] = ~(layer2_outputs[3390]);
    assign outputs[1236] = ~(layer2_outputs[8095]) | (layer2_outputs[3058]);
    assign outputs[1237] = (layer2_outputs[2839]) & ~(layer2_outputs[6982]);
    assign outputs[1238] = (layer2_outputs[28]) ^ (layer2_outputs[7689]);
    assign outputs[1239] = (layer2_outputs[8004]) ^ (layer2_outputs[7559]);
    assign outputs[1240] = ~(layer2_outputs[9619]);
    assign outputs[1241] = (layer2_outputs[2787]) & (layer2_outputs[7721]);
    assign outputs[1242] = ~(layer2_outputs[3196]);
    assign outputs[1243] = ~(layer2_outputs[3301]);
    assign outputs[1244] = (layer2_outputs[11596]) ^ (layer2_outputs[4757]);
    assign outputs[1245] = ~(layer2_outputs[12155]);
    assign outputs[1246] = ~((layer2_outputs[9921]) ^ (layer2_outputs[84]));
    assign outputs[1247] = (layer2_outputs[11531]) & (layer2_outputs[10452]);
    assign outputs[1248] = layer2_outputs[2742];
    assign outputs[1249] = ~(layer2_outputs[4388]) | (layer2_outputs[6798]);
    assign outputs[1250] = ~(layer2_outputs[10342]) | (layer2_outputs[2090]);
    assign outputs[1251] = ~((layer2_outputs[6630]) ^ (layer2_outputs[11429]));
    assign outputs[1252] = ~(layer2_outputs[8282]);
    assign outputs[1253] = (layer2_outputs[10900]) ^ (layer2_outputs[3353]);
    assign outputs[1254] = ~(layer2_outputs[8234]);
    assign outputs[1255] = ~(layer2_outputs[3822]) | (layer2_outputs[3384]);
    assign outputs[1256] = ~((layer2_outputs[9503]) | (layer2_outputs[5944]));
    assign outputs[1257] = ~(layer2_outputs[1786]);
    assign outputs[1258] = (layer2_outputs[7831]) | (layer2_outputs[696]);
    assign outputs[1259] = layer2_outputs[7735];
    assign outputs[1260] = ~(layer2_outputs[9406]);
    assign outputs[1261] = (layer2_outputs[5853]) ^ (layer2_outputs[8442]);
    assign outputs[1262] = (layer2_outputs[11067]) | (layer2_outputs[8498]);
    assign outputs[1263] = ~(layer2_outputs[1255]);
    assign outputs[1264] = ~((layer2_outputs[8817]) ^ (layer2_outputs[357]));
    assign outputs[1265] = ~(layer2_outputs[1883]);
    assign outputs[1266] = ~((layer2_outputs[10728]) ^ (layer2_outputs[11787]));
    assign outputs[1267] = (layer2_outputs[3566]) | (layer2_outputs[2074]);
    assign outputs[1268] = ~(layer2_outputs[10514]);
    assign outputs[1269] = ~(layer2_outputs[4088]);
    assign outputs[1270] = (layer2_outputs[4501]) & ~(layer2_outputs[12729]);
    assign outputs[1271] = (layer2_outputs[11957]) & ~(layer2_outputs[11216]);
    assign outputs[1272] = ~(layer2_outputs[9481]) | (layer2_outputs[8164]);
    assign outputs[1273] = ~((layer2_outputs[2829]) ^ (layer2_outputs[3634]));
    assign outputs[1274] = ~(layer2_outputs[5423]);
    assign outputs[1275] = (layer2_outputs[9823]) & (layer2_outputs[1709]);
    assign outputs[1276] = ~(layer2_outputs[1986]);
    assign outputs[1277] = ~(layer2_outputs[2903]);
    assign outputs[1278] = layer2_outputs[10630];
    assign outputs[1279] = (layer2_outputs[7641]) ^ (layer2_outputs[701]);
    assign outputs[1280] = (layer2_outputs[1851]) ^ (layer2_outputs[4266]);
    assign outputs[1281] = ~((layer2_outputs[7225]) | (layer2_outputs[8351]));
    assign outputs[1282] = (layer2_outputs[11478]) & ~(layer2_outputs[10389]);
    assign outputs[1283] = ~(layer2_outputs[178]);
    assign outputs[1284] = (layer2_outputs[3265]) & ~(layer2_outputs[2368]);
    assign outputs[1285] = ~((layer2_outputs[2323]) ^ (layer2_outputs[10024]));
    assign outputs[1286] = layer2_outputs[147];
    assign outputs[1287] = layer2_outputs[11618];
    assign outputs[1288] = (layer2_outputs[5616]) & (layer2_outputs[11786]);
    assign outputs[1289] = layer2_outputs[7609];
    assign outputs[1290] = (layer2_outputs[5733]) & ~(layer2_outputs[9521]);
    assign outputs[1291] = ~(layer2_outputs[10707]);
    assign outputs[1292] = ~(layer2_outputs[6407]);
    assign outputs[1293] = ~((layer2_outputs[2784]) ^ (layer2_outputs[7913]));
    assign outputs[1294] = (layer2_outputs[7777]) ^ (layer2_outputs[8181]);
    assign outputs[1295] = layer2_outputs[2953];
    assign outputs[1296] = layer2_outputs[10489];
    assign outputs[1297] = ~((layer2_outputs[7930]) ^ (layer2_outputs[541]));
    assign outputs[1298] = (layer2_outputs[4372]) & (layer2_outputs[11422]);
    assign outputs[1299] = (layer2_outputs[12659]) & ~(layer2_outputs[234]);
    assign outputs[1300] = (layer2_outputs[1478]) ^ (layer2_outputs[107]);
    assign outputs[1301] = ~((layer2_outputs[5447]) ^ (layer2_outputs[4778]));
    assign outputs[1302] = ~((layer2_outputs[11396]) ^ (layer2_outputs[7950]));
    assign outputs[1303] = ~((layer2_outputs[7126]) ^ (layer2_outputs[12217]));
    assign outputs[1304] = ~((layer2_outputs[8065]) | (layer2_outputs[5805]));
    assign outputs[1305] = ~((layer2_outputs[3053]) | (layer2_outputs[2720]));
    assign outputs[1306] = ~((layer2_outputs[8671]) ^ (layer2_outputs[10251]));
    assign outputs[1307] = ~((layer2_outputs[8123]) | (layer2_outputs[5312]));
    assign outputs[1308] = ~(layer2_outputs[9965]);
    assign outputs[1309] = layer2_outputs[1810];
    assign outputs[1310] = layer2_outputs[12781];
    assign outputs[1311] = (layer2_outputs[8192]) & ~(layer2_outputs[8048]);
    assign outputs[1312] = ~(layer2_outputs[910]);
    assign outputs[1313] = (layer2_outputs[6842]) ^ (layer2_outputs[5629]);
    assign outputs[1314] = ~((layer2_outputs[11238]) ^ (layer2_outputs[12138]));
    assign outputs[1315] = ~((layer2_outputs[5677]) ^ (layer2_outputs[6067]));
    assign outputs[1316] = ~((layer2_outputs[417]) ^ (layer2_outputs[11866]));
    assign outputs[1317] = (layer2_outputs[9008]) ^ (layer2_outputs[7458]);
    assign outputs[1318] = layer2_outputs[5862];
    assign outputs[1319] = ~((layer2_outputs[12642]) & (layer2_outputs[3503]));
    assign outputs[1320] = ~(layer2_outputs[1462]) | (layer2_outputs[5632]);
    assign outputs[1321] = (layer2_outputs[10450]) & (layer2_outputs[6445]);
    assign outputs[1322] = layer2_outputs[9362];
    assign outputs[1323] = ~((layer2_outputs[2236]) ^ (layer2_outputs[4295]));
    assign outputs[1324] = (layer2_outputs[7539]) & (layer2_outputs[7610]);
    assign outputs[1325] = (layer2_outputs[686]) ^ (layer2_outputs[12701]);
    assign outputs[1326] = ~((layer2_outputs[4566]) & (layer2_outputs[969]));
    assign outputs[1327] = (layer2_outputs[5175]) & ~(layer2_outputs[10750]);
    assign outputs[1328] = ~(layer2_outputs[8990]);
    assign outputs[1329] = layer2_outputs[12505];
    assign outputs[1330] = (layer2_outputs[9212]) ^ (layer2_outputs[12497]);
    assign outputs[1331] = ~((layer2_outputs[5109]) & (layer2_outputs[9371]));
    assign outputs[1332] = ~(layer2_outputs[8870]);
    assign outputs[1333] = ~((layer2_outputs[7606]) ^ (layer2_outputs[10649]));
    assign outputs[1334] = ~(layer2_outputs[3275]);
    assign outputs[1335] = (layer2_outputs[1232]) & ~(layer2_outputs[2434]);
    assign outputs[1336] = ~(layer2_outputs[2735]);
    assign outputs[1337] = ~(layer2_outputs[734]);
    assign outputs[1338] = ~(layer2_outputs[9622]);
    assign outputs[1339] = ~((layer2_outputs[10624]) ^ (layer2_outputs[12711]));
    assign outputs[1340] = ~(layer2_outputs[6347]);
    assign outputs[1341] = (layer2_outputs[8242]) & ~(layer2_outputs[3593]);
    assign outputs[1342] = ~((layer2_outputs[9024]) | (layer2_outputs[1183]));
    assign outputs[1343] = ~((layer2_outputs[7431]) ^ (layer2_outputs[4913]));
    assign outputs[1344] = ~(layer2_outputs[7044]);
    assign outputs[1345] = ~((layer2_outputs[3633]) ^ (layer2_outputs[9460]));
    assign outputs[1346] = layer2_outputs[5421];
    assign outputs[1347] = layer2_outputs[5365];
    assign outputs[1348] = layer2_outputs[2627];
    assign outputs[1349] = layer2_outputs[12734];
    assign outputs[1350] = layer2_outputs[10862];
    assign outputs[1351] = (layer2_outputs[12188]) ^ (layer2_outputs[12582]);
    assign outputs[1352] = layer2_outputs[6773];
    assign outputs[1353] = (layer2_outputs[3517]) ^ (layer2_outputs[2501]);
    assign outputs[1354] = ~(layer2_outputs[3181]);
    assign outputs[1355] = (layer2_outputs[11476]) ^ (layer2_outputs[4779]);
    assign outputs[1356] = layer2_outputs[4180];
    assign outputs[1357] = ~((layer2_outputs[5933]) | (layer2_outputs[8603]));
    assign outputs[1358] = ~(layer2_outputs[7290]) | (layer2_outputs[8774]);
    assign outputs[1359] = ~(layer2_outputs[10750]);
    assign outputs[1360] = (layer2_outputs[6774]) & (layer2_outputs[1814]);
    assign outputs[1361] = (layer2_outputs[1758]) ^ (layer2_outputs[4856]);
    assign outputs[1362] = ~(layer2_outputs[8563]) | (layer2_outputs[1030]);
    assign outputs[1363] = ~((layer2_outputs[451]) | (layer2_outputs[8054]));
    assign outputs[1364] = ~(layer2_outputs[2451]);
    assign outputs[1365] = ~((layer2_outputs[5411]) | (layer2_outputs[5755]));
    assign outputs[1366] = (layer2_outputs[9361]) & ~(layer2_outputs[5681]);
    assign outputs[1367] = layer2_outputs[4013];
    assign outputs[1368] = ~((layer2_outputs[6389]) | (layer2_outputs[4532]));
    assign outputs[1369] = (layer2_outputs[7147]) & ~(layer2_outputs[11569]);
    assign outputs[1370] = (layer2_outputs[6411]) & ~(layer2_outputs[5503]);
    assign outputs[1371] = layer2_outputs[11113];
    assign outputs[1372] = ~((layer2_outputs[10839]) ^ (layer2_outputs[6088]));
    assign outputs[1373] = layer2_outputs[3078];
    assign outputs[1374] = ~((layer2_outputs[7615]) ^ (layer2_outputs[5082]));
    assign outputs[1375] = (layer2_outputs[5695]) & ~(layer2_outputs[7557]);
    assign outputs[1376] = ~((layer2_outputs[9446]) ^ (layer2_outputs[6544]));
    assign outputs[1377] = (layer2_outputs[8736]) | (layer2_outputs[2208]);
    assign outputs[1378] = ~((layer2_outputs[4312]) ^ (layer2_outputs[1444]));
    assign outputs[1379] = ~((layer2_outputs[3523]) | (layer2_outputs[5103]));
    assign outputs[1380] = (layer2_outputs[6671]) & ~(layer2_outputs[1507]);
    assign outputs[1381] = layer2_outputs[159];
    assign outputs[1382] = (layer2_outputs[5601]) ^ (layer2_outputs[1361]);
    assign outputs[1383] = ~(layer2_outputs[11973]);
    assign outputs[1384] = (layer2_outputs[11295]) ^ (layer2_outputs[9103]);
    assign outputs[1385] = (layer2_outputs[137]) ^ (layer2_outputs[10185]);
    assign outputs[1386] = ~((layer2_outputs[7350]) ^ (layer2_outputs[10104]));
    assign outputs[1387] = ~(layer2_outputs[4424]);
    assign outputs[1388] = ~((layer2_outputs[1015]) ^ (layer2_outputs[9009]));
    assign outputs[1389] = ~(layer2_outputs[6649]);
    assign outputs[1390] = ~((layer2_outputs[1833]) & (layer2_outputs[6345]));
    assign outputs[1391] = ~((layer2_outputs[7103]) | (layer2_outputs[1261]));
    assign outputs[1392] = ~(layer2_outputs[5174]);
    assign outputs[1393] = (layer2_outputs[10874]) & (layer2_outputs[5985]);
    assign outputs[1394] = (layer2_outputs[7619]) ^ (layer2_outputs[5363]);
    assign outputs[1395] = ~((layer2_outputs[11589]) ^ (layer2_outputs[6663]));
    assign outputs[1396] = ~(layer2_outputs[11698]);
    assign outputs[1397] = (layer2_outputs[4904]) & ~(layer2_outputs[2420]);
    assign outputs[1398] = layer2_outputs[11179];
    assign outputs[1399] = ~((layer2_outputs[9834]) ^ (layer2_outputs[569]));
    assign outputs[1400] = (layer2_outputs[9651]) & (layer2_outputs[56]);
    assign outputs[1401] = layer2_outputs[5302];
    assign outputs[1402] = ~(layer2_outputs[10549]) | (layer2_outputs[10833]);
    assign outputs[1403] = ~(layer2_outputs[12542]);
    assign outputs[1404] = ~(layer2_outputs[6910]);
    assign outputs[1405] = (layer2_outputs[5911]) & ~(layer2_outputs[7086]);
    assign outputs[1406] = ~((layer2_outputs[10315]) ^ (layer2_outputs[10816]));
    assign outputs[1407] = layer2_outputs[2224];
    assign outputs[1408] = ~((layer2_outputs[10180]) ^ (layer2_outputs[2660]));
    assign outputs[1409] = (layer2_outputs[8695]) & ~(layer2_outputs[9348]);
    assign outputs[1410] = ~(layer2_outputs[8011]);
    assign outputs[1411] = layer2_outputs[6534];
    assign outputs[1412] = ~((layer2_outputs[1306]) ^ (layer2_outputs[5986]));
    assign outputs[1413] = ~(layer2_outputs[2059]);
    assign outputs[1414] = ~(layer2_outputs[8624]) | (layer2_outputs[2286]);
    assign outputs[1415] = ~(layer2_outputs[11198]);
    assign outputs[1416] = (layer2_outputs[7076]) & (layer2_outputs[11217]);
    assign outputs[1417] = ~((layer2_outputs[3158]) & (layer2_outputs[914]));
    assign outputs[1418] = layer2_outputs[11052];
    assign outputs[1419] = (layer2_outputs[5634]) & ~(layer2_outputs[748]);
    assign outputs[1420] = ~((layer2_outputs[7874]) & (layer2_outputs[10951]));
    assign outputs[1421] = ~((layer2_outputs[2840]) ^ (layer2_outputs[1790]));
    assign outputs[1422] = ~(layer2_outputs[2025]);
    assign outputs[1423] = (layer2_outputs[1273]) & ~(layer2_outputs[334]);
    assign outputs[1424] = (layer2_outputs[2184]) ^ (layer2_outputs[2231]);
    assign outputs[1425] = ~(layer2_outputs[4852]);
    assign outputs[1426] = (layer2_outputs[11879]) & ~(layer2_outputs[4014]);
    assign outputs[1427] = ~((layer2_outputs[11735]) | (layer2_outputs[8770]));
    assign outputs[1428] = ~((layer2_outputs[6059]) | (layer2_outputs[10419]));
    assign outputs[1429] = (layer2_outputs[7105]) ^ (layer2_outputs[4585]);
    assign outputs[1430] = ~(layer2_outputs[11160]);
    assign outputs[1431] = layer2_outputs[3667];
    assign outputs[1432] = ~((layer2_outputs[20]) ^ (layer2_outputs[1331]));
    assign outputs[1433] = ~(layer2_outputs[4042]) | (layer2_outputs[9842]);
    assign outputs[1434] = (layer2_outputs[10319]) ^ (layer2_outputs[5335]);
    assign outputs[1435] = layer2_outputs[4077];
    assign outputs[1436] = (layer2_outputs[12001]) & (layer2_outputs[3280]);
    assign outputs[1437] = layer2_outputs[6693];
    assign outputs[1438] = (layer2_outputs[10045]) & ~(layer2_outputs[3999]);
    assign outputs[1439] = (layer2_outputs[10966]) ^ (layer2_outputs[8748]);
    assign outputs[1440] = ~((layer2_outputs[9420]) | (layer2_outputs[3033]));
    assign outputs[1441] = (layer2_outputs[5119]) & ~(layer2_outputs[1564]);
    assign outputs[1442] = layer2_outputs[2876];
    assign outputs[1443] = layer2_outputs[3977];
    assign outputs[1444] = layer2_outputs[9656];
    assign outputs[1445] = layer2_outputs[5823];
    assign outputs[1446] = (layer2_outputs[10960]) & ~(layer2_outputs[11313]);
    assign outputs[1447] = (layer2_outputs[9558]) & ~(layer2_outputs[58]);
    assign outputs[1448] = layer2_outputs[5541];
    assign outputs[1449] = (layer2_outputs[8217]) ^ (layer2_outputs[11168]);
    assign outputs[1450] = (layer2_outputs[11922]) ^ (layer2_outputs[8885]);
    assign outputs[1451] = (layer2_outputs[12085]) & ~(layer2_outputs[4322]);
    assign outputs[1452] = ~(layer2_outputs[4886]);
    assign outputs[1453] = ~((layer2_outputs[5006]) ^ (layer2_outputs[12009]));
    assign outputs[1454] = (layer2_outputs[4071]) ^ (layer2_outputs[5265]);
    assign outputs[1455] = ~(layer2_outputs[1691]);
    assign outputs[1456] = (layer2_outputs[11733]) | (layer2_outputs[3263]);
    assign outputs[1457] = layer2_outputs[1560];
    assign outputs[1458] = (layer2_outputs[5372]) ^ (layer2_outputs[5740]);
    assign outputs[1459] = (layer2_outputs[3343]) ^ (layer2_outputs[9128]);
    assign outputs[1460] = (layer2_outputs[10147]) ^ (layer2_outputs[12067]);
    assign outputs[1461] = (layer2_outputs[2614]) & ~(layer2_outputs[3599]);
    assign outputs[1462] = (layer2_outputs[9681]) & (layer2_outputs[8608]);
    assign outputs[1463] = (layer2_outputs[8671]) & (layer2_outputs[5428]);
    assign outputs[1464] = ~((layer2_outputs[6421]) ^ (layer2_outputs[9947]));
    assign outputs[1465] = ~((layer2_outputs[7860]) ^ (layer2_outputs[1936]));
    assign outputs[1466] = ~(layer2_outputs[12528]);
    assign outputs[1467] = ~((layer2_outputs[11280]) | (layer2_outputs[10778]));
    assign outputs[1468] = (layer2_outputs[2960]) ^ (layer2_outputs[12082]);
    assign outputs[1469] = (layer2_outputs[10152]) ^ (layer2_outputs[9195]);
    assign outputs[1470] = ~(layer2_outputs[3170]);
    assign outputs[1471] = ~((layer2_outputs[7877]) ^ (layer2_outputs[2752]));
    assign outputs[1472] = ~(layer2_outputs[2506]);
    assign outputs[1473] = ~(layer2_outputs[1103]);
    assign outputs[1474] = ~((layer2_outputs[8989]) | (layer2_outputs[4291]));
    assign outputs[1475] = (layer2_outputs[958]) & ~(layer2_outputs[801]);
    assign outputs[1476] = ~((layer2_outputs[10713]) ^ (layer2_outputs[288]));
    assign outputs[1477] = ~((layer2_outputs[3227]) ^ (layer2_outputs[255]));
    assign outputs[1478] = (layer2_outputs[9758]) & (layer2_outputs[12087]);
    assign outputs[1479] = (layer2_outputs[3754]) & (layer2_outputs[9858]);
    assign outputs[1480] = ~((layer2_outputs[12207]) ^ (layer2_outputs[8074]));
    assign outputs[1481] = ~((layer2_outputs[459]) ^ (layer2_outputs[6955]));
    assign outputs[1482] = (layer2_outputs[7155]) ^ (layer2_outputs[7818]);
    assign outputs[1483] = ~((layer2_outputs[8571]) ^ (layer2_outputs[9926]));
    assign outputs[1484] = ~((layer2_outputs[3129]) ^ (layer2_outputs[9228]));
    assign outputs[1485] = ~(layer2_outputs[11905]);
    assign outputs[1486] = layer2_outputs[9845];
    assign outputs[1487] = 1'b0;
    assign outputs[1488] = (layer2_outputs[8354]) ^ (layer2_outputs[5639]);
    assign outputs[1489] = layer2_outputs[12461];
    assign outputs[1490] = (layer2_outputs[3805]) & ~(layer2_outputs[8469]);
    assign outputs[1491] = (layer2_outputs[2572]) & ~(layer2_outputs[11485]);
    assign outputs[1492] = layer2_outputs[3019];
    assign outputs[1493] = (layer2_outputs[8211]) & ~(layer2_outputs[10258]);
    assign outputs[1494] = layer2_outputs[6145];
    assign outputs[1495] = (layer2_outputs[5309]) & ~(layer2_outputs[149]);
    assign outputs[1496] = ~(layer2_outputs[3382]);
    assign outputs[1497] = (layer2_outputs[2654]) ^ (layer2_outputs[689]);
    assign outputs[1498] = ~(layer2_outputs[8768]);
    assign outputs[1499] = ~(layer2_outputs[9368]);
    assign outputs[1500] = layer2_outputs[8929];
    assign outputs[1501] = ~((layer2_outputs[323]) & (layer2_outputs[2159]));
    assign outputs[1502] = (layer2_outputs[11361]) & ~(layer2_outputs[5815]);
    assign outputs[1503] = (layer2_outputs[9016]) | (layer2_outputs[4896]);
    assign outputs[1504] = ~(layer2_outputs[3322]);
    assign outputs[1505] = ~((layer2_outputs[11591]) | (layer2_outputs[5638]));
    assign outputs[1506] = layer2_outputs[221];
    assign outputs[1507] = (layer2_outputs[7343]) & ~(layer2_outputs[290]);
    assign outputs[1508] = ~((layer2_outputs[1230]) ^ (layer2_outputs[10425]));
    assign outputs[1509] = (layer2_outputs[8987]) ^ (layer2_outputs[2459]);
    assign outputs[1510] = ~(layer2_outputs[698]);
    assign outputs[1511] = (layer2_outputs[6963]) ^ (layer2_outputs[12778]);
    assign outputs[1512] = ~(layer2_outputs[11174]);
    assign outputs[1513] = ~(layer2_outputs[3717]);
    assign outputs[1514] = layer2_outputs[4665];
    assign outputs[1515] = layer2_outputs[8503];
    assign outputs[1516] = ~((layer2_outputs[6611]) | (layer2_outputs[8117]));
    assign outputs[1517] = layer2_outputs[874];
    assign outputs[1518] = layer2_outputs[4942];
    assign outputs[1519] = ~((layer2_outputs[5731]) | (layer2_outputs[3875]));
    assign outputs[1520] = (layer2_outputs[6096]) & ~(layer2_outputs[11815]);
    assign outputs[1521] = ~((layer2_outputs[4409]) ^ (layer2_outputs[6541]));
    assign outputs[1522] = ~(layer2_outputs[3715]);
    assign outputs[1523] = ~(layer2_outputs[5831]);
    assign outputs[1524] = layer2_outputs[4471];
    assign outputs[1525] = (layer2_outputs[1358]) | (layer2_outputs[10933]);
    assign outputs[1526] = (layer2_outputs[1971]) & (layer2_outputs[10740]);
    assign outputs[1527] = (layer2_outputs[12745]) ^ (layer2_outputs[7561]);
    assign outputs[1528] = ~(layer2_outputs[5703]);
    assign outputs[1529] = ~((layer2_outputs[5429]) ^ (layer2_outputs[7653]));
    assign outputs[1530] = ~((layer2_outputs[1611]) ^ (layer2_outputs[8937]));
    assign outputs[1531] = ~(layer2_outputs[8205]);
    assign outputs[1532] = ~((layer2_outputs[8405]) ^ (layer2_outputs[962]));
    assign outputs[1533] = layer2_outputs[7601];
    assign outputs[1534] = ~((layer2_outputs[5893]) ^ (layer2_outputs[4681]));
    assign outputs[1535] = (layer2_outputs[7202]) ^ (layer2_outputs[2015]);
    assign outputs[1536] = (layer2_outputs[2024]) & ~(layer2_outputs[2343]);
    assign outputs[1537] = layer2_outputs[12662];
    assign outputs[1538] = ~((layer2_outputs[653]) ^ (layer2_outputs[6650]));
    assign outputs[1539] = (layer2_outputs[7057]) & ~(layer2_outputs[5010]);
    assign outputs[1540] = layer2_outputs[9866];
    assign outputs[1541] = ~((layer2_outputs[6384]) ^ (layer2_outputs[8138]));
    assign outputs[1542] = layer2_outputs[3043];
    assign outputs[1543] = ~((layer2_outputs[2524]) | (layer2_outputs[9542]));
    assign outputs[1544] = ~(layer2_outputs[11290]);
    assign outputs[1545] = ~((layer2_outputs[9606]) ^ (layer2_outputs[1514]));
    assign outputs[1546] = ~((layer2_outputs[4257]) ^ (layer2_outputs[10936]));
    assign outputs[1547] = layer2_outputs[6780];
    assign outputs[1548] = (layer2_outputs[7317]) & ~(layer2_outputs[12129]);
    assign outputs[1549] = ~((layer2_outputs[4404]) ^ (layer2_outputs[11117]));
    assign outputs[1550] = (layer2_outputs[2871]) & ~(layer2_outputs[523]);
    assign outputs[1551] = layer2_outputs[312];
    assign outputs[1552] = (layer2_outputs[12297]) ^ (layer2_outputs[2768]);
    assign outputs[1553] = (layer2_outputs[3692]) | (layer2_outputs[2520]);
    assign outputs[1554] = layer2_outputs[10054];
    assign outputs[1555] = (layer2_outputs[7720]) ^ (layer2_outputs[11798]);
    assign outputs[1556] = (layer2_outputs[9259]) & ~(layer2_outputs[7809]);
    assign outputs[1557] = (layer2_outputs[11121]) & ~(layer2_outputs[1541]);
    assign outputs[1558] = ~(layer2_outputs[10327]);
    assign outputs[1559] = layer2_outputs[11636];
    assign outputs[1560] = ~(layer2_outputs[4676]);
    assign outputs[1561] = (layer2_outputs[1023]) & ~(layer2_outputs[9806]);
    assign outputs[1562] = ~((layer2_outputs[901]) ^ (layer2_outputs[1803]));
    assign outputs[1563] = ~(layer2_outputs[1754]);
    assign outputs[1564] = (layer2_outputs[3859]) & ~(layer2_outputs[821]);
    assign outputs[1565] = layer2_outputs[2503];
    assign outputs[1566] = ~(layer2_outputs[5025]);
    assign outputs[1567] = ~(layer2_outputs[1926]);
    assign outputs[1568] = (layer2_outputs[12212]) ^ (layer2_outputs[8704]);
    assign outputs[1569] = (layer2_outputs[5084]) & ~(layer2_outputs[11751]);
    assign outputs[1570] = ~(layer2_outputs[4945]) | (layer2_outputs[12325]);
    assign outputs[1571] = (layer2_outputs[3870]) & ~(layer2_outputs[2197]);
    assign outputs[1572] = (layer2_outputs[1683]) & (layer2_outputs[3809]);
    assign outputs[1573] = layer2_outputs[4302];
    assign outputs[1574] = layer2_outputs[44];
    assign outputs[1575] = (layer2_outputs[4213]) & (layer2_outputs[9718]);
    assign outputs[1576] = (layer2_outputs[3947]) | (layer2_outputs[6266]);
    assign outputs[1577] = ~(layer2_outputs[1944]);
    assign outputs[1578] = (layer2_outputs[6486]) & (layer2_outputs[1706]);
    assign outputs[1579] = ~((layer2_outputs[9938]) | (layer2_outputs[161]));
    assign outputs[1580] = ~(layer2_outputs[4878]);
    assign outputs[1581] = ~((layer2_outputs[9791]) ^ (layer2_outputs[12272]));
    assign outputs[1582] = (layer2_outputs[8546]) ^ (layer2_outputs[5055]);
    assign outputs[1583] = ~(layer2_outputs[1906]);
    assign outputs[1584] = ~(layer2_outputs[945]);
    assign outputs[1585] = ~(layer2_outputs[1895]);
    assign outputs[1586] = (layer2_outputs[11112]) | (layer2_outputs[5818]);
    assign outputs[1587] = ~((layer2_outputs[8089]) ^ (layer2_outputs[67]));
    assign outputs[1588] = ~(layer2_outputs[4566]);
    assign outputs[1589] = ~(layer2_outputs[4722]);
    assign outputs[1590] = ~((layer2_outputs[4176]) ^ (layer2_outputs[1783]));
    assign outputs[1591] = (layer2_outputs[7616]) & ~(layer2_outputs[9827]);
    assign outputs[1592] = layer2_outputs[4796];
    assign outputs[1593] = ~(layer2_outputs[8821]);
    assign outputs[1594] = layer2_outputs[12002];
    assign outputs[1595] = layer2_outputs[7209];
    assign outputs[1596] = ~((layer2_outputs[10138]) ^ (layer2_outputs[3112]));
    assign outputs[1597] = ~(layer2_outputs[2578]);
    assign outputs[1598] = ~((layer2_outputs[109]) ^ (layer2_outputs[10320]));
    assign outputs[1599] = layer2_outputs[10453];
    assign outputs[1600] = ~((layer2_outputs[5413]) | (layer2_outputs[8536]));
    assign outputs[1601] = layer2_outputs[9501];
    assign outputs[1602] = (layer2_outputs[3068]) | (layer2_outputs[4718]);
    assign outputs[1603] = layer2_outputs[3782];
    assign outputs[1604] = ~(layer2_outputs[2342]);
    assign outputs[1605] = ~(layer2_outputs[2403]);
    assign outputs[1606] = (layer2_outputs[9528]) & (layer2_outputs[53]);
    assign outputs[1607] = layer2_outputs[12324];
    assign outputs[1608] = ~(layer2_outputs[6356]);
    assign outputs[1609] = ~((layer2_outputs[9393]) | (layer2_outputs[3832]));
    assign outputs[1610] = ~(layer2_outputs[11769]);
    assign outputs[1611] = ~(layer2_outputs[8152]);
    assign outputs[1612] = ~((layer2_outputs[7334]) | (layer2_outputs[2741]));
    assign outputs[1613] = ~(layer2_outputs[12449]) | (layer2_outputs[442]);
    assign outputs[1614] = (layer2_outputs[1665]) & ~(layer2_outputs[7590]);
    assign outputs[1615] = ~((layer2_outputs[596]) ^ (layer2_outputs[7777]));
    assign outputs[1616] = layer2_outputs[3548];
    assign outputs[1617] = layer2_outputs[8303];
    assign outputs[1618] = (layer2_outputs[8568]) & (layer2_outputs[6839]);
    assign outputs[1619] = ~((layer2_outputs[11358]) ^ (layer2_outputs[10324]));
    assign outputs[1620] = ~(layer2_outputs[2373]) | (layer2_outputs[832]);
    assign outputs[1621] = (layer2_outputs[6621]) & ~(layer2_outputs[10773]);
    assign outputs[1622] = ~(layer2_outputs[3071]);
    assign outputs[1623] = ~((layer2_outputs[11556]) ^ (layer2_outputs[9810]));
    assign outputs[1624] = ~(layer2_outputs[12775]);
    assign outputs[1625] = (layer2_outputs[5616]) ^ (layer2_outputs[5941]);
    assign outputs[1626] = (layer2_outputs[4323]) | (layer2_outputs[6473]);
    assign outputs[1627] = layer2_outputs[3606];
    assign outputs[1628] = (layer2_outputs[5073]) & (layer2_outputs[9932]);
    assign outputs[1629] = layer2_outputs[8454];
    assign outputs[1630] = (layer2_outputs[9165]) & ~(layer2_outputs[2000]);
    assign outputs[1631] = (layer2_outputs[12007]) ^ (layer2_outputs[6774]);
    assign outputs[1632] = layer2_outputs[8100];
    assign outputs[1633] = ~(layer2_outputs[7569]);
    assign outputs[1634] = (layer2_outputs[9609]) & ~(layer2_outputs[2325]);
    assign outputs[1635] = (layer2_outputs[5482]) ^ (layer2_outputs[11336]);
    assign outputs[1636] = ~(layer2_outputs[6408]) | (layer2_outputs[2416]);
    assign outputs[1637] = layer2_outputs[10047];
    assign outputs[1638] = ~((layer2_outputs[12140]) ^ (layer2_outputs[12520]));
    assign outputs[1639] = (layer2_outputs[970]) & (layer2_outputs[7209]);
    assign outputs[1640] = ~((layer2_outputs[10974]) ^ (layer2_outputs[8504]));
    assign outputs[1641] = (layer2_outputs[6580]) ^ (layer2_outputs[1376]);
    assign outputs[1642] = (layer2_outputs[8848]) ^ (layer2_outputs[2466]);
    assign outputs[1643] = ~(layer2_outputs[10759]);
    assign outputs[1644] = layer2_outputs[10506];
    assign outputs[1645] = ~((layer2_outputs[8925]) & (layer2_outputs[10166]));
    assign outputs[1646] = ~((layer2_outputs[358]) ^ (layer2_outputs[11269]));
    assign outputs[1647] = (layer2_outputs[578]) & (layer2_outputs[7520]);
    assign outputs[1648] = layer2_outputs[8336];
    assign outputs[1649] = ~(layer2_outputs[4579]);
    assign outputs[1650] = (layer2_outputs[9658]) ^ (layer2_outputs[9705]);
    assign outputs[1651] = layer2_outputs[7834];
    assign outputs[1652] = ~(layer2_outputs[1160]);
    assign outputs[1653] = ~((layer2_outputs[6759]) ^ (layer2_outputs[5774]));
    assign outputs[1654] = ~((layer2_outputs[8407]) ^ (layer2_outputs[11865]));
    assign outputs[1655] = ~((layer2_outputs[12079]) ^ (layer2_outputs[11360]));
    assign outputs[1656] = ~(layer2_outputs[12158]);
    assign outputs[1657] = ~((layer2_outputs[2470]) | (layer2_outputs[1500]));
    assign outputs[1658] = ~(layer2_outputs[4759]);
    assign outputs[1659] = ~(layer2_outputs[6890]);
    assign outputs[1660] = ~(layer2_outputs[10829]);
    assign outputs[1661] = (layer2_outputs[9237]) & ~(layer2_outputs[12006]);
    assign outputs[1662] = ~((layer2_outputs[2004]) ^ (layer2_outputs[2127]));
    assign outputs[1663] = (layer2_outputs[3289]) & (layer2_outputs[12366]);
    assign outputs[1664] = ~((layer2_outputs[7563]) | (layer2_outputs[6190]));
    assign outputs[1665] = (layer2_outputs[2002]) | (layer2_outputs[4378]);
    assign outputs[1666] = ~(layer2_outputs[7340]);
    assign outputs[1667] = ~(layer2_outputs[1299]);
    assign outputs[1668] = ~(layer2_outputs[3676]);
    assign outputs[1669] = ~(layer2_outputs[12012]);
    assign outputs[1670] = (layer2_outputs[2541]) & (layer2_outputs[10112]);
    assign outputs[1671] = (layer2_outputs[10320]) ^ (layer2_outputs[6103]);
    assign outputs[1672] = (layer2_outputs[11026]) & ~(layer2_outputs[4265]);
    assign outputs[1673] = ~(layer2_outputs[6648]);
    assign outputs[1674] = ~((layer2_outputs[9164]) ^ (layer2_outputs[1881]));
    assign outputs[1675] = (layer2_outputs[12521]) & ~(layer2_outputs[6739]);
    assign outputs[1676] = ~(layer2_outputs[6480]);
    assign outputs[1677] = ~(layer2_outputs[12572]);
    assign outputs[1678] = layer2_outputs[1883];
    assign outputs[1679] = (layer2_outputs[9732]) ^ (layer2_outputs[7640]);
    assign outputs[1680] = layer2_outputs[6086];
    assign outputs[1681] = (layer2_outputs[2034]) & (layer2_outputs[7878]);
    assign outputs[1682] = ~((layer2_outputs[10648]) ^ (layer2_outputs[2877]));
    assign outputs[1683] = (layer2_outputs[941]) & ~(layer2_outputs[1538]);
    assign outputs[1684] = (layer2_outputs[3816]) | (layer2_outputs[11629]);
    assign outputs[1685] = ~((layer2_outputs[8359]) & (layer2_outputs[8714]));
    assign outputs[1686] = (layer2_outputs[5159]) & (layer2_outputs[8387]);
    assign outputs[1687] = ~(layer2_outputs[8119]);
    assign outputs[1688] = ~(layer2_outputs[1299]);
    assign outputs[1689] = (layer2_outputs[1998]) & ~(layer2_outputs[9517]);
    assign outputs[1690] = layer2_outputs[9099];
    assign outputs[1691] = ~(layer2_outputs[3719]);
    assign outputs[1692] = ~(layer2_outputs[470]);
    assign outputs[1693] = ~(layer2_outputs[1461]);
    assign outputs[1694] = layer2_outputs[8600];
    assign outputs[1695] = ~((layer2_outputs[4017]) ^ (layer2_outputs[2403]));
    assign outputs[1696] = (layer2_outputs[11354]) ^ (layer2_outputs[12550]);
    assign outputs[1697] = ~((layer2_outputs[4051]) | (layer2_outputs[8945]));
    assign outputs[1698] = ~(layer2_outputs[7352]);
    assign outputs[1699] = ~((layer2_outputs[5891]) | (layer2_outputs[4970]));
    assign outputs[1700] = ~(layer2_outputs[3668]);
    assign outputs[1701] = ~((layer2_outputs[5087]) | (layer2_outputs[702]));
    assign outputs[1702] = ~(layer2_outputs[3834]);
    assign outputs[1703] = ~((layer2_outputs[2712]) | (layer2_outputs[11331]));
    assign outputs[1704] = ~((layer2_outputs[9837]) ^ (layer2_outputs[922]));
    assign outputs[1705] = (layer2_outputs[10252]) & ~(layer2_outputs[11856]);
    assign outputs[1706] = ~((layer2_outputs[1447]) ^ (layer2_outputs[4980]));
    assign outputs[1707] = layer2_outputs[124];
    assign outputs[1708] = layer2_outputs[11152];
    assign outputs[1709] = (layer2_outputs[8327]) & ~(layer2_outputs[1563]);
    assign outputs[1710] = (layer2_outputs[9714]) | (layer2_outputs[2696]);
    assign outputs[1711] = (layer2_outputs[3366]) & ~(layer2_outputs[2409]);
    assign outputs[1712] = ~(layer2_outputs[4885]);
    assign outputs[1713] = (layer2_outputs[1252]) & ~(layer2_outputs[9180]);
    assign outputs[1714] = layer2_outputs[7388];
    assign outputs[1715] = ~(layer2_outputs[11914]);
    assign outputs[1716] = layer2_outputs[12351];
    assign outputs[1717] = ~(layer2_outputs[12453]);
    assign outputs[1718] = layer2_outputs[12668];
    assign outputs[1719] = (layer2_outputs[11399]) & (layer2_outputs[7491]);
    assign outputs[1720] = ~((layer2_outputs[507]) ^ (layer2_outputs[6961]));
    assign outputs[1721] = ~((layer2_outputs[3333]) | (layer2_outputs[11033]));
    assign outputs[1722] = (layer2_outputs[6978]) & (layer2_outputs[3942]);
    assign outputs[1723] = (layer2_outputs[8220]) ^ (layer2_outputs[11205]);
    assign outputs[1724] = (layer2_outputs[10871]) ^ (layer2_outputs[11757]);
    assign outputs[1725] = ~(layer2_outputs[1943]);
    assign outputs[1726] = ~(layer2_outputs[1512]);
    assign outputs[1727] = (layer2_outputs[1611]) & ~(layer2_outputs[1274]);
    assign outputs[1728] = layer2_outputs[9046];
    assign outputs[1729] = ~(layer2_outputs[3438]);
    assign outputs[1730] = (layer2_outputs[2603]) ^ (layer2_outputs[12177]);
    assign outputs[1731] = layer2_outputs[10008];
    assign outputs[1732] = (layer2_outputs[8664]) & (layer2_outputs[4826]);
    assign outputs[1733] = layer2_outputs[4113];
    assign outputs[1734] = ~(layer2_outputs[8997]);
    assign outputs[1735] = (layer2_outputs[3016]) ^ (layer2_outputs[868]);
    assign outputs[1736] = (layer2_outputs[5010]) ^ (layer2_outputs[447]);
    assign outputs[1737] = layer2_outputs[3576];
    assign outputs[1738] = ~(layer2_outputs[8036]);
    assign outputs[1739] = ~(layer2_outputs[12050]);
    assign outputs[1740] = layer2_outputs[2619];
    assign outputs[1741] = layer2_outputs[10377];
    assign outputs[1742] = ~((layer2_outputs[1780]) & (layer2_outputs[8983]));
    assign outputs[1743] = (layer2_outputs[11832]) & (layer2_outputs[2371]);
    assign outputs[1744] = ~((layer2_outputs[7621]) ^ (layer2_outputs[7369]));
    assign outputs[1745] = (layer2_outputs[7691]) ^ (layer2_outputs[10968]);
    assign outputs[1746] = ~((layer2_outputs[1537]) ^ (layer2_outputs[11083]));
    assign outputs[1747] = ~((layer2_outputs[7177]) | (layer2_outputs[9074]));
    assign outputs[1748] = layer2_outputs[11472];
    assign outputs[1749] = ~((layer2_outputs[11873]) ^ (layer2_outputs[497]));
    assign outputs[1750] = (layer2_outputs[4597]) ^ (layer2_outputs[8474]);
    assign outputs[1751] = 1'b1;
    assign outputs[1752] = ~((layer2_outputs[1788]) ^ (layer2_outputs[5990]));
    assign outputs[1753] = ~(layer2_outputs[5065]);
    assign outputs[1754] = layer2_outputs[4072];
    assign outputs[1755] = ~(layer2_outputs[11253]);
    assign outputs[1756] = ~((layer2_outputs[3108]) | (layer2_outputs[5689]));
    assign outputs[1757] = (layer2_outputs[9222]) & (layer2_outputs[6082]);
    assign outputs[1758] = ~((layer2_outputs[8899]) ^ (layer2_outputs[1828]));
    assign outputs[1759] = ~(layer2_outputs[7818]);
    assign outputs[1760] = layer2_outputs[5242];
    assign outputs[1761] = ~((layer2_outputs[1058]) ^ (layer2_outputs[2548]));
    assign outputs[1762] = ~(layer2_outputs[6141]);
    assign outputs[1763] = layer2_outputs[7161];
    assign outputs[1764] = ~((layer2_outputs[4740]) | (layer2_outputs[6654]));
    assign outputs[1765] = ~(layer2_outputs[352]);
    assign outputs[1766] = (layer2_outputs[10149]) & (layer2_outputs[8303]);
    assign outputs[1767] = ~(layer2_outputs[10088]);
    assign outputs[1768] = (layer2_outputs[6011]) & (layer2_outputs[9556]);
    assign outputs[1769] = ~(layer2_outputs[10901]);
    assign outputs[1770] = (layer2_outputs[10101]) ^ (layer2_outputs[5094]);
    assign outputs[1771] = ~((layer2_outputs[7066]) ^ (layer2_outputs[5193]));
    assign outputs[1772] = (layer2_outputs[4975]) & (layer2_outputs[6206]);
    assign outputs[1773] = (layer2_outputs[4403]) & (layer2_outputs[7219]);
    assign outputs[1774] = ~((layer2_outputs[8782]) ^ (layer2_outputs[6628]));
    assign outputs[1775] = ~((layer2_outputs[7465]) ^ (layer2_outputs[9485]));
    assign outputs[1776] = ~(layer2_outputs[11930]);
    assign outputs[1777] = layer2_outputs[9239];
    assign outputs[1778] = layer2_outputs[3327];
    assign outputs[1779] = ~((layer2_outputs[10398]) ^ (layer2_outputs[6310]));
    assign outputs[1780] = (layer2_outputs[4700]) ^ (layer2_outputs[9455]);
    assign outputs[1781] = (layer2_outputs[1762]) ^ (layer2_outputs[1794]);
    assign outputs[1782] = (layer2_outputs[2353]) & ~(layer2_outputs[11563]);
    assign outputs[1783] = (layer2_outputs[6446]) ^ (layer2_outputs[2407]);
    assign outputs[1784] = ~(layer2_outputs[11928]);
    assign outputs[1785] = ~((layer2_outputs[157]) ^ (layer2_outputs[11887]));
    assign outputs[1786] = ~((layer2_outputs[6259]) | (layer2_outputs[9058]));
    assign outputs[1787] = ~(layer2_outputs[12162]);
    assign outputs[1788] = ~((layer2_outputs[3356]) | (layer2_outputs[5830]));
    assign outputs[1789] = ~(layer2_outputs[5717]);
    assign outputs[1790] = (layer2_outputs[2613]) ^ (layer2_outputs[1433]);
    assign outputs[1791] = (layer2_outputs[3771]) & ~(layer2_outputs[1697]);
    assign outputs[1792] = ~((layer2_outputs[11099]) | (layer2_outputs[4911]));
    assign outputs[1793] = layer2_outputs[2284];
    assign outputs[1794] = ~((layer2_outputs[272]) | (layer2_outputs[11093]));
    assign outputs[1795] = (layer2_outputs[3825]) & ~(layer2_outputs[12397]);
    assign outputs[1796] = (layer2_outputs[7485]) & (layer2_outputs[12741]);
    assign outputs[1797] = layer2_outputs[3177];
    assign outputs[1798] = (layer2_outputs[4774]) ^ (layer2_outputs[885]);
    assign outputs[1799] = (layer2_outputs[8095]) ^ (layer2_outputs[6642]);
    assign outputs[1800] = (layer2_outputs[1094]) ^ (layer2_outputs[6108]);
    assign outputs[1801] = ~((layer2_outputs[5155]) | (layer2_outputs[105]));
    assign outputs[1802] = (layer2_outputs[11938]) ^ (layer2_outputs[7225]);
    assign outputs[1803] = ~(layer2_outputs[5209]);
    assign outputs[1804] = ~(layer2_outputs[2172]);
    assign outputs[1805] = layer2_outputs[6421];
    assign outputs[1806] = ~((layer2_outputs[12315]) ^ (layer2_outputs[9187]));
    assign outputs[1807] = ~((layer2_outputs[10942]) | (layer2_outputs[8140]));
    assign outputs[1808] = layer2_outputs[12147];
    assign outputs[1809] = (layer2_outputs[742]) & ~(layer2_outputs[1866]);
    assign outputs[1810] = ~(layer2_outputs[1472]);
    assign outputs[1811] = ~(layer2_outputs[8252]);
    assign outputs[1812] = ~(layer2_outputs[6150]);
    assign outputs[1813] = (layer2_outputs[5981]) ^ (layer2_outputs[7421]);
    assign outputs[1814] = layer2_outputs[6621];
    assign outputs[1815] = ~(layer2_outputs[6656]);
    assign outputs[1816] = (layer2_outputs[1123]) ^ (layer2_outputs[9512]);
    assign outputs[1817] = (layer2_outputs[9389]) & ~(layer2_outputs[11689]);
    assign outputs[1818] = ~(layer2_outputs[1046]);
    assign outputs[1819] = (layer2_outputs[875]) ^ (layer2_outputs[12621]);
    assign outputs[1820] = ~(layer2_outputs[7017]) | (layer2_outputs[3366]);
    assign outputs[1821] = (layer2_outputs[5048]) ^ (layer2_outputs[11932]);
    assign outputs[1822] = ~((layer2_outputs[9188]) ^ (layer2_outputs[11420]));
    assign outputs[1823] = ~((layer2_outputs[7781]) | (layer2_outputs[3547]));
    assign outputs[1824] = (layer2_outputs[653]) & ~(layer2_outputs[1919]);
    assign outputs[1825] = ~((layer2_outputs[2443]) | (layer2_outputs[162]));
    assign outputs[1826] = ~((layer2_outputs[8417]) | (layer2_outputs[2054]));
    assign outputs[1827] = ~((layer2_outputs[10704]) | (layer2_outputs[9140]));
    assign outputs[1828] = ~(layer2_outputs[2692]);
    assign outputs[1829] = (layer2_outputs[10744]) ^ (layer2_outputs[5797]);
    assign outputs[1830] = ~((layer2_outputs[1400]) ^ (layer2_outputs[6691]));
    assign outputs[1831] = ~((layer2_outputs[8550]) ^ (layer2_outputs[7957]));
    assign outputs[1832] = layer2_outputs[5957];
    assign outputs[1833] = ~((layer2_outputs[1347]) | (layer2_outputs[11060]));
    assign outputs[1834] = layer2_outputs[3539];
    assign outputs[1835] = ~(layer2_outputs[3589]);
    assign outputs[1836] = ~(layer2_outputs[5369]);
    assign outputs[1837] = ~((layer2_outputs[7403]) ^ (layer2_outputs[4214]));
    assign outputs[1838] = layer2_outputs[8092];
    assign outputs[1839] = ~(layer2_outputs[1948]);
    assign outputs[1840] = ~((layer2_outputs[1401]) | (layer2_outputs[11886]));
    assign outputs[1841] = layer2_outputs[974];
    assign outputs[1842] = layer2_outputs[2693];
    assign outputs[1843] = ~(layer2_outputs[3574]);
    assign outputs[1844] = layer2_outputs[12573];
    assign outputs[1845] = layer2_outputs[7149];
    assign outputs[1846] = ~(layer2_outputs[516]);
    assign outputs[1847] = ~((layer2_outputs[1894]) ^ (layer2_outputs[758]));
    assign outputs[1848] = ~((layer2_outputs[3231]) ^ (layer2_outputs[5980]));
    assign outputs[1849] = ~(layer2_outputs[10476]);
    assign outputs[1850] = layer2_outputs[5564];
    assign outputs[1851] = (layer2_outputs[7804]) & (layer2_outputs[11187]);
    assign outputs[1852] = layer2_outputs[9646];
    assign outputs[1853] = layer2_outputs[7614];
    assign outputs[1854] = ~(layer2_outputs[1552]);
    assign outputs[1855] = (layer2_outputs[8052]) & (layer2_outputs[8588]);
    assign outputs[1856] = layer2_outputs[9014];
    assign outputs[1857] = layer2_outputs[10791];
    assign outputs[1858] = (layer2_outputs[9926]) ^ (layer2_outputs[6428]);
    assign outputs[1859] = ~((layer2_outputs[5261]) ^ (layer2_outputs[10762]));
    assign outputs[1860] = layer2_outputs[12502];
    assign outputs[1861] = (layer2_outputs[11131]) & (layer2_outputs[10681]);
    assign outputs[1862] = ~((layer2_outputs[4450]) ^ (layer2_outputs[4346]));
    assign outputs[1863] = (layer2_outputs[10187]) & (layer2_outputs[1266]);
    assign outputs[1864] = (layer2_outputs[9161]) & ~(layer2_outputs[11822]);
    assign outputs[1865] = layer2_outputs[9398];
    assign outputs[1866] = (layer2_outputs[3481]) ^ (layer2_outputs[7774]);
    assign outputs[1867] = ~((layer2_outputs[1590]) | (layer2_outputs[10014]));
    assign outputs[1868] = ~(layer2_outputs[420]);
    assign outputs[1869] = ~((layer2_outputs[1121]) | (layer2_outputs[1848]));
    assign outputs[1870] = layer2_outputs[6125];
    assign outputs[1871] = ~((layer2_outputs[1919]) ^ (layer2_outputs[10749]));
    assign outputs[1872] = ~(layer2_outputs[1010]);
    assign outputs[1873] = (layer2_outputs[6679]) ^ (layer2_outputs[325]);
    assign outputs[1874] = (layer2_outputs[7573]) ^ (layer2_outputs[5782]);
    assign outputs[1875] = ~((layer2_outputs[4246]) ^ (layer2_outputs[12072]));
    assign outputs[1876] = (layer2_outputs[7125]) & ~(layer2_outputs[9083]);
    assign outputs[1877] = ~((layer2_outputs[11507]) ^ (layer2_outputs[3065]));
    assign outputs[1878] = ~(layer2_outputs[691]);
    assign outputs[1879] = layer2_outputs[2828];
    assign outputs[1880] = ~(layer2_outputs[1310]);
    assign outputs[1881] = (layer2_outputs[1487]) & ~(layer2_outputs[7454]);
    assign outputs[1882] = ~(layer2_outputs[7337]);
    assign outputs[1883] = (layer2_outputs[7262]) & (layer2_outputs[12201]);
    assign outputs[1884] = (layer2_outputs[2663]) ^ (layer2_outputs[766]);
    assign outputs[1885] = ~((layer2_outputs[11695]) ^ (layer2_outputs[8524]));
    assign outputs[1886] = ~(layer2_outputs[7440]) | (layer2_outputs[1850]);
    assign outputs[1887] = ~(layer2_outputs[3890]);
    assign outputs[1888] = ~((layer2_outputs[9686]) ^ (layer2_outputs[6495]));
    assign outputs[1889] = (layer2_outputs[12084]) ^ (layer2_outputs[11335]);
    assign outputs[1890] = ~((layer2_outputs[3705]) ^ (layer2_outputs[4537]));
    assign outputs[1891] = (layer2_outputs[5221]) & ~(layer2_outputs[3189]);
    assign outputs[1892] = layer2_outputs[12587];
    assign outputs[1893] = ~(layer2_outputs[10763]);
    assign outputs[1894] = (layer2_outputs[431]) & (layer2_outputs[5748]);
    assign outputs[1895] = (layer2_outputs[1952]) & ~(layer2_outputs[10084]);
    assign outputs[1896] = (layer2_outputs[9643]) | (layer2_outputs[4211]);
    assign outputs[1897] = ~(layer2_outputs[6827]) | (layer2_outputs[6493]);
    assign outputs[1898] = ~((layer2_outputs[7182]) ^ (layer2_outputs[562]));
    assign outputs[1899] = ~(layer2_outputs[266]);
    assign outputs[1900] = (layer2_outputs[12666]) ^ (layer2_outputs[6037]);
    assign outputs[1901] = ~((layer2_outputs[10490]) | (layer2_outputs[7657]));
    assign outputs[1902] = (layer2_outputs[4379]) & ~(layer2_outputs[8751]);
    assign outputs[1903] = (layer2_outputs[2072]) ^ (layer2_outputs[1255]);
    assign outputs[1904] = ~(layer2_outputs[9485]);
    assign outputs[1905] = (layer2_outputs[10936]) ^ (layer2_outputs[2522]);
    assign outputs[1906] = ~(layer2_outputs[4006]);
    assign outputs[1907] = ~((layer2_outputs[2760]) | (layer2_outputs[4643]));
    assign outputs[1908] = ~((layer2_outputs[11561]) ^ (layer2_outputs[2322]));
    assign outputs[1909] = ~((layer2_outputs[6001]) | (layer2_outputs[684]));
    assign outputs[1910] = ~((layer2_outputs[11625]) | (layer2_outputs[2834]));
    assign outputs[1911] = (layer2_outputs[11982]) & ~(layer2_outputs[10080]);
    assign outputs[1912] = layer2_outputs[12567];
    assign outputs[1913] = ~((layer2_outputs[1834]) ^ (layer2_outputs[3524]));
    assign outputs[1914] = (layer2_outputs[10731]) ^ (layer2_outputs[5700]);
    assign outputs[1915] = (layer2_outputs[2710]) & ~(layer2_outputs[4673]);
    assign outputs[1916] = ~(layer2_outputs[4880]);
    assign outputs[1917] = ~(layer2_outputs[10737]);
    assign outputs[1918] = ~(layer2_outputs[983]);
    assign outputs[1919] = ~(layer2_outputs[12122]);
    assign outputs[1920] = layer2_outputs[7827];
    assign outputs[1921] = ~(layer2_outputs[10663]);
    assign outputs[1922] = layer2_outputs[7574];
    assign outputs[1923] = (layer2_outputs[9865]) ^ (layer2_outputs[10446]);
    assign outputs[1924] = ~((layer2_outputs[4172]) | (layer2_outputs[9859]));
    assign outputs[1925] = ~((layer2_outputs[10441]) ^ (layer2_outputs[8594]));
    assign outputs[1926] = layer2_outputs[5256];
    assign outputs[1927] = ~((layer2_outputs[11477]) ^ (layer2_outputs[12224]));
    assign outputs[1928] = ~(layer2_outputs[2961]);
    assign outputs[1929] = ~(layer2_outputs[2087]);
    assign outputs[1930] = (layer2_outputs[12764]) & ~(layer2_outputs[7099]);
    assign outputs[1931] = (layer2_outputs[4341]) & ~(layer2_outputs[9208]);
    assign outputs[1932] = ~((layer2_outputs[2685]) | (layer2_outputs[10087]));
    assign outputs[1933] = (layer2_outputs[12750]) & ~(layer2_outputs[9837]);
    assign outputs[1934] = ~((layer2_outputs[8850]) ^ (layer2_outputs[11938]));
    assign outputs[1935] = (layer2_outputs[7919]) ^ (layer2_outputs[2840]);
    assign outputs[1936] = layer2_outputs[4816];
    assign outputs[1937] = ~((layer2_outputs[9292]) ^ (layer2_outputs[7178]));
    assign outputs[1938] = ~((layer2_outputs[1108]) ^ (layer2_outputs[8159]));
    assign outputs[1939] = layer2_outputs[10651];
    assign outputs[1940] = layer2_outputs[12238];
    assign outputs[1941] = ~(layer2_outputs[9476]);
    assign outputs[1942] = (layer2_outputs[2596]) ^ (layer2_outputs[242]);
    assign outputs[1943] = ~((layer2_outputs[10231]) ^ (layer2_outputs[8946]));
    assign outputs[1944] = (layer2_outputs[8609]) ^ (layer2_outputs[9152]);
    assign outputs[1945] = (layer2_outputs[11803]) & (layer2_outputs[8855]);
    assign outputs[1946] = layer2_outputs[3367];
    assign outputs[1947] = (layer2_outputs[3702]) ^ (layer2_outputs[3063]);
    assign outputs[1948] = ~((layer2_outputs[3368]) ^ (layer2_outputs[12434]));
    assign outputs[1949] = layer2_outputs[995];
    assign outputs[1950] = ~(layer2_outputs[7693]);
    assign outputs[1951] = ~((layer2_outputs[12009]) ^ (layer2_outputs[7103]));
    assign outputs[1952] = (layer2_outputs[6355]) ^ (layer2_outputs[11061]);
    assign outputs[1953] = layer2_outputs[1526];
    assign outputs[1954] = ~((layer2_outputs[5974]) | (layer2_outputs[4759]));
    assign outputs[1955] = (layer2_outputs[7432]) & ~(layer2_outputs[1833]);
    assign outputs[1956] = ~(layer2_outputs[7890]);
    assign outputs[1957] = (layer2_outputs[7441]) & ~(layer2_outputs[2461]);
    assign outputs[1958] = ~((layer2_outputs[1999]) ^ (layer2_outputs[8310]));
    assign outputs[1959] = layer2_outputs[6970];
    assign outputs[1960] = ~((layer2_outputs[6191]) | (layer2_outputs[7942]));
    assign outputs[1961] = ~(layer2_outputs[3236]);
    assign outputs[1962] = ~(layer2_outputs[297]);
    assign outputs[1963] = layer2_outputs[7525];
    assign outputs[1964] = ~(layer2_outputs[7708]);
    assign outputs[1965] = ~((layer2_outputs[11801]) & (layer2_outputs[5390]));
    assign outputs[1966] = ~((layer2_outputs[77]) ^ (layer2_outputs[6836]));
    assign outputs[1967] = ~(layer2_outputs[8821]);
    assign outputs[1968] = ~((layer2_outputs[8597]) ^ (layer2_outputs[5291]));
    assign outputs[1969] = layer2_outputs[9588];
    assign outputs[1970] = (layer2_outputs[9866]) ^ (layer2_outputs[754]);
    assign outputs[1971] = ~(layer2_outputs[9796]);
    assign outputs[1972] = ~((layer2_outputs[1349]) ^ (layer2_outputs[3713]));
    assign outputs[1973] = ~(layer2_outputs[4252]);
    assign outputs[1974] = ~((layer2_outputs[8356]) | (layer2_outputs[714]));
    assign outputs[1975] = ~((layer2_outputs[5456]) & (layer2_outputs[5099]));
    assign outputs[1976] = ~((layer2_outputs[10368]) ^ (layer2_outputs[6748]));
    assign outputs[1977] = ~(layer2_outputs[9935]);
    assign outputs[1978] = layer2_outputs[4782];
    assign outputs[1979] = (layer2_outputs[2438]) & (layer2_outputs[9890]);
    assign outputs[1980] = layer2_outputs[8804];
    assign outputs[1981] = (layer2_outputs[4982]) & ~(layer2_outputs[2581]);
    assign outputs[1982] = ~((layer2_outputs[5515]) ^ (layer2_outputs[1525]));
    assign outputs[1983] = ~((layer2_outputs[436]) ^ (layer2_outputs[4708]));
    assign outputs[1984] = ~(layer2_outputs[4526]);
    assign outputs[1985] = (layer2_outputs[4770]) & (layer2_outputs[4230]);
    assign outputs[1986] = ~((layer2_outputs[4825]) | (layer2_outputs[2130]));
    assign outputs[1987] = (layer2_outputs[3403]) ^ (layer2_outputs[4939]);
    assign outputs[1988] = ~(layer2_outputs[1448]);
    assign outputs[1989] = ~(layer2_outputs[3384]) | (layer2_outputs[7775]);
    assign outputs[1990] = ~((layer2_outputs[9405]) ^ (layer2_outputs[5669]));
    assign outputs[1991] = (layer2_outputs[10865]) ^ (layer2_outputs[9474]);
    assign outputs[1992] = ~(layer2_outputs[8213]);
    assign outputs[1993] = ~((layer2_outputs[12207]) ^ (layer2_outputs[4987]));
    assign outputs[1994] = ~((layer2_outputs[2754]) ^ (layer2_outputs[121]));
    assign outputs[1995] = layer2_outputs[8388];
    assign outputs[1996] = (layer2_outputs[10049]) & ~(layer2_outputs[861]);
    assign outputs[1997] = (layer2_outputs[11797]) ^ (layer2_outputs[2041]);
    assign outputs[1998] = ~(layer2_outputs[11048]);
    assign outputs[1999] = layer2_outputs[8921];
    assign outputs[2000] = ~(layer2_outputs[7735]);
    assign outputs[2001] = ~((layer2_outputs[5676]) | (layer2_outputs[10428]));
    assign outputs[2002] = ~((layer2_outputs[1697]) | (layer2_outputs[7001]));
    assign outputs[2003] = layer2_outputs[4951];
    assign outputs[2004] = ~(layer2_outputs[8195]);
    assign outputs[2005] = ~(layer2_outputs[2157]);
    assign outputs[2006] = layer2_outputs[1092];
    assign outputs[2007] = (layer2_outputs[8355]) & ~(layer2_outputs[3257]);
    assign outputs[2008] = ~((layer2_outputs[9107]) | (layer2_outputs[6724]));
    assign outputs[2009] = ~(layer2_outputs[1063]);
    assign outputs[2010] = (layer2_outputs[5326]) & ~(layer2_outputs[4407]);
    assign outputs[2011] = ~(layer2_outputs[1604]);
    assign outputs[2012] = ~((layer2_outputs[8145]) | (layer2_outputs[7992]));
    assign outputs[2013] = ~(layer2_outputs[4886]);
    assign outputs[2014] = layer2_outputs[6068];
    assign outputs[2015] = ~(layer2_outputs[3150]);
    assign outputs[2016] = (layer2_outputs[5608]) & ~(layer2_outputs[1464]);
    assign outputs[2017] = (layer2_outputs[6861]) & ~(layer2_outputs[4831]);
    assign outputs[2018] = ~((layer2_outputs[83]) | (layer2_outputs[11465]));
    assign outputs[2019] = ~(layer2_outputs[11456]);
    assign outputs[2020] = layer2_outputs[9870];
    assign outputs[2021] = ~(layer2_outputs[11885]) | (layer2_outputs[9953]);
    assign outputs[2022] = layer2_outputs[1435];
    assign outputs[2023] = ~((layer2_outputs[1276]) | (layer2_outputs[528]));
    assign outputs[2024] = (layer2_outputs[6271]) ^ (layer2_outputs[12231]);
    assign outputs[2025] = ~(layer2_outputs[5076]);
    assign outputs[2026] = ~((layer2_outputs[10206]) | (layer2_outputs[7439]));
    assign outputs[2027] = layer2_outputs[4060];
    assign outputs[2028] = (layer2_outputs[7982]) ^ (layer2_outputs[7521]);
    assign outputs[2029] = layer2_outputs[4242];
    assign outputs[2030] = ~((layer2_outputs[1394]) ^ (layer2_outputs[7602]));
    assign outputs[2031] = (layer2_outputs[7112]) & ~(layer2_outputs[4468]);
    assign outputs[2032] = ~(layer2_outputs[12570]);
    assign outputs[2033] = (layer2_outputs[8149]) ^ (layer2_outputs[664]);
    assign outputs[2034] = layer2_outputs[4950];
    assign outputs[2035] = layer2_outputs[3554];
    assign outputs[2036] = layer2_outputs[5440];
    assign outputs[2037] = ~((layer2_outputs[3915]) | (layer2_outputs[6654]));
    assign outputs[2038] = ~((layer2_outputs[11659]) ^ (layer2_outputs[6768]));
    assign outputs[2039] = ~((layer2_outputs[284]) | (layer2_outputs[12625]));
    assign outputs[2040] = layer2_outputs[9785];
    assign outputs[2041] = ~(layer2_outputs[6448]);
    assign outputs[2042] = ~(layer2_outputs[10156]);
    assign outputs[2043] = ~((layer2_outputs[5144]) | (layer2_outputs[2942]));
    assign outputs[2044] = (layer2_outputs[4704]) & ~(layer2_outputs[10050]);
    assign outputs[2045] = (layer2_outputs[10585]) ^ (layer2_outputs[59]);
    assign outputs[2046] = ~((layer2_outputs[215]) ^ (layer2_outputs[9840]));
    assign outputs[2047] = ~(layer2_outputs[4866]);
    assign outputs[2048] = (layer2_outputs[9204]) & ~(layer2_outputs[11958]);
    assign outputs[2049] = layer2_outputs[6852];
    assign outputs[2050] = (layer2_outputs[5952]) ^ (layer2_outputs[12733]);
    assign outputs[2051] = (layer2_outputs[9853]) ^ (layer2_outputs[11357]);
    assign outputs[2052] = layer2_outputs[1673];
    assign outputs[2053] = ~((layer2_outputs[5026]) | (layer2_outputs[7655]));
    assign outputs[2054] = layer2_outputs[11788];
    assign outputs[2055] = ~(layer2_outputs[8275]);
    assign outputs[2056] = ~(layer2_outputs[11366]);
    assign outputs[2057] = (layer2_outputs[3632]) & ~(layer2_outputs[4220]);
    assign outputs[2058] = ~(layer2_outputs[6554]);
    assign outputs[2059] = layer2_outputs[749];
    assign outputs[2060] = ~((layer2_outputs[1176]) ^ (layer2_outputs[10976]));
    assign outputs[2061] = ~(layer2_outputs[3741]);
    assign outputs[2062] = (layer2_outputs[5409]) & (layer2_outputs[3985]);
    assign outputs[2063] = (layer2_outputs[3545]) & ~(layer2_outputs[11291]);
    assign outputs[2064] = (layer2_outputs[2446]) & (layer2_outputs[751]);
    assign outputs[2065] = layer2_outputs[5605];
    assign outputs[2066] = ~(layer2_outputs[5274]);
    assign outputs[2067] = (layer2_outputs[11835]) ^ (layer2_outputs[2481]);
    assign outputs[2068] = ~((layer2_outputs[799]) & (layer2_outputs[3729]));
    assign outputs[2069] = ~((layer2_outputs[12121]) | (layer2_outputs[6522]));
    assign outputs[2070] = ~((layer2_outputs[2326]) | (layer2_outputs[6609]));
    assign outputs[2071] = ~((layer2_outputs[10546]) ^ (layer2_outputs[6995]));
    assign outputs[2072] = ~((layer2_outputs[5910]) ^ (layer2_outputs[5863]));
    assign outputs[2073] = layer2_outputs[9615];
    assign outputs[2074] = layer2_outputs[10440];
    assign outputs[2075] = (layer2_outputs[4609]) & (layer2_outputs[4469]);
    assign outputs[2076] = (layer2_outputs[6099]) & ~(layer2_outputs[385]);
    assign outputs[2077] = (layer2_outputs[965]) ^ (layer2_outputs[9399]);
    assign outputs[2078] = layer2_outputs[8270];
    assign outputs[2079] = (layer2_outputs[6413]) & (layer2_outputs[11728]);
    assign outputs[2080] = ~(layer2_outputs[8413]);
    assign outputs[2081] = ~((layer2_outputs[6562]) | (layer2_outputs[11775]));
    assign outputs[2082] = layer2_outputs[6129];
    assign outputs[2083] = layer2_outputs[1815];
    assign outputs[2084] = (layer2_outputs[4560]) ^ (layer2_outputs[8507]);
    assign outputs[2085] = layer2_outputs[12065];
    assign outputs[2086] = (layer2_outputs[4084]) & ~(layer2_outputs[580]);
    assign outputs[2087] = ~(layer2_outputs[5015]);
    assign outputs[2088] = (layer2_outputs[4318]) & ~(layer2_outputs[8569]);
    assign outputs[2089] = layer2_outputs[6091];
    assign outputs[2090] = ~(layer2_outputs[6212]);
    assign outputs[2091] = (layer2_outputs[7428]) ^ (layer2_outputs[2893]);
    assign outputs[2092] = (layer2_outputs[4961]) & (layer2_outputs[8786]);
    assign outputs[2093] = (layer2_outputs[8400]) & ~(layer2_outputs[12163]);
    assign outputs[2094] = ~((layer2_outputs[6767]) ^ (layer2_outputs[11651]));
    assign outputs[2095] = ~(layer2_outputs[6316]);
    assign outputs[2096] = layer2_outputs[180];
    assign outputs[2097] = ~((layer2_outputs[4486]) ^ (layer2_outputs[4442]));
    assign outputs[2098] = ~((layer2_outputs[10123]) ^ (layer2_outputs[1718]));
    assign outputs[2099] = ~((layer2_outputs[4191]) ^ (layer2_outputs[8527]));
    assign outputs[2100] = (layer2_outputs[4045]) ^ (layer2_outputs[10694]);
    assign outputs[2101] = layer2_outputs[4384];
    assign outputs[2102] = layer2_outputs[9772];
    assign outputs[2103] = ~((layer2_outputs[11973]) | (layer2_outputs[5785]));
    assign outputs[2104] = ~(layer2_outputs[11134]);
    assign outputs[2105] = ~(layer2_outputs[7582]);
    assign outputs[2106] = ~((layer2_outputs[2043]) ^ (layer2_outputs[3592]));
    assign outputs[2107] = ~((layer2_outputs[11909]) ^ (layer2_outputs[1643]));
    assign outputs[2108] = ~((layer2_outputs[11751]) ^ (layer2_outputs[7656]));
    assign outputs[2109] = (layer2_outputs[4960]) & (layer2_outputs[8627]);
    assign outputs[2110] = (layer2_outputs[4097]) & ~(layer2_outputs[6529]);
    assign outputs[2111] = (layer2_outputs[4721]) | (layer2_outputs[5618]);
    assign outputs[2112] = layer2_outputs[3259];
    assign outputs[2113] = (layer2_outputs[8249]) & ~(layer2_outputs[1001]);
    assign outputs[2114] = (layer2_outputs[6675]) & ~(layer2_outputs[5982]);
    assign outputs[2115] = (layer2_outputs[12427]) | (layer2_outputs[9249]);
    assign outputs[2116] = ~(layer2_outputs[6714]);
    assign outputs[2117] = ~(layer2_outputs[1664]);
    assign outputs[2118] = layer2_outputs[9362];
    assign outputs[2119] = ~((layer2_outputs[10806]) ^ (layer2_outputs[9083]));
    assign outputs[2120] = (layer2_outputs[3208]) & (layer2_outputs[9398]);
    assign outputs[2121] = ~((layer2_outputs[4937]) | (layer2_outputs[11791]));
    assign outputs[2122] = layer2_outputs[8844];
    assign outputs[2123] = layer2_outputs[1153];
    assign outputs[2124] = (layer2_outputs[8625]) & ~(layer2_outputs[4236]);
    assign outputs[2125] = layer2_outputs[11561];
    assign outputs[2126] = ~(layer2_outputs[4339]);
    assign outputs[2127] = ~(layer2_outputs[7897]);
    assign outputs[2128] = ~((layer2_outputs[12769]) ^ (layer2_outputs[2275]));
    assign outputs[2129] = ~((layer2_outputs[8143]) ^ (layer2_outputs[423]));
    assign outputs[2130] = (layer2_outputs[2366]) ^ (layer2_outputs[820]);
    assign outputs[2131] = ~((layer2_outputs[5854]) ^ (layer2_outputs[11034]));
    assign outputs[2132] = ~((layer2_outputs[5148]) | (layer2_outputs[5812]));
    assign outputs[2133] = ~((layer2_outputs[8621]) ^ (layer2_outputs[5393]));
    assign outputs[2134] = (layer2_outputs[9052]) ^ (layer2_outputs[6322]);
    assign outputs[2135] = ~(layer2_outputs[9936]);
    assign outputs[2136] = (layer2_outputs[9148]) & ~(layer2_outputs[11066]);
    assign outputs[2137] = (layer2_outputs[7139]) & ~(layer2_outputs[1415]);
    assign outputs[2138] = ~((layer2_outputs[6356]) ^ (layer2_outputs[10482]));
    assign outputs[2139] = ~(layer2_outputs[10704]);
    assign outputs[2140] = ~(layer2_outputs[4301]);
    assign outputs[2141] = ~((layer2_outputs[1287]) ^ (layer2_outputs[5619]));
    assign outputs[2142] = (layer2_outputs[4844]) & ~(layer2_outputs[747]);
    assign outputs[2143] = (layer2_outputs[8783]) & (layer2_outputs[4427]);
    assign outputs[2144] = ~((layer2_outputs[4048]) ^ (layer2_outputs[4600]));
    assign outputs[2145] = ~(layer2_outputs[10226]);
    assign outputs[2146] = ~((layer2_outputs[6197]) ^ (layer2_outputs[583]));
    assign outputs[2147] = (layer2_outputs[9464]) ^ (layer2_outputs[4092]);
    assign outputs[2148] = (layer2_outputs[10365]) | (layer2_outputs[8189]);
    assign outputs[2149] = layer2_outputs[3816];
    assign outputs[2150] = (layer2_outputs[5998]) & (layer2_outputs[6289]);
    assign outputs[2151] = (layer2_outputs[9809]) & ~(layer2_outputs[4518]);
    assign outputs[2152] = layer2_outputs[6559];
    assign outputs[2153] = ~(layer2_outputs[8956]) | (layer2_outputs[3383]);
    assign outputs[2154] = ~(layer2_outputs[3578]);
    assign outputs[2155] = ~(layer2_outputs[536]);
    assign outputs[2156] = ~((layer2_outputs[7156]) | (layer2_outputs[5167]));
    assign outputs[2157] = ~((layer2_outputs[898]) | (layer2_outputs[3605]));
    assign outputs[2158] = (layer2_outputs[1728]) ^ (layer2_outputs[10003]);
    assign outputs[2159] = ~(layer2_outputs[6844]);
    assign outputs[2160] = ~((layer2_outputs[5842]) ^ (layer2_outputs[12026]));
    assign outputs[2161] = ~((layer2_outputs[2848]) ^ (layer2_outputs[2187]));
    assign outputs[2162] = layer2_outputs[4984];
    assign outputs[2163] = (layer2_outputs[1781]) & ~(layer2_outputs[10298]);
    assign outputs[2164] = (layer2_outputs[7500]) ^ (layer2_outputs[12374]);
    assign outputs[2165] = (layer2_outputs[4773]) & ~(layer2_outputs[2622]);
    assign outputs[2166] = ~(layer2_outputs[11676]);
    assign outputs[2167] = ~((layer2_outputs[1842]) ^ (layer2_outputs[1441]));
    assign outputs[2168] = (layer2_outputs[11193]) | (layer2_outputs[5468]);
    assign outputs[2169] = (layer2_outputs[5521]) & ~(layer2_outputs[11764]);
    assign outputs[2170] = ~(layer2_outputs[9630]);
    assign outputs[2171] = (layer2_outputs[10958]) ^ (layer2_outputs[6986]);
    assign outputs[2172] = ~((layer2_outputs[5165]) ^ (layer2_outputs[7758]));
    assign outputs[2173] = layer2_outputs[2586];
    assign outputs[2174] = ~(layer2_outputs[8212]);
    assign outputs[2175] = (layer2_outputs[5993]) ^ (layer2_outputs[3020]);
    assign outputs[2176] = ~((layer2_outputs[10719]) | (layer2_outputs[12153]));
    assign outputs[2177] = (layer2_outputs[2021]) & ~(layer2_outputs[8329]);
    assign outputs[2178] = (layer2_outputs[3632]) & (layer2_outputs[177]);
    assign outputs[2179] = (layer2_outputs[12661]) & ~(layer2_outputs[12676]);
    assign outputs[2180] = layer2_outputs[1772];
    assign outputs[2181] = layer2_outputs[4792];
    assign outputs[2182] = (layer2_outputs[305]) & ~(layer2_outputs[6043]);
    assign outputs[2183] = (layer2_outputs[1826]) & ~(layer2_outputs[6355]);
    assign outputs[2184] = ~(layer2_outputs[2319]);
    assign outputs[2185] = ~((layer2_outputs[10475]) ^ (layer2_outputs[5986]));
    assign outputs[2186] = (layer2_outputs[2162]) ^ (layer2_outputs[9242]);
    assign outputs[2187] = layer2_outputs[3514];
    assign outputs[2188] = ~(layer2_outputs[1702]);
    assign outputs[2189] = ~(layer2_outputs[9104]);
    assign outputs[2190] = (layer2_outputs[8670]) ^ (layer2_outputs[12689]);
    assign outputs[2191] = (layer2_outputs[5425]) ^ (layer2_outputs[921]);
    assign outputs[2192] = ~(layer2_outputs[2391]);
    assign outputs[2193] = layer2_outputs[3067];
    assign outputs[2194] = layer2_outputs[6556];
    assign outputs[2195] = ~((layer2_outputs[4601]) ^ (layer2_outputs[5097]));
    assign outputs[2196] = ~(layer2_outputs[1872]);
    assign outputs[2197] = (layer2_outputs[3029]) ^ (layer2_outputs[3443]);
    assign outputs[2198] = (layer2_outputs[10369]) ^ (layer2_outputs[3701]);
    assign outputs[2199] = (layer2_outputs[8294]) & (layer2_outputs[2555]);
    assign outputs[2200] = (layer2_outputs[10279]) & ~(layer2_outputs[3135]);
    assign outputs[2201] = ~(layer2_outputs[6546]);
    assign outputs[2202] = ~(layer2_outputs[12754]);
    assign outputs[2203] = ~(layer2_outputs[4578]);
    assign outputs[2204] = (layer2_outputs[5852]) & ~(layer2_outputs[1865]);
    assign outputs[2205] = layer2_outputs[2318];
    assign outputs[2206] = ~(layer2_outputs[2189]);
    assign outputs[2207] = (layer2_outputs[12790]) & ~(layer2_outputs[3560]);
    assign outputs[2208] = ~((layer2_outputs[10034]) ^ (layer2_outputs[9996]));
    assign outputs[2209] = (layer2_outputs[10621]) ^ (layer2_outputs[5775]);
    assign outputs[2210] = layer2_outputs[11736];
    assign outputs[2211] = ~(layer2_outputs[1990]) | (layer2_outputs[10019]);
    assign outputs[2212] = layer2_outputs[8539];
    assign outputs[2213] = ~(layer2_outputs[398]);
    assign outputs[2214] = (layer2_outputs[10049]) & ~(layer2_outputs[12137]);
    assign outputs[2215] = ~((layer2_outputs[7018]) ^ (layer2_outputs[5122]));
    assign outputs[2216] = (layer2_outputs[4041]) & (layer2_outputs[6560]);
    assign outputs[2217] = (layer2_outputs[11574]) & ~(layer2_outputs[96]);
    assign outputs[2218] = (layer2_outputs[233]) ^ (layer2_outputs[11077]);
    assign outputs[2219] = ~(layer2_outputs[8665]);
    assign outputs[2220] = ~(layer2_outputs[12175]);
    assign outputs[2221] = layer2_outputs[12471];
    assign outputs[2222] = (layer2_outputs[12498]) & (layer2_outputs[10918]);
    assign outputs[2223] = (layer2_outputs[2599]) & ~(layer2_outputs[2575]);
    assign outputs[2224] = (layer2_outputs[11098]) ^ (layer2_outputs[11668]);
    assign outputs[2225] = (layer2_outputs[4317]) ^ (layer2_outputs[11203]);
    assign outputs[2226] = layer2_outputs[2119];
    assign outputs[2227] = ~(layer2_outputs[3900]);
    assign outputs[2228] = ~(layer2_outputs[10919]);
    assign outputs[2229] = ~((layer2_outputs[2504]) | (layer2_outputs[8762]));
    assign outputs[2230] = (layer2_outputs[3199]) ^ (layer2_outputs[8691]);
    assign outputs[2231] = ~(layer2_outputs[8666]);
    assign outputs[2232] = ~(layer2_outputs[12559]);
    assign outputs[2233] = (layer2_outputs[1722]) & ~(layer2_outputs[10602]);
    assign outputs[2234] = (layer2_outputs[8779]) & ~(layer2_outputs[4662]);
    assign outputs[2235] = (layer2_outputs[6391]) & ~(layer2_outputs[7201]);
    assign outputs[2236] = (layer2_outputs[5427]) & (layer2_outputs[10058]);
    assign outputs[2237] = (layer2_outputs[2222]) & (layer2_outputs[8532]);
    assign outputs[2238] = ~(layer2_outputs[12215]);
    assign outputs[2239] = (layer2_outputs[5354]) ^ (layer2_outputs[8020]);
    assign outputs[2240] = ~(layer2_outputs[8517]);
    assign outputs[2241] = (layer2_outputs[8364]) & ~(layer2_outputs[4352]);
    assign outputs[2242] = (layer2_outputs[1172]) ^ (layer2_outputs[12024]);
    assign outputs[2243] = ~(layer2_outputs[3708]);
    assign outputs[2244] = (layer2_outputs[3120]) & ~(layer2_outputs[6921]);
    assign outputs[2245] = ~(layer2_outputs[12389]);
    assign outputs[2246] = (layer2_outputs[401]) & ~(layer2_outputs[4671]);
    assign outputs[2247] = (layer2_outputs[10264]) ^ (layer2_outputs[239]);
    assign outputs[2248] = (layer2_outputs[271]) & ~(layer2_outputs[11533]);
    assign outputs[2249] = layer2_outputs[5599];
    assign outputs[2250] = ~((layer2_outputs[10112]) ^ (layer2_outputs[11344]));
    assign outputs[2251] = layer2_outputs[5049];
    assign outputs[2252] = ~(layer2_outputs[4441]);
    assign outputs[2253] = ~(layer2_outputs[11040]);
    assign outputs[2254] = layer2_outputs[3838];
    assign outputs[2255] = ~(layer2_outputs[9614]);
    assign outputs[2256] = (layer2_outputs[7824]) & ~(layer2_outputs[7864]);
    assign outputs[2257] = ~(layer2_outputs[3407]);
    assign outputs[2258] = ~(layer2_outputs[7706]);
    assign outputs[2259] = ~(layer2_outputs[8676]);
    assign outputs[2260] = ~(layer2_outputs[1381]);
    assign outputs[2261] = layer2_outputs[5597];
    assign outputs[2262] = (layer2_outputs[7107]) & ~(layer2_outputs[8759]);
    assign outputs[2263] = layer2_outputs[7403];
    assign outputs[2264] = ~((layer2_outputs[1608]) ^ (layer2_outputs[2886]));
    assign outputs[2265] = (layer2_outputs[2117]) ^ (layer2_outputs[1906]);
    assign outputs[2266] = (layer2_outputs[5210]) ^ (layer2_outputs[7000]);
    assign outputs[2267] = (layer2_outputs[1032]) ^ (layer2_outputs[6302]);
    assign outputs[2268] = ~((layer2_outputs[6387]) ^ (layer2_outputs[4289]));
    assign outputs[2269] = (layer2_outputs[5561]) & (layer2_outputs[10386]);
    assign outputs[2270] = layer2_outputs[1576];
    assign outputs[2271] = ~((layer2_outputs[10561]) ^ (layer2_outputs[8913]));
    assign outputs[2272] = ~(layer2_outputs[12145]);
    assign outputs[2273] = ~((layer2_outputs[5435]) ^ (layer2_outputs[1247]));
    assign outputs[2274] = (layer2_outputs[2447]) ^ (layer2_outputs[5294]);
    assign outputs[2275] = layer2_outputs[12201];
    assign outputs[2276] = (layer2_outputs[10184]) ^ (layer2_outputs[2405]);
    assign outputs[2277] = ~((layer2_outputs[2093]) ^ (layer2_outputs[1004]));
    assign outputs[2278] = ~((layer2_outputs[4522]) ^ (layer2_outputs[5945]));
    assign outputs[2279] = ~(layer2_outputs[11795]);
    assign outputs[2280] = (layer2_outputs[8749]) ^ (layer2_outputs[2005]);
    assign outputs[2281] = (layer2_outputs[12495]) | (layer2_outputs[8427]);
    assign outputs[2282] = (layer2_outputs[11270]) ^ (layer2_outputs[4576]);
    assign outputs[2283] = layer2_outputs[1031];
    assign outputs[2284] = (layer2_outputs[1847]) | (layer2_outputs[2576]);
    assign outputs[2285] = ~(layer2_outputs[7297]) | (layer2_outputs[8251]);
    assign outputs[2286] = (layer2_outputs[1847]) | (layer2_outputs[4044]);
    assign outputs[2287] = ~((layer2_outputs[5392]) | (layer2_outputs[5312]));
    assign outputs[2288] = layer2_outputs[11276];
    assign outputs[2289] = ~(layer2_outputs[5194]);
    assign outputs[2290] = layer2_outputs[6863];
    assign outputs[2291] = layer2_outputs[10434];
    assign outputs[2292] = (layer2_outputs[12731]) & (layer2_outputs[6669]);
    assign outputs[2293] = (layer2_outputs[12454]) ^ (layer2_outputs[7391]);
    assign outputs[2294] = (layer2_outputs[1594]) & (layer2_outputs[8269]);
    assign outputs[2295] = (layer2_outputs[5323]) ^ (layer2_outputs[12576]);
    assign outputs[2296] = layer2_outputs[6326];
    assign outputs[2297] = ~((layer2_outputs[5646]) & (layer2_outputs[11149]));
    assign outputs[2298] = (layer2_outputs[5178]) ^ (layer2_outputs[126]);
    assign outputs[2299] = (layer2_outputs[7908]) ^ (layer2_outputs[5082]);
    assign outputs[2300] = (layer2_outputs[737]) & (layer2_outputs[3902]);
    assign outputs[2301] = layer2_outputs[658];
    assign outputs[2302] = layer2_outputs[9656];
    assign outputs[2303] = layer2_outputs[826];
    assign outputs[2304] = (layer2_outputs[3749]) ^ (layer2_outputs[82]);
    assign outputs[2305] = ~(layer2_outputs[11056]);
    assign outputs[2306] = ~(layer2_outputs[11960]);
    assign outputs[2307] = (layer2_outputs[2154]) ^ (layer2_outputs[10568]);
    assign outputs[2308] = (layer2_outputs[2616]) ^ (layer2_outputs[11823]);
    assign outputs[2309] = ~(layer2_outputs[1161]);
    assign outputs[2310] = ~(layer2_outputs[8477]);
    assign outputs[2311] = (layer2_outputs[3203]) ^ (layer2_outputs[9407]);
    assign outputs[2312] = ~((layer2_outputs[859]) ^ (layer2_outputs[8514]));
    assign outputs[2313] = (layer2_outputs[1293]) & (layer2_outputs[1886]);
    assign outputs[2314] = ~((layer2_outputs[5426]) ^ (layer2_outputs[11192]));
    assign outputs[2315] = layer2_outputs[8567];
    assign outputs[2316] = ~((layer2_outputs[3341]) & (layer2_outputs[1270]));
    assign outputs[2317] = (layer2_outputs[3807]) & (layer2_outputs[7149]);
    assign outputs[2318] = layer2_outputs[10926];
    assign outputs[2319] = ~(layer2_outputs[3380]);
    assign outputs[2320] = (layer2_outputs[4034]) ^ (layer2_outputs[2013]);
    assign outputs[2321] = (layer2_outputs[11639]) ^ (layer2_outputs[1603]);
    assign outputs[2322] = layer2_outputs[1470];
    assign outputs[2323] = ~((layer2_outputs[9373]) ^ (layer2_outputs[9098]));
    assign outputs[2324] = ~(layer2_outputs[5297]);
    assign outputs[2325] = (layer2_outputs[7675]) ^ (layer2_outputs[4211]);
    assign outputs[2326] = layer2_outputs[8361];
    assign outputs[2327] = ~(layer2_outputs[3376]);
    assign outputs[2328] = layer2_outputs[5715];
    assign outputs[2329] = ~(layer2_outputs[1373]);
    assign outputs[2330] = (layer2_outputs[5522]) & ~(layer2_outputs[169]);
    assign outputs[2331] = (layer2_outputs[6753]) & ~(layer2_outputs[8730]);
    assign outputs[2332] = (layer2_outputs[576]) ^ (layer2_outputs[2045]);
    assign outputs[2333] = layer2_outputs[9105];
    assign outputs[2334] = layer2_outputs[8740];
    assign outputs[2335] = ~((layer2_outputs[6279]) | (layer2_outputs[7195]));
    assign outputs[2336] = (layer2_outputs[3688]) & ~(layer2_outputs[2341]);
    assign outputs[2337] = (layer2_outputs[9339]) & (layer2_outputs[3436]);
    assign outputs[2338] = ~((layer2_outputs[42]) ^ (layer2_outputs[6188]));
    assign outputs[2339] = ~(layer2_outputs[3099]);
    assign outputs[2340] = (layer2_outputs[12029]) ^ (layer2_outputs[9363]);
    assign outputs[2341] = ~(layer2_outputs[9367]);
    assign outputs[2342] = (layer2_outputs[8629]) & (layer2_outputs[9311]);
    assign outputs[2343] = layer2_outputs[8341];
    assign outputs[2344] = ~(layer2_outputs[11298]);
    assign outputs[2345] = (layer2_outputs[4029]) ^ (layer2_outputs[8460]);
    assign outputs[2346] = layer2_outputs[9946];
    assign outputs[2347] = (layer2_outputs[6093]) & (layer2_outputs[1456]);
    assign outputs[2348] = ~(layer2_outputs[11037]);
    assign outputs[2349] = ~(layer2_outputs[11526]);
    assign outputs[2350] = layer2_outputs[10566];
    assign outputs[2351] = layer2_outputs[6232];
    assign outputs[2352] = ~(layer2_outputs[12241]);
    assign outputs[2353] = (layer2_outputs[11903]) ^ (layer2_outputs[11819]);
    assign outputs[2354] = ~(layer2_outputs[12485]);
    assign outputs[2355] = ~((layer2_outputs[8945]) | (layer2_outputs[11606]));
    assign outputs[2356] = layer2_outputs[12502];
    assign outputs[2357] = layer2_outputs[12048];
    assign outputs[2358] = ~(layer2_outputs[4645]);
    assign outputs[2359] = (layer2_outputs[12782]) ^ (layer2_outputs[4872]);
    assign outputs[2360] = ~((layer2_outputs[8134]) | (layer2_outputs[4593]));
    assign outputs[2361] = (layer2_outputs[5486]) & ~(layer2_outputs[6730]);
    assign outputs[2362] = (layer2_outputs[8907]) ^ (layer2_outputs[11311]);
    assign outputs[2363] = ~(layer2_outputs[9020]);
    assign outputs[2364] = layer2_outputs[257];
    assign outputs[2365] = ~(layer2_outputs[1457]);
    assign outputs[2366] = (layer2_outputs[1393]) & ~(layer2_outputs[733]);
    assign outputs[2367] = (layer2_outputs[11437]) & ~(layer2_outputs[8046]);
    assign outputs[2368] = layer2_outputs[7060];
    assign outputs[2369] = ~((layer2_outputs[6819]) ^ (layer2_outputs[7453]));
    assign outputs[2370] = ~(layer2_outputs[8072]);
    assign outputs[2371] = (layer2_outputs[9119]) & ~(layer2_outputs[1992]);
    assign outputs[2372] = (layer2_outputs[11601]) & ~(layer2_outputs[10860]);
    assign outputs[2373] = (layer2_outputs[2527]) ^ (layer2_outputs[1707]);
    assign outputs[2374] = layer2_outputs[4264];
    assign outputs[2375] = (layer2_outputs[3479]) & ~(layer2_outputs[4955]);
    assign outputs[2376] = ~((layer2_outputs[7475]) ^ (layer2_outputs[1915]));
    assign outputs[2377] = ~((layer2_outputs[3851]) | (layer2_outputs[10602]));
    assign outputs[2378] = (layer2_outputs[8286]) & ~(layer2_outputs[647]);
    assign outputs[2379] = (layer2_outputs[3554]) & ~(layer2_outputs[57]);
    assign outputs[2380] = (layer2_outputs[11605]) & (layer2_outputs[1814]);
    assign outputs[2381] = ~((layer2_outputs[9382]) ^ (layer2_outputs[5030]));
    assign outputs[2382] = ~(layer2_outputs[8853]);
    assign outputs[2383] = (layer2_outputs[4076]) ^ (layer2_outputs[5598]);
    assign outputs[2384] = ~((layer2_outputs[8155]) | (layer2_outputs[6317]));
    assign outputs[2385] = (layer2_outputs[3980]) & ~(layer2_outputs[12050]);
    assign outputs[2386] = (layer2_outputs[9835]) & ~(layer2_outputs[11002]);
    assign outputs[2387] = (layer2_outputs[4359]) ^ (layer2_outputs[12163]);
    assign outputs[2388] = ~(layer2_outputs[1492]);
    assign outputs[2389] = layer2_outputs[11713];
    assign outputs[2390] = (layer2_outputs[9244]) & ~(layer2_outputs[4336]);
    assign outputs[2391] = (layer2_outputs[4267]) ^ (layer2_outputs[10624]);
    assign outputs[2392] = ~((layer2_outputs[5399]) & (layer2_outputs[10606]));
    assign outputs[2393] = (layer2_outputs[5]) & (layer2_outputs[9941]);
    assign outputs[2394] = ~((layer2_outputs[11186]) | (layer2_outputs[4286]));
    assign outputs[2395] = (layer2_outputs[5014]) & ~(layer2_outputs[10866]);
    assign outputs[2396] = layer2_outputs[9566];
    assign outputs[2397] = ~(layer2_outputs[2276]);
    assign outputs[2398] = ~(layer2_outputs[7730]);
    assign outputs[2399] = ~((layer2_outputs[7361]) | (layer2_outputs[1000]));
    assign outputs[2400] = layer2_outputs[3565];
    assign outputs[2401] = ~((layer2_outputs[12114]) ^ (layer2_outputs[12421]));
    assign outputs[2402] = layer2_outputs[10078];
    assign outputs[2403] = (layer2_outputs[7691]) & ~(layer2_outputs[733]);
    assign outputs[2404] = ~(layer2_outputs[10214]);
    assign outputs[2405] = ~(layer2_outputs[9041]);
    assign outputs[2406] = (layer2_outputs[9281]) | (layer2_outputs[11715]);
    assign outputs[2407] = (layer2_outputs[5991]) & ~(layer2_outputs[9725]);
    assign outputs[2408] = ~(layer2_outputs[10635]);
    assign outputs[2409] = (layer2_outputs[4028]) | (layer2_outputs[11220]);
    assign outputs[2410] = ~(layer2_outputs[11660]);
    assign outputs[2411] = ~(layer2_outputs[928]);
    assign outputs[2412] = layer2_outputs[10228];
    assign outputs[2413] = ~((layer2_outputs[2227]) | (layer2_outputs[11464]));
    assign outputs[2414] = ~(layer2_outputs[11927]);
    assign outputs[2415] = (layer2_outputs[5168]) ^ (layer2_outputs[10917]);
    assign outputs[2416] = (layer2_outputs[7424]) & ~(layer2_outputs[1317]);
    assign outputs[2417] = ~(layer2_outputs[9213]);
    assign outputs[2418] = ~(layer2_outputs[5125]);
    assign outputs[2419] = (layer2_outputs[5664]) & ~(layer2_outputs[10701]);
    assign outputs[2420] = ~(layer2_outputs[10160]);
    assign outputs[2421] = layer2_outputs[10044];
    assign outputs[2422] = ~(layer2_outputs[5303]) | (layer2_outputs[10261]);
    assign outputs[2423] = ~(layer2_outputs[10428]);
    assign outputs[2424] = layer2_outputs[6660];
    assign outputs[2425] = ~(layer2_outputs[6856]);
    assign outputs[2426] = (layer2_outputs[8636]) ^ (layer2_outputs[2584]);
    assign outputs[2427] = (layer2_outputs[574]) ^ (layer2_outputs[5827]);
    assign outputs[2428] = ~(layer2_outputs[2791]);
    assign outputs[2429] = (layer2_outputs[11740]) & ~(layer2_outputs[6085]);
    assign outputs[2430] = (layer2_outputs[11401]) & ~(layer2_outputs[9729]);
    assign outputs[2431] = ~((layer2_outputs[8910]) | (layer2_outputs[9554]));
    assign outputs[2432] = ~(layer2_outputs[5090]);
    assign outputs[2433] = ~(layer2_outputs[10989]);
    assign outputs[2434] = layer2_outputs[2924];
    assign outputs[2435] = layer2_outputs[10758];
    assign outputs[2436] = (layer2_outputs[2673]) ^ (layer2_outputs[9287]);
    assign outputs[2437] = ~((layer2_outputs[9520]) | (layer2_outputs[5884]));
    assign outputs[2438] = (layer2_outputs[8825]) & ~(layer2_outputs[10523]);
    assign outputs[2439] = layer2_outputs[3486];
    assign outputs[2440] = (layer2_outputs[6946]) & ~(layer2_outputs[5609]);
    assign outputs[2441] = (layer2_outputs[639]) & ~(layer2_outputs[1257]);
    assign outputs[2442] = ~(layer2_outputs[9900]);
    assign outputs[2443] = (layer2_outputs[6637]) ^ (layer2_outputs[8699]);
    assign outputs[2444] = ~(layer2_outputs[5956]);
    assign outputs[2445] = 1'b0;
    assign outputs[2446] = layer2_outputs[5551];
    assign outputs[2447] = (layer2_outputs[8310]) ^ (layer2_outputs[11557]);
    assign outputs[2448] = ~(layer2_outputs[11767]) | (layer2_outputs[9752]);
    assign outputs[2449] = ~((layer2_outputs[3267]) ^ (layer2_outputs[6542]));
    assign outputs[2450] = ~((layer2_outputs[11070]) ^ (layer2_outputs[4771]));
    assign outputs[2451] = (layer2_outputs[5905]) & ~(layer2_outputs[691]);
    assign outputs[2452] = ~((layer2_outputs[10738]) | (layer2_outputs[3693]));
    assign outputs[2453] = (layer2_outputs[7371]) ^ (layer2_outputs[6515]);
    assign outputs[2454] = (layer2_outputs[1917]) & (layer2_outputs[3597]);
    assign outputs[2455] = ~(layer2_outputs[12033]);
    assign outputs[2456] = ~((layer2_outputs[12023]) ^ (layer2_outputs[619]));
    assign outputs[2457] = (layer2_outputs[9634]) & (layer2_outputs[852]);
    assign outputs[2458] = ~((layer2_outputs[12005]) ^ (layer2_outputs[1410]));
    assign outputs[2459] = (layer2_outputs[7752]) & (layer2_outputs[5995]);
    assign outputs[2460] = layer2_outputs[9655];
    assign outputs[2461] = (layer2_outputs[9788]) | (layer2_outputs[1679]);
    assign outputs[2462] = ~(layer2_outputs[6344]) | (layer2_outputs[1655]);
    assign outputs[2463] = ~(layer2_outputs[12168]);
    assign outputs[2464] = layer2_outputs[775];
    assign outputs[2465] = (layer2_outputs[12725]) & (layer2_outputs[6161]);
    assign outputs[2466] = layer2_outputs[2569];
    assign outputs[2467] = layer2_outputs[6469];
    assign outputs[2468] = ~(layer2_outputs[10176]);
    assign outputs[2469] = layer2_outputs[3173];
    assign outputs[2470] = ~((layer2_outputs[3834]) | (layer2_outputs[2456]));
    assign outputs[2471] = (layer2_outputs[10656]) & ~(layer2_outputs[4080]);
    assign outputs[2472] = (layer2_outputs[6866]) & ~(layer2_outputs[8620]);
    assign outputs[2473] = ~(layer2_outputs[9886]);
    assign outputs[2474] = layer2_outputs[5374];
    assign outputs[2475] = layer2_outputs[3043];
    assign outputs[2476] = (layer2_outputs[5944]) & ~(layer2_outputs[8967]);
    assign outputs[2477] = ~(layer2_outputs[695]);
    assign outputs[2478] = ~(layer2_outputs[12006]);
    assign outputs[2479] = ~((layer2_outputs[361]) ^ (layer2_outputs[3435]));
    assign outputs[2480] = (layer2_outputs[1009]) & ~(layer2_outputs[7186]);
    assign outputs[2481] = ~(layer2_outputs[10387]);
    assign outputs[2482] = (layer2_outputs[12281]) ^ (layer2_outputs[12104]);
    assign outputs[2483] = (layer2_outputs[3092]) ^ (layer2_outputs[12447]);
    assign outputs[2484] = (layer2_outputs[11444]) ^ (layer2_outputs[9105]);
    assign outputs[2485] = (layer2_outputs[8652]) & ~(layer2_outputs[8153]);
    assign outputs[2486] = (layer2_outputs[6113]) ^ (layer2_outputs[9899]);
    assign outputs[2487] = (layer2_outputs[3738]) & ~(layer2_outputs[3756]);
    assign outputs[2488] = (layer2_outputs[11020]) ^ (layer2_outputs[6892]);
    assign outputs[2489] = ~((layer2_outputs[2792]) ^ (layer2_outputs[4947]));
    assign outputs[2490] = (layer2_outputs[1644]) & ~(layer2_outputs[8058]);
    assign outputs[2491] = (layer2_outputs[8811]) & ~(layer2_outputs[11935]);
    assign outputs[2492] = (layer2_outputs[11969]) ^ (layer2_outputs[1739]);
    assign outputs[2493] = ~(layer2_outputs[11711]);
    assign outputs[2494] = ~(layer2_outputs[4142]);
    assign outputs[2495] = (layer2_outputs[10706]) & (layer2_outputs[3889]);
    assign outputs[2496] = ~((layer2_outputs[9949]) ^ (layer2_outputs[991]));
    assign outputs[2497] = ~((layer2_outputs[11594]) ^ (layer2_outputs[8077]));
    assign outputs[2498] = ~((layer2_outputs[11325]) | (layer2_outputs[5030]));
    assign outputs[2499] = (layer2_outputs[2725]) ^ (layer2_outputs[2245]);
    assign outputs[2500] = (layer2_outputs[6838]) & ~(layer2_outputs[5136]);
    assign outputs[2501] = ~((layer2_outputs[7682]) ^ (layer2_outputs[8896]));
    assign outputs[2502] = layer2_outputs[8948];
    assign outputs[2503] = ~(layer2_outputs[9351]);
    assign outputs[2504] = ~((layer2_outputs[5197]) ^ (layer2_outputs[11339]));
    assign outputs[2505] = ~(layer2_outputs[10955]);
    assign outputs[2506] = ~(layer2_outputs[2487]);
    assign outputs[2507] = layer2_outputs[6772];
    assign outputs[2508] = ~((layer2_outputs[3054]) ^ (layer2_outputs[1845]));
    assign outputs[2509] = ~((layer2_outputs[7902]) | (layer2_outputs[6904]));
    assign outputs[2510] = (layer2_outputs[6406]) & ~(layer2_outputs[7178]);
    assign outputs[2511] = ~((layer2_outputs[12278]) ^ (layer2_outputs[7074]));
    assign outputs[2512] = ~((layer2_outputs[2124]) ^ (layer2_outputs[1104]));
    assign outputs[2513] = (layer2_outputs[2149]) & ~(layer2_outputs[4809]);
    assign outputs[2514] = ~((layer2_outputs[3010]) | (layer2_outputs[4502]));
    assign outputs[2515] = ~(layer2_outputs[9424]);
    assign outputs[2516] = (layer2_outputs[7085]) & (layer2_outputs[4076]);
    assign outputs[2517] = layer2_outputs[7703];
    assign outputs[2518] = (layer2_outputs[10074]) & ~(layer2_outputs[1171]);
    assign outputs[2519] = ~((layer2_outputs[4523]) ^ (layer2_outputs[6510]));
    assign outputs[2520] = layer2_outputs[12613];
    assign outputs[2521] = ~((layer2_outputs[2291]) ^ (layer2_outputs[3746]));
    assign outputs[2522] = ~(layer2_outputs[2206]);
    assign outputs[2523] = (layer2_outputs[6506]) ^ (layer2_outputs[705]);
    assign outputs[2524] = layer2_outputs[10238];
    assign outputs[2525] = ~((layer2_outputs[2899]) ^ (layer2_outputs[6935]));
    assign outputs[2526] = layer2_outputs[38];
    assign outputs[2527] = ~(layer2_outputs[10277]);
    assign outputs[2528] = (layer2_outputs[8169]) & ~(layer2_outputs[11612]);
    assign outputs[2529] = (layer2_outputs[8075]) ^ (layer2_outputs[6937]);
    assign outputs[2530] = layer2_outputs[8739];
    assign outputs[2531] = (layer2_outputs[8562]) ^ (layer2_outputs[2708]);
    assign outputs[2532] = layer2_outputs[7698];
    assign outputs[2533] = (layer2_outputs[1745]) ^ (layer2_outputs[3938]);
    assign outputs[2534] = ~((layer2_outputs[3912]) ^ (layer2_outputs[8818]));
    assign outputs[2535] = layer2_outputs[4689];
    assign outputs[2536] = layer2_outputs[203];
    assign outputs[2537] = ~((layer2_outputs[2350]) & (layer2_outputs[3470]));
    assign outputs[2538] = ~((layer2_outputs[2173]) | (layer2_outputs[8158]));
    assign outputs[2539] = (layer2_outputs[4412]) & ~(layer2_outputs[9699]);
    assign outputs[2540] = ~((layer2_outputs[470]) & (layer2_outputs[1070]));
    assign outputs[2541] = layer2_outputs[6751];
    assign outputs[2542] = ~((layer2_outputs[4022]) ^ (layer2_outputs[9719]));
    assign outputs[2543] = (layer2_outputs[9879]) ^ (layer2_outputs[3494]);
    assign outputs[2544] = layer2_outputs[5242];
    assign outputs[2545] = ~((layer2_outputs[503]) ^ (layer2_outputs[10460]));
    assign outputs[2546] = layer2_outputs[3942];
    assign outputs[2547] = ~(layer2_outputs[3715]) | (layer2_outputs[7527]);
    assign outputs[2548] = ~((layer2_outputs[1817]) ^ (layer2_outputs[5753]));
    assign outputs[2549] = (layer2_outputs[4246]) ^ (layer2_outputs[10992]);
    assign outputs[2550] = ~((layer2_outputs[11282]) | (layer2_outputs[748]));
    assign outputs[2551] = ~((layer2_outputs[1088]) ^ (layer2_outputs[3187]));
    assign outputs[2552] = (layer2_outputs[5149]) ^ (layer2_outputs[36]);
    assign outputs[2553] = ~((layer2_outputs[9363]) ^ (layer2_outputs[4608]));
    assign outputs[2554] = layer2_outputs[5112];
    assign outputs[2555] = ~((layer2_outputs[6447]) ^ (layer2_outputs[10487]));
    assign outputs[2556] = ~((layer2_outputs[2369]) ^ (layer2_outputs[10162]));
    assign outputs[2557] = ~(layer2_outputs[11382]);
    assign outputs[2558] = layer2_outputs[7509];
    assign outputs[2559] = ~(layer2_outputs[11620]);
    assign outputs[2560] = ~(layer2_outputs[7056]);
    assign outputs[2561] = layer2_outputs[9161];
    assign outputs[2562] = ~((layer2_outputs[11194]) ^ (layer2_outputs[4170]));
    assign outputs[2563] = (layer2_outputs[4406]) & (layer2_outputs[10265]);
    assign outputs[2564] = ~(layer2_outputs[7807]) | (layer2_outputs[491]);
    assign outputs[2565] = ~(layer2_outputs[11094]);
    assign outputs[2566] = layer2_outputs[3000];
    assign outputs[2567] = ~((layer2_outputs[7395]) ^ (layer2_outputs[11946]));
    assign outputs[2568] = (layer2_outputs[1167]) ^ (layer2_outputs[2732]);
    assign outputs[2569] = ~(layer2_outputs[6594]);
    assign outputs[2570] = layer2_outputs[3925];
    assign outputs[2571] = ~(layer2_outputs[1206]) | (layer2_outputs[10447]);
    assign outputs[2572] = ~(layer2_outputs[1653]);
    assign outputs[2573] = layer2_outputs[1172];
    assign outputs[2574] = ~((layer2_outputs[11950]) & (layer2_outputs[1532]));
    assign outputs[2575] = (layer2_outputs[886]) & (layer2_outputs[7852]);
    assign outputs[2576] = ~((layer2_outputs[1474]) ^ (layer2_outputs[5973]));
    assign outputs[2577] = ~((layer2_outputs[3491]) ^ (layer2_outputs[3242]));
    assign outputs[2578] = ~(layer2_outputs[11106]);
    assign outputs[2579] = ~(layer2_outputs[9156]) | (layer2_outputs[2052]);
    assign outputs[2580] = ~(layer2_outputs[1179]);
    assign outputs[2581] = (layer2_outputs[8239]) | (layer2_outputs[9753]);
    assign outputs[2582] = layer2_outputs[6353];
    assign outputs[2583] = (layer2_outputs[1841]) | (layer2_outputs[732]);
    assign outputs[2584] = ~(layer2_outputs[6157]);
    assign outputs[2585] = ~((layer2_outputs[3443]) ^ (layer2_outputs[2788]));
    assign outputs[2586] = ~(layer2_outputs[2851]);
    assign outputs[2587] = ~(layer2_outputs[10835]) | (layer2_outputs[2714]);
    assign outputs[2588] = (layer2_outputs[12412]) ^ (layer2_outputs[7994]);
    assign outputs[2589] = ~((layer2_outputs[5966]) ^ (layer2_outputs[3595]));
    assign outputs[2590] = layer2_outputs[7174];
    assign outputs[2591] = ~(layer2_outputs[10458]);
    assign outputs[2592] = ~(layer2_outputs[9084]);
    assign outputs[2593] = ~(layer2_outputs[2870]);
    assign outputs[2594] = ~(layer2_outputs[5338]) | (layer2_outputs[6552]);
    assign outputs[2595] = ~(layer2_outputs[2586]);
    assign outputs[2596] = layer2_outputs[648];
    assign outputs[2597] = layer2_outputs[4808];
    assign outputs[2598] = (layer2_outputs[12121]) & ~(layer2_outputs[10040]);
    assign outputs[2599] = ~(layer2_outputs[1937]);
    assign outputs[2600] = ~(layer2_outputs[7124]);
    assign outputs[2601] = ~((layer2_outputs[7960]) | (layer2_outputs[1338]));
    assign outputs[2602] = ~((layer2_outputs[7184]) ^ (layer2_outputs[6809]));
    assign outputs[2603] = ~(layer2_outputs[8291]);
    assign outputs[2604] = ~((layer2_outputs[9174]) ^ (layer2_outputs[3052]));
    assign outputs[2605] = (layer2_outputs[7454]) ^ (layer2_outputs[1712]);
    assign outputs[2606] = ~(layer2_outputs[8077]) | (layer2_outputs[5602]);
    assign outputs[2607] = layer2_outputs[3222];
    assign outputs[2608] = ~(layer2_outputs[4455]);
    assign outputs[2609] = layer2_outputs[8638];
    assign outputs[2610] = ~(layer2_outputs[3713]) | (layer2_outputs[519]);
    assign outputs[2611] = (layer2_outputs[354]) ^ (layer2_outputs[3933]);
    assign outputs[2612] = (layer2_outputs[9510]) & (layer2_outputs[9973]);
    assign outputs[2613] = ~((layer2_outputs[6828]) ^ (layer2_outputs[2887]));
    assign outputs[2614] = (layer2_outputs[10820]) & ~(layer2_outputs[1292]);
    assign outputs[2615] = ~((layer2_outputs[8771]) ^ (layer2_outputs[12491]));
    assign outputs[2616] = ~(layer2_outputs[53]);
    assign outputs[2617] = layer2_outputs[7556];
    assign outputs[2618] = ~((layer2_outputs[6160]) | (layer2_outputs[9583]));
    assign outputs[2619] = ~(layer2_outputs[9538]);
    assign outputs[2620] = ~((layer2_outputs[3402]) ^ (layer2_outputs[618]));
    assign outputs[2621] = layer2_outputs[6523];
    assign outputs[2622] = layer2_outputs[1868];
    assign outputs[2623] = (layer2_outputs[6154]) ^ (layer2_outputs[5548]);
    assign outputs[2624] = ~((layer2_outputs[3304]) ^ (layer2_outputs[7394]));
    assign outputs[2625] = layer2_outputs[5004];
    assign outputs[2626] = (layer2_outputs[3151]) | (layer2_outputs[2217]);
    assign outputs[2627] = ~(layer2_outputs[1229]);
    assign outputs[2628] = ~(layer2_outputs[7558]);
    assign outputs[2629] = (layer2_outputs[10657]) ^ (layer2_outputs[11267]);
    assign outputs[2630] = layer2_outputs[4483];
    assign outputs[2631] = ~(layer2_outputs[2481]);
    assign outputs[2632] = ~(layer2_outputs[4231]);
    assign outputs[2633] = layer2_outputs[4592];
    assign outputs[2634] = (layer2_outputs[11867]) ^ (layer2_outputs[9659]);
    assign outputs[2635] = ~(layer2_outputs[4258]);
    assign outputs[2636] = layer2_outputs[12587];
    assign outputs[2637] = ~((layer2_outputs[12683]) ^ (layer2_outputs[6701]));
    assign outputs[2638] = layer2_outputs[6041];
    assign outputs[2639] = ~(layer2_outputs[2253]);
    assign outputs[2640] = ~(layer2_outputs[11265]);
    assign outputs[2641] = ~((layer2_outputs[12312]) ^ (layer2_outputs[7853]));
    assign outputs[2642] = layer2_outputs[9195];
    assign outputs[2643] = ~((layer2_outputs[3600]) ^ (layer2_outputs[7020]));
    assign outputs[2644] = ~(layer2_outputs[12578]);
    assign outputs[2645] = ~(layer2_outputs[3265]) | (layer2_outputs[2131]);
    assign outputs[2646] = layer2_outputs[12146];
    assign outputs[2647] = ~((layer2_outputs[558]) ^ (layer2_outputs[9436]));
    assign outputs[2648] = ~(layer2_outputs[1726]);
    assign outputs[2649] = ~(layer2_outputs[5990]);
    assign outputs[2650] = (layer2_outputs[8195]) & ~(layer2_outputs[2068]);
    assign outputs[2651] = ~(layer2_outputs[6734]);
    assign outputs[2652] = ~((layer2_outputs[6569]) ^ (layer2_outputs[7943]));
    assign outputs[2653] = ~(layer2_outputs[8060]) | (layer2_outputs[3487]);
    assign outputs[2654] = ~(layer2_outputs[9340]) | (layer2_outputs[11566]);
    assign outputs[2655] = layer2_outputs[11915];
    assign outputs[2656] = (layer2_outputs[9964]) | (layer2_outputs[10941]);
    assign outputs[2657] = ~(layer2_outputs[8824]);
    assign outputs[2658] = ~(layer2_outputs[9766]);
    assign outputs[2659] = ~(layer2_outputs[11418]);
    assign outputs[2660] = ~(layer2_outputs[11992]);
    assign outputs[2661] = (layer2_outputs[1511]) & ~(layer2_outputs[146]);
    assign outputs[2662] = ~((layer2_outputs[3076]) ^ (layer2_outputs[11383]));
    assign outputs[2663] = ~((layer2_outputs[2192]) ^ (layer2_outputs[11272]));
    assign outputs[2664] = ~((layer2_outputs[1286]) ^ (layer2_outputs[723]));
    assign outputs[2665] = (layer2_outputs[918]) | (layer2_outputs[2480]);
    assign outputs[2666] = (layer2_outputs[3245]) ^ (layer2_outputs[2211]);
    assign outputs[2667] = layer2_outputs[11386];
    assign outputs[2668] = layer2_outputs[5002];
    assign outputs[2669] = ~(layer2_outputs[7088]);
    assign outputs[2670] = ~(layer2_outputs[2136]);
    assign outputs[2671] = ~(layer2_outputs[10531]);
    assign outputs[2672] = (layer2_outputs[5938]) ^ (layer2_outputs[6321]);
    assign outputs[2673] = layer2_outputs[4698];
    assign outputs[2674] = ~(layer2_outputs[1600]);
    assign outputs[2675] = layer2_outputs[7793];
    assign outputs[2676] = ~(layer2_outputs[3851]);
    assign outputs[2677] = (layer2_outputs[6662]) ^ (layer2_outputs[12644]);
    assign outputs[2678] = ~((layer2_outputs[1154]) ^ (layer2_outputs[8960]));
    assign outputs[2679] = ~(layer2_outputs[4714]) | (layer2_outputs[8822]);
    assign outputs[2680] = ~(layer2_outputs[8284]) | (layer2_outputs[3496]);
    assign outputs[2681] = (layer2_outputs[2805]) ^ (layer2_outputs[566]);
    assign outputs[2682] = layer2_outputs[12518];
    assign outputs[2683] = ~((layer2_outputs[12706]) ^ (layer2_outputs[7059]));
    assign outputs[2684] = ~(layer2_outputs[6111]);
    assign outputs[2685] = ~(layer2_outputs[10961]);
    assign outputs[2686] = ~(layer2_outputs[11564]);
    assign outputs[2687] = (layer2_outputs[1445]) & (layer2_outputs[6968]);
    assign outputs[2688] = layer2_outputs[9294];
    assign outputs[2689] = ~(layer2_outputs[6571]);
    assign outputs[2690] = layer2_outputs[4188];
    assign outputs[2691] = (layer2_outputs[2973]) ^ (layer2_outputs[2559]);
    assign outputs[2692] = ~(layer2_outputs[7796]);
    assign outputs[2693] = (layer2_outputs[6807]) ^ (layer2_outputs[750]);
    assign outputs[2694] = layer2_outputs[2032];
    assign outputs[2695] = layer2_outputs[9421];
    assign outputs[2696] = ~((layer2_outputs[10692]) & (layer2_outputs[7637]));
    assign outputs[2697] = ~(layer2_outputs[9723]);
    assign outputs[2698] = ~((layer2_outputs[8891]) & (layer2_outputs[12486]));
    assign outputs[2699] = layer2_outputs[10332];
    assign outputs[2700] = (layer2_outputs[3164]) | (layer2_outputs[10454]);
    assign outputs[2701] = (layer2_outputs[8334]) & (layer2_outputs[10580]);
    assign outputs[2702] = ~(layer2_outputs[4292]) | (layer2_outputs[11530]);
    assign outputs[2703] = (layer2_outputs[1003]) & (layer2_outputs[9198]);
    assign outputs[2704] = ~((layer2_outputs[10605]) ^ (layer2_outputs[3810]));
    assign outputs[2705] = layer2_outputs[4663];
    assign outputs[2706] = layer2_outputs[11607];
    assign outputs[2707] = ~(layer2_outputs[2308]);
    assign outputs[2708] = (layer2_outputs[11239]) | (layer2_outputs[10190]);
    assign outputs[2709] = ~(layer2_outputs[9863]) | (layer2_outputs[604]);
    assign outputs[2710] = ~(layer2_outputs[7733]);
    assign outputs[2711] = ~(layer2_outputs[5639]);
    assign outputs[2712] = ~(layer2_outputs[2615]);
    assign outputs[2713] = ~(layer2_outputs[7182]);
    assign outputs[2714] = ~(layer2_outputs[8482]);
    assign outputs[2715] = layer2_outputs[11405];
    assign outputs[2716] = layer2_outputs[3967];
    assign outputs[2717] = ~((layer2_outputs[1756]) ^ (layer2_outputs[7549]));
    assign outputs[2718] = (layer2_outputs[3532]) | (layer2_outputs[4811]);
    assign outputs[2719] = (layer2_outputs[8118]) & ~(layer2_outputs[11488]);
    assign outputs[2720] = ~(layer2_outputs[7464]);
    assign outputs[2721] = ~((layer2_outputs[11390]) & (layer2_outputs[1994]));
    assign outputs[2722] = layer2_outputs[4616];
    assign outputs[2723] = layer2_outputs[12660];
    assign outputs[2724] = ~((layer2_outputs[6271]) ^ (layer2_outputs[3704]));
    assign outputs[2725] = layer2_outputs[7422];
    assign outputs[2726] = ~(layer2_outputs[9486]);
    assign outputs[2727] = layer2_outputs[2553];
    assign outputs[2728] = ~(layer2_outputs[1189]);
    assign outputs[2729] = ~((layer2_outputs[2380]) ^ (layer2_outputs[3325]));
    assign outputs[2730] = layer2_outputs[2043];
    assign outputs[2731] = layer2_outputs[9166];
    assign outputs[2732] = layer2_outputs[12099];
    assign outputs[2733] = ~(layer2_outputs[12206]);
    assign outputs[2734] = ~(layer2_outputs[3065]);
    assign outputs[2735] = (layer2_outputs[6086]) ^ (layer2_outputs[12242]);
    assign outputs[2736] = ~(layer2_outputs[889]);
    assign outputs[2737] = ~(layer2_outputs[6943]);
    assign outputs[2738] = ~((layer2_outputs[2408]) | (layer2_outputs[3678]));
    assign outputs[2739] = (layer2_outputs[3844]) & (layer2_outputs[8113]);
    assign outputs[2740] = layer2_outputs[12398];
    assign outputs[2741] = (layer2_outputs[476]) ^ (layer2_outputs[10599]);
    assign outputs[2742] = ~(layer2_outputs[6538]);
    assign outputs[2743] = layer2_outputs[1964];
    assign outputs[2744] = ~((layer2_outputs[8938]) ^ (layer2_outputs[11858]));
    assign outputs[2745] = (layer2_outputs[5325]) ^ (layer2_outputs[10529]);
    assign outputs[2746] = layer2_outputs[3550];
    assign outputs[2747] = ~(layer2_outputs[4831]);
    assign outputs[2748] = ~((layer2_outputs[3971]) | (layer2_outputs[874]));
    assign outputs[2749] = layer2_outputs[7704];
    assign outputs[2750] = ~((layer2_outputs[12157]) & (layer2_outputs[23]));
    assign outputs[2751] = ~((layer2_outputs[11965]) ^ (layer2_outputs[8930]));
    assign outputs[2752] = layer2_outputs[5428];
    assign outputs[2753] = ~((layer2_outputs[6865]) ^ (layer2_outputs[5403]));
    assign outputs[2754] = layer2_outputs[3744];
    assign outputs[2755] = ~(layer2_outputs[381]);
    assign outputs[2756] = ~(layer2_outputs[4276]);
    assign outputs[2757] = ~(layer2_outputs[7469]);
    assign outputs[2758] = (layer2_outputs[12077]) & (layer2_outputs[6797]);
    assign outputs[2759] = (layer2_outputs[3011]) | (layer2_outputs[1829]);
    assign outputs[2760] = layer2_outputs[4005];
    assign outputs[2761] = layer2_outputs[7188];
    assign outputs[2762] = ~(layer2_outputs[12520]) | (layer2_outputs[11633]);
    assign outputs[2763] = (layer2_outputs[11765]) & ~(layer2_outputs[4574]);
    assign outputs[2764] = layer2_outputs[1638];
    assign outputs[2765] = layer2_outputs[5766];
    assign outputs[2766] = ~((layer2_outputs[5036]) ^ (layer2_outputs[12404]));
    assign outputs[2767] = ~((layer2_outputs[8867]) & (layer2_outputs[10132]));
    assign outputs[2768] = (layer2_outputs[9808]) & ~(layer2_outputs[1303]);
    assign outputs[2769] = ~(layer2_outputs[2906]) | (layer2_outputs[3559]);
    assign outputs[2770] = ~((layer2_outputs[175]) | (layer2_outputs[8829]));
    assign outputs[2771] = ~(layer2_outputs[3225]);
    assign outputs[2772] = (layer2_outputs[4404]) & ~(layer2_outputs[6154]);
    assign outputs[2773] = ~(layer2_outputs[6551]);
    assign outputs[2774] = ~((layer2_outputs[4657]) ^ (layer2_outputs[10837]));
    assign outputs[2775] = ~(layer2_outputs[5510]) | (layer2_outputs[4187]);
    assign outputs[2776] = (layer2_outputs[6574]) & ~(layer2_outputs[10156]);
    assign outputs[2777] = ~(layer2_outputs[4495]);
    assign outputs[2778] = ~(layer2_outputs[1244]);
    assign outputs[2779] = (layer2_outputs[1155]) ^ (layer2_outputs[9764]);
    assign outputs[2780] = ~(layer2_outputs[8703]) | (layer2_outputs[9211]);
    assign outputs[2781] = ~((layer2_outputs[5492]) ^ (layer2_outputs[62]));
    assign outputs[2782] = ~((layer2_outputs[3169]) ^ (layer2_outputs[3446]));
    assign outputs[2783] = ~((layer2_outputs[10376]) ^ (layer2_outputs[2958]));
    assign outputs[2784] = ~(layer2_outputs[5661]);
    assign outputs[2785] = ~(layer2_outputs[8918]) | (layer2_outputs[6531]);
    assign outputs[2786] = ~(layer2_outputs[5374]);
    assign outputs[2787] = (layer2_outputs[5808]) ^ (layer2_outputs[9811]);
    assign outputs[2788] = layer2_outputs[5393];
    assign outputs[2789] = layer2_outputs[8500];
    assign outputs[2790] = layer2_outputs[7955];
    assign outputs[2791] = (layer2_outputs[5041]) & (layer2_outputs[7738]);
    assign outputs[2792] = (layer2_outputs[7547]) | (layer2_outputs[4786]);
    assign outputs[2793] = ~(layer2_outputs[7678]);
    assign outputs[2794] = layer2_outputs[3306];
    assign outputs[2795] = ~((layer2_outputs[4482]) ^ (layer2_outputs[9732]));
    assign outputs[2796] = layer2_outputs[380];
    assign outputs[2797] = layer2_outputs[6287];
    assign outputs[2798] = layer2_outputs[1470];
    assign outputs[2799] = layer2_outputs[9590];
    assign outputs[2800] = layer2_outputs[5714];
    assign outputs[2801] = ~(layer2_outputs[6498]);
    assign outputs[2802] = (layer2_outputs[8302]) & ~(layer2_outputs[2376]);
    assign outputs[2803] = layer2_outputs[9592];
    assign outputs[2804] = ~(layer2_outputs[4561]);
    assign outputs[2805] = (layer2_outputs[1364]) ^ (layer2_outputs[3249]);
    assign outputs[2806] = ~(layer2_outputs[10944]) | (layer2_outputs[6290]);
    assign outputs[2807] = layer2_outputs[8032];
    assign outputs[2808] = ~(layer2_outputs[12057]);
    assign outputs[2809] = (layer2_outputs[2635]) & (layer2_outputs[11585]);
    assign outputs[2810] = ~(layer2_outputs[5069]);
    assign outputs[2811] = ~((layer2_outputs[197]) ^ (layer2_outputs[9746]));
    assign outputs[2812] = ~(layer2_outputs[2688]);
    assign outputs[2813] = ~(layer2_outputs[6042]) | (layer2_outputs[8725]);
    assign outputs[2814] = (layer2_outputs[8332]) ^ (layer2_outputs[7312]);
    assign outputs[2815] = layer2_outputs[7823];
    assign outputs[2816] = ~(layer2_outputs[230]);
    assign outputs[2817] = ~(layer2_outputs[759]) | (layer2_outputs[6027]);
    assign outputs[2818] = ~((layer2_outputs[1375]) ^ (layer2_outputs[2723]));
    assign outputs[2819] = (layer2_outputs[10204]) | (layer2_outputs[6826]);
    assign outputs[2820] = (layer2_outputs[7890]) ^ (layer2_outputs[11930]);
    assign outputs[2821] = (layer2_outputs[11146]) & ~(layer2_outputs[8238]);
    assign outputs[2822] = layer2_outputs[4394];
    assign outputs[2823] = (layer2_outputs[5579]) ^ (layer2_outputs[2841]);
    assign outputs[2824] = (layer2_outputs[9251]) | (layer2_outputs[11738]);
    assign outputs[2825] = layer2_outputs[3178];
    assign outputs[2826] = ~(layer2_outputs[9766]);
    assign outputs[2827] = ~((layer2_outputs[11395]) & (layer2_outputs[5676]));
    assign outputs[2828] = (layer2_outputs[12631]) & ~(layer2_outputs[9399]);
    assign outputs[2829] = ~((layer2_outputs[12079]) & (layer2_outputs[8160]));
    assign outputs[2830] = ~(layer2_outputs[2637]);
    assign outputs[2831] = ~(layer2_outputs[2280]);
    assign outputs[2832] = ~((layer2_outputs[6452]) ^ (layer2_outputs[1624]));
    assign outputs[2833] = ~(layer2_outputs[12491]);
    assign outputs[2834] = ~(layer2_outputs[5200]);
    assign outputs[2835] = ~(layer2_outputs[9341]);
    assign outputs[2836] = (layer2_outputs[3969]) ^ (layer2_outputs[3417]);
    assign outputs[2837] = ~(layer2_outputs[7531]) | (layer2_outputs[3976]);
    assign outputs[2838] = (layer2_outputs[1774]) | (layer2_outputs[5690]);
    assign outputs[2839] = (layer2_outputs[861]) | (layer2_outputs[6619]);
    assign outputs[2840] = layer2_outputs[6849];
    assign outputs[2841] = ~((layer2_outputs[320]) ^ (layer2_outputs[4378]));
    assign outputs[2842] = ~(layer2_outputs[3602]);
    assign outputs[2843] = ~(layer2_outputs[6352]);
    assign outputs[2844] = ~(layer2_outputs[833]);
    assign outputs[2845] = ~(layer2_outputs[5868]);
    assign outputs[2846] = layer2_outputs[11739];
    assign outputs[2847] = ~(layer2_outputs[3048]) | (layer2_outputs[9768]);
    assign outputs[2848] = ~(layer2_outputs[1285]);
    assign outputs[2849] = layer2_outputs[1547];
    assign outputs[2850] = ~(layer2_outputs[1466]);
    assign outputs[2851] = (layer2_outputs[12306]) ^ (layer2_outputs[3620]);
    assign outputs[2852] = layer2_outputs[9566];
    assign outputs[2853] = ~(layer2_outputs[11999]);
    assign outputs[2854] = layer2_outputs[7863];
    assign outputs[2855] = ~((layer2_outputs[7185]) ^ (layer2_outputs[9452]));
    assign outputs[2856] = layer2_outputs[9235];
    assign outputs[2857] = layer2_outputs[320];
    assign outputs[2858] = (layer2_outputs[4000]) & (layer2_outputs[4052]);
    assign outputs[2859] = ~((layer2_outputs[5302]) ^ (layer2_outputs[11294]));
    assign outputs[2860] = ~((layer2_outputs[7158]) ^ (layer2_outputs[8846]));
    assign outputs[2861] = ~((layer2_outputs[10757]) ^ (layer2_outputs[3614]));
    assign outputs[2862] = ~((layer2_outputs[5972]) ^ (layer2_outputs[12571]));
    assign outputs[2863] = layer2_outputs[5859];
    assign outputs[2864] = ~((layer2_outputs[6149]) ^ (layer2_outputs[10230]));
    assign outputs[2865] = ~(layer2_outputs[6318]);
    assign outputs[2866] = ~(layer2_outputs[854]);
    assign outputs[2867] = ~((layer2_outputs[1386]) ^ (layer2_outputs[8265]));
    assign outputs[2868] = layer2_outputs[9122];
    assign outputs[2869] = ~((layer2_outputs[11698]) ^ (layer2_outputs[8033]));
    assign outputs[2870] = (layer2_outputs[8234]) & ~(layer2_outputs[9094]);
    assign outputs[2871] = layer2_outputs[8024];
    assign outputs[2872] = (layer2_outputs[3587]) & ~(layer2_outputs[10021]);
    assign outputs[2873] = layer2_outputs[1294];
    assign outputs[2874] = (layer2_outputs[9773]) ^ (layer2_outputs[11910]);
    assign outputs[2875] = ~(layer2_outputs[2659]);
    assign outputs[2876] = ~(layer2_outputs[6003]);
    assign outputs[2877] = ~(layer2_outputs[12575]) | (layer2_outputs[794]);
    assign outputs[2878] = ~((layer2_outputs[10973]) & (layer2_outputs[7148]));
    assign outputs[2879] = layer2_outputs[11711];
    assign outputs[2880] = layer2_outputs[3294];
    assign outputs[2881] = layer2_outputs[9448];
    assign outputs[2882] = (layer2_outputs[4356]) | (layer2_outputs[4616]);
    assign outputs[2883] = layer2_outputs[4869];
    assign outputs[2884] = layer2_outputs[11823];
    assign outputs[2885] = layer2_outputs[12087];
    assign outputs[2886] = (layer2_outputs[7583]) ^ (layer2_outputs[4921]);
    assign outputs[2887] = ~((layer2_outputs[3421]) ^ (layer2_outputs[4998]));
    assign outputs[2888] = ~((layer2_outputs[2725]) ^ (layer2_outputs[6528]));
    assign outputs[2889] = ~(layer2_outputs[1330]);
    assign outputs[2890] = ~((layer2_outputs[896]) & (layer2_outputs[8273]));
    assign outputs[2891] = ~(layer2_outputs[12293]);
    assign outputs[2892] = ~(layer2_outputs[9930]) | (layer2_outputs[480]);
    assign outputs[2893] = layer2_outputs[1687];
    assign outputs[2894] = layer2_outputs[11208];
    assign outputs[2895] = ~((layer2_outputs[10952]) & (layer2_outputs[10360]));
    assign outputs[2896] = (layer2_outputs[7314]) & ~(layer2_outputs[6320]);
    assign outputs[2897] = (layer2_outputs[9536]) & ~(layer2_outputs[1265]);
    assign outputs[2898] = (layer2_outputs[11154]) ^ (layer2_outputs[1607]);
    assign outputs[2899] = layer2_outputs[3396];
    assign outputs[2900] = ~(layer2_outputs[2951]);
    assign outputs[2901] = (layer2_outputs[9269]) ^ (layer2_outputs[12562]);
    assign outputs[2902] = ~(layer2_outputs[7858]);
    assign outputs[2903] = layer2_outputs[610];
    assign outputs[2904] = layer2_outputs[4059];
    assign outputs[2905] = ~((layer2_outputs[1673]) ^ (layer2_outputs[2128]));
    assign outputs[2906] = ~(layer2_outputs[10335]);
    assign outputs[2907] = ~(layer2_outputs[3857]);
    assign outputs[2908] = (layer2_outputs[1082]) ^ (layer2_outputs[10027]);
    assign outputs[2909] = (layer2_outputs[8185]) ^ (layer2_outputs[11431]);
    assign outputs[2910] = (layer2_outputs[8905]) ^ (layer2_outputs[4918]);
    assign outputs[2911] = ~((layer2_outputs[9835]) ^ (layer2_outputs[11374]));
    assign outputs[2912] = ~((layer2_outputs[9746]) | (layer2_outputs[4199]));
    assign outputs[2913] = ~(layer2_outputs[10426]) | (layer2_outputs[7842]);
    assign outputs[2914] = ~(layer2_outputs[3689]);
    assign outputs[2915] = layer2_outputs[10683];
    assign outputs[2916] = ~(layer2_outputs[8508]);
    assign outputs[2917] = (layer2_outputs[8070]) & ~(layer2_outputs[11497]);
    assign outputs[2918] = ~(layer2_outputs[1838]);
    assign outputs[2919] = (layer2_outputs[3681]) ^ (layer2_outputs[3877]);
    assign outputs[2920] = layer2_outputs[4585];
    assign outputs[2921] = layer2_outputs[9325];
    assign outputs[2922] = layer2_outputs[8012];
    assign outputs[2923] = (layer2_outputs[5455]) ^ (layer2_outputs[3788]);
    assign outputs[2924] = layer2_outputs[6900];
    assign outputs[2925] = ~((layer2_outputs[2979]) ^ (layer2_outputs[7571]));
    assign outputs[2926] = layer2_outputs[11042];
    assign outputs[2927] = ~(layer2_outputs[12544]);
    assign outputs[2928] = ~((layer2_outputs[3846]) ^ (layer2_outputs[8331]));
    assign outputs[2929] = ~((layer2_outputs[6454]) | (layer2_outputs[9278]));
    assign outputs[2930] = layer2_outputs[6278];
    assign outputs[2931] = ~((layer2_outputs[4650]) ^ (layer2_outputs[2215]));
    assign outputs[2932] = ~(layer2_outputs[12655]);
    assign outputs[2933] = ~(layer2_outputs[6966]);
    assign outputs[2934] = layer2_outputs[1758];
    assign outputs[2935] = ~(layer2_outputs[8927]);
    assign outputs[2936] = ~(layer2_outputs[912]);
    assign outputs[2937] = (layer2_outputs[1747]) & ~(layer2_outputs[11285]);
    assign outputs[2938] = (layer2_outputs[9219]) ^ (layer2_outputs[5628]);
    assign outputs[2939] = layer2_outputs[10984];
    assign outputs[2940] = layer2_outputs[6189];
    assign outputs[2941] = ~((layer2_outputs[10118]) ^ (layer2_outputs[6796]));
    assign outputs[2942] = ~(layer2_outputs[1418]);
    assign outputs[2943] = ~(layer2_outputs[9022]);
    assign outputs[2944] = layer2_outputs[1044];
    assign outputs[2945] = ~(layer2_outputs[4665]);
    assign outputs[2946] = layer2_outputs[1694];
    assign outputs[2947] = ~((layer2_outputs[11884]) ^ (layer2_outputs[2019]));
    assign outputs[2948] = layer2_outputs[1735];
    assign outputs[2949] = ~(layer2_outputs[11107]);
    assign outputs[2950] = ~(layer2_outputs[1209]);
    assign outputs[2951] = ~(layer2_outputs[12580]);
    assign outputs[2952] = ~(layer2_outputs[8351]);
    assign outputs[2953] = ~(layer2_outputs[10348]);
    assign outputs[2954] = ~(layer2_outputs[3439]);
    assign outputs[2955] = layer2_outputs[6999];
    assign outputs[2956] = ~(layer2_outputs[12037]);
    assign outputs[2957] = layer2_outputs[2633];
    assign outputs[2958] = ~(layer2_outputs[11992]);
    assign outputs[2959] = ~(layer2_outputs[10821]);
    assign outputs[2960] = layer2_outputs[909];
    assign outputs[2961] = (layer2_outputs[8401]) ^ (layer2_outputs[1357]);
    assign outputs[2962] = ~((layer2_outputs[8771]) ^ (layer2_outputs[316]));
    assign outputs[2963] = layer2_outputs[6341];
    assign outputs[2964] = layer2_outputs[10776];
    assign outputs[2965] = layer2_outputs[513];
    assign outputs[2966] = layer2_outputs[7537];
    assign outputs[2967] = ~(layer2_outputs[2351]);
    assign outputs[2968] = (layer2_outputs[2676]) & (layer2_outputs[7938]);
    assign outputs[2969] = (layer2_outputs[240]) ^ (layer2_outputs[6718]);
    assign outputs[2970] = layer2_outputs[11348];
    assign outputs[2971] = layer2_outputs[7422];
    assign outputs[2972] = ~(layer2_outputs[588]);
    assign outputs[2973] = ~(layer2_outputs[1726]);
    assign outputs[2974] = ~((layer2_outputs[10484]) ^ (layer2_outputs[9442]));
    assign outputs[2975] = (layer2_outputs[8968]) ^ (layer2_outputs[9771]);
    assign outputs[2976] = ~(layer2_outputs[4521]);
    assign outputs[2977] = ~(layer2_outputs[7971]);
    assign outputs[2978] = ~(layer2_outputs[7876]);
    assign outputs[2979] = ~((layer2_outputs[10472]) ^ (layer2_outputs[9964]));
    assign outputs[2980] = ~(layer2_outputs[7466]);
    assign outputs[2981] = ~(layer2_outputs[11872]);
    assign outputs[2982] = ~(layer2_outputs[4750]);
    assign outputs[2983] = ~(layer2_outputs[12770]);
    assign outputs[2984] = ~(layer2_outputs[2357]);
    assign outputs[2985] = ~(layer2_outputs[11127]);
    assign outputs[2986] = layer2_outputs[1510];
    assign outputs[2987] = layer2_outputs[939];
    assign outputs[2988] = layer2_outputs[11334];
    assign outputs[2989] = ~(layer2_outputs[3986]);
    assign outputs[2990] = layer2_outputs[10256];
    assign outputs[2991] = layer2_outputs[3519];
    assign outputs[2992] = layer2_outputs[4269];
    assign outputs[2993] = ~((layer2_outputs[3643]) ^ (layer2_outputs[1134]));
    assign outputs[2994] = layer2_outputs[12382];
    assign outputs[2995] = ~(layer2_outputs[10397]) | (layer2_outputs[4548]);
    assign outputs[2996] = ~((layer2_outputs[11054]) ^ (layer2_outputs[6105]));
    assign outputs[2997] = ~(layer2_outputs[8835]);
    assign outputs[2998] = (layer2_outputs[5970]) ^ (layer2_outputs[1056]);
    assign outputs[2999] = ~(layer2_outputs[9928]);
    assign outputs[3000] = layer2_outputs[3906];
    assign outputs[3001] = ~((layer2_outputs[8049]) ^ (layer2_outputs[7675]));
    assign outputs[3002] = ~((layer2_outputs[9814]) & (layer2_outputs[1280]));
    assign outputs[3003] = ~(layer2_outputs[3426]);
    assign outputs[3004] = (layer2_outputs[8903]) & ~(layer2_outputs[5369]);
    assign outputs[3005] = ~(layer2_outputs[1112]);
    assign outputs[3006] = ~(layer2_outputs[11508]);
    assign outputs[3007] = ~((layer2_outputs[33]) ^ (layer2_outputs[1801]));
    assign outputs[3008] = (layer2_outputs[816]) ^ (layer2_outputs[10924]);
    assign outputs[3009] = (layer2_outputs[8335]) & ~(layer2_outputs[1304]);
    assign outputs[3010] = layer2_outputs[4959];
    assign outputs[3011] = ~(layer2_outputs[3776]);
    assign outputs[3012] = ~(layer2_outputs[1466]);
    assign outputs[3013] = ~(layer2_outputs[12138]);
    assign outputs[3014] = ~(layer2_outputs[9981]);
    assign outputs[3015] = ~(layer2_outputs[11884]);
    assign outputs[3016] = (layer2_outputs[10875]) ^ (layer2_outputs[4350]);
    assign outputs[3017] = (layer2_outputs[362]) | (layer2_outputs[6451]);
    assign outputs[3018] = layer2_outputs[8445];
    assign outputs[3019] = layer2_outputs[1662];
    assign outputs[3020] = ~(layer2_outputs[8227]);
    assign outputs[3021] = ~((layer2_outputs[637]) ^ (layer2_outputs[7263]));
    assign outputs[3022] = (layer2_outputs[11395]) ^ (layer2_outputs[1432]);
    assign outputs[3023] = layer2_outputs[11302];
    assign outputs[3024] = (layer2_outputs[12297]) | (layer2_outputs[12733]);
    assign outputs[3025] = (layer2_outputs[10322]) ^ (layer2_outputs[4295]);
    assign outputs[3026] = layer2_outputs[5208];
    assign outputs[3027] = ~(layer2_outputs[1490]);
    assign outputs[3028] = ~(layer2_outputs[5807]);
    assign outputs[3029] = ~(layer2_outputs[10358]) | (layer2_outputs[6895]);
    assign outputs[3030] = layer2_outputs[3720];
    assign outputs[3031] = layer2_outputs[11648];
    assign outputs[3032] = (layer2_outputs[7236]) & ~(layer2_outputs[2827]);
    assign outputs[3033] = ~(layer2_outputs[10165]) | (layer2_outputs[6094]);
    assign outputs[3034] = ~(layer2_outputs[9450]) | (layer2_outputs[4537]);
    assign outputs[3035] = layer2_outputs[11090];
    assign outputs[3036] = ~((layer2_outputs[5452]) ^ (layer2_outputs[5219]));
    assign outputs[3037] = layer2_outputs[5508];
    assign outputs[3038] = ~(layer2_outputs[5604]);
    assign outputs[3039] = layer2_outputs[8377];
    assign outputs[3040] = ~(layer2_outputs[4420]);
    assign outputs[3041] = ~(layer2_outputs[10489]);
    assign outputs[3042] = (layer2_outputs[7378]) & ~(layer2_outputs[11267]);
    assign outputs[3043] = ~(layer2_outputs[8416]) | (layer2_outputs[6680]);
    assign outputs[3044] = layer2_outputs[12664];
    assign outputs[3045] = (layer2_outputs[5790]) & (layer2_outputs[5914]);
    assign outputs[3046] = layer2_outputs[9494];
    assign outputs[3047] = layer2_outputs[8172];
    assign outputs[3048] = layer2_outputs[11818];
    assign outputs[3049] = layer2_outputs[7514];
    assign outputs[3050] = ~(layer2_outputs[8484]);
    assign outputs[3051] = ~(layer2_outputs[10821]);
    assign outputs[3052] = ~(layer2_outputs[11109]);
    assign outputs[3053] = layer2_outputs[4049];
    assign outputs[3054] = ~(layer2_outputs[10923]);
    assign outputs[3055] = ~(layer2_outputs[9761]);
    assign outputs[3056] = (layer2_outputs[3640]) & ~(layer2_outputs[11394]);
    assign outputs[3057] = layer2_outputs[10977];
    assign outputs[3058] = ~((layer2_outputs[9148]) ^ (layer2_outputs[12299]));
    assign outputs[3059] = (layer2_outputs[11367]) ^ (layer2_outputs[1096]);
    assign outputs[3060] = ~(layer2_outputs[7459]);
    assign outputs[3061] = layer2_outputs[703];
    assign outputs[3062] = (layer2_outputs[2902]) ^ (layer2_outputs[1367]);
    assign outputs[3063] = ~((layer2_outputs[4456]) ^ (layer2_outputs[10398]));
    assign outputs[3064] = (layer2_outputs[378]) ^ (layer2_outputs[8002]);
    assign outputs[3065] = layer2_outputs[457];
    assign outputs[3066] = ~(layer2_outputs[10600]);
    assign outputs[3067] = ~((layer2_outputs[12296]) ^ (layer2_outputs[9080]));
    assign outputs[3068] = (layer2_outputs[4431]) & (layer2_outputs[9808]);
    assign outputs[3069] = (layer2_outputs[9035]) | (layer2_outputs[7632]);
    assign outputs[3070] = ~(layer2_outputs[11521]);
    assign outputs[3071] = layer2_outputs[5812];
    assign outputs[3072] = layer2_outputs[337];
    assign outputs[3073] = layer2_outputs[10317];
    assign outputs[3074] = ~(layer2_outputs[8957]);
    assign outputs[3075] = (layer2_outputs[2322]) & ~(layer2_outputs[8927]);
    assign outputs[3076] = (layer2_outputs[3319]) | (layer2_outputs[6239]);
    assign outputs[3077] = ~(layer2_outputs[6269]);
    assign outputs[3078] = layer2_outputs[7388];
    assign outputs[3079] = (layer2_outputs[2693]) ^ (layer2_outputs[5065]);
    assign outputs[3080] = ~(layer2_outputs[3833]);
    assign outputs[3081] = layer2_outputs[9977];
    assign outputs[3082] = ~(layer2_outputs[5811]) | (layer2_outputs[4002]);
    assign outputs[3083] = layer2_outputs[11370];
    assign outputs[3084] = (layer2_outputs[8868]) ^ (layer2_outputs[4725]);
    assign outputs[3085] = (layer2_outputs[5786]) ^ (layer2_outputs[7705]);
    assign outputs[3086] = (layer2_outputs[5325]) | (layer2_outputs[7962]);
    assign outputs[3087] = layer2_outputs[3119];
    assign outputs[3088] = ~(layer2_outputs[6002]);
    assign outputs[3089] = ~(layer2_outputs[8000]);
    assign outputs[3090] = layer2_outputs[5364];
    assign outputs[3091] = ~(layer2_outputs[3094]);
    assign outputs[3092] = ~(layer2_outputs[6696]);
    assign outputs[3093] = ~((layer2_outputs[3159]) & (layer2_outputs[1334]));
    assign outputs[3094] = layer2_outputs[3949];
    assign outputs[3095] = (layer2_outputs[2779]) & (layer2_outputs[3995]);
    assign outputs[3096] = ~(layer2_outputs[10859]);
    assign outputs[3097] = ~(layer2_outputs[8542]);
    assign outputs[3098] = ~(layer2_outputs[3354]);
    assign outputs[3099] = layer2_outputs[2552];
    assign outputs[3100] = ~(layer2_outputs[3040]);
    assign outputs[3101] = (layer2_outputs[7575]) | (layer2_outputs[968]);
    assign outputs[3102] = ~(layer2_outputs[11662]);
    assign outputs[3103] = ~(layer2_outputs[6709]);
    assign outputs[3104] = (layer2_outputs[9762]) | (layer2_outputs[6968]);
    assign outputs[3105] = (layer2_outputs[7635]) | (layer2_outputs[6741]);
    assign outputs[3106] = (layer2_outputs[11602]) & ~(layer2_outputs[1797]);
    assign outputs[3107] = ~(layer2_outputs[7371]);
    assign outputs[3108] = ~(layer2_outputs[3118]) | (layer2_outputs[3947]);
    assign outputs[3109] = ~((layer2_outputs[6803]) ^ (layer2_outputs[5897]));
    assign outputs[3110] = layer2_outputs[1882];
    assign outputs[3111] = ~(layer2_outputs[1377]);
    assign outputs[3112] = (layer2_outputs[2708]) ^ (layer2_outputs[11439]);
    assign outputs[3113] = ~((layer2_outputs[990]) ^ (layer2_outputs[6187]));
    assign outputs[3114] = (layer2_outputs[2016]) | (layer2_outputs[5029]);
    assign outputs[3115] = (layer2_outputs[2121]) ^ (layer2_outputs[2710]);
    assign outputs[3116] = (layer2_outputs[8604]) & ~(layer2_outputs[11949]);
    assign outputs[3117] = layer2_outputs[5571];
    assign outputs[3118] = ~(layer2_outputs[11554]);
    assign outputs[3119] = (layer2_outputs[1412]) & ~(layer2_outputs[1518]);
    assign outputs[3120] = layer2_outputs[8789];
    assign outputs[3121] = layer2_outputs[12144];
    assign outputs[3122] = ~(layer2_outputs[11787]);
    assign outputs[3123] = ~(layer2_outputs[9807]);
    assign outputs[3124] = ~(layer2_outputs[8350]);
    assign outputs[3125] = ~(layer2_outputs[9169]);
    assign outputs[3126] = ~((layer2_outputs[5232]) | (layer2_outputs[9381]));
    assign outputs[3127] = ~(layer2_outputs[4223]);
    assign outputs[3128] = ~(layer2_outputs[5102]) | (layer2_outputs[1701]);
    assign outputs[3129] = (layer2_outputs[5221]) ^ (layer2_outputs[5800]);
    assign outputs[3130] = (layer2_outputs[582]) ^ (layer2_outputs[6470]);
    assign outputs[3131] = ~((layer2_outputs[4122]) & (layer2_outputs[2600]));
    assign outputs[3132] = layer2_outputs[3955];
    assign outputs[3133] = layer2_outputs[1856];
    assign outputs[3134] = layer2_outputs[5844];
    assign outputs[3135] = ~(layer2_outputs[5494]) | (layer2_outputs[10732]);
    assign outputs[3136] = layer2_outputs[1655];
    assign outputs[3137] = ~((layer2_outputs[11821]) | (layer2_outputs[7089]));
    assign outputs[3138] = layer2_outputs[2217];
    assign outputs[3139] = layer2_outputs[11888];
    assign outputs[3140] = ~(layer2_outputs[4929]);
    assign outputs[3141] = layer2_outputs[4797];
    assign outputs[3142] = ~(layer2_outputs[8949]);
    assign outputs[3143] = ~(layer2_outputs[2892]);
    assign outputs[3144] = ~(layer2_outputs[11421]) | (layer2_outputs[10317]);
    assign outputs[3145] = ~(layer2_outputs[962]);
    assign outputs[3146] = ~(layer2_outputs[9832]);
    assign outputs[3147] = ~((layer2_outputs[646]) ^ (layer2_outputs[7611]));
    assign outputs[3148] = layer2_outputs[12310];
    assign outputs[3149] = layer2_outputs[1459];
    assign outputs[3150] = ~(layer2_outputs[3520]);
    assign outputs[3151] = layer2_outputs[9523];
    assign outputs[3152] = (layer2_outputs[2362]) & ~(layer2_outputs[5793]);
    assign outputs[3153] = ~(layer2_outputs[1106]);
    assign outputs[3154] = ~(layer2_outputs[9993]);
    assign outputs[3155] = layer2_outputs[2022];
    assign outputs[3156] = (layer2_outputs[3411]) ^ (layer2_outputs[12136]);
    assign outputs[3157] = layer2_outputs[3549];
    assign outputs[3158] = layer2_outputs[9989];
    assign outputs[3159] = ~((layer2_outputs[2628]) & (layer2_outputs[8598]));
    assign outputs[3160] = ~((layer2_outputs[1341]) ^ (layer2_outputs[8580]));
    assign outputs[3161] = layer2_outputs[5452];
    assign outputs[3162] = layer2_outputs[909];
    assign outputs[3163] = layer2_outputs[7585];
    assign outputs[3164] = (layer2_outputs[11473]) & (layer2_outputs[1429]);
    assign outputs[3165] = (layer2_outputs[5672]) & ~(layer2_outputs[12039]);
    assign outputs[3166] = layer2_outputs[10768];
    assign outputs[3167] = ~(layer2_outputs[4780]);
    assign outputs[3168] = layer2_outputs[5654];
    assign outputs[3169] = ~((layer2_outputs[8328]) ^ (layer2_outputs[11714]));
    assign outputs[3170] = (layer2_outputs[1330]) ^ (layer2_outputs[7934]);
    assign outputs[3171] = ~(layer2_outputs[29]) | (layer2_outputs[9787]);
    assign outputs[3172] = (layer2_outputs[2956]) ^ (layer2_outputs[6801]);
    assign outputs[3173] = ~((layer2_outputs[802]) & (layer2_outputs[7215]));
    assign outputs[3174] = ~(layer2_outputs[4235]);
    assign outputs[3175] = layer2_outputs[5253];
    assign outputs[3176] = (layer2_outputs[8139]) ^ (layer2_outputs[10042]);
    assign outputs[3177] = ~((layer2_outputs[11003]) | (layer2_outputs[370]));
    assign outputs[3178] = ~((layer2_outputs[3960]) ^ (layer2_outputs[12708]));
    assign outputs[3179] = ~(layer2_outputs[10066]);
    assign outputs[3180] = ~((layer2_outputs[9930]) & (layer2_outputs[12263]));
    assign outputs[3181] = ~((layer2_outputs[1526]) ^ (layer2_outputs[11917]));
    assign outputs[3182] = layer2_outputs[2472];
    assign outputs[3183] = layer2_outputs[7375];
    assign outputs[3184] = ~(layer2_outputs[9241]);
    assign outputs[3185] = layer2_outputs[694];
    assign outputs[3186] = layer2_outputs[2299];
    assign outputs[3187] = ~((layer2_outputs[3427]) ^ (layer2_outputs[2434]));
    assign outputs[3188] = ~(layer2_outputs[4444]);
    assign outputs[3189] = ~(layer2_outputs[5726]) | (layer2_outputs[11475]);
    assign outputs[3190] = ~(layer2_outputs[4594]) | (layer2_outputs[355]);
    assign outputs[3191] = ~((layer2_outputs[7151]) | (layer2_outputs[4867]));
    assign outputs[3192] = layer2_outputs[720];
    assign outputs[3193] = ~(layer2_outputs[260]);
    assign outputs[3194] = ~(layer2_outputs[7872]);
    assign outputs[3195] = ~(layer2_outputs[8683]) | (layer2_outputs[3045]);
    assign outputs[3196] = ~(layer2_outputs[1313]);
    assign outputs[3197] = layer2_outputs[10175];
    assign outputs[3198] = ~(layer2_outputs[5857]);
    assign outputs[3199] = layer2_outputs[737];
    assign outputs[3200] = layer2_outputs[7261];
    assign outputs[3201] = ~(layer2_outputs[1921]);
    assign outputs[3202] = layer2_outputs[1282];
    assign outputs[3203] = ~(layer2_outputs[10146]);
    assign outputs[3204] = layer2_outputs[7882];
    assign outputs[3205] = ~(layer2_outputs[2261]);
    assign outputs[3206] = ~((layer2_outputs[10134]) & (layer2_outputs[1629]));
    assign outputs[3207] = ~(layer2_outputs[3216]);
    assign outputs[3208] = ~(layer2_outputs[5034]);
    assign outputs[3209] = layer2_outputs[2946];
    assign outputs[3210] = (layer2_outputs[8314]) ^ (layer2_outputs[11471]);
    assign outputs[3211] = (layer2_outputs[1727]) & ~(layer2_outputs[8223]);
    assign outputs[3212] = layer2_outputs[9603];
    assign outputs[3213] = ~((layer2_outputs[4194]) ^ (layer2_outputs[8144]));
    assign outputs[3214] = ~(layer2_outputs[32]);
    assign outputs[3215] = ~((layer2_outputs[2918]) ^ (layer2_outputs[1763]));
    assign outputs[3216] = ~(layer2_outputs[3568]);
    assign outputs[3217] = ~(layer2_outputs[200]);
    assign outputs[3218] = (layer2_outputs[5924]) ^ (layer2_outputs[2167]);
    assign outputs[3219] = layer2_outputs[10379];
    assign outputs[3220] = (layer2_outputs[1484]) ^ (layer2_outputs[8713]);
    assign outputs[3221] = ~(layer2_outputs[4160]) | (layer2_outputs[11396]);
    assign outputs[3222] = layer2_outputs[11713];
    assign outputs[3223] = (layer2_outputs[7865]) | (layer2_outputs[3148]);
    assign outputs[3224] = ~(layer2_outputs[2248]);
    assign outputs[3225] = ~(layer2_outputs[2443]);
    assign outputs[3226] = ~(layer2_outputs[5828]) | (layer2_outputs[10621]);
    assign outputs[3227] = ~((layer2_outputs[6208]) & (layer2_outputs[5005]));
    assign outputs[3228] = ~((layer2_outputs[6683]) ^ (layer2_outputs[8431]));
    assign outputs[3229] = layer2_outputs[11900];
    assign outputs[3230] = (layer2_outputs[12738]) & ~(layer2_outputs[1133]);
    assign outputs[3231] = ~(layer2_outputs[95]);
    assign outputs[3232] = ~(layer2_outputs[7647]);
    assign outputs[3233] = ~(layer2_outputs[4365]) | (layer2_outputs[3731]);
    assign outputs[3234] = ~(layer2_outputs[12130]);
    assign outputs[3235] = layer2_outputs[275];
    assign outputs[3236] = ~(layer2_outputs[2802]);
    assign outputs[3237] = layer2_outputs[2778];
    assign outputs[3238] = layer2_outputs[4363];
    assign outputs[3239] = layer2_outputs[7168];
    assign outputs[3240] = layer2_outputs[10693];
    assign outputs[3241] = ~(layer2_outputs[3264]) | (layer2_outputs[3522]);
    assign outputs[3242] = layer2_outputs[696];
    assign outputs[3243] = ~(layer2_outputs[2241]);
    assign outputs[3244] = ~((layer2_outputs[4900]) | (layer2_outputs[9774]));
    assign outputs[3245] = ~((layer2_outputs[3978]) ^ (layer2_outputs[9676]));
    assign outputs[3246] = layer2_outputs[6102];
    assign outputs[3247] = ~(layer2_outputs[2323]);
    assign outputs[3248] = (layer2_outputs[7183]) & ~(layer2_outputs[11682]);
    assign outputs[3249] = ~(layer2_outputs[1135]);
    assign outputs[3250] = layer2_outputs[8823];
    assign outputs[3251] = layer2_outputs[10128];
    assign outputs[3252] = ~((layer2_outputs[4402]) & (layer2_outputs[10755]));
    assign outputs[3253] = ~((layer2_outputs[9301]) & (layer2_outputs[7292]));
    assign outputs[3254] = ~((layer2_outputs[12003]) ^ (layer2_outputs[6763]));
    assign outputs[3255] = ~(layer2_outputs[2611]) | (layer2_outputs[10966]);
    assign outputs[3256] = ~(layer2_outputs[831]) | (layer2_outputs[6795]);
    assign outputs[3257] = (layer2_outputs[4962]) ^ (layer2_outputs[4108]);
    assign outputs[3258] = ~(layer2_outputs[1421]);
    assign outputs[3259] = layer2_outputs[10948];
    assign outputs[3260] = ~((layer2_outputs[11852]) | (layer2_outputs[5880]));
    assign outputs[3261] = ~((layer2_outputs[7763]) & (layer2_outputs[6630]));
    assign outputs[3262] = layer2_outputs[11848];
    assign outputs[3263] = layer2_outputs[9564];
    assign outputs[3264] = (layer2_outputs[3563]) ^ (layer2_outputs[6197]);
    assign outputs[3265] = (layer2_outputs[3707]) | (layer2_outputs[3532]);
    assign outputs[3266] = ~(layer2_outputs[7517]) | (layer2_outputs[140]);
    assign outputs[3267] = layer2_outputs[3283];
    assign outputs[3268] = ~(layer2_outputs[1438]);
    assign outputs[3269] = layer2_outputs[8399];
    assign outputs[3270] = ~(layer2_outputs[7866]);
    assign outputs[3271] = ~(layer2_outputs[6688]);
    assign outputs[3272] = layer2_outputs[4631];
    assign outputs[3273] = ~(layer2_outputs[1594]);
    assign outputs[3274] = ~(layer2_outputs[11528]);
    assign outputs[3275] = ~(layer2_outputs[8014]);
    assign outputs[3276] = ~((layer2_outputs[7487]) & (layer2_outputs[12164]));
    assign outputs[3277] = ~((layer2_outputs[11790]) | (layer2_outputs[3392]));
    assign outputs[3278] = layer2_outputs[8337];
    assign outputs[3279] = ~((layer2_outputs[8511]) ^ (layer2_outputs[8602]));
    assign outputs[3280] = ~((layer2_outputs[135]) ^ (layer2_outputs[6475]));
    assign outputs[3281] = layer2_outputs[1584];
    assign outputs[3282] = layer2_outputs[1296];
    assign outputs[3283] = layer2_outputs[6302];
    assign outputs[3284] = ~(layer2_outputs[1088]);
    assign outputs[3285] = (layer2_outputs[5313]) | (layer2_outputs[6054]);
    assign outputs[3286] = layer2_outputs[4278];
    assign outputs[3287] = ~(layer2_outputs[4227]);
    assign outputs[3288] = layer2_outputs[3538];
    assign outputs[3289] = (layer2_outputs[6098]) & (layer2_outputs[484]);
    assign outputs[3290] = layer2_outputs[5667];
    assign outputs[3291] = (layer2_outputs[9005]) ^ (layer2_outputs[6757]);
    assign outputs[3292] = layer2_outputs[484];
    assign outputs[3293] = ~(layer2_outputs[6581]) | (layer2_outputs[12054]);
    assign outputs[3294] = ~((layer2_outputs[12172]) | (layer2_outputs[856]));
    assign outputs[3295] = (layer2_outputs[5559]) ^ (layer2_outputs[9822]);
    assign outputs[3296] = ~(layer2_outputs[4596]);
    assign outputs[3297] = ~(layer2_outputs[3002]);
    assign outputs[3298] = ~(layer2_outputs[7173]);
    assign outputs[3299] = ~(layer2_outputs[6926]);
    assign outputs[3300] = layer2_outputs[2184];
    assign outputs[3301] = (layer2_outputs[1873]) & ~(layer2_outputs[3700]);
    assign outputs[3302] = ~(layer2_outputs[10200]);
    assign outputs[3303] = ~(layer2_outputs[8649]);
    assign outputs[3304] = ~(layer2_outputs[1669]);
    assign outputs[3305] = ~(layer2_outputs[1483]);
    assign outputs[3306] = (layer2_outputs[1515]) ^ (layer2_outputs[7651]);
    assign outputs[3307] = (layer2_outputs[9296]) ^ (layer2_outputs[937]);
    assign outputs[3308] = (layer2_outputs[4461]) ^ (layer2_outputs[11926]);
    assign outputs[3309] = layer2_outputs[5113];
    assign outputs[3310] = ~((layer2_outputs[4011]) & (layer2_outputs[9646]));
    assign outputs[3311] = ~((layer2_outputs[298]) ^ (layer2_outputs[12192]));
    assign outputs[3312] = layer2_outputs[8656];
    assign outputs[3313] = ~(layer2_outputs[11230]) | (layer2_outputs[9631]);
    assign outputs[3314] = ~(layer2_outputs[9914]) | (layer2_outputs[4902]);
    assign outputs[3315] = layer2_outputs[634];
    assign outputs[3316] = layer2_outputs[9128];
    assign outputs[3317] = (layer2_outputs[9207]) ^ (layer2_outputs[10930]);
    assign outputs[3318] = ~(layer2_outputs[10396]) | (layer2_outputs[2428]);
    assign outputs[3319] = ~(layer2_outputs[2854]);
    assign outputs[3320] = (layer2_outputs[4502]) & ~(layer2_outputs[4872]);
    assign outputs[3321] = ~(layer2_outputs[739]);
    assign outputs[3322] = layer2_outputs[7019];
    assign outputs[3323] = (layer2_outputs[6066]) ^ (layer2_outputs[11275]);
    assign outputs[3324] = (layer2_outputs[11356]) & ~(layer2_outputs[12487]);
    assign outputs[3325] = layer2_outputs[2817];
    assign outputs[3326] = ~(layer2_outputs[8473]);
    assign outputs[3327] = ~(layer2_outputs[11158]);
    assign outputs[3328] = layer2_outputs[1459];
    assign outputs[3329] = ~(layer2_outputs[3431]);
    assign outputs[3330] = layer2_outputs[3539];
    assign outputs[3331] = ~((layer2_outputs[487]) & (layer2_outputs[6247]));
    assign outputs[3332] = (layer2_outputs[9456]) ^ (layer2_outputs[3769]);
    assign outputs[3333] = layer2_outputs[3230];
    assign outputs[3334] = ~((layer2_outputs[1743]) ^ (layer2_outputs[3205]));
    assign outputs[3335] = ~(layer2_outputs[11745]);
    assign outputs[3336] = layer2_outputs[2150];
    assign outputs[3337] = layer2_outputs[7625];
    assign outputs[3338] = ~(layer2_outputs[6286]) | (layer2_outputs[5177]);
    assign outputs[3339] = ~(layer2_outputs[1982]);
    assign outputs[3340] = ~(layer2_outputs[5151]) | (layer2_outputs[2476]);
    assign outputs[3341] = layer2_outputs[420];
    assign outputs[3342] = ~((layer2_outputs[193]) ^ (layer2_outputs[5556]));
    assign outputs[3343] = layer2_outputs[4099];
    assign outputs[3344] = ~(layer2_outputs[8523]);
    assign outputs[3345] = ~(layer2_outputs[9897]);
    assign outputs[3346] = layer2_outputs[903];
    assign outputs[3347] = ~((layer2_outputs[4802]) | (layer2_outputs[2926]));
    assign outputs[3348] = ~((layer2_outputs[1173]) ^ (layer2_outputs[6533]));
    assign outputs[3349] = ~(layer2_outputs[10777]);
    assign outputs[3350] = (layer2_outputs[7389]) ^ (layer2_outputs[5758]);
    assign outputs[3351] = layer2_outputs[2272];
    assign outputs[3352] = (layer2_outputs[2252]) ^ (layer2_outputs[4396]);
    assign outputs[3353] = layer2_outputs[11304];
    assign outputs[3354] = ~((layer2_outputs[3979]) ^ (layer2_outputs[8654]));
    assign outputs[3355] = ~(layer2_outputs[11508]);
    assign outputs[3356] = layer2_outputs[4183];
    assign outputs[3357] = ~(layer2_outputs[7765]);
    assign outputs[3358] = ~(layer2_outputs[7006]) | (layer2_outputs[2480]);
    assign outputs[3359] = (layer2_outputs[5465]) & ~(layer2_outputs[2657]);
    assign outputs[3360] = ~((layer2_outputs[795]) & (layer2_outputs[11452]));
    assign outputs[3361] = layer2_outputs[4983];
    assign outputs[3362] = ~(layer2_outputs[11109]);
    assign outputs[3363] = layer2_outputs[6057];
    assign outputs[3364] = ~(layer2_outputs[8130]);
    assign outputs[3365] = ~(layer2_outputs[9912]) | (layer2_outputs[7136]);
    assign outputs[3366] = layer2_outputs[3876];
    assign outputs[3367] = (layer2_outputs[11056]) ^ (layer2_outputs[5322]);
    assign outputs[3368] = (layer2_outputs[1516]) & (layer2_outputs[3027]);
    assign outputs[3369] = ~(layer2_outputs[3894]);
    assign outputs[3370] = ~(layer2_outputs[6615]);
    assign outputs[3371] = layer2_outputs[7416];
    assign outputs[3372] = layer2_outputs[11901];
    assign outputs[3373] = layer2_outputs[5919];
    assign outputs[3374] = layer2_outputs[9003];
    assign outputs[3375] = layer2_outputs[3881];
    assign outputs[3376] = (layer2_outputs[5936]) ^ (layer2_outputs[445]);
    assign outputs[3377] = ~((layer2_outputs[9840]) ^ (layer2_outputs[1343]));
    assign outputs[3378] = layer2_outputs[10542];
    assign outputs[3379] = ~(layer2_outputs[310]);
    assign outputs[3380] = (layer2_outputs[4302]) ^ (layer2_outputs[3307]);
    assign outputs[3381] = ~((layer2_outputs[7267]) & (layer2_outputs[9539]));
    assign outputs[3382] = layer2_outputs[5606];
    assign outputs[3383] = ~((layer2_outputs[12634]) | (layer2_outputs[4682]));
    assign outputs[3384] = ~(layer2_outputs[2695]) | (layer2_outputs[4498]);
    assign outputs[3385] = layer2_outputs[8204];
    assign outputs[3386] = ~((layer2_outputs[6936]) ^ (layer2_outputs[2333]));
    assign outputs[3387] = (layer2_outputs[12641]) & ~(layer2_outputs[2989]);
    assign outputs[3388] = layer2_outputs[4966];
    assign outputs[3389] = ~(layer2_outputs[4539]);
    assign outputs[3390] = ~((layer2_outputs[3334]) ^ (layer2_outputs[6149]));
    assign outputs[3391] = ~(layer2_outputs[8944]) | (layer2_outputs[3745]);
    assign outputs[3392] = (layer2_outputs[4233]) ^ (layer2_outputs[9256]);
    assign outputs[3393] = (layer2_outputs[5044]) & ~(layer2_outputs[7550]);
    assign outputs[3394] = layer2_outputs[10673];
    assign outputs[3395] = layer2_outputs[12730];
    assign outputs[3396] = ~(layer2_outputs[5263]);
    assign outputs[3397] = ~(layer2_outputs[4353]) | (layer2_outputs[2986]);
    assign outputs[3398] = layer2_outputs[4483];
    assign outputs[3399] = layer2_outputs[1358];
    assign outputs[3400] = (layer2_outputs[2119]) ^ (layer2_outputs[6717]);
    assign outputs[3401] = ~(layer2_outputs[10056]);
    assign outputs[3402] = ~(layer2_outputs[2695]);
    assign outputs[3403] = ~(layer2_outputs[1054]);
    assign outputs[3404] = ~(layer2_outputs[8772]);
    assign outputs[3405] = ~(layer2_outputs[7744]);
    assign outputs[3406] = (layer2_outputs[7072]) & (layer2_outputs[9707]);
    assign outputs[3407] = layer2_outputs[9488];
    assign outputs[3408] = ~(layer2_outputs[2535]);
    assign outputs[3409] = (layer2_outputs[9707]) & ~(layer2_outputs[11444]);
    assign outputs[3410] = ~(layer2_outputs[10424]);
    assign outputs[3411] = ~(layer2_outputs[6216]);
    assign outputs[3412] = ~(layer2_outputs[1331]);
    assign outputs[3413] = ~(layer2_outputs[5008]) | (layer2_outputs[9472]);
    assign outputs[3414] = layer2_outputs[10295];
    assign outputs[3415] = ~(layer2_outputs[659]);
    assign outputs[3416] = (layer2_outputs[8681]) ^ (layer2_outputs[10136]);
    assign outputs[3417] = layer2_outputs[4338];
    assign outputs[3418] = (layer2_outputs[7051]) ^ (layer2_outputs[11709]);
    assign outputs[3419] = ~(layer2_outputs[6627]);
    assign outputs[3420] = (layer2_outputs[1546]) ^ (layer2_outputs[2937]);
    assign outputs[3421] = layer2_outputs[4454];
    assign outputs[3422] = layer2_outputs[4345];
    assign outputs[3423] = ~(layer2_outputs[7590]);
    assign outputs[3424] = layer2_outputs[4416];
    assign outputs[3425] = ~(layer2_outputs[4276]);
    assign outputs[3426] = (layer2_outputs[6451]) | (layer2_outputs[3810]);
    assign outputs[3427] = ~(layer2_outputs[5721]) | (layer2_outputs[8047]);
    assign outputs[3428] = ~((layer2_outputs[11712]) ^ (layer2_outputs[5422]));
    assign outputs[3429] = ~(layer2_outputs[7368]);
    assign outputs[3430] = (layer2_outputs[1609]) ^ (layer2_outputs[7393]);
    assign outputs[3431] = layer2_outputs[6545];
    assign outputs[3432] = layer2_outputs[7084];
    assign outputs[3433] = ~(layer2_outputs[820]);
    assign outputs[3434] = ~((layer2_outputs[11169]) & (layer2_outputs[12337]));
    assign outputs[3435] = ~(layer2_outputs[392]);
    assign outputs[3436] = ~(layer2_outputs[5407]);
    assign outputs[3437] = ~((layer2_outputs[11245]) ^ (layer2_outputs[7434]));
    assign outputs[3438] = (layer2_outputs[3674]) ^ (layer2_outputs[8014]);
    assign outputs[3439] = (layer2_outputs[130]) ^ (layer2_outputs[9756]);
    assign outputs[3440] = ~(layer2_outputs[8145]);
    assign outputs[3441] = layer2_outputs[11234];
    assign outputs[3442] = layer2_outputs[10731];
    assign outputs[3443] = ~(layer2_outputs[6409]);
    assign outputs[3444] = ~(layer2_outputs[1717]);
    assign outputs[3445] = ~(layer2_outputs[5306]) | (layer2_outputs[12381]);
    assign outputs[3446] = layer2_outputs[1419];
    assign outputs[3447] = (layer2_outputs[2691]) ^ (layer2_outputs[7915]);
    assign outputs[3448] = ~(layer2_outputs[10515]) | (layer2_outputs[12712]);
    assign outputs[3449] = (layer2_outputs[5501]) | (layer2_outputs[3792]);
    assign outputs[3450] = ~(layer2_outputs[10159]);
    assign outputs[3451] = ~(layer2_outputs[11479]);
    assign outputs[3452] = ~(layer2_outputs[7301]);
    assign outputs[3453] = (layer2_outputs[2842]) ^ (layer2_outputs[6610]);
    assign outputs[3454] = layer2_outputs[9224];
    assign outputs[3455] = ~(layer2_outputs[8412]);
    assign outputs[3456] = (layer2_outputs[11565]) ^ (layer2_outputs[7552]);
    assign outputs[3457] = layer2_outputs[8612];
    assign outputs[3458] = layer2_outputs[6942];
    assign outputs[3459] = ~(layer2_outputs[3569]);
    assign outputs[3460] = ~((layer2_outputs[11459]) ^ (layer2_outputs[6314]));
    assign outputs[3461] = ~(layer2_outputs[11761]);
    assign outputs[3462] = (layer2_outputs[11368]) ^ (layer2_outputs[8139]);
    assign outputs[3463] = layer2_outputs[6273];
    assign outputs[3464] = (layer2_outputs[8166]) & ~(layer2_outputs[8637]);
    assign outputs[3465] = layer2_outputs[2580];
    assign outputs[3466] = ~(layer2_outputs[63]);
    assign outputs[3467] = layer2_outputs[4806];
    assign outputs[3468] = ~((layer2_outputs[10680]) | (layer2_outputs[860]));
    assign outputs[3469] = layer2_outputs[5035];
    assign outputs[3470] = ~(layer2_outputs[10593]) | (layer2_outputs[9048]);
    assign outputs[3471] = ~(layer2_outputs[6333]);
    assign outputs[3472] = ~(layer2_outputs[10891]);
    assign outputs[3473] = ~((layer2_outputs[8787]) & (layer2_outputs[8099]));
    assign outputs[3474] = ~(layer2_outputs[6311]);
    assign outputs[3475] = ~(layer2_outputs[5701]);
    assign outputs[3476] = layer2_outputs[3088];
    assign outputs[3477] = (layer2_outputs[5791]) ^ (layer2_outputs[9555]);
    assign outputs[3478] = layer2_outputs[9721];
    assign outputs[3479] = (layer2_outputs[7430]) & ~(layer2_outputs[3197]);
    assign outputs[3480] = ~((layer2_outputs[3453]) | (layer2_outputs[9285]));
    assign outputs[3481] = ~(layer2_outputs[12269]) | (layer2_outputs[1723]);
    assign outputs[3482] = ~(layer2_outputs[4087]);
    assign outputs[3483] = ~((layer2_outputs[8208]) & (layer2_outputs[11586]));
    assign outputs[3484] = layer2_outputs[585];
    assign outputs[3485] = ~(layer2_outputs[4840]);
    assign outputs[3486] = (layer2_outputs[587]) & (layer2_outputs[4924]);
    assign outputs[3487] = ~((layer2_outputs[8131]) ^ (layer2_outputs[11423]));
    assign outputs[3488] = layer2_outputs[9320];
    assign outputs[3489] = ~(layer2_outputs[12748]);
    assign outputs[3490] = layer2_outputs[9144];
    assign outputs[3491] = ~(layer2_outputs[12578]) | (layer2_outputs[10170]);
    assign outputs[3492] = layer2_outputs[10754];
    assign outputs[3493] = ~(layer2_outputs[9457]);
    assign outputs[3494] = (layer2_outputs[11224]) | (layer2_outputs[5422]);
    assign outputs[3495] = layer2_outputs[9321];
    assign outputs[3496] = ~((layer2_outputs[4975]) ^ (layer2_outputs[10445]));
    assign outputs[3497] = ~((layer2_outputs[7648]) & (layer2_outputs[369]));
    assign outputs[3498] = layer2_outputs[1671];
    assign outputs[3499] = ~(layer2_outputs[6632]);
    assign outputs[3500] = ~(layer2_outputs[7610]);
    assign outputs[3501] = layer2_outputs[4742];
    assign outputs[3502] = layer2_outputs[4163];
    assign outputs[3503] = ~(layer2_outputs[12774]) | (layer2_outputs[9090]);
    assign outputs[3504] = (layer2_outputs[6263]) ^ (layer2_outputs[10533]);
    assign outputs[3505] = layer2_outputs[1635];
    assign outputs[3506] = layer2_outputs[8001];
    assign outputs[3507] = (layer2_outputs[12256]) ^ (layer2_outputs[4249]);
    assign outputs[3508] = ~(layer2_outputs[5706]);
    assign outputs[3509] = layer2_outputs[1346];
    assign outputs[3510] = (layer2_outputs[8366]) ^ (layer2_outputs[33]);
    assign outputs[3511] = (layer2_outputs[10508]) & ~(layer2_outputs[221]);
    assign outputs[3512] = ~(layer2_outputs[2138]);
    assign outputs[3513] = ~(layer2_outputs[1575]);
    assign outputs[3514] = ~((layer2_outputs[2894]) ^ (layer2_outputs[5215]));
    assign outputs[3515] = layer2_outputs[8191];
    assign outputs[3516] = layer2_outputs[12637];
    assign outputs[3517] = (layer2_outputs[8875]) | (layer2_outputs[4065]);
    assign outputs[3518] = (layer2_outputs[6323]) & ~(layer2_outputs[7313]);
    assign outputs[3519] = layer2_outputs[1777];
    assign outputs[3520] = ~((layer2_outputs[1259]) ^ (layer2_outputs[4898]));
    assign outputs[3521] = (layer2_outputs[10689]) & ~(layer2_outputs[2656]);
    assign outputs[3522] = ~((layer2_outputs[219]) & (layer2_outputs[100]));
    assign outputs[3523] = ~((layer2_outputs[556]) ^ (layer2_outputs[5558]));
    assign outputs[3524] = layer2_outputs[2622];
    assign outputs[3525] = ~((layer2_outputs[603]) ^ (layer2_outputs[4812]));
    assign outputs[3526] = ~(layer2_outputs[11425]);
    assign outputs[3527] = (layer2_outputs[8079]) ^ (layer2_outputs[1325]);
    assign outputs[3528] = layer2_outputs[8167];
    assign outputs[3529] = (layer2_outputs[3655]) | (layer2_outputs[4952]);
    assign outputs[3530] = ~(layer2_outputs[12298]);
    assign outputs[3531] = layer2_outputs[8876];
    assign outputs[3532] = ~(layer2_outputs[6345]);
    assign outputs[3533] = layer2_outputs[7852];
    assign outputs[3534] = layer2_outputs[11652];
    assign outputs[3535] = ~(layer2_outputs[6661]);
    assign outputs[3536] = layer2_outputs[11296];
    assign outputs[3537] = ~((layer2_outputs[4818]) & (layer2_outputs[2885]));
    assign outputs[3538] = layer2_outputs[610];
    assign outputs[3539] = ~(layer2_outputs[11029]);
    assign outputs[3540] = ~(layer2_outputs[2463]);
    assign outputs[3541] = layer2_outputs[8309];
    assign outputs[3542] = layer2_outputs[4623];
    assign outputs[3543] = (layer2_outputs[9790]) & ~(layer2_outputs[6163]);
    assign outputs[3544] = (layer2_outputs[2934]) ^ (layer2_outputs[1369]);
    assign outputs[3545] = ~((layer2_outputs[4934]) & (layer2_outputs[12400]));
    assign outputs[3546] = ~(layer2_outputs[2233]);
    assign outputs[3547] = (layer2_outputs[10429]) ^ (layer2_outputs[12012]);
    assign outputs[3548] = ~(layer2_outputs[7160]);
    assign outputs[3549] = (layer2_outputs[10316]) | (layer2_outputs[10153]);
    assign outputs[3550] = (layer2_outputs[5207]) ^ (layer2_outputs[3859]);
    assign outputs[3551] = (layer2_outputs[5023]) | (layer2_outputs[5753]);
    assign outputs[3552] = layer2_outputs[11731];
    assign outputs[3553] = (layer2_outputs[2316]) ^ (layer2_outputs[11926]);
    assign outputs[3554] = (layer2_outputs[5074]) ^ (layer2_outputs[46]);
    assign outputs[3555] = layer2_outputs[8718];
    assign outputs[3556] = ~(layer2_outputs[6526]);
    assign outputs[3557] = ~((layer2_outputs[5433]) & (layer2_outputs[911]));
    assign outputs[3558] = (layer2_outputs[5397]) & (layer2_outputs[4019]);
    assign outputs[3559] = ~((layer2_outputs[6237]) ^ (layer2_outputs[9878]));
    assign outputs[3560] = (layer2_outputs[2700]) & (layer2_outputs[8687]);
    assign outputs[3561] = ~(layer2_outputs[4207]);
    assign outputs[3562] = layer2_outputs[4830];
    assign outputs[3563] = ~(layer2_outputs[1674]);
    assign outputs[3564] = layer2_outputs[3667];
    assign outputs[3565] = layer2_outputs[8525];
    assign outputs[3566] = ~(layer2_outputs[11948]);
    assign outputs[3567] = (layer2_outputs[918]) ^ (layer2_outputs[12567]);
    assign outputs[3568] = layer2_outputs[8541];
    assign outputs[3569] = (layer2_outputs[4358]) ^ (layer2_outputs[11877]);
    assign outputs[3570] = layer2_outputs[12183];
    assign outputs[3571] = layer2_outputs[10970];
    assign outputs[3572] = ~(layer2_outputs[4153]);
    assign outputs[3573] = ~(layer2_outputs[615]);
    assign outputs[3574] = ~(layer2_outputs[11150]) | (layer2_outputs[1971]);
    assign outputs[3575] = layer2_outputs[11346];
    assign outputs[3576] = (layer2_outputs[5555]) & (layer2_outputs[7036]);
    assign outputs[3577] = ~(layer2_outputs[7896]);
    assign outputs[3578] = layer2_outputs[11547];
    assign outputs[3579] = ~(layer2_outputs[6906]);
    assign outputs[3580] = (layer2_outputs[8126]) & ~(layer2_outputs[665]);
    assign outputs[3581] = layer2_outputs[8086];
    assign outputs[3582] = ~(layer2_outputs[6522]);
    assign outputs[3583] = layer2_outputs[1328];
    assign outputs[3584] = layer2_outputs[10553];
    assign outputs[3585] = ~((layer2_outputs[4593]) ^ (layer2_outputs[7120]));
    assign outputs[3586] = (layer2_outputs[2796]) ^ (layer2_outputs[7669]);
    assign outputs[3587] = ~(layer2_outputs[1703]);
    assign outputs[3588] = ~(layer2_outputs[10009]);
    assign outputs[3589] = layer2_outputs[11137];
    assign outputs[3590] = (layer2_outputs[9813]) ^ (layer2_outputs[12720]);
    assign outputs[3591] = ~(layer2_outputs[11209]);
    assign outputs[3592] = ~(layer2_outputs[2713]) | (layer2_outputs[4530]);
    assign outputs[3593] = (layer2_outputs[10120]) | (layer2_outputs[7514]);
    assign outputs[3594] = layer2_outputs[2890];
    assign outputs[3595] = (layer2_outputs[11476]) ^ (layer2_outputs[2302]);
    assign outputs[3596] = (layer2_outputs[1733]) ^ (layer2_outputs[567]);
    assign outputs[3597] = layer2_outputs[8823];
    assign outputs[3598] = ~((layer2_outputs[5525]) & (layer2_outputs[3980]));
    assign outputs[3599] = layer2_outputs[5395];
    assign outputs[3600] = ~((layer2_outputs[12548]) | (layer2_outputs[9484]));
    assign outputs[3601] = layer2_outputs[11235];
    assign outputs[3602] = layer2_outputs[6246];
    assign outputs[3603] = (layer2_outputs[3198]) & (layer2_outputs[4814]);
    assign outputs[3604] = ~(layer2_outputs[11091]);
    assign outputs[3605] = (layer2_outputs[594]) ^ (layer2_outputs[9726]);
    assign outputs[3606] = (layer2_outputs[9470]) ^ (layer2_outputs[5188]);
    assign outputs[3607] = layer2_outputs[6123];
    assign outputs[3608] = layer2_outputs[11277];
    assign outputs[3609] = (layer2_outputs[6392]) ^ (layer2_outputs[10522]);
    assign outputs[3610] = ~(layer2_outputs[2396]);
    assign outputs[3611] = ~(layer2_outputs[9307]);
    assign outputs[3612] = ~(layer2_outputs[2016]);
    assign outputs[3613] = ~((layer2_outputs[3866]) & (layer2_outputs[7771]));
    assign outputs[3614] = (layer2_outputs[11893]) ^ (layer2_outputs[4571]);
    assign outputs[3615] = (layer2_outputs[5034]) ^ (layer2_outputs[8836]);
    assign outputs[3616] = (layer2_outputs[2021]) | (layer2_outputs[6606]);
    assign outputs[3617] = ~(layer2_outputs[11397]);
    assign outputs[3618] = layer2_outputs[1232];
    assign outputs[3619] = layer2_outputs[10031];
    assign outputs[3620] = layer2_outputs[2483];
    assign outputs[3621] = (layer2_outputs[10657]) ^ (layer2_outputs[4218]);
    assign outputs[3622] = (layer2_outputs[11007]) & ~(layer2_outputs[11280]);
    assign outputs[3623] = ~(layer2_outputs[6889]);
    assign outputs[3624] = (layer2_outputs[11084]) ^ (layer2_outputs[4072]);
    assign outputs[3625] = layer2_outputs[12643];
    assign outputs[3626] = (layer2_outputs[11376]) ^ (layer2_outputs[932]);
    assign outputs[3627] = layer2_outputs[7473];
    assign outputs[3628] = layer2_outputs[5657];
    assign outputs[3629] = (layer2_outputs[6365]) & ~(layer2_outputs[4331]);
    assign outputs[3630] = ~(layer2_outputs[1518]);
    assign outputs[3631] = ~(layer2_outputs[9254]);
    assign outputs[3632] = ~(layer2_outputs[2108]);
    assign outputs[3633] = ~(layer2_outputs[5431]);
    assign outputs[3634] = ~((layer2_outputs[10675]) & (layer2_outputs[2967]));
    assign outputs[3635] = layer2_outputs[10609];
    assign outputs[3636] = ~((layer2_outputs[6953]) ^ (layer2_outputs[2359]));
    assign outputs[3637] = ~(layer2_outputs[8393]);
    assign outputs[3638] = ~(layer2_outputs[7529]) | (layer2_outputs[2719]);
    assign outputs[3639] = ~(layer2_outputs[9955]) | (layer2_outputs[6112]);
    assign outputs[3640] = layer2_outputs[12769];
    assign outputs[3641] = (layer2_outputs[11255]) | (layer2_outputs[7506]);
    assign outputs[3642] = (layer2_outputs[10476]) ^ (layer2_outputs[11716]);
    assign outputs[3643] = (layer2_outputs[803]) & (layer2_outputs[12064]);
    assign outputs[3644] = ~((layer2_outputs[9333]) & (layer2_outputs[10232]));
    assign outputs[3645] = ~(layer2_outputs[3936]);
    assign outputs[3646] = (layer2_outputs[3283]) | (layer2_outputs[1142]);
    assign outputs[3647] = ~(layer2_outputs[8548]);
    assign outputs[3648] = layer2_outputs[9295];
    assign outputs[3649] = layer2_outputs[287];
    assign outputs[3650] = ~((layer2_outputs[11343]) ^ (layer2_outputs[7801]));
    assign outputs[3651] = (layer2_outputs[3778]) & (layer2_outputs[7325]);
    assign outputs[3652] = layer2_outputs[11600];
    assign outputs[3653] = ~(layer2_outputs[7719]);
    assign outputs[3654] = ~(layer2_outputs[7944]);
    assign outputs[3655] = (layer2_outputs[9910]) ^ (layer2_outputs[7460]);
    assign outputs[3656] = ~((layer2_outputs[7954]) ^ (layer2_outputs[3365]));
    assign outputs[3657] = layer2_outputs[9444];
    assign outputs[3658] = ~(layer2_outputs[10182]);
    assign outputs[3659] = (layer2_outputs[8392]) ^ (layer2_outputs[3724]);
    assign outputs[3660] = ~(layer2_outputs[597]);
    assign outputs[3661] = ~(layer2_outputs[6725]) | (layer2_outputs[5922]);
    assign outputs[3662] = ~(layer2_outputs[6448]);
    assign outputs[3663] = ~(layer2_outputs[4539]);
    assign outputs[3664] = ~(layer2_outputs[2742]);
    assign outputs[3665] = layer2_outputs[3719];
    assign outputs[3666] = ~(layer2_outputs[3332]);
    assign outputs[3667] = layer2_outputs[7320];
    assign outputs[3668] = layer2_outputs[4440];
    assign outputs[3669] = ~(layer2_outputs[920]) | (layer2_outputs[11447]);
    assign outputs[3670] = (layer2_outputs[12125]) ^ (layer2_outputs[7911]);
    assign outputs[3671] = ~(layer2_outputs[621]);
    assign outputs[3672] = (layer2_outputs[2188]) & (layer2_outputs[1362]);
    assign outputs[3673] = layer2_outputs[10718];
    assign outputs[3674] = ~(layer2_outputs[12745]);
    assign outputs[3675] = layer2_outputs[883];
    assign outputs[3676] = ~(layer2_outputs[786]) | (layer2_outputs[7635]);
    assign outputs[3677] = ~(layer2_outputs[612]);
    assign outputs[3678] = (layer2_outputs[1165]) ^ (layer2_outputs[8063]);
    assign outputs[3679] = ~(layer2_outputs[6835]);
    assign outputs[3680] = layer2_outputs[9651];
    assign outputs[3681] = (layer2_outputs[9288]) ^ (layer2_outputs[7296]);
    assign outputs[3682] = layer2_outputs[2673];
    assign outputs[3683] = layer2_outputs[9536];
    assign outputs[3684] = layer2_outputs[1766];
    assign outputs[3685] = (layer2_outputs[4987]) & ~(layer2_outputs[955]);
    assign outputs[3686] = (layer2_outputs[12722]) ^ (layer2_outputs[5972]);
    assign outputs[3687] = ~(layer2_outputs[11023]);
    assign outputs[3688] = layer2_outputs[4056];
    assign outputs[3689] = ~(layer2_outputs[12380]) | (layer2_outputs[780]);
    assign outputs[3690] = layer2_outputs[3210];
    assign outputs[3691] = ~(layer2_outputs[7087]) | (layer2_outputs[10965]);
    assign outputs[3692] = (layer2_outputs[4592]) & ~(layer2_outputs[2595]);
    assign outputs[3693] = ~(layer2_outputs[8248]);
    assign outputs[3694] = layer2_outputs[2872];
    assign outputs[3695] = (layer2_outputs[1278]) & (layer2_outputs[11807]);
    assign outputs[3696] = (layer2_outputs[2807]) ^ (layer2_outputs[6299]);
    assign outputs[3697] = ~((layer2_outputs[1531]) & (layer2_outputs[1444]));
    assign outputs[3698] = layer2_outputs[6798];
    assign outputs[3699] = (layer2_outputs[9087]) ^ (layer2_outputs[3292]);
    assign outputs[3700] = ~(layer2_outputs[3537]);
    assign outputs[3701] = ~(layer2_outputs[5110]);
    assign outputs[3702] = layer2_outputs[11144];
    assign outputs[3703] = (layer2_outputs[8630]) | (layer2_outputs[3091]);
    assign outputs[3704] = ~((layer2_outputs[5076]) ^ (layer2_outputs[3772]));
    assign outputs[3705] = ~(layer2_outputs[3869]);
    assign outputs[3706] = layer2_outputs[4220];
    assign outputs[3707] = (layer2_outputs[967]) ^ (layer2_outputs[2036]);
    assign outputs[3708] = ~(layer2_outputs[3553]);
    assign outputs[3709] = layer2_outputs[2919];
    assign outputs[3710] = (layer2_outputs[4969]) ^ (layer2_outputs[5237]);
    assign outputs[3711] = layer2_outputs[4341];
    assign outputs[3712] = ~((layer2_outputs[9394]) ^ (layer2_outputs[3919]));
    assign outputs[3713] = ~(layer2_outputs[9666]);
    assign outputs[3714] = layer2_outputs[11188];
    assign outputs[3715] = layer2_outputs[10571];
    assign outputs[3716] = layer2_outputs[9977];
    assign outputs[3717] = layer2_outputs[2352];
    assign outputs[3718] = layer2_outputs[9268];
    assign outputs[3719] = ~(layer2_outputs[7344]);
    assign outputs[3720] = ~((layer2_outputs[2029]) ^ (layer2_outputs[5522]));
    assign outputs[3721] = layer2_outputs[1713];
    assign outputs[3722] = ~(layer2_outputs[7598]);
    assign outputs[3723] = (layer2_outputs[5692]) ^ (layer2_outputs[3762]);
    assign outputs[3724] = (layer2_outputs[2134]) | (layer2_outputs[5961]);
    assign outputs[3725] = ~(layer2_outputs[11913]);
    assign outputs[3726] = ~((layer2_outputs[2430]) & (layer2_outputs[4528]));
    assign outputs[3727] = ~(layer2_outputs[4776]);
    assign outputs[3728] = (layer2_outputs[4547]) ^ (layer2_outputs[3513]);
    assign outputs[3729] = (layer2_outputs[1648]) | (layer2_outputs[8023]);
    assign outputs[3730] = layer2_outputs[959];
    assign outputs[3731] = layer2_outputs[11776];
    assign outputs[3732] = layer2_outputs[4971];
    assign outputs[3733] = (layer2_outputs[7136]) & ~(layer2_outputs[9040]);
    assign outputs[3734] = ~(layer2_outputs[12458]);
    assign outputs[3735] = ~(layer2_outputs[8773]);
    assign outputs[3736] = layer2_outputs[6487];
    assign outputs[3737] = layer2_outputs[2971];
    assign outputs[3738] = ~((layer2_outputs[10665]) ^ (layer2_outputs[7043]));
    assign outputs[3739] = (layer2_outputs[2263]) & ~(layer2_outputs[2265]);
    assign outputs[3740] = (layer2_outputs[6974]) ^ (layer2_outputs[6794]);
    assign outputs[3741] = ~(layer2_outputs[10011]);
    assign outputs[3742] = layer2_outputs[4876];
    assign outputs[3743] = ~(layer2_outputs[4584]);
    assign outputs[3744] = (layer2_outputs[7197]) ^ (layer2_outputs[7030]);
    assign outputs[3745] = ~(layer2_outputs[9794]);
    assign outputs[3746] = layer2_outputs[5472];
    assign outputs[3747] = ~(layer2_outputs[11705]);
    assign outputs[3748] = ~(layer2_outputs[9482]);
    assign outputs[3749] = layer2_outputs[6672];
    assign outputs[3750] = ~(layer2_outputs[6623]);
    assign outputs[3751] = (layer2_outputs[9974]) ^ (layer2_outputs[10682]);
    assign outputs[3752] = ~(layer2_outputs[8405]);
    assign outputs[3753] = ~((layer2_outputs[7609]) ^ (layer2_outputs[1294]));
    assign outputs[3754] = (layer2_outputs[11626]) ^ (layer2_outputs[3401]);
    assign outputs[3755] = ~(layer2_outputs[987]);
    assign outputs[3756] = ~((layer2_outputs[3679]) | (layer2_outputs[1513]));
    assign outputs[3757] = ~(layer2_outputs[9825]);
    assign outputs[3758] = layer2_outputs[9722];
    assign outputs[3759] = ~(layer2_outputs[11814]) | (layer2_outputs[12059]);
    assign outputs[3760] = ~((layer2_outputs[2896]) ^ (layer2_outputs[10496]));
    assign outputs[3761] = layer2_outputs[7519];
    assign outputs[3762] = layer2_outputs[12356];
    assign outputs[3763] = layer2_outputs[2569];
    assign outputs[3764] = ~((layer2_outputs[295]) ^ (layer2_outputs[1808]));
    assign outputs[3765] = ~(layer2_outputs[11461]);
    assign outputs[3766] = ~(layer2_outputs[7469]) | (layer2_outputs[774]);
    assign outputs[3767] = ~(layer2_outputs[5923]);
    assign outputs[3768] = ~(layer2_outputs[5795]);
    assign outputs[3769] = ~((layer2_outputs[3023]) ^ (layer2_outputs[12584]));
    assign outputs[3770] = layer2_outputs[12651];
    assign outputs[3771] = (layer2_outputs[1484]) ^ (layer2_outputs[6867]);
    assign outputs[3772] = ~((layer2_outputs[9670]) ^ (layer2_outputs[11222]));
    assign outputs[3773] = ~((layer2_outputs[12000]) & (layer2_outputs[4030]));
    assign outputs[3774] = layer2_outputs[12279];
    assign outputs[3775] = (layer2_outputs[1884]) ^ (layer2_outputs[11180]);
    assign outputs[3776] = layer2_outputs[8466];
    assign outputs[3777] = layer2_outputs[8212];
    assign outputs[3778] = ~(layer2_outputs[4479]);
    assign outputs[3779] = ~(layer2_outputs[3872]);
    assign outputs[3780] = layer2_outputs[7276];
    assign outputs[3781] = ~(layer2_outputs[2755]);
    assign outputs[3782] = layer2_outputs[11096];
    assign outputs[3783] = layer2_outputs[4655];
    assign outputs[3784] = ~(layer2_outputs[12181]) | (layer2_outputs[5754]);
    assign outputs[3785] = ~((layer2_outputs[11156]) ^ (layer2_outputs[2306]));
    assign outputs[3786] = ~(layer2_outputs[4426]);
    assign outputs[3787] = ~(layer2_outputs[4432]);
    assign outputs[3788] = ~(layer2_outputs[1573]);
    assign outputs[3789] = ~(layer2_outputs[4161]);
    assign outputs[3790] = ~(layer2_outputs[7229]) | (layer2_outputs[1666]);
    assign outputs[3791] = (layer2_outputs[9543]) & ~(layer2_outputs[6398]);
    assign outputs[3792] = ~(layer2_outputs[1263]);
    assign outputs[3793] = layer2_outputs[505];
    assign outputs[3794] = (layer2_outputs[2644]) & ~(layer2_outputs[5071]);
    assign outputs[3795] = ~(layer2_outputs[11202]);
    assign outputs[3796] = layer2_outputs[2163];
    assign outputs[3797] = ~(layer2_outputs[2865]);
    assign outputs[3798] = (layer2_outputs[3208]) ^ (layer2_outputs[10694]);
    assign outputs[3799] = (layer2_outputs[8337]) & ~(layer2_outputs[6932]);
    assign outputs[3800] = layer2_outputs[2763];
    assign outputs[3801] = ~((layer2_outputs[2234]) ^ (layer2_outputs[10421]));
    assign outputs[3802] = layer2_outputs[5928];
    assign outputs[3803] = ~((layer2_outputs[3087]) ^ (layer2_outputs[4572]));
    assign outputs[3804] = ~(layer2_outputs[486]) | (layer2_outputs[12259]);
    assign outputs[3805] = ~((layer2_outputs[3815]) ^ (layer2_outputs[12473]));
    assign outputs[3806] = ~(layer2_outputs[3786]);
    assign outputs[3807] = ~(layer2_outputs[3104]);
    assign outputs[3808] = ~((layer2_outputs[6821]) ^ (layer2_outputs[8170]));
    assign outputs[3809] = ~(layer2_outputs[9286]);
    assign outputs[3810] = (layer2_outputs[7166]) ^ (layer2_outputs[7038]);
    assign outputs[3811] = ~(layer2_outputs[5040]) | (layer2_outputs[10964]);
    assign outputs[3812] = ~(layer2_outputs[9469]);
    assign outputs[3813] = layer2_outputs[3670];
    assign outputs[3814] = layer2_outputs[10063];
    assign outputs[3815] = ~(layer2_outputs[10887]) | (layer2_outputs[4412]);
    assign outputs[3816] = ~((layer2_outputs[2212]) ^ (layer2_outputs[8251]));
    assign outputs[3817] = ~((layer2_outputs[5077]) ^ (layer2_outputs[249]));
    assign outputs[3818] = ~(layer2_outputs[5829]) | (layer2_outputs[8650]);
    assign outputs[3819] = ~(layer2_outputs[7008]);
    assign outputs[3820] = ~((layer2_outputs[10277]) & (layer2_outputs[3362]));
    assign outputs[3821] = ~(layer2_outputs[6318]);
    assign outputs[3822] = ~(layer2_outputs[8148]);
    assign outputs[3823] = layer2_outputs[48];
    assign outputs[3824] = (layer2_outputs[4859]) ^ (layer2_outputs[2195]);
    assign outputs[3825] = ~(layer2_outputs[4443]);
    assign outputs[3826] = ~(layer2_outputs[12036]);
    assign outputs[3827] = (layer2_outputs[2080]) ^ (layer2_outputs[8050]);
    assign outputs[3828] = ~(layer2_outputs[4529]);
    assign outputs[3829] = (layer2_outputs[5341]) ^ (layer2_outputs[1109]);
    assign outputs[3830] = ~(layer2_outputs[943]);
    assign outputs[3831] = layer2_outputs[1782];
    assign outputs[3832] = ~(layer2_outputs[10737]) | (layer2_outputs[3047]);
    assign outputs[3833] = ~(layer2_outputs[7132]);
    assign outputs[3834] = (layer2_outputs[3068]) | (layer2_outputs[411]);
    assign outputs[3835] = layer2_outputs[7958];
    assign outputs[3836] = ~(layer2_outputs[6593]) | (layer2_outputs[9554]);
    assign outputs[3837] = ~(layer2_outputs[7996]);
    assign outputs[3838] = layer2_outputs[2242];
    assign outputs[3839] = ~(layer2_outputs[12313]);
    assign outputs[3840] = (layer2_outputs[5056]) & (layer2_outputs[618]);
    assign outputs[3841] = ~(layer2_outputs[12313]);
    assign outputs[3842] = layer2_outputs[4737];
    assign outputs[3843] = layer2_outputs[4175];
    assign outputs[3844] = ~((layer2_outputs[5984]) & (layer2_outputs[12703]));
    assign outputs[3845] = layer2_outputs[12194];
    assign outputs[3846] = ~((layer2_outputs[8315]) ^ (layer2_outputs[6397]));
    assign outputs[3847] = ~((layer2_outputs[3893]) ^ (layer2_outputs[3853]));
    assign outputs[3848] = (layer2_outputs[3145]) ^ (layer2_outputs[10092]);
    assign outputs[3849] = ~((layer2_outputs[4687]) ^ (layer2_outputs[7932]));
    assign outputs[3850] = layer2_outputs[7080];
    assign outputs[3851] = ~(layer2_outputs[6201]);
    assign outputs[3852] = layer2_outputs[2057];
    assign outputs[3853] = ~(layer2_outputs[11895]);
    assign outputs[3854] = ~((layer2_outputs[9174]) ^ (layer2_outputs[6041]));
    assign outputs[3855] = layer2_outputs[11311];
    assign outputs[3856] = (layer2_outputs[6605]) & (layer2_outputs[8811]);
    assign outputs[3857] = ~(layer2_outputs[5135]);
    assign outputs[3858] = layer2_outputs[2691];
    assign outputs[3859] = layer2_outputs[7];
    assign outputs[3860] = ~(layer2_outputs[1262]);
    assign outputs[3861] = layer2_outputs[7033];
    assign outputs[3862] = ~((layer2_outputs[6964]) ^ (layer2_outputs[3829]));
    assign outputs[3863] = layer2_outputs[7330];
    assign outputs[3864] = ~(layer2_outputs[11975]);
    assign outputs[3865] = layer2_outputs[1296];
    assign outputs[3866] = ~((layer2_outputs[7799]) ^ (layer2_outputs[4401]));
    assign outputs[3867] = ~(layer2_outputs[9982]);
    assign outputs[3868] = (layer2_outputs[6169]) ^ (layer2_outputs[6221]);
    assign outputs[3869] = layer2_outputs[3506];
    assign outputs[3870] = layer2_outputs[7098];
    assign outputs[3871] = ~(layer2_outputs[4371]);
    assign outputs[3872] = layer2_outputs[5651];
    assign outputs[3873] = layer2_outputs[10880];
    assign outputs[3874] = (layer2_outputs[6766]) ^ (layer2_outputs[1184]);
    assign outputs[3875] = layer2_outputs[4970];
    assign outputs[3876] = ~(layer2_outputs[12504]);
    assign outputs[3877] = ~(layer2_outputs[11776]);
    assign outputs[3878] = ~((layer2_outputs[6103]) | (layer2_outputs[5723]));
    assign outputs[3879] = ~(layer2_outputs[3126]);
    assign outputs[3880] = ~(layer2_outputs[10329]) | (layer2_outputs[7800]);
    assign outputs[3881] = (layer2_outputs[10818]) ^ (layer2_outputs[11919]);
    assign outputs[3882] = ~(layer2_outputs[3380]) | (layer2_outputs[6307]);
    assign outputs[3883] = ~(layer2_outputs[8375]);
    assign outputs[3884] = ~(layer2_outputs[10883]);
    assign outputs[3885] = (layer2_outputs[12244]) | (layer2_outputs[11747]);
    assign outputs[3886] = layer2_outputs[11020];
    assign outputs[3887] = ~(layer2_outputs[6978]);
    assign outputs[3888] = ~((layer2_outputs[6194]) | (layer2_outputs[7251]));
    assign outputs[3889] = layer2_outputs[3165];
    assign outputs[3890] = ~((layer2_outputs[4427]) ^ (layer2_outputs[12568]));
    assign outputs[3891] = (layer2_outputs[9797]) ^ (layer2_outputs[8958]);
    assign outputs[3892] = (layer2_outputs[11316]) & ~(layer2_outputs[4856]);
    assign outputs[3893] = ~((layer2_outputs[2721]) ^ (layer2_outputs[11596]));
    assign outputs[3894] = layer2_outputs[12705];
    assign outputs[3895] = (layer2_outputs[2141]) & ~(layer2_outputs[5921]);
    assign outputs[3896] = layer2_outputs[5284];
    assign outputs[3897] = ~((layer2_outputs[2709]) ^ (layer2_outputs[2193]));
    assign outputs[3898] = ~(layer2_outputs[7060]);
    assign outputs[3899] = layer2_outputs[1041];
    assign outputs[3900] = ~(layer2_outputs[9839]);
    assign outputs[3901] = (layer2_outputs[9820]) ^ (layer2_outputs[5471]);
    assign outputs[3902] = layer2_outputs[5965];
    assign outputs[3903] = ~(layer2_outputs[5653]);
    assign outputs[3904] = layer2_outputs[3331];
    assign outputs[3905] = ~(layer2_outputs[9193]);
    assign outputs[3906] = layer2_outputs[12659];
    assign outputs[3907] = ~((layer2_outputs[12487]) ^ (layer2_outputs[1103]));
    assign outputs[3908] = layer2_outputs[3347];
    assign outputs[3909] = ~((layer2_outputs[6876]) ^ (layer2_outputs[10412]));
    assign outputs[3910] = layer2_outputs[11157];
    assign outputs[3911] = (layer2_outputs[1589]) & (layer2_outputs[4315]);
    assign outputs[3912] = (layer2_outputs[740]) ^ (layer2_outputs[3159]);
    assign outputs[3913] = (layer2_outputs[7639]) | (layer2_outputs[11918]);
    assign outputs[3914] = ~(layer2_outputs[313]);
    assign outputs[3915] = (layer2_outputs[9209]) ^ (layer2_outputs[11042]);
    assign outputs[3916] = layer2_outputs[4327];
    assign outputs[3917] = (layer2_outputs[12099]) & ~(layer2_outputs[6220]);
    assign outputs[3918] = (layer2_outputs[5333]) & ~(layer2_outputs[8482]);
    assign outputs[3919] = ~(layer2_outputs[10394]);
    assign outputs[3920] = layer2_outputs[8572];
    assign outputs[3921] = layer2_outputs[10722];
    assign outputs[3922] = ~(layer2_outputs[2385]);
    assign outputs[3923] = ~(layer2_outputs[3086]);
    assign outputs[3924] = ~(layer2_outputs[3468]);
    assign outputs[3925] = ~(layer2_outputs[7408]);
    assign outputs[3926] = layer2_outputs[9132];
    assign outputs[3927] = layer2_outputs[2200];
    assign outputs[3928] = ~(layer2_outputs[2336]);
    assign outputs[3929] = layer2_outputs[10557];
    assign outputs[3930] = ~((layer2_outputs[6019]) ^ (layer2_outputs[10532]));
    assign outputs[3931] = (layer2_outputs[5120]) ^ (layer2_outputs[8098]);
    assign outputs[3932] = ~((layer2_outputs[3956]) ^ (layer2_outputs[11916]));
    assign outputs[3933] = (layer2_outputs[6400]) ^ (layer2_outputs[11310]);
    assign outputs[3934] = ~((layer2_outputs[7830]) ^ (layer2_outputs[6134]));
    assign outputs[3935] = (layer2_outputs[11558]) ^ (layer2_outputs[1711]);
    assign outputs[3936] = ~(layer2_outputs[7983]);
    assign outputs[3937] = (layer2_outputs[1558]) ^ (layer2_outputs[5220]);
    assign outputs[3938] = ~(layer2_outputs[5600]);
    assign outputs[3939] = ~((layer2_outputs[6559]) ^ (layer2_outputs[12361]));
    assign outputs[3940] = ~(layer2_outputs[2919]);
    assign outputs[3941] = (layer2_outputs[8354]) ^ (layer2_outputs[1399]);
    assign outputs[3942] = layer2_outputs[6537];
    assign outputs[3943] = ~((layer2_outputs[9950]) ^ (layer2_outputs[440]));
    assign outputs[3944] = (layer2_outputs[7284]) ^ (layer2_outputs[3397]);
    assign outputs[3945] = ~((layer2_outputs[12482]) ^ (layer2_outputs[8473]));
    assign outputs[3946] = (layer2_outputs[1319]) & ~(layer2_outputs[12765]);
    assign outputs[3947] = (layer2_outputs[12038]) & ~(layer2_outputs[8404]);
    assign outputs[3948] = layer2_outputs[5704];
    assign outputs[3949] = ~((layer2_outputs[7665]) ^ (layer2_outputs[6491]));
    assign outputs[3950] = ~(layer2_outputs[6523]);
    assign outputs[3951] = ~(layer2_outputs[12717]);
    assign outputs[3952] = ~((layer2_outputs[12102]) ^ (layer2_outputs[9278]));
    assign outputs[3953] = ~(layer2_outputs[9659]);
    assign outputs[3954] = layer2_outputs[5519];
    assign outputs[3955] = ~(layer2_outputs[8246]);
    assign outputs[3956] = ~((layer2_outputs[10575]) | (layer2_outputs[1527]));
    assign outputs[3957] = ~(layer2_outputs[2686]);
    assign outputs[3958] = layer2_outputs[10388];
    assign outputs[3959] = ~(layer2_outputs[12488]) | (layer2_outputs[10123]);
    assign outputs[3960] = layer2_outputs[791];
    assign outputs[3961] = ~(layer2_outputs[537]) | (layer2_outputs[235]);
    assign outputs[3962] = layer2_outputs[11531];
    assign outputs[3963] = ~(layer2_outputs[12536]);
    assign outputs[3964] = ~((layer2_outputs[4330]) | (layer2_outputs[10855]));
    assign outputs[3965] = ~((layer2_outputs[442]) ^ (layer2_outputs[11009]));
    assign outputs[3966] = ~(layer2_outputs[6794]);
    assign outputs[3967] = ~(layer2_outputs[5695]);
    assign outputs[3968] = ~((layer2_outputs[11290]) ^ (layer2_outputs[6980]));
    assign outputs[3969] = ~((layer2_outputs[4787]) ^ (layer2_outputs[2884]));
    assign outputs[3970] = layer2_outputs[12013];
    assign outputs[3971] = ~(layer2_outputs[4309]);
    assign outputs[3972] = (layer2_outputs[3266]) ^ (layer2_outputs[7486]);
    assign outputs[3973] = layer2_outputs[9459];
    assign outputs[3974] = ~(layer2_outputs[8936]) | (layer2_outputs[11469]);
    assign outputs[3975] = layer2_outputs[10885];
    assign outputs[3976] = ~((layer2_outputs[4841]) & (layer2_outputs[10073]));
    assign outputs[3977] = ~(layer2_outputs[9599]) | (layer2_outputs[8506]);
    assign outputs[3978] = ~(layer2_outputs[7470]);
    assign outputs[3979] = ~(layer2_outputs[97]);
    assign outputs[3980] = (layer2_outputs[8780]) & ~(layer2_outputs[2026]);
    assign outputs[3981] = layer2_outputs[301];
    assign outputs[3982] = layer2_outputs[6644];
    assign outputs[3983] = ~(layer2_outputs[3896]);
    assign outputs[3984] = layer2_outputs[3623];
    assign outputs[3985] = layer2_outputs[11844];
    assign outputs[3986] = layer2_outputs[11897];
    assign outputs[3987] = ~((layer2_outputs[10931]) ^ (layer2_outputs[11934]));
    assign outputs[3988] = (layer2_outputs[866]) & (layer2_outputs[6068]);
    assign outputs[3989] = ~((layer2_outputs[4508]) | (layer2_outputs[2324]));
    assign outputs[3990] = (layer2_outputs[11768]) ^ (layer2_outputs[2495]);
    assign outputs[3991] = ~((layer2_outputs[8973]) ^ (layer2_outputs[6547]));
    assign outputs[3992] = ~(layer2_outputs[12165]);
    assign outputs[3993] = layer2_outputs[12507];
    assign outputs[3994] = (layer2_outputs[9983]) & ~(layer2_outputs[6288]);
    assign outputs[3995] = layer2_outputs[2605];
    assign outputs[3996] = ~(layer2_outputs[8554]);
    assign outputs[3997] = ~(layer2_outputs[4490]);
    assign outputs[3998] = (layer2_outputs[4426]) | (layer2_outputs[12754]);
    assign outputs[3999] = (layer2_outputs[3218]) & (layer2_outputs[8492]);
    assign outputs[4000] = (layer2_outputs[12171]) & (layer2_outputs[12747]);
    assign outputs[4001] = ~(layer2_outputs[1635]);
    assign outputs[4002] = layer2_outputs[9393];
    assign outputs[4003] = (layer2_outputs[7595]) ^ (layer2_outputs[9735]);
    assign outputs[4004] = (layer2_outputs[3865]) & (layer2_outputs[3844]);
    assign outputs[4005] = (layer2_outputs[1581]) ^ (layer2_outputs[10854]);
    assign outputs[4006] = ~(layer2_outputs[6241]);
    assign outputs[4007] = layer2_outputs[3815];
    assign outputs[4008] = ~(layer2_outputs[7465]);
    assign outputs[4009] = layer2_outputs[10957];
    assign outputs[4010] = ~(layer2_outputs[6886]);
    assign outputs[4011] = ~(layer2_outputs[10474]) | (layer2_outputs[672]);
    assign outputs[4012] = layer2_outputs[5828];
    assign outputs[4013] = ~(layer2_outputs[10202]);
    assign outputs[4014] = (layer2_outputs[7330]) & ~(layer2_outputs[112]);
    assign outputs[4015] = layer2_outputs[10089];
    assign outputs[4016] = layer2_outputs[8925];
    assign outputs[4017] = layer2_outputs[9844];
    assign outputs[4018] = layer2_outputs[2757];
    assign outputs[4019] = (layer2_outputs[421]) ^ (layer2_outputs[8203]);
    assign outputs[4020] = (layer2_outputs[7872]) ^ (layer2_outputs[8494]);
    assign outputs[4021] = (layer2_outputs[4944]) ^ (layer2_outputs[8322]);
    assign outputs[4022] = (layer2_outputs[8839]) & ~(layer2_outputs[1659]);
    assign outputs[4023] = ~(layer2_outputs[9411]);
    assign outputs[4024] = ~(layer2_outputs[10217]);
    assign outputs[4025] = ~(layer2_outputs[8988]);
    assign outputs[4026] = ~(layer2_outputs[10995]);
    assign outputs[4027] = ~(layer2_outputs[450]);
    assign outputs[4028] = (layer2_outputs[3508]) ^ (layer2_outputs[8267]);
    assign outputs[4029] = ~((layer2_outputs[1678]) ^ (layer2_outputs[3593]));
    assign outputs[4030] = (layer2_outputs[3511]) ^ (layer2_outputs[492]);
    assign outputs[4031] = layer2_outputs[8837];
    assign outputs[4032] = ~(layer2_outputs[2292]);
    assign outputs[4033] = ~(layer2_outputs[3793]);
    assign outputs[4034] = (layer2_outputs[6498]) | (layer2_outputs[311]);
    assign outputs[4035] = layer2_outputs[2714];
    assign outputs[4036] = layer2_outputs[12735];
    assign outputs[4037] = (layer2_outputs[10366]) & ~(layer2_outputs[10631]);
    assign outputs[4038] = ~(layer2_outputs[4136]);
    assign outputs[4039] = ~((layer2_outputs[7907]) ^ (layer2_outputs[12066]));
    assign outputs[4040] = (layer2_outputs[3570]) & (layer2_outputs[5336]);
    assign outputs[4041] = (layer2_outputs[10116]) & ~(layer2_outputs[2823]);
    assign outputs[4042] = ~((layer2_outputs[493]) ^ (layer2_outputs[80]));
    assign outputs[4043] = layer2_outputs[164];
    assign outputs[4044] = ~(layer2_outputs[4898]);
    assign outputs[4045] = ~(layer2_outputs[8736]) | (layer2_outputs[4740]);
    assign outputs[4046] = ~((layer2_outputs[8841]) ^ (layer2_outputs[6842]));
    assign outputs[4047] = layer2_outputs[7714];
    assign outputs[4048] = (layer2_outputs[2444]) ^ (layer2_outputs[4903]);
    assign outputs[4049] = layer2_outputs[5955];
    assign outputs[4050] = (layer2_outputs[3082]) ^ (layer2_outputs[3628]);
    assign outputs[4051] = ~(layer2_outputs[692]);
    assign outputs[4052] = (layer2_outputs[7753]) ^ (layer2_outputs[6332]);
    assign outputs[4053] = ~(layer2_outputs[1002]);
    assign outputs[4054] = (layer2_outputs[370]) | (layer2_outputs[436]);
    assign outputs[4055] = (layer2_outputs[1040]) ^ (layer2_outputs[12379]);
    assign outputs[4056] = ~(layer2_outputs[12185]) | (layer2_outputs[9140]);
    assign outputs[4057] = layer2_outputs[9302];
    assign outputs[4058] = ~(layer2_outputs[5652]);
    assign outputs[4059] = layer2_outputs[3673];
    assign outputs[4060] = ~(layer2_outputs[8640]);
    assign outputs[4061] = (layer2_outputs[1989]) ^ (layer2_outputs[8306]);
    assign outputs[4062] = layer2_outputs[10574];
    assign outputs[4063] = ~(layer2_outputs[5107]);
    assign outputs[4064] = ~((layer2_outputs[8576]) | (layer2_outputs[1914]));
    assign outputs[4065] = (layer2_outputs[9902]) & ~(layer2_outputs[2950]);
    assign outputs[4066] = ~(layer2_outputs[2529]);
    assign outputs[4067] = layer2_outputs[5565];
    assign outputs[4068] = layer2_outputs[1799];
    assign outputs[4069] = ~((layer2_outputs[4348]) ^ (layer2_outputs[9167]));
    assign outputs[4070] = ~((layer2_outputs[8733]) ^ (layer2_outputs[6987]));
    assign outputs[4071] = ~((layer2_outputs[11688]) ^ (layer2_outputs[10803]));
    assign outputs[4072] = (layer2_outputs[2273]) ^ (layer2_outputs[9786]);
    assign outputs[4073] = (layer2_outputs[12320]) & ~(layer2_outputs[9500]);
    assign outputs[4074] = layer2_outputs[2314];
    assign outputs[4075] = ~((layer2_outputs[9202]) ^ (layer2_outputs[9715]));
    assign outputs[4076] = (layer2_outputs[1787]) ^ (layer2_outputs[2340]);
    assign outputs[4077] = (layer2_outputs[10034]) & ~(layer2_outputs[10143]);
    assign outputs[4078] = (layer2_outputs[12062]) ^ (layer2_outputs[3848]);
    assign outputs[4079] = (layer2_outputs[7105]) ^ (layer2_outputs[982]);
    assign outputs[4080] = (layer2_outputs[7897]) & ~(layer2_outputs[11837]);
    assign outputs[4081] = ~(layer2_outputs[1759]);
    assign outputs[4082] = layer2_outputs[5124];
    assign outputs[4083] = (layer2_outputs[4457]) & ~(layer2_outputs[2432]);
    assign outputs[4084] = ~((layer2_outputs[2694]) & (layer2_outputs[991]));
    assign outputs[4085] = layer2_outputs[2804];
    assign outputs[4086] = (layer2_outputs[1327]) ^ (layer2_outputs[11435]);
    assign outputs[4087] = ~((layer2_outputs[6380]) & (layer2_outputs[2696]));
    assign outputs[4088] = ~((layer2_outputs[72]) ^ (layer2_outputs[1701]));
    assign outputs[4089] = ~(layer2_outputs[12198]);
    assign outputs[4090] = ~(layer2_outputs[9581]);
    assign outputs[4091] = ~(layer2_outputs[1676]);
    assign outputs[4092] = (layer2_outputs[12552]) | (layer2_outputs[557]);
    assign outputs[4093] = (layer2_outputs[7493]) ^ (layer2_outputs[10655]);
    assign outputs[4094] = (layer2_outputs[9153]) & ~(layer2_outputs[12474]);
    assign outputs[4095] = (layer2_outputs[2903]) & (layer2_outputs[2328]);
    assign outputs[4096] = (layer2_outputs[1198]) ^ (layer2_outputs[10753]);
    assign outputs[4097] = (layer2_outputs[9369]) & (layer2_outputs[11996]);
    assign outputs[4098] = ~((layer2_outputs[8919]) & (layer2_outputs[6383]));
    assign outputs[4099] = ~((layer2_outputs[4533]) ^ (layer2_outputs[3744]));
    assign outputs[4100] = ~(layer2_outputs[12399]) | (layer2_outputs[5359]);
    assign outputs[4101] = ~((layer2_outputs[11829]) ^ (layer2_outputs[9378]));
    assign outputs[4102] = layer2_outputs[8426];
    assign outputs[4103] = layer2_outputs[6933];
    assign outputs[4104] = (layer2_outputs[4897]) ^ (layer2_outputs[6180]);
    assign outputs[4105] = ~(layer2_outputs[3890]);
    assign outputs[4106] = ~(layer2_outputs[5414]);
    assign outputs[4107] = ~(layer2_outputs[3962]);
    assign outputs[4108] = ~((layer2_outputs[5349]) ^ (layer2_outputs[5129]));
    assign outputs[4109] = layer2_outputs[7505];
    assign outputs[4110] = (layer2_outputs[5395]) & ~(layer2_outputs[1876]);
    assign outputs[4111] = ~(layer2_outputs[4047]);
    assign outputs[4112] = ~(layer2_outputs[10792]);
    assign outputs[4113] = ~((layer2_outputs[4174]) ^ (layer2_outputs[10590]));
    assign outputs[4114] = layer2_outputs[8950];
    assign outputs[4115] = ~(layer2_outputs[1147]);
    assign outputs[4116] = (layer2_outputs[12774]) & (layer2_outputs[11028]);
    assign outputs[4117] = layer2_outputs[5713];
    assign outputs[4118] = ~((layer2_outputs[5629]) ^ (layer2_outputs[2196]));
    assign outputs[4119] = (layer2_outputs[274]) ^ (layer2_outputs[6476]);
    assign outputs[4120] = (layer2_outputs[1734]) ^ (layer2_outputs[5768]);
    assign outputs[4121] = layer2_outputs[12716];
    assign outputs[4122] = layer2_outputs[5111];
    assign outputs[4123] = ~(layer2_outputs[8712]) | (layer2_outputs[3738]);
    assign outputs[4124] = layer2_outputs[6403];
    assign outputs[4125] = layer2_outputs[7002];
    assign outputs[4126] = layer2_outputs[9183];
    assign outputs[4127] = (layer2_outputs[10919]) ^ (layer2_outputs[11955]);
    assign outputs[4128] = (layer2_outputs[10105]) ^ (layer2_outputs[12532]);
    assign outputs[4129] = (layer2_outputs[8034]) & (layer2_outputs[471]);
    assign outputs[4130] = ~(layer2_outputs[1874]);
    assign outputs[4131] = ~(layer2_outputs[8199]);
    assign outputs[4132] = (layer2_outputs[10513]) ^ (layer2_outputs[6473]);
    assign outputs[4133] = (layer2_outputs[11071]) & ~(layer2_outputs[3425]);
    assign outputs[4134] = layer2_outputs[2528];
    assign outputs[4135] = layer2_outputs[7064];
    assign outputs[4136] = ~((layer2_outputs[12387]) | (layer2_outputs[2515]));
    assign outputs[4137] = layer2_outputs[12680];
    assign outputs[4138] = (layer2_outputs[8541]) & (layer2_outputs[2964]);
    assign outputs[4139] = layer2_outputs[5977];
    assign outputs[4140] = (layer2_outputs[10090]) ^ (layer2_outputs[7786]);
    assign outputs[4141] = (layer2_outputs[3611]) | (layer2_outputs[11496]);
    assign outputs[4142] = layer2_outputs[10111];
    assign outputs[4143] = layer2_outputs[7053];
    assign outputs[4144] = ~(layer2_outputs[9036]);
    assign outputs[4145] = ~((layer2_outputs[8930]) ^ (layer2_outputs[6665]));
    assign outputs[4146] = (layer2_outputs[3321]) ^ (layer2_outputs[11023]);
    assign outputs[4147] = layer2_outputs[1592];
    assign outputs[4148] = ~(layer2_outputs[5311]);
    assign outputs[4149] = layer2_outputs[10877];
    assign outputs[4150] = layer2_outputs[5350];
    assign outputs[4151] = (layer2_outputs[12246]) ^ (layer2_outputs[12220]);
    assign outputs[4152] = ~(layer2_outputs[7235]) | (layer2_outputs[188]);
    assign outputs[4153] = ~(layer2_outputs[12462]);
    assign outputs[4154] = ~(layer2_outputs[2207]);
    assign outputs[4155] = (layer2_outputs[3681]) & ~(layer2_outputs[5367]);
    assign outputs[4156] = layer2_outputs[7026];
    assign outputs[4157] = ~((layer2_outputs[10362]) ^ (layer2_outputs[8686]));
    assign outputs[4158] = ~(layer2_outputs[8009]);
    assign outputs[4159] = ~(layer2_outputs[8010]);
    assign outputs[4160] = layer2_outputs[594];
    assign outputs[4161] = (layer2_outputs[117]) ^ (layer2_outputs[1258]);
    assign outputs[4162] = (layer2_outputs[549]) & (layer2_outputs[1476]);
    assign outputs[4163] = ~(layer2_outputs[2140]);
    assign outputs[4164] = layer2_outputs[12445];
    assign outputs[4165] = ~(layer2_outputs[6165]) | (layer2_outputs[5234]);
    assign outputs[4166] = (layer2_outputs[1670]) & ~(layer2_outputs[12464]);
    assign outputs[4167] = layer2_outputs[4434];
    assign outputs[4168] = (layer2_outputs[11279]) ^ (layer2_outputs[10270]);
    assign outputs[4169] = (layer2_outputs[6299]) ^ (layer2_outputs[446]);
    assign outputs[4170] = ~(layer2_outputs[4063]);
    assign outputs[4171] = layer2_outputs[9789];
    assign outputs[4172] = (layer2_outputs[7807]) ^ (layer2_outputs[10556]);
    assign outputs[4173] = layer2_outputs[2943];
    assign outputs[4174] = ~(layer2_outputs[7776]);
    assign outputs[4175] = ~((layer2_outputs[89]) ^ (layer2_outputs[2709]));
    assign outputs[4176] = ~(layer2_outputs[6113]);
    assign outputs[4177] = ~((layer2_outputs[3860]) & (layer2_outputs[5980]));
    assign outputs[4178] = ~(layer2_outputs[4729]) | (layer2_outputs[2001]);
    assign outputs[4179] = layer2_outputs[549];
    assign outputs[4180] = layer2_outputs[7040];
    assign outputs[4181] = (layer2_outputs[3921]) ^ (layer2_outputs[4205]);
    assign outputs[4182] = ~(layer2_outputs[2044]);
    assign outputs[4183] = ~(layer2_outputs[3905]);
    assign outputs[4184] = ~(layer2_outputs[3895]);
    assign outputs[4185] = layer2_outputs[10639];
    assign outputs[4186] = (layer2_outputs[6744]) ^ (layer2_outputs[3511]);
    assign outputs[4187] = ~(layer2_outputs[7204]) | (layer2_outputs[7813]);
    assign outputs[4188] = layer2_outputs[3104];
    assign outputs[4189] = ~(layer2_outputs[233]);
    assign outputs[4190] = layer2_outputs[12616];
    assign outputs[4191] = ~(layer2_outputs[9625]);
    assign outputs[4192] = ~((layer2_outputs[11968]) | (layer2_outputs[11026]));
    assign outputs[4193] = layer2_outputs[1483];
    assign outputs[4194] = (layer2_outputs[500]) ^ (layer2_outputs[251]);
    assign outputs[4195] = layer2_outputs[10983];
    assign outputs[4196] = ~(layer2_outputs[4680]);
    assign outputs[4197] = (layer2_outputs[125]) & ~(layer2_outputs[3655]);
    assign outputs[4198] = ~(layer2_outputs[6471]);
    assign outputs[4199] = layer2_outputs[8065];
    assign outputs[4200] = layer2_outputs[5122];
    assign outputs[4201] = (layer2_outputs[12467]) & (layer2_outputs[3110]);
    assign outputs[4202] = layer2_outputs[232];
    assign outputs[4203] = ~((layer2_outputs[4551]) ^ (layer2_outputs[8232]));
    assign outputs[4204] = ~((layer2_outputs[11972]) ^ (layer2_outputs[4621]));
    assign outputs[4205] = layer2_outputs[6816];
    assign outputs[4206] = ~((layer2_outputs[5257]) | (layer2_outputs[9222]));
    assign outputs[4207] = ~(layer2_outputs[10103]);
    assign outputs[4208] = layer2_outputs[1631];
    assign outputs[4209] = layer2_outputs[8975];
    assign outputs[4210] = layer2_outputs[7373];
    assign outputs[4211] = ~((layer2_outputs[3108]) | (layer2_outputs[7634]));
    assign outputs[4212] = (layer2_outputs[12255]) ^ (layer2_outputs[10124]);
    assign outputs[4213] = layer2_outputs[10839];
    assign outputs[4214] = ~(layer2_outputs[10687]) | (layer2_outputs[1223]);
    assign outputs[4215] = layer2_outputs[8102];
    assign outputs[4216] = (layer2_outputs[3204]) ^ (layer2_outputs[5696]);
    assign outputs[4217] = ~((layer2_outputs[3856]) | (layer2_outputs[7671]));
    assign outputs[4218] = layer2_outputs[2969];
    assign outputs[4219] = ~((layer2_outputs[7857]) ^ (layer2_outputs[4810]));
    assign outputs[4220] = ~(layer2_outputs[7412]);
    assign outputs[4221] = ~(layer2_outputs[80]);
    assign outputs[4222] = layer2_outputs[5852];
    assign outputs[4223] = ~((layer2_outputs[7889]) ^ (layer2_outputs[3648]));
    assign outputs[4224] = (layer2_outputs[11256]) & (layer2_outputs[8153]);
    assign outputs[4225] = layer2_outputs[9078];
    assign outputs[4226] = layer2_outputs[9668];
    assign outputs[4227] = layer2_outputs[4626];
    assign outputs[4228] = (layer2_outputs[7987]) ^ (layer2_outputs[11506]);
    assign outputs[4229] = (layer2_outputs[8882]) ^ (layer2_outputs[8635]);
    assign outputs[4230] = layer2_outputs[10711];
    assign outputs[4231] = ~(layer2_outputs[12336]);
    assign outputs[4232] = layer2_outputs[2341];
    assign outputs[4233] = layer2_outputs[280];
    assign outputs[4234] = ~((layer2_outputs[9795]) ^ (layer2_outputs[6898]));
    assign outputs[4235] = (layer2_outputs[4074]) ^ (layer2_outputs[8184]);
    assign outputs[4236] = layer2_outputs[3213];
    assign outputs[4237] = ~(layer2_outputs[9806]);
    assign outputs[4238] = (layer2_outputs[3767]) ^ (layer2_outputs[6864]);
    assign outputs[4239] = ~(layer2_outputs[8785]);
    assign outputs[4240] = (layer2_outputs[7450]) ^ (layer2_outputs[5106]);
    assign outputs[4241] = ~((layer2_outputs[4050]) ^ (layer2_outputs[9687]));
    assign outputs[4242] = (layer2_outputs[10110]) ^ (layer2_outputs[20]);
    assign outputs[4243] = layer2_outputs[11266];
    assign outputs[4244] = layer2_outputs[11778];
    assign outputs[4245] = (layer2_outputs[10096]) ^ (layer2_outputs[6320]);
    assign outputs[4246] = ~(layer2_outputs[10276]);
    assign outputs[4247] = ~(layer2_outputs[7181]);
    assign outputs[4248] = (layer2_outputs[708]) ^ (layer2_outputs[1394]);
    assign outputs[4249] = ~(layer2_outputs[7106]);
    assign outputs[4250] = layer2_outputs[5305];
    assign outputs[4251] = ~(layer2_outputs[1933]);
    assign outputs[4252] = ~((layer2_outputs[11719]) ^ (layer2_outputs[4743]));
    assign outputs[4253] = layer2_outputs[6913];
    assign outputs[4254] = ~(layer2_outputs[11792]);
    assign outputs[4255] = (layer2_outputs[897]) ^ (layer2_outputs[4743]);
    assign outputs[4256] = ~(layer2_outputs[7847]);
    assign outputs[4257] = (layer2_outputs[7900]) & ~(layer2_outputs[12526]);
    assign outputs[4258] = ~(layer2_outputs[6453]);
    assign outputs[4259] = ~(layer2_outputs[12105]);
    assign outputs[4260] = layer2_outputs[4393];
    assign outputs[4261] = layer2_outputs[2707];
    assign outputs[4262] = ~(layer2_outputs[11514]);
    assign outputs[4263] = ~((layer2_outputs[4534]) ^ (layer2_outputs[3774]));
    assign outputs[4264] = ~(layer2_outputs[10879]);
    assign outputs[4265] = (layer2_outputs[11371]) ^ (layer2_outputs[1806]);
    assign outputs[4266] = ~((layer2_outputs[10652]) ^ (layer2_outputs[2972]));
    assign outputs[4267] = ~((layer2_outputs[6080]) | (layer2_outputs[9129]));
    assign outputs[4268] = layer2_outputs[11628];
    assign outputs[4269] = ~((layer2_outputs[3690]) ^ (layer2_outputs[12317]));
    assign outputs[4270] = layer2_outputs[1664];
    assign outputs[4271] = layer2_outputs[11047];
    assign outputs[4272] = layer2_outputs[606];
    assign outputs[4273] = (layer2_outputs[11608]) ^ (layer2_outputs[2583]);
    assign outputs[4274] = layer2_outputs[10071];
    assign outputs[4275] = ~((layer2_outputs[4415]) ^ (layer2_outputs[4191]));
    assign outputs[4276] = layer2_outputs[3871];
    assign outputs[4277] = (layer2_outputs[5053]) & ~(layer2_outputs[5538]);
    assign outputs[4278] = ~(layer2_outputs[2609]);
    assign outputs[4279] = (layer2_outputs[4012]) & (layer2_outputs[7438]);
    assign outputs[4280] = (layer2_outputs[7681]) ^ (layer2_outputs[4687]);
    assign outputs[4281] = ~(layer2_outputs[4920]);
    assign outputs[4282] = (layer2_outputs[2486]) | (layer2_outputs[583]);
    assign outputs[4283] = ~((layer2_outputs[11859]) ^ (layer2_outputs[4353]));
    assign outputs[4284] = ~((layer2_outputs[1602]) ^ (layer2_outputs[2360]));
    assign outputs[4285] = layer2_outputs[8407];
    assign outputs[4286] = (layer2_outputs[6074]) ^ (layer2_outputs[9711]);
    assign outputs[4287] = ~(layer2_outputs[11159]);
    assign outputs[4288] = layer2_outputs[8162];
    assign outputs[4289] = (layer2_outputs[9657]) ^ (layer2_outputs[10783]);
    assign outputs[4290] = (layer2_outputs[12200]) ^ (layer2_outputs[5218]);
    assign outputs[4291] = layer2_outputs[9618];
    assign outputs[4292] = layer2_outputs[9349];
    assign outputs[4293] = ~(layer2_outputs[10338]);
    assign outputs[4294] = ~((layer2_outputs[2772]) ^ (layer2_outputs[4219]));
    assign outputs[4295] = (layer2_outputs[10212]) | (layer2_outputs[8727]);
    assign outputs[4296] = (layer2_outputs[5720]) ^ (layer2_outputs[1579]);
    assign outputs[4297] = layer2_outputs[6859];
    assign outputs[4298] = layer2_outputs[1017];
    assign outputs[4299] = layer2_outputs[12514];
    assign outputs[4300] = (layer2_outputs[6133]) & ~(layer2_outputs[2923]);
    assign outputs[4301] = ~(layer2_outputs[7355]);
    assign outputs[4302] = (layer2_outputs[4400]) ^ (layer2_outputs[5098]);
    assign outputs[4303] = ~(layer2_outputs[11578]);
    assign outputs[4304] = ~((layer2_outputs[2704]) & (layer2_outputs[11851]));
    assign outputs[4305] = ~(layer2_outputs[10488]);
    assign outputs[4306] = (layer2_outputs[10876]) ^ (layer2_outputs[1364]);
    assign outputs[4307] = (layer2_outputs[1808]) ^ (layer2_outputs[8519]);
    assign outputs[4308] = (layer2_outputs[9635]) | (layer2_outputs[5708]);
    assign outputs[4309] = layer2_outputs[6722];
    assign outputs[4310] = ~(layer2_outputs[2553]);
    assign outputs[4311] = layer2_outputs[2151];
    assign outputs[4312] = (layer2_outputs[2204]) ^ (layer2_outputs[4167]);
    assign outputs[4313] = ~(layer2_outputs[1297]);
    assign outputs[4314] = ~(layer2_outputs[1904]) | (layer2_outputs[4249]);
    assign outputs[4315] = ~(layer2_outputs[713]);
    assign outputs[4316] = ~(layer2_outputs[5483]);
    assign outputs[4317] = (layer2_outputs[11407]) | (layer2_outputs[5507]);
    assign outputs[4318] = layer2_outputs[8933];
    assign outputs[4319] = ~(layer2_outputs[1920]);
    assign outputs[4320] = ~(layer2_outputs[11999]);
    assign outputs[4321] = ~((layer2_outputs[8893]) ^ (layer2_outputs[5804]));
    assign outputs[4322] = (layer2_outputs[2681]) & ~(layer2_outputs[12613]);
    assign outputs[4323] = layer2_outputs[1021];
    assign outputs[4324] = ~(layer2_outputs[8135]);
    assign outputs[4325] = ~(layer2_outputs[3173]);
    assign outputs[4326] = layer2_outputs[893];
    assign outputs[4327] = layer2_outputs[5021];
    assign outputs[4328] = layer2_outputs[4627];
    assign outputs[4329] = ~(layer2_outputs[12481]);
    assign outputs[4330] = layer2_outputs[587];
    assign outputs[4331] = (layer2_outputs[6854]) & ~(layer2_outputs[930]);
    assign outputs[4332] = ~((layer2_outputs[3071]) ^ (layer2_outputs[8632]));
    assign outputs[4333] = layer2_outputs[7262];
    assign outputs[4334] = ~((layer2_outputs[12082]) ^ (layer2_outputs[8061]));
    assign outputs[4335] = ~(layer2_outputs[4590]);
    assign outputs[4336] = ~((layer2_outputs[9259]) ^ (layer2_outputs[10304]));
    assign outputs[4337] = layer2_outputs[3418];
    assign outputs[4338] = (layer2_outputs[8678]) & ~(layer2_outputs[5821]);
    assign outputs[4339] = ~((layer2_outputs[7064]) ^ (layer2_outputs[7281]));
    assign outputs[4340] = layer2_outputs[6698];
    assign outputs[4341] = (layer2_outputs[4510]) ^ (layer2_outputs[8299]);
    assign outputs[4342] = layer2_outputs[12583];
    assign outputs[4343] = ~(layer2_outputs[2722]);
    assign outputs[4344] = ~(layer2_outputs[5532]);
    assign outputs[4345] = ~((layer2_outputs[9310]) ^ (layer2_outputs[2816]));
    assign outputs[4346] = (layer2_outputs[5179]) ^ (layer2_outputs[2464]);
    assign outputs[4347] = ~(layer2_outputs[1064]);
    assign outputs[4348] = layer2_outputs[4121];
    assign outputs[4349] = (layer2_outputs[10986]) ^ (layer2_outputs[4340]);
    assign outputs[4350] = (layer2_outputs[1745]) | (layer2_outputs[9450]);
    assign outputs[4351] = ~(layer2_outputs[11603]);
    assign outputs[4352] = layer2_outputs[7155];
    assign outputs[4353] = (layer2_outputs[6810]) ^ (layer2_outputs[11242]);
    assign outputs[4354] = (layer2_outputs[12675]) & ~(layer2_outputs[4666]);
    assign outputs[4355] = layer2_outputs[7757];
    assign outputs[4356] = layer2_outputs[8142];
    assign outputs[4357] = ~(layer2_outputs[8078]);
    assign outputs[4358] = layer2_outputs[8016];
    assign outputs[4359] = (layer2_outputs[12552]) | (layer2_outputs[9936]);
    assign outputs[4360] = ~(layer2_outputs[10678]) | (layer2_outputs[10439]);
    assign outputs[4361] = (layer2_outputs[6869]) ^ (layer2_outputs[1658]);
    assign outputs[4362] = ~(layer2_outputs[4333]) | (layer2_outputs[8235]);
    assign outputs[4363] = layer2_outputs[8549];
    assign outputs[4364] = ~((layer2_outputs[5326]) ^ (layer2_outputs[7629]));
    assign outputs[4365] = ~((layer2_outputs[12228]) ^ (layer2_outputs[2518]));
    assign outputs[4366] = ~(layer2_outputs[9803]);
    assign outputs[4367] = (layer2_outputs[5875]) ^ (layer2_outputs[8788]);
    assign outputs[4368] = (layer2_outputs[12736]) ^ (layer2_outputs[3485]);
    assign outputs[4369] = ~((layer2_outputs[11240]) ^ (layer2_outputs[109]));
    assign outputs[4370] = ~(layer2_outputs[293]);
    assign outputs[4371] = ~(layer2_outputs[3433]) | (layer2_outputs[4879]);
    assign outputs[4372] = ~(layer2_outputs[6233]);
    assign outputs[4373] = ~((layer2_outputs[1545]) ^ (layer2_outputs[846]));
    assign outputs[4374] = ~(layer2_outputs[1011]);
    assign outputs[4375] = layer2_outputs[11113];
    assign outputs[4376] = (layer2_outputs[1085]) ^ (layer2_outputs[11595]);
    assign outputs[4377] = layer2_outputs[10727];
    assign outputs[4378] = layer2_outputs[7411];
    assign outputs[4379] = ~((layer2_outputs[7556]) & (layer2_outputs[10431]));
    assign outputs[4380] = ~(layer2_outputs[7250]);
    assign outputs[4381] = (layer2_outputs[5849]) | (layer2_outputs[333]);
    assign outputs[4382] = (layer2_outputs[4926]) ^ (layer2_outputs[2841]);
    assign outputs[4383] = ~((layer2_outputs[7346]) ^ (layer2_outputs[9160]));
    assign outputs[4384] = ~(layer2_outputs[5154]);
    assign outputs[4385] = layer2_outputs[933];
    assign outputs[4386] = (layer2_outputs[11247]) ^ (layer2_outputs[5610]);
    assign outputs[4387] = ~(layer2_outputs[4410]);
    assign outputs[4388] = ~((layer2_outputs[4473]) ^ (layer2_outputs[10361]));
    assign outputs[4389] = ~(layer2_outputs[12597]);
    assign outputs[4390] = ~(layer2_outputs[7614]);
    assign outputs[4391] = layer2_outputs[728];
    assign outputs[4392] = ~((layer2_outputs[1612]) ^ (layer2_outputs[6938]));
    assign outputs[4393] = (layer2_outputs[5396]) ^ (layer2_outputs[12205]);
    assign outputs[4394] = (layer2_outputs[8481]) & ~(layer2_outputs[11968]);
    assign outputs[4395] = layer2_outputs[10804];
    assign outputs[4396] = ~(layer2_outputs[4224]);
    assign outputs[4397] = (layer2_outputs[4360]) & ~(layer2_outputs[4783]);
    assign outputs[4398] = ~(layer2_outputs[1366]) | (layer2_outputs[623]);
    assign outputs[4399] = (layer2_outputs[5347]) ^ (layer2_outputs[6535]);
    assign outputs[4400] = layer2_outputs[3200];
    assign outputs[4401] = ~((layer2_outputs[3728]) & (layer2_outputs[10661]));
    assign outputs[4402] = ~(layer2_outputs[10548]);
    assign outputs[4403] = ~((layer2_outputs[8269]) | (layer2_outputs[5592]));
    assign outputs[4404] = ~(layer2_outputs[538]);
    assign outputs[4405] = (layer2_outputs[3743]) & ~(layer2_outputs[635]);
    assign outputs[4406] = ~((layer2_outputs[8890]) ^ (layer2_outputs[4425]));
    assign outputs[4407] = layer2_outputs[6789];
    assign outputs[4408] = layer2_outputs[7920];
    assign outputs[4409] = layer2_outputs[11413];
    assign outputs[4410] = ~(layer2_outputs[6667]);
    assign outputs[4411] = layer2_outputs[600];
    assign outputs[4412] = layer2_outputs[11736];
    assign outputs[4413] = ~(layer2_outputs[6538]);
    assign outputs[4414] = layer2_outputs[7824];
    assign outputs[4415] = (layer2_outputs[10287]) ^ (layer2_outputs[5727]);
    assign outputs[4416] = ~(layer2_outputs[8674]);
    assign outputs[4417] = (layer2_outputs[10896]) ^ (layer2_outputs[6070]);
    assign outputs[4418] = ~(layer2_outputs[10280]);
    assign outputs[4419] = layer2_outputs[11916];
    assign outputs[4420] = ~((layer2_outputs[7837]) ^ (layer2_outputs[2564]));
    assign outputs[4421] = ~((layer2_outputs[1668]) ^ (layer2_outputs[10796]));
    assign outputs[4422] = ~(layer2_outputs[12533]);
    assign outputs[4423] = (layer2_outputs[2174]) & (layer2_outputs[5198]);
    assign outputs[4424] = layer2_outputs[7666];
    assign outputs[4425] = layer2_outputs[11463];
    assign outputs[4426] = ~(layer2_outputs[5798]);
    assign outputs[4427] = layer2_outputs[9535];
    assign outputs[4428] = ~(layer2_outputs[8906]);
    assign outputs[4429] = (layer2_outputs[2536]) & (layer2_outputs[3997]);
    assign outputs[4430] = (layer2_outputs[9454]) & (layer2_outputs[988]);
    assign outputs[4431] = layer2_outputs[3500];
    assign outputs[4432] = ~(layer2_outputs[7429]);
    assign outputs[4433] = ~(layer2_outputs[4768]);
    assign outputs[4434] = (layer2_outputs[7714]) & (layer2_outputs[11844]);
    assign outputs[4435] = (layer2_outputs[9927]) & ~(layer2_outputs[11692]);
    assign outputs[4436] = ~((layer2_outputs[2830]) ^ (layer2_outputs[373]));
    assign outputs[4437] = (layer2_outputs[4491]) ^ (layer2_outputs[4880]);
    assign outputs[4438] = layer2_outputs[679];
    assign outputs[4439] = ~((layer2_outputs[3595]) ^ (layer2_outputs[11637]));
    assign outputs[4440] = layer2_outputs[12411];
    assign outputs[4441] = ~((layer2_outputs[3637]) | (layer2_outputs[10559]));
    assign outputs[4442] = ~(layer2_outputs[10076]);
    assign outputs[4443] = ~(layer2_outputs[7021]) | (layer2_outputs[9273]);
    assign outputs[4444] = ~(layer2_outputs[2390]) | (layer2_outputs[607]);
    assign outputs[4445] = layer2_outputs[7729];
    assign outputs[4446] = ~(layer2_outputs[6844]) | (layer2_outputs[215]);
    assign outputs[4447] = (layer2_outputs[500]) & (layer2_outputs[2784]);
    assign outputs[4448] = ~(layer2_outputs[4319]);
    assign outputs[4449] = ~(layer2_outputs[5534]);
    assign outputs[4450] = ~(layer2_outputs[3324]);
    assign outputs[4451] = layer2_outputs[12448];
    assign outputs[4452] = ~(layer2_outputs[6893]);
    assign outputs[4453] = layer2_outputs[8308];
    assign outputs[4454] = ~((layer2_outputs[3415]) ^ (layer2_outputs[11725]));
    assign outputs[4455] = layer2_outputs[3549];
    assign outputs[4456] = ~(layer2_outputs[5233]);
    assign outputs[4457] = (layer2_outputs[12670]) & (layer2_outputs[2067]);
    assign outputs[4458] = ~(layer2_outputs[48]);
    assign outputs[4459] = layer2_outputs[6588];
    assign outputs[4460] = (layer2_outputs[7035]) ^ (layer2_outputs[11749]);
    assign outputs[4461] = ~((layer2_outputs[6306]) ^ (layer2_outputs[1619]));
    assign outputs[4462] = (layer2_outputs[8]) ^ (layer2_outputs[3201]);
    assign outputs[4463] = (layer2_outputs[1212]) & ~(layer2_outputs[2264]);
    assign outputs[4464] = (layer2_outputs[2965]) ^ (layer2_outputs[7581]);
    assign outputs[4465] = ~((layer2_outputs[12060]) ^ (layer2_outputs[10259]));
    assign outputs[4466] = layer2_outputs[1706];
    assign outputs[4467] = layer2_outputs[10070];
    assign outputs[4468] = ~((layer2_outputs[3044]) ^ (layer2_outputs[3586]));
    assign outputs[4469] = ~((layer2_outputs[4741]) ^ (layer2_outputs[1458]));
    assign outputs[4470] = layer2_outputs[4417];
    assign outputs[4471] = (layer2_outputs[5045]) & ~(layer2_outputs[11942]);
    assign outputs[4472] = (layer2_outputs[9194]) & (layer2_outputs[7383]);
    assign outputs[4473] = (layer2_outputs[1522]) & ~(layer2_outputs[1569]);
    assign outputs[4474] = ~((layer2_outputs[3097]) ^ (layer2_outputs[1718]));
    assign outputs[4475] = ~(layer2_outputs[10297]);
    assign outputs[4476] = ~(layer2_outputs[2718]);
    assign outputs[4477] = (layer2_outputs[356]) ^ (layer2_outputs[10697]);
    assign outputs[4478] = ~((layer2_outputs[11745]) ^ (layer2_outputs[2386]));
    assign outputs[4479] = layer2_outputs[12161];
    assign outputs[4480] = ~(layer2_outputs[5667]);
    assign outputs[4481] = (layer2_outputs[9541]) & (layer2_outputs[6502]);
    assign outputs[4482] = layer2_outputs[3656];
    assign outputs[4483] = ~(layer2_outputs[9770]) | (layer2_outputs[1125]);
    assign outputs[4484] = ~(layer2_outputs[5113]);
    assign outputs[4485] = ~((layer2_outputs[6441]) ^ (layer2_outputs[8788]));
    assign outputs[4486] = layer2_outputs[329];
    assign outputs[4487] = ~(layer2_outputs[12103]);
    assign outputs[4488] = ~(layer2_outputs[8566]);
    assign outputs[4489] = ~(layer2_outputs[8728]);
    assign outputs[4490] = (layer2_outputs[3037]) ^ (layer2_outputs[11923]);
    assign outputs[4491] = (layer2_outputs[11840]) ^ (layer2_outputs[9390]);
    assign outputs[4492] = ~(layer2_outputs[10210]);
    assign outputs[4493] = layer2_outputs[3469];
    assign outputs[4494] = (layer2_outputs[3165]) ^ (layer2_outputs[7003]);
    assign outputs[4495] = layer2_outputs[10566];
    assign outputs[4496] = (layer2_outputs[942]) ^ (layer2_outputs[940]);
    assign outputs[4497] = layer2_outputs[1257];
    assign outputs[4498] = (layer2_outputs[11212]) ^ (layer2_outputs[4959]);
    assign outputs[4499] = ~((layer2_outputs[765]) ^ (layer2_outputs[9060]));
    assign outputs[4500] = layer2_outputs[927];
    assign outputs[4501] = ~((layer2_outputs[3358]) ^ (layer2_outputs[7218]));
    assign outputs[4502] = (layer2_outputs[2753]) & ~(layer2_outputs[11969]);
    assign outputs[4503] = layer2_outputs[6783];
    assign outputs[4504] = (layer2_outputs[6867]) | (layer2_outputs[7667]);
    assign outputs[4505] = (layer2_outputs[1288]) ^ (layer2_outputs[5645]);
    assign outputs[4506] = ~(layer2_outputs[8123]);
    assign outputs[4507] = ~(layer2_outputs[12046]);
    assign outputs[4508] = ~((layer2_outputs[11779]) & (layer2_outputs[138]));
    assign outputs[4509] = ~(layer2_outputs[11551]);
    assign outputs[4510] = ~((layer2_outputs[1025]) | (layer2_outputs[9999]));
    assign outputs[4511] = (layer2_outputs[7663]) | (layer2_outputs[10495]);
    assign outputs[4512] = ~(layer2_outputs[5832]);
    assign outputs[4513] = ~(layer2_outputs[4181]);
    assign outputs[4514] = (layer2_outputs[8228]) & ~(layer2_outputs[4990]);
    assign outputs[4515] = ~((layer2_outputs[4961]) | (layer2_outputs[2284]));
    assign outputs[4516] = ~(layer2_outputs[12526]);
    assign outputs[4517] = layer2_outputs[7918];
    assign outputs[4518] = ~(layer2_outputs[11936]);
    assign outputs[4519] = ~(layer2_outputs[10521]) | (layer2_outputs[12312]);
    assign outputs[4520] = ~(layer2_outputs[4089]);
    assign outputs[4521] = ~(layer2_outputs[10530]);
    assign outputs[4522] = ~((layer2_outputs[2950]) | (layer2_outputs[956]));
    assign outputs[4523] = layer2_outputs[5816];
    assign outputs[4524] = ~(layer2_outputs[10641]);
    assign outputs[4525] = ~((layer2_outputs[32]) ^ (layer2_outputs[9887]));
    assign outputs[4526] = (layer2_outputs[10180]) & ~(layer2_outputs[6758]);
    assign outputs[4527] = ~(layer2_outputs[6612]);
    assign outputs[4528] = ~(layer2_outputs[6108]);
    assign outputs[4529] = (layer2_outputs[1469]) ^ (layer2_outputs[5970]);
    assign outputs[4530] = (layer2_outputs[418]) ^ (layer2_outputs[2800]);
    assign outputs[4531] = ~(layer2_outputs[10697]) | (layer2_outputs[2675]);
    assign outputs[4532] = ~((layer2_outputs[9470]) ^ (layer2_outputs[12266]));
    assign outputs[4533] = ~(layer2_outputs[483]);
    assign outputs[4534] = layer2_outputs[5732];
    assign outputs[4535] = (layer2_outputs[1816]) & (layer2_outputs[4627]);
    assign outputs[4536] = ~(layer2_outputs[6678]);
    assign outputs[4537] = (layer2_outputs[6000]) & (layer2_outputs[12795]);
    assign outputs[4538] = layer2_outputs[12078];
    assign outputs[4539] = ~(layer2_outputs[1636]);
    assign outputs[4540] = (layer2_outputs[4398]) | (layer2_outputs[10244]);
    assign outputs[4541] = layer2_outputs[9366];
    assign outputs[4542] = (layer2_outputs[5134]) & ~(layer2_outputs[12080]);
    assign outputs[4543] = layer2_outputs[646];
    assign outputs[4544] = ~(layer2_outputs[8359]);
    assign outputs[4545] = (layer2_outputs[6245]) ^ (layer2_outputs[2478]);
    assign outputs[4546] = ~(layer2_outputs[4635]);
    assign outputs[4547] = layer2_outputs[8757];
    assign outputs[4548] = ~((layer2_outputs[11782]) ^ (layer2_outputs[811]));
    assign outputs[4549] = ~(layer2_outputs[7646]);
    assign outputs[4550] = (layer2_outputs[4598]) ^ (layer2_outputs[8425]);
    assign outputs[4551] = ~((layer2_outputs[672]) ^ (layer2_outputs[2885]));
    assign outputs[4552] = ~(layer2_outputs[7646]);
    assign outputs[4553] = ~(layer2_outputs[2065]);
    assign outputs[4554] = (layer2_outputs[9589]) ^ (layer2_outputs[10197]);
    assign outputs[4555] = (layer2_outputs[2487]) ^ (layer2_outputs[2442]);
    assign outputs[4556] = (layer2_outputs[10962]) & ~(layer2_outputs[7742]);
    assign outputs[4557] = ~(layer2_outputs[1998]);
    assign outputs[4558] = (layer2_outputs[2704]) ^ (layer2_outputs[2653]);
    assign outputs[4559] = ~(layer2_outputs[12015]);
    assign outputs[4560] = (layer2_outputs[1219]) & ~(layer2_outputs[4148]);
    assign outputs[4561] = layer2_outputs[855];
    assign outputs[4562] = layer2_outputs[6890];
    assign outputs[4563] = ~((layer2_outputs[1354]) ^ (layer2_outputs[815]));
    assign outputs[4564] = (layer2_outputs[12445]) & ~(layer2_outputs[10771]);
    assign outputs[4565] = ~(layer2_outputs[1207]);
    assign outputs[4566] = ~(layer2_outputs[11568]);
    assign outputs[4567] = layer2_outputs[12365];
    assign outputs[4568] = ~((layer2_outputs[1759]) ^ (layer2_outputs[10608]));
    assign outputs[4569] = layer2_outputs[6177];
    assign outputs[4570] = layer2_outputs[7845];
    assign outputs[4571] = (layer2_outputs[8705]) ^ (layer2_outputs[2809]);
    assign outputs[4572] = ~(layer2_outputs[11087]);
    assign outputs[4573] = ~(layer2_outputs[7171]);
    assign outputs[4574] = ~(layer2_outputs[1935]);
    assign outputs[4575] = layer2_outputs[3448];
    assign outputs[4576] = ~((layer2_outputs[2377]) ^ (layer2_outputs[5900]));
    assign outputs[4577] = ~((layer2_outputs[8254]) ^ (layer2_outputs[747]));
    assign outputs[4578] = ~(layer2_outputs[2671]) | (layer2_outputs[1742]);
    assign outputs[4579] = layer2_outputs[7168];
    assign outputs[4580] = (layer2_outputs[4294]) ^ (layer2_outputs[9879]);
    assign outputs[4581] = ~(layer2_outputs[4450]) | (layer2_outputs[2811]);
    assign outputs[4582] = ~(layer2_outputs[9291]);
    assign outputs[4583] = ~((layer2_outputs[12034]) ^ (layer2_outputs[3495]));
    assign outputs[4584] = ~((layer2_outputs[7600]) & (layer2_outputs[5546]));
    assign outputs[4585] = ~(layer2_outputs[10876]);
    assign outputs[4586] = ~(layer2_outputs[12428]);
    assign outputs[4587] = ~(layer2_outputs[2076]);
    assign outputs[4588] = ~((layer2_outputs[9890]) ^ (layer2_outputs[1863]));
    assign outputs[4589] = ~(layer2_outputs[8992]);
    assign outputs[4590] = layer2_outputs[5184];
    assign outputs[4591] = (layer2_outputs[6777]) ^ (layer2_outputs[1142]);
    assign outputs[4592] = ~((layer2_outputs[9649]) | (layer2_outputs[9134]));
    assign outputs[4593] = (layer2_outputs[8411]) ^ (layer2_outputs[12494]);
    assign outputs[4594] = (layer2_outputs[4836]) & ~(layer2_outputs[6346]);
    assign outputs[4595] = layer2_outputs[9330];
    assign outputs[4596] = ~((layer2_outputs[10206]) ^ (layer2_outputs[4717]));
    assign outputs[4597] = (layer2_outputs[2280]) | (layer2_outputs[894]);
    assign outputs[4598] = (layer2_outputs[9922]) & (layer2_outputs[3221]);
    assign outputs[4599] = ~(layer2_outputs[2793]);
    assign outputs[4600] = (layer2_outputs[10119]) & ~(layer2_outputs[1668]);
    assign outputs[4601] = layer2_outputs[600];
    assign outputs[4602] = ~(layer2_outputs[8501]);
    assign outputs[4603] = (layer2_outputs[4733]) ^ (layer2_outputs[6222]);
    assign outputs[4604] = layer2_outputs[11978];
    assign outputs[4605] = (layer2_outputs[11237]) & ~(layer2_outputs[11062]);
    assign outputs[4606] = ~((layer2_outputs[1309]) ^ (layer2_outputs[4765]));
    assign outputs[4607] = layer2_outputs[4814];
    assign outputs[4608] = ~((layer2_outputs[2515]) ^ (layer2_outputs[6151]));
    assign outputs[4609] = layer2_outputs[5163];
    assign outputs[4610] = ~((layer2_outputs[5626]) ^ (layer2_outputs[9640]));
    assign outputs[4611] = ~(layer2_outputs[11568]);
    assign outputs[4612] = (layer2_outputs[4655]) & ~(layer2_outputs[3515]);
    assign outputs[4613] = ~(layer2_outputs[3583]);
    assign outputs[4614] = (layer2_outputs[9479]) ^ (layer2_outputs[11932]);
    assign outputs[4615] = layer2_outputs[6859];
    assign outputs[4616] = (layer2_outputs[2304]) ^ (layer2_outputs[5824]);
    assign outputs[4617] = layer2_outputs[8649];
    assign outputs[4618] = layer2_outputs[6945];
    assign outputs[4619] = ~((layer2_outputs[10395]) ^ (layer2_outputs[810]));
    assign outputs[4620] = (layer2_outputs[3663]) ^ (layer2_outputs[7028]);
    assign outputs[4621] = ~(layer2_outputs[5846]);
    assign outputs[4622] = ~((layer2_outputs[5950]) ^ (layer2_outputs[8201]));
    assign outputs[4623] = (layer2_outputs[2092]) & ~(layer2_outputs[3695]);
    assign outputs[4624] = layer2_outputs[495];
    assign outputs[4625] = (layer2_outputs[4217]) ^ (layer2_outputs[9192]);
    assign outputs[4626] = ~((layer2_outputs[11073]) ^ (layer2_outputs[4577]));
    assign outputs[4627] = layer2_outputs[7449];
    assign outputs[4628] = ~(layer2_outputs[4449]);
    assign outputs[4629] = (layer2_outputs[10357]) ^ (layer2_outputs[1182]);
    assign outputs[4630] = ~((layer2_outputs[6691]) ^ (layer2_outputs[1729]));
    assign outputs[4631] = layer2_outputs[4310];
    assign outputs[4632] = ~((layer2_outputs[8646]) ^ (layer2_outputs[756]));
    assign outputs[4633] = ~(layer2_outputs[1573]);
    assign outputs[4634] = ~(layer2_outputs[1251]) | (layer2_outputs[3293]);
    assign outputs[4635] = (layer2_outputs[6005]) & ~(layer2_outputs[11761]);
    assign outputs[4636] = ~((layer2_outputs[6922]) ^ (layer2_outputs[3271]));
    assign outputs[4637] = ~(layer2_outputs[2630]);
    assign outputs[4638] = ~(layer2_outputs[7923]);
    assign outputs[4639] = ~(layer2_outputs[4807]);
    assign outputs[4640] = layer2_outputs[4579];
    assign outputs[4641] = ~(layer2_outputs[7758]);
    assign outputs[4642] = ~(layer2_outputs[11529]);
    assign outputs[4643] = layer2_outputs[12229];
    assign outputs[4644] = ~(layer2_outputs[11574]);
    assign outputs[4645] = ~(layer2_outputs[2060]);
    assign outputs[4646] = (layer2_outputs[2756]) ^ (layer2_outputs[7949]);
    assign outputs[4647] = layer2_outputs[11449];
    assign outputs[4648] = layer2_outputs[9784];
    assign outputs[4649] = ~((layer2_outputs[4542]) | (layer2_outputs[10691]));
    assign outputs[4650] = ~((layer2_outputs[4210]) ^ (layer2_outputs[8414]));
    assign outputs[4651] = ~((layer2_outputs[4451]) | (layer2_outputs[4159]));
    assign outputs[4652] = ~(layer2_outputs[10135]) | (layer2_outputs[12732]);
    assign outputs[4653] = ~((layer2_outputs[7832]) ^ (layer2_outputs[11464]));
    assign outputs[4654] = ~(layer2_outputs[5795]);
    assign outputs[4655] = layer2_outputs[2233];
    assign outputs[4656] = layer2_outputs[8590];
    assign outputs[4657] = layer2_outputs[7623];
    assign outputs[4658] = ~(layer2_outputs[4200]);
    assign outputs[4659] = ~(layer2_outputs[1945]);
    assign outputs[4660] = ~((layer2_outputs[4475]) ^ (layer2_outputs[7854]));
    assign outputs[4661] = ~(layer2_outputs[12048]) | (layer2_outputs[9123]);
    assign outputs[4662] = layer2_outputs[6028];
    assign outputs[4663] = ~((layer2_outputs[11900]) ^ (layer2_outputs[7685]));
    assign outputs[4664] = layer2_outputs[9073];
    assign outputs[4665] = layer2_outputs[6733];
    assign outputs[4666] = ~(layer2_outputs[10314]);
    assign outputs[4667] = ~(layer2_outputs[9085]);
    assign outputs[4668] = ~((layer2_outputs[6230]) ^ (layer2_outputs[4999]));
    assign outputs[4669] = (layer2_outputs[5036]) ^ (layer2_outputs[3334]);
    assign outputs[4670] = (layer2_outputs[5564]) | (layer2_outputs[7033]);
    assign outputs[4671] = layer2_outputs[5372];
    assign outputs[4672] = ~(layer2_outputs[11707]);
    assign outputs[4673] = layer2_outputs[11297];
    assign outputs[4674] = ~((layer2_outputs[9348]) ^ (layer2_outputs[7175]));
    assign outputs[4675] = ~((layer2_outputs[10433]) ^ (layer2_outputs[11796]));
    assign outputs[4676] = ~(layer2_outputs[2074]);
    assign outputs[4677] = (layer2_outputs[12370]) ^ (layer2_outputs[11116]);
    assign outputs[4678] = (layer2_outputs[10539]) ^ (layer2_outputs[145]);
    assign outputs[4679] = ~(layer2_outputs[2436]) | (layer2_outputs[10561]);
    assign outputs[4680] = layer2_outputs[10004];
    assign outputs[4681] = ~((layer2_outputs[12780]) ^ (layer2_outputs[2307]));
    assign outputs[4682] = ~(layer2_outputs[2469]) | (layer2_outputs[10491]);
    assign outputs[4683] = layer2_outputs[4553];
    assign outputs[4684] = ~(layer2_outputs[9742]) | (layer2_outputs[3964]);
    assign outputs[4685] = (layer2_outputs[1034]) ^ (layer2_outputs[7107]);
    assign outputs[4686] = (layer2_outputs[2988]) & ~(layer2_outputs[6607]);
    assign outputs[4687] = ~(layer2_outputs[4830]);
    assign outputs[4688] = ~(layer2_outputs[7811]);
    assign outputs[4689] = ~(layer2_outputs[3069]) | (layer2_outputs[10888]);
    assign outputs[4690] = ~(layer2_outputs[8836]);
    assign outputs[4691] = (layer2_outputs[4500]) ^ (layer2_outputs[9391]);
    assign outputs[4692] = ~(layer2_outputs[2952]) | (layer2_outputs[4435]);
    assign outputs[4693] = ~(layer2_outputs[6357]) | (layer2_outputs[12635]);
    assign outputs[4694] = ~(layer2_outputs[3585]);
    assign outputs[4695] = ~(layer2_outputs[5490]);
    assign outputs[4696] = (layer2_outputs[1491]) ^ (layer2_outputs[11813]);
    assign outputs[4697] = ~(layer2_outputs[10947]);
    assign outputs[4698] = layer2_outputs[8330];
    assign outputs[4699] = ~(layer2_outputs[10528]);
    assign outputs[4700] = ~((layer2_outputs[1818]) ^ (layer2_outputs[4789]));
    assign outputs[4701] = ~((layer2_outputs[425]) ^ (layer2_outputs[11634]));
    assign outputs[4702] = (layer2_outputs[12646]) & ~(layer2_outputs[7621]);
    assign outputs[4703] = layer2_outputs[3483];
    assign outputs[4704] = ~(layer2_outputs[8011]);
    assign outputs[4705] = ~(layer2_outputs[3965]);
    assign outputs[4706] = layer2_outputs[4795];
    assign outputs[4707] = ~(layer2_outputs[2169]);
    assign outputs[4708] = layer2_outputs[10949];
    assign outputs[4709] = layer2_outputs[5222];
    assign outputs[4710] = layer2_outputs[10596];
    assign outputs[4711] = ~(layer2_outputs[5963]);
    assign outputs[4712] = layer2_outputs[4256];
    assign outputs[4713] = ~((layer2_outputs[3886]) ^ (layer2_outputs[9583]));
    assign outputs[4714] = layer2_outputs[6396];
    assign outputs[4715] = ~(layer2_outputs[10225]);
    assign outputs[4716] = layer2_outputs[1021];
    assign outputs[4717] = ~((layer2_outputs[7492]) ^ (layer2_outputs[9229]));
    assign outputs[4718] = ~(layer2_outputs[10644]);
    assign outputs[4719] = ~(layer2_outputs[1542]);
    assign outputs[4720] = ~(layer2_outputs[4948]);
    assign outputs[4721] = (layer2_outputs[188]) & ~(layer2_outputs[4023]);
    assign outputs[4722] = ~(layer2_outputs[9579]) | (layer2_outputs[3074]);
    assign outputs[4723] = layer2_outputs[9332];
    assign outputs[4724] = ~(layer2_outputs[11353]) | (layer2_outputs[3297]);
    assign outputs[4725] = ~(layer2_outputs[8257]);
    assign outputs[4726] = ~(layer2_outputs[5664]) | (layer2_outputs[4925]);
    assign outputs[4727] = (layer2_outputs[1958]) ^ (layer2_outputs[7378]);
    assign outputs[4728] = ~((layer2_outputs[11817]) ^ (layer2_outputs[1055]));
    assign outputs[4729] = (layer2_outputs[2724]) & ~(layer2_outputs[4433]);
    assign outputs[4730] = ~(layer2_outputs[4953]);
    assign outputs[4731] = (layer2_outputs[8677]) & (layer2_outputs[96]);
    assign outputs[4732] = ~(layer2_outputs[5594]);
    assign outputs[4733] = ~((layer2_outputs[540]) ^ (layer2_outputs[9461]));
    assign outputs[4734] = layer2_outputs[327];
    assign outputs[4735] = layer2_outputs[674];
    assign outputs[4736] = layer2_outputs[5557];
    assign outputs[4737] = ~(layer2_outputs[3854]);
    assign outputs[4738] = layer2_outputs[10753];
    assign outputs[4739] = ~(layer2_outputs[6061]);
    assign outputs[4740] = layer2_outputs[2786];
    assign outputs[4741] = layer2_outputs[12253];
    assign outputs[4742] = ~((layer2_outputs[6507]) ^ (layer2_outputs[7207]));
    assign outputs[4743] = layer2_outputs[1100];
    assign outputs[4744] = ~((layer2_outputs[7909]) ^ (layer2_outputs[11114]));
    assign outputs[4745] = ~(layer2_outputs[4198]) | (layer2_outputs[1478]);
    assign outputs[4746] = layer2_outputs[981];
    assign outputs[4747] = (layer2_outputs[3116]) ^ (layer2_outputs[4307]);
    assign outputs[4748] = ~(layer2_outputs[2618]);
    assign outputs[4749] = (layer2_outputs[1208]) ^ (layer2_outputs[722]);
    assign outputs[4750] = (layer2_outputs[8266]) ^ (layer2_outputs[3642]);
    assign outputs[4751] = (layer2_outputs[4038]) & ~(layer2_outputs[11100]);
    assign outputs[4752] = ~((layer2_outputs[4503]) ^ (layer2_outputs[1173]));
    assign outputs[4753] = ~(layer2_outputs[1151]) | (layer2_outputs[1960]);
    assign outputs[4754] = layer2_outputs[12786];
    assign outputs[4755] = layer2_outputs[12755];
    assign outputs[4756] = ~((layer2_outputs[9693]) ^ (layer2_outputs[10432]));
    assign outputs[4757] = ~(layer2_outputs[11975]);
    assign outputs[4758] = ~(layer2_outputs[7958]);
    assign outputs[4759] = layer2_outputs[1822];
    assign outputs[4760] = layer2_outputs[3434];
    assign outputs[4761] = (layer2_outputs[10906]) & ~(layer2_outputs[3087]);
    assign outputs[4762] = ~(layer2_outputs[5307]);
    assign outputs[4763] = ~(layer2_outputs[5838]);
    assign outputs[4764] = ~((layer2_outputs[9956]) ^ (layer2_outputs[557]));
    assign outputs[4765] = (layer2_outputs[5518]) & (layer2_outputs[11963]);
    assign outputs[4766] = layer2_outputs[3175];
    assign outputs[4767] = ~(layer2_outputs[3515]);
    assign outputs[4768] = ~(layer2_outputs[8056]);
    assign outputs[4769] = ~((layer2_outputs[12790]) & (layer2_outputs[473]));
    assign outputs[4770] = ~((layer2_outputs[8642]) ^ (layer2_outputs[7778]));
    assign outputs[4771] = layer2_outputs[2525];
    assign outputs[4772] = layer2_outputs[7633];
    assign outputs[4773] = (layer2_outputs[4279]) ^ (layer2_outputs[12359]);
    assign outputs[4774] = layer2_outputs[6914];
    assign outputs[4775] = ~((layer2_outputs[1371]) ^ (layer2_outputs[4735]));
    assign outputs[4776] = layer2_outputs[5707];
    assign outputs[4777] = layer2_outputs[8252];
    assign outputs[4778] = ~((layer2_outputs[4532]) ^ (layer2_outputs[8808]));
    assign outputs[4779] = ~(layer2_outputs[7381]);
    assign outputs[4780] = ~(layer2_outputs[8858]);
    assign outputs[4781] = layer2_outputs[8054];
    assign outputs[4782] = (layer2_outputs[10715]) & (layer2_outputs[6102]);
    assign outputs[4783] = ~(layer2_outputs[5380]);
    assign outputs[4784] = (layer2_outputs[11486]) & ~(layer2_outputs[5746]);
    assign outputs[4785] = (layer2_outputs[8161]) ^ (layer2_outputs[9230]);
    assign outputs[4786] = layer2_outputs[10326];
    assign outputs[4787] = layer2_outputs[9225];
    assign outputs[4788] = ~(layer2_outputs[12348]);
    assign outputs[4789] = layer2_outputs[4821];
    assign outputs[4790] = (layer2_outputs[5445]) ^ (layer2_outputs[1181]);
    assign outputs[4791] = ~(layer2_outputs[3854]);
    assign outputs[4792] = (layer2_outputs[4749]) & (layer2_outputs[10804]);
    assign outputs[4793] = ~(layer2_outputs[5192]);
    assign outputs[4794] = ~((layer2_outputs[12222]) & (layer2_outputs[7654]));
    assign outputs[4795] = ~((layer2_outputs[1647]) ^ (layer2_outputs[1755]));
    assign outputs[4796] = layer2_outputs[4205];
    assign outputs[4797] = ~(layer2_outputs[6051]);
    assign outputs[4798] = (layer2_outputs[10208]) ^ (layer2_outputs[3475]);
    assign outputs[4799] = layer2_outputs[10971];
    assign outputs[4800] = (layer2_outputs[9072]) ^ (layer2_outputs[162]);
    assign outputs[4801] = layer2_outputs[7873];
    assign outputs[4802] = layer2_outputs[12675];
    assign outputs[4803] = ~(layer2_outputs[6282]);
    assign outputs[4804] = layer2_outputs[11937];
    assign outputs[4805] = layer2_outputs[6329];
    assign outputs[4806] = ~((layer2_outputs[10834]) ^ (layer2_outputs[7264]));
    assign outputs[4807] = ~(layer2_outputs[7265]);
    assign outputs[4808] = layer2_outputs[5320];
    assign outputs[4809] = (layer2_outputs[11443]) ^ (layer2_outputs[11907]);
    assign outputs[4810] = (layer2_outputs[11468]) ^ (layer2_outputs[2908]);
    assign outputs[4811] = ~((layer2_outputs[12667]) ^ (layer2_outputs[11522]));
    assign outputs[4812] = (layer2_outputs[8118]) & (layer2_outputs[12220]);
    assign outputs[4813] = layer2_outputs[6182];
    assign outputs[4814] = layer2_outputs[10068];
    assign outputs[4815] = layer2_outputs[1886];
    assign outputs[4816] = (layer2_outputs[9921]) & ~(layer2_outputs[118]);
    assign outputs[4817] = ~(layer2_outputs[7279]);
    assign outputs[4818] = layer2_outputs[8463];
    assign outputs[4819] = (layer2_outputs[1557]) ^ (layer2_outputs[4756]);
    assign outputs[4820] = (layer2_outputs[9449]) ^ (layer2_outputs[9516]);
    assign outputs[4821] = ~((layer2_outputs[286]) | (layer2_outputs[6127]));
    assign outputs[4822] = ~(layer2_outputs[1436]);
    assign outputs[4823] = layer2_outputs[2451];
    assign outputs[4824] = (layer2_outputs[11843]) ^ (layer2_outputs[2925]);
    assign outputs[4825] = ~(layer2_outputs[11724]) | (layer2_outputs[2220]);
    assign outputs[4826] = layer2_outputs[5968];
    assign outputs[4827] = layer2_outputs[12679];
    assign outputs[4828] = ~(layer2_outputs[3327]);
    assign outputs[4829] = layer2_outputs[11756];
    assign outputs[4830] = ~(layer2_outputs[9381]);
    assign outputs[4831] = layer2_outputs[5412];
    assign outputs[4832] = ~(layer2_outputs[1857]);
    assign outputs[4833] = layer2_outputs[3157];
    assign outputs[4834] = layer2_outputs[5495];
    assign outputs[4835] = ~((layer2_outputs[7244]) | (layer2_outputs[7783]));
    assign outputs[4836] = (layer2_outputs[543]) & (layer2_outputs[5528]);
    assign outputs[4837] = ~((layer2_outputs[11895]) ^ (layer2_outputs[5788]));
    assign outputs[4838] = (layer2_outputs[5255]) | (layer2_outputs[2983]);
    assign outputs[4839] = layer2_outputs[4349];
    assign outputs[4840] = layer2_outputs[5924];
    assign outputs[4841] = layer2_outputs[2025];
    assign outputs[4842] = ~(layer2_outputs[2612]);
    assign outputs[4843] = ~((layer2_outputs[4118]) & (layer2_outputs[8581]));
    assign outputs[4844] = (layer2_outputs[2442]) & (layer2_outputs[2333]);
    assign outputs[4845] = ~((layer2_outputs[1985]) | (layer2_outputs[300]));
    assign outputs[4846] = ~(layer2_outputs[2071]);
    assign outputs[4847] = (layer2_outputs[9736]) ^ (layer2_outputs[4397]);
    assign outputs[4848] = (layer2_outputs[8416]) ^ (layer2_outputs[9471]);
    assign outputs[4849] = ~(layer2_outputs[11335]);
    assign outputs[4850] = ~((layer2_outputs[2863]) ^ (layer2_outputs[6112]));
    assign outputs[4851] = layer2_outputs[1617];
    assign outputs[4852] = ~(layer2_outputs[10154]);
    assign outputs[4853] = ~((layer2_outputs[11710]) & (layer2_outputs[2432]));
    assign outputs[4854] = layer2_outputs[8737];
    assign outputs[4855] = ~((layer2_outputs[5400]) ^ (layer2_outputs[10309]));
    assign outputs[4856] = layer2_outputs[5058];
    assign outputs[4857] = ~(layer2_outputs[9563]);
    assign outputs[4858] = (layer2_outputs[7697]) & (layer2_outputs[7420]);
    assign outputs[4859] = ~(layer2_outputs[8660]) | (layer2_outputs[4842]);
    assign outputs[4860] = (layer2_outputs[3273]) ^ (layer2_outputs[338]);
    assign outputs[4861] = ~(layer2_outputs[2088]);
    assign outputs[4862] = (layer2_outputs[9693]) | (layer2_outputs[7180]);
    assign outputs[4863] = (layer2_outputs[668]) ^ (layer2_outputs[10686]);
    assign outputs[4864] = layer2_outputs[2308];
    assign outputs[4865] = layer2_outputs[10751];
    assign outputs[4866] = ~((layer2_outputs[4203]) ^ (layer2_outputs[3944]));
    assign outputs[4867] = (layer2_outputs[11408]) | (layer2_outputs[11140]);
    assign outputs[4868] = layer2_outputs[11281];
    assign outputs[4869] = layer2_outputs[6682];
    assign outputs[4870] = ~(layer2_outputs[7737]);
    assign outputs[4871] = layer2_outputs[9643];
    assign outputs[4872] = ~(layer2_outputs[6638]);
    assign outputs[4873] = layer2_outputs[3768];
    assign outputs[4874] = ~(layer2_outputs[4177]);
    assign outputs[4875] = ~((layer2_outputs[4642]) ^ (layer2_outputs[841]));
    assign outputs[4876] = layer2_outputs[4586];
    assign outputs[4877] = ~(layer2_outputs[6640]);
    assign outputs[4878] = ~((layer2_outputs[9546]) ^ (layer2_outputs[7603]));
    assign outputs[4879] = (layer2_outputs[9465]) ^ (layer2_outputs[5287]);
    assign outputs[4880] = ~((layer2_outputs[10834]) & (layer2_outputs[10629]));
    assign outputs[4881] = ~(layer2_outputs[12439]) | (layer2_outputs[10004]);
    assign outputs[4882] = ~(layer2_outputs[8447]);
    assign outputs[4883] = (layer2_outputs[5801]) & ~(layer2_outputs[12257]);
    assign outputs[4884] = ~((layer2_outputs[5523]) ^ (layer2_outputs[7560]));
    assign outputs[4885] = ~(layer2_outputs[795]);
    assign outputs[4886] = (layer2_outputs[6741]) ^ (layer2_outputs[1119]);
    assign outputs[4887] = (layer2_outputs[7532]) | (layer2_outputs[4515]);
    assign outputs[4888] = ~(layer2_outputs[779]);
    assign outputs[4889] = ~(layer2_outputs[6463]);
    assign outputs[4890] = (layer2_outputs[9794]) & ~(layer2_outputs[11453]);
    assign outputs[4891] = layer2_outputs[11642];
    assign outputs[4892] = ~(layer2_outputs[5926]) | (layer2_outputs[10047]);
    assign outputs[4893] = ~(layer2_outputs[6065]);
    assign outputs[4894] = ~((layer2_outputs[8638]) ^ (layer2_outputs[7965]));
    assign outputs[4895] = ~(layer2_outputs[2387]);
    assign outputs[4896] = layer2_outputs[220];
    assign outputs[4897] = ~(layer2_outputs[6875]);
    assign outputs[4898] = layer2_outputs[6];
    assign outputs[4899] = (layer2_outputs[5821]) ^ (layer2_outputs[6998]);
    assign outputs[4900] = layer2_outputs[8280];
    assign outputs[4901] = layer2_outputs[5528];
    assign outputs[4902] = (layer2_outputs[5919]) ^ (layer2_outputs[12186]);
    assign outputs[4903] = layer2_outputs[9368];
    assign outputs[4904] = layer2_outputs[2978];
    assign outputs[4905] = ~(layer2_outputs[1089]);
    assign outputs[4906] = (layer2_outputs[5788]) ^ (layer2_outputs[3444]);
    assign outputs[4907] = ~((layer2_outputs[12517]) & (layer2_outputs[5180]));
    assign outputs[4908] = layer2_outputs[9884];
    assign outputs[4909] = layer2_outputs[4234];
    assign outputs[4910] = ~((layer2_outputs[2976]) ^ (layer2_outputs[6304]));
    assign outputs[4911] = layer2_outputs[1199];
    assign outputs[4912] = ~(layer2_outputs[12335]);
    assign outputs[4913] = (layer2_outputs[949]) | (layer2_outputs[4411]);
    assign outputs[4914] = (layer2_outputs[3064]) | (layer2_outputs[7495]);
    assign outputs[4915] = (layer2_outputs[5454]) & (layer2_outputs[5234]);
    assign outputs[4916] = ~(layer2_outputs[1460]);
    assign outputs[4917] = layer2_outputs[5197];
    assign outputs[4918] = ~((layer2_outputs[4675]) ^ (layer2_outputs[2593]));
    assign outputs[4919] = ~(layer2_outputs[5467]);
    assign outputs[4920] = (layer2_outputs[26]) ^ (layer2_outputs[1837]);
    assign outputs[4921] = (layer2_outputs[1032]) & (layer2_outputs[2692]);
    assign outputs[4922] = ~(layer2_outputs[9688]) | (layer2_outputs[10169]);
    assign outputs[4923] = (layer2_outputs[4282]) ^ (layer2_outputs[7042]);
    assign outputs[4924] = (layer2_outputs[2374]) & ~(layer2_outputs[12402]);
    assign outputs[4925] = ~((layer2_outputs[12573]) ^ (layer2_outputs[10017]));
    assign outputs[4926] = ~(layer2_outputs[11646]);
    assign outputs[4927] = (layer2_outputs[2602]) & ~(layer2_outputs[2665]);
    assign outputs[4928] = ~(layer2_outputs[5204]);
    assign outputs[4929] = layer2_outputs[4626];
    assign outputs[4930] = layer2_outputs[9631];
    assign outputs[4931] = (layer2_outputs[11413]) & (layer2_outputs[1283]);
    assign outputs[4932] = (layer2_outputs[66]) & ~(layer2_outputs[9567]);
    assign outputs[4933] = (layer2_outputs[8675]) ^ (layer2_outputs[7268]);
    assign outputs[4934] = layer2_outputs[5125];
    assign outputs[4935] = ~(layer2_outputs[8706]);
    assign outputs[4936] = (layer2_outputs[1267]) ^ (layer2_outputs[816]);
    assign outputs[4937] = layer2_outputs[11881];
    assign outputs[4938] = ~(layer2_outputs[651]) | (layer2_outputs[2]);
    assign outputs[4939] = ~(layer2_outputs[8807]);
    assign outputs[4940] = (layer2_outputs[4218]) ^ (layer2_outputs[2528]);
    assign outputs[4941] = (layer2_outputs[432]) ^ (layer2_outputs[4978]);
    assign outputs[4942] = ~((layer2_outputs[1819]) ^ (layer2_outputs[6889]));
    assign outputs[4943] = ~((layer2_outputs[12779]) ^ (layer2_outputs[10781]));
    assign outputs[4944] = layer2_outputs[11324];
    assign outputs[4945] = ~(layer2_outputs[11346]);
    assign outputs[4946] = layer2_outputs[9139];
    assign outputs[4947] = layer2_outputs[12756];
    assign outputs[4948] = layer2_outputs[4057];
    assign outputs[4949] = (layer2_outputs[5636]) ^ (layer2_outputs[1704]);
    assign outputs[4950] = layer2_outputs[10649];
    assign outputs[4951] = ~((layer2_outputs[7072]) & (layer2_outputs[7576]));
    assign outputs[4952] = ~(layer2_outputs[6901]);
    assign outputs[4953] = ~(layer2_outputs[3687]);
    assign outputs[4954] = ~(layer2_outputs[3720]);
    assign outputs[4955] = layer2_outputs[430];
    assign outputs[4956] = layer2_outputs[6217];
    assign outputs[4957] = (layer2_outputs[5346]) ^ (layer2_outputs[12057]);
    assign outputs[4958] = ~((layer2_outputs[11076]) & (layer2_outputs[9462]));
    assign outputs[4959] = (layer2_outputs[4672]) & ~(layer2_outputs[3733]);
    assign outputs[4960] = (layer2_outputs[8952]) ^ (layer2_outputs[10892]);
    assign outputs[4961] = ~(layer2_outputs[12290]);
    assign outputs[4962] = (layer2_outputs[3035]) & ~(layer2_outputs[7726]);
    assign outputs[4963] = (layer2_outputs[2052]) & ~(layer2_outputs[6670]);
    assign outputs[4964] = ~(layer2_outputs[1245]);
    assign outputs[4965] = ~((layer2_outputs[7414]) ^ (layer2_outputs[10945]));
    assign outputs[4966] = ~(layer2_outputs[7102]);
    assign outputs[4967] = ~(layer2_outputs[2989]);
    assign outputs[4968] = ~(layer2_outputs[8226]);
    assign outputs[4969] = (layer2_outputs[8019]) ^ (layer2_outputs[551]);
    assign outputs[4970] = ~(layer2_outputs[421]);
    assign outputs[4971] = ~(layer2_outputs[8986]) | (layer2_outputs[5663]);
    assign outputs[4972] = layer2_outputs[1333];
    assign outputs[4973] = ~((layer2_outputs[7759]) | (layer2_outputs[6071]));
    assign outputs[4974] = ~(layer2_outputs[11562]);
    assign outputs[4975] = (layer2_outputs[1387]) & ~(layer2_outputs[12628]);
    assign outputs[4976] = (layer2_outputs[4845]) & ~(layer2_outputs[407]);
    assign outputs[4977] = layer2_outputs[5338];
    assign outputs[4978] = layer2_outputs[6423];
    assign outputs[4979] = (layer2_outputs[5134]) & (layer2_outputs[7487]);
    assign outputs[4980] = ~(layer2_outputs[10716]);
    assign outputs[4981] = layer2_outputs[792];
    assign outputs[4982] = ~((layer2_outputs[7826]) ^ (layer2_outputs[2347]));
    assign outputs[4983] = layer2_outputs[4027];
    assign outputs[4984] = ~((layer2_outputs[772]) | (layer2_outputs[10513]));
    assign outputs[4985] = ~((layer2_outputs[359]) | (layer2_outputs[6224]));
    assign outputs[4986] = (layer2_outputs[5943]) ^ (layer2_outputs[12543]);
    assign outputs[4987] = ~(layer2_outputs[7509]);
    assign outputs[4988] = layer2_outputs[3367];
    assign outputs[4989] = layer2_outputs[11971];
    assign outputs[4990] = ~(layer2_outputs[268]) | (layer2_outputs[9021]);
    assign outputs[4991] = ~(layer2_outputs[9376]);
    assign outputs[4992] = layer2_outputs[8810];
    assign outputs[4993] = ~(layer2_outputs[3802]);
    assign outputs[4994] = layer2_outputs[2980];
    assign outputs[4995] = layer2_outputs[5506];
    assign outputs[4996] = layer2_outputs[2544];
    assign outputs[4997] = layer2_outputs[3440];
    assign outputs[4998] = ~((layer2_outputs[10497]) ^ (layer2_outputs[199]));
    assign outputs[4999] = ~(layer2_outputs[3453]);
    assign outputs[5000] = (layer2_outputs[1236]) & ~(layer2_outputs[11550]);
    assign outputs[5001] = layer2_outputs[3132];
    assign outputs[5002] = ~((layer2_outputs[12761]) | (layer2_outputs[7256]));
    assign outputs[5003] = (layer2_outputs[149]) ^ (layer2_outputs[2311]);
    assign outputs[5004] = ~(layer2_outputs[9697]) | (layer2_outputs[12720]);
    assign outputs[5005] = layer2_outputs[8417];
    assign outputs[5006] = layer2_outputs[3017];
    assign outputs[5007] = layer2_outputs[4150];
    assign outputs[5008] = layer2_outputs[12273];
    assign outputs[5009] = (layer2_outputs[201]) ^ (layer2_outputs[5746]);
    assign outputs[5010] = ~((layer2_outputs[9772]) ^ (layer2_outputs[5908]));
    assign outputs[5011] = (layer2_outputs[4480]) ^ (layer2_outputs[8288]);
    assign outputs[5012] = layer2_outputs[6104];
    assign outputs[5013] = layer2_outputs[10382];
    assign outputs[5014] = ~((layer2_outputs[857]) ^ (layer2_outputs[10235]));
    assign outputs[5015] = ~(layer2_outputs[905]);
    assign outputs[5016] = ~(layer2_outputs[6082]);
    assign outputs[5017] = (layer2_outputs[10623]) & ~(layer2_outputs[5204]);
    assign outputs[5018] = ~(layer2_outputs[727]);
    assign outputs[5019] = (layer2_outputs[1677]) ^ (layer2_outputs[5427]);
    assign outputs[5020] = (layer2_outputs[7548]) & ~(layer2_outputs[5516]);
    assign outputs[5021] = (layer2_outputs[7277]) ^ (layer2_outputs[3540]);
    assign outputs[5022] = (layer2_outputs[265]) & (layer2_outputs[3391]);
    assign outputs[5023] = layer2_outputs[5584];
    assign outputs[5024] = ~(layer2_outputs[3792]);
    assign outputs[5025] = ~((layer2_outputs[12164]) | (layer2_outputs[881]));
    assign outputs[5026] = (layer2_outputs[11051]) ^ (layer2_outputs[455]);
    assign outputs[5027] = layer2_outputs[1250];
    assign outputs[5028] = ~(layer2_outputs[9489]);
    assign outputs[5029] = ~(layer2_outputs[2083]);
    assign outputs[5030] = (layer2_outputs[9040]) ^ (layer2_outputs[8378]);
    assign outputs[5031] = (layer2_outputs[11522]) ^ (layer2_outputs[2234]);
    assign outputs[5032] = (layer2_outputs[254]) ^ (layer2_outputs[7510]);
    assign outputs[5033] = layer2_outputs[10646];
    assign outputs[5034] = layer2_outputs[9239];
    assign outputs[5035] = layer2_outputs[1480];
    assign outputs[5036] = (layer2_outputs[6385]) & ~(layer2_outputs[5096]);
    assign outputs[5037] = ~(layer2_outputs[12233]);
    assign outputs[5038] = layer2_outputs[612];
    assign outputs[5039] = layer2_outputs[12268];
    assign outputs[5040] = (layer2_outputs[4014]) ^ (layer2_outputs[7972]);
    assign outputs[5041] = layer2_outputs[8507];
    assign outputs[5042] = (layer2_outputs[7407]) & ~(layer2_outputs[5470]);
    assign outputs[5043] = layer2_outputs[10983];
    assign outputs[5044] = (layer2_outputs[12298]) ^ (layer2_outputs[7498]);
    assign outputs[5045] = ~(layer2_outputs[1876]);
    assign outputs[5046] = (layer2_outputs[7766]) & ~(layer2_outputs[7280]);
    assign outputs[5047] = ~((layer2_outputs[5022]) ^ (layer2_outputs[3698]));
    assign outputs[5048] = ~(layer2_outputs[7385]);
    assign outputs[5049] = layer2_outputs[5596];
    assign outputs[5050] = ~(layer2_outputs[1901]);
    assign outputs[5051] = layer2_outputs[12053];
    assign outputs[5052] = layer2_outputs[7402];
    assign outputs[5053] = (layer2_outputs[11985]) | (layer2_outputs[3710]);
    assign outputs[5054] = ~(layer2_outputs[9096]);
    assign outputs[5055] = ~((layer2_outputs[7152]) ^ (layer2_outputs[9888]));
    assign outputs[5056] = ~(layer2_outputs[10534]);
    assign outputs[5057] = ~((layer2_outputs[9082]) | (layer2_outputs[2909]));
    assign outputs[5058] = layer2_outputs[8810];
    assign outputs[5059] = layer2_outputs[4079];
    assign outputs[5060] = layer2_outputs[10253];
    assign outputs[5061] = layer2_outputs[10447];
    assign outputs[5062] = (layer2_outputs[9813]) ^ (layer2_outputs[1166]);
    assign outputs[5063] = ~((layer2_outputs[12340]) | (layer2_outputs[6512]));
    assign outputs[5064] = layer2_outputs[9855];
    assign outputs[5065] = ~(layer2_outputs[8332]);
    assign outputs[5066] = layer2_outputs[10745];
    assign outputs[5067] = layer2_outputs[2984];
    assign outputs[5068] = layer2_outputs[8398];
    assign outputs[5069] = layer2_outputs[6336];
    assign outputs[5070] = layer2_outputs[10714];
    assign outputs[5071] = ~(layer2_outputs[12080]);
    assign outputs[5072] = layer2_outputs[4602];
    assign outputs[5073] = ~(layer2_outputs[9090]);
    assign outputs[5074] = ~(layer2_outputs[5430]);
    assign outputs[5075] = ~((layer2_outputs[7772]) ^ (layer2_outputs[1529]));
    assign outputs[5076] = layer2_outputs[10340];
    assign outputs[5077] = ~(layer2_outputs[12309]);
    assign outputs[5078] = (layer2_outputs[12019]) ^ (layer2_outputs[3612]);
    assign outputs[5079] = layer2_outputs[10199];
    assign outputs[5080] = (layer2_outputs[7031]) & (layer2_outputs[2649]);
    assign outputs[5081] = ~(layer2_outputs[250]);
    assign outputs[5082] = ~(layer2_outputs[9136]);
    assign outputs[5083] = (layer2_outputs[8642]) & (layer2_outputs[7352]);
    assign outputs[5084] = layer2_outputs[201];
    assign outputs[5085] = (layer2_outputs[2149]) ^ (layer2_outputs[2591]);
    assign outputs[5086] = ~((layer2_outputs[3155]) ^ (layer2_outputs[5241]));
    assign outputs[5087] = ~(layer2_outputs[579]);
    assign outputs[5088] = (layer2_outputs[11316]) & ~(layer2_outputs[5896]);
    assign outputs[5089] = ~((layer2_outputs[3682]) ^ (layer2_outputs[7779]));
    assign outputs[5090] = ~(layer2_outputs[9307]);
    assign outputs[5091] = (layer2_outputs[11983]) ^ (layer2_outputs[11273]);
    assign outputs[5092] = ~(layer2_outputs[12346]);
    assign outputs[5093] = layer2_outputs[11666];
    assign outputs[5094] = ~(layer2_outputs[8163]);
    assign outputs[5095] = (layer2_outputs[2133]) & ~(layer2_outputs[8662]);
    assign outputs[5096] = ~((layer2_outputs[8174]) ^ (layer2_outputs[11980]));
    assign outputs[5097] = (layer2_outputs[2087]) & ~(layer2_outputs[9781]);
    assign outputs[5098] = ~(layer2_outputs[9217]);
    assign outputs[5099] = layer2_outputs[1713];
    assign outputs[5100] = ~(layer2_outputs[11967]) | (layer2_outputs[7790]);
    assign outputs[5101] = ~(layer2_outputs[3488]);
    assign outputs[5102] = layer2_outputs[7160];
    assign outputs[5103] = (layer2_outputs[3433]) ^ (layer2_outputs[1159]);
    assign outputs[5104] = layer2_outputs[6328];
    assign outputs[5105] = (layer2_outputs[7081]) ^ (layer2_outputs[7835]);
    assign outputs[5106] = ~(layer2_outputs[9035]);
    assign outputs[5107] = ~(layer2_outputs[10091]);
    assign outputs[5108] = ~((layer2_outputs[12360]) ^ (layer2_outputs[8892]));
    assign outputs[5109] = layer2_outputs[4828];
    assign outputs[5110] = ~((layer2_outputs[10057]) ^ (layer2_outputs[6851]));
    assign outputs[5111] = ~(layer2_outputs[2664]);
    assign outputs[5112] = ~(layer2_outputs[11773]);
    assign outputs[5113] = layer2_outputs[7009];
    assign outputs[5114] = layer2_outputs[5831];
    assign outputs[5115] = ~(layer2_outputs[6616]);
    assign outputs[5116] = layer2_outputs[12723];
    assign outputs[5117] = ~(layer2_outputs[204]);
    assign outputs[5118] = ~(layer2_outputs[3134]);
    assign outputs[5119] = (layer2_outputs[6508]) ^ (layer2_outputs[8545]);
    assign outputs[5120] = ~((layer2_outputs[12238]) | (layer2_outputs[8886]));
    assign outputs[5121] = (layer2_outputs[6668]) ^ (layer2_outputs[7295]);
    assign outputs[5122] = layer2_outputs[4767];
    assign outputs[5123] = layer2_outputs[3229];
    assign outputs[5124] = ~(layer2_outputs[10517]);
    assign outputs[5125] = layer2_outputs[10225];
    assign outputs[5126] = layer2_outputs[1033];
    assign outputs[5127] = ~(layer2_outputs[261]);
    assign outputs[5128] = ~(layer2_outputs[5061]);
    assign outputs[5129] = ~(layer2_outputs[3113]);
    assign outputs[5130] = ~((layer2_outputs[4152]) ^ (layer2_outputs[3958]));
    assign outputs[5131] = (layer2_outputs[8924]) | (layer2_outputs[1072]);
    assign outputs[5132] = (layer2_outputs[10943]) ^ (layer2_outputs[6265]);
    assign outputs[5133] = ~(layer2_outputs[1368]);
    assign outputs[5134] = (layer2_outputs[6276]) ^ (layer2_outputs[6520]);
    assign outputs[5135] = layer2_outputs[9749];
    assign outputs[5136] = ~(layer2_outputs[9149]) | (layer2_outputs[6490]);
    assign outputs[5137] = (layer2_outputs[8058]) ^ (layer2_outputs[3933]);
    assign outputs[5138] = ~((layer2_outputs[9377]) ^ (layer2_outputs[648]));
    assign outputs[5139] = layer2_outputs[1750];
    assign outputs[5140] = (layer2_outputs[3342]) ^ (layer2_outputs[7097]);
    assign outputs[5141] = (layer2_outputs[5922]) ^ (layer2_outputs[11401]);
    assign outputs[5142] = layer2_outputs[8633];
    assign outputs[5143] = ~((layer2_outputs[12531]) ^ (layer2_outputs[4188]));
    assign outputs[5144] = (layer2_outputs[6032]) & (layer2_outputs[11190]);
    assign outputs[5145] = (layer2_outputs[11511]) & ~(layer2_outputs[11633]);
    assign outputs[5146] = layer2_outputs[12609];
    assign outputs[5147] = layer2_outputs[6038];
    assign outputs[5148] = (layer2_outputs[3546]) ^ (layer2_outputs[3361]);
    assign outputs[5149] = ~((layer2_outputs[694]) | (layer2_outputs[12269]));
    assign outputs[5150] = ~((layer2_outputs[4588]) ^ (layer2_outputs[819]));
    assign outputs[5151] = (layer2_outputs[3228]) ^ (layer2_outputs[3624]);
    assign outputs[5152] = (layer2_outputs[12767]) ^ (layer2_outputs[7320]);
    assign outputs[5153] = (layer2_outputs[11044]) ^ (layer2_outputs[5044]);
    assign outputs[5154] = ~(layer2_outputs[5890]);
    assign outputs[5155] = ~(layer2_outputs[5699]) | (layer2_outputs[12765]);
    assign outputs[5156] = (layer2_outputs[11171]) ^ (layer2_outputs[5093]);
    assign outputs[5157] = (layer2_outputs[5649]) ^ (layer2_outputs[7640]);
    assign outputs[5158] = layer2_outputs[10855];
    assign outputs[5159] = ~((layer2_outputs[11201]) | (layer2_outputs[8312]));
    assign outputs[5160] = ~(layer2_outputs[850]);
    assign outputs[5161] = (layer2_outputs[10505]) ^ (layer2_outputs[2624]);
    assign outputs[5162] = (layer2_outputs[12749]) ^ (layer2_outputs[3829]);
    assign outputs[5163] = ~(layer2_outputs[8453]) | (layer2_outputs[8361]);
    assign outputs[5164] = ~(layer2_outputs[5440]);
    assign outputs[5165] = (layer2_outputs[1196]) ^ (layer2_outputs[3573]);
    assign outputs[5166] = ~((layer2_outputs[5081]) & (layer2_outputs[7046]));
    assign outputs[5167] = ~(layer2_outputs[517]);
    assign outputs[5168] = ~((layer2_outputs[7702]) | (layer2_outputs[4884]));
    assign outputs[5169] = ~(layer2_outputs[4953]);
    assign outputs[5170] = layer2_outputs[474];
    assign outputs[5171] = (layer2_outputs[8573]) ^ (layer2_outputs[5194]);
    assign outputs[5172] = (layer2_outputs[5001]) ^ (layer2_outputs[6592]);
    assign outputs[5173] = ~(layer2_outputs[10477]);
    assign outputs[5174] = ~(layer2_outputs[2138]);
    assign outputs[5175] = ~((layer2_outputs[10833]) | (layer2_outputs[7695]));
    assign outputs[5176] = layer2_outputs[10812];
    assign outputs[5177] = ~(layer2_outputs[7019]);
    assign outputs[5178] = ~(layer2_outputs[6912]);
    assign outputs[5179] = ~(layer2_outputs[7724]);
    assign outputs[5180] = layer2_outputs[5451];
    assign outputs[5181] = layer2_outputs[2258];
    assign outputs[5182] = (layer2_outputs[11211]) ^ (layer2_outputs[5796]);
    assign outputs[5183] = (layer2_outputs[6936]) ^ (layer2_outputs[10042]);
    assign outputs[5184] = layer2_outputs[10993];
    assign outputs[5185] = ~((layer2_outputs[9441]) ^ (layer2_outputs[6031]));
    assign outputs[5186] = ~(layer2_outputs[3864]);
    assign outputs[5187] = (layer2_outputs[11696]) ^ (layer2_outputs[3233]);
    assign outputs[5188] = layer2_outputs[12753];
    assign outputs[5189] = ~(layer2_outputs[3716]);
    assign outputs[5190] = layer2_outputs[6995];
    assign outputs[5191] = (layer2_outputs[8619]) & (layer2_outputs[12598]);
    assign outputs[5192] = layer2_outputs[7701];
    assign outputs[5193] = ~(layer2_outputs[5156]);
    assign outputs[5194] = layer2_outputs[10022];
    assign outputs[5195] = (layer2_outputs[3613]) ^ (layer2_outputs[1961]);
    assign outputs[5196] = (layer2_outputs[5334]) ^ (layer2_outputs[7592]);
    assign outputs[5197] = (layer2_outputs[757]) ^ (layer2_outputs[2098]);
    assign outputs[5198] = ~(layer2_outputs[4575]);
    assign outputs[5199] = ~(layer2_outputs[5291]);
    assign outputs[5200] = ~(layer2_outputs[1516]);
    assign outputs[5201] = ~(layer2_outputs[510]);
    assign outputs[5202] = ~(layer2_outputs[8419]);
    assign outputs[5203] = layer2_outputs[5778];
    assign outputs[5204] = layer2_outputs[8943];
    assign outputs[5205] = ~(layer2_outputs[7568]);
    assign outputs[5206] = (layer2_outputs[12544]) ^ (layer2_outputs[10274]);
    assign outputs[5207] = ~(layer2_outputs[52]);
    assign outputs[5208] = ~(layer2_outputs[602]) | (layer2_outputs[9686]);
    assign outputs[5209] = ~(layer2_outputs[7137]);
    assign outputs[5210] = ~(layer2_outputs[3754]);
    assign outputs[5211] = layer2_outputs[9101];
    assign outputs[5212] = ~(layer2_outputs[6447]);
    assign outputs[5213] = ~(layer2_outputs[12038]);
    assign outputs[5214] = ~((layer2_outputs[7246]) ^ (layer2_outputs[3908]));
    assign outputs[5215] = layer2_outputs[12454];
    assign outputs[5216] = ~((layer2_outputs[5330]) ^ (layer2_outputs[1380]));
    assign outputs[5217] = ~(layer2_outputs[8173]) | (layer2_outputs[9456]);
    assign outputs[5218] = (layer2_outputs[5925]) ^ (layer2_outputs[10598]);
    assign outputs[5219] = ~(layer2_outputs[2702]);
    assign outputs[5220] = ~(layer2_outputs[378]);
    assign outputs[5221] = layer2_outputs[946];
    assign outputs[5222] = (layer2_outputs[7425]) | (layer2_outputs[10174]);
    assign outputs[5223] = ~((layer2_outputs[7232]) ^ (layer2_outputs[4271]));
    assign outputs[5224] = layer2_outputs[3838];
    assign outputs[5225] = layer2_outputs[8326];
    assign outputs[5226] = ~((layer2_outputs[11200]) ^ (layer2_outputs[8546]));
    assign outputs[5227] = ~((layer2_outputs[1914]) ^ (layer2_outputs[8304]));
    assign outputs[5228] = layer2_outputs[7650];
    assign outputs[5229] = ~(layer2_outputs[4172]);
    assign outputs[5230] = layer2_outputs[12652];
    assign outputs[5231] = layer2_outputs[7408];
    assign outputs[5232] = ~(layer2_outputs[12650]);
    assign outputs[5233] = ~(layer2_outputs[3006]);
    assign outputs[5234] = ~((layer2_outputs[8466]) & (layer2_outputs[1062]));
    assign outputs[5235] = (layer2_outputs[7]) & ~(layer2_outputs[10169]);
    assign outputs[5236] = (layer2_outputs[10721]) & ~(layer2_outputs[319]);
    assign outputs[5237] = ~((layer2_outputs[1019]) & (layer2_outputs[997]));
    assign outputs[5238] = layer2_outputs[7249];
    assign outputs[5239] = ~((layer2_outputs[8015]) ^ (layer2_outputs[6089]));
    assign outputs[5240] = ~((layer2_outputs[1554]) ^ (layer2_outputs[8883]));
    assign outputs[5241] = layer2_outputs[7957];
    assign outputs[5242] = ~(layer2_outputs[3861]);
    assign outputs[5243] = ~(layer2_outputs[8920]) | (layer2_outputs[661]);
    assign outputs[5244] = layer2_outputs[3690];
    assign outputs[5245] = ~(layer2_outputs[4736]) | (layer2_outputs[3659]);
    assign outputs[5246] = ~(layer2_outputs[10747]);
    assign outputs[5247] = layer2_outputs[7922];
    assign outputs[5248] = ~(layer2_outputs[1967]);
    assign outputs[5249] = ~(layer2_outputs[8129]) | (layer2_outputs[7237]);
    assign outputs[5250] = (layer2_outputs[1633]) & (layer2_outputs[12459]);
    assign outputs[5251] = layer2_outputs[2499];
    assign outputs[5252] = layer2_outputs[7927];
    assign outputs[5253] = ~(layer2_outputs[10746]);
    assign outputs[5254] = ~(layer2_outputs[12440]) | (layer2_outputs[6728]);
    assign outputs[5255] = layer2_outputs[2398];
    assign outputs[5256] = ~((layer2_outputs[4025]) & (layer2_outputs[8467]));
    assign outputs[5257] = layer2_outputs[116];
    assign outputs[5258] = layer2_outputs[12235];
    assign outputs[5259] = ~(layer2_outputs[2473]) | (layer2_outputs[7370]);
    assign outputs[5260] = (layer2_outputs[10122]) | (layer2_outputs[5923]);
    assign outputs[5261] = layer2_outputs[2721];
    assign outputs[5262] = ~(layer2_outputs[9719]);
    assign outputs[5263] = ~(layer2_outputs[8769]);
    assign outputs[5264] = ~(layer2_outputs[11078]);
    assign outputs[5265] = layer2_outputs[9314];
    assign outputs[5266] = ~(layer2_outputs[11223]) | (layer2_outputs[724]);
    assign outputs[5267] = layer2_outputs[7409];
    assign outputs[5268] = ~(layer2_outputs[9016]);
    assign outputs[5269] = ~((layer2_outputs[101]) ^ (layer2_outputs[5058]));
    assign outputs[5270] = (layer2_outputs[8516]) & (layer2_outputs[325]);
    assign outputs[5271] = ~(layer2_outputs[6342]);
    assign outputs[5272] = ~((layer2_outputs[12400]) ^ (layer2_outputs[1495]));
    assign outputs[5273] = layer2_outputs[376];
    assign outputs[5274] = (layer2_outputs[4652]) ^ (layer2_outputs[11584]);
    assign outputs[5275] = ~(layer2_outputs[10312]) | (layer2_outputs[1785]);
    assign outputs[5276] = layer2_outputs[9545];
    assign outputs[5277] = ~(layer2_outputs[4342]);
    assign outputs[5278] = (layer2_outputs[4659]) | (layer2_outputs[10922]);
    assign outputs[5279] = ~(layer2_outputs[7683]) | (layer2_outputs[8913]);
    assign outputs[5280] = ~(layer2_outputs[9172]);
    assign outputs[5281] = (layer2_outputs[183]) ^ (layer2_outputs[3179]);
    assign outputs[5282] = ~(layer2_outputs[7638]);
    assign outputs[5283] = ~((layer2_outputs[4557]) ^ (layer2_outputs[8288]));
    assign outputs[5284] = (layer2_outputs[6384]) ^ (layer2_outputs[5931]);
    assign outputs[5285] = layer2_outputs[5764];
    assign outputs[5286] = (layer2_outputs[6703]) & (layer2_outputs[7087]);
    assign outputs[5287] = ~(layer2_outputs[8453]);
    assign outputs[5288] = (layer2_outputs[4470]) ^ (layer2_outputs[6873]);
    assign outputs[5289] = ~((layer2_outputs[7751]) ^ (layer2_outputs[232]));
    assign outputs[5290] = layer2_outputs[8439];
    assign outputs[5291] = ~(layer2_outputs[6294]);
    assign outputs[5292] = ~((layer2_outputs[2957]) ^ (layer2_outputs[3215]));
    assign outputs[5293] = layer2_outputs[11130];
    assign outputs[5294] = (layer2_outputs[11065]) ^ (layer2_outputs[6225]);
    assign outputs[5295] = ~(layer2_outputs[12752]);
    assign outputs[5296] = ~(layer2_outputs[5008]);
    assign outputs[5297] = ~(layer2_outputs[8813]);
    assign outputs[5298] = ~(layer2_outputs[283]);
    assign outputs[5299] = ~(layer2_outputs[7063]);
    assign outputs[5300] = ~(layer2_outputs[3835]);
    assign outputs[5301] = ~((layer2_outputs[8151]) ^ (layer2_outputs[5760]));
    assign outputs[5302] = ~(layer2_outputs[3077]);
    assign outputs[5303] = layer2_outputs[10062];
    assign outputs[5304] = layer2_outputs[1273];
    assign outputs[5305] = (layer2_outputs[11012]) | (layer2_outputs[5068]);
    assign outputs[5306] = ~((layer2_outputs[8035]) ^ (layer2_outputs[1315]));
    assign outputs[5307] = (layer2_outputs[11856]) ^ (layer2_outputs[4924]);
    assign outputs[5308] = layer2_outputs[2290];
    assign outputs[5309] = layer2_outputs[2664];
    assign outputs[5310] = layer2_outputs[3653];
    assign outputs[5311] = ~((layer2_outputs[6425]) ^ (layer2_outputs[7894]));
    assign outputs[5312] = (layer2_outputs[1942]) & ~(layer2_outputs[2143]);
    assign outputs[5313] = (layer2_outputs[11004]) ^ (layer2_outputs[9313]);
    assign outputs[5314] = (layer2_outputs[4567]) & (layer2_outputs[11147]);
    assign outputs[5315] = ~((layer2_outputs[1493]) | (layer2_outputs[548]));
    assign outputs[5316] = layer2_outputs[10422];
    assign outputs[5317] = layer2_outputs[11175];
    assign outputs[5318] = layer2_outputs[4090];
    assign outputs[5319] = ~(layer2_outputs[8520]);
    assign outputs[5320] = layer2_outputs[718];
    assign outputs[5321] = (layer2_outputs[8611]) & ~(layer2_outputs[3840]);
    assign outputs[5322] = (layer2_outputs[10819]) ^ (layer2_outputs[9965]);
    assign outputs[5323] = ~(layer2_outputs[9696]);
    assign outputs[5324] = (layer2_outputs[4565]) ^ (layer2_outputs[3571]);
    assign outputs[5325] = layer2_outputs[9627];
    assign outputs[5326] = layer2_outputs[10978];
    assign outputs[5327] = ~(layer2_outputs[11547]);
    assign outputs[5328] = layer2_outputs[8634];
    assign outputs[5329] = (layer2_outputs[6338]) ^ (layer2_outputs[561]);
    assign outputs[5330] = ~(layer2_outputs[4104]);
    assign outputs[5331] = ~(layer2_outputs[645]);
    assign outputs[5332] = (layer2_outputs[1404]) ^ (layer2_outputs[1620]);
    assign outputs[5333] = ~((layer2_outputs[227]) ^ (layer2_outputs[8825]));
    assign outputs[5334] = (layer2_outputs[11414]) | (layer2_outputs[1334]);
    assign outputs[5335] = layer2_outputs[4897];
    assign outputs[5336] = layer2_outputs[9629];
    assign outputs[5337] = (layer2_outputs[5598]) & (layer2_outputs[7243]);
    assign outputs[5338] = layer2_outputs[10484];
    assign outputs[5339] = (layer2_outputs[7756]) ^ (layer2_outputs[1328]);
    assign outputs[5340] = ~(layer2_outputs[10081]);
    assign outputs[5341] = (layer2_outputs[8632]) ^ (layer2_outputs[2202]);
    assign outputs[5342] = layer2_outputs[5187];
    assign outputs[5343] = ~((layer2_outputs[2927]) ^ (layer2_outputs[9345]));
    assign outputs[5344] = ~((layer2_outputs[8002]) | (layer2_outputs[2712]));
    assign outputs[5345] = (layer2_outputs[3650]) & ~(layer2_outputs[8133]);
    assign outputs[5346] = ~(layer2_outputs[2220]);
    assign outputs[5347] = layer2_outputs[6438];
    assign outputs[5348] = ~((layer2_outputs[4730]) ^ (layer2_outputs[2837]));
    assign outputs[5349] = ~(layer2_outputs[6305]);
    assign outputs[5350] = layer2_outputs[5989];
    assign outputs[5351] = ~(layer2_outputs[5699]);
    assign outputs[5352] = ~(layer2_outputs[8859]);
    assign outputs[5353] = (layer2_outputs[1952]) & ~(layer2_outputs[8000]);
    assign outputs[5354] = layer2_outputs[7906];
    assign outputs[5355] = ~(layer2_outputs[1326]);
    assign outputs[5356] = layer2_outputs[11378];
    assign outputs[5357] = layer2_outputs[5730];
    assign outputs[5358] = ~(layer2_outputs[2384]);
    assign outputs[5359] = ~(layer2_outputs[12602]);
    assign outputs[5360] = ~(layer2_outputs[3333]) | (layer2_outputs[1469]);
    assign outputs[5361] = layer2_outputs[2382];
    assign outputs[5362] = ~(layer2_outputs[3317]);
    assign outputs[5363] = (layer2_outputs[11289]) ^ (layer2_outputs[46]);
    assign outputs[5364] = ~(layer2_outputs[1268]);
    assign outputs[5365] = ~(layer2_outputs[9600]) | (layer2_outputs[8346]);
    assign outputs[5366] = ~(layer2_outputs[8372]);
    assign outputs[5367] = (layer2_outputs[12506]) & ~(layer2_outputs[191]);
    assign outputs[5368] = ~((layer2_outputs[9331]) ^ (layer2_outputs[7300]));
    assign outputs[5369] = layer2_outputs[2358];
    assign outputs[5370] = layer2_outputs[11111];
    assign outputs[5371] = ~(layer2_outputs[904]);
    assign outputs[5372] = ~(layer2_outputs[3374]);
    assign outputs[5373] = ~((layer2_outputs[9480]) ^ (layer2_outputs[10167]));
    assign outputs[5374] = ~((layer2_outputs[2770]) ^ (layer2_outputs[1059]));
    assign outputs[5375] = (layer2_outputs[8805]) & ~(layer2_outputs[9426]);
    assign outputs[5376] = ~(layer2_outputs[5962]);
    assign outputs[5377] = ~((layer2_outputs[7012]) | (layer2_outputs[5662]));
    assign outputs[5378] = (layer2_outputs[885]) ^ (layer2_outputs[5913]);
    assign outputs[5379] = (layer2_outputs[2987]) & (layer2_outputs[1070]);
    assign outputs[5380] = layer2_outputs[3082];
    assign outputs[5381] = layer2_outputs[8190];
    assign outputs[5382] = ~(layer2_outputs[6110]);
    assign outputs[5383] = layer2_outputs[6137];
    assign outputs[5384] = ~(layer2_outputs[4357]);
    assign outputs[5385] = layer2_outputs[5632];
    assign outputs[5386] = layer2_outputs[4870];
    assign outputs[5387] = layer2_outputs[6199];
    assign outputs[5388] = (layer2_outputs[6181]) & ~(layer2_outputs[8229]);
    assign outputs[5389] = ~(layer2_outputs[5859]);
    assign outputs[5390] = ~(layer2_outputs[725]);
    assign outputs[5391] = ~((layer2_outputs[9602]) ^ (layer2_outputs[5841]));
    assign outputs[5392] = ~((layer2_outputs[8833]) & (layer2_outputs[10766]));
    assign outputs[5393] = layer2_outputs[5932];
    assign outputs[5394] = (layer2_outputs[539]) | (layer2_outputs[7725]);
    assign outputs[5395] = (layer2_outputs[8273]) ^ (layer2_outputs[10710]);
    assign outputs[5396] = (layer2_outputs[11344]) ^ (layer2_outputs[4607]);
    assign outputs[5397] = ~(layer2_outputs[12284]);
    assign outputs[5398] = ~(layer2_outputs[5324]);
    assign outputs[5399] = ~(layer2_outputs[11]) | (layer2_outputs[11950]);
    assign outputs[5400] = layer2_outputs[6425];
    assign outputs[5401] = ~(layer2_outputs[2496]);
    assign outputs[5402] = ~(layer2_outputs[9106]);
    assign outputs[5403] = ~(layer2_outputs[8802]) | (layer2_outputs[6225]);
    assign outputs[5404] = (layer2_outputs[5770]) & ~(layer2_outputs[12353]);
    assign outputs[5405] = ~((layer2_outputs[10182]) | (layer2_outputs[9500]));
    assign outputs[5406] = (layer2_outputs[5253]) ^ (layer2_outputs[5199]);
    assign outputs[5407] = ~(layer2_outputs[10321]);
    assign outputs[5408] = ~((layer2_outputs[11086]) ^ (layer2_outputs[810]));
    assign outputs[5409] = ~(layer2_outputs[11314]);
    assign outputs[5410] = (layer2_outputs[10048]) ^ (layer2_outputs[10642]);
    assign outputs[5411] = ~((layer2_outputs[7451]) ^ (layer2_outputs[2438]));
    assign outputs[5412] = (layer2_outputs[223]) ^ (layer2_outputs[5344]);
    assign outputs[5413] = ~(layer2_outputs[12660]);
    assign outputs[5414] = ~(layer2_outputs[2039]);
    assign outputs[5415] = ~(layer2_outputs[2734]);
    assign outputs[5416] = layer2_outputs[2825];
    assign outputs[5417] = layer2_outputs[7963];
    assign outputs[5418] = (layer2_outputs[295]) ^ (layer2_outputs[12337]);
    assign outputs[5419] = ~(layer2_outputs[343]);
    assign outputs[5420] = ~(layer2_outputs[3345]);
    assign outputs[5421] = ~((layer2_outputs[6625]) & (layer2_outputs[2999]));
    assign outputs[5422] = ~(layer2_outputs[7662]);
    assign outputs[5423] = (layer2_outputs[10867]) ^ (layer2_outputs[8112]);
    assign outputs[5424] = ~(layer2_outputs[1302]) | (layer2_outputs[598]);
    assign outputs[5425] = ~((layer2_outputs[9990]) ^ (layer2_outputs[5589]));
    assign outputs[5426] = ~(layer2_outputs[5777]) | (layer2_outputs[11080]);
    assign outputs[5427] = (layer2_outputs[6486]) | (layer2_outputs[12472]);
    assign outputs[5428] = layer2_outputs[12296];
    assign outputs[5429] = ~(layer2_outputs[3139]);
    assign outputs[5430] = layer2_outputs[11763];
    assign outputs[5431] = (layer2_outputs[4739]) & ~(layer2_outputs[2509]);
    assign outputs[5432] = ~(layer2_outputs[4558]);
    assign outputs[5433] = layer2_outputs[2647];
    assign outputs[5434] = layer2_outputs[12174];
    assign outputs[5435] = ~((layer2_outputs[7627]) | (layer2_outputs[2193]));
    assign outputs[5436] = layer2_outputs[6381];
    assign outputs[5437] = (layer2_outputs[4194]) | (layer2_outputs[7162]);
    assign outputs[5438] = ~(layer2_outputs[12444]);
    assign outputs[5439] = (layer2_outputs[8859]) ^ (layer2_outputs[11303]);
    assign outputs[5440] = (layer2_outputs[797]) & ~(layer2_outputs[4169]);
    assign outputs[5441] = layer2_outputs[3393];
    assign outputs[5442] = ~(layer2_outputs[3016]);
    assign outputs[5443] = (layer2_outputs[1186]) & (layer2_outputs[9586]);
    assign outputs[5444] = (layer2_outputs[12332]) & ~(layer2_outputs[4594]);
    assign outputs[5445] = ~(layer2_outputs[5215]);
    assign outputs[5446] = layer2_outputs[12143];
    assign outputs[5447] = layer2_outputs[1421];
    assign outputs[5448] = layer2_outputs[10807];
    assign outputs[5449] = ~(layer2_outputs[11096]);
    assign outputs[5450] = layer2_outputs[3760];
    assign outputs[5451] = (layer2_outputs[4387]) ^ (layer2_outputs[10685]);
    assign outputs[5452] = layer2_outputs[1260];
    assign outputs[5453] = layer2_outputs[6325];
    assign outputs[5454] = layer2_outputs[2453];
    assign outputs[5455] = (layer2_outputs[2402]) ^ (layer2_outputs[4746]);
    assign outputs[5456] = ~(layer2_outputs[8847]) | (layer2_outputs[1090]);
    assign outputs[5457] = ~(layer2_outputs[6496]);
    assign outputs[5458] = layer2_outputs[12410];
    assign outputs[5459] = layer2_outputs[10109];
    assign outputs[5460] = ~(layer2_outputs[4251]) | (layer2_outputs[7372]);
    assign outputs[5461] = layer2_outputs[4477];
    assign outputs[5462] = ~(layer2_outputs[10216]);
    assign outputs[5463] = ~((layer2_outputs[11642]) & (layer2_outputs[4986]));
    assign outputs[5464] = ~(layer2_outputs[4466]);
    assign outputs[5465] = ~((layer2_outputs[6426]) | (layer2_outputs[4906]));
    assign outputs[5466] = (layer2_outputs[12760]) & ~(layer2_outputs[1986]);
    assign outputs[5467] = ~(layer2_outputs[10811]);
    assign outputs[5468] = layer2_outputs[7976];
    assign outputs[5469] = (layer2_outputs[622]) ^ (layer2_outputs[3800]);
    assign outputs[5470] = ~((layer2_outputs[103]) ^ (layer2_outputs[12762]));
    assign outputs[5471] = ~((layer2_outputs[1045]) ^ (layer2_outputs[2421]));
    assign outputs[5472] = ~(layer2_outputs[5527]);
    assign outputs[5473] = ~(layer2_outputs[10231]);
    assign outputs[5474] = ~(layer2_outputs[11771]);
    assign outputs[5475] = layer2_outputs[3556];
    assign outputs[5476] = layer2_outputs[11364];
    assign outputs[5477] = (layer2_outputs[6124]) & (layer2_outputs[2062]);
    assign outputs[5478] = ~(layer2_outputs[3112]);
    assign outputs[5479] = ~(layer2_outputs[4951]);
    assign outputs[5480] = ~((layer2_outputs[5665]) ^ (layer2_outputs[6454]));
    assign outputs[5481] = ~(layer2_outputs[6860]);
    assign outputs[5482] = (layer2_outputs[9542]) & ~(layer2_outputs[11226]);
    assign outputs[5483] = layer2_outputs[10603];
    assign outputs[5484] = layer2_outputs[5601];
    assign outputs[5485] = layer2_outputs[12474];
    assign outputs[5486] = ~(layer2_outputs[8386]) | (layer2_outputs[4173]);
    assign outputs[5487] = ~((layer2_outputs[9116]) ^ (layer2_outputs[10291]));
    assign outputs[5488] = ~(layer2_outputs[4256]);
    assign outputs[5489] = layer2_outputs[2981];
    assign outputs[5490] = ~(layer2_outputs[4189]);
    assign outputs[5491] = layer2_outputs[10849];
    assign outputs[5492] = ~(layer2_outputs[9721]);
    assign outputs[5493] = ~((layer2_outputs[9358]) ^ (layer2_outputs[5855]));
    assign outputs[5494] = (layer2_outputs[9115]) & ~(layer2_outputs[10219]);
    assign outputs[5495] = ~(layer2_outputs[10165]) | (layer2_outputs[1802]);
    assign outputs[5496] = ~(layer2_outputs[11521]);
    assign outputs[5497] = ~((layer2_outputs[265]) ^ (layer2_outputs[6014]));
    assign outputs[5498] = ~(layer2_outputs[3618]);
    assign outputs[5499] = ~(layer2_outputs[799]);
    assign outputs[5500] = (layer2_outputs[5893]) ^ (layer2_outputs[9850]);
    assign outputs[5501] = ~(layer2_outputs[374]);
    assign outputs[5502] = (layer2_outputs[7100]) ^ (layer2_outputs[6058]);
    assign outputs[5503] = layer2_outputs[12300];
    assign outputs[5504] = ~((layer2_outputs[8025]) ^ (layer2_outputs[1742]));
    assign outputs[5505] = (layer2_outputs[5833]) ^ (layer2_outputs[5550]);
    assign outputs[5506] = (layer2_outputs[5767]) ^ (layer2_outputs[9432]);
    assign outputs[5507] = ~((layer2_outputs[10742]) ^ (layer2_outputs[7014]));
    assign outputs[5508] = (layer2_outputs[4080]) | (layer2_outputs[10577]);
    assign outputs[5509] = layer2_outputs[11372];
    assign outputs[5510] = (layer2_outputs[9093]) ^ (layer2_outputs[10310]);
    assign outputs[5511] = (layer2_outputs[7803]) & (layer2_outputs[11119]);
    assign outputs[5512] = ~(layer2_outputs[10700]);
    assign outputs[5513] = layer2_outputs[3730];
    assign outputs[5514] = (layer2_outputs[7390]) & ~(layer2_outputs[5137]);
    assign outputs[5515] = (layer2_outputs[11055]) & (layer2_outputs[122]);
    assign outputs[5516] = ~(layer2_outputs[5588]) | (layer2_outputs[1862]);
    assign outputs[5517] = layer2_outputs[8021];
    assign outputs[5518] = (layer2_outputs[390]) ^ (layer2_outputs[6133]);
    assign outputs[5519] = layer2_outputs[9645];
    assign outputs[5520] = ~(layer2_outputs[11174]);
    assign outputs[5521] = layer2_outputs[8230];
    assign outputs[5522] = layer2_outputs[2122];
    assign outputs[5523] = ~(layer2_outputs[512]);
    assign outputs[5524] = ~((layer2_outputs[11665]) ^ (layer2_outputs[3747]));
    assign outputs[5525] = ~(layer2_outputs[1461]);
    assign outputs[5526] = (layer2_outputs[3758]) ^ (layer2_outputs[10770]);
    assign outputs[5527] = (layer2_outputs[10303]) ^ (layer2_outputs[6837]);
    assign outputs[5528] = (layer2_outputs[3960]) & (layer2_outputs[12388]);
    assign outputs[5529] = layer2_outputs[1616];
    assign outputs[5530] = layer2_outputs[6418];
    assign outputs[5531] = ~((layer2_outputs[12252]) | (layer2_outputs[10113]));
    assign outputs[5532] = (layer2_outputs[2849]) & (layer2_outputs[2293]);
    assign outputs[5533] = ~((layer2_outputs[2671]) & (layer2_outputs[12190]));
    assign outputs[5534] = ~((layer2_outputs[2352]) ^ (layer2_outputs[12549]));
    assign outputs[5535] = ~(layer2_outputs[11324]);
    assign outputs[5536] = layer2_outputs[4911];
    assign outputs[5537] = (layer2_outputs[3335]) & (layer2_outputs[8358]);
    assign outputs[5538] = ~(layer2_outputs[23]);
    assign outputs[5539] = layer2_outputs[1642];
    assign outputs[5540] = ~(layer2_outputs[3146]);
    assign outputs[5541] = (layer2_outputs[1623]) ^ (layer2_outputs[6134]);
    assign outputs[5542] = ~((layer2_outputs[1405]) & (layer2_outputs[11014]));
    assign outputs[5543] = (layer2_outputs[4214]) ^ (layer2_outputs[8985]);
    assign outputs[5544] = ~(layer2_outputs[988]);
    assign outputs[5545] = layer2_outputs[775];
    assign outputs[5546] = ~((layer2_outputs[8169]) ^ (layer2_outputs[2272]));
    assign outputs[5547] = ~(layer2_outputs[1747]) | (layer2_outputs[11638]);
    assign outputs[5548] = (layer2_outputs[10073]) | (layer2_outputs[8257]);
    assign outputs[5549] = layer2_outputs[6132];
    assign outputs[5550] = ~(layer2_outputs[3321]);
    assign outputs[5551] = layer2_outputs[3723];
    assign outputs[5552] = ~(layer2_outputs[8530]);
    assign outputs[5553] = ~(layer2_outputs[5553]);
    assign outputs[5554] = layer2_outputs[10143];
    assign outputs[5555] = ~((layer2_outputs[2105]) ^ (layer2_outputs[12095]));
    assign outputs[5556] = ~(layer2_outputs[4670]) | (layer2_outputs[11172]);
    assign outputs[5557] = layer2_outputs[1575];
    assign outputs[5558] = ~(layer2_outputs[627]);
    assign outputs[5559] = ~(layer2_outputs[11585]);
    assign outputs[5560] = layer2_outputs[5054];
    assign outputs[5561] = (layer2_outputs[208]) ^ (layer2_outputs[1149]);
    assign outputs[5562] = ~(layer2_outputs[4403]);
    assign outputs[5563] = layer2_outputs[11801];
    assign outputs[5564] = ~(layer2_outputs[2316]);
    assign outputs[5565] = (layer2_outputs[6802]) & ~(layer2_outputs[1793]);
    assign outputs[5566] = (layer2_outputs[6337]) ^ (layer2_outputs[6673]);
    assign outputs[5567] = layer2_outputs[10524];
    assign outputs[5568] = (layer2_outputs[1654]) ^ (layer2_outputs[7711]);
    assign outputs[5569] = ~(layer2_outputs[2384]);
    assign outputs[5570] = layer2_outputs[11922];
    assign outputs[5571] = layer2_outputs[6685];
    assign outputs[5572] = ~(layer2_outputs[1841]);
    assign outputs[5573] = layer2_outputs[8580];
    assign outputs[5574] = layer2_outputs[4561];
    assign outputs[5575] = ~((layer2_outputs[206]) ^ (layer2_outputs[472]));
    assign outputs[5576] = ~(layer2_outputs[12075]);
    assign outputs[5577] = ~(layer2_outputs[8770]);
    assign outputs[5578] = ~((layer2_outputs[2635]) ^ (layer2_outputs[6139]));
    assign outputs[5579] = ~(layer2_outputs[3820]);
    assign outputs[5580] = layer2_outputs[6107];
    assign outputs[5581] = ~((layer2_outputs[8197]) ^ (layer2_outputs[6762]));
    assign outputs[5582] = (layer2_outputs[185]) ^ (layer2_outputs[4024]);
    assign outputs[5583] = ~(layer2_outputs[7738]) | (layer2_outputs[5246]);
    assign outputs[5584] = (layer2_outputs[8619]) & (layer2_outputs[688]);
    assign outputs[5585] = ~(layer2_outputs[7369]);
    assign outputs[5586] = (layer2_outputs[1126]) ^ (layer2_outputs[4086]);
    assign outputs[5587] = ~((layer2_outputs[8442]) ^ (layer2_outputs[8727]));
    assign outputs[5588] = ~(layer2_outputs[9954]);
    assign outputs[5589] = ~(layer2_outputs[5536]);
    assign outputs[5590] = layer2_outputs[4933];
    assign outputs[5591] = layer2_outputs[5818];
    assign outputs[5592] = layer2_outputs[1719];
    assign outputs[5593] = ~((layer2_outputs[8776]) | (layer2_outputs[1191]));
    assign outputs[5594] = ~(layer2_outputs[7309]);
    assign outputs[5595] = ~((layer2_outputs[3268]) ^ (layer2_outputs[8752]));
    assign outputs[5596] = (layer2_outputs[8380]) ^ (layer2_outputs[1384]);
    assign outputs[5597] = ~(layer2_outputs[12568]);
    assign outputs[5598] = ~(layer2_outputs[7227]);
    assign outputs[5599] = layer2_outputs[1941];
    assign outputs[5600] = (layer2_outputs[4976]) & ~(layer2_outputs[2077]);
    assign outputs[5601] = ~((layer2_outputs[2505]) ^ (layer2_outputs[10695]));
    assign outputs[5602] = ~(layer2_outputs[8088]);
    assign outputs[5603] = ~((layer2_outputs[11466]) ^ (layer2_outputs[363]));
    assign outputs[5604] = (layer2_outputs[5988]) ^ (layer2_outputs[8713]);
    assign outputs[5605] = ~((layer2_outputs[3847]) ^ (layer2_outputs[10736]));
    assign outputs[5606] = layer2_outputs[6886];
    assign outputs[5607] = layer2_outputs[3318];
    assign outputs[5608] = (layer2_outputs[1570]) ^ (layer2_outputs[2312]);
    assign outputs[5609] = layer2_outputs[5187];
    assign outputs[5610] = ~(layer2_outputs[2839]) | (layer2_outputs[1856]);
    assign outputs[5611] = ~(layer2_outputs[3180]);
    assign outputs[5612] = ~(layer2_outputs[9958]);
    assign outputs[5613] = ~((layer2_outputs[4526]) ^ (layer2_outputs[1619]));
    assign outputs[5614] = ~(layer2_outputs[7986]);
    assign outputs[5615] = (layer2_outputs[4118]) ^ (layer2_outputs[11218]);
    assign outputs[5616] = layer2_outputs[10881];
    assign outputs[5617] = (layer2_outputs[3409]) ^ (layer2_outputs[3094]);
    assign outputs[5618] = ~(layer2_outputs[2345]);
    assign outputs[5619] = ~(layer2_outputs[274]) | (layer2_outputs[5752]);
    assign outputs[5620] = ~(layer2_outputs[6779]);
    assign outputs[5621] = layer2_outputs[12342];
    assign outputs[5622] = (layer2_outputs[10087]) ^ (layer2_outputs[1320]);
    assign outputs[5623] = ~((layer2_outputs[84]) & (layer2_outputs[8955]));
    assign outputs[5624] = (layer2_outputs[524]) ^ (layer2_outputs[613]);
    assign outputs[5625] = layer2_outputs[4440];
    assign outputs[5626] = (layer2_outputs[5935]) ^ (layer2_outputs[9372]);
    assign outputs[5627] = (layer2_outputs[1229]) & (layer2_outputs[461]);
    assign outputs[5628] = ~((layer2_outputs[4021]) ^ (layer2_outputs[8556]));
    assign outputs[5629] = ~(layer2_outputs[1751]);
    assign outputs[5630] = ~(layer2_outputs[10985]);
    assign outputs[5631] = ~((layer2_outputs[11209]) ^ (layer2_outputs[1016]));
    assign outputs[5632] = (layer2_outputs[3378]) ^ (layer2_outputs[9234]);
    assign outputs[5633] = (layer2_outputs[12170]) ^ (layer2_outputs[12742]);
    assign outputs[5634] = layer2_outputs[10129];
    assign outputs[5635] = ~((layer2_outputs[6390]) ^ (layer2_outputs[301]));
    assign outputs[5636] = (layer2_outputs[1231]) ^ (layer2_outputs[10684]);
    assign outputs[5637] = layer2_outputs[10183];
    assign outputs[5638] = ~(layer2_outputs[8391]);
    assign outputs[5639] = ~(layer2_outputs[2171]);
    assign outputs[5640] = ~(layer2_outputs[4494]);
    assign outputs[5641] = (layer2_outputs[9759]) & ~(layer2_outputs[9432]);
    assign outputs[5642] = ~(layer2_outputs[11939]);
    assign outputs[5643] = ~((layer2_outputs[11613]) | (layer2_outputs[2959]));
    assign outputs[5644] = ~((layer2_outputs[1810]) ^ (layer2_outputs[9611]));
    assign outputs[5645] = ~(layer2_outputs[6512]);
    assign outputs[5646] = ~((layer2_outputs[7154]) ^ (layer2_outputs[7377]));
    assign outputs[5647] = ~(layer2_outputs[1391]);
    assign outputs[5648] = (layer2_outputs[2889]) ^ (layer2_outputs[10140]);
    assign outputs[5649] = ~(layer2_outputs[3180]);
    assign outputs[5650] = (layer2_outputs[6736]) & (layer2_outputs[5304]);
    assign outputs[5651] = layer2_outputs[7083];
    assign outputs[5652] = ~((layer2_outputs[5442]) ^ (layer2_outputs[309]));
    assign outputs[5653] = (layer2_outputs[6787]) ^ (layer2_outputs[11035]);
    assign outputs[5654] = ~(layer2_outputs[259]);
    assign outputs[5655] = layer2_outputs[3669];
    assign outputs[5656] = ~(layer2_outputs[108]);
    assign outputs[5657] = ~(layer2_outputs[1975]);
    assign outputs[5658] = ~(layer2_outputs[9110]);
    assign outputs[5659] = ~(layer2_outputs[9076]);
    assign outputs[5660] = layer2_outputs[4861];
    assign outputs[5661] = layer2_outputs[195];
    assign outputs[5662] = layer2_outputs[10910];
    assign outputs[5663] = layer2_outputs[11330];
    assign outputs[5664] = ~((layer2_outputs[3790]) & (layer2_outputs[10824]));
    assign outputs[5665] = (layer2_outputs[3590]) & ~(layer2_outputs[8299]);
    assign outputs[5666] = layer2_outputs[8960];
    assign outputs[5667] = ~((layer2_outputs[10209]) ^ (layer2_outputs[10016]));
    assign outputs[5668] = layer2_outputs[5329];
    assign outputs[5669] = layer2_outputs[8041];
    assign outputs[5670] = ~((layer2_outputs[12090]) ^ (layer2_outputs[1811]));
    assign outputs[5671] = layer2_outputs[4496];
    assign outputs[5672] = layer2_outputs[3730];
    assign outputs[5673] = (layer2_outputs[9395]) ^ (layer2_outputs[5227]);
    assign outputs[5674] = ~(layer2_outputs[577]);
    assign outputs[5675] = layer2_outputs[1288];
    assign outputs[5676] = ~(layer2_outputs[4728]);
    assign outputs[5677] = layer2_outputs[5559];
    assign outputs[5678] = ~(layer2_outputs[7819]);
    assign outputs[5679] = (layer2_outputs[11117]) & ~(layer2_outputs[6729]);
    assign outputs[5680] = (layer2_outputs[3215]) & (layer2_outputs[12433]);
    assign outputs[5681] = ~(layer2_outputs[2754]);
    assign outputs[5682] = ~(layer2_outputs[7069]);
    assign outputs[5683] = (layer2_outputs[11350]) & (layer2_outputs[72]);
    assign outputs[5684] = (layer2_outputs[12421]) ^ (layer2_outputs[6822]);
    assign outputs[5685] = ~((layer2_outputs[8177]) ^ (layer2_outputs[11536]));
    assign outputs[5686] = ~(layer2_outputs[9206]);
    assign outputs[5687] = ~((layer2_outputs[9041]) | (layer2_outputs[3429]));
    assign outputs[5688] = layer2_outputs[2064];
    assign outputs[5689] = ~(layer2_outputs[4157]);
    assign outputs[5690] = ~(layer2_outputs[3966]);
    assign outputs[5691] = (layer2_outputs[2195]) ^ (layer2_outputs[10851]);
    assign outputs[5692] = ~((layer2_outputs[5199]) ^ (layer2_outputs[11673]));
    assign outputs[5693] = ~(layer2_outputs[2538]) | (layer2_outputs[12681]);
    assign outputs[5694] = ~(layer2_outputs[544]);
    assign outputs[5695] = ~(layer2_outputs[4512]);
    assign outputs[5696] = ~(layer2_outputs[7473]);
    assign outputs[5697] = layer2_outputs[1590];
    assign outputs[5698] = ~((layer2_outputs[11891]) ^ (layer2_outputs[4263]));
    assign outputs[5699] = (layer2_outputs[7756]) ^ (layer2_outputs[3884]);
    assign outputs[5700] = layer2_outputs[6051];
    assign outputs[5701] = ~(layer2_outputs[9896]);
    assign outputs[5702] = layer2_outputs[11249];
    assign outputs[5703] = (layer2_outputs[6879]) ^ (layer2_outputs[7125]);
    assign outputs[5704] = (layer2_outputs[7006]) ^ (layer2_outputs[4863]);
    assign outputs[5705] = layer2_outputs[8721];
    assign outputs[5706] = ~(layer2_outputs[2812]);
    assign outputs[5707] = ~(layer2_outputs[9504]);
    assign outputs[5708] = ~((layer2_outputs[5819]) | (layer2_outputs[6848]));
    assign outputs[5709] = ~(layer2_outputs[3350]);
    assign outputs[5710] = ~((layer2_outputs[11271]) ^ (layer2_outputs[3205]));
    assign outputs[5711] = layer2_outputs[7305];
    assign outputs[5712] = ~(layer2_outputs[3371]);
    assign outputs[5713] = ~(layer2_outputs[2971]);
    assign outputs[5714] = layer2_outputs[2396];
    assign outputs[5715] = ~(layer2_outputs[4782]);
    assign outputs[5716] = ~(layer2_outputs[7694]);
    assign outputs[5717] = ~(layer2_outputs[8683]);
    assign outputs[5718] = layer2_outputs[11658];
    assign outputs[5719] = layer2_outputs[1435];
    assign outputs[5720] = ~(layer2_outputs[7975]);
    assign outputs[5721] = ~((layer2_outputs[1968]) ^ (layer2_outputs[176]));
    assign outputs[5722] = ~(layer2_outputs[3128]);
    assign outputs[5723] = ~(layer2_outputs[5021]);
    assign outputs[5724] = (layer2_outputs[12706]) | (layer2_outputs[1262]);
    assign outputs[5725] = layer2_outputs[11063];
    assign outputs[5726] = ~(layer2_outputs[60]);
    assign outputs[5727] = ~(layer2_outputs[1185]);
    assign outputs[5728] = layer2_outputs[5280];
    assign outputs[5729] = ~(layer2_outputs[9375]);
    assign outputs[5730] = (layer2_outputs[8048]) | (layer2_outputs[5931]);
    assign outputs[5731] = layer2_outputs[8828];
    assign outputs[5732] = (layer2_outputs[11402]) ^ (layer2_outputs[4063]);
    assign outputs[5733] = layer2_outputs[5558];
    assign outputs[5734] = ~(layer2_outputs[1617]);
    assign outputs[5735] = (layer2_outputs[3639]) ^ (layer2_outputs[7273]);
    assign outputs[5736] = ~(layer2_outputs[11747]);
    assign outputs[5737] = ~(layer2_outputs[6913]);
    assign outputs[5738] = ~(layer2_outputs[9527]);
    assign outputs[5739] = ~((layer2_outputs[2899]) ^ (layer2_outputs[5205]));
    assign outputs[5740] = ~(layer2_outputs[5250]);
    assign outputs[5741] = layer2_outputs[4219];
    assign outputs[5742] = ~(layer2_outputs[11091]);
    assign outputs[5743] = (layer2_outputs[10886]) ^ (layer2_outputs[1303]);
    assign outputs[5744] = ~(layer2_outputs[12377]);
    assign outputs[5745] = ~(layer2_outputs[11032]);
    assign outputs[5746] = ~((layer2_outputs[7243]) ^ (layer2_outputs[11388]));
    assign outputs[5747] = ~(layer2_outputs[4610]);
    assign outputs[5748] = layer2_outputs[4132];
    assign outputs[5749] = layer2_outputs[12058];
    assign outputs[5750] = (layer2_outputs[8937]) & ~(layer2_outputs[1597]);
    assign outputs[5751] = layer2_outputs[3675];
    assign outputs[5752] = layer2_outputs[6411];
    assign outputs[5753] = ~(layer2_outputs[6303]);
    assign outputs[5754] = ~((layer2_outputs[1908]) | (layer2_outputs[11367]));
    assign outputs[5755] = ~((layer2_outputs[7745]) ^ (layer2_outputs[5637]));
    assign outputs[5756] = (layer2_outputs[6405]) | (layer2_outputs[1336]);
    assign outputs[5757] = ~(layer2_outputs[12305]);
    assign outputs[5758] = layer2_outputs[11410];
    assign outputs[5759] = layer2_outputs[1973];
    assign outputs[5760] = ~((layer2_outputs[11941]) | (layer2_outputs[8871]));
    assign outputs[5761] = (layer2_outputs[6300]) ^ (layer2_outputs[8734]);
    assign outputs[5762] = ~((layer2_outputs[7655]) & (layer2_outputs[7192]));
    assign outputs[5763] = (layer2_outputs[5532]) & ~(layer2_outputs[8797]);
    assign outputs[5764] = layer2_outputs[6777];
    assign outputs[5765] = ~(layer2_outputs[1276]);
    assign outputs[5766] = layer2_outputs[11511];
    assign outputs[5767] = (layer2_outputs[4947]) ^ (layer2_outputs[6297]);
    assign outputs[5768] = ~((layer2_outputs[4731]) ^ (layer2_outputs[11309]));
    assign outputs[5769] = ~(layer2_outputs[5620]);
    assign outputs[5770] = (layer2_outputs[10820]) ^ (layer2_outputs[6248]);
    assign outputs[5771] = (layer2_outputs[10874]) ^ (layer2_outputs[2136]);
    assign outputs[5772] = ~((layer2_outputs[7115]) ^ (layer2_outputs[6714]));
    assign outputs[5773] = layer2_outputs[9761];
    assign outputs[5774] = (layer2_outputs[10650]) & (layer2_outputs[3416]);
    assign outputs[5775] = ~(layer2_outputs[6731]);
    assign outputs[5776] = layer2_outputs[8639];
    assign outputs[5777] = ~(layer2_outputs[7668]);
    assign outputs[5778] = ~(layer2_outputs[7393]) | (layer2_outputs[6293]);
    assign outputs[5779] = ~((layer2_outputs[8174]) ^ (layer2_outputs[8151]));
    assign outputs[5780] = (layer2_outputs[3819]) ^ (layer2_outputs[12355]);
    assign outputs[5781] = layer2_outputs[1890];
    assign outputs[5782] = ~((layer2_outputs[9592]) | (layer2_outputs[5259]));
    assign outputs[5783] = layer2_outputs[323];
    assign outputs[5784] = (layer2_outputs[3007]) ^ (layer2_outputs[7548]);
    assign outputs[5785] = (layer2_outputs[4965]) ^ (layer2_outputs[669]);
    assign outputs[5786] = ~(layer2_outputs[9202]) | (layer2_outputs[10544]);
    assign outputs[5787] = ~(layer2_outputs[8621]);
    assign outputs[5788] = ~(layer2_outputs[11555]) | (layer2_outputs[8271]);
    assign outputs[5789] = layer2_outputs[11351];
    assign outputs[5790] = layer2_outputs[7362];
    assign outputs[5791] = layer2_outputs[2690];
    assign outputs[5792] = ~(layer2_outputs[4736]) | (layer2_outputs[1632]);
    assign outputs[5793] = layer2_outputs[3387];
    assign outputs[5794] = layer2_outputs[6148];
    assign outputs[5795] = (layer2_outputs[3999]) | (layer2_outputs[2837]);
    assign outputs[5796] = ~(layer2_outputs[1212]);
    assign outputs[5797] = (layer2_outputs[12372]) ^ (layer2_outputs[10178]);
    assign outputs[5798] = layer2_outputs[9939];
    assign outputs[5799] = ~(layer2_outputs[12135]);
    assign outputs[5800] = layer2_outputs[713];
    assign outputs[5801] = (layer2_outputs[11549]) ^ (layer2_outputs[10927]);
    assign outputs[5802] = (layer2_outputs[11902]) ^ (layer2_outputs[6142]);
    assign outputs[5803] = layer2_outputs[8287];
    assign outputs[5804] = (layer2_outputs[2833]) & (layer2_outputs[5867]);
    assign outputs[5805] = layer2_outputs[3753];
    assign outputs[5806] = layer2_outputs[3057];
    assign outputs[5807] = (layer2_outputs[10009]) & ~(layer2_outputs[3049]);
    assign outputs[5808] = ~(layer2_outputs[4078]);
    assign outputs[5809] = (layer2_outputs[6332]) ^ (layer2_outputs[9913]);
    assign outputs[5810] = ~(layer2_outputs[9246]) | (layer2_outputs[1226]);
    assign outputs[5811] = layer2_outputs[7237];
    assign outputs[5812] = layer2_outputs[8221];
    assign outputs[5813] = layer2_outputs[8154];
    assign outputs[5814] = layer2_outputs[8790];
    assign outputs[5815] = ~((layer2_outputs[4184]) ^ (layer2_outputs[7690]));
    assign outputs[5816] = ~((layer2_outputs[12004]) & (layer2_outputs[4991]));
    assign outputs[5817] = ~((layer2_outputs[2102]) ^ (layer2_outputs[7194]));
    assign outputs[5818] = ~(layer2_outputs[3151]);
    assign outputs[5819] = (layer2_outputs[4103]) & ~(layer2_outputs[3817]);
    assign outputs[5820] = ~((layer2_outputs[10696]) ^ (layer2_outputs[10998]));
    assign outputs[5821] = (layer2_outputs[8344]) ^ (layer2_outputs[1413]);
    assign outputs[5822] = ~(layer2_outputs[302]);
    assign outputs[5823] = layer2_outputs[9972];
    assign outputs[5824] = layer2_outputs[9472];
    assign outputs[5825] = layer2_outputs[4703];
    assign outputs[5826] = ~((layer2_outputs[384]) ^ (layer2_outputs[2494]));
    assign outputs[5827] = ~(layer2_outputs[9279]);
    assign outputs[5828] = ~(layer2_outputs[8068]);
    assign outputs[5829] = (layer2_outputs[2449]) ^ (layer2_outputs[4166]);
    assign outputs[5830] = ~(layer2_outputs[2674]);
    assign outputs[5831] = ~(layer2_outputs[9004]);
    assign outputs[5832] = (layer2_outputs[2844]) ^ (layer2_outputs[12243]);
    assign outputs[5833] = ~(layer2_outputs[5521]);
    assign outputs[5834] = (layer2_outputs[6965]) ^ (layer2_outputs[6947]);
    assign outputs[5835] = (layer2_outputs[10012]) | (layer2_outputs[907]);
    assign outputs[5836] = ~((layer2_outputs[60]) ^ (layer2_outputs[2355]));
    assign outputs[5837] = ~((layer2_outputs[2262]) | (layer2_outputs[8138]));
    assign outputs[5838] = (layer2_outputs[790]) & ~(layer2_outputs[1523]);
    assign outputs[5839] = ~(layer2_outputs[598]) | (layer2_outputs[3236]);
    assign outputs[5840] = layer2_outputs[5288];
    assign outputs[5841] = (layer2_outputs[9947]) & (layer2_outputs[1238]);
    assign outputs[5842] = ~(layer2_outputs[10749]);
    assign outputs[5843] = layer2_outputs[4832];
    assign outputs[5844] = ~(layer2_outputs[6764]);
    assign outputs[5845] = ~(layer2_outputs[6742]);
    assign outputs[5846] = layer2_outputs[7464];
    assign outputs[5847] = ~(layer2_outputs[1503]);
    assign outputs[5848] = ~(layer2_outputs[12420]);
    assign outputs[5849] = ~(layer2_outputs[8039]);
    assign outputs[5850] = ~(layer2_outputs[10841]);
    assign outputs[5851] = layer2_outputs[2103];
    assign outputs[5852] = layer2_outputs[535];
    assign outputs[5853] = layer2_outputs[6938];
    assign outputs[5854] = (layer2_outputs[12663]) ^ (layer2_outputs[6989]);
    assign outputs[5855] = ~(layer2_outputs[12413]);
    assign outputs[5856] = ~((layer2_outputs[3765]) ^ (layer2_outputs[895]));
    assign outputs[5857] = layer2_outputs[3545];
    assign outputs[5858] = ~(layer2_outputs[2200]);
    assign outputs[5859] = (layer2_outputs[5310]) | (layer2_outputs[10779]);
    assign outputs[5860] = ~(layer2_outputs[6833]);
    assign outputs[5861] = ~(layer2_outputs[3928]);
    assign outputs[5862] = layer2_outputs[8024];
    assign outputs[5863] = ~(layer2_outputs[3422]);
    assign outputs[5864] = ~(layer2_outputs[6170]);
    assign outputs[5865] = ~((layer2_outputs[8083]) ^ (layer2_outputs[12658]));
    assign outputs[5866] = ~(layer2_outputs[4631]) | (layer2_outputs[8749]);
    assign outputs[5867] = (layer2_outputs[8794]) ^ (layer2_outputs[3091]);
    assign outputs[5868] = ~((layer2_outputs[1178]) ^ (layer2_outputs[9701]));
    assign outputs[5869] = layer2_outputs[3473];
    assign outputs[5870] = ~((layer2_outputs[2142]) & (layer2_outputs[6564]));
    assign outputs[5871] = ~(layer2_outputs[564]);
    assign outputs[5872] = layer2_outputs[2294];
    assign outputs[5873] = (layer2_outputs[166]) | (layer2_outputs[2783]);
    assign outputs[5874] = (layer2_outputs[4005]) ^ (layer2_outputs[12453]);
    assign outputs[5875] = layer2_outputs[3562];
    assign outputs[5876] = ~(layer2_outputs[9515]);
    assign outputs[5877] = layer2_outputs[3];
    assign outputs[5878] = layer2_outputs[5806];
    assign outputs[5879] = ~(layer2_outputs[6950]) | (layer2_outputs[8543]);
    assign outputs[5880] = ~(layer2_outputs[8464]);
    assign outputs[5881] = ~(layer2_outputs[5579]) | (layer2_outputs[8673]);
    assign outputs[5882] = layer2_outputs[4745];
    assign outputs[5883] = ~(layer2_outputs[11520]);
    assign outputs[5884] = ~(layer2_outputs[3284]);
    assign outputs[5885] = ~(layer2_outputs[5769]);
    assign outputs[5886] = ~(layer2_outputs[12698]);
    assign outputs[5887] = layer2_outputs[12515];
    assign outputs[5888] = (layer2_outputs[6080]) & ~(layer2_outputs[2565]);
    assign outputs[5889] = ~((layer2_outputs[11471]) ^ (layer2_outputs[9978]));
    assign outputs[5890] = ~((layer2_outputs[12074]) ^ (layer2_outputs[2570]));
    assign outputs[5891] = ~((layer2_outputs[8644]) ^ (layer2_outputs[584]));
    assign outputs[5892] = ~((layer2_outputs[6147]) ^ (layer2_outputs[4151]));
    assign outputs[5893] = ~((layer2_outputs[12572]) ^ (layer2_outputs[11234]));
    assign outputs[5894] = ~(layer2_outputs[9249]) | (layer2_outputs[6501]);
    assign outputs[5895] = ~(layer2_outputs[10696]);
    assign outputs[5896] = ~(layer2_outputs[12670]);
    assign outputs[5897] = (layer2_outputs[9007]) & ~(layer2_outputs[2277]);
    assign outputs[5898] = (layer2_outputs[7171]) | (layer2_outputs[1724]);
    assign outputs[5899] = ~(layer2_outputs[1318]) | (layer2_outputs[381]);
    assign outputs[5900] = layer2_outputs[11341];
    assign outputs[5901] = layer2_outputs[7030];
    assign outputs[5902] = ~((layer2_outputs[7817]) | (layer2_outputs[6363]));
    assign outputs[5903] = layer2_outputs[6418];
    assign outputs[5904] = ~(layer2_outputs[10763]);
    assign outputs[5905] = (layer2_outputs[5854]) ^ (layer2_outputs[7140]);
    assign outputs[5906] = layer2_outputs[662];
    assign outputs[5907] = ~(layer2_outputs[12311]);
    assign outputs[5908] = layer2_outputs[9750];
    assign outputs[5909] = (layer2_outputs[8196]) ^ (layer2_outputs[12508]);
    assign outputs[5910] = (layer2_outputs[5000]) & ~(layer2_outputs[6153]);
    assign outputs[5911] = layer2_outputs[277];
    assign outputs[5912] = (layer2_outputs[9754]) & ~(layer2_outputs[2925]);
    assign outputs[5913] = (layer2_outputs[1]) ^ (layer2_outputs[10838]);
    assign outputs[5914] = layer2_outputs[1178];
    assign outputs[5915] = (layer2_outputs[9756]) & ~(layer2_outputs[1643]);
    assign outputs[5916] = layer2_outputs[5435];
    assign outputs[5917] = ~((layer2_outputs[443]) ^ (layer2_outputs[1253]));
    assign outputs[5918] = (layer2_outputs[3412]) ^ (layer2_outputs[6662]);
    assign outputs[5919] = layer2_outputs[35];
    assign outputs[5920] = layer2_outputs[2479];
    assign outputs[5921] = layer2_outputs[6652];
    assign outputs[5922] = layer2_outputs[5214];
    assign outputs[5923] = (layer2_outputs[7974]) ^ (layer2_outputs[2588]);
    assign outputs[5924] = ~(layer2_outputs[494]);
    assign outputs[5925] = ~(layer2_outputs[3594]);
    assign outputs[5926] = ~(layer2_outputs[271]) | (layer2_outputs[2146]);
    assign outputs[5927] = layer2_outputs[6760];
    assign outputs[5928] = ~(layer2_outputs[8170]);
    assign outputs[5929] = ~((layer2_outputs[10451]) ^ (layer2_outputs[11181]));
    assign outputs[5930] = ~(layer2_outputs[8253]) | (layer2_outputs[3445]);
    assign outputs[5931] = layer2_outputs[11726];
    assign outputs[5932] = ~(layer2_outputs[12657]);
    assign outputs[5933] = layer2_outputs[12124];
    assign outputs[5934] = layer2_outputs[9094];
    assign outputs[5935] = layer2_outputs[5494];
    assign outputs[5936] = (layer2_outputs[6399]) | (layer2_outputs[9437]);
    assign outputs[5937] = layer2_outputs[9411];
    assign outputs[5938] = ~(layer2_outputs[367]) | (layer2_outputs[4752]);
    assign outputs[5939] = ~((layer2_outputs[4146]) ^ (layer2_outputs[3356]));
    assign outputs[5940] = ~((layer2_outputs[9416]) ^ (layer2_outputs[10454]));
    assign outputs[5941] = (layer2_outputs[6462]) & ~(layer2_outputs[4527]);
    assign outputs[5942] = ~(layer2_outputs[1132]);
    assign outputs[5943] = ~((layer2_outputs[10318]) ^ (layer2_outputs[3867]));
    assign outputs[5944] = ~(layer2_outputs[2342]);
    assign outputs[5945] = ~(layer2_outputs[4748]);
    assign outputs[5946] = layer2_outputs[7132];
    assign outputs[5947] = layer2_outputs[2956];
    assign outputs[5948] = layer2_outputs[6549];
    assign outputs[5949] = ~((layer2_outputs[93]) | (layer2_outputs[8485]));
    assign outputs[5950] = ~((layer2_outputs[6366]) ^ (layer2_outputs[7870]));
    assign outputs[5951] = layer2_outputs[10918];
    assign outputs[5952] = (layer2_outputs[228]) & ~(layer2_outputs[7137]);
    assign outputs[5953] = ~(layer2_outputs[7928]);
    assign outputs[5954] = (layer2_outputs[2424]) & ~(layer2_outputs[957]);
    assign outputs[5955] = ~((layer2_outputs[9309]) ^ (layer2_outputs[3404]));
    assign outputs[5956] = ~(layer2_outputs[2675]);
    assign outputs[5957] = (layer2_outputs[606]) | (layer2_outputs[12360]);
    assign outputs[5958] = ~(layer2_outputs[340]);
    assign outputs[5959] = ~(layer2_outputs[7543]);
    assign outputs[5960] = ~(layer2_outputs[4131]);
    assign outputs[5961] = layer2_outputs[794];
    assign outputs[5962] = (layer2_outputs[832]) ^ (layer2_outputs[10830]);
    assign outputs[5963] = layer2_outputs[10466];
    assign outputs[5964] = layer2_outputs[9893];
    assign outputs[5965] = ~((layer2_outputs[1219]) ^ (layer2_outputs[9669]));
    assign outputs[5966] = ~((layer2_outputs[10861]) ^ (layer2_outputs[9549]));
    assign outputs[5967] = layer2_outputs[9915];
    assign outputs[5968] = ~((layer2_outputs[12145]) ^ (layer2_outputs[7327]));
    assign outputs[5969] = (layer2_outputs[205]) ^ (layer2_outputs[7238]);
    assign outputs[5970] = layer2_outputs[7215];
    assign outputs[5971] = ~((layer2_outputs[5502]) & (layer2_outputs[10878]));
    assign outputs[5972] = (layer2_outputs[4298]) ^ (layer2_outputs[7564]);
    assign outputs[5973] = layer2_outputs[11584];
    assign outputs[5974] = ~((layer2_outputs[4129]) ^ (layer2_outputs[4967]));
    assign outputs[5975] = layer2_outputs[6782];
    assign outputs[5976] = ~(layer2_outputs[9403]);
    assign outputs[5977] = ~(layer2_outputs[2017]);
    assign outputs[5978] = ~(layer2_outputs[1964]);
    assign outputs[5979] = ~((layer2_outputs[12059]) ^ (layer2_outputs[1534]));
    assign outputs[5980] = ~(layer2_outputs[10267]);
    assign outputs[5981] = ~(layer2_outputs[11402]);
    assign outputs[5982] = ~(layer2_outputs[8750]);
    assign outputs[5983] = ~(layer2_outputs[4033]);
    assign outputs[5984] = layer2_outputs[11693];
    assign outputs[5985] = ~(layer2_outputs[8974]) | (layer2_outputs[5001]);
    assign outputs[5986] = ~((layer2_outputs[4428]) ^ (layer2_outputs[5582]));
    assign outputs[5987] = (layer2_outputs[4921]) ^ (layer2_outputs[9525]);
    assign outputs[5988] = layer2_outputs[11349];
    assign outputs[5989] = (layer2_outputs[1087]) ^ (layer2_outputs[158]);
    assign outputs[5990] = layer2_outputs[6878];
    assign outputs[5991] = ~((layer2_outputs[9304]) ^ (layer2_outputs[9588]));
    assign outputs[5992] = (layer2_outputs[10146]) & ~(layer2_outputs[8488]);
    assign outputs[5993] = (layer2_outputs[4004]) & ~(layer2_outputs[4642]);
    assign outputs[5994] = ~(layer2_outputs[5173]);
    assign outputs[5995] = layer2_outputs[8135];
    assign outputs[5996] = ~(layer2_outputs[9946]);
    assign outputs[5997] = ~(layer2_outputs[9728]) | (layer2_outputs[429]);
    assign outputs[5998] = layer2_outputs[6361];
    assign outputs[5999] = ~(layer2_outputs[6811]);
    assign outputs[6000] = layer2_outputs[9467];
    assign outputs[6001] = ~(layer2_outputs[7708]);
    assign outputs[6002] = layer2_outputs[6148];
    assign outputs[6003] = layer2_outputs[6771];
    assign outputs[6004] = (layer2_outputs[913]) & ~(layer2_outputs[7791]);
    assign outputs[6005] = (layer2_outputs[2506]) ^ (layer2_outputs[10103]);
    assign outputs[6006] = ~(layer2_outputs[5264]);
    assign outputs[6007] = ~((layer2_outputs[3189]) ^ (layer2_outputs[4638]));
    assign outputs[6008] = layer2_outputs[4855];
    assign outputs[6009] = layer2_outputs[12488];
    assign outputs[6010] = ~(layer2_outputs[1001]);
    assign outputs[6011] = layer2_outputs[49];
    assign outputs[6012] = ~(layer2_outputs[1093]);
    assign outputs[6013] = layer2_outputs[6458];
    assign outputs[6014] = (layer2_outputs[12258]) & ~(layer2_outputs[10478]);
    assign outputs[6015] = (layer2_outputs[3887]) ^ (layer2_outputs[547]);
    assign outputs[6016] = ~(layer2_outputs[886]);
    assign outputs[6017] = ~(layer2_outputs[8947]) | (layer2_outputs[2941]);
    assign outputs[6018] = ~(layer2_outputs[9823]);
    assign outputs[6019] = layer2_outputs[12047];
    assign outputs[6020] = ~((layer2_outputs[10969]) ^ (layer2_outputs[8668]));
    assign outputs[6021] = ~(layer2_outputs[10986]);
    assign outputs[6022] = layer2_outputs[7045];
    assign outputs[6023] = layer2_outputs[4956];
    assign outputs[6024] = ~((layer2_outputs[10071]) ^ (layer2_outputs[712]));
    assign outputs[6025] = (layer2_outputs[11313]) ^ (layer2_outputs[10852]);
    assign outputs[6026] = ~(layer2_outputs[3195]);
    assign outputs[6027] = ~(layer2_outputs[3213]);
    assign outputs[6028] = ~(layer2_outputs[1007]);
    assign outputs[6029] = ~(layer2_outputs[10652]);
    assign outputs[6030] = (layer2_outputs[6427]) ^ (layer2_outputs[11732]);
    assign outputs[6031] = ~((layer2_outputs[6020]) | (layer2_outputs[12334]));
    assign outputs[6032] = ~(layer2_outputs[1006]);
    assign outputs[6033] = ~(layer2_outputs[11611]);
    assign outputs[6034] = ~((layer2_outputs[8167]) ^ (layer2_outputs[9907]));
    assign outputs[6035] = layer2_outputs[6589];
    assign outputs[6036] = ~(layer2_outputs[1807]);
    assign outputs[6037] = ~(layer2_outputs[4652]);
    assign outputs[6038] = ~((layer2_outputs[4608]) ^ (layer2_outputs[5555]));
    assign outputs[6039] = layer2_outputs[9380];
    assign outputs[6040] = ~(layer2_outputs[3906]);
    assign outputs[6041] = layer2_outputs[3669];
    assign outputs[6042] = ~(layer2_outputs[8467]);
    assign outputs[6043] = ~((layer2_outputs[4154]) ^ (layer2_outputs[4116]));
    assign outputs[6044] = layer2_outputs[7927];
    assign outputs[6045] = ~((layer2_outputs[7427]) | (layer2_outputs[1570]));
    assign outputs[6046] = ~(layer2_outputs[11771]) | (layer2_outputs[3671]);
    assign outputs[6047] = ~(layer2_outputs[7658]);
    assign outputs[6048] = ~(layer2_outputs[11017]);
    assign outputs[6049] = ~((layer2_outputs[7579]) ^ (layer2_outputs[3913]));
    assign outputs[6050] = (layer2_outputs[11529]) & (layer2_outputs[10520]);
    assign outputs[6051] = ~(layer2_outputs[11133]);
    assign outputs[6052] = layer2_outputs[263];
    assign outputs[6053] = layer2_outputs[7437];
    assign outputs[6054] = layer2_outputs[1982];
    assign outputs[6055] = layer2_outputs[6851];
    assign outputs[6056] = (layer2_outputs[5883]) & (layer2_outputs[9283]);
    assign outputs[6057] = layer2_outputs[12597];
    assign outputs[6058] = ~(layer2_outputs[5032]);
    assign outputs[6059] = (layer2_outputs[145]) ^ (layer2_outputs[12270]);
    assign outputs[6060] = ~((layer2_outputs[1282]) ^ (layer2_outputs[1280]));
    assign outputs[6061] = ~(layer2_outputs[590]);
    assign outputs[6062] = ~(layer2_outputs[12716]);
    assign outputs[6063] = (layer2_outputs[10052]) & ~(layer2_outputs[12041]);
    assign outputs[6064] = ~(layer2_outputs[3090]);
    assign outputs[6065] = layer2_outputs[3896];
    assign outputs[6066] = ~(layer2_outputs[1370]);
    assign outputs[6067] = (layer2_outputs[10847]) ^ (layer2_outputs[994]);
    assign outputs[6068] = ~((layer2_outputs[2745]) ^ (layer2_outputs[9549]));
    assign outputs[6069] = ~((layer2_outputs[8931]) ^ (layer2_outputs[7244]));
    assign outputs[6070] = ~((layer2_outputs[9895]) ^ (layer2_outputs[11705]));
    assign outputs[6071] = ~(layer2_outputs[3140]);
    assign outputs[6072] = layer2_outputs[2126];
    assign outputs[6073] = ~(layer2_outputs[2510]);
    assign outputs[6074] = (layer2_outputs[6441]) & ~(layer2_outputs[6814]);
    assign outputs[6075] = layer2_outputs[914];
    assign outputs[6076] = ~((layer2_outputs[6719]) | (layer2_outputs[5682]));
    assign outputs[6077] = ~((layer2_outputs[10939]) ^ (layer2_outputs[11472]));
    assign outputs[6078] = layer2_outputs[388];
    assign outputs[6079] = layer2_outputs[236];
    assign outputs[6080] = ~((layer2_outputs[9883]) ^ (layer2_outputs[7791]));
    assign outputs[6081] = (layer2_outputs[11073]) ^ (layer2_outputs[11068]);
    assign outputs[6082] = layer2_outputs[12288];
    assign outputs[6083] = (layer2_outputs[5554]) ^ (layer2_outputs[154]);
    assign outputs[6084] = ~(layer2_outputs[6090]);
    assign outputs[6085] = (layer2_outputs[5063]) | (layer2_outputs[7350]);
    assign outputs[6086] = ~(layer2_outputs[4646]);
    assign outputs[6087] = (layer2_outputs[741]) ^ (layer2_outputs[7169]);
    assign outputs[6088] = layer2_outputs[3761];
    assign outputs[6089] = layer2_outputs[4333];
    assign outputs[6090] = (layer2_outputs[7360]) ^ (layer2_outputs[12525]);
    assign outputs[6091] = ~(layer2_outputs[6205]);
    assign outputs[6092] = ~(layer2_outputs[845]);
    assign outputs[6093] = layer2_outputs[9315];
    assign outputs[6094] = ~(layer2_outputs[788]);
    assign outputs[6095] = ~((layer2_outputs[5498]) ^ (layer2_outputs[12314]));
    assign outputs[6096] = layer2_outputs[8767];
    assign outputs[6097] = layer2_outputs[5778];
    assign outputs[6098] = ~(layer2_outputs[12271]);
    assign outputs[6099] = layer2_outputs[1565];
    assign outputs[6100] = ~(layer2_outputs[3263]);
    assign outputs[6101] = layer2_outputs[11080];
    assign outputs[6102] = ~(layer2_outputs[68]);
    assign outputs[6103] = layer2_outputs[394];
    assign outputs[6104] = ~(layer2_outputs[7079]);
    assign outputs[6105] = ~(layer2_outputs[4845]);
    assign outputs[6106] = ~(layer2_outputs[499]);
    assign outputs[6107] = ~((layer2_outputs[3526]) ^ (layer2_outputs[10628]));
    assign outputs[6108] = ~(layer2_outputs[1843]);
    assign outputs[6109] = layer2_outputs[8575];
    assign outputs[6110] = (layer2_outputs[3276]) ^ (layer2_outputs[6296]);
    assign outputs[6111] = layer2_outputs[10415];
    assign outputs[6112] = layer2_outputs[12369];
    assign outputs[6113] = ~(layer2_outputs[9309]);
    assign outputs[6114] = ~(layer2_outputs[12682]);
    assign outputs[6115] = ~((layer2_outputs[565]) | (layer2_outputs[515]));
    assign outputs[6116] = ~((layer2_outputs[1994]) ^ (layer2_outputs[1572]));
    assign outputs[6117] = (layer2_outputs[6349]) & ~(layer2_outputs[9223]);
    assign outputs[6118] = ~((layer2_outputs[5117]) ^ (layer2_outputs[5887]));
    assign outputs[6119] = ~((layer2_outputs[5771]) ^ (layer2_outputs[5299]));
    assign outputs[6120] = layer2_outputs[1127];
    assign outputs[6121] = layer2_outputs[8091];
    assign outputs[6122] = (layer2_outputs[8317]) | (layer2_outputs[6434]);
    assign outputs[6123] = ~(layer2_outputs[8594]);
    assign outputs[6124] = (layer2_outputs[7952]) & (layer2_outputs[11679]);
    assign outputs[6125] = ~(layer2_outputs[5927]) | (layer2_outputs[4848]);
    assign outputs[6126] = ~((layer2_outputs[1117]) ^ (layer2_outputs[8614]));
    assign outputs[6127] = ~(layer2_outputs[7446]);
    assign outputs[6128] = layer2_outputs[9370];
    assign outputs[6129] = ~(layer2_outputs[396]);
    assign outputs[6130] = (layer2_outputs[12500]) ^ (layer2_outputs[8071]);
    assign outputs[6131] = ~(layer2_outputs[52]);
    assign outputs[6132] = (layer2_outputs[189]) & (layer2_outputs[9282]);
    assign outputs[6133] = (layer2_outputs[10650]) & ~(layer2_outputs[11603]);
    assign outputs[6134] = (layer2_outputs[4381]) ^ (layer2_outputs[2163]);
    assign outputs[6135] = layer2_outputs[1804];
    assign outputs[6136] = layer2_outputs[3693];
    assign outputs[6137] = ~(layer2_outputs[3330]);
    assign outputs[6138] = ~((layer2_outputs[2039]) & (layer2_outputs[11043]));
    assign outputs[6139] = layer2_outputs[964];
    assign outputs[6140] = (layer2_outputs[321]) & (layer2_outputs[9552]);
    assign outputs[6141] = (layer2_outputs[3783]) ^ (layer2_outputs[9126]);
    assign outputs[6142] = layer2_outputs[6349];
    assign outputs[6143] = (layer2_outputs[5787]) ^ (layer2_outputs[1024]);
    assign outputs[6144] = ~((layer2_outputs[9142]) | (layer2_outputs[6788]));
    assign outputs[6145] = (layer2_outputs[6174]) | (layer2_outputs[567]);
    assign outputs[6146] = ~((layer2_outputs[12037]) | (layer2_outputs[3993]));
    assign outputs[6147] = ~(layer2_outputs[8338]);
    assign outputs[6148] = ~((layer2_outputs[44]) ^ (layer2_outputs[4395]));
    assign outputs[6149] = (layer2_outputs[12208]) ^ (layer2_outputs[209]);
    assign outputs[6150] = ~(layer2_outputs[4108]);
    assign outputs[6151] = (layer2_outputs[4359]) ^ (layer2_outputs[2009]);
    assign outputs[6152] = ~((layer2_outputs[2375]) ^ (layer2_outputs[824]));
    assign outputs[6153] = ~(layer2_outputs[512]);
    assign outputs[6154] = layer2_outputs[6865];
    assign outputs[6155] = (layer2_outputs[3553]) | (layer2_outputs[9049]);
    assign outputs[6156] = ~(layer2_outputs[10526]);
    assign outputs[6157] = layer2_outputs[2571];
    assign outputs[6158] = ~((layer2_outputs[6053]) ^ (layer2_outputs[11142]));
    assign outputs[6159] = ~((layer2_outputs[8419]) | (layer2_outputs[7457]));
    assign outputs[6160] = layer2_outputs[615];
    assign outputs[6161] = ~(layer2_outputs[1431]);
    assign outputs[6162] = layer2_outputs[10299];
    assign outputs[6163] = ~((layer2_outputs[11727]) & (layer2_outputs[12179]));
    assign outputs[6164] = (layer2_outputs[8963]) ^ (layer2_outputs[1660]);
    assign outputs[6165] = ~((layer2_outputs[2547]) ^ (layer2_outputs[7492]));
    assign outputs[6166] = ~(layer2_outputs[673]) | (layer2_outputs[515]);
    assign outputs[6167] = layer2_outputs[4927];
    assign outputs[6168] = ~(layer2_outputs[11979]);
    assign outputs[6169] = (layer2_outputs[12692]) ^ (layer2_outputs[6516]);
    assign outputs[6170] = ~(layer2_outputs[8396]);
    assign outputs[6171] = (layer2_outputs[640]) ^ (layer2_outputs[9831]);
    assign outputs[6172] = ~((layer2_outputs[9931]) & (layer2_outputs[6176]));
    assign outputs[6173] = layer2_outputs[6702];
    assign outputs[6174] = (layer2_outputs[11120]) ^ (layer2_outputs[9776]);
    assign outputs[6175] = ~(layer2_outputs[12477]);
    assign outputs[6176] = (layer2_outputs[1885]) ^ (layer2_outputs[852]);
    assign outputs[6177] = (layer2_outputs[5798]) ^ (layer2_outputs[1149]);
    assign outputs[6178] = ~(layer2_outputs[11281]);
    assign outputs[6179] = (layer2_outputs[1624]) & ~(layer2_outputs[9317]);
    assign outputs[6180] = ~(layer2_outputs[4038]);
    assign outputs[6181] = ~(layer2_outputs[12338]);
    assign outputs[6182] = layer2_outputs[7447];
    assign outputs[6183] = ~(layer2_outputs[2279]);
    assign outputs[6184] = layer2_outputs[9181];
    assign outputs[6185] = (layer2_outputs[12566]) ^ (layer2_outputs[9952]);
    assign outputs[6186] = (layer2_outputs[8168]) & (layer2_outputs[450]);
    assign outputs[6187] = layer2_outputs[4549];
    assign outputs[6188] = ~(layer2_outputs[8570]);
    assign outputs[6189] = layer2_outputs[6132];
    assign outputs[6190] = ~(layer2_outputs[5145]) | (layer2_outputs[2343]);
    assign outputs[6191] = layer2_outputs[5166];
    assign outputs[6192] = ~((layer2_outputs[4801]) ^ (layer2_outputs[8509]));
    assign outputs[6193] = ~(layer2_outputs[3998]);
    assign outputs[6194] = ~((layer2_outputs[6824]) ^ (layer2_outputs[54]));
    assign outputs[6195] = ~((layer2_outputs[4678]) ^ (layer2_outputs[1233]));
    assign outputs[6196] = ~(layer2_outputs[4865]);
    assign outputs[6197] = ~(layer2_outputs[2454]);
    assign outputs[6198] = ~((layer2_outputs[7751]) | (layer2_outputs[7090]));
    assign outputs[6199] = ~(layer2_outputs[6715]);
    assign outputs[6200] = ~(layer2_outputs[11661]);
    assign outputs[6201] = ~(layer2_outputs[5519]);
    assign outputs[6202] = ~(layer2_outputs[5444]) | (layer2_outputs[5358]);
    assign outputs[6203] = (layer2_outputs[11331]) ^ (layer2_outputs[8805]);
    assign outputs[6204] = ~(layer2_outputs[1249]);
    assign outputs[6205] = ~(layer2_outputs[3724]);
    assign outputs[6206] = layer2_outputs[7275];
    assign outputs[6207] = ~(layer2_outputs[4321]);
    assign outputs[6208] = (layer2_outputs[8661]) & (layer2_outputs[8957]);
    assign outputs[6209] = ~((layer2_outputs[561]) ^ (layer2_outputs[5772]));
    assign outputs[6210] = ~(layer2_outputs[652]);
    assign outputs[6211] = layer2_outputs[1206];
    assign outputs[6212] = (layer2_outputs[2125]) ^ (layer2_outputs[12674]);
    assign outputs[6213] = layer2_outputs[11989];
    assign outputs[6214] = layer2_outputs[806];
    assign outputs[6215] = ~(layer2_outputs[11967]);
    assign outputs[6216] = ~(layer2_outputs[847]);
    assign outputs[6217] = ~(layer2_outputs[5565]);
    assign outputs[6218] = (layer2_outputs[8605]) ^ (layer2_outputs[7049]);
    assign outputs[6219] = (layer2_outputs[4813]) ^ (layer2_outputs[4062]);
    assign outputs[6220] = ~(layer2_outputs[6586]);
    assign outputs[6221] = ~((layer2_outputs[4615]) ^ (layer2_outputs[9728]));
    assign outputs[6222] = ~(layer2_outputs[11706]);
    assign outputs[6223] = layer2_outputs[12218];
    assign outputs[6224] = ~(layer2_outputs[6357]);
    assign outputs[6225] = (layer2_outputs[11239]) ^ (layer2_outputs[8178]);
    assign outputs[6226] = layer2_outputs[9353];
    assign outputs[6227] = layer2_outputs[9265];
    assign outputs[6228] = ~(layer2_outputs[6431]);
    assign outputs[6229] = layer2_outputs[4111];
    assign outputs[6230] = layer2_outputs[6203];
    assign outputs[6231] = ~((layer2_outputs[10575]) & (layer2_outputs[4241]));
    assign outputs[6232] = (layer2_outputs[9503]) | (layer2_outputs[3653]);
    assign outputs[6233] = ~(layer2_outputs[4254]);
    assign outputs[6234] = ~(layer2_outputs[11233]);
    assign outputs[6235] = ~(layer2_outputs[11125]);
    assign outputs[6236] = layer2_outputs[1439];
    assign outputs[6237] = ~(layer2_outputs[8063]);
    assign outputs[6238] = ~(layer2_outputs[5418]) | (layer2_outputs[1911]);
    assign outputs[6239] = layer2_outputs[9857];
    assign outputs[6240] = ~((layer2_outputs[10100]) ^ (layer2_outputs[12562]));
    assign outputs[6241] = ~(layer2_outputs[3186]);
    assign outputs[6242] = ~(layer2_outputs[11000]) | (layer2_outputs[2900]);
    assign outputs[6243] = ~(layer2_outputs[10160]);
    assign outputs[6244] = ~((layer2_outputs[160]) | (layer2_outputs[9776]));
    assign outputs[6245] = ~((layer2_outputs[10343]) | (layer2_outputs[4098]));
    assign outputs[6246] = ~(layer2_outputs[8228]);
    assign outputs[6247] = ~(layer2_outputs[6284]);
    assign outputs[6248] = (layer2_outputs[12044]) ^ (layer2_outputs[4489]);
    assign outputs[6249] = (layer2_outputs[5037]) ^ (layer2_outputs[4879]);
    assign outputs[6250] = ~(layer2_outputs[2816]);
    assign outputs[6251] = ~((layer2_outputs[9158]) & (layer2_outputs[6792]));
    assign outputs[6252] = layer2_outputs[2005];
    assign outputs[6253] = layer2_outputs[7587];
    assign outputs[6254] = ~((layer2_outputs[3658]) ^ (layer2_outputs[7946]));
    assign outputs[6255] = (layer2_outputs[5857]) ^ (layer2_outputs[6578]);
    assign outputs[6256] = layer2_outputs[8759];
    assign outputs[6257] = (layer2_outputs[2144]) | (layer2_outputs[6260]);
    assign outputs[6258] = layer2_outputs[7933];
    assign outputs[6259] = ~((layer2_outputs[7436]) ^ (layer2_outputs[410]));
    assign outputs[6260] = ~(layer2_outputs[7359]);
    assign outputs[6261] = ~(layer2_outputs[6326]);
    assign outputs[6262] = layer2_outputs[9457];
    assign outputs[6263] = (layer2_outputs[2558]) ^ (layer2_outputs[10562]);
    assign outputs[6264] = ~((layer2_outputs[4914]) ^ (layer2_outputs[141]));
    assign outputs[6265] = ~(layer2_outputs[4940]);
    assign outputs[6266] = ~((layer2_outputs[968]) ^ (layer2_outputs[5955]));
    assign outputs[6267] = ~(layer2_outputs[10934]);
    assign outputs[6268] = ~(layer2_outputs[8396]);
    assign outputs[6269] = layer2_outputs[6107];
    assign outputs[6270] = layer2_outputs[9057];
    assign outputs[6271] = layer2_outputs[8831];
    assign outputs[6272] = ~(layer2_outputs[6419]) | (layer2_outputs[11675]);
    assign outputs[6273] = (layer2_outputs[2517]) ^ (layer2_outputs[3580]);
    assign outputs[6274] = ~(layer2_outputs[7538]);
    assign outputs[6275] = (layer2_outputs[631]) & ~(layer2_outputs[9626]);
    assign outputs[6276] = ~((layer2_outputs[9258]) ^ (layer2_outputs[11446]));
    assign outputs[6277] = layer2_outputs[11567];
    assign outputs[6278] = ~((layer2_outputs[9612]) & (layer2_outputs[11397]));
    assign outputs[6279] = ~(layer2_outputs[11168]);
    assign outputs[6280] = (layer2_outputs[8953]) & ~(layer2_outputs[11236]);
    assign outputs[6281] = ~(layer2_outputs[5331]);
    assign outputs[6282] = ~(layer2_outputs[9284]);
    assign outputs[6283] = (layer2_outputs[3009]) ^ (layer2_outputs[5712]);
    assign outputs[6284] = layer2_outputs[6770];
    assign outputs[6285] = ~((layer2_outputs[6449]) ^ (layer2_outputs[8592]));
    assign outputs[6286] = layer2_outputs[1108];
    assign outputs[6287] = (layer2_outputs[8435]) ^ (layer2_outputs[552]);
    assign outputs[6288] = (layer2_outputs[10873]) ^ (layer2_outputs[5158]);
    assign outputs[6289] = ~((layer2_outputs[5864]) | (layer2_outputs[2889]));
    assign outputs[6290] = (layer2_outputs[8881]) ^ (layer2_outputs[10063]);
    assign outputs[6291] = ~(layer2_outputs[11286]);
    assign outputs[6292] = layer2_outputs[7673];
    assign outputs[6293] = (layer2_outputs[5600]) ^ (layer2_outputs[3454]);
    assign outputs[6294] = layer2_outputs[2887];
    assign outputs[6295] = ~((layer2_outputs[9663]) ^ (layer2_outputs[10061]));
    assign outputs[6296] = (layer2_outputs[9714]) | (layer2_outputs[3766]);
    assign outputs[6297] = layer2_outputs[10423];
    assign outputs[6298] = (layer2_outputs[12361]) ^ (layer2_outputs[9039]);
    assign outputs[6299] = layer2_outputs[5063];
    assign outputs[6300] = ~(layer2_outputs[5236]);
    assign outputs[6301] = layer2_outputs[6961];
    assign outputs[6302] = (layer2_outputs[11381]) ^ (layer2_outputs[6533]);
    assign outputs[6303] = layer2_outputs[5176];
    assign outputs[6304] = ~(layer2_outputs[3517]);
    assign outputs[6305] = ~(layer2_outputs[11890]);
    assign outputs[6306] = ~(layer2_outputs[9635]);
    assign outputs[6307] = ~(layer2_outputs[1445]);
    assign outputs[6308] = ~(layer2_outputs[47]);
    assign outputs[6309] = (layer2_outputs[12272]) | (layer2_outputs[7315]);
    assign outputs[6310] = ~((layer2_outputs[6657]) ^ (layer2_outputs[6747]));
    assign outputs[6311] = layer2_outputs[9716];
    assign outputs[6312] = ~(layer2_outputs[9295]);
    assign outputs[6313] = layer2_outputs[3992];
    assign outputs[6314] = ~((layer2_outputs[11697]) ^ (layer2_outputs[5825]));
    assign outputs[6315] = ~((layer2_outputs[1950]) ^ (layer2_outputs[2864]));
    assign outputs[6316] = ~(layer2_outputs[1036]);
    assign outputs[6317] = layer2_outputs[11954];
    assign outputs[6318] = ~((layer2_outputs[10352]) ^ (layer2_outputs[6122]));
    assign outputs[6319] = ~(layer2_outputs[8353]);
    assign outputs[6320] = ~((layer2_outputs[7455]) | (layer2_outputs[9025]));
    assign outputs[6321] = (layer2_outputs[3084]) ^ (layer2_outputs[10653]);
    assign outputs[6322] = (layer2_outputs[5945]) ^ (layer2_outputs[3042]);
    assign outputs[6323] = layer2_outputs[5438];
    assign outputs[6324] = ~(layer2_outputs[5488]) | (layer2_outputs[8978]);
    assign outputs[6325] = layer2_outputs[5633];
    assign outputs[6326] = ~(layer2_outputs[644]);
    assign outputs[6327] = layer2_outputs[8037];
    assign outputs[6328] = layer2_outputs[5352];
    assign outputs[6329] = layer2_outputs[12489];
    assign outputs[6330] = (layer2_outputs[5092]) & ~(layer2_outputs[11659]);
    assign outputs[6331] = ~((layer2_outputs[7401]) ^ (layer2_outputs[7011]));
    assign outputs[6332] = ~((layer2_outputs[893]) ^ (layer2_outputs[8592]));
    assign outputs[6333] = ~((layer2_outputs[4165]) ^ (layer2_outputs[2766]));
    assign outputs[6334] = ~(layer2_outputs[4764]);
    assign outputs[6335] = ~(layer2_outputs[3339]);
    assign outputs[6336] = ~(layer2_outputs[9163]);
    assign outputs[6337] = (layer2_outputs[2311]) ^ (layer2_outputs[2028]);
    assign outputs[6338] = ~(layer2_outputs[4355]);
    assign outputs[6339] = ~(layer2_outputs[10956]);
    assign outputs[6340] = (layer2_outputs[7667]) & ~(layer2_outputs[1657]);
    assign outputs[6341] = layer2_outputs[1818];
    assign outputs[6342] = ~((layer2_outputs[5569]) ^ (layer2_outputs[4291]));
    assign outputs[6343] = ~(layer2_outputs[66]);
    assign outputs[6344] = ~(layer2_outputs[1015]);
    assign outputs[6345] = ~((layer2_outputs[10030]) ^ (layer2_outputs[7622]));
    assign outputs[6346] = (layer2_outputs[3413]) ^ (layer2_outputs[2304]);
    assign outputs[6347] = ~(layer2_outputs[1014]);
    assign outputs[6348] = (layer2_outputs[5608]) ^ (layer2_outputs[2433]);
    assign outputs[6349] = ~(layer2_outputs[6765]);
    assign outputs[6350] = layer2_outputs[7338];
    assign outputs[6351] = (layer2_outputs[4335]) & (layer2_outputs[8646]);
    assign outputs[6352] = ~(layer2_outputs[1934]);
    assign outputs[6353] = ~(layer2_outputs[5623]);
    assign outputs[6354] = ~(layer2_outputs[12438]);
    assign outputs[6355] = (layer2_outputs[4690]) ^ (layer2_outputs[11368]);
    assign outputs[6356] = ~((layer2_outputs[6663]) ^ (layer2_outputs[5516]));
    assign outputs[6357] = ~(layer2_outputs[10963]);
    assign outputs[6358] = (layer2_outputs[12134]) ^ (layer2_outputs[9091]);
    assign outputs[6359] = ~(layer2_outputs[5613]) | (layer2_outputs[3233]);
    assign outputs[6360] = layer2_outputs[4710];
    assign outputs[6361] = layer2_outputs[6660];
    assign outputs[6362] = ~(layer2_outputs[4068]);
    assign outputs[6363] = layer2_outputs[7804];
    assign outputs[6364] = layer2_outputs[5748];
    assign outputs[6365] = ~((layer2_outputs[11408]) ^ (layer2_outputs[11172]));
    assign outputs[6366] = ~(layer2_outputs[10464]);
    assign outputs[6367] = layer2_outputs[2425];
    assign outputs[6368] = ~(layer2_outputs[6731]);
    assign outputs[6369] = ~(layer2_outputs[6276]);
    assign outputs[6370] = ~(layer2_outputs[1081]);
    assign outputs[6371] = (layer2_outputs[835]) & ~(layer2_outputs[1783]);
    assign outputs[6372] = layer2_outputs[400];
    assign outputs[6373] = layer2_outputs[6485];
    assign outputs[6374] = layer2_outputs[8900];
    assign outputs[6375] = ~(layer2_outputs[8827]);
    assign outputs[6376] = ~(layer2_outputs[1536]);
    assign outputs[6377] = (layer2_outputs[12734]) ^ (layer2_outputs[7276]);
    assign outputs[6378] = ~(layer2_outputs[1158]);
    assign outputs[6379] = layer2_outputs[4495];
    assign outputs[6380] = (layer2_outputs[9875]) ^ (layer2_outputs[12154]);
    assign outputs[6381] = layer2_outputs[2246];
    assign outputs[6382] = (layer2_outputs[4753]) | (layer2_outputs[12647]);
    assign outputs[6383] = ~((layer2_outputs[10564]) ^ (layer2_outputs[11296]));
    assign outputs[6384] = layer2_outputs[3803];
    assign outputs[6385] = layer2_outputs[7061];
    assign outputs[6386] = layer2_outputs[1169];
    assign outputs[6387] = ~((layer2_outputs[9484]) ^ (layer2_outputs[3930]));
    assign outputs[6388] = ~(layer2_outputs[2991]);
    assign outputs[6389] = layer2_outputs[10913];
    assign outputs[6390] = layer2_outputs[8832];
    assign outputs[6391] = layer2_outputs[5103];
    assign outputs[6392] = ~(layer2_outputs[12184]) | (layer2_outputs[12270]);
    assign outputs[6393] = ~(layer2_outputs[1308]);
    assign outputs[6394] = ~((layer2_outputs[7853]) ^ (layer2_outputs[3869]));
    assign outputs[6395] = layer2_outputs[11826];
    assign outputs[6396] = (layer2_outputs[11448]) & ~(layer2_outputs[5837]);
    assign outputs[6397] = ~(layer2_outputs[6840]);
    assign outputs[6398] = ~((layer2_outputs[9559]) | (layer2_outputs[5252]));
    assign outputs[6399] = ~((layer2_outputs[1763]) ^ (layer2_outputs[1450]));
    assign outputs[6400] = layer2_outputs[2104];
    assign outputs[6401] = (layer2_outputs[9557]) | (layer2_outputs[105]);
    assign outputs[6402] = ~(layer2_outputs[12415]);
    assign outputs[6403] = layer2_outputs[8565];
    assign outputs[6404] = layer2_outputs[4686];
    assign outputs[6405] = layer2_outputs[9317];
    assign outputs[6406] = ~((layer2_outputs[11857]) & (layer2_outputs[7050]));
    assign outputs[6407] = (layer2_outputs[4325]) ^ (layer2_outputs[5371]);
    assign outputs[6408] = ~(layer2_outputs[7410]);
    assign outputs[6409] = layer2_outputs[1382];
    assign outputs[6410] = ~((layer2_outputs[10852]) ^ (layer2_outputs[11970]));
    assign outputs[6411] = ~(layer2_outputs[2054]);
    assign outputs[6412] = layer2_outputs[8161];
    assign outputs[6413] = ~(layer2_outputs[12226]);
    assign outputs[6414] = ~((layer2_outputs[12340]) ^ (layer2_outputs[7630]));
    assign outputs[6415] = ~(layer2_outputs[11192]);
    assign outputs[6416] = ~((layer2_outputs[12189]) ^ (layer2_outputs[4408]));
    assign outputs[6417] = ~(layer2_outputs[3385]);
    assign outputs[6418] = ~(layer2_outputs[11225]);
    assign outputs[6419] = ~(layer2_outputs[9444]);
    assign outputs[6420] = (layer2_outputs[8006]) ^ (layer2_outputs[8547]);
    assign outputs[6421] = (layer2_outputs[8882]) ^ (layer2_outputs[5386]);
    assign outputs[6422] = ~(layer2_outputs[7467]);
    assign outputs[6423] = layer2_outputs[8990];
    assign outputs[6424] = ~(layer2_outputs[3170]);
    assign outputs[6425] = layer2_outputs[4764];
    assign outputs[6426] = ~((layer2_outputs[873]) | (layer2_outputs[11970]));
    assign outputs[6427] = ~(layer2_outputs[10390]) | (layer2_outputs[8216]);
    assign outputs[6428] = layer2_outputs[974];
    assign outputs[6429] = ~(layer2_outputs[3743]);
    assign outputs[6430] = layer2_outputs[6827];
    assign outputs[6431] = ~(layer2_outputs[10543]);
    assign outputs[6432] = layer2_outputs[11742];
    assign outputs[6433] = ~(layer2_outputs[10800]);
    assign outputs[6434] = ~((layer2_outputs[107]) ^ (layer2_outputs[3160]));
    assign outputs[6435] = layer2_outputs[6796];
    assign outputs[6436] = (layer2_outputs[3592]) & ~(layer2_outputs[3664]);
    assign outputs[6437] = ~((layer2_outputs[1402]) ^ (layer2_outputs[1956]));
    assign outputs[6438] = ~((layer2_outputs[8107]) ^ (layer2_outputs[7450]));
    assign outputs[6439] = ~(layer2_outputs[5822]) | (layer2_outputs[9633]);
    assign outputs[6440] = ~(layer2_outputs[8495]);
    assign outputs[6441] = (layer2_outputs[9114]) & ~(layer2_outputs[1750]);
    assign outputs[6442] = layer2_outputs[9280];
    assign outputs[6443] = ~((layer2_outputs[7500]) & (layer2_outputs[1124]));
    assign outputs[6444] = ~(layer2_outputs[2051]) | (layer2_outputs[3522]);
    assign outputs[6445] = ~(layer2_outputs[2003]);
    assign outputs[6446] = (layer2_outputs[10653]) ^ (layer2_outputs[10457]);
    assign outputs[6447] = ~(layer2_outputs[4632]);
    assign outputs[6448] = (layer2_outputs[5811]) ^ (layer2_outputs[11332]);
    assign outputs[6449] = layer2_outputs[12103];
    assign outputs[6450] = ~((layer2_outputs[8194]) ^ (layer2_outputs[6249]));
    assign outputs[6451] = layer2_outputs[9418];
    assign outputs[6452] = ~(layer2_outputs[9537]);
    assign outputs[6453] = ~(layer2_outputs[11116]);
    assign outputs[6454] = ~(layer2_outputs[2774]);
    assign outputs[6455] = layer2_outputs[8820];
    assign outputs[6456] = layer2_outputs[8321];
    assign outputs[6457] = ~((layer2_outputs[12354]) ^ (layer2_outputs[2617]));
    assign outputs[6458] = layer2_outputs[486];
    assign outputs[6459] = layer2_outputs[7010];
    assign outputs[6460] = (layer2_outputs[5381]) ^ (layer2_outputs[8083]);
    assign outputs[6461] = layer2_outputs[11959];
    assign outputs[6462] = ~(layer2_outputs[4920]);
    assign outputs[6463] = layer2_outputs[2229];
    assign outputs[6464] = layer2_outputs[5279];
    assign outputs[6465] = ~(layer2_outputs[9971]) | (layer2_outputs[10325]);
    assign outputs[6466] = ~((layer2_outputs[2143]) ^ (layer2_outputs[1099]));
    assign outputs[6467] = (layer2_outputs[1416]) & (layer2_outputs[1429]);
    assign outputs[6468] = ~((layer2_outputs[6811]) ^ (layer2_outputs[11868]));
    assign outputs[6469] = ~(layer2_outputs[9575]);
    assign outputs[6470] = layer2_outputs[5892];
    assign outputs[6471] = (layer2_outputs[4417]) ^ (layer2_outputs[501]);
    assign outputs[6472] = ~(layer2_outputs[1494]);
    assign outputs[6473] = (layer2_outputs[6156]) & (layer2_outputs[8313]);
    assign outputs[6474] = ~(layer2_outputs[3779]);
    assign outputs[6475] = ~((layer2_outputs[9162]) ^ (layer2_outputs[10502]));
    assign outputs[6476] = layer2_outputs[5423];
    assign outputs[6477] = (layer2_outputs[9574]) ^ (layer2_outputs[10604]);
    assign outputs[6478] = (layer2_outputs[8379]) ^ (layer2_outputs[12702]);
    assign outputs[6479] = layer2_outputs[908];
    assign outputs[6480] = ~(layer2_outputs[12126]);
    assign outputs[6481] = layer2_outputs[669];
    assign outputs[6482] = ~(layer2_outputs[2514]);
    assign outputs[6483] = ~((layer2_outputs[3830]) ^ (layer2_outputs[11925]));
    assign outputs[6484] = (layer2_outputs[10869]) | (layer2_outputs[5478]);
    assign outputs[6485] = (layer2_outputs[6617]) ^ (layer2_outputs[7716]);
    assign outputs[6486] = ~(layer2_outputs[281]) | (layer2_outputs[11389]);
    assign outputs[6487] = layer2_outputs[11490];
    assign outputs[6488] = ~(layer2_outputs[10379]);
    assign outputs[6489] = layer2_outputs[9043];
    assign outputs[6490] = ~((layer2_outputs[2274]) ^ (layer2_outputs[2]));
    assign outputs[6491] = ~(layer2_outputs[11252]);
    assign outputs[6492] = layer2_outputs[3382];
    assign outputs[6493] = ~(layer2_outputs[12040]);
    assign outputs[6494] = layer2_outputs[1628];
    assign outputs[6495] = ~((layer2_outputs[2392]) ^ (layer2_outputs[1817]));
    assign outputs[6496] = layer2_outputs[9274];
    assign outputs[6497] = ~((layer2_outputs[8021]) & (layer2_outputs[6925]));
    assign outputs[6498] = ~(layer2_outputs[12586]);
    assign outputs[6499] = (layer2_outputs[11781]) & ~(layer2_outputs[5911]);
    assign outputs[6500] = ~(layer2_outputs[3795]);
    assign outputs[6501] = ~(layer2_outputs[8686]);
    assign outputs[6502] = layer2_outputs[1512];
    assign outputs[6503] = ~((layer2_outputs[12170]) ^ (layer2_outputs[1468]));
    assign outputs[6504] = (layer2_outputs[3777]) & ~(layer2_outputs[5130]);
    assign outputs[6505] = layer2_outputs[4936];
    assign outputs[6506] = ~((layer2_outputs[1605]) ^ (layer2_outputs[9545]));
    assign outputs[6507] = layer2_outputs[7190];
    assign outputs[6508] = layer2_outputs[2199];
    assign outputs[6509] = layer2_outputs[1661];
    assign outputs[6510] = layer2_outputs[315];
    assign outputs[6511] = layer2_outputs[6823];
    assign outputs[6512] = layer2_outputs[4313];
    assign outputs[6513] = (layer2_outputs[3299]) ^ (layer2_outputs[2040]);
    assign outputs[6514] = (layer2_outputs[7903]) & ~(layer2_outputs[7329]);
    assign outputs[6515] = ~((layer2_outputs[4996]) & (layer2_outputs[9665]));
    assign outputs[6516] = layer2_outputs[11095];
    assign outputs[6517] = layer2_outputs[6316];
    assign outputs[6518] = ~((layer2_outputs[10622]) ^ (layer2_outputs[1456]));
    assign outputs[6519] = ~(layer2_outputs[6382]);
    assign outputs[6520] = ~((layer2_outputs[8390]) ^ (layer2_outputs[5027]));
    assign outputs[6521] = ~(layer2_outputs[7329]);
    assign outputs[6522] = layer2_outputs[6833];
    assign outputs[6523] = ~(layer2_outputs[11164]);
    assign outputs[6524] = ~((layer2_outputs[5148]) ^ (layer2_outputs[7181]));
    assign outputs[6525] = ~((layer2_outputs[4146]) ^ (layer2_outputs[1000]));
    assign outputs[6526] = layer2_outputs[6223];
    assign outputs[6527] = (layer2_outputs[10364]) | (layer2_outputs[8094]);
    assign outputs[6528] = ~(layer2_outputs[10507]);
    assign outputs[6529] = ~(layer2_outputs[10025]) | (layer2_outputs[4391]);
    assign outputs[6530] = ~(layer2_outputs[8817]) | (layer2_outputs[11251]);
    assign outputs[6531] = ~((layer2_outputs[10829]) ^ (layer2_outputs[3769]));
    assign outputs[6532] = ~(layer2_outputs[9167]);
    assign outputs[6533] = ~((layer2_outputs[3855]) ^ (layer2_outputs[9852]));
    assign outputs[6534] = layer2_outputs[3241];
    assign outputs[6535] = (layer2_outputs[2063]) & (layer2_outputs[10932]);
    assign outputs[6536] = ~((layer2_outputs[3450]) ^ (layer2_outputs[4402]));
    assign outputs[6537] = ~((layer2_outputs[4487]) ^ (layer2_outputs[845]));
    assign outputs[6538] = ~(layer2_outputs[5012]);
    assign outputs[6539] = layer2_outputs[1102];
    assign outputs[6540] = (layer2_outputs[5697]) ^ (layer2_outputs[4046]);
    assign outputs[6541] = layer2_outputs[8889];
    assign outputs[6542] = ~(layer2_outputs[2027]);
    assign outputs[6543] = (layer2_outputs[3288]) ^ (layer2_outputs[5813]);
    assign outputs[6544] = (layer2_outputs[3836]) & ~(layer2_outputs[6071]);
    assign outputs[6545] = ~(layer2_outputs[11869]) | (layer2_outputs[7058]);
    assign outputs[6546] = layer2_outputs[7367];
    assign outputs[6547] = layer2_outputs[245];
    assign outputs[6548] = ~(layer2_outputs[2774]);
    assign outputs[6549] = (layer2_outputs[1027]) ^ (layer2_outputs[12721]);
    assign outputs[6550] = layer2_outputs[654];
    assign outputs[6551] = ~(layer2_outputs[1910]);
    assign outputs[6552] = (layer2_outputs[2238]) ^ (layer2_outputs[12484]);
    assign outputs[6553] = layer2_outputs[1121];
    assign outputs[6554] = ~(layer2_outputs[7341]);
    assign outputs[6555] = (layer2_outputs[5747]) & ~(layer2_outputs[1417]);
    assign outputs[6556] = ~(layer2_outputs[10343]) | (layer2_outputs[9315]);
    assign outputs[6557] = (layer2_outputs[640]) ^ (layer2_outputs[9059]);
    assign outputs[6558] = layer2_outputs[9671];
    assign outputs[6559] = ~(layer2_outputs[8954]);
    assign outputs[6560] = ~(layer2_outputs[11482]);
    assign outputs[6561] = ~(layer2_outputs[6327]);
    assign outputs[6562] = ~(layer2_outputs[12024]);
    assign outputs[6563] = ~(layer2_outputs[950]);
    assign outputs[6564] = layer2_outputs[7665];
    assign outputs[6565] = ~(layer2_outputs[1322]);
    assign outputs[6566] = ~(layer2_outputs[3675]);
    assign outputs[6567] = (layer2_outputs[229]) ^ (layer2_outputs[3781]);
    assign outputs[6568] = ~(layer2_outputs[134]);
    assign outputs[6569] = ~(layer2_outputs[9352]) | (layer2_outputs[11114]);
    assign outputs[6570] = layer2_outputs[7232];
    assign outputs[6571] = ~((layer2_outputs[1923]) ^ (layer2_outputs[9227]));
    assign outputs[6572] = ~(layer2_outputs[987]);
    assign outputs[6573] = layer2_outputs[11800];
    assign outputs[6574] = layer2_outputs[10761];
    assign outputs[6575] = ~((layer2_outputs[8547]) ^ (layer2_outputs[10064]));
    assign outputs[6576] = ~(layer2_outputs[1153]) | (layer2_outputs[10310]);
    assign outputs[6577] = layer2_outputs[4262];
    assign outputs[6578] = layer2_outputs[10164];
    assign outputs[6579] = (layer2_outputs[9851]) ^ (layer2_outputs[755]);
    assign outputs[6580] = layer2_outputs[1245];
    assign outputs[6581] = ~(layer2_outputs[1577]);
    assign outputs[6582] = ~((layer2_outputs[5421]) ^ (layer2_outputs[2856]));
    assign outputs[6583] = layer2_outputs[5640];
    assign outputs[6584] = layer2_outputs[5275];
    assign outputs[6585] = (layer2_outputs[1579]) ^ (layer2_outputs[6764]);
    assign outputs[6586] = ~(layer2_outputs[2832]);
    assign outputs[6587] = (layer2_outputs[12737]) ^ (layer2_outputs[9254]);
    assign outputs[6588] = (layer2_outputs[7479]) ^ (layer2_outputs[9396]);
    assign outputs[6589] = layer2_outputs[5301];
    assign outputs[6590] = ~(layer2_outputs[11833]);
    assign outputs[6591] = (layer2_outputs[10094]) & ~(layer2_outputs[4996]);
    assign outputs[6592] = (layer2_outputs[9386]) ^ (layer2_outputs[6734]);
    assign outputs[6593] = (layer2_outputs[7978]) ^ (layer2_outputs[5363]);
    assign outputs[6594] = ~((layer2_outputs[10756]) ^ (layer2_outputs[2144]));
    assign outputs[6595] = ~((layer2_outputs[3126]) ^ (layer2_outputs[605]));
    assign outputs[6596] = layer2_outputs[5738];
    assign outputs[6597] = layer2_outputs[2378];
    assign outputs[6598] = ~(layer2_outputs[10507]);
    assign outputs[6599] = (layer2_outputs[8895]) ^ (layer2_outputs[50]);
    assign outputs[6600] = ~(layer2_outputs[11817]);
    assign outputs[6601] = (layer2_outputs[9113]) ^ (layer2_outputs[3060]);
    assign outputs[6602] = (layer2_outputs[1948]) & ~(layer2_outputs[12159]);
    assign outputs[6603] = layer2_outputs[3472];
    assign outputs[6604] = (layer2_outputs[3347]) ^ (layer2_outputs[868]);
    assign outputs[6605] = (layer2_outputs[5889]) ^ (layer2_outputs[4366]);
    assign outputs[6606] = (layer2_outputs[8424]) & (layer2_outputs[8149]);
    assign outputs[6607] = (layer2_outputs[7206]) ^ (layer2_outputs[1413]);
    assign outputs[6608] = layer2_outputs[4466];
    assign outputs[6609] = layer2_outputs[8425];
    assign outputs[6610] = (layer2_outputs[10108]) ^ (layer2_outputs[3722]);
    assign outputs[6611] = ~(layer2_outputs[6073]);
    assign outputs[6612] = ~(layer2_outputs[12061]);
    assign outputs[6613] = layer2_outputs[10394];
    assign outputs[6614] = layer2_outputs[7001];
    assign outputs[6615] = layer2_outputs[7015];
    assign outputs[6616] = ~(layer2_outputs[6970]);
    assign outputs[6617] = ~((layer2_outputs[10664]) | (layer2_outputs[6075]));
    assign outputs[6618] = layer2_outputs[9532];
    assign outputs[6619] = (layer2_outputs[128]) ^ (layer2_outputs[6260]);
    assign outputs[6620] = ~((layer2_outputs[5535]) | (layer2_outputs[5635]));
    assign outputs[6621] = (layer2_outputs[11919]) | (layer2_outputs[2815]);
    assign outputs[6622] = (layer2_outputs[3370]) & (layer2_outputs[12122]);
    assign outputs[6623] = ~(layer2_outputs[2768]);
    assign outputs[6624] = ~(layer2_outputs[3668]);
    assign outputs[6625] = (layer2_outputs[3460]) ^ (layer2_outputs[6949]);
    assign outputs[6626] = (layer2_outputs[9200]) | (layer2_outputs[11777]);
    assign outputs[6627] = ~(layer2_outputs[4884]);
    assign outputs[6628] = layer2_outputs[9155];
    assign outputs[6629] = (layer2_outputs[12364]) ^ (layer2_outputs[7660]);
    assign outputs[6630] = ~(layer2_outputs[2064]);
    assign outputs[6631] = layer2_outputs[7687];
    assign outputs[6632] = layer2_outputs[9551];
    assign outputs[6633] = ~(layer2_outputs[17]);
    assign outputs[6634] = layer2_outputs[7037];
    assign outputs[6635] = layer2_outputs[11943];
    assign outputs[6636] = (layer2_outputs[7792]) & ~(layer2_outputs[8382]);
    assign outputs[6637] = layer2_outputs[8484];
    assign outputs[6638] = ~(layer2_outputs[3210]) | (layer2_outputs[0]);
    assign outputs[6639] = (layer2_outputs[4506]) & (layer2_outputs[7153]);
    assign outputs[6640] = ~((layer2_outputs[3541]) & (layer2_outputs[2520]));
    assign outputs[6641] = ~((layer2_outputs[9099]) | (layer2_outputs[3289]));
    assign outputs[6642] = layer2_outputs[10860];
    assign outputs[6643] = (layer2_outputs[2595]) ^ (layer2_outputs[7195]);
    assign outputs[6644] = (layer2_outputs[11754]) ^ (layer2_outputs[8993]);
    assign outputs[6645] = ~((layer2_outputs[1135]) ^ (layer2_outputs[6957]));
    assign outputs[6646] = (layer2_outputs[7380]) ^ (layer2_outputs[5390]);
    assign outputs[6647] = ~(layer2_outputs[5416]) | (layer2_outputs[9483]);
    assign outputs[6648] = layer2_outputs[10843];
    assign outputs[6649] = ~(layer2_outputs[1035]);
    assign outputs[6650] = layer2_outputs[4691];
    assign outputs[6651] = ~(layer2_outputs[10033]);
    assign outputs[6652] = ~((layer2_outputs[4485]) & (layer2_outputs[10894]));
    assign outputs[6653] = ~(layer2_outputs[4275]);
    assign outputs[6654] = ~((layer2_outputs[6613]) ^ (layer2_outputs[1360]));
    assign outputs[6655] = layer2_outputs[10223];
    assign outputs[6656] = layer2_outputs[2415];
    assign outputs[6657] = ~(layer2_outputs[10664]);
    assign outputs[6658] = ~(layer2_outputs[2951]);
    assign outputs[6659] = ~(layer2_outputs[3437]);
    assign outputs[6660] = layer2_outputs[7741];
    assign outputs[6661] = ~(layer2_outputs[2643]);
    assign outputs[6662] = layer2_outputs[3904];
    assign outputs[6663] = layer2_outputs[10339];
    assign outputs[6664] = (layer2_outputs[9243]) & (layer2_outputs[5874]);
    assign outputs[6665] = (layer2_outputs[4158]) ^ (layer2_outputs[9173]);
    assign outputs[6666] = ~(layer2_outputs[9849]) | (layer2_outputs[6002]);
    assign outputs[6667] = layer2_outputs[11352];
    assign outputs[6668] = layer2_outputs[867];
    assign outputs[6669] = (layer2_outputs[11718]) ^ (layer2_outputs[6146]);
    assign outputs[6670] = layer2_outputs[9191];
    assign outputs[6671] = layer2_outputs[11451];
    assign outputs[6672] = ~((layer2_outputs[5224]) ^ (layer2_outputs[12305]));
    assign outputs[6673] = ~((layer2_outputs[4183]) | (layer2_outputs[9541]));
    assign outputs[6674] = (layer2_outputs[11536]) ^ (layer2_outputs[3013]);
    assign outputs[6675] = (layer2_outputs[3061]) & ~(layer2_outputs[9294]);
    assign outputs[6676] = (layer2_outputs[11729]) ^ (layer2_outputs[1286]);
    assign outputs[6677] = layer2_outputs[10611];
    assign outputs[6678] = layer2_outputs[2677];
    assign outputs[6679] = layer2_outputs[7862];
    assign outputs[6680] = ~((layer2_outputs[1076]) ^ (layer2_outputs[12707]));
    assign outputs[6681] = ~(layer2_outputs[5228]);
    assign outputs[6682] = ~(layer2_outputs[625]) | (layer2_outputs[9400]);
    assign outputs[6683] = layer2_outputs[3610];
    assign outputs[6684] = (layer2_outputs[7433]) ^ (layer2_outputs[2596]);
    assign outputs[6685] = (layer2_outputs[1983]) & (layer2_outputs[1476]);
    assign outputs[6686] = ~(layer2_outputs[4437]);
    assign outputs[6687] = ~(layer2_outputs[2916]);
    assign outputs[6688] = layer2_outputs[4257];
    assign outputs[6689] = ~((layer2_outputs[15]) ^ (layer2_outputs[3945]));
    assign outputs[6690] = (layer2_outputs[10706]) ^ (layer2_outputs[6901]);
    assign outputs[6691] = ~(layer2_outputs[3400]);
    assign outputs[6692] = ~(layer2_outputs[844]);
    assign outputs[6693] = ~(layer2_outputs[1738]);
    assign outputs[6694] = (layer2_outputs[1711]) & ~(layer2_outputs[12083]);
    assign outputs[6695] = ~(layer2_outputs[5887]);
    assign outputs[6696] = ~((layer2_outputs[12240]) | (layer2_outputs[5477]));
    assign outputs[6697] = layer2_outputs[4229];
    assign outputs[6698] = (layer2_outputs[12436]) & ~(layer2_outputs[9708]);
    assign outputs[6699] = ~(layer2_outputs[12388]);
    assign outputs[6700] = (layer2_outputs[4051]) ^ (layer2_outputs[2941]);
    assign outputs[6701] = (layer2_outputs[6495]) ^ (layer2_outputs[2814]);
    assign outputs[6702] = (layer2_outputs[5789]) ^ (layer2_outputs[3245]);
    assign outputs[6703] = layer2_outputs[4578];
    assign outputs[6704] = ~((layer2_outputs[4836]) ^ (layer2_outputs[1018]));
    assign outputs[6705] = ~(layer2_outputs[5410]);
    assign outputs[6706] = ~(layer2_outputs[2294]);
    assign outputs[6707] = layer2_outputs[9520];
    assign outputs[6708] = ~((layer2_outputs[11071]) & (layer2_outputs[1180]));
    assign outputs[6709] = (layer2_outputs[6152]) ^ (layer2_outputs[11349]);
    assign outputs[6710] = layer2_outputs[9940];
    assign outputs[6711] = (layer2_outputs[6959]) & ~(layer2_outputs[3697]);
    assign outputs[6712] = (layer2_outputs[4342]) ^ (layer2_outputs[4900]);
    assign outputs[6713] = ~((layer2_outputs[4297]) ^ (layer2_outputs[4574]));
    assign outputs[6714] = ~((layer2_outputs[3008]) ^ (layer2_outputs[12350]));
    assign outputs[6715] = ~(layer2_outputs[5475]);
    assign outputs[6716] = (layer2_outputs[3168]) ^ (layer2_outputs[12010]);
    assign outputs[6717] = layer2_outputs[4089];
    assign outputs[6718] = (layer2_outputs[1878]) & ~(layer2_outputs[526]);
    assign outputs[6719] = layer2_outputs[1901];
    assign outputs[6720] = ~((layer2_outputs[8512]) ^ (layer2_outputs[9262]));
    assign outputs[6721] = layer2_outputs[2065];
    assign outputs[6722] = ~(layer2_outputs[10571]);
    assign outputs[6723] = ~((layer2_outputs[3363]) ^ (layer2_outputs[1133]));
    assign outputs[6724] = ~(layer2_outputs[1492]);
    assign outputs[6725] = ~(layer2_outputs[10567]);
    assign outputs[6726] = ~(layer2_outputs[4865]);
    assign outputs[6727] = (layer2_outputs[3338]) | (layer2_outputs[1653]);
    assign outputs[6728] = layer2_outputs[9968];
    assign outputs[6729] = ~((layer2_outputs[11680]) ^ (layer2_outputs[3447]));
    assign outputs[6730] = ~(layer2_outputs[3166]);
    assign outputs[6731] = ~(layer2_outputs[2423]);
    assign outputs[6732] = (layer2_outputs[5882]) & ~(layer2_outputs[12724]);
    assign outputs[6733] = (layer2_outputs[11947]) ^ (layer2_outputs[9726]);
    assign outputs[6734] = layer2_outputs[7892];
    assign outputs[6735] = ~(layer2_outputs[1920]) | (layer2_outputs[5864]);
    assign outputs[6736] = layer2_outputs[3493];
    assign outputs[6737] = (layer2_outputs[1793]) | (layer2_outputs[1281]);
    assign outputs[6738] = layer2_outputs[11206];
    assign outputs[6739] = layer2_outputs[11592];
    assign outputs[6740] = ~(layer2_outputs[7093]);
    assign outputs[6741] = (layer2_outputs[12168]) & ~(layer2_outputs[9565]);
    assign outputs[6742] = ~(layer2_outputs[7533]) | (layer2_outputs[3230]);
    assign outputs[6743] = ~((layer2_outputs[12791]) ^ (layer2_outputs[5132]));
    assign outputs[6744] = ~(layer2_outputs[5471]);
    assign outputs[6745] = layer2_outputs[10420];
    assign outputs[6746] = layer2_outputs[3073];
    assign outputs[6747] = layer2_outputs[1502];
    assign outputs[6748] = (layer2_outputs[3819]) ^ (layer2_outputs[5866]);
    assign outputs[6749] = ~(layer2_outputs[11517]);
    assign outputs[6750] = ~(layer2_outputs[10280]);
    assign outputs[6751] = ~((layer2_outputs[10774]) & (layer2_outputs[7907]));
    assign outputs[6752] = ~(layer2_outputs[6623]);
    assign outputs[6753] = layer2_outputs[3877];
    assign outputs[6754] = ~((layer2_outputs[7028]) ^ (layer2_outputs[9826]));
    assign outputs[6755] = layer2_outputs[2199];
    assign outputs[6756] = ~(layer2_outputs[3323]);
    assign outputs[6757] = layer2_outputs[3017];
    assign outputs[6758] = layer2_outputs[6542];
    assign outputs[6759] = ~(layer2_outputs[333]);
    assign outputs[6760] = (layer2_outputs[2716]) ^ (layer2_outputs[5331]);
    assign outputs[6761] = ~(layer2_outputs[5950]) | (layer2_outputs[7216]);
    assign outputs[6762] = ~((layer2_outputs[329]) ^ (layer2_outputs[5673]));
    assign outputs[6763] = layer2_outputs[8399];
    assign outputs[6764] = (layer2_outputs[1502]) & ~(layer2_outputs[3036]);
    assign outputs[6765] = ~(layer2_outputs[8535]);
    assign outputs[6766] = (layer2_outputs[10082]) | (layer2_outputs[5982]);
    assign outputs[6767] = ~(layer2_outputs[9530]);
    assign outputs[6768] = (layer2_outputs[1737]) ^ (layer2_outputs[3696]);
    assign outputs[6769] = layer2_outputs[5771];
    assign outputs[6770] = ~((layer2_outputs[257]) ^ (layer2_outputs[9909]));
    assign outputs[6771] = (layer2_outputs[3420]) ^ (layer2_outputs[2730]);
    assign outputs[6772] = ~(layer2_outputs[9316]);
    assign outputs[6773] = ~(layer2_outputs[917]);
    assign outputs[6774] = (layer2_outputs[6758]) ^ (layer2_outputs[5378]);
    assign outputs[6775] = ~(layer2_outputs[6695]);
    assign outputs[6776] = ~(layer2_outputs[6574]);
    assign outputs[6777] = (layer2_outputs[9654]) & ~(layer2_outputs[1104]);
    assign outputs[6778] = ~(layer2_outputs[1947]);
    assign outputs[6779] = ~((layer2_outputs[2672]) & (layer2_outputs[2017]));
    assign outputs[6780] = layer2_outputs[10135];
    assign outputs[6781] = (layer2_outputs[8919]) & ~(layer2_outputs[11366]);
    assign outputs[6782] = ~(layer2_outputs[5384]) | (layer2_outputs[3527]);
    assign outputs[6783] = layer2_outputs[9392];
    assign outputs[6784] = (layer2_outputs[10334]) ^ (layer2_outputs[819]);
    assign outputs[6785] = ~(layer2_outputs[7542]);
    assign outputs[6786] = layer2_outputs[6401];
    assign outputs[6787] = ~(layer2_outputs[7952]);
    assign outputs[6788] = ~(layer2_outputs[156]);
    assign outputs[6789] = ~(layer2_outputs[1116]);
    assign outputs[6790] = (layer2_outputs[3883]) ^ (layer2_outputs[11822]);
    assign outputs[6791] = ~(layer2_outputs[6916]);
    assign outputs[6792] = (layer2_outputs[4330]) & ~(layer2_outputs[10329]);
    assign outputs[6793] = (layer2_outputs[12171]) & (layer2_outputs[2879]);
    assign outputs[6794] = ~((layer2_outputs[3956]) ^ (layer2_outputs[1422]));
    assign outputs[6795] = (layer2_outputs[8456]) ^ (layer2_outputs[4030]);
    assign outputs[6796] = (layer2_outputs[8207]) & ~(layer2_outputs[7289]);
    assign outputs[6797] = ~(layer2_outputs[7213]);
    assign outputs[6798] = ~(layer2_outputs[760]);
    assign outputs[6799] = layer2_outputs[4738];
    assign outputs[6800] = layer2_outputs[10788];
    assign outputs[6801] = (layer2_outputs[10591]) & (layer2_outputs[3389]);
    assign outputs[6802] = ~(layer2_outputs[5016]);
    assign outputs[6803] = ~(layer2_outputs[10242]);
    assign outputs[6804] = layer2_outputs[5722];
    assign outputs[6805] = ~(layer2_outputs[7021]) | (layer2_outputs[9735]);
    assign outputs[6806] = layer2_outputs[10483];
    assign outputs[6807] = ~(layer2_outputs[1825]);
    assign outputs[6808] = layer2_outputs[10810];
    assign outputs[6809] = (layer2_outputs[4852]) ^ (layer2_outputs[8745]);
    assign outputs[6810] = ~((layer2_outputs[5848]) ^ (layer2_outputs[3567]));
    assign outputs[6811] = (layer2_outputs[1488]) ^ (layer2_outputs[3500]);
    assign outputs[6812] = ~(layer2_outputs[11842]);
    assign outputs[6813] = (layer2_outputs[2931]) & ~(layer2_outputs[6707]);
    assign outputs[6814] = ~(layer2_outputs[4981]);
    assign outputs[6815] = ~(layer2_outputs[3096]);
    assign outputs[6816] = layer2_outputs[768];
    assign outputs[6817] = ~(layer2_outputs[10751]);
    assign outputs[6818] = ~(layer2_outputs[10939]) | (layer2_outputs[2106]);
    assign outputs[6819] = ~(layer2_outputs[7546]);
    assign outputs[6820] = layer2_outputs[11935];
    assign outputs[6821] = ~((layer2_outputs[6537]) & (layer2_outputs[5637]));
    assign outputs[6822] = (layer2_outputs[11208]) ^ (layer2_outputs[5895]);
    assign outputs[6823] = layer2_outputs[5164];
    assign outputs[6824] = ~(layer2_outputs[10724]) | (layer2_outputs[1208]);
    assign outputs[6825] = layer2_outputs[9351];
    assign outputs[6826] = layer2_outputs[7015];
    assign outputs[6827] = (layer2_outputs[2381]) ^ (layer2_outputs[9306]);
    assign outputs[6828] = ~(layer2_outputs[9460]) | (layer2_outputs[9153]);
    assign outputs[6829] = layer2_outputs[1751];
    assign outputs[6830] = ~((layer2_outputs[6804]) & (layer2_outputs[7979]));
    assign outputs[6831] = ~(layer2_outputs[1378]);
    assign outputs[6832] = (layer2_outputs[3193]) ^ (layer2_outputs[6159]);
    assign outputs[6833] = ~(layer2_outputs[3083]);
    assign outputs[6834] = layer2_outputs[10368];
    assign outputs[6835] = ~((layer2_outputs[1430]) ^ (layer2_outputs[10563]));
    assign outputs[6836] = layer2_outputs[1767];
    assign outputs[6837] = ~(layer2_outputs[9339]) | (layer2_outputs[4784]);
    assign outputs[6838] = ~((layer2_outputs[11432]) ^ (layer2_outputs[1839]));
    assign outputs[6839] = ~(layer2_outputs[12766]);
    assign outputs[6840] = layer2_outputs[10870];
    assign outputs[6841] = ~(layer2_outputs[2204]);
    assign outputs[6842] = layer2_outputs[7944];
    assign outputs[6843] = (layer2_outputs[8994]) ^ (layer2_outputs[7025]);
    assign outputs[6844] = (layer2_outputs[7594]) & ~(layer2_outputs[9237]);
    assign outputs[6845] = ~((layer2_outputs[789]) & (layer2_outputs[1205]));
    assign outputs[6846] = (layer2_outputs[8253]) ^ (layer2_outputs[1789]);
    assign outputs[6847] = (layer2_outputs[5638]) & ~(layer2_outputs[1316]);
    assign outputs[6848] = ~((layer2_outputs[11793]) ^ (layer2_outputs[146]));
    assign outputs[6849] = ~((layer2_outputs[1773]) ^ (layer2_outputs[9159]));
    assign outputs[6850] = ~((layer2_outputs[3101]) & (layer2_outputs[6045]));
    assign outputs[6851] = ~((layer2_outputs[9877]) | (layer2_outputs[1339]));
    assign outputs[6852] = (layer2_outputs[3892]) | (layer2_outputs[6969]);
    assign outputs[6853] = ~(layer2_outputs[10897]);
    assign outputs[6854] = layer2_outputs[4428];
    assign outputs[6855] = ~(layer2_outputs[2441]);
    assign outputs[6856] = layer2_outputs[1017];
    assign outputs[6857] = ~(layer2_outputs[1980]);
    assign outputs[6858] = ~((layer2_outputs[7929]) ^ (layer2_outputs[127]));
    assign outputs[6859] = layer2_outputs[10057];
    assign outputs[6860] = ~((layer2_outputs[5091]) | (layer2_outputs[12068]));
    assign outputs[6861] = layer2_outputs[2162];
    assign outputs[6862] = ~((layer2_outputs[1571]) ^ (layer2_outputs[9412]));
    assign outputs[6863] = ~(layer2_outputs[2514]);
    assign outputs[6864] = ~(layer2_outputs[8609]);
    assign outputs[6865] = (layer2_outputs[7338]) ^ (layer2_outputs[3640]);
    assign outputs[6866] = ~(layer2_outputs[2046]);
    assign outputs[6867] = (layer2_outputs[2105]) & ~(layer2_outputs[1482]);
    assign outputs[6868] = layer2_outputs[12372];
    assign outputs[6869] = ~(layer2_outputs[5418]);
    assign outputs[6870] = ~((layer2_outputs[10338]) ^ (layer2_outputs[839]));
    assign outputs[6871] = ~((layer2_outputs[5361]) ^ (layer2_outputs[4390]));
    assign outputs[6872] = (layer2_outputs[2318]) ^ (layer2_outputs[8720]);
    assign outputs[6873] = ~(layer2_outputs[8979]);
    assign outputs[6874] = (layer2_outputs[8875]) | (layer2_outputs[12511]);
    assign outputs[6875] = (layer2_outputs[4895]) ^ (layer2_outputs[11059]);
    assign outputs[6876] = ~((layer2_outputs[10501]) ^ (layer2_outputs[6034]));
    assign outputs[6877] = ~(layer2_outputs[3541]);
    assign outputs[6878] = ~((layer2_outputs[12684]) ^ (layer2_outputs[9144]));
    assign outputs[6879] = ~(layer2_outputs[10013]);
    assign outputs[6880] = (layer2_outputs[11871]) ^ (layer2_outputs[6872]);
    assign outputs[6881] = layer2_outputs[6556];
    assign outputs[6882] = ~(layer2_outputs[10514]);
    assign outputs[6883] = (layer2_outputs[1698]) ^ (layer2_outputs[8224]);
    assign outputs[6884] = (layer2_outputs[7792]) & ~(layer2_outputs[7719]);
    assign outputs[6885] = ~(layer2_outputs[4543]);
    assign outputs[6886] = ~(layer2_outputs[6799]);
    assign outputs[6887] = (layer2_outputs[11103]) | (layer2_outputs[6175]);
    assign outputs[6888] = (layer2_outputs[6762]) & (layer2_outputs[1532]);
    assign outputs[6889] = layer2_outputs[4600];
    assign outputs[6890] = ~((layer2_outputs[9082]) ^ (layer2_outputs[4581]));
    assign outputs[6891] = ~(layer2_outputs[4973]);
    assign outputs[6892] = ~((layer2_outputs[8137]) ^ (layer2_outputs[8685]));
    assign outputs[6893] = ~((layer2_outputs[5709]) & (layer2_outputs[1157]));
    assign outputs[6894] = ~(layer2_outputs[3562]);
    assign outputs[6895] = layer2_outputs[3275];
    assign outputs[6896] = ~(layer2_outputs[3992]);
    assign outputs[6897] = ~((layer2_outputs[1359]) ^ (layer2_outputs[4963]));
    assign outputs[6898] = layer2_outputs[2228];
    assign outputs[6899] = ~((layer2_outputs[11820]) ^ (layer2_outputs[6568]));
    assign outputs[6900] = ~(layer2_outputs[10581]);
    assign outputs[6901] = ~(layer2_outputs[8188]);
    assign outputs[6902] = layer2_outputs[9679];
    assign outputs[6903] = (layer2_outputs[4126]) ^ (layer2_outputs[12017]);
    assign outputs[6904] = layer2_outputs[1279];
    assign outputs[6905] = (layer2_outputs[5074]) ^ (layer2_outputs[5170]);
    assign outputs[6906] = layer2_outputs[10646];
    assign outputs[6907] = ~((layer2_outputs[715]) ^ (layer2_outputs[1544]));
    assign outputs[6908] = layer2_outputs[8129];
    assign outputs[6909] = layer2_outputs[10786];
    assign outputs[6910] = layer2_outputs[2165];
    assign outputs[6911] = ~(layer2_outputs[9620]);
    assign outputs[6912] = layer2_outputs[9355];
    assign outputs[6913] = layer2_outputs[5684];
    assign outputs[6914] = ~(layer2_outputs[10487]);
    assign outputs[6915] = (layer2_outputs[8141]) & ~(layer2_outputs[5755]);
    assign outputs[6916] = layer2_outputs[6836];
    assign outputs[6917] = (layer2_outputs[1689]) ^ (layer2_outputs[9680]);
    assign outputs[6918] = (layer2_outputs[7412]) ^ (layer2_outputs[10813]);
    assign outputs[6919] = ~((layer2_outputs[6267]) ^ (layer2_outputs[11002]));
    assign outputs[6920] = ~((layer2_outputs[7731]) | (layer2_outputs[522]));
    assign outputs[6921] = ~(layer2_outputs[1639]);
    assign outputs[6922] = ~(layer2_outputs[6482]);
    assign outputs[6923] = ~(layer2_outputs[4943]);
    assign outputs[6924] = (layer2_outputs[3863]) ^ (layer2_outputs[8490]);
    assign outputs[6925] = (layer2_outputs[8112]) & ~(layer2_outputs[6450]);
    assign outputs[6926] = ~((layer2_outputs[827]) & (layer2_outputs[8628]));
    assign outputs[6927] = ~(layer2_outputs[5050]);
    assign outputs[6928] = ~(layer2_outputs[641]);
    assign outputs[6929] = ~((layer2_outputs[1962]) ^ (layer2_outputs[5151]));
    assign outputs[6930] = (layer2_outputs[10730]) ^ (layer2_outputs[9577]);
    assign outputs[6931] = (layer2_outputs[2535]) ^ (layer2_outputs[1477]);
    assign outputs[6932] = layer2_outputs[958];
    assign outputs[6933] = ~(layer2_outputs[1268]);
    assign outputs[6934] = layer2_outputs[3069];
    assign outputs[6935] = (layer2_outputs[12144]) & ~(layer2_outputs[7366]);
    assign outputs[6936] = ~(layer2_outputs[12776]);
    assign outputs[6937] = (layer2_outputs[570]) ^ (layer2_outputs[7660]);
    assign outputs[6938] = layer2_outputs[5985];
    assign outputs[6939] = layer2_outputs[9527];
    assign outputs[6940] = (layer2_outputs[1693]) ^ (layer2_outputs[7102]);
    assign outputs[6941] = (layer2_outputs[61]) ^ (layer2_outputs[2375]);
    assign outputs[6942] = layer2_outputs[8985];
    assign outputs[6943] = layer2_outputs[2344];
    assign outputs[6944] = (layer2_outputs[1249]) | (layer2_outputs[11838]);
    assign outputs[6945] = (layer2_outputs[695]) ^ (layer2_outputs[699]);
    assign outputs[6946] = layer2_outputs[6046];
    assign outputs[6947] = layer2_outputs[2560];
    assign outputs[6948] = layer2_outputs[5305];
    assign outputs[6949] = layer2_outputs[5783];
    assign outputs[6950] = ~((layer2_outputs[4651]) ^ (layer2_outputs[7504]));
    assign outputs[6951] = (layer2_outputs[6021]) | (layer2_outputs[6919]);
    assign outputs[6952] = layer2_outputs[12545];
    assign outputs[6953] = ~(layer2_outputs[2061]) | (layer2_outputs[6664]);
    assign outputs[6954] = ~(layer2_outputs[5181]);
    assign outputs[6955] = layer2_outputs[6223];
    assign outputs[6956] = (layer2_outputs[3376]) ^ (layer2_outputs[1981]);
    assign outputs[6957] = (layer2_outputs[9165]) & ~(layer2_outputs[11525]);
    assign outputs[6958] = ~(layer2_outputs[6312]);
    assign outputs[6959] = layer2_outputs[2315];
    assign outputs[6960] = layer2_outputs[5476];
    assign outputs[6961] = ~(layer2_outputs[2213]);
    assign outputs[6962] = ~(layer2_outputs[2235]);
    assign outputs[6963] = layer2_outputs[11943];
    assign outputs[6964] = ~((layer2_outputs[1119]) ^ (layer2_outputs[3045]));
    assign outputs[6965] = ~(layer2_outputs[3490]);
    assign outputs[6966] = (layer2_outputs[435]) ^ (layer2_outputs[1600]);
    assign outputs[6967] = layer2_outputs[8754];
    assign outputs[6968] = ~(layer2_outputs[7650]);
    assign outputs[6969] = layer2_outputs[4826];
    assign outputs[6970] = ~(layer2_outputs[5295]);
    assign outputs[6971] = layer2_outputs[11428];
    assign outputs[6972] = ~(layer2_outputs[11848]);
    assign outputs[6973] = ~((layer2_outputs[1055]) ^ (layer2_outputs[9028]));
    assign outputs[6974] = layer2_outputs[6468];
    assign outputs[6975] = (layer2_outputs[7717]) ^ (layer2_outputs[1016]);
    assign outputs[6976] = layer2_outputs[8413];
    assign outputs[6977] = ~(layer2_outputs[3295]);
    assign outputs[6978] = ~(layer2_outputs[10479]);
    assign outputs[6979] = ~((layer2_outputs[2129]) & (layer2_outputs[7086]));
    assign outputs[6980] = ~((layer2_outputs[4033]) | (layer2_outputs[12126]));
    assign outputs[6981] = (layer2_outputs[2798]) ^ (layer2_outputs[1917]);
    assign outputs[6982] = ~((layer2_outputs[3001]) | (layer2_outputs[9369]));
    assign outputs[6983] = ~(layer2_outputs[1569]);
    assign outputs[6984] = ~(layer2_outputs[6278]);
    assign outputs[6985] = ~((layer2_outputs[4907]) ^ (layer2_outputs[8705]));
    assign outputs[6986] = ~((layer2_outputs[5038]) & (layer2_outputs[11211]));
    assign outputs[6987] = ~((layer2_outputs[5067]) ^ (layer2_outputs[4511]));
    assign outputs[6988] = layer2_outputs[863];
    assign outputs[6989] = ~((layer2_outputs[11765]) ^ (layer2_outputs[3474]));
    assign outputs[6990] = (layer2_outputs[7670]) & ~(layer2_outputs[979]);
    assign outputs[6991] = ~((layer2_outputs[7166]) ^ (layer2_outputs[6863]));
    assign outputs[6992] = layer2_outputs[2164];
    assign outputs[6993] = layer2_outputs[3564];
    assign outputs[6994] = (layer2_outputs[8180]) ^ (layer2_outputs[7812]);
    assign outputs[6995] = layer2_outputs[2908];
    assign outputs[6996] = layer2_outputs[5404];
    assign outputs[6997] = layer2_outputs[199];
    assign outputs[6998] = ~(layer2_outputs[11041]);
    assign outputs[6999] = ~(layer2_outputs[11869]) | (layer2_outputs[4300]);
    assign outputs[7000] = ~(layer2_outputs[3893]);
    assign outputs[7001] = ~(layer2_outputs[2546]);
    assign outputs[7002] = ~(layer2_outputs[6070]);
    assign outputs[7003] = ~((layer2_outputs[8311]) ^ (layer2_outputs[10211]));
    assign outputs[7004] = ~(layer2_outputs[12056]);
    assign outputs[7005] = (layer2_outputs[8187]) ^ (layer2_outputs[626]);
    assign outputs[7006] = ~((layer2_outputs[10594]) ^ (layer2_outputs[11151]));
    assign outputs[7007] = ~((layer2_outputs[11986]) ^ (layer2_outputs[2106]));
    assign outputs[7008] = ~((layer2_outputs[3466]) & (layer2_outputs[10392]));
    assign outputs[7009] = (layer2_outputs[5300]) & (layer2_outputs[6861]);
    assign outputs[7010] = (layer2_outputs[2735]) | (layer2_outputs[8643]);
    assign outputs[7011] = layer2_outputs[6857];
    assign outputs[7012] = layer2_outputs[7278];
    assign outputs[7013] = (layer2_outputs[7633]) ^ (layer2_outputs[11436]);
    assign outputs[7014] = ~((layer2_outputs[5737]) ^ (layer2_outputs[7486]));
    assign outputs[7015] = layer2_outputs[5262];
    assign outputs[7016] = layer2_outputs[7482];
    assign outputs[7017] = (layer2_outputs[236]) & ~(layer2_outputs[11532]);
    assign outputs[7018] = ~(layer2_outputs[11081]);
    assign outputs[7019] = layer2_outputs[2702];
    assign outputs[7020] = (layer2_outputs[3682]) ^ (layer2_outputs[1712]);
    assign outputs[7021] = ~(layer2_outputs[1284]) | (layer2_outputs[3337]);
    assign outputs[7022] = (layer2_outputs[588]) ^ (layer2_outputs[8799]);
    assign outputs[7023] = ~((layer2_outputs[11075]) | (layer2_outputs[1253]));
    assign outputs[7024] = ~(layer2_outputs[3773]) | (layer2_outputs[11036]);
    assign outputs[7025] = layer2_outputs[6331];
    assign outputs[7026] = layer2_outputs[6325];
    assign outputs[7027] = (layer2_outputs[1769]) | (layer2_outputs[955]);
    assign outputs[7028] = ~(layer2_outputs[10136]);
    assign outputs[7029] = layer2_outputs[5463];
    assign outputs[7030] = layer2_outputs[12591];
    assign outputs[7031] = layer2_outputs[10991];
    assign outputs[7032] = layer2_outputs[12678];
    assign outputs[7033] = (layer2_outputs[3342]) ^ (layer2_outputs[10404]);
    assign outputs[7034] = layer2_outputs[2115];
    assign outputs[7035] = (layer2_outputs[11677]) & ~(layer2_outputs[763]);
    assign outputs[7036] = ~(layer2_outputs[12000]);
    assign outputs[7037] = layer2_outputs[9177];
    assign outputs[7038] = ~((layer2_outputs[11034]) ^ (layer2_outputs[1482]));
    assign outputs[7039] = ~(layer2_outputs[3833]);
    assign outputs[7040] = layer2_outputs[5102];
    assign outputs[7041] = ~(layer2_outputs[9531]);
    assign outputs[7042] = ~(layer2_outputs[3850]);
    assign outputs[7043] = (layer2_outputs[7805]) & ~(layer2_outputs[8690]);
    assign outputs[7044] = layer2_outputs[1383];
    assign outputs[7045] = ~(layer2_outputs[7133]) | (layer2_outputs[9860]);
    assign outputs[7046] = ~((layer2_outputs[6029]) ^ (layer2_outputs[10782]));
    assign outputs[7047] = (layer2_outputs[12346]) ^ (layer2_outputs[1379]);
    assign outputs[7048] = layer2_outputs[2612];
    assign outputs[7049] = layer2_outputs[10792];
    assign outputs[7050] = ~(layer2_outputs[8863]);
    assign outputs[7051] = ~((layer2_outputs[10593]) | (layer2_outputs[11512]));
    assign outputs[7052] = ~((layer2_outputs[5878]) | (layer2_outputs[11436]));
    assign outputs[7053] = (layer2_outputs[1959]) | (layer2_outputs[4963]);
    assign outputs[7054] = ~(layer2_outputs[12542]);
    assign outputs[7055] = ~(layer2_outputs[5899]);
    assign outputs[7056] = layer2_outputs[12396];
    assign outputs[7057] = ~(layer2_outputs[2107]);
    assign outputs[7058] = layer2_outputs[9366];
    assign outputs[7059] = layer2_outputs[4558];
    assign outputs[7060] = layer2_outputs[2237];
    assign outputs[7061] = (layer2_outputs[5053]) & ~(layer2_outputs[10927]);
    assign outputs[7062] = ~((layer2_outputs[5617]) ^ (layer2_outputs[1403]));
    assign outputs[7063] = layer2_outputs[11430];
    assign outputs[7064] = ~(layer2_outputs[1114]);
    assign outputs[7065] = (layer2_outputs[5258]) & (layer2_outputs[12322]);
    assign outputs[7066] = ~((layer2_outputs[9159]) ^ (layer2_outputs[12588]));
    assign outputs[7067] = layer2_outputs[10996];
    assign outputs[7068] = ~((layer2_outputs[11815]) ^ (layer2_outputs[6793]));
    assign outputs[7069] = ~(layer2_outputs[10921]);
    assign outputs[7070] = (layer2_outputs[3525]) & ~(layer2_outputs[11655]);
    assign outputs[7071] = ~(layer2_outputs[12040]);
    assign outputs[7072] = (layer2_outputs[11708]) | (layer2_outputs[5953]);
    assign outputs[7073] = (layer2_outputs[5085]) ^ (layer2_outputs[6739]);
    assign outputs[7074] = (layer2_outputs[3527]) ^ (layer2_outputs[5759]);
    assign outputs[7075] = ~(layer2_outputs[2522]);
    assign outputs[7076] = (layer2_outputs[3282]) ^ (layer2_outputs[9562]);
    assign outputs[7077] = ~(layer2_outputs[4145]);
    assign outputs[7078] = layer2_outputs[9891];
    assign outputs[7079] = layer2_outputs[8689];
    assign outputs[7080] = ~(layer2_outputs[8264]) | (layer2_outputs[9446]);
    assign outputs[7081] = ~(layer2_outputs[9401]);
    assign outputs[7082] = (layer2_outputs[5264]) & (layer2_outputs[2843]);
    assign outputs[7083] = layer2_outputs[4101];
    assign outputs[7084] = ~((layer2_outputs[9802]) ^ (layer2_outputs[2245]));
    assign outputs[7085] = (layer2_outputs[5728]) ^ (layer2_outputs[931]);
    assign outputs[7086] = ~((layer2_outputs[5232]) | (layer2_outputs[11297]));
    assign outputs[7087] = ~(layer2_outputs[10316]);
    assign outputs[7088] = (layer2_outputs[210]) & ~(layer2_outputs[2226]);
    assign outputs[7089] = (layer2_outputs[11433]) ^ (layer2_outputs[10608]);
    assign outputs[7090] = ~(layer2_outputs[2650]);
    assign outputs[7091] = (layer2_outputs[8432]) | (layer2_outputs[8647]);
    assign outputs[7092] = ~(layer2_outputs[270]);
    assign outputs[7093] = ~((layer2_outputs[11183]) ^ (layer2_outputs[1652]));
    assign outputs[7094] = layer2_outputs[3298];
    assign outputs[7095] = layer2_outputs[10857];
    assign outputs[7096] = ~((layer2_outputs[2282]) ^ (layer2_outputs[4248]));
    assign outputs[7097] = ~(layer2_outputs[38]);
    assign outputs[7098] = ~((layer2_outputs[12608]) ^ (layer2_outputs[5902]));
    assign outputs[7099] = ~(layer2_outputs[8731]);
    assign outputs[7100] = ~((layer2_outputs[203]) ^ (layer2_outputs[10361]));
    assign outputs[7101] = ~(layer2_outputs[5160]);
    assign outputs[7102] = (layer2_outputs[3261]) ^ (layer2_outputs[12525]);
    assign outputs[7103] = (layer2_outputs[12537]) ^ (layer2_outputs[7606]);
    assign outputs[7104] = ~((layer2_outputs[1274]) ^ (layer2_outputs[2706]));
    assign outputs[7105] = ~(layer2_outputs[3383]);
    assign outputs[7106] = ~(layer2_outputs[4238]);
    assign outputs[7107] = ~(layer2_outputs[3491]);
    assign outputs[7108] = layer2_outputs[1976];
    assign outputs[7109] = layer2_outputs[7483];
    assign outputs[7110] = (layer2_outputs[751]) ^ (layer2_outputs[4788]);
    assign outputs[7111] = (layer2_outputs[8493]) & (layer2_outputs[10420]);
    assign outputs[7112] = layer2_outputs[10319];
    assign outputs[7113] = (layer2_outputs[10911]) ^ (layer2_outputs[1704]);
    assign outputs[7114] = ~((layer2_outputs[3507]) & (layer2_outputs[10908]));
    assign outputs[7115] = ~((layer2_outputs[7208]) ^ (layer2_outputs[5011]));
    assign outputs[7116] = ~((layer2_outputs[4400]) ^ (layer2_outputs[3285]));
    assign outputs[7117] = ~((layer2_outputs[4628]) ^ (layer2_outputs[10943]));
    assign outputs[7118] = (layer2_outputs[1559]) ^ (layer2_outputs[7574]);
    assign outputs[7119] = (layer2_outputs[3029]) ^ (layer2_outputs[11362]);
    assign outputs[7120] = ~(layer2_outputs[2669]);
    assign outputs[7121] = layer2_outputs[12799];
    assign outputs[7122] = layer2_outputs[12450];
    assign outputs[7123] = ~((layer2_outputs[6309]) ^ (layer2_outputs[5480]));
    assign outputs[7124] = (layer2_outputs[7780]) | (layer2_outputs[523]);
    assign outputs[7125] = ~(layer2_outputs[7981]);
    assign outputs[7126] = ~((layer2_outputs[12469]) ^ (layer2_outputs[10868]));
    assign outputs[7127] = ~(layer2_outputs[6273]);
    assign outputs[7128] = layer2_outputs[1112];
    assign outputs[7129] = layer2_outputs[10798];
    assign outputs[7130] = layer2_outputs[4047];
    assign outputs[7131] = ~(layer2_outputs[2917]);
    assign outputs[7132] = ~((layer2_outputs[4066]) ^ (layer2_outputs[2554]));
    assign outputs[7133] = layer2_outputs[4864];
    assign outputs[7134] = (layer2_outputs[11570]) | (layer2_outputs[6334]);
    assign outputs[7135] = ~(layer2_outputs[5939]);
    assign outputs[7136] = ~(layer2_outputs[10643]);
    assign outputs[7137] = ~(layer2_outputs[10174]);
    assign outputs[7138] = (layer2_outputs[9720]) & ~(layer2_outputs[12626]);
    assign outputs[7139] = ~(layer2_outputs[10126]);
    assign outputs[7140] = layer2_outputs[117];
    assign outputs[7141] = ~((layer2_outputs[9906]) ^ (layer2_outputs[9629]));
    assign outputs[7142] = ~(layer2_outputs[534]);
    assign outputs[7143] = ~((layer2_outputs[3596]) ^ (layer2_outputs[2795]));
    assign outputs[7144] = (layer2_outputs[8795]) & ~(layer2_outputs[12795]);
    assign outputs[7145] = (layer2_outputs[2869]) ^ (layer2_outputs[879]);
    assign outputs[7146] = layer2_outputs[3529];
    assign outputs[7147] = ~(layer2_outputs[9261]);
    assign outputs[7148] = (layer2_outputs[1201]) | (layer2_outputs[1320]);
    assign outputs[7149] = layer2_outputs[7073];
    assign outputs[7150] = (layer2_outputs[595]) & (layer2_outputs[3103]);
    assign outputs[7151] = (layer2_outputs[12285]) & (layer2_outputs[12560]);
    assign outputs[7152] = ~((layer2_outputs[1972]) ^ (layer2_outputs[879]));
    assign outputs[7153] = layer2_outputs[994];
    assign outputs[7154] = (layer2_outputs[4012]) & (layer2_outputs[1925]);
    assign outputs[7155] = ~(layer2_outputs[6115]) | (layer2_outputs[11144]);
    assign outputs[7156] = layer2_outputs[2557];
    assign outputs[7157] = ~(layer2_outputs[9647]);
    assign outputs[7158] = layer2_outputs[773];
    assign outputs[7159] = ~(layer2_outputs[11318]);
    assign outputs[7160] = ~((layer2_outputs[3194]) ^ (layer2_outputs[6504]));
    assign outputs[7161] = layer2_outputs[9429];
    assign outputs[7162] = ~((layer2_outputs[1265]) ^ (layer2_outputs[5624]));
    assign outputs[7163] = layer2_outputs[6021];
    assign outputs[7164] = layer2_outputs[1007];
    assign outputs[7165] = (layer2_outputs[10495]) ^ (layer2_outputs[5419]);
    assign outputs[7166] = layer2_outputs[10028];
    assign outputs[7167] = layer2_outputs[1414];
    assign outputs[7168] = (layer2_outputs[4184]) ^ (layer2_outputs[3943]);
    assign outputs[7169] = ~((layer2_outputs[3394]) ^ (layer2_outputs[5574]));
    assign outputs[7170] = ~(layer2_outputs[681]);
    assign outputs[7171] = layer2_outputs[12617];
    assign outputs[7172] = ~((layer2_outputs[12744]) ^ (layer2_outputs[3278]));
    assign outputs[7173] = ~((layer2_outputs[12262]) & (layer2_outputs[1379]));
    assign outputs[7174] = (layer2_outputs[2486]) | (layer2_outputs[12466]);
    assign outputs[7175] = ~((layer2_outputs[6632]) ^ (layer2_outputs[10678]));
    assign outputs[7176] = ~(layer2_outputs[3437]) | (layer2_outputs[10796]);
    assign outputs[7177] = (layer2_outputs[8976]) ^ (layer2_outputs[12222]);
    assign outputs[7178] = ~(layer2_outputs[6810]);
    assign outputs[7179] = layer2_outputs[5656];
    assign outputs[7180] = ~(layer2_outputs[39]);
    assign outputs[7181] = ~((layer2_outputs[11264]) ^ (layer2_outputs[9595]));
    assign outputs[7182] = layer2_outputs[2915];
    assign outputs[7183] = ~(layer2_outputs[11594]);
    assign outputs[7184] = ~(layer2_outputs[1961]);
    assign outputs[7185] = ~(layer2_outputs[136]);
    assign outputs[7186] = ~((layer2_outputs[7413]) ^ (layer2_outputs[1266]));
    assign outputs[7187] = (layer2_outputs[7200]) ^ (layer2_outputs[2773]);
    assign outputs[7188] = (layer2_outputs[5669]) ^ (layer2_outputs[6689]);
    assign outputs[7189] = layer2_outputs[7541];
    assign outputs[7190] = layer2_outputs[6352];
    assign outputs[7191] = (layer2_outputs[8143]) ^ (layer2_outputs[12250]);
    assign outputs[7192] = ~(layer2_outputs[5350]);
    assign outputs[7193] = (layer2_outputs[5115]) ^ (layer2_outputs[12739]);
    assign outputs[7194] = ~(layer2_outputs[3516]);
    assign outputs[7195] = (layer2_outputs[1272]) ^ (layer2_outputs[7567]);
    assign outputs[7196] = ~((layer2_outputs[11560]) ^ (layer2_outputs[5457]));
    assign outputs[7197] = ~((layer2_outputs[12275]) ^ (layer2_outputs[5585]));
    assign outputs[7198] = layer2_outputs[11248];
    assign outputs[7199] = layer2_outputs[6286];
    assign outputs[7200] = layer2_outputs[2317];
    assign outputs[7201] = ~((layer2_outputs[57]) ^ (layer2_outputs[2594]));
    assign outputs[7202] = (layer2_outputs[8091]) | (layer2_outputs[8082]);
    assign outputs[7203] = layer2_outputs[9903];
    assign outputs[7204] = ~((layer2_outputs[9227]) | (layer2_outputs[11255]));
    assign outputs[7205] = ~(layer2_outputs[1344]);
    assign outputs[7206] = (layer2_outputs[2965]) ^ (layer2_outputs[5544]);
    assign outputs[7207] = ~((layer2_outputs[11880]) | (layer2_outputs[8617]));
    assign outputs[7208] = ~((layer2_outputs[1078]) ^ (layer2_outputs[10199]));
    assign outputs[7209] = ~(layer2_outputs[6928]);
    assign outputs[7210] = (layer2_outputs[11067]) | (layer2_outputs[3929]);
    assign outputs[7211] = layer2_outputs[171];
    assign outputs[7212] = ~(layer2_outputs[12243]);
    assign outputs[7213] = (layer2_outputs[5706]) & ~(layer2_outputs[182]);
    assign outputs[7214] = layer2_outputs[10114];
    assign outputs[7215] = ~(layer2_outputs[4478]);
    assign outputs[7216] = ~(layer2_outputs[1923]);
    assign outputs[7217] = ~(layer2_outputs[2777]);
    assign outputs[7218] = ~(layer2_outputs[10294]);
    assign outputs[7219] = ~(layer2_outputs[5619]) | (layer2_outputs[12685]);
    assign outputs[7220] = ~(layer2_outputs[9038]);
    assign outputs[7221] = (layer2_outputs[11685]) ^ (layer2_outputs[4204]);
    assign outputs[7222] = layer2_outputs[6675];
    assign outputs[7223] = ~((layer2_outputs[2185]) ^ (layer2_outputs[8934]));
    assign outputs[7224] = ~(layer2_outputs[4781]);
    assign outputs[7225] = ~(layer2_outputs[8389]);
    assign outputs[7226] = (layer2_outputs[1360]) ^ (layer2_outputs[6838]);
    assign outputs[7227] = layer2_outputs[8724];
    assign outputs[7228] = ~((layer2_outputs[9512]) & (layer2_outputs[1140]));
    assign outputs[7229] = (layer2_outputs[1727]) ^ (layer2_outputs[9179]);
    assign outputs[7230] = (layer2_outputs[2994]) ^ (layer2_outputs[4676]);
    assign outputs[7231] = layer2_outputs[12072];
    assign outputs[7232] = (layer2_outputs[5714]) ^ (layer2_outputs[1443]);
    assign outputs[7233] = (layer2_outputs[2542]) ^ (layer2_outputs[11201]);
    assign outputs[7234] = layer2_outputs[4817];
    assign outputs[7235] = (layer2_outputs[1629]) & (layer2_outputs[2378]);
    assign outputs[7236] = layer2_outputs[6412];
    assign outputs[7237] = (layer2_outputs[7869]) & ~(layer2_outputs[2101]);
    assign outputs[7238] = (layer2_outputs[4840]) ^ (layer2_outputs[2485]);
    assign outputs[7239] = ~((layer2_outputs[5321]) ^ (layer2_outputs[4210]));
    assign outputs[7240] = ~(layer2_outputs[4683]);
    assign outputs[7241] = layer2_outputs[4905];
    assign outputs[7242] = (layer2_outputs[856]) ^ (layer2_outputs[3684]);
    assign outputs[7243] = layer2_outputs[7007];
    assign outputs[7244] = ~(layer2_outputs[6417]);
    assign outputs[7245] = ~(layer2_outputs[9792]);
    assign outputs[7246] = layer2_outputs[9809];
    assign outputs[7247] = (layer2_outputs[1717]) | (layer2_outputs[10660]);
    assign outputs[7248] = (layer2_outputs[506]) ^ (layer2_outputs[3063]);
    assign outputs[7249] = ~(layer2_outputs[1784]);
    assign outputs[7250] = ~(layer2_outputs[2207]);
    assign outputs[7251] = (layer2_outputs[29]) ^ (layer2_outputs[12160]);
    assign outputs[7252] = (layer2_outputs[1761]) ^ (layer2_outputs[8961]);
    assign outputs[7253] = ~(layer2_outputs[2978]);
    assign outputs[7254] = (layer2_outputs[9886]) ^ (layer2_outputs[7593]);
    assign outputs[7255] = layer2_outputs[8216];
    assign outputs[7256] = layer2_outputs[9538];
    assign outputs[7257] = ~(layer2_outputs[4531]);
    assign outputs[7258] = ~(layer2_outputs[7275]);
    assign outputs[7259] = (layer2_outputs[8732]) & (layer2_outputs[10386]);
    assign outputs[7260] = layer2_outputs[6990];
    assign outputs[7261] = (layer2_outputs[6106]) & (layer2_outputs[4965]);
    assign outputs[7262] = layer2_outputs[3973];
    assign outputs[7263] = layer2_outputs[7937];
    assign outputs[7264] = (layer2_outputs[1667]) ^ (layer2_outputs[4305]);
    assign outputs[7265] = layer2_outputs[12228];
    assign outputs[7266] = ~((layer2_outputs[5561]) & (layer2_outputs[5613]));
    assign outputs[7267] = ~(layer2_outputs[7542]);
    assign outputs[7268] = (layer2_outputs[6116]) & ~(layer2_outputs[6620]);
    assign outputs[7269] = (layer2_outputs[11984]) ^ (layer2_outputs[7567]);
    assign outputs[7270] = layer2_outputs[11227];
    assign outputs[7271] = (layer2_outputs[2263]) | (layer2_outputs[3346]);
    assign outputs[7272] = ~(layer2_outputs[6916]);
    assign outputs[7273] = (layer2_outputs[10268]) ^ (layer2_outputs[8284]);
    assign outputs[7274] = ~(layer2_outputs[10228]);
    assign outputs[7275] = (layer2_outputs[5742]) ^ (layer2_outputs[7999]);
    assign outputs[7276] = ~(layer2_outputs[12331]);
    assign outputs[7277] = layer2_outputs[630];
    assign outputs[7278] = ~(layer2_outputs[485]) | (layer2_outputs[850]);
    assign outputs[7279] = layer2_outputs[3652];
    assign outputs[7280] = ~((layer2_outputs[4311]) ^ (layer2_outputs[749]));
    assign outputs[7281] = ~((layer2_outputs[5707]) ^ (layer2_outputs[11283]));
    assign outputs[7282] = ~((layer2_outputs[9276]) | (layer2_outputs[5329]));
    assign outputs[7283] = ~((layer2_outputs[2132]) | (layer2_outputs[678]));
    assign outputs[7284] = ~(layer2_outputs[11640]);
    assign outputs[7285] = ~(layer2_outputs[2647]);
    assign outputs[7286] = ~(layer2_outputs[1097]);
    assign outputs[7287] = layer2_outputs[9561];
    assign outputs[7288] = (layer2_outputs[2733]) ^ (layer2_outputs[8263]);
    assign outputs[7289] = ~(layer2_outputs[11743]);
    assign outputs[7290] = ~(layer2_outputs[1023]);
    assign outputs[7291] = ~((layer2_outputs[12191]) ^ (layer2_outputs[8331]));
    assign outputs[7292] = (layer2_outputs[11982]) ^ (layer2_outputs[9407]);
    assign outputs[7293] = layer2_outputs[7222];
    assign outputs[7294] = ~((layer2_outputs[792]) ^ (layer2_outputs[12516]));
    assign outputs[7295] = layer2_outputs[12732];
    assign outputs[7296] = layer2_outputs[12358];
    assign outputs[7297] = ~((layer2_outputs[4693]) ^ (layer2_outputs[8961]));
    assign outputs[7298] = (layer2_outputs[539]) ^ (layer2_outputs[6251]);
    assign outputs[7299] = (layer2_outputs[3296]) ^ (layer2_outputs[8125]);
    assign outputs[7300] = ~(layer2_outputs[7082]);
    assign outputs[7301] = (layer2_outputs[4647]) & ~(layer2_outputs[4820]);
    assign outputs[7302] = layer2_outputs[1240];
    assign outputs[7303] = ~((layer2_outputs[9189]) ^ (layer2_outputs[299]));
    assign outputs[7304] = (layer2_outputs[5781]) ^ (layer2_outputs[5115]);
    assign outputs[7305] = ~(layer2_outputs[8533]);
    assign outputs[7306] = ~((layer2_outputs[4018]) & (layer2_outputs[12627]));
    assign outputs[7307] = layer2_outputs[7392];
    assign outputs[7308] = ~((layer2_outputs[10144]) ^ (layer2_outputs[11484]));
    assign outputs[7309] = layer2_outputs[3863];
    assign outputs[7310] = (layer2_outputs[9182]) ^ (layer2_outputs[1576]);
    assign outputs[7311] = ~((layer2_outputs[8637]) ^ (layer2_outputs[12496]));
    assign outputs[7312] = (layer2_outputs[10526]) ^ (layer2_outputs[3621]);
    assign outputs[7313] = (layer2_outputs[5314]) ^ (layer2_outputs[5185]);
    assign outputs[7314] = (layer2_outputs[6006]) | (layer2_outputs[530]);
    assign outputs[7315] = ~((layer2_outputs[6317]) & (layer2_outputs[2033]));
    assign outputs[7316] = (layer2_outputs[11920]) | (layer2_outputs[9713]);
    assign outputs[7317] = layer2_outputs[9077];
    assign outputs[7318] = ~(layer2_outputs[8336]);
    assign outputs[7319] = layer2_outputs[187];
    assign outputs[7320] = (layer2_outputs[12435]) ^ (layer2_outputs[12385]);
    assign outputs[7321] = (layer2_outputs[2680]) & ~(layer2_outputs[4525]);
    assign outputs[7322] = (layer2_outputs[2259]) ^ (layer2_outputs[5202]);
    assign outputs[7323] = (layer2_outputs[10247]) & ~(layer2_outputs[11480]);
    assign outputs[7324] = (layer2_outputs[3868]) ^ (layer2_outputs[3032]);
    assign outputs[7325] = ~(layer2_outputs[5055]);
    assign outputs[7326] = layer2_outputs[11866];
    assign outputs[7327] = layer2_outputs[4131];
    assign outputs[7328] = layer2_outputs[8040];
    assign outputs[7329] = layer2_outputs[7067];
    assign outputs[7330] = (layer2_outputs[2437]) ^ (layer2_outputs[2648]);
    assign outputs[7331] = (layer2_outputs[614]) & ~(layer2_outputs[5856]);
    assign outputs[7332] = ~(layer2_outputs[4839]);
    assign outputs[7333] = layer2_outputs[9737];
    assign outputs[7334] = ~((layer2_outputs[12148]) ^ (layer2_outputs[3073]));
    assign outputs[7335] = (layer2_outputs[4015]) ^ (layer2_outputs[11488]);
    assign outputs[7336] = layer2_outputs[12403];
    assign outputs[7337] = ~((layer2_outputs[1409]) & (layer2_outputs[4496]));
    assign outputs[7338] = layer2_outputs[5313];
    assign outputs[7339] = layer2_outputs[7016];
    assign outputs[7340] = (layer2_outputs[3120]) ^ (layer2_outputs[7881]);
    assign outputs[7341] = ~(layer2_outputs[4363]);
    assign outputs[7342] = ~(layer2_outputs[5971]);
    assign outputs[7343] = ~((layer2_outputs[5663]) ^ (layer2_outputs[566]));
    assign outputs[7344] = layer2_outputs[7471];
    assign outputs[7345] = ~(layer2_outputs[11870]);
    assign outputs[7346] = layer2_outputs[5099];
    assign outputs[7347] = (layer2_outputs[9896]) ^ (layer2_outputs[4972]);
    assign outputs[7348] = ~(layer2_outputs[11081]);
    assign outputs[7349] = ~(layer2_outputs[10173]);
    assign outputs[7350] = ~(layer2_outputs[12710]);
    assign outputs[7351] = ~(layer2_outputs[7631]);
    assign outputs[7352] = ~(layer2_outputs[6367]);
    assign outputs[7353] = ~((layer2_outputs[5144]) ^ (layer2_outputs[5047]));
    assign outputs[7354] = ~(layer2_outputs[4555]);
    assign outputs[7355] = ~((layer2_outputs[1601]) ^ (layer2_outputs[6442]));
    assign outputs[7356] = layer2_outputs[5510];
    assign outputs[7357] = ~((layer2_outputs[12533]) ^ (layer2_outputs[5142]));
    assign outputs[7358] = ~(layer2_outputs[11292]);
    assign outputs[7359] = layer2_outputs[2993];
    assign outputs[7360] = ~(layer2_outputs[3442]);
    assign outputs[7361] = layer2_outputs[11478];
    assign outputs[7362] = ~((layer2_outputs[10455]) ^ (layer2_outputs[3358]));
    assign outputs[7363] = ~((layer2_outputs[11146]) & (layer2_outputs[6484]));
    assign outputs[7364] = layer2_outputs[10344];
    assign outputs[7365] = layer2_outputs[12260];
    assign outputs[7366] = layer2_outputs[4990];
    assign outputs[7367] = (layer2_outputs[818]) ^ (layer2_outputs[977]);
    assign outputs[7368] = ~(layer2_outputs[6534]);
    assign outputs[7369] = (layer2_outputs[9797]) ^ (layer2_outputs[12107]);
    assign outputs[7370] = (layer2_outputs[3106]) & ~(layer2_outputs[3752]);
    assign outputs[7371] = layer2_outputs[7385];
    assign outputs[7372] = (layer2_outputs[4237]) & ~(layer2_outputs[639]);
    assign outputs[7373] = ~(layer2_outputs[12539]);
    assign outputs[7374] = layer2_outputs[10288];
    assign outputs[7375] = layer2_outputs[6499];
    assign outputs[7376] = ~((layer2_outputs[11827]) | (layer2_outputs[3332]));
    assign outputs[7377] = (layer2_outputs[10995]) ^ (layer2_outputs[3067]);
    assign outputs[7378] = layer2_outputs[4411];
    assign outputs[7379] = layer2_outputs[3880];
    assign outputs[7380] = ~((layer2_outputs[2954]) ^ (layer2_outputs[5960]));
    assign outputs[7381] = ~((layer2_outputs[3482]) ^ (layer2_outputs[7143]));
    assign outputs[7382] = layer2_outputs[4654];
    assign outputs[7383] = (layer2_outputs[9945]) ^ (layer2_outputs[12639]);
    assign outputs[7384] = ~(layer2_outputs[11616]);
    assign outputs[7385] = ~(layer2_outputs[9427]);
    assign outputs[7386] = ~((layer2_outputs[7511]) ^ (layer2_outputs[864]));
    assign outputs[7387] = (layer2_outputs[2507]) ^ (layer2_outputs[3534]);
    assign outputs[7388] = layer2_outputs[7968];
    assign outputs[7389] = ~(layer2_outputs[11785]);
    assign outputs[7390] = ~(layer2_outputs[12255]);
    assign outputs[7391] = (layer2_outputs[1821]) & ~(layer2_outputs[3664]);
    assign outputs[7392] = ~(layer2_outputs[10890]) | (layer2_outputs[4668]);
    assign outputs[7393] = (layer2_outputs[9957]) ^ (layer2_outputs[7503]);
    assign outputs[7394] = ~(layer2_outputs[9748]);
    assign outputs[7395] = (layer2_outputs[6909]) ^ (layer2_outputs[711]);
    assign outputs[7396] = layer2_outputs[10198];
    assign outputs[7397] = ~(layer2_outputs[5195]) | (layer2_outputs[1657]);
    assign outputs[7398] = (layer2_outputs[2743]) & (layer2_outputs[11690]);
    assign outputs[7399] = ~((layer2_outputs[7091]) ^ (layer2_outputs[9924]));
    assign outputs[7400] = (layer2_outputs[10815]) ^ (layer2_outputs[11515]);
    assign outputs[7401] = ~((layer2_outputs[7321]) ^ (layer2_outputs[4422]));
    assign outputs[7402] = layer2_outputs[1485];
    assign outputs[7403] = layer2_outputs[10980];
    assign outputs[7404] = ~(layer2_outputs[6771]);
    assign outputs[7405] = layer2_outputs[5382];
    assign outputs[7406] = layer2_outputs[9988];
    assign outputs[7407] = layer2_outputs[6372];
    assign outputs[7408] = ~(layer2_outputs[3096]);
    assign outputs[7409] = ~(layer2_outputs[10773]);
    assign outputs[7410] = ~(layer2_outputs[6808]);
    assign outputs[7411] = ~((layer2_outputs[6850]) ^ (layer2_outputs[11834]));
    assign outputs[7412] = (layer2_outputs[4785]) ^ (layer2_outputs[9421]);
    assign outputs[7413] = ~(layer2_outputs[8962]);
    assign outputs[7414] = ~(layer2_outputs[1555]) | (layer2_outputs[7697]);
    assign outputs[7415] = ~((layer2_outputs[9534]) & (layer2_outputs[5946]));
    assign outputs[7416] = ~(layer2_outputs[10795]);
    assign outputs[7417] = ~(layer2_outputs[4969]) | (layer2_outputs[8301]);
    assign outputs[7418] = ~(layer2_outputs[8422]);
    assign outputs[7419] = ~(layer2_outputs[2764]);
    assign outputs[7420] = (layer2_outputs[7075]) & ~(layer2_outputs[699]);
    assign outputs[7421] = (layer2_outputs[9025]) ^ (layer2_outputs[7876]);
    assign outputs[7422] = ~(layer2_outputs[2266]);
    assign outputs[7423] = layer2_outputs[10887];
    assign outputs[7424] = (layer2_outputs[11833]) ^ (layer2_outputs[3477]);
    assign outputs[7425] = layer2_outputs[62];
    assign outputs[7426] = ~(layer2_outputs[5244]);
    assign outputs[7427] = layer2_outputs[5250];
    assign outputs[7428] = ~(layer2_outputs[2209]);
    assign outputs[7429] = layer2_outputs[245];
    assign outputs[7430] = (layer2_outputs[3305]) | (layer2_outputs[6644]);
    assign outputs[7431] = (layer2_outputs[2392]) ^ (layer2_outputs[8742]);
    assign outputs[7432] = ~(layer2_outputs[11905]);
    assign outputs[7433] = layer2_outputs[11622];
    assign outputs[7434] = (layer2_outputs[4739]) & ~(layer2_outputs[1715]);
    assign outputs[7435] = ~(layer2_outputs[1929]);
    assign outputs[7436] = ~((layer2_outputs[9226]) & (layer2_outputs[11052]));
    assign outputs[7437] = layer2_outputs[6170];
    assign outputs[7438] = layer2_outputs[11390];
    assign outputs[7439] = layer2_outputs[10046];
    assign outputs[7440] = (layer2_outputs[8189]) ^ (layer2_outputs[12219]);
    assign outputs[7441] = (layer2_outputs[3313]) | (layer2_outputs[912]);
    assign outputs[7442] = (layer2_outputs[3763]) ^ (layer2_outputs[3317]);
    assign outputs[7443] = (layer2_outputs[2244]) ^ (layer2_outputs[5794]);
    assign outputs[7444] = (layer2_outputs[7340]) & (layer2_outputs[7724]);
    assign outputs[7445] = (layer2_outputs[10041]) | (layer2_outputs[4797]);
    assign outputs[7446] = ~(layer2_outputs[6461]);
    assign outputs[7447] = ~(layer2_outputs[8657]);
    assign outputs[7448] = ~(layer2_outputs[4292]) | (layer2_outputs[10569]);
    assign outputs[7449] = ~(layer2_outputs[10897]);
    assign outputs[7450] = ~((layer2_outputs[9359]) ^ (layer2_outputs[2416]));
    assign outputs[7451] = layer2_outputs[7318];
    assign outputs[7452] = ~(layer2_outputs[5230]);
    assign outputs[7453] = ~((layer2_outputs[8576]) ^ (layer2_outputs[5357]));
    assign outputs[7454] = ~(layer2_outputs[8962]);
    assign outputs[7455] = ~(layer2_outputs[9993]);
    assign outputs[7456] = (layer2_outputs[6711]) ^ (layer2_outputs[9653]);
    assign outputs[7457] = ~(layer2_outputs[5231]);
    assign outputs[7458] = ~(layer2_outputs[3721]);
    assign outputs[7459] = ~((layer2_outputs[5214]) & (layer2_outputs[10144]));
    assign outputs[7460] = ~(layer2_outputs[3927]);
    assign outputs[7461] = layer2_outputs[4360];
    assign outputs[7462] = ~((layer2_outputs[8524]) ^ (layer2_outputs[798]));
    assign outputs[7463] = (layer2_outputs[2583]) ^ (layer2_outputs[2711]);
    assign outputs[7464] = ~(layer2_outputs[12432]);
    assign outputs[7465] = ~(layer2_outputs[8286]);
    assign outputs[7466] = (layer2_outputs[4591]) & ~(layer2_outputs[3979]);
    assign outputs[7467] = (layer2_outputs[6749]) ^ (layer2_outputs[3641]);
    assign outputs[7468] = (layer2_outputs[514]) ^ (layer2_outputs[424]);
    assign outputs[7469] = layer2_outputs[5692];
    assign outputs[7470] = (layer2_outputs[8036]) ^ (layer2_outputs[5824]);
    assign outputs[7471] = ~((layer2_outputs[11995]) | (layer2_outputs[2556]));
    assign outputs[7472] = layer2_outputs[37];
    assign outputs[7473] = ~(layer2_outputs[10762]) | (layer2_outputs[3186]);
    assign outputs[7474] = ~((layer2_outputs[12344]) ^ (layer2_outputs[2621]));
    assign outputs[7475] = layer2_outputs[6637];
    assign outputs[7476] = (layer2_outputs[5245]) ^ (layer2_outputs[842]);
    assign outputs[7477] = (layer2_outputs[2880]) & (layer2_outputs[4319]);
    assign outputs[7478] = ~((layer2_outputs[8171]) & (layer2_outputs[10823]));
    assign outputs[7479] = layer2_outputs[3248];
    assign outputs[7480] = layer2_outputs[11032];
    assign outputs[7481] = ~(layer2_outputs[4794]);
    assign outputs[7482] = layer2_outputs[8444];
    assign outputs[7483] = (layer2_outputs[5631]) & ~(layer2_outputs[11503]);
    assign outputs[7484] = ~((layer2_outputs[8585]) ^ (layer2_outputs[12753]));
    assign outputs[7485] = ~(layer2_outputs[5126]);
    assign outputs[7486] = ~((layer2_outputs[5273]) ^ (layer2_outputs[12151]));
    assign outputs[7487] = ~(layer2_outputs[913]) | (layer2_outputs[11715]);
    assign outputs[7488] = ~(layer2_outputs[9616]);
    assign outputs[7489] = (layer2_outputs[11892]) ^ (layer2_outputs[8983]);
    assign outputs[7490] = ~(layer2_outputs[6695]);
    assign outputs[7491] = layer2_outputs[453];
    assign outputs[7492] = layer2_outputs[4878];
    assign outputs[7493] = layer2_outputs[12606];
    assign outputs[7494] = (layer2_outputs[11347]) ^ (layer2_outputs[7964]);
    assign outputs[7495] = layer2_outputs[9738];
    assign outputs[7496] = ~((layer2_outputs[5490]) | (layer2_outputs[4968]));
    assign outputs[7497] = layer2_outputs[4444];
    assign outputs[7498] = layer2_outputs[8115];
    assign outputs[7499] = (layer2_outputs[7399]) ^ (layer2_outputs[3398]);
    assign outputs[7500] = (layer2_outputs[4100]) & ~(layer2_outputs[9343]);
    assign outputs[7501] = ~(layer2_outputs[6899]);
    assign outputs[7502] = ~((layer2_outputs[5025]) ^ (layer2_outputs[3050]));
    assign outputs[7503] = ~((layer2_outputs[5110]) ^ (layer2_outputs[3221]));
    assign outputs[7504] = ~((layer2_outputs[9650]) ^ (layer2_outputs[3401]));
    assign outputs[7505] = layer2_outputs[4035];
    assign outputs[7506] = ~(layer2_outputs[10179]) | (layer2_outputs[6716]);
    assign outputs[7507] = layer2_outputs[11764];
    assign outputs[7508] = ~(layer2_outputs[253]);
    assign outputs[7509] = layer2_outputs[3860];
    assign outputs[7510] = layer2_outputs[6819];
    assign outputs[7511] = ~((layer2_outputs[10813]) ^ (layer2_outputs[8448]));
    assign outputs[7512] = ~(layer2_outputs[12407]);
    assign outputs[7513] = ~((layer2_outputs[3997]) ^ (layer2_outputs[6081]));
    assign outputs[7514] = ~((layer2_outputs[1311]) ^ (layer2_outputs[4667]));
    assign outputs[7515] = layer2_outputs[11987];
    assign outputs[7516] = layer2_outputs[710];
    assign outputs[7517] = (layer2_outputs[4414]) ^ (layer2_outputs[8201]);
    assign outputs[7518] = (layer2_outputs[1508]) ^ (layer2_outputs[3981]);
    assign outputs[7519] = ~((layer2_outputs[2814]) & (layer2_outputs[6301]));
    assign outputs[7520] = ~((layer2_outputs[11630]) ^ (layer2_outputs[690]));
    assign outputs[7521] = ~(layer2_outputs[5457]);
    assign outputs[7522] = ~(layer2_outputs[4178]);
    assign outputs[7523] = (layer2_outputs[11980]) ^ (layer2_outputs[231]);
    assign outputs[7524] = layer2_outputs[12036];
    assign outputs[7525] = (layer2_outputs[607]) & ~(layer2_outputs[12051]);
    assign outputs[7526] = layer2_outputs[532];
    assign outputs[7527] = (layer2_outputs[8352]) ^ (layer2_outputs[1049]);
    assign outputs[7528] = layer2_outputs[12663];
    assign outputs[7529] = (layer2_outputs[12794]) ^ (layer2_outputs[7901]);
    assign outputs[7530] = ~(layer2_outputs[6131]);
    assign outputs[7531] = ~(layer2_outputs[5840]) | (layer2_outputs[11484]);
    assign outputs[7532] = layer2_outputs[8321];
    assign outputs[7533] = ~((layer2_outputs[7916]) ^ (layer2_outputs[2495]));
    assign outputs[7534] = ~(layer2_outputs[5524]);
    assign outputs[7535] = ~((layer2_outputs[741]) ^ (layer2_outputs[9443]));
    assign outputs[7536] = layer2_outputs[649];
    assign outputs[7537] = ~((layer2_outputs[10545]) ^ (layer2_outputs[5412]));
    assign outputs[7538] = (layer2_outputs[6227]) & ~(layer2_outputs[3639]);
    assign outputs[7539] = ~(layer2_outputs[3878]);
    assign outputs[7540] = ~(layer2_outputs[8276]);
    assign outputs[7541] = ~((layer2_outputs[1510]) ^ (layer2_outputs[2361]));
    assign outputs[7542] = layer2_outputs[444];
    assign outputs[7543] = ~(layer2_outputs[3523]);
    assign outputs[7544] = ~((layer2_outputs[11131]) ^ (layer2_outputs[7799]));
    assign outputs[7545] = ~(layer2_outputs[11347]) | (layer2_outputs[54]);
    assign outputs[7546] = (layer2_outputs[10806]) ^ (layer2_outputs[8993]);
    assign outputs[7547] = ~(layer2_outputs[10107]);
    assign outputs[7548] = ~((layer2_outputs[1018]) ^ (layer2_outputs[12224]));
    assign outputs[7549] = ~(layer2_outputs[4844]);
    assign outputs[7550] = layer2_outputs[4621];
    assign outputs[7551] = layer2_outputs[6969];
    assign outputs[7552] = layer2_outputs[4429];
    assign outputs[7553] = layer2_outputs[2344];
    assign outputs[7554] = (layer2_outputs[3775]) ^ (layer2_outputs[545]);
    assign outputs[7555] = ~(layer2_outputs[8116]);
    assign outputs[7556] = layer2_outputs[6759];
    assign outputs[7557] = (layer2_outputs[1167]) ^ (layer2_outputs[4125]);
    assign outputs[7558] = ~(layer2_outputs[10658]) | (layer2_outputs[1427]);
    assign outputs[7559] = ~(layer2_outputs[8534]);
    assign outputs[7560] = ~(layer2_outputs[5265]);
    assign outputs[7561] = ~((layer2_outputs[11153]) ^ (layer2_outputs[7335]));
    assign outputs[7562] = (layer2_outputs[418]) ^ (layer2_outputs[1443]);
    assign outputs[7563] = (layer2_outputs[1905]) ^ (layer2_outputs[9465]);
    assign outputs[7564] = ~(layer2_outputs[7536]);
    assign outputs[7565] = ~(layer2_outputs[3797]);
    assign outputs[7566] = (layer2_outputs[9242]) & ~(layer2_outputs[11519]);
    assign outputs[7567] = layer2_outputs[2737];
    assign outputs[7568] = ~(layer2_outputs[9618]);
    assign outputs[7569] = layer2_outputs[12681];
    assign outputs[7570] = ~((layer2_outputs[5396]) ^ (layer2_outputs[2098]));
    assign outputs[7571] = ~(layer2_outputs[8400]);
    assign outputs[7572] = (layer2_outputs[7308]) ^ (layer2_outputs[3022]);
    assign outputs[7573] = ~(layer2_outputs[9387]);
    assign outputs[7574] = ~(layer2_outputs[1024]) | (layer2_outputs[10219]);
    assign outputs[7575] = layer2_outputs[9968];
    assign outputs[7576] = ~(layer2_outputs[8055]);
    assign outputs[7577] = (layer2_outputs[3501]) ^ (layer2_outputs[7228]);
    assign outputs[7578] = ~(layer2_outputs[10002]) | (layer2_outputs[4668]);
    assign outputs[7579] = (layer2_outputs[7333]) ^ (layer2_outputs[12722]);
    assign outputs[7580] = layer2_outputs[11336];
    assign outputs[7581] = ~(layer2_outputs[11187]);
    assign outputs[7582] = layer2_outputs[11443];
    assign outputs[7583] = ~(layer2_outputs[8812]);
    assign outputs[7584] = layer2_outputs[8851];
    assign outputs[7585] = ~(layer2_outputs[12785]);
    assign outputs[7586] = (layer2_outputs[8403]) ^ (layer2_outputs[948]);
    assign outputs[7587] = layer2_outputs[4288];
    assign outputs[7588] = ~((layer2_outputs[10735]) & (layer2_outputs[5878]));
    assign outputs[7589] = ~((layer2_outputs[11489]) ^ (layer2_outputs[3740]));
    assign outputs[7590] = ~(layer2_outputs[9581]);
    assign outputs[7591] = layer2_outputs[11082];
    assign outputs[7592] = ~((layer2_outputs[6509]) & (layer2_outputs[7887]));
    assign outputs[7593] = ~((layer2_outputs[1372]) & (layer2_outputs[9911]));
    assign outputs[7594] = ~(layer2_outputs[1493]) | (layer2_outputs[6587]);
    assign outputs[7595] = ~((layer2_outputs[10950]) & (layer2_outputs[2012]));
    assign outputs[7596] = ~(layer2_outputs[6977]) | (layer2_outputs[12132]);
    assign outputs[7597] = layer2_outputs[7435];
    assign outputs[7598] = layer2_outputs[12092];
    assign outputs[7599] = ~(layer2_outputs[4901]);
    assign outputs[7600] = ~(layer2_outputs[8517]);
    assign outputs[7601] = ~(layer2_outputs[8037]);
    assign outputs[7602] = (layer2_outputs[9383]) ^ (layer2_outputs[4699]);
    assign outputs[7603] = ~(layer2_outputs[6951]);
    assign outputs[7604] = (layer2_outputs[7865]) & (layer2_outputs[9591]);
    assign outputs[7605] = ~(layer2_outputs[10956]);
    assign outputs[7606] = layer2_outputs[3959];
    assign outputs[7607] = layer2_outputs[12005];
    assign outputs[7608] = layer2_outputs[12789];
    assign outputs[7609] = layer2_outputs[11904];
    assign outputs[7610] = (layer2_outputs[6967]) ^ (layer2_outputs[2205]);
    assign outputs[7611] = (layer2_outputs[8792]) & ~(layer2_outputs[5697]);
    assign outputs[7612] = ~((layer2_outputs[3853]) | (layer2_outputs[6832]));
    assign outputs[7613] = (layer2_outputs[8084]) ^ (layer2_outputs[1634]);
    assign outputs[7614] = ~(layer2_outputs[6927]);
    assign outputs[7615] = ~(layer2_outputs[11170]);
    assign outputs[7616] = ~(layer2_outputs[7426]);
    assign outputs[7617] = layer2_outputs[9034];
    assign outputs[7618] = (layer2_outputs[7083]) ^ (layer2_outputs[8542]);
    assign outputs[7619] = ~((layer2_outputs[1813]) ^ (layer2_outputs[6907]));
    assign outputs[7620] = ~(layer2_outputs[11746]);
    assign outputs[7621] = (layer2_outputs[5853]) ^ (layer2_outputs[10043]);
    assign outputs[7622] = ~((layer2_outputs[7537]) & (layer2_outputs[10503]));
    assign outputs[7623] = ~((layer2_outputs[5568]) ^ (layer2_outputs[4084]));
    assign outputs[7624] = layer2_outputs[10798];
    assign outputs[7625] = ~(layer2_outputs[8670]);
    assign outputs[7626] = layer2_outputs[4997];
    assign outputs[7627] = (layer2_outputs[9605]) ^ (layer2_outputs[9634]);
    assign outputs[7628] = (layer2_outputs[6704]) ^ (layer2_outputs[4250]);
    assign outputs[7629] = layer2_outputs[1053];
    assign outputs[7630] = layer2_outputs[732];
    assign outputs[7631] = layer2_outputs[577];
    assign outputs[7632] = (layer2_outputs[1501]) ^ (layer2_outputs[5093]);
    assign outputs[7633] = (layer2_outputs[11593]) & ~(layer2_outputs[3750]);
    assign outputs[7634] = (layer2_outputs[5018]) ^ (layer2_outputs[430]);
    assign outputs[7635] = ~(layer2_outputs[3924]);
    assign outputs[7636] = layer2_outputs[673];
    assign outputs[7637] = (layer2_outputs[10400]) ^ (layer2_outputs[9166]);
    assign outputs[7638] = ~(layer2_outputs[2389]);
    assign outputs[7639] = (layer2_outputs[5458]) ^ (layer2_outputs[10026]);
    assign outputs[7640] = (layer2_outputs[9992]) & ~(layer2_outputs[4771]);
    assign outputs[7641] = (layer2_outputs[6295]) ^ (layer2_outputs[1820]);
    assign outputs[7642] = (layer2_outputs[4401]) ^ (layer2_outputs[10474]);
    assign outputs[7643] = (layer2_outputs[11700]) ^ (layer2_outputs[11149]);
    assign outputs[7644] = ~(layer2_outputs[4670]);
    assign outputs[7645] = (layer2_outputs[7721]) & ~(layer2_outputs[1732]);
    assign outputs[7646] = layer2_outputs[3430];
    assign outputs[7647] = layer2_outputs[9206];
    assign outputs[7648] = (layer2_outputs[10072]) ^ (layer2_outputs[9012]);
    assign outputs[7649] = layer2_outputs[2510];
    assign outputs[7650] = (layer2_outputs[1863]) ^ (layer2_outputs[11780]);
    assign outputs[7651] = ~((layer2_outputs[10845]) | (layer2_outputs[1188]));
    assign outputs[7652] = ~((layer2_outputs[9327]) ^ (layer2_outputs[4491]));
    assign outputs[7653] = layer2_outputs[3354];
    assign outputs[7654] = (layer2_outputs[5710]) & ~(layer2_outputs[1729]);
    assign outputs[7655] = ~(layer2_outputs[8353]);
    assign outputs[7656] = (layer2_outputs[1626]) & ~(layer2_outputs[4544]);
    assign outputs[7657] = layer2_outputs[11526];
    assign outputs[7658] = ~((layer2_outputs[6909]) ^ (layer2_outputs[12202]));
    assign outputs[7659] = layer2_outputs[7849];
    assign outputs[7660] = ~((layer2_outputs[3088]) ^ (layer2_outputs[9214]));
    assign outputs[7661] = (layer2_outputs[5281]) ^ (layer2_outputs[10121]);
    assign outputs[7662] = ~((layer2_outputs[1256]) ^ (layer2_outputs[5734]));
    assign outputs[7663] = ~(layer2_outputs[2485]);
    assign outputs[7664] = ~(layer2_outputs[8349]);
    assign outputs[7665] = layer2_outputs[8763];
    assign outputs[7666] = layer2_outputs[8813];
    assign outputs[7667] = layer2_outputs[11703];
    assign outputs[7668] = layer2_outputs[12501];
    assign outputs[7669] = layer2_outputs[1659];
    assign outputs[7670] = ~(layer2_outputs[11261]) | (layer2_outputs[6868]);
    assign outputs[7671] = ~((layer2_outputs[1560]) ^ (layer2_outputs[2232]));
    assign outputs[7672] = (layer2_outputs[7943]) & ~(layer2_outputs[6306]);
    assign outputs[7673] = ~(layer2_outputs[10051]) | (layer2_outputs[11903]);
    assign outputs[7674] = layer2_outputs[12216];
    assign outputs[7675] = ~((layer2_outputs[4445]) ^ (layer2_outputs[5059]));
    assign outputs[7676] = ~(layer2_outputs[11384]);
    assign outputs[7677] = layer2_outputs[10889];
    assign outputs[7678] = layer2_outputs[9898];
    assign outputs[7679] = ~(layer2_outputs[7703]);
    assign outputs[7680] = layer2_outputs[9212];
    assign outputs[7681] = layer2_outputs[10775];
    assign outputs[7682] = ~(layer2_outputs[1933]);
    assign outputs[7683] = (layer2_outputs[2928]) ^ (layer2_outputs[6847]);
    assign outputs[7684] = layer2_outputs[11767];
    assign outputs[7685] = layer2_outputs[5029];
    assign outputs[7686] = layer2_outputs[6376];
    assign outputs[7687] = ~(layer2_outputs[6178]);
    assign outputs[7688] = layer2_outputs[5152];
    assign outputs[7689] = ~(layer2_outputs[10130]);
    assign outputs[7690] = ~(layer2_outputs[413]);
    assign outputs[7691] = ~(layer2_outputs[7908]);
    assign outputs[7692] = ~(layer2_outputs[2239]);
    assign outputs[7693] = ~(layer2_outputs[9286]) | (layer2_outputs[7248]);
    assign outputs[7694] = ~(layer2_outputs[7511]) | (layer2_outputs[551]);
    assign outputs[7695] = (layer2_outputs[7419]) ^ (layer2_outputs[5895]);
    assign outputs[7696] = ~((layer2_outputs[12385]) & (layer2_outputs[823]));
    assign outputs[7697] = layer2_outputs[6487];
    assign outputs[7698] = layer2_outputs[12509];
    assign outputs[7699] = (layer2_outputs[1939]) & (layer2_outputs[100]);
    assign outputs[7700] = ~(layer2_outputs[11962]);
    assign outputs[7701] = (layer2_outputs[1452]) ^ (layer2_outputs[3911]);
    assign outputs[7702] = (layer2_outputs[6872]) & ~(layer2_outputs[4563]);
    assign outputs[7703] = ~(layer2_outputs[4421]);
    assign outputs[7704] = layer2_outputs[4281];
    assign outputs[7705] = ~(layer2_outputs[5710]);
    assign outputs[7706] = (layer2_outputs[4039]) & ~(layer2_outputs[4082]);
    assign outputs[7707] = layer2_outputs[4405];
    assign outputs[7708] = ~(layer2_outputs[3156]);
    assign outputs[7709] = layer2_outputs[10610];
    assign outputs[7710] = layer2_outputs[10952];
    assign outputs[7711] = layer2_outputs[4791];
    assign outputs[7712] = layer2_outputs[12530];
    assign outputs[7713] = (layer2_outputs[1213]) & ~(layer2_outputs[5092]);
    assign outputs[7714] = (layer2_outputs[9934]) ^ (layer2_outputs[218]);
    assign outputs[7715] = ~(layer2_outputs[2331]);
    assign outputs[7716] = layer2_outputs[6334];
    assign outputs[7717] = layer2_outputs[1972];
    assign outputs[7718] = layer2_outputs[2354];
    assign outputs[7719] = ~(layer2_outputs[4766]);
    assign outputs[7720] = layer2_outputs[6846];
    assign outputs[7721] = ~((layer2_outputs[11750]) & (layer2_outputs[2668]));
    assign outputs[7722] = ~(layer2_outputs[5729]) | (layer2_outputs[12467]);
    assign outputs[7723] = ~((layer2_outputs[36]) ^ (layer2_outputs[6437]));
    assign outputs[7724] = ~(layer2_outputs[12519]);
    assign outputs[7725] = (layer2_outputs[11623]) & ~(layer2_outputs[11743]);
    assign outputs[7726] = ~((layer2_outputs[8890]) ^ (layer2_outputs[4298]));
    assign outputs[7727] = layer2_outputs[12219];
    assign outputs[7728] = (layer2_outputs[6391]) & (layer2_outputs[10619]);
    assign outputs[7729] = layer2_outputs[7365];
    assign outputs[7730] = ~(layer2_outputs[12455]);
    assign outputs[7731] = ~(layer2_outputs[8831]);
    assign outputs[7732] = ~((layer2_outputs[3257]) ^ (layer2_outputs[12152]));
    assign outputs[7733] = layer2_outputs[4169];
    assign outputs[7734] = ~(layer2_outputs[8558]);
    assign outputs[7735] = (layer2_outputs[8535]) & ~(layer2_outputs[8371]);
    assign outputs[7736] = ~(layer2_outputs[6549]);
    assign outputs[7737] = ~(layer2_outputs[11161]);
    assign outputs[7738] = ~(layer2_outputs[10248]);
    assign outputs[7739] = layer2_outputs[7271];
    assign outputs[7740] = ~(layer2_outputs[4112]);
    assign outputs[7741] = ~(layer2_outputs[3577]);
    assign outputs[7742] = ~((layer2_outputs[5615]) ^ (layer2_outputs[6168]));
    assign outputs[7743] = layer2_outputs[7784];
    assign outputs[7744] = (layer2_outputs[12710]) & (layer2_outputs[267]);
    assign outputs[7745] = ~(layer2_outputs[2858]) | (layer2_outputs[8980]);
    assign outputs[7746] = layer2_outputs[702];
    assign outputs[7747] = layer2_outputs[1029];
    assign outputs[7748] = layer2_outputs[4912];
    assign outputs[7749] = layer2_outputs[590];
    assign outputs[7750] = (layer2_outputs[11773]) & (layer2_outputs[4995]);
    assign outputs[7751] = ~(layer2_outputs[11537]);
    assign outputs[7752] = ~((layer2_outputs[3528]) ^ (layer2_outputs[4633]));
    assign outputs[7753] = ~(layer2_outputs[6848]);
    assign outputs[7754] = layer2_outputs[11688];
    assign outputs[7755] = (layer2_outputs[414]) ^ (layer2_outputs[4945]);
    assign outputs[7756] = ~(layer2_outputs[9805]);
    assign outputs[7757] = layer2_outputs[4821];
    assign outputs[7758] = ~(layer2_outputs[4480]);
    assign outputs[7759] = ~((layer2_outputs[9575]) | (layer2_outputs[3124]));
    assign outputs[7760] = layer2_outputs[6536];
    assign outputs[7761] = ~(layer2_outputs[11400]) | (layer2_outputs[1848]);
    assign outputs[7762] = ~(layer2_outputs[10853]);
    assign outputs[7763] = ~((layer2_outputs[9347]) ^ (layer2_outputs[11836]));
    assign outputs[7764] = layer2_outputs[8057];
    assign outputs[7765] = layer2_outputs[10370];
    assign outputs[7766] = layer2_outputs[10418];
    assign outputs[7767] = layer2_outputs[3647];
    assign outputs[7768] = layer2_outputs[8685];
    assign outputs[7769] = layer2_outputs[3921];
    assign outputs[7770] = layer2_outputs[6440];
    assign outputs[7771] = ~((layer2_outputs[219]) ^ (layer2_outputs[4514]));
    assign outputs[7772] = (layer2_outputs[1061]) & ~(layer2_outputs[9758]);
    assign outputs[7773] = ~(layer2_outputs[8318]);
    assign outputs[7774] = ~(layer2_outputs[6263]) | (layer2_outputs[3740]);
    assign outputs[7775] = (layer2_outputs[10380]) & ~(layer2_outputs[12610]);
    assign outputs[7776] = ~((layer2_outputs[2370]) & (layer2_outputs[6275]));
    assign outputs[7777] = (layer2_outputs[10824]) & ~(layer2_outputs[4982]);
    assign outputs[7778] = layer2_outputs[3767];
    assign outputs[7779] = ~(layer2_outputs[6587]);
    assign outputs[7780] = layer2_outputs[6780];
    assign outputs[7781] = (layer2_outputs[94]) ^ (layer2_outputs[483]);
    assign outputs[7782] = layer2_outputs[6613];
    assign outputs[7783] = ~(layer2_outputs[5437]);
    assign outputs[7784] = ~((layer2_outputs[7796]) ^ (layer2_outputs[4530]));
    assign outputs[7785] = ~(layer2_outputs[1002]);
    assign outputs[7786] = ~(layer2_outputs[4503]);
    assign outputs[7787] = ~(layer2_outputs[10431]);
    assign outputs[7788] = ~(layer2_outputs[11602]);
    assign outputs[7789] = ~(layer2_outputs[11556]);
    assign outputs[7790] = ~(layer2_outputs[10536]);
    assign outputs[7791] = layer2_outputs[330];
    assign outputs[7792] = ~(layer2_outputs[12294]);
    assign outputs[7793] = ~(layer2_outputs[8013]) | (layer2_outputs[2186]);
    assign outputs[7794] = ~(layer2_outputs[9825]);
    assign outputs[7795] = layer2_outputs[12404];
    assign outputs[7796] = layer2_outputs[6460];
    assign outputs[7797] = ~(layer2_outputs[11944]);
    assign outputs[7798] = layer2_outputs[12391];
    assign outputs[7799] = (layer2_outputs[11921]) ^ (layer2_outputs[9253]);
    assign outputs[7800] = (layer2_outputs[1069]) ^ (layer2_outputs[305]);
    assign outputs[7801] = layer2_outputs[9523];
    assign outputs[7802] = layer2_outputs[8365];
    assign outputs[7803] = (layer2_outputs[4769]) ^ (layer2_outputs[8838]);
    assign outputs[7804] = (layer2_outputs[3365]) ^ (layer2_outputs[5283]);
    assign outputs[7805] = (layer2_outputs[10190]) & ~(layer2_outputs[3887]);
    assign outputs[7806] = ~(layer2_outputs[12394]);
    assign outputs[7807] = ~(layer2_outputs[884]);
    assign outputs[7808] = layer2_outputs[12427];
    assign outputs[7809] = ~(layer2_outputs[4147]);
    assign outputs[7810] = (layer2_outputs[11027]) & ~(layer2_outputs[9736]);
    assign outputs[7811] = layer2_outputs[5967];
    assign outputs[7812] = ~((layer2_outputs[8682]) | (layer2_outputs[6167]));
    assign outputs[7813] = (layer2_outputs[3222]) & (layer2_outputs[8857]);
    assign outputs[7814] = layer2_outputs[1561];
    assign outputs[7815] = (layer2_outputs[2379]) ^ (layer2_outputs[1362]);
    assign outputs[7816] = ~((layer2_outputs[3051]) ^ (layer2_outputs[3277]));
    assign outputs[7817] = (layer2_outputs[9419]) & ~(layer2_outputs[752]);
    assign outputs[7818] = ~((layer2_outputs[2666]) & (layer2_outputs[1367]));
    assign outputs[7819] = (layer2_outputs[6931]) & ~(layer2_outputs[2115]);
    assign outputs[7820] = (layer2_outputs[1587]) & ~(layer2_outputs[12555]);
    assign outputs[7821] = ~((layer2_outputs[7510]) ^ (layer2_outputs[7561]));
    assign outputs[7822] = ~(layer2_outputs[7468]);
    assign outputs[7823] = layer2_outputs[7418];
    assign outputs[7824] = ~(layer2_outputs[12638]);
    assign outputs[7825] = ~(layer2_outputs[5726]);
    assign outputs[7826] = ~(layer2_outputs[437]) | (layer2_outputs[11741]);
    assign outputs[7827] = ~(layer2_outputs[5192]);
    assign outputs[7828] = layer2_outputs[3351];
    assign outputs[7829] = ~(layer2_outputs[6141]);
    assign outputs[7830] = (layer2_outputs[9763]) & ~(layer2_outputs[2226]);
    assign outputs[7831] = layer2_outputs[12120];
    assign outputs[7832] = ~(layer2_outputs[12111]);
    assign outputs[7833] = ~((layer2_outputs[4284]) & (layer2_outputs[7298]));
    assign outputs[7834] = ~((layer2_outputs[12755]) ^ (layer2_outputs[8559]));
    assign outputs[7835] = layer2_outputs[9293];
    assign outputs[7836] = ~((layer2_outputs[5340]) | (layer2_outputs[12289]));
    assign outputs[7837] = (layer2_outputs[11805]) & (layer2_outputs[2470]);
    assign outputs[7838] = layer2_outputs[19];
    assign outputs[7839] = (layer2_outputs[1195]) | (layer2_outputs[2825]);
    assign outputs[7840] = (layer2_outputs[11898]) & (layer2_outputs[7346]);
    assign outputs[7841] = (layer2_outputs[6670]) ^ (layer2_outputs[6063]);
    assign outputs[7842] = ~(layer2_outputs[1725]);
    assign outputs[7843] = (layer2_outputs[8456]) ^ (layer2_outputs[8061]);
    assign outputs[7844] = ~((layer2_outputs[12106]) ^ (layer2_outputs[9559]));
    assign outputs[7845] = ~(layer2_outputs[1588]);
    assign outputs[7846] = layer2_outputs[7299];
    assign outputs[7847] = ~((layer2_outputs[10761]) ^ (layer2_outputs[194]));
    assign outputs[7848] = ~(layer2_outputs[7924]);
    assign outputs[7849] = layer2_outputs[1561];
    assign outputs[7850] = ~(layer2_outputs[5687]);
    assign outputs[7851] = (layer2_outputs[2579]) ^ (layer2_outputs[858]);
    assign outputs[7852] = layer2_outputs[336];
    assign outputs[7853] = ~(layer2_outputs[5998]);
    assign outputs[7854] = ~((layer2_outputs[4949]) ^ (layer2_outputs[5995]));
    assign outputs[7855] = layer2_outputs[11613];
    assign outputs[7856] = (layer2_outputs[1424]) & ~(layer2_outputs[1152]);
    assign outputs[7857] = layer2_outputs[4719];
    assign outputs[7858] = ~((layer2_outputs[9184]) ^ (layer2_outputs[12674]));
    assign outputs[7859] = ~((layer2_outputs[8767]) & (layer2_outputs[6768]));
    assign outputs[7860] = layer2_outputs[11483];
    assign outputs[7861] = ~(layer2_outputs[738]) | (layer2_outputs[2354]);
    assign outputs[7862] = (layer2_outputs[5370]) & ~(layer2_outputs[9507]);
    assign outputs[7863] = layer2_outputs[4028];
    assign outputs[7864] = layer2_outputs[6788];
    assign outputs[7865] = layer2_outputs[11333];
    assign outputs[7866] = layer2_outputs[7129];
    assign outputs[7867] = (layer2_outputs[12530]) | (layer2_outputs[11577]);
    assign outputs[7868] = ~((layer2_outputs[3331]) ^ (layer2_outputs[3249]));
    assign outputs[7869] = layer2_outputs[591];
    assign outputs[7870] = layer2_outputs[9584];
    assign outputs[7871] = layer2_outputs[3037];
    assign outputs[7872] = ~(layer2_outputs[8335]);
    assign outputs[7873] = layer2_outputs[899];
    assign outputs[7874] = ~(layer2_outputs[7380]);
    assign outputs[7875] = (layer2_outputs[8519]) & (layer2_outputs[11972]);
    assign outputs[7876] = ~(layer2_outputs[7755]);
    assign outputs[7877] = ~(layer2_outputs[11850]);
    assign outputs[7878] = layer2_outputs[1834];
    assign outputs[7879] = (layer2_outputs[8422]) | (layer2_outputs[4346]);
    assign outputs[7880] = ~(layer2_outputs[6793]);
    assign outputs[7881] = layer2_outputs[6823];
    assign outputs[7882] = ~((layer2_outputs[11503]) ^ (layer2_outputs[11078]));
    assign outputs[7883] = ~(layer2_outputs[2422]);
    assign outputs[7884] = layer2_outputs[2533];
    assign outputs[7885] = (layer2_outputs[2824]) ^ (layer2_outputs[8043]);
    assign outputs[7886] = (layer2_outputs[9718]) & ~(layer2_outputs[7620]);
    assign outputs[7887] = layer2_outputs[193];
    assign outputs[7888] = layer2_outputs[11759];
    assign outputs[7889] = (layer2_outputs[9558]) & (layer2_outputs[11181]);
    assign outputs[7890] = ~(layer2_outputs[6564]);
    assign outputs[7891] = ~(layer2_outputs[4448]);
    assign outputs[7892] = ~((layer2_outputs[12676]) ^ (layer2_outputs[4915]));
    assign outputs[7893] = (layer2_outputs[11513]) & ~(layer2_outputs[8564]);
    assign outputs[7894] = (layer2_outputs[1528]) ^ (layer2_outputs[1216]);
    assign outputs[7895] = ~((layer2_outputs[10721]) ^ (layer2_outputs[5871]));
    assign outputs[7896] = ~(layer2_outputs[2279]);
    assign outputs[7897] = ~((layer2_outputs[10831]) | (layer2_outputs[9395]));
    assign outputs[7898] = ~((layer2_outputs[1028]) ^ (layer2_outputs[1300]));
    assign outputs[7899] = ~(layer2_outputs[2130]) | (layer2_outputs[2298]);
    assign outputs[7900] = ~(layer2_outputs[6664]);
    assign outputs[7901] = ~(layer2_outputs[9458]);
    assign outputs[7902] = ~(layer2_outputs[7386]);
    assign outputs[7903] = ~(layer2_outputs[1236]);
    assign outputs[7904] = layer2_outputs[700];
    assign outputs[7905] = ~(layer2_outputs[2617]);
    assign outputs[7906] = (layer2_outputs[8857]) & (layer2_outputs[7405]);
    assign outputs[7907] = ~(layer2_outputs[12612]);
    assign outputs[7908] = (layer2_outputs[12216]) ^ (layer2_outputs[11050]);
    assign outputs[7909] = ~((layer2_outputs[3054]) | (layer2_outputs[4525]));
    assign outputs[7910] = ~(layer2_outputs[7187]);
    assign outputs[7911] = ~((layer2_outputs[5780]) ^ (layer2_outputs[1488]));
    assign outputs[7912] = ~(layer2_outputs[9218]);
    assign outputs[7913] = ~(layer2_outputs[4559]);
    assign outputs[7914] = ~(layer2_outputs[11270]);
    assign outputs[7915] = ~(layer2_outputs[8499]);
    assign outputs[7916] = layer2_outputs[9244];
    assign outputs[7917] = layer2_outputs[6440];
    assign outputs[7918] = layer2_outputs[6014];
    assign outputs[7919] = ~(layer2_outputs[12539]);
    assign outputs[7920] = ~(layer2_outputs[3798]);
    assign outputs[7921] = ~(layer2_outputs[5992]);
    assign outputs[7922] = layer2_outputs[3174];
    assign outputs[7923] = ~(layer2_outputs[8171]) | (layer2_outputs[9045]);
    assign outputs[7924] = layer2_outputs[1217];
    assign outputs[7925] = ~(layer2_outputs[4520]);
    assign outputs[7926] = ~(layer2_outputs[5462]);
    assign outputs[7927] = ~(layer2_outputs[8897]);
    assign outputs[7928] = ~(layer2_outputs[4372]);
    assign outputs[7929] = layer2_outputs[5118];
    assign outputs[7930] = (layer2_outputs[11927]) & ~(layer2_outputs[9120]);
    assign outputs[7931] = ~((layer2_outputs[6236]) ^ (layer2_outputs[11728]));
    assign outputs[7932] = ~(layer2_outputs[10756]);
    assign outputs[7933] = ~(layer2_outputs[9504]);
    assign outputs[7934] = layer2_outputs[11305];
    assign outputs[7935] = ~(layer2_outputs[6439]);
    assign outputs[7936] = ~((layer2_outputs[7134]) & (layer2_outputs[8259]));
    assign outputs[7937] = ~(layer2_outputs[1465]);
    assign outputs[7938] = ~(layer2_outputs[8915]) | (layer2_outputs[837]);
    assign outputs[7939] = layer2_outputs[11572];
    assign outputs[7940] = ~((layer2_outputs[9948]) | (layer2_outputs[5190]));
    assign outputs[7941] = layer2_outputs[6687];
    assign outputs[7942] = ~(layer2_outputs[5185]) | (layer2_outputs[12503]);
    assign outputs[7943] = (layer2_outputs[10263]) & ~(layer2_outputs[7969]);
    assign outputs[7944] = layer2_outputs[5858];
    assign outputs[7945] = ~(layer2_outputs[7707]);
    assign outputs[7946] = layer2_outputs[10271];
    assign outputs[7947] = ~((layer2_outputs[12]) ^ (layer2_outputs[11977]));
    assign outputs[7948] = layer2_outputs[7316];
    assign outputs[7949] = layer2_outputs[1139];
    assign outputs[7950] = (layer2_outputs[954]) & ~(layer2_outputs[6118]);
    assign outputs[7951] = layer2_outputs[12649];
    assign outputs[7952] = layer2_outputs[9283];
    assign outputs[7953] = ~(layer2_outputs[4919]);
    assign outputs[7954] = (layer2_outputs[11572]) & ~(layer2_outputs[9880]);
    assign outputs[7955] = ~(layer2_outputs[10951]);
    assign outputs[7956] = (layer2_outputs[12521]) ^ (layer2_outputs[6576]);
    assign outputs[7957] = layer2_outputs[3481];
    assign outputs[7958] = ~(layer2_outputs[11010]);
    assign outputs[7959] = ~((layer2_outputs[3385]) ^ (layer2_outputs[1138]));
    assign outputs[7960] = ~(layer2_outputs[11129]) | (layer2_outputs[1129]);
    assign outputs[7961] = ~(layer2_outputs[4109]);
    assign outputs[7962] = layer2_outputs[2258];
    assign outputs[7963] = (layer2_outputs[12760]) & (layer2_outputs[5590]);
    assign outputs[7964] = ~(layer2_outputs[4613]);
    assign outputs[7965] = ~(layer2_outputs[5965]);
    assign outputs[7966] = (layer2_outputs[10920]) ^ (layer2_outputs[9913]);
    assign outputs[7967] = ~((layer2_outputs[11506]) ^ (layer2_outputs[4980]));
    assign outputs[7968] = ~(layer2_outputs[7967]);
    assign outputs[7969] = (layer2_outputs[6803]) & (layer2_outputs[5777]);
    assign outputs[7970] = ~((layer2_outputs[5190]) | (layer2_outputs[2048]));
    assign outputs[7971] = ~(layer2_outputs[2404]);
    assign outputs[7972] = layer2_outputs[2067];
    assign outputs[7973] = ~(layer2_outputs[1487]);
    assign outputs[7974] = layer2_outputs[10333];
    assign outputs[7975] = layer2_outputs[8858];
    assign outputs[7976] = 1'b0;
    assign outputs[7977] = ~(layer2_outputs[10766]);
    assign outputs[7978] = layer2_outputs[8661];
    assign outputs[7979] = layer2_outputs[12336];
    assign outputs[7980] = ~(layer2_outputs[8243]);
    assign outputs[7981] = layer2_outputs[4892];
    assign outputs[7982] = (layer2_outputs[10592]) ^ (layer2_outputs[7074]);
    assign outputs[7983] = ~(layer2_outputs[11978]);
    assign outputs[7984] = ~(layer2_outputs[6544]);
    assign outputs[7985] = ~(layer2_outputs[2777]);
    assign outputs[7986] = layer2_outputs[7601];
    assign outputs[7987] = layer2_outputs[10066];
    assign outputs[7988] = ~(layer2_outputs[9194]);
    assign outputs[7989] = (layer2_outputs[8854]) ^ (layer2_outputs[8028]);
    assign outputs[7990] = (layer2_outputs[11450]) & ~(layer2_outputs[5282]);
    assign outputs[7991] = (layer2_outputs[285]) & (layer2_outputs[8465]);
    assign outputs[7992] = ~(layer2_outputs[9847]);
    assign outputs[7993] = ~((layer2_outputs[3600]) & (layer2_outputs[855]));
    assign outputs[7994] = ~((layer2_outputs[8510]) ^ (layer2_outputs[8433]));
    assign outputs[7995] = layer2_outputs[10257];
    assign outputs[7996] = layer2_outputs[589];
    assign outputs[7997] = (layer2_outputs[11811]) | (layer2_outputs[9065]);
    assign outputs[7998] = (layer2_outputs[10471]) & ~(layer2_outputs[8244]);
    assign outputs[7999] = ~(layer2_outputs[5431]);
    assign outputs[8000] = (layer2_outputs[3651]) ^ (layer2_outputs[8656]);
    assign outputs[8001] = layer2_outputs[12574];
    assign outputs[8002] = layer2_outputs[11447];
    assign outputs[8003] = ~((layer2_outputs[3280]) ^ (layer2_outputs[7355]));
    assign outputs[8004] = ~(layer2_outputs[537]) | (layer2_outputs[11587]);
    assign outputs[8005] = ~(layer2_outputs[5937]);
    assign outputs[8006] = layer2_outputs[939];
    assign outputs[8007] = layer2_outputs[12044];
    assign outputs[8008] = layer2_outputs[950];
    assign outputs[8009] = (layer2_outputs[7770]) & ~(layer2_outputs[5803]);
    assign outputs[8010] = layer2_outputs[332];
    assign outputs[8011] = ~((layer2_outputs[5260]) ^ (layer2_outputs[2114]));
    assign outputs[8012] = ~((layer2_outputs[517]) | (layer2_outputs[8623]));
    assign outputs[8013] = ~(layer2_outputs[132]);
    assign outputs[8014] = ~(layer2_outputs[310]);
    assign outputs[8015] = layer2_outputs[1184];
    assign outputs[8016] = ~(layer2_outputs[2512]);
    assign outputs[8017] = layer2_outputs[4780];
    assign outputs[8018] = ~(layer2_outputs[224]);
    assign outputs[8019] = ~(layer2_outputs[746]);
    assign outputs[8020] = ~(layer2_outputs[5651]) | (layer2_outputs[6622]);
    assign outputs[8021] = ~((layer2_outputs[11481]) ^ (layer2_outputs[1993]));
    assign outputs[8022] = layer2_outputs[5293];
    assign outputs[8023] = ~(layer2_outputs[11598]);
    assign outputs[8024] = (layer2_outputs[11273]) ^ (layer2_outputs[1441]);
    assign outputs[8025] = ~(layer2_outputs[2751]) | (layer2_outputs[11063]);
    assign outputs[8026] = ~(layer2_outputs[663]);
    assign outputs[8027] = ~((layer2_outputs[4541]) ^ (layer2_outputs[5545]));
    assign outputs[8028] = layer2_outputs[6188];
    assign outputs[8029] = ~(layer2_outputs[5780]) | (layer2_outputs[9297]);
    assign outputs[8030] = ~(layer2_outputs[7671]);
    assign outputs[8031] = ~(layer2_outputs[12609]);
    assign outputs[8032] = ~(layer2_outputs[1943]);
    assign outputs[8033] = ~((layer2_outputs[7452]) ^ (layer2_outputs[3913]));
    assign outputs[8034] = ~(layer2_outputs[3451]);
    assign outputs[8035] = layer2_outputs[2910];
    assign outputs[8036] = ~(layer2_outputs[7652]);
    assign outputs[8037] = layer2_outputs[8027];
    assign outputs[8038] = ~((layer2_outputs[263]) | (layer2_outputs[12431]));
    assign outputs[8039] = layer2_outputs[11639];
    assign outputs[8040] = ~(layer2_outputs[5469]);
    assign outputs[8041] = ~(layer2_outputs[8039]);
    assign outputs[8042] = ~(layer2_outputs[8255]);
    assign outputs[8043] = (layer2_outputs[5483]) & ~(layer2_outputs[502]);
    assign outputs[8044] = layer2_outputs[8210];
    assign outputs[8045] = ~(layer2_outputs[9335]);
    assign outputs[8046] = ~(layer2_outputs[8988]);
    assign outputs[8047] = ~((layer2_outputs[7349]) | (layer2_outputs[3846]));
    assign outputs[8048] = ~(layer2_outputs[9054]);
    assign outputs[8049] = ~(layer2_outputs[1823]);
    assign outputs[8050] = layer2_outputs[1495];
    assign outputs[8051] = layer2_outputs[1311];
    assign outputs[8052] = ~(layer2_outputs[6264]);
    assign outputs[8053] = layer2_outputs[3622];
    assign outputs[8054] = ~((layer2_outputs[8271]) ^ (layer2_outputs[781]));
    assign outputs[8055] = (layer2_outputs[10077]) & ~(layer2_outputs[11379]);
    assign outputs[8056] = ~(layer2_outputs[12292]);
    assign outputs[8057] = ~(layer2_outputs[11233]);
    assign outputs[8058] = ~(layer2_outputs[6364]);
    assign outputs[8059] = (layer2_outputs[10298]) & (layer2_outputs[2018]);
    assign outputs[8060] = layer2_outputs[9740];
    assign outputs[8061] = (layer2_outputs[2534]) ^ (layer2_outputs[5425]);
    assign outputs[8062] = (layer2_outputs[7000]) & ~(layer2_outputs[2256]);
    assign outputs[8063] = ~(layer2_outputs[9121]);
    assign outputs[8064] = ~(layer2_outputs[2112]);
    assign outputs[8065] = layer2_outputs[675];
    assign outputs[8066] = ~((layer2_outputs[10365]) ^ (layer2_outputs[348]));
    assign outputs[8067] = ~(layer2_outputs[1692]);
    assign outputs[8068] = layer2_outputs[2954];
    assign outputs[8069] = ~(layer2_outputs[8998]);
    assign outputs[8070] = ~(layer2_outputs[524]);
    assign outputs[8071] = ~((layer2_outputs[9953]) & (layer2_outputs[2502]));
    assign outputs[8072] = (layer2_outputs[3944]) & (layer2_outputs[10163]);
    assign outputs[8073] = (layer2_outputs[12008]) ^ (layer2_outputs[8555]);
    assign outputs[8074] = layer2_outputs[1708];
    assign outputs[8075] = ~(layer2_outputs[7788]);
    assign outputs[8076] = (layer2_outputs[4212]) & ~(layer2_outputs[6007]);
    assign outputs[8077] = ~(layer2_outputs[5701]);
    assign outputs[8078] = layer2_outputs[4004];
    assign outputs[8079] = ~((layer2_outputs[770]) | (layer2_outputs[7259]));
    assign outputs[8080] = (layer2_outputs[8636]) ^ (layer2_outputs[7286]);
    assign outputs[8081] = ~(layer2_outputs[1949]);
    assign outputs[8082] = ~(layer2_outputs[9557]);
    assign outputs[8083] = ~(layer2_outputs[4591]);
    assign outputs[8084] = layer2_outputs[490];
    assign outputs[8085] = ~((layer2_outputs[4154]) | (layer2_outputs[3264]));
    assign outputs[8086] = layer2_outputs[10958];
    assign outputs[8087] = layer2_outputs[7470];
    assign outputs[8088] = ~(layer2_outputs[9066]);
    assign outputs[8089] = layer2_outputs[5533];
    assign outputs[8090] = (layer2_outputs[6655]) ^ (layer2_outputs[11359]);
    assign outputs[8091] = ~(layer2_outputs[9139]);
    assign outputs[8092] = (layer2_outputs[4162]) & ~(layer2_outputs[6754]);
    assign outputs[8093] = (layer2_outputs[2770]) & (layer2_outputs[3262]);
    assign outputs[8094] = ~(layer2_outputs[5822]);
    assign outputs[8095] = layer2_outputs[8903];
    assign outputs[8096] = (layer2_outputs[11220]) & ~(layer2_outputs[7455]);
    assign outputs[8097] = layer2_outputs[9961];
    assign outputs[8098] = ~((layer2_outputs[8994]) ^ (layer2_outputs[9220]));
    assign outputs[8099] = layer2_outputs[2599];
    assign outputs[8100] = ~(layer2_outputs[11462]);
    assign outputs[8101] = layer2_outputs[9240];
    assign outputs[8102] = layer2_outputs[1300];
    assign outputs[8103] = layer2_outputs[6048];
    assign outputs[8104] = ~((layer2_outputs[7518]) ^ (layer2_outputs[11976]));
    assign outputs[8105] = layer2_outputs[9158];
    assign outputs[8106] = layer2_outputs[6469];
    assign outputs[8107] = ~(layer2_outputs[12577]);
    assign outputs[8108] = ~((layer2_outputs[7604]) ^ (layer2_outputs[2731]));
    assign outputs[8109] = (layer2_outputs[12077]) ^ (layer2_outputs[6707]);
    assign outputs[8110] = layer2_outputs[779];
    assign outputs[8111] = (layer2_outputs[2862]) & (layer2_outputs[2436]);
    assign outputs[8112] = layer2_outputs[11445];
    assign outputs[8113] = ~(layer2_outputs[7761]);
    assign outputs[8114] = (layer2_outputs[7353]) & (layer2_outputs[7989]);
    assign outputs[8115] = ~((layer2_outputs[1353]) ^ (layer2_outputs[8320]));
    assign outputs[8116] = layer2_outputs[11778];
    assign outputs[8117] = layer2_outputs[2892];
    assign outputs[8118] = layer2_outputs[2577];
    assign outputs[8119] = layer2_outputs[8183];
    assign outputs[8120] = ~(layer2_outputs[2444]) | (layer2_outputs[2281]);
    assign outputs[8121] = ~(layer2_outputs[12289]);
    assign outputs[8122] = ~((layer2_outputs[4199]) ^ (layer2_outputs[12047]));
    assign outputs[8123] = ~(layer2_outputs[5229]);
    assign outputs[8124] = (layer2_outputs[6213]) ^ (layer2_outputs[7476]);
    assign outputs[8125] = (layer2_outputs[7302]) & ~(layer2_outputs[10723]);
    assign outputs[8126] = ~(layer2_outputs[1081]);
    assign outputs[8127] = ~((layer2_outputs[2967]) ^ (layer2_outputs[5314]));
    assign outputs[8128] = ~(layer2_outputs[9875]);
    assign outputs[8129] = ~(layer2_outputs[2632]);
    assign outputs[8130] = layer2_outputs[12694];
    assign outputs[8131] = layer2_outputs[6144];
    assign outputs[8132] = (layer2_outputs[10619]) & ~(layer2_outputs[10778]);
    assign outputs[8133] = (layer2_outputs[8147]) & (layer2_outputs[8691]);
    assign outputs[8134] = (layer2_outputs[629]) & ~(layer2_outputs[4549]);
    assign outputs[8135] = ~((layer2_outputs[3314]) | (layer2_outputs[111]));
    assign outputs[8136] = ~(layer2_outputs[1406]);
    assign outputs[8137] = ~(layer2_outputs[10567]);
    assign outputs[8138] = ~(layer2_outputs[5087]);
    assign outputs[8139] = ~(layer2_outputs[7972]);
    assign outputs[8140] = ~(layer2_outputs[8293]);
    assign outputs[8141] = layer2_outputs[4832];
    assign outputs[8142] = ~((layer2_outputs[6388]) ^ (layer2_outputs[1271]));
    assign outputs[8143] = (layer2_outputs[9723]) & ~(layer2_outputs[11341]);
    assign outputs[8144] = ~(layer2_outputs[3599]);
    assign outputs[8145] = (layer2_outputs[1061]) & ~(layer2_outputs[12383]);
    assign outputs[8146] = layer2_outputs[4569];
    assign outputs[8147] = ~(layer2_outputs[4049]);
    assign outputs[8148] = ~(layer2_outputs[10516]);
    assign outputs[8149] = layer2_outputs[3488];
    assign outputs[8150] = layer2_outputs[8948];
    assign outputs[8151] = ~(layer2_outputs[3269]);
    assign outputs[8152] = layer2_outputs[6887];
    assign outputs[8153] = ~(layer2_outputs[11537]);
    assign outputs[8154] = (layer2_outputs[1625]) & ~(layer2_outputs[5]);
    assign outputs[8155] = ~(layer2_outputs[5484]);
    assign outputs[8156] = ~(layer2_outputs[4545]);
    assign outputs[8157] = layer2_outputs[2440];
    assign outputs[8158] = ~((layer2_outputs[9984]) ^ (layer2_outputs[1350]));
    assign outputs[8159] = ~(layer2_outputs[7167]);
    assign outputs[8160] = (layer2_outputs[10289]) | (layer2_outputs[8562]);
    assign outputs[8161] = ~(layer2_outputs[4605]);
    assign outputs[8162] = ~(layer2_outputs[942]);
    assign outputs[8163] = ~(layer2_outputs[823]);
    assign outputs[8164] = (layer2_outputs[5912]) & ~(layer2_outputs[12416]);
    assign outputs[8165] = ~(layer2_outputs[7438]);
    assign outputs[8166] = ~(layer2_outputs[454]);
    assign outputs[8167] = ~((layer2_outputs[9213]) | (layer2_outputs[3494]));
    assign outputs[8168] = ~(layer2_outputs[7810]);
    assign outputs[8169] = ~(layer2_outputs[10555]) | (layer2_outputs[3288]);
    assign outputs[8170] = ~(layer2_outputs[4149]);
    assign outputs[8171] = layer2_outputs[5529];
    assign outputs[8172] = ~((layer2_outputs[2519]) & (layer2_outputs[12748]));
    assign outputs[8173] = layer2_outputs[9474];
    assign outputs[8174] = layer2_outputs[8157];
    assign outputs[8175] = ~(layer2_outputs[10673]);
    assign outputs[8176] = (layer2_outputs[3485]) & ~(layer2_outputs[2366]);
    assign outputs[8177] = ~(layer2_outputs[212]);
    assign outputs[8178] = layer2_outputs[4748];
    assign outputs[8179] = (layer2_outputs[9306]) ^ (layer2_outputs[10399]);
    assign outputs[8180] = ~(layer2_outputs[6230]);
    assign outputs[8181] = (layer2_outputs[3779]) ^ (layer2_outputs[12431]);
    assign outputs[8182] = ~(layer2_outputs[12192]);
    assign outputs[8183] = ~(layer2_outputs[6885]) | (layer2_outputs[12375]);
    assign outputs[8184] = ~((layer2_outputs[1415]) | (layer2_outputs[2209]));
    assign outputs[8185] = ~(layer2_outputs[4766]);
    assign outputs[8186] = layer2_outputs[3635];
    assign outputs[8187] = layer2_outputs[7080];
    assign outputs[8188] = (layer2_outputs[1852]) & ~(layer2_outputs[11730]);
    assign outputs[8189] = ~((layer2_outputs[1197]) ^ (layer2_outputs[7785]));
    assign outputs[8190] = ~(layer2_outputs[1663]);
    assign outputs[8191] = layer2_outputs[1067];
    assign outputs[8192] = ~(layer2_outputs[511]);
    assign outputs[8193] = (layer2_outputs[6923]) & (layer2_outputs[7058]);
    assign outputs[8194] = layer2_outputs[1622];
    assign outputs[8195] = (layer2_outputs[12570]) ^ (layer2_outputs[10538]);
    assign outputs[8196] = ~(layer2_outputs[8707]);
    assign outputs[8197] = layer2_outputs[2645];
    assign outputs[8198] = ~((layer2_outputs[3803]) ^ (layer2_outputs[11008]));
    assign outputs[8199] = ~(layer2_outputs[605]);
    assign outputs[8200] = layer2_outputs[8134];
    assign outputs[8201] = ~(layer2_outputs[4419]);
    assign outputs[8202] = (layer2_outputs[2332]) ^ (layer2_outputs[11240]);
    assign outputs[8203] = ~(layer2_outputs[6222]);
    assign outputs[8204] = ~((layer2_outputs[3629]) ^ (layer2_outputs[2037]));
    assign outputs[8205] = (layer2_outputs[7104]) & ~(layer2_outputs[10723]);
    assign outputs[8206] = ~(layer2_outputs[5691]);
    assign outputs[8207] = ~((layer2_outputs[978]) ^ (layer2_outputs[1230]));
    assign outputs[8208] = layer2_outputs[10330];
    assign outputs[8209] = layer2_outputs[9830];
    assign outputs[8210] = ~((layer2_outputs[4541]) ^ (layer2_outputs[1307]));
    assign outputs[8211] = ~((layer2_outputs[12110]) ^ (layer2_outputs[887]));
    assign outputs[8212] = (layer2_outputs[7383]) & ~(layer2_outputs[8430]);
    assign outputs[8213] = layer2_outputs[11740];
    assign outputs[8214] = (layer2_outputs[12308]) | (layer2_outputs[1829]);
    assign outputs[8215] = (layer2_outputs[1938]) ^ (layer2_outputs[5013]);
    assign outputs[8216] = layer2_outputs[1472];
    assign outputs[8217] = ~(layer2_outputs[5736]);
    assign outputs[8218] = (layer2_outputs[3864]) ^ (layer2_outputs[5702]);
    assign outputs[8219] = layer2_outputs[4815];
    assign outputs[8220] = ~(layer2_outputs[7448]);
    assign outputs[8221] = ~((layer2_outputs[10699]) ^ (layer2_outputs[2810]));
    assign outputs[8222] = ~(layer2_outputs[2657]);
    assign outputs[8223] = ~(layer2_outputs[10999]);
    assign outputs[8224] = layer2_outputs[11697];
    assign outputs[8225] = layer2_outputs[5660];
    assign outputs[8226] = ~(layer2_outputs[1182]);
    assign outputs[8227] = ~(layer2_outputs[8991]);
    assign outputs[8228] = ~((layer2_outputs[8737]) ^ (layer2_outputs[768]));
    assign outputs[8229] = ~(layer2_outputs[5244]);
    assign outputs[8230] = (layer2_outputs[4976]) & (layer2_outputs[6016]);
    assign outputs[8231] = layer2_outputs[3172];
    assign outputs[8232] = ~(layer2_outputs[10518]);
    assign outputs[8233] = layer2_outputs[6262];
    assign outputs[8234] = layer2_outputs[9021];
    assign outputs[8235] = ~((layer2_outputs[6503]) & (layer2_outputs[8154]));
    assign outputs[8236] = layer2_outputs[2044];
    assign outputs[8237] = (layer2_outputs[5213]) | (layer2_outputs[12182]);
    assign outputs[8238] = layer2_outputs[6189];
    assign outputs[8239] = ~(layer2_outputs[10349]);
    assign outputs[8240] = ~(layer2_outputs[4796]);
    assign outputs[8241] = ~(layer2_outputs[3619]);
    assign outputs[8242] = ~(layer2_outputs[1778]);
    assign outputs[8243] = layer2_outputs[9208];
    assign outputs[8244] = (layer2_outputs[2531]) & (layer2_outputs[3645]);
    assign outputs[8245] = layer2_outputs[9175];
    assign outputs[8246] = ~((layer2_outputs[880]) ^ (layer2_outputs[1693]));
    assign outputs[8247] = ~(layer2_outputs[7769]);
    assign outputs[8248] = ~(layer2_outputs[4035]);
    assign outputs[8249] = (layer2_outputs[7471]) & (layer2_outputs[10373]);
    assign outputs[8250] = ~(layer2_outputs[2794]);
    assign outputs[8251] = ~(layer2_outputs[12607]);
    assign outputs[8252] = ~(layer2_outputs[2030]);
    assign outputs[8253] = ~(layer2_outputs[4123]);
    assign outputs[8254] = ~(layer2_outputs[4542]);
    assign outputs[8255] = ~(layer2_outputs[10765]);
    assign outputs[8256] = layer2_outputs[2580];
    assign outputs[8257] = (layer2_outputs[12010]) | (layer2_outputs[1084]);
    assign outputs[8258] = layer2_outputs[1988];
    assign outputs[8259] = ~((layer2_outputs[12323]) & (layer2_outputs[8777]));
    assign outputs[8260] = ~((layer2_outputs[1705]) ^ (layer2_outputs[5120]));
    assign outputs[8261] = ~(layer2_outputs[7315]);
    assign outputs[8262] = layer2_outputs[1449];
    assign outputs[8263] = ~(layer2_outputs[2906]);
    assign outputs[8264] = layer2_outputs[10266];
    assign outputs[8265] = ~(layer2_outputs[12088]);
    assign outputs[8266] = layer2_outputs[4576];
    assign outputs[8267] = ~(layer2_outputs[5560]);
    assign outputs[8268] = layer2_outputs[3882];
    assign outputs[8269] = ~((layer2_outputs[2446]) ^ (layer2_outputs[12362]));
    assign outputs[8270] = (layer2_outputs[6524]) & (layer2_outputs[6573]);
    assign outputs[8271] = ~(layer2_outputs[9458]);
    assign outputs[8272] = ~(layer2_outputs[2521]);
    assign outputs[8273] = ~((layer2_outputs[5562]) | (layer2_outputs[9009]));
    assign outputs[8274] = (layer2_outputs[6155]) ^ (layer2_outputs[1193]);
    assign outputs[8275] = ~(layer2_outputs[6353]);
    assign outputs[8276] = ~((layer2_outputs[11000]) ^ (layer2_outputs[9180]));
    assign outputs[8277] = ~(layer2_outputs[7821]);
    assign outputs[8278] = layer2_outputs[589];
    assign outputs[8279] = (layer2_outputs[4127]) & ~(layer2_outputs[3714]);
    assign outputs[8280] = ~(layer2_outputs[5254]);
    assign outputs[8281] = (layer2_outputs[10293]) ^ (layer2_outputs[2457]);
    assign outputs[8282] = layer2_outputs[2962];
    assign outputs[8283] = layer2_outputs[4681];
    assign outputs[8284] = (layer2_outputs[651]) & ~(layer2_outputs[2660]);
    assign outputs[8285] = ~(layer2_outputs[6860]);
    assign outputs[8286] = (layer2_outputs[476]) ^ (layer2_outputs[10886]);
    assign outputs[8287] = layer2_outputs[6330];
    assign outputs[8288] = layer2_outputs[11931];
    assign outputs[8289] = layer2_outputs[11578];
    assign outputs[8290] = ~(layer2_outputs[5910]);
    assign outputs[8291] = ~(layer2_outputs[6883]);
    assign outputs[8292] = ~(layer2_outputs[1060]);
    assign outputs[8293] = ~((layer2_outputs[2604]) ^ (layer2_outputs[3885]));
    assign outputs[8294] = (layer2_outputs[6359]) & ~(layer2_outputs[4820]);
    assign outputs[8295] = (layer2_outputs[1064]) ^ (layer2_outputs[10554]);
    assign outputs[8296] = ~(layer2_outputs[8478]);
    assign outputs[8297] = layer2_outputs[351];
    assign outputs[8298] = (layer2_outputs[7135]) & ~(layer2_outputs[6494]);
    assign outputs[8299] = ~(layer2_outputs[1238]);
    assign outputs[8300] = layer2_outputs[8283];
    assign outputs[8301] = (layer2_outputs[4357]) & ~(layer2_outputs[5316]);
    assign outputs[8302] = (layer2_outputs[2876]) ^ (layer2_outputs[3931]);
    assign outputs[8303] = ~(layer2_outputs[7716]) | (layer2_outputs[11038]);
    assign outputs[8304] = ~((layer2_outputs[2289]) ^ (layer2_outputs[8743]));
    assign outputs[8305] = layer2_outputs[7095];
    assign outputs[8306] = ~(layer2_outputs[5276]);
    assign outputs[8307] = ~((layer2_outputs[3031]) ^ (layer2_outputs[8316]));
    assign outputs[8308] = layer2_outputs[11516];
    assign outputs[8309] = ~(layer2_outputs[2148]);
    assign outputs[8310] = ~(layer2_outputs[5562]);
    assign outputs[8311] = ~(layer2_outputs[9910]);
    assign outputs[8312] = layer2_outputs[3839];
    assign outputs[8313] = (layer2_outputs[782]) & (layer2_outputs[9739]);
    assign outputs[8314] = ~(layer2_outputs[4647]);
    assign outputs[8315] = ~(layer2_outputs[7569]);
    assign outputs[8316] = ~((layer2_outputs[10674]) ^ (layer2_outputs[12640]));
    assign outputs[8317] = ~(layer2_outputs[7057]);
    assign outputs[8318] = (layer2_outputs[10086]) ^ (layer2_outputs[77]);
    assign outputs[8319] = ~(layer2_outputs[9344]);
    assign outputs[8320] = ~(layer2_outputs[5917]);
    assign outputs[8321] = layer2_outputs[9675];
    assign outputs[8322] = (layer2_outputs[5886]) & ~(layer2_outputs[4793]);
    assign outputs[8323] = layer2_outputs[5606];
    assign outputs[8324] = ~(layer2_outputs[10780]);
    assign outputs[8325] = layer2_outputs[6818];
    assign outputs[8326] = (layer2_outputs[1]) ^ (layer2_outputs[6829]);
    assign outputs[8327] = ~(layer2_outputs[8023]);
    assign outputs[8328] = ~((layer2_outputs[12341]) ^ (layer2_outputs[1039]));
    assign outputs[8329] = (layer2_outputs[5207]) & ~(layer2_outputs[3557]);
    assign outputs[8330] = ~(layer2_outputs[3085]);
    assign outputs[8331] = layer2_outputs[6047];
    assign outputs[8332] = ~((layer2_outputs[194]) ^ (layer2_outputs[6147]));
    assign outputs[8333] = (layer2_outputs[1902]) ^ (layer2_outputs[5020]);
    assign outputs[8334] = layer2_outputs[5679];
    assign outputs[8335] = ~(layer2_outputs[5080]);
    assign outputs[8336] = ~(layer2_outputs[553]);
    assign outputs[8337] = ~(layer2_outputs[3415]);
    assign outputs[8338] = ~(layer2_outputs[2450]) | (layer2_outputs[10547]);
    assign outputs[8339] = layer2_outputs[9812];
    assign outputs[8340] = ~(layer2_outputs[10479]);
    assign outputs[8341] = ~((layer2_outputs[12394]) | (layer2_outputs[8015]));
    assign outputs[8342] = layer2_outputs[9790];
    assign outputs[8343] = layer2_outputs[7642];
    assign outputs[8344] = ~((layer2_outputs[12175]) | (layer2_outputs[172]));
    assign outputs[8345] = ~(layer2_outputs[8652]);
    assign outputs[8346] = (layer2_outputs[10693]) & ~(layer2_outputs[7800]);
    assign outputs[8347] = ~(layer2_outputs[8208]);
    assign outputs[8348] = ~((layer2_outputs[6656]) | (layer2_outputs[7559]));
    assign outputs[8349] = (layer2_outputs[8180]) & ~(layer2_outputs[3145]);
    assign outputs[8350] = ~(layer2_outputs[2385]);
    assign outputs[8351] = (layer2_outputs[6194]) ^ (layer2_outputs[3142]);
    assign outputs[8352] = ~(layer2_outputs[12363]) | (layer2_outputs[10005]);
    assign outputs[8353] = ~(layer2_outputs[411]);
    assign outputs[8354] = ~((layer2_outputs[2490]) ^ (layer2_outputs[8202]));
    assign outputs[8355] = ~(layer2_outputs[7121]);
    assign outputs[8356] = (layer2_outputs[499]) & (layer2_outputs[3258]);
    assign outputs[8357] = ~(layer2_outputs[9670]);
    assign outputs[8358] = layer2_outputs[6428];
    assign outputs[8359] = layer2_outputs[10738];
    assign outputs[8360] = ~(layer2_outputs[1109]);
    assign outputs[8361] = ~(layer2_outputs[4128]);
    assign outputs[8362] = ~(layer2_outputs[5172]);
    assign outputs[8363] = layer2_outputs[451];
    assign outputs[8364] = layer2_outputs[7709];
    assign outputs[8365] = ~(layer2_outputs[98]);
    assign outputs[8366] = ~(layer2_outputs[2652]);
    assign outputs[8367] = layer2_outputs[9894];
    assign outputs[8368] = (layer2_outputs[8198]) & (layer2_outputs[2996]);
    assign outputs[8369] = (layer2_outputs[11683]) & ~(layer2_outputs[11808]);
    assign outputs[8370] = layer2_outputs[7809];
    assign outputs[8371] = (layer2_outputs[7407]) & ~(layer2_outputs[5183]);
    assign outputs[8372] = (layer2_outputs[632]) ^ (layer2_outputs[12237]);
    assign outputs[8373] = ~(layer2_outputs[6185]);
    assign outputs[8374] = ~(layer2_outputs[2738]);
    assign outputs[8375] = layer2_outputs[10636];
    assign outputs[8376] = (layer2_outputs[7672]) & ~(layer2_outputs[2551]);
    assign outputs[8377] = (layer2_outputs[17]) & ~(layer2_outputs[5007]);
    assign outputs[8378] = ~(layer2_outputs[10837]);
    assign outputs[8379] = (layer2_outputs[641]) & ~(layer2_outputs[11810]);
    assign outputs[8380] = (layer2_outputs[1651]) & ~(layer2_outputs[8276]);
    assign outputs[8381] = layer2_outputs[11540];
    assign outputs[8382] = ~(layer2_outputs[3118]);
    assign outputs[8383] = ~(layer2_outputs[2758]);
    assign outputs[8384] = layer2_outputs[3862];
    assign outputs[8385] = ~(layer2_outputs[10167]);
    assign outputs[8386] = (layer2_outputs[3530]) ^ (layer2_outputs[8402]);
    assign outputs[8387] = (layer2_outputs[11804]) & ~(layer2_outputs[10850]);
    assign outputs[8388] = (layer2_outputs[8830]) & ~(layer2_outputs[1892]);
    assign outputs[8389] = ~((layer2_outputs[10315]) & (layer2_outputs[9018]));
    assign outputs[8390] = (layer2_outputs[1225]) ^ (layer2_outputs[3110]);
    assign outputs[8391] = layer2_outputs[1390];
    assign outputs[8392] = ~(layer2_outputs[7158]);
    assign outputs[8393] = ~(layer2_outputs[8471]);
    assign outputs[8394] = layer2_outputs[9621];
    assign outputs[8395] = (layer2_outputs[5749]) & (layer2_outputs[6215]);
    assign outputs[8396] = (layer2_outputs[2190]) ^ (layer2_outputs[1467]);
    assign outputs[8397] = layer2_outputs[11289];
    assign outputs[8398] = ~(layer2_outputs[1116]);
    assign outputs[8399] = ~(layer2_outputs[383]);
    assign outputs[8400] = ~(layer2_outputs[1631]);
    assign outputs[8401] = ~(layer2_outputs[2328]);
    assign outputs[8402] = ~(layer2_outputs[7204]) | (layer2_outputs[3660]);
    assign outputs[8403] = (layer2_outputs[6354]) ^ (layer2_outputs[9705]);
    assign outputs[8404] = (layer2_outputs[10471]) & ~(layer2_outputs[5624]);
    assign outputs[8405] = (layer2_outputs[12028]) & ~(layer2_outputs[6705]);
    assign outputs[8406] = ~(layer2_outputs[12443]);
    assign outputs[8407] = (layer2_outputs[8267]) ^ (layer2_outputs[12236]);
    assign outputs[8408] = ~(layer2_outputs[10305]);
    assign outputs[8409] = (layer2_outputs[12279]) & (layer2_outputs[5391]);
    assign outputs[8410] = layer2_outputs[2401];
    assign outputs[8411] = ~((layer2_outputs[2638]) ^ (layer2_outputs[11224]));
    assign outputs[8412] = ~(layer2_outputs[11553]);
    assign outputs[8413] = ~(layer2_outputs[7860]);
    assign outputs[8414] = layer2_outputs[10634];
    assign outputs[8415] = ~((layer2_outputs[9547]) ^ (layer2_outputs[532]));
    assign outputs[8416] = ~((layer2_outputs[5466]) ^ (layer2_outputs[6718]));
    assign outputs[8417] = layer2_outputs[7065];
    assign outputs[8418] = ~((layer2_outputs[9092]) ^ (layer2_outputs[7515]));
    assign outputs[8419] = ~((layer2_outputs[8322]) & (layer2_outputs[8272]));
    assign outputs[8420] = layer2_outputs[259];
    assign outputs[8421] = ~(layer2_outputs[7157]);
    assign outputs[8422] = (layer2_outputs[3395]) ^ (layer2_outputs[734]);
    assign outputs[8423] = layer2_outputs[10734];
    assign outputs[8424] = (layer2_outputs[337]) & ~(layer2_outputs[11165]);
    assign outputs[8425] = ~(layer2_outputs[8496]) | (layer2_outputs[1148]);
    assign outputs[8426] = layer2_outputs[4903];
    assign outputs[8427] = ~(layer2_outputs[10224]) | (layer2_outputs[1058]);
    assign outputs[8428] = layer2_outputs[12784];
    assign outputs[8429] = ~(layer2_outputs[1663]) | (layer2_outputs[6028]);
    assign outputs[8430] = ~((layer2_outputs[6594]) ^ (layer2_outputs[345]));
    assign outputs[8431] = (layer2_outputs[578]) & ~(layer2_outputs[11107]);
    assign outputs[8432] = (layer2_outputs[4858]) & (layer2_outputs[11509]);
    assign outputs[8433] = ~(layer2_outputs[2613]);
    assign outputs[8434] = (layer2_outputs[8434]) & ~(layer2_outputs[5926]);
    assign outputs[8435] = ~(layer2_outputs[5056]);
    assign outputs[8436] = layer2_outputs[4479];
    assign outputs[8437] = (layer2_outputs[4925]) | (layer2_outputs[6800]);
    assign outputs[8438] = (layer2_outputs[3256]) & (layer2_outputs[2541]);
    assign outputs[8439] = (layer2_outputs[6776]) & (layer2_outputs[3946]);
    assign outputs[8440] = layer2_outputs[11118];
    assign outputs[8441] = (layer2_outputs[12319]) ^ (layer2_outputs[6322]);
    assign outputs[8442] = ~(layer2_outputs[12401]) | (layer2_outputs[12614]);
    assign outputs[8443] = ~((layer2_outputs[12266]) ^ (layer2_outputs[2213]));
    assign outputs[8444] = ~(layer2_outputs[6394]);
    assign outputs[8445] = layer2_outputs[10353];
    assign outputs[8446] = ~(layer2_outputs[9689]);
    assign outputs[8447] = (layer2_outputs[8664]) & (layer2_outputs[2698]);
    assign outputs[8448] = layer2_outputs[9889];
    assign outputs[8449] = ~((layer2_outputs[5038]) ^ (layer2_outputs[11934]));
    assign outputs[8450] = ~(layer2_outputs[9323]);
    assign outputs[8451] = (layer2_outputs[5577]) ^ (layer2_outputs[9300]);
    assign outputs[8452] = (layer2_outputs[6596]) & (layer2_outputs[7768]);
    assign outputs[8453] = layer2_outputs[7534];
    assign outputs[8454] = (layer2_outputs[7522]) & ~(layer2_outputs[9235]);
    assign outputs[8455] = ~(layer2_outputs[4657]);
    assign outputs[8456] = ~(layer2_outputs[5223]) | (layer2_outputs[1610]);
    assign outputs[8457] = ~(layer2_outputs[6641]) | (layer2_outputs[10674]);
    assign outputs[8458] = (layer2_outputs[12628]) ^ (layer2_outputs[7684]);
    assign outputs[8459] = ~(layer2_outputs[776]);
    assign outputs[8460] = ~(layer2_outputs[12719]);
    assign outputs[8461] = layer2_outputs[5191];
    assign outputs[8462] = ~((layer2_outputs[1210]) ^ (layer2_outputs[11210]));
    assign outputs[8463] = layer2_outputs[1080];
    assign outputs[8464] = (layer2_outputs[3994]) & (layer2_outputs[9476]);
    assign outputs[8465] = layer2_outputs[6330];
    assign outputs[8466] = ~(layer2_outputs[4851]);
    assign outputs[8467] = ~(layer2_outputs[7563]);
    assign outputs[8468] = (layer2_outputs[9354]) & ~(layer2_outputs[10568]);
    assign outputs[8469] = layer2_outputs[5203];
    assign outputs[8470] = layer2_outputs[2577];
    assign outputs[8471] = (layer2_outputs[12515]) & ~(layer2_outputs[999]);
    assign outputs[8472] = ~(layer2_outputs[12392]);
    assign outputs[8473] = layer2_outputs[2670];
    assign outputs[8474] = (layer2_outputs[2170]) ^ (layer2_outputs[4337]);
    assign outputs[8475] = ~(layer2_outputs[5595]);
    assign outputs[8476] = layer2_outputs[5967];
    assign outputs[8477] = ~(layer2_outputs[6015]);
    assign outputs[8478] = layer2_outputs[4459];
    assign outputs[8479] = layer2_outputs[3192];
    assign outputs[8480] = ~(layer2_outputs[1335]);
    assign outputs[8481] = (layer2_outputs[5877]) ^ (layer2_outputs[8881]);
    assign outputs[8482] = (layer2_outputs[6880]) ^ (layer2_outputs[4509]);
    assign outputs[8483] = layer2_outputs[9119];
    assign outputs[8484] = layer2_outputs[3535];
    assign outputs[8485] = ~(layer2_outputs[6456]);
    assign outputs[8486] = ~(layer2_outputs[11246]);
    assign outputs[8487] = ~(layer2_outputs[2407]) | (layer2_outputs[12174]);
    assign outputs[8488] = (layer2_outputs[609]) ^ (layer2_outputs[10324]);
    assign outputs[8489] = layer2_outputs[2812];
    assign outputs[8490] = ~(layer2_outputs[6862]);
    assign outputs[8491] = ~(layer2_outputs[770]);
    assign outputs[8492] = layer2_outputs[2498];
    assign outputs[8493] = ~((layer2_outputs[2668]) ^ (layer2_outputs[10911]));
    assign outputs[8494] = ~((layer2_outputs[1944]) ^ (layer2_outputs[10287]));
    assign outputs[8495] = ~((layer2_outputs[12136]) | (layer2_outputs[993]));
    assign outputs[8496] = ~(layer2_outputs[543]);
    assign outputs[8497] = (layer2_outputs[1416]) ^ (layer2_outputs[4589]);
    assign outputs[8498] = ~(layer2_outputs[4478]);
    assign outputs[8499] = (layer2_outputs[10257]) ^ (layer2_outputs[9438]);
    assign outputs[8500] = (layer2_outputs[5466]) & (layer2_outputs[4116]);
    assign outputs[8501] = ~(layer2_outputs[9436]);
    assign outputs[8502] = (layer2_outputs[1630]) | (layer2_outputs[5602]);
    assign outputs[8503] = ~(layer2_outputs[2159]);
    assign outputs[8504] = (layer2_outputs[69]) & ~(layer2_outputs[10131]);
    assign outputs[8505] = ~(layer2_outputs[11403]);
    assign outputs[8506] = (layer2_outputs[683]) & (layer2_outputs[155]);
    assign outputs[8507] = ~((layer2_outputs[6598]) ^ (layer2_outputs[7259]));
    assign outputs[8508] = ~((layer2_outputs[5511]) ^ (layer2_outputs[1650]));
    assign outputs[8509] = ~(layer2_outputs[11535]);
    assign outputs[8510] = layer2_outputs[2560];
    assign outputs[8511] = (layer2_outputs[5833]) ^ (layer2_outputs[3652]);
    assign outputs[8512] = ~(layer2_outputs[3254]);
    assign outputs[8513] = layer2_outputs[8677];
    assign outputs[8514] = ~((layer2_outputs[719]) ^ (layer2_outputs[1305]));
    assign outputs[8515] = layer2_outputs[3561];
    assign outputs[8516] = layer2_outputs[7285];
    assign outputs[8517] = layer2_outputs[3839];
    assign outputs[8518] = ~((layer2_outputs[5665]) ^ (layer2_outputs[3388]));
    assign outputs[8519] = (layer2_outputs[3867]) ^ (layer2_outputs[11726]);
    assign outputs[8520] = ~((layer2_outputs[6674]) ^ (layer2_outputs[11775]));
    assign outputs[8521] = layer2_outputs[10928];
    assign outputs[8522] = (layer2_outputs[6087]) & ~(layer2_outputs[9971]);
    assign outputs[8523] = ~(layer2_outputs[7795]);
    assign outputs[8524] = ~(layer2_outputs[2488]);
    assign outputs[8525] = ~(layer2_outputs[7368]);
    assign outputs[8526] = (layer2_outputs[2327]) ^ (layer2_outputs[3284]);
    assign outputs[8527] = layer2_outputs[11427];
    assign outputs[8528] = layer2_outputs[11931];
    assign outputs[8529] = layer2_outputs[5094];
    assign outputs[8530] = (layer2_outputs[12435]) ^ (layer2_outputs[6324]);
    assign outputs[8531] = ~(layer2_outputs[9350]) | (layer2_outputs[11333]);
    assign outputs[8532] = layer2_outputs[4705];
    assign outputs[8533] = ~(layer2_outputs[12693]);
    assign outputs[8534] = (layer2_outputs[9697]) ^ (layer2_outputs[8904]);
    assign outputs[8535] = layer2_outputs[1689];
    assign outputs[8536] = ~(layer2_outputs[6703]) | (layer2_outputs[7395]);
    assign outputs[8537] = layer2_outputs[3308];
    assign outputs[8538] = layer2_outputs[853];
    assign outputs[8539] = layer2_outputs[4705];
    assign outputs[8540] = (layer2_outputs[10501]) & (layer2_outputs[7875]);
    assign outputs[8541] = ~((layer2_outputs[12615]) ^ (layer2_outputs[8630]));
    assign outputs[8542] = (layer2_outputs[867]) & (layer2_outputs[8934]);
    assign outputs[8543] = layer2_outputs[9091];
    assign outputs[8544] = ~(layer2_outputs[10189]);
    assign outputs[8545] = layer2_outputs[7196];
    assign outputs[8546] = ~((layer2_outputs[11161]) | (layer2_outputs[10391]));
    assign outputs[8547] = ~(layer2_outputs[1152]);
    assign outputs[8548] = (layer2_outputs[12214]) & ~(layer2_outputs[9975]);
    assign outputs[8549] = ~((layer2_outputs[929]) ^ (layer2_outputs[6784]));
    assign outputs[8550] = layer2_outputs[8843];
    assign outputs[8551] = ~(layer2_outputs[10659]);
    assign outputs[8552] = layer2_outputs[427];
    assign outputs[8553] = ~(layer2_outputs[10623]);
    assign outputs[8554] = layer2_outputs[7078];
    assign outputs[8555] = ~(layer2_outputs[4434]);
    assign outputs[8556] = (layer2_outputs[3757]) ^ (layer2_outputs[7955]);
    assign outputs[8557] = ~(layer2_outputs[3609]);
    assign outputs[8558] = (layer2_outputs[39]) & ~(layer2_outputs[3450]);
    assign outputs[8559] = (layer2_outputs[5070]) & (layer2_outputs[11301]);
    assign outputs[8560] = ~((layer2_outputs[10592]) ^ (layer2_outputs[2589]));
    assign outputs[8561] = ~((layer2_outputs[1215]) ^ (layer2_outputs[6888]));
    assign outputs[8562] = layer2_outputs[2212];
    assign outputs[8563] = ~(layer2_outputs[11260]);
    assign outputs[8564] = ~(layer2_outputs[7288]);
    assign outputs[8565] = (layer2_outputs[6024]) & (layer2_outputs[12739]);
    assign outputs[8566] = (layer2_outputs[11479]) ^ (layer2_outputs[10462]);
    assign outputs[8567] = layer2_outputs[3231];
    assign outputs[8568] = layer2_outputs[11274];
    assign outputs[8569] = ~(layer2_outputs[5459]);
    assign outputs[8570] = ~((layer2_outputs[12510]) | (layer2_outputs[5914]));
    assign outputs[8571] = layer2_outputs[764];
    assign outputs[8572] = ~((layer2_outputs[2614]) & (layer2_outputs[8387]));
    assign outputs[8573] = ~(layer2_outputs[7553]) | (layer2_outputs[10473]);
    assign outputs[8574] = (layer2_outputs[1566]) & ~(layer2_outputs[6475]);
    assign outputs[8575] = ~(layer2_outputs[7235]) | (layer2_outputs[5905]);
    assign outputs[8576] = ~(layer2_outputs[8558]);
    assign outputs[8577] = (layer2_outputs[5803]) ^ (layer2_outputs[687]);
    assign outputs[8578] = ~(layer2_outputs[168]) | (layer2_outputs[34]);
    assign outputs[8579] = ~(layer2_outputs[6840]);
    assign outputs[8580] = ~(layer2_outputs[10552]);
    assign outputs[8581] = (layer2_outputs[9]) & (layer2_outputs[5979]);
    assign outputs[8582] = (layer2_outputs[12142]) ^ (layer2_outputs[1481]);
    assign outputs[8583] = (layer2_outputs[1939]) | (layer2_outputs[9597]);
    assign outputs[8584] = (layer2_outputs[8604]) & ~(layer2_outputs[1543]);
    assign outputs[8585] = (layer2_outputs[9068]) & (layer2_outputs[12117]);
    assign outputs[8586] = layer2_outputs[11583];
    assign outputs[8587] = ~(layer2_outputs[7916]);
    assign outputs[8588] = (layer2_outputs[1187]) ^ (layer2_outputs[11687]);
    assign outputs[8589] = ~(layer2_outputs[1191]);
    assign outputs[8590] = ~(layer2_outputs[3801]);
    assign outputs[8591] = ~(layer2_outputs[10068]);
    assign outputs[8592] = layer2_outputs[11118];
    assign outputs[8593] = ~(layer2_outputs[575]);
    assign outputs[8594] = layer2_outputs[3400];
    assign outputs[8595] = layer2_outputs[5449];
    assign outputs[8596] = (layer2_outputs[4280]) & (layer2_outputs[3459]);
    assign outputs[8597] = layer2_outputs[2933];
    assign outputs[8598] = ~(layer2_outputs[5482]);
    assign outputs[8599] = layer2_outputs[5958];
    assign outputs[8600] = layer2_outputs[11302];
    assign outputs[8601] = layer2_outputs[9602];
    assign outputs[8602] = ~(layer2_outputs[7998]);
    assign outputs[8603] = ~((layer2_outputs[8928]) ^ (layer2_outputs[10625]));
    assign outputs[8604] = layer2_outputs[12364];
    assign outputs[8605] = (layer2_outputs[9682]) & ~(layer2_outputs[9053]);
    assign outputs[8606] = ~(layer2_outputs[1554]);
    assign outputs[8607] = ~((layer2_outputs[2291]) ^ (layer2_outputs[8824]));
    assign outputs[8608] = layer2_outputs[6025];
    assign outputs[8609] = (layer2_outputs[11092]) ^ (layer2_outputs[12633]);
    assign outputs[8610] = ~((layer2_outputs[9942]) & (layer2_outputs[1838]));
    assign outputs[8611] = layer2_outputs[187];
    assign outputs[8612] = layer2_outputs[9160];
    assign outputs[8613] = layer2_outputs[5830];
    assign outputs[8614] = ~((layer2_outputs[4003]) | (layer2_outputs[9610]));
    assign outputs[8615] = ~(layer2_outputs[3970]);
    assign outputs[8616] = layer2_outputs[6374];
    assign outputs[8617] = ~(layer2_outputs[3542]);
    assign outputs[8618] = ~((layer2_outputs[4449]) ^ (layer2_outputs[1275]));
    assign outputs[8619] = layer2_outputs[9419];
    assign outputs[8620] = (layer2_outputs[6106]) & ~(layer2_outputs[8146]);
    assign outputs[8621] = ~((layer2_outputs[4695]) ^ (layer2_outputs[10335]));
    assign outputs[8622] = ~(layer2_outputs[12647]);
    assign outputs[8623] = ~((layer2_outputs[6617]) | (layer2_outputs[6210]));
    assign outputs[8624] = (layer2_outputs[1113]) ^ (layer2_outputs[5975]);
    assign outputs[8625] = ~(layer2_outputs[1324]);
    assign outputs[8626] = ~(layer2_outputs[12619]) | (layer2_outputs[276]);
    assign outputs[8627] = ~(layer2_outputs[9232]);
    assign outputs[8628] = layer2_outputs[11376];
    assign outputs[8629] = ~(layer2_outputs[2773]);
    assign outputs[8630] = ~(layer2_outputs[6439]);
    assign outputs[8631] = layer2_outputs[3191];
    assign outputs[8632] = ~((layer2_outputs[4803]) ^ (layer2_outputs[4023]));
    assign outputs[8633] = layer2_outputs[12061];
    assign outputs[8634] = (layer2_outputs[6200]) & ~(layer2_outputs[8106]);
    assign outputs[8635] = ~(layer2_outputs[4351]);
    assign outputs[8636] = ~(layer2_outputs[3149]) | (layer2_outputs[10270]);
    assign outputs[8637] = ~((layer2_outputs[11796]) | (layer2_outputs[459]));
    assign outputs[8638] = layer2_outputs[2181];
    assign outputs[8639] = layer2_outputs[9729];
    assign outputs[8640] = ~(layer2_outputs[7748]);
    assign outputs[8641] = layer2_outputs[5650];
    assign outputs[8642] = ~(layer2_outputs[10570]);
    assign outputs[8643] = ~((layer2_outputs[10171]) & (layer2_outputs[2563]));
    assign outputs[8644] = ~((layer2_outputs[2399]) & (layer2_outputs[2538]));
    assign outputs[8645] = ~((layer2_outputs[4387]) ^ (layer2_outputs[12498]));
    assign outputs[8646] = layer2_outputs[4130];
    assign outputs[8647] = ~(layer2_outputs[2679]);
    assign outputs[8648] = (layer2_outputs[2069]) ^ (layer2_outputs[5718]);
    assign outputs[8649] = layer2_outputs[2483];
    assign outputs[8650] = ~(layer2_outputs[3139]);
    assign outputs[8651] = ~(layer2_outputs[8584]);
    assign outputs[8652] = layer2_outputs[3552];
    assign outputs[8653] = layer2_outputs[10015];
    assign outputs[8654] = ~(layer2_outputs[2471]);
    assign outputs[8655] = ~(layer2_outputs[8833]);
    assign outputs[8656] = ~(layer2_outputs[5106]);
    assign outputs[8657] = ~(layer2_outputs[11643]) | (layer2_outputs[2746]);
    assign outputs[8658] = layer2_outputs[3601];
    assign outputs[8659] = ~((layer2_outputs[12348]) ^ (layer2_outputs[99]));
    assign outputs[8660] = (layer2_outputs[11295]) ^ (layer2_outputs[10455]);
    assign outputs[8661] = ~(layer2_outputs[6684]);
    assign outputs[8662] = ~(layer2_outputs[3438]);
    assign outputs[8663] = layer2_outputs[5235];
    assign outputs[8664] = ~(layer2_outputs[1295]);
    assign outputs[8665] = ~(layer2_outputs[12589]);
    assign outputs[8666] = (layer2_outputs[10331]) & ~(layer2_outputs[9232]);
    assign outputs[8667] = ~(layer2_outputs[4849]);
    assign outputs[8668] = layer2_outputs[3499];
    assign outputs[8669] = ~(layer2_outputs[5694]) | (layer2_outputs[11753]);
    assign outputs[8670] = (layer2_outputs[12786]) | (layer2_outputs[12387]);
    assign outputs[8671] = layer2_outputs[9771];
    assign outputs[8672] = layer2_outputs[6052];
    assign outputs[8673] = ~((layer2_outputs[10532]) ^ (layer2_outputs[8514]));
    assign outputs[8674] = layer2_outputs[8250];
    assign outputs[8675] = ~(layer2_outputs[8523]);
    assign outputs[8676] = ~(layer2_outputs[8816]);
    assign outputs[8677] = ~((layer2_outputs[3778]) ^ (layer2_outputs[10758]));
    assign outputs[8678] = (layer2_outputs[1147]) ^ (layer2_outputs[8110]);
    assign outputs[8679] = (layer2_outputs[10735]) & ~(layer2_outputs[1588]);
    assign outputs[8680] = ~(layer2_outputs[2590]);
    assign outputs[8681] = layer2_outputs[4815];
    assign outputs[8682] = ~(layer2_outputs[8437]);
    assign outputs[8683] = layer2_outputs[2575];
    assign outputs[8684] = layer2_outputs[4971];
    assign outputs[8685] = layer2_outputs[3948];
    assign outputs[8686] = ~((layer2_outputs[4778]) ^ (layer2_outputs[1879]));
    assign outputs[8687] = ~(layer2_outputs[10236]);
    assign outputs[8688] = ~(layer2_outputs[9769]);
    assign outputs[8689] = (layer2_outputs[12104]) ^ (layer2_outputs[12073]);
    assign outputs[8690] = (layer2_outputs[632]) & (layer2_outputs[5354]);
    assign outputs[8691] = ~(layer2_outputs[4301]);
    assign outputs[8692] = (layer2_outputs[3026]) & ~(layer2_outputs[12188]);
    assign outputs[8693] = ~((layer2_outputs[5901]) | (layer2_outputs[1122]));
    assign outputs[8694] = layer2_outputs[2981];
    assign outputs[8695] = layer2_outputs[9281];
    assign outputs[8696] = layer2_outputs[527];
    assign outputs[8697] = ~(layer2_outputs[8508]);
    assign outputs[8698] = ~((layer2_outputs[1228]) ^ (layer2_outputs[7427]));
    assign outputs[8699] = ~(layer2_outputs[12311]);
    assign outputs[8700] = (layer2_outputs[12652]) & (layer2_outputs[10550]);
    assign outputs[8701] = layer2_outputs[10527];
    assign outputs[8702] = ~((layer2_outputs[9744]) | (layer2_outputs[8489]));
    assign outputs[8703] = (layer2_outputs[3765]) & ~(layer2_outputs[8844]);
    assign outputs[8704] = ~(layer2_outputs[2459]);
    assign outputs[8705] = ~(layer2_outputs[1912]);
    assign outputs[8706] = layer2_outputs[8064];
    assign outputs[8707] = layer2_outputs[7240];
    assign outputs[8708] = layer2_outputs[7798];
    assign outputs[8709] = ~(layer2_outputs[8398]) | (layer2_outputs[10938]);
    assign outputs[8710] = layer2_outputs[6653];
    assign outputs[8711] = ~(layer2_outputs[12455]);
    assign outputs[8712] = (layer2_outputs[863]) & (layer2_outputs[6696]);
    assign outputs[8713] = layer2_outputs[8917];
    assign outputs[8714] = layer2_outputs[4974];
    assign outputs[8715] = ~((layer2_outputs[7636]) | (layer2_outputs[6238]));
    assign outputs[8716] = (layer2_outputs[1377]) ^ (layer2_outputs[3024]);
    assign outputs[8717] = (layer2_outputs[2031]) & ~(layer2_outputs[4398]);
    assign outputs[8718] = layer2_outputs[6994];
    assign outputs[8719] = ~((layer2_outputs[1246]) ^ (layer2_outputs[1969]));
    assign outputs[8720] = layer2_outputs[3097];
    assign outputs[8721] = layer2_outputs[12173];
    assign outputs[8722] = ~(layer2_outputs[841]);
    assign outputs[8723] = layer2_outputs[10741];
    assign outputs[8724] = ~(layer2_outputs[7825]);
    assign outputs[8725] = ~(layer2_outputs[1821]);
    assign outputs[8726] = (layer2_outputs[8540]) ^ (layer2_outputs[3193]);
    assign outputs[8727] = ~((layer2_outputs[464]) ^ (layer2_outputs[12191]));
    assign outputs[8728] = (layer2_outputs[8914]) & (layer2_outputs[2435]);
    assign outputs[8729] = layer2_outputs[12787];
    assign outputs[8730] = ~(layer2_outputs[6924]);
    assign outputs[8731] = layer2_outputs[4159];
    assign outputs[8732] = layer2_outputs[5518];
    assign outputs[8733] = layer2_outputs[4685];
    assign outputs[8734] = ~(layer2_outputs[2230]);
    assign outputs[8735] = ~(layer2_outputs[2249]);
    assign outputs[8736] = ~(layer2_outputs[6502]);
    assign outputs[8737] = layer2_outputs[5474];
    assign outputs[8738] = layer2_outputs[3457];
    assign outputs[8739] = (layer2_outputs[8800]) ^ (layer2_outputs[1150]);
    assign outputs[8740] = (layer2_outputs[8395]) & ~(layer2_outputs[1647]);
    assign outputs[8741] = (layer2_outputs[9279]) & ~(layer2_outputs[6971]);
    assign outputs[8742] = (layer2_outputs[8092]) | (layer2_outputs[8579]);
    assign outputs[8743] = layer2_outputs[693];
    assign outputs[8744] = ~(layer2_outputs[3711]);
    assign outputs[8745] = layer2_outputs[6040];
    assign outputs[8746] = layer2_outputs[1065];
    assign outputs[8747] = layer2_outputs[10075];
    assign outputs[8748] = (layer2_outputs[12058]) & (layer2_outputs[12071]);
    assign outputs[8749] = ~(layer2_outputs[4453]);
    assign outputs[8750] = (layer2_outputs[11738]) | (layer2_outputs[3680]);
    assign outputs[8751] = ~(layer2_outputs[5266]);
    assign outputs[8752] = ~((layer2_outputs[3201]) | (layer2_outputs[7055]));
    assign outputs[8753] = ~((layer2_outputs[2606]) ^ (layer2_outputs[6472]));
    assign outputs[8754] = ~((layer2_outputs[2893]) ^ (layer2_outputs[7192]));
    assign outputs[8755] = (layer2_outputs[1369]) & ~(layer2_outputs[9623]);
    assign outputs[8756] = ~(layer2_outputs[2808]);
    assign outputs[8757] = ~(layer2_outputs[1503]);
    assign outputs[8758] = (layer2_outputs[90]) ^ (layer2_outputs[11544]);
    assign outputs[8759] = ~(layer2_outputs[239]);
    assign outputs[8760] = layer2_outputs[7753];
    assign outputs[8761] = layer2_outputs[7522];
    assign outputs[8762] = ~(layer2_outputs[3923]) | (layer2_outputs[4804]);
    assign outputs[8763] = ~((layer2_outputs[2883]) ^ (layer2_outputs[9453]));
    assign outputs[8764] = layer2_outputs[4952];
    assign outputs[8765] = ~(layer2_outputs[12217]);
    assign outputs[8766] = ~((layer2_outputs[11832]) ^ (layer2_outputs[7138]));
    assign outputs[8767] = ~(layer2_outputs[216]);
    assign outputs[8768] = ~(layer2_outputs[9711]);
    assign outputs[8769] = (layer2_outputs[4989]) & ~(layer2_outputs[9881]);
    assign outputs[8770] = ~(layer2_outputs[8684]);
    assign outputs[8771] = layer2_outputs[944];
    assign outputs[8772] = ~((layer2_outputs[1123]) ^ (layer2_outputs[12147]));
    assign outputs[8773] = layer2_outputs[9997];
    assign outputs[8774] = layer2_outputs[11799];
    assign outputs[8775] = ~((layer2_outputs[6571]) ^ (layer2_outputs[6813]));
    assign outputs[8776] = (layer2_outputs[520]) ^ (layer2_outputs[12250]);
    assign outputs[8777] = layer2_outputs[4887];
    assign outputs[8778] = ~(layer2_outputs[5765]);
    assign outputs[8779] = (layer2_outputs[5290]) & ~(layer2_outputs[8408]);
    assign outputs[8780] = (layer2_outputs[11283]) ^ (layer2_outputs[9267]);
    assign outputs[8781] = (layer2_outputs[1596]) ^ (layer2_outputs[4837]);
    assign outputs[8782] = ~(layer2_outputs[11971]);
    assign outputs[8783] = ~(layer2_outputs[3301]);
    assign outputs[8784] = ~(layer2_outputs[324]);
    assign outputs[8785] = (layer2_outputs[3926]) ^ (layer2_outputs[10433]);
    assign outputs[8786] = ~(layer2_outputs[10836]);
    assign outputs[8787] = layer2_outputs[12002];
    assign outputs[8788] = ~((layer2_outputs[11933]) ^ (layer2_outputs[12645]));
    assign outputs[8789] = (layer2_outputs[7031]) ^ (layer2_outputs[7140]);
    assign outputs[8790] = ~((layer2_outputs[12195]) | (layer2_outputs[10011]));
    assign outputs[8791] = layer2_outputs[7303];
    assign outputs[8792] = ~(layer2_outputs[6489]);
    assign outputs[8793] = ~((layer2_outputs[1860]) ^ (layer2_outputs[2191]));
    assign outputs[8794] = layer2_outputs[9648];
    assign outputs[8795] = (layer2_outputs[7012]) ^ (layer2_outputs[9757]);
    assign outputs[8796] = ~((layer2_outputs[2230]) ^ (layer2_outputs[9787]));
    assign outputs[8797] = (layer2_outputs[7827]) & ~(layer2_outputs[592]);
    assign outputs[8798] = ~(layer2_outputs[7956]);
    assign outputs[8799] = layer2_outputs[12505];
    assign outputs[8800] = (layer2_outputs[7356]) ^ (layer2_outputs[2974]);
    assign outputs[8801] = layer2_outputs[9124];
    assign outputs[8802] = ~(layer2_outputs[4904]) | (layer2_outputs[371]);
    assign outputs[8803] = ~((layer2_outputs[9493]) ^ (layer2_outputs[2194]));
    assign outputs[8804] = ~((layer2_outputs[12306]) ^ (layer2_outputs[12384]));
    assign outputs[8805] = ~((layer2_outputs[12232]) ^ (layer2_outputs[9147]));
    assign outputs[8806] = layer2_outputs[12101];
    assign outputs[8807] = layer2_outputs[5402];
    assign outputs[8808] = ~(layer2_outputs[383]);
    assign outputs[8809] = ~(layer2_outputs[8334]);
    assign outputs[8810] = layer2_outputs[6187];
    assign outputs[8811] = (layer2_outputs[10980]) & ~(layer2_outputs[7591]);
    assign outputs[8812] = ~(layer2_outputs[3556]);
    assign outputs[8813] = layer2_outputs[6162];
    assign outputs[8814] = ~(layer2_outputs[7351]);
    assign outputs[8815] = layer2_outputs[1792];
    assign outputs[8816] = layer2_outputs[2888];
    assign outputs[8817] = (layer2_outputs[2830]) & (layer2_outputs[4991]);
    assign outputs[8818] = ~(layer2_outputs[12460]);
    assign outputs[8819] = (layer2_outputs[8847]) ^ (layer2_outputs[6540]);
    assign outputs[8820] = ~(layer2_outputs[5540]);
    assign outputs[8821] = layer2_outputs[7905];
    assign outputs[8822] = (layer2_outputs[12408]) ^ (layer2_outputs[10791]);
    assign outputs[8823] = ~(layer2_outputs[3550]);
    assign outputs[8824] = ~(layer2_outputs[11084]);
    assign outputs[8825] = layer2_outputs[645];
    assign outputs[8826] = ~(layer2_outputs[4493]);
    assign outputs[8827] = layer2_outputs[690];
    assign outputs[8828] = layer2_outputs[1641];
    assign outputs[8829] = ~(layer2_outputs[7163]);
    assign outputs[8830] = ~(layer2_outputs[678]);
    assign outputs[8831] = ~((layer2_outputs[2424]) ^ (layer2_outputs[10881]));
    assign outputs[8832] = (layer2_outputs[6156]) & ~(layer2_outputs[773]);
    assign outputs[8833] = ~(layer2_outputs[6975]);
    assign outputs[8834] = ~(layer2_outputs[9424]);
    assign outputs[8835] = layer2_outputs[5165];
    assign outputs[8836] = ~(layer2_outputs[8877]);
    assign outputs[8837] = layer2_outputs[3386];
    assign outputs[8838] = ~(layer2_outputs[2942]);
    assign outputs[8839] = (layer2_outputs[6874]) & (layer2_outputs[3758]);
    assign outputs[8840] = ~((layer2_outputs[2061]) | (layer2_outputs[8966]));
    assign outputs[8841] = layer2_outputs[4148];
    assign outputs[8842] = layer2_outputs[11720];
    assign outputs[8843] = (layer2_outputs[8613]) ^ (layer2_outputs[830]);
    assign outputs[8844] = ~(layer2_outputs[7296]) | (layer2_outputs[11657]);
    assign outputs[8845] = ~(layer2_outputs[9141]) | (layer2_outputs[3086]);
    assign outputs[8846] = ~((layer2_outputs[4603]) ^ (layer2_outputs[8518]));
    assign outputs[8847] = layer2_outputs[6712];
    assign outputs[8848] = layer2_outputs[1467];
    assign outputs[8849] = ~((layer2_outputs[7428]) ^ (layer2_outputs[2567]));
    assign outputs[8850] = ~(layer2_outputs[11962]);
    assign outputs[8851] = layer2_outputs[4883];
    assign outputs[8852] = (layer2_outputs[5641]) ^ (layer2_outputs[3868]);
    assign outputs[8853] = layer2_outputs[11317];
    assign outputs[8854] = ~(layer2_outputs[7253]) | (layer2_outputs[4212]);
    assign outputs[8855] = ~(layer2_outputs[731]);
    assign outputs[8856] = layer2_outputs[11742];
    assign outputs[8857] = (layer2_outputs[3766]) ^ (layer2_outputs[4995]);
    assign outputs[8858] = ~((layer2_outputs[11329]) ^ (layer2_outputs[2736]));
    assign outputs[8859] = ~((layer2_outputs[6829]) | (layer2_outputs[809]));
    assign outputs[8860] = (layer2_outputs[7433]) ^ (layer2_outputs[7444]);
    assign outputs[8861] = ~(layer2_outputs[12032]);
    assign outputs[8862] = layer2_outputs[6595];
    assign outputs[8863] = layer2_outputs[2381];
    assign outputs[8864] = (layer2_outputs[12617]) ^ (layer2_outputs[10647]);
    assign outputs[8865] = ~((layer2_outputs[825]) ^ (layer2_outputs[2955]));
    assign outputs[8866] = layer2_outputs[5612];
    assign outputs[8867] = (layer2_outputs[6049]) ^ (layer2_outputs[11426]);
    assign outputs[8868] = layer2_outputs[10296];
    assign outputs[8869] = ~(layer2_outputs[1455]);
    assign outputs[8870] = layer2_outputs[6488];
    assign outputs[8871] = ~(layer2_outputs[12447]);
    assign outputs[8872] = ~(layer2_outputs[7481]);
    assign outputs[8873] = ~((layer2_outputs[3759]) ^ (layer2_outputs[2765]));
    assign outputs[8874] = ~((layer2_outputs[4361]) ^ (layer2_outputs[5702]));
    assign outputs[8875] = ~(layer2_outputs[10148]);
    assign outputs[8876] = layer2_outputs[8373];
    assign outputs[8877] = layer2_outputs[4653];
    assign outputs[8878] = (layer2_outputs[3636]) & ~(layer2_outputs[11246]);
    assign outputs[8879] = layer2_outputs[292];
    assign outputs[8880] = ~(layer2_outputs[546]);
    assign outputs[8881] = ~(layer2_outputs[5999]);
    assign outputs[8882] = layer2_outputs[11470];
    assign outputs[8883] = layer2_outputs[6040];
    assign outputs[8884] = layer2_outputs[8030];
    assign outputs[8885] = layer2_outputs[9185];
    assign outputs[8886] = layer2_outputs[9972];
    assign outputs[8887] = ~((layer2_outputs[2390]) ^ (layer2_outputs[8498]));
    assign outputs[8888] = (layer2_outputs[8101]) & (layer2_outputs[7699]);
    assign outputs[8889] = (layer2_outputs[2530]) ^ (layer2_outputs[3704]);
    assign outputs[8890] = ~(layer2_outputs[7210]);
    assign outputs[8891] = ~(layer2_outputs[11998]);
    assign outputs[8892] = layer2_outputs[6676];
    assign outputs[8893] = ~(layer2_outputs[11655]);
    assign outputs[8894] = layer2_outputs[7300];
    assign outputs[8895] = ~((layer2_outputs[12511]) | (layer2_outputs[115]));
    assign outputs[8896] = (layer2_outputs[9528]) & (layer2_outputs[5851]);
    assign outputs[8897] = ~(layer2_outputs[616]);
    assign outputs[8898] = ~(layer2_outputs[7996]);
    assign outputs[8899] = ~(layer2_outputs[7448]);
    assign outputs[8900] = (layer2_outputs[8512]) & ~(layer2_outputs[6390]);
    assign outputs[8901] = ~(layer2_outputs[3808]);
    assign outputs[8902] = (layer2_outputs[7415]) ^ (layer2_outputs[8104]);
    assign outputs[8903] = (layer2_outputs[6980]) ^ (layer2_outputs[5407]);
    assign outputs[8904] = layer2_outputs[5847];
    assign outputs[8905] = (layer2_outputs[2550]) & ~(layer2_outputs[3735]);
    assign outputs[8906] = ~(layer2_outputs[6828]) | (layer2_outputs[6463]);
    assign outputs[8907] = ~((layer2_outputs[12278]) ^ (layer2_outputs[6520]));
    assign outputs[8908] = (layer2_outputs[10777]) | (layer2_outputs[3594]);
    assign outputs[8909] = ~(layer2_outputs[4460]) | (layer2_outputs[8032]);
    assign outputs[8910] = ~(layer2_outputs[111]);
    assign outputs[8911] = ~(layer2_outputs[12457]);
    assign outputs[8912] = ~(layer2_outputs[10375]);
    assign outputs[8913] = ~((layer2_outputs[2222]) | (layer2_outputs[120]));
    assign outputs[8914] = layer2_outputs[9704];
    assign outputs[8915] = ~((layer2_outputs[5153]) ^ (layer2_outputs[3929]));
    assign outputs[8916] = ~(layer2_outputs[3850]);
    assign outputs[8917] = (layer2_outputs[278]) & ~(layer2_outputs[554]);
    assign outputs[8918] = ~(layer2_outputs[6477]);
    assign outputs[8919] = ~(layer2_outputs[12100]);
    assign outputs[8920] = ~((layer2_outputs[10282]) ^ (layer2_outputs[207]));
    assign outputs[8921] = layer2_outputs[4241];
    assign outputs[8922] = ~(layer2_outputs[12042]);
    assign outputs[8923] = ~(layer2_outputs[2642]);
    assign outputs[8924] = ~(layer2_outputs[5124]);
    assign outputs[8925] = ~(layer2_outputs[7277]) | (layer2_outputs[434]);
    assign outputs[8926] = (layer2_outputs[11231]) ^ (layer2_outputs[7840]);
    assign outputs[8927] = ~(layer2_outputs[11263]);
    assign outputs[8928] = ~(layer2_outputs[3103]);
    assign outputs[8929] = layer2_outputs[10842];
    assign outputs[8930] = ~((layer2_outputs[6442]) ^ (layer2_outputs[1909]));
    assign outputs[8931] = ~(layer2_outputs[9507]);
    assign outputs[8932] = ~(layer2_outputs[5384]);
    assign outputs[8933] = ~(layer2_outputs[3303]);
    assign outputs[8934] = ~(layer2_outputs[1997]);
    assign outputs[8935] = ~((layer2_outputs[6122]) | (layer2_outputs[1787]));
    assign outputs[8936] = layer2_outputs[1957];
    assign outputs[8937] = ~(layer2_outputs[7456]);
    assign outputs[8938] = ~(layer2_outputs[6403]);
    assign outputs[8939] = layer2_outputs[8784];
    assign outputs[8940] = ~(layer2_outputs[2011]);
    assign outputs[8941] = ~(layer2_outputs[2761]);
    assign outputs[8942] = (layer2_outputs[6033]) ^ (layer2_outputs[5738]);
    assign outputs[8943] = (layer2_outputs[6536]) & ~(layer2_outputs[2421]);
    assign outputs[8944] = ~((layer2_outputs[4888]) | (layer2_outputs[9487]));
    assign outputs[8945] = ~(layer2_outputs[8146]);
    assign outputs[8946] = (layer2_outputs[8764]) & ~(layer2_outputs[10640]);
    assign outputs[8947] = ~(layer2_outputs[4166]);
    assign outputs[8948] = (layer2_outputs[339]) & ~(layer2_outputs[3279]);
    assign outputs[8949] = ~(layer2_outputs[6500]);
    assign outputs[8950] = ~((layer2_outputs[3526]) | (layer2_outputs[8865]));
    assign outputs[8951] = layer2_outputs[6142];
    assign outputs[8952] = ~(layer2_outputs[10780]);
    assign outputs[8953] = ~((layer2_outputs[8260]) ^ (layer2_outputs[7467]));
    assign outputs[8954] = layer2_outputs[8347];
    assign outputs[8955] = ~(layer2_outputs[7032]);
    assign outputs[8956] = (layer2_outputs[11287]) & (layer2_outputs[2982]);
    assign outputs[8957] = layer2_outputs[1946];
    assign outputs[8958] = (layer2_outputs[10364]) | (layer2_outputs[3558]);
    assign outputs[8959] = ~(layer2_outputs[12703]);
    assign outputs[8960] = (layer2_outputs[3520]) ^ (layer2_outputs[3371]);
    assign outputs[8961] = layer2_outputs[508];
    assign outputs[8962] = layer2_outputs[9060];
    assign outputs[8963] = layer2_outputs[7765];
    assign outputs[8964] = (layer2_outputs[11523]) ^ (layer2_outputs[10825]);
    assign outputs[8965] = ~(layer2_outputs[11486]) | (layer2_outputs[6335]);
    assign outputs[8966] = ~(layer2_outputs[697]);
    assign outputs[8967] = ~((layer2_outputs[1140]) ^ (layer2_outputs[7358]));
    assign outputs[8968] = (layer2_outputs[12757]) & ~(layer2_outputs[9621]);
    assign outputs[8969] = (layer2_outputs[11354]) & ~(layer2_outputs[11802]);
    assign outputs[8970] = ~(layer2_outputs[1940]);
    assign outputs[8971] = ~((layer2_outputs[7649]) ^ (layer2_outputs[1538]));
    assign outputs[8972] = (layer2_outputs[11684]) ^ (layer2_outputs[3963]);
    assign outputs[8973] = (layer2_outputs[8537]) ^ (layer2_outputs[10246]);
    assign outputs[8974] = layer2_outputs[965];
    assign outputs[8975] = ~((layer2_outputs[198]) & (layer2_outputs[3939]));
    assign outputs[8976] = (layer2_outputs[3083]) ^ (layer2_outputs[8680]);
    assign outputs[8977] = layer2_outputs[8888];
    assign outputs[8978] = layer2_outputs[7299];
    assign outputs[8979] = (layer2_outputs[11595]) & ~(layer2_outputs[7984]);
    assign outputs[8980] = ~(layer2_outputs[5869]);
    assign outputs[8981] = (layer2_outputs[3048]) ^ (layer2_outputs[11115]);
    assign outputs[8982] = layer2_outputs[9118];
    assign outputs[8983] = (layer2_outputs[2315]) & ~(layer2_outputs[2497]);
    assign outputs[8984] = layer2_outputs[2198];
    assign outputs[8985] = layer2_outputs[11991];
    assign outputs[8986] = ~(layer2_outputs[3587]);
    assign outputs[8987] = (layer2_outputs[8793]) & ~(layer2_outputs[10157]);
    assign outputs[8988] = (layer2_outputs[5552]) ^ (layer2_outputs[5786]);
    assign outputs[8989] = layer2_outputs[12020];
    assign outputs[8990] = ~(layer2_outputs[8339]);
    assign outputs[8991] = ~(layer2_outputs[9498]) | (layer2_outputs[5127]);
    assign outputs[8992] = (layer2_outputs[474]) | (layer2_outputs[1372]);
    assign outputs[8993] = (layer2_outputs[3650]) ^ (layer2_outputs[12218]);
    assign outputs[8994] = ~(layer2_outputs[1716]);
    assign outputs[8995] = layer2_outputs[9344];
    assign outputs[8996] = ~(layer2_outputs[4296]);
    assign outputs[8997] = (layer2_outputs[6745]) & (layer2_outputs[925]);
    assign outputs[8998] = ~((layer2_outputs[9155]) ^ (layer2_outputs[2069]));
    assign outputs[8999] = layer2_outputs[9442];
    assign outputs[9000] = ~(layer2_outputs[6253]) | (layer2_outputs[1386]);
    assign outputs[9001] = ~((layer2_outputs[6233]) ^ (layer2_outputs[9383]));
    assign outputs[9002] = ~(layer2_outputs[8912]);
    assign outputs[9003] = layer2_outputs[3399];
    assign outputs[9004] = ~((layer2_outputs[5762]) | (layer2_outputs[10726]));
    assign outputs[9005] = layer2_outputs[10975];
    assign outputs[9006] = ~(layer2_outputs[801]);
    assign outputs[9007] = ~((layer2_outputs[10218]) ^ (layer2_outputs[8615]));
    assign outputs[9008] = layer2_outputs[8577];
    assign outputs[9009] = (layer2_outputs[6847]) ^ (layer2_outputs[1562]);
    assign outputs[9010] = (layer2_outputs[4546]) & ~(layer2_outputs[5883]);
    assign outputs[9011] = ~(layer2_outputs[3959]);
    assign outputs[9012] = layer2_outputs[10882];
    assign outputs[9013] = layer2_outputs[3806];
    assign outputs[9014] = ~((layer2_outputs[2244]) & (layer2_outputs[2933]));
    assign outputs[9015] = (layer2_outputs[12013]) & ~(layer2_outputs[11619]);
    assign outputs[9016] = layer2_outputs[9255];
    assign outputs[9017] = ~(layer2_outputs[1519]);
    assign outputs[9018] = (layer2_outputs[11202]) & ~(layer2_outputs[1601]);
    assign outputs[9019] = ~(layer2_outputs[10031]);
    assign outputs[9020] = (layer2_outputs[6982]) & ~(layer2_outputs[4102]);
    assign outputs[9021] = (layer2_outputs[1313]) & ~(layer2_outputs[5398]);
    assign outputs[9022] = ~(layer2_outputs[10083]);
    assign outputs[9023] = layer2_outputs[3495];
    assign outputs[9024] = layer2_outputs[7766];
    assign outputs[9025] = ~(layer2_outputs[10611]);
    assign outputs[9026] = ~(layer2_outputs[12276]);
    assign outputs[9027] = ~(layer2_outputs[1571]);
    assign outputs[9028] = ~(layer2_outputs[8976]);
    assign outputs[9029] = ~(layer2_outputs[3691]);
    assign outputs[9030] = ~((layer2_outputs[2594]) | (layer2_outputs[9209]));
    assign outputs[9031] = ~(layer2_outputs[8780]);
    assign outputs[9032] = ~((layer2_outputs[1115]) ^ (layer2_outputs[2460]));
    assign outputs[9033] = layer2_outputs[7797];
    assign outputs[9034] = ~(layer2_outputs[7245]);
    assign outputs[9035] = ~(layer2_outputs[6093]);
    assign outputs[9036] = ~(layer2_outputs[9796]);
    assign outputs[9037] = (layer2_outputs[1627]) ^ (layer2_outputs[10286]);
    assign outputs[9038] = ~(layer2_outputs[6496]);
    assign outputs[9039] = (layer2_outputs[9066]) | (layer2_outputs[1603]);
    assign outputs[9040] = ~((layer2_outputs[8367]) ^ (layer2_outputs[12527]));
    assign outputs[9041] = ~((layer2_outputs[6290]) ^ (layer2_outputs[4465]));
    assign outputs[9042] = layer2_outputs[2687];
    assign outputs[9043] = ~(layer2_outputs[3117]);
    assign outputs[9044] = ~(layer2_outputs[12169]);
    assign outputs[9045] = ~(layer2_outputs[9818]) | (layer2_outputs[2140]);
    assign outputs[9046] = (layer2_outputs[6083]) & (layer2_outputs[9106]);
    assign outputs[9047] = layer2_outputs[3974];
    assign outputs[9048] = (layer2_outputs[5523]) ^ (layer2_outputs[2884]);
    assign outputs[9049] = (layer2_outputs[9970]) ^ (layer2_outputs[553]);
    assign outputs[9050] = ~(layer2_outputs[6783]);
    assign outputs[9051] = ~(layer2_outputs[11509]);
    assign outputs[9052] = ~(layer2_outputs[4535]);
    assign outputs[9053] = ~(layer2_outputs[9032]);
    assign outputs[9054] = ~(layer2_outputs[2501]);
    assign outputs[9055] = layer2_outputs[8657];
    assign outputs[9056] = (layer2_outputs[5891]) ^ (layer2_outputs[6732]);
    assign outputs[9057] = (layer2_outputs[1223]) & ~(layer2_outputs[6633]);
    assign outputs[9058] = ~(layer2_outputs[1359]);
    assign outputs[9059] = ~((layer2_outputs[2476]) ^ (layer2_outputs[1535]));
    assign outputs[9060] = ~(layer2_outputs[4582]);
    assign outputs[9061] = ~(layer2_outputs[2722]);
    assign outputs[9062] = ~((layer2_outputs[4986]) ^ (layer2_outputs[6618]));
    assign outputs[9063] = ~(layer2_outputs[8200]);
    assign outputs[9064] = ~((layer2_outputs[7245]) ^ (layer2_outputs[12261]));
    assign outputs[9065] = (layer2_outputs[12777]) ^ (layer2_outputs[5472]);
    assign outputs[9066] = layer2_outputs[8327];
    assign outputs[9067] = ~(layer2_outputs[10101]);
    assign outputs[9068] = (layer2_outputs[4988]) & ~(layer2_outputs[10341]);
    assign outputs[9069] = ~((layer2_outputs[7005]) ^ (layer2_outputs[11340]));
    assign outputs[9070] = layer2_outputs[9694];
    assign outputs[9071] = layer2_outputs[1978];
    assign outputs[9072] = layer2_outputs[8451];
    assign outputs[9073] = ~((layer2_outputs[7054]) & (layer2_outputs[209]));
    assign outputs[9074] = layer2_outputs[6787];
    assign outputs[9075] = (layer2_outputs[9386]) & ~(layer2_outputs[5337]);
    assign outputs[9076] = ~(layer2_outputs[6573]);
    assign outputs[9077] = layer2_outputs[3312];
    assign outputs[9078] = ~((layer2_outputs[10663]) | (layer2_outputs[3490]));
    assign outputs[9079] = layer2_outputs[986];
    assign outputs[9080] = ~(layer2_outputs[10559]) | (layer2_outputs[8563]);
    assign outputs[9081] = (layer2_outputs[4040]) ^ (layer2_outputs[6991]);
    assign outputs[9082] = (layer2_outputs[7723]) & ~(layer2_outputs[5286]);
    assign outputs[9083] = layer2_outputs[1033];
    assign outputs[9084] = ~(layer2_outputs[1013]);
    assign outputs[9085] = ~(layer2_outputs[11907]);
    assign outputs[9086] = ~(layer2_outputs[478]);
    assign outputs[9087] = ~(layer2_outputs[9402]);
    assign outputs[9088] = (layer2_outputs[9019]) ^ (layer2_outputs[91]);
    assign outputs[9089] = ~(layer2_outputs[10533]);
    assign outputs[9090] = layer2_outputs[2637];
    assign outputs[9091] = (layer2_outputs[10372]) & ~(layer2_outputs[7733]);
    assign outputs[9092] = ~(layer2_outputs[3319]);
    assign outputs[9093] = layer2_outputs[10375];
    assign outputs[9094] = ~(layer2_outputs[12309]);
    assign outputs[9095] = ~(layer2_outputs[12762]) | (layer2_outputs[11097]);
    assign outputs[9096] = ~(layer2_outputs[1259]);
    assign outputs[9097] = layer2_outputs[9904];
    assign outputs[9098] = ~(layer2_outputs[1218]);
    assign outputs[9099] = ~(layer2_outputs[11044]);
    assign outputs[9100] = layer2_outputs[7410];
    assign outputs[9101] = ~(layer2_outputs[3328]);
    assign outputs[9102] = ~(layer2_outputs[5582]);
    assign outputs[9103] = ~(layer2_outputs[12247]);
    assign outputs[9104] = ~(layer2_outputs[2992]);
    assign outputs[9105] = layer2_outputs[2875];
    assign outputs[9106] = (layer2_outputs[813]) & ~(layer2_outputs[314]);
    assign outputs[9107] = (layer2_outputs[1748]) & ~(layer2_outputs[6685]);
    assign outputs[9108] = ~((layer2_outputs[7293]) ^ (layer2_outputs[4811]));
    assign outputs[9109] = layer2_outputs[6934];
    assign outputs[9110] = ~(layer2_outputs[10020]);
    assign outputs[9111] = layer2_outputs[1927];
    assign outputs[9112] = (layer2_outputs[5432]) ^ (layer2_outputs[8560]);
    assign outputs[9113] = ~(layer2_outputs[262]);
    assign outputs[9114] = (layer2_outputs[5560]) ^ (layer2_outputs[8019]);
    assign outputs[9115] = ~((layer2_outputs[12107]) | (layer2_outputs[6983]));
    assign outputs[9116] = (layer2_outputs[7309]) | (layer2_outputs[2408]);
    assign outputs[9117] = ~(layer2_outputs[1431]);
    assign outputs[9118] = layer2_outputs[7797];
    assign outputs[9119] = (layer2_outputs[4105]) | (layer2_outputs[3831]);
    assign outputs[9120] = ~(layer2_outputs[10128]);
    assign outputs[9121] = (layer2_outputs[8765]) & (layer2_outputs[6445]);
    assign outputs[9122] = ~((layer2_outputs[4436]) | (layer2_outputs[307]));
    assign outputs[9123] = layer2_outputs[11222];
    assign outputs[9124] = ~(layer2_outputs[3171]);
    assign outputs[9125] = ~((layer2_outputs[4458]) ^ (layer2_outputs[11452]));
    assign outputs[9126] = ~((layer2_outputs[5415]) ^ (layer2_outputs[7879]));
    assign outputs[9127] = layer2_outputs[10442];
    assign outputs[9128] = (layer2_outputs[12540]) ^ (layer2_outputs[11217]);
    assign outputs[9129] = ~((layer2_outputs[3059]) ^ (layer2_outputs[5298]));
    assign outputs[9130] = ~(layer2_outputs[891]);
    assign outputs[9131] = ~((layer2_outputs[4202]) ^ (layer2_outputs[11454]));
    assign outputs[9132] = layer2_outputs[4658];
    assign outputs[9133] = layer2_outputs[6259];
    assign outputs[9134] = ~((layer2_outputs[7694]) ^ (layer2_outputs[7995]));
    assign outputs[9135] = ~(layer2_outputs[2002]);
    assign outputs[9136] = ~(layer2_outputs[7026]);
    assign outputs[9137] = (layer2_outputs[2667]) ^ (layer2_outputs[7750]);
    assign outputs[9138] = ~(layer2_outputs[4992]);
    assign outputs[9139] = ~(layer2_outputs[4383]);
    assign outputs[9140] = ~((layer2_outputs[8814]) ^ (layer2_outputs[11393]));
    assign outputs[9141] = ~((layer2_outputs[12267]) ^ (layer2_outputs[1186]));
    assign outputs[9142] = ~(layer2_outputs[9293]);
    assign outputs[9143] = layer2_outputs[6284];
    assign outputs[9144] = ~((layer2_outputs[8475]) ^ (layer2_outputs[4557]));
    assign outputs[9145] = ~(layer2_outputs[5343]);
    assign outputs[9146] = ~(layer2_outputs[5075]);
    assign outputs[9147] = layer2_outputs[8111];
    assign outputs[9148] = layer2_outputs[4465];
    assign outputs[9149] = ~(layer2_outputs[5556]);
    assign outputs[9150] = ~(layer2_outputs[12271]) | (layer2_outputs[8186]);
    assign outputs[9151] = layer2_outputs[5670];
    assign outputs[9152] = (layer2_outputs[6781]) ^ (layer2_outputs[9055]);
    assign outputs[9153] = ~(layer2_outputs[12287]);
    assign outputs[9154] = ~((layer2_outputs[9176]) ^ (layer2_outputs[10104]));
    assign outputs[9155] = ~(layer2_outputs[8488]);
    assign outputs[9156] = layer2_outputs[12323];
    assign outputs[9157] = (layer2_outputs[6235]) ^ (layer2_outputs[1672]);
    assign outputs[9158] = ~(layer2_outputs[10346]);
    assign outputs[9159] = ~(layer2_outputs[8397]);
    assign outputs[9160] = ~(layer2_outputs[10534]);
    assign outputs[9161] = ~(layer2_outputs[599]) | (layer2_outputs[5575]);
    assign outputs[9162] = ~(layer2_outputs[192]);
    assign outputs[9163] = (layer2_outputs[12689]) & (layer2_outputs[857]);
    assign outputs[9164] = ~(layer2_outputs[4026]) | (layer2_outputs[10355]);
    assign outputs[9165] = ~(layer2_outputs[5238]);
    assign outputs[9166] = ~((layer2_outputs[5346]) ^ (layer2_outputs[1099]));
    assign outputs[9167] = ~((layer2_outputs[3336]) ^ (layer2_outputs[5023]));
    assign outputs[9168] = layer2_outputs[10383];
    assign outputs[9169] = layer2_outputs[11111];
    assign outputs[9170] = ~(layer2_outputs[2570]);
    assign outputs[9171] = (layer2_outputs[5517]) ^ (layer2_outputs[11005]);
    assign outputs[9172] = ~(layer2_outputs[8701]);
    assign outputs[9173] = (layer2_outputs[3489]) & ~(layer2_outputs[9412]);
    assign outputs[9174] = ~(layer2_outputs[908]);
    assign outputs[9175] = ~(layer2_outputs[8794]);
    assign outputs[9176] = layer2_outputs[6435];
    assign outputs[9177] = layer2_outputs[296];
    assign outputs[9178] = ~(layer2_outputs[1402]);
    assign outputs[9179] = (layer2_outputs[12673]) ^ (layer2_outputs[10451]);
    assign outputs[9180] = (layer2_outputs[2859]) & (layer2_outputs[2473]);
    assign outputs[9181] = ~(layer2_outputs[11474]);
    assign outputs[9182] = ~(layer2_outputs[9793]);
    assign outputs[9183] = ~(layer2_outputs[11327]);
    assign outputs[9184] = ~((layer2_outputs[6715]) ^ (layer2_outputs[4822]));
    assign outputs[9185] = layer2_outputs[2847];
    assign outputs[9186] = ~((layer2_outputs[11624]) ^ (layer2_outputs[3909]));
    assign outputs[9187] = (layer2_outputs[8798]) & ~(layer2_outputs[946]);
    assign outputs[9188] = (layer2_outputs[9044]) ^ (layer2_outputs[3644]);
    assign outputs[9189] = layer2_outputs[3270];
    assign outputs[9190] = layer2_outputs[2118];
    assign outputs[9191] = (layer2_outputs[10504]) ^ (layer2_outputs[11795]);
    assign outputs[9192] = (layer2_outputs[4358]) & ~(layer2_outputs[5256]);
    assign outputs[9193] = layer2_outputs[1312];
    assign outputs[9194] = (layer2_outputs[12480]) & ~(layer2_outputs[306]);
    assign outputs[9195] = (layer2_outputs[7094]) & (layer2_outputs[4160]);
    assign outputs[9196] = ~(layer2_outputs[3814]);
    assign outputs[9197] = ~(layer2_outputs[1951]);
    assign outputs[9198] = layer2_outputs[1110];
    assign outputs[9199] = ~(layer2_outputs[8434]);
    assign outputs[9200] = (layer2_outputs[9943]) & ~(layer2_outputs[10449]);
    assign outputs[9201] = (layer2_outputs[1335]) & (layer2_outputs[6947]);
    assign outputs[9202] = ~((layer2_outputs[8319]) ^ (layer2_outputs[7969]));
    assign outputs[9203] = layer2_outputs[3375];
    assign outputs[9204] = (layer2_outputs[3218]) & ~(layer2_outputs[7988]);
    assign outputs[9205] = layer2_outputs[11269];
    assign outputs[9206] = ~(layer2_outputs[5022]);
    assign outputs[9207] = (layer2_outputs[8789]) & ~(layer2_outputs[8540]);
    assign outputs[9208] = layer2_outputs[12624];
    assign outputs[9209] = ~((layer2_outputs[11626]) ^ (layer2_outputs[504]));
    assign outputs[9210] = ~(layer2_outputs[4069]);
    assign outputs[9211] = ~(layer2_outputs[3953]);
    assign outputs[9212] = ~((layer2_outputs[1513]) | (layer2_outputs[9423]));
    assign outputs[9213] = layer2_outputs[230];
    assign outputs[9214] = layer2_outputs[1978];
    assign outputs[9215] = ~(layer2_outputs[2071]);
    assign outputs[9216] = (layer2_outputs[898]) | (layer2_outputs[4910]);
    assign outputs[9217] = layer2_outputs[12767];
    assign outputs[9218] = ~(layer2_outputs[3171]);
    assign outputs[9219] = (layer2_outputs[10242]) ^ (layer2_outputs[10125]);
    assign outputs[9220] = (layer2_outputs[5913]) ^ (layer2_outputs[2593]);
    assign outputs[9221] = (layer2_outputs[670]) | (layer2_outputs[10809]);
    assign outputs[9222] = layer2_outputs[9370];
    assign outputs[9223] = layer2_outputs[10709];
    assign outputs[9224] = ~(layer2_outputs[6584]);
    assign outputs[9225] = ~(layer2_outputs[6018]);
    assign outputs[9226] = ~((layer2_outputs[3206]) & (layer2_outputs[3302]));
    assign outputs[9227] = ~((layer2_outputs[6219]) ^ (layer2_outputs[12492]));
    assign outputs[9228] = (layer2_outputs[5784]) & ~(layer2_outputs[5800]);
    assign outputs[9229] = ~(layer2_outputs[8333]);
    assign outputs[9230] = layer2_outputs[1291];
    assign outputs[9231] = layer2_outputs[7055];
    assign outputs[9232] = ~((layer2_outputs[1246]) ^ (layer2_outputs[7896]));
    assign outputs[9233] = ~(layer2_outputs[865]);
    assign outputs[9234] = layer2_outputs[2757];
    assign outputs[9235] = ~(layer2_outputs[328]);
    assign outputs[9236] = ~(layer2_outputs[3305]);
    assign outputs[9237] = ~((layer2_outputs[11614]) | (layer2_outputs[10216]));
    assign outputs[9238] = ~(layer2_outputs[8116]) | (layer2_outputs[5368]);
    assign outputs[9239] = ~(layer2_outputs[1388]);
    assign outputs[9240] = ~(layer2_outputs[8210]) | (layer2_outputs[1397]);
    assign outputs[9241] = (layer2_outputs[2654]) | (layer2_outputs[106]);
    assign outputs[9242] = ~(layer2_outputs[9271]);
    assign outputs[9243] = ~((layer2_outputs[1598]) ^ (layer2_outputs[11162]));
    assign outputs[9244] = (layer2_outputs[2070]) & ~(layer2_outputs[7802]);
    assign outputs[9245] = ~(layer2_outputs[6939]);
    assign outputs[9246] = ~(layer2_outputs[12752]);
    assign outputs[9247] = ~(layer2_outputs[5317]) | (layer2_outputs[4134]);
    assign outputs[9248] = layer2_outputs[5277];
    assign outputs[9249] = layer2_outputs[9962];
    assign outputs[9250] = ~((layer2_outputs[8226]) | (layer2_outputs[11045]));
    assign outputs[9251] = layer2_outputs[7535];
    assign outputs[9252] = ~(layer2_outputs[4492]);
    assign outputs[9253] = layer2_outputs[10771];
    assign outputs[9254] = layer2_outputs[3897];
    assign outputs[9255] = ~(layer2_outputs[4977]);
    assign outputs[9256] = ~(layer2_outputs[8098]);
    assign outputs[9257] = ~(layer2_outputs[7664]);
    assign outputs[9258] = layer2_outputs[7523];
    assign outputs[9259] = (layer2_outputs[4917]) ^ (layer2_outputs[8997]);
    assign outputs[9260] = ~((layer2_outputs[7625]) | (layer2_outputs[11482]));
    assign outputs[9261] = (layer2_outputs[11565]) ^ (layer2_outputs[4649]);
    assign outputs[9262] = (layer2_outputs[7763]) ^ (layer2_outputs[11812]);
    assign outputs[9263] = ~(layer2_outputs[8840]);
    assign outputs[9264] = ~((layer2_outputs[3579]) ^ (layer2_outputs[5983]));
    assign outputs[9265] = ~((layer2_outputs[2574]) ^ (layer2_outputs[5576]));
    assign outputs[9266] = (layer2_outputs[8319]) ^ (layer2_outputs[10994]);
    assign outputs[9267] = (layer2_outputs[11540]) ^ (layer2_outputs[4233]);
    assign outputs[9268] = (layer2_outputs[494]) & (layer2_outputs[8213]);
    assign outputs[9269] = (layer2_outputs[6121]) ^ (layer2_outputs[3219]);
    assign outputs[9270] = ~(layer2_outputs[11965]);
    assign outputs[9271] = ~((layer2_outputs[6344]) | (layer2_outputs[4712]));
    assign outputs[9272] = ~(layer2_outputs[8631]) | (layer2_outputs[6585]);
    assign outputs[9273] = (layer2_outputs[397]) ^ (layer2_outputs[373]);
    assign outputs[9274] = layer2_outputs[2278];
    assign outputs[9275] = ~((layer2_outputs[5790]) ^ (layer2_outputs[1272]));
    assign outputs[9276] = ~(layer2_outputs[3077]);
    assign outputs[9277] = (layer2_outputs[3207]) ^ (layer2_outputs[5928]);
    assign outputs[9278] = ~(layer2_outputs[5161]);
    assign outputs[9279] = (layer2_outputs[5932]) & ~(layer2_outputs[4688]);
    assign outputs[9280] = ~((layer2_outputs[8490]) ^ (layer2_outputs[8711]));
    assign outputs[9281] = (layer2_outputs[848]) ^ (layer2_outputs[10727]);
    assign outputs[9282] = layer2_outputs[12583];
    assign outputs[9283] = ~(layer2_outputs[509]);
    assign outputs[9284] = ~((layer2_outputs[7034]) ^ (layer2_outputs[969]));
    assign outputs[9285] = (layer2_outputs[1457]) & (layer2_outputs[11103]);
    assign outputs[9286] = layer2_outputs[7727];
    assign outputs[9287] = ~((layer2_outputs[6450]) ^ (layer2_outputs[5724]));
    assign outputs[9288] = ~(layer2_outputs[10052]);
    assign outputs[9289] = ~((layer2_outputs[2419]) ^ (layer2_outputs[11762]));
    assign outputs[9290] = layer2_outputs[3240];
    assign outputs[9291] = layer2_outputs[12003];
    assign outputs[9292] = ~((layer2_outputs[12156]) ^ (layer2_outputs[11863]));
    assign outputs[9293] = ~(layer2_outputs[5150]);
    assign outputs[9294] = (layer2_outputs[5035]) & ~(layer2_outputs[2562]);
    assign outputs[9295] = layer2_outputs[7773];
    assign outputs[9296] = layer2_outputs[9000];
    assign outputs[9297] = ~(layer2_outputs[9703]);
    assign outputs[9298] = layer2_outputs[9314];
    assign outputs[9299] = (layer2_outputs[2361]) & (layer2_outputs[2452]);
    assign outputs[9300] = layer2_outputs[10793];
    assign outputs[9301] = ~(layer2_outputs[745]) | (layer2_outputs[5949]);
    assign outputs[9302] = ~(layer2_outputs[7476]);
    assign outputs[9303] = layer2_outputs[11710];
    assign outputs[9304] = layer2_outputs[8235];
    assign outputs[9305] = (layer2_outputs[12441]) ^ (layer2_outputs[11849]);
    assign outputs[9306] = ~(layer2_outputs[246]);
    assign outputs[9307] = ~(layer2_outputs[490]);
    assign outputs[9308] = ~(layer2_outputs[2835]);
    assign outputs[9309] = layer2_outputs[5157];
    assign outputs[9310] = ~(layer2_outputs[9853]);
    assign outputs[9311] = ~((layer2_outputs[6527]) ^ (layer2_outputs[6408]));
    assign outputs[9312] = ~(layer2_outputs[6586]);
    assign outputs[9313] = layer2_outputs[1602];
    assign outputs[9314] = (layer2_outputs[6812]) ^ (layer2_outputs[12197]);
    assign outputs[9315] = (layer2_outputs[11085]) ^ (layer2_outputs[2139]);
    assign outputs[9316] = ~((layer2_outputs[2928]) ^ (layer2_outputs[8038]));
    assign outputs[9317] = (layer2_outputs[11204]) ^ (layer2_outputs[9262]);
    assign outputs[9318] = ~((layer2_outputs[11589]) ^ (layer2_outputs[11816]));
    assign outputs[9319] = ~((layer2_outputs[438]) & (layer2_outputs[2502]));
    assign outputs[9320] = ~(layer2_outputs[6773]);
    assign outputs[9321] = ~(layer2_outputs[2484]);
    assign outputs[9322] = ~((layer2_outputs[1548]) ^ (layer2_outputs[5563]));
    assign outputs[9323] = (layer2_outputs[3324]) | (layer2_outputs[11956]);
    assign outputs[9324] = layer2_outputs[11414];
    assign outputs[9325] = ~(layer2_outputs[9550]);
    assign outputs[9326] = layer2_outputs[9502];
    assign outputs[9327] = layer2_outputs[2468];
    assign outputs[9328] = layer2_outputs[6389];
    assign outputs[9329] = (layer2_outputs[10312]) ^ (layer2_outputs[604]);
    assign outputs[9330] = ~(layer2_outputs[3117]);
    assign outputs[9331] = ~((layer2_outputs[5940]) & (layer2_outputs[8908]));
    assign outputs[9332] = (layer2_outputs[7712]) ^ (layer2_outputs[6184]);
    assign outputs[9333] = (layer2_outputs[2913]) ^ (layer2_outputs[9760]);
    assign outputs[9334] = ~((layer2_outputs[8130]) ^ (layer2_outputs[3028]));
    assign outputs[9335] = ~((layer2_outputs[11828]) ^ (layer2_outputs[3728]));
    assign outputs[9336] = ~((layer2_outputs[4009]) ^ (layer2_outputs[10425]));
    assign outputs[9337] = (layer2_outputs[12444]) ^ (layer2_outputs[2758]);
    assign outputs[9338] = ~((layer2_outputs[5101]) & (layer2_outputs[8119]));
    assign outputs[9339] = (layer2_outputs[10498]) & ~(layer2_outputs[2780]);
    assign outputs[9340] = ~((layer2_outputs[5441]) ^ (layer2_outputs[5918]));
    assign outputs[9341] = ~(layer2_outputs[368]);
    assign outputs[9342] = layer2_outputs[286];
    assign outputs[9343] = layer2_outputs[3357];
    assign outputs[9344] = ~((layer2_outputs[9300]) ^ (layer2_outputs[3447]));
    assign outputs[9345] = layer2_outputs[4141];
    assign outputs[9346] = layer2_outputs[5789];
    assign outputs[9347] = ~(layer2_outputs[4482]);
    assign outputs[9348] = ~(layer2_outputs[4964]);
    assign outputs[9349] = ~(layer2_outputs[9062]);
    assign outputs[9350] = ~((layer2_outputs[181]) ^ (layer2_outputs[3359]));
    assign outputs[9351] = (layer2_outputs[11952]) & ~(layer2_outputs[5813]);
    assign outputs[9352] = ~((layer2_outputs[2610]) ^ (layer2_outputs[1052]));
    assign outputs[9353] = ~((layer2_outputs[5424]) | (layer2_outputs[1993]));
    assign outputs[9354] = (layer2_outputs[2606]) ^ (layer2_outputs[2944]);
    assign outputs[9355] = ~((layer2_outputs[12143]) ^ (layer2_outputs[9108]));
    assign outputs[9356] = ~(layer2_outputs[9571]);
    assign outputs[9357] = (layer2_outputs[1800]) & ~(layer2_outputs[4833]);
    assign outputs[9358] = ~(layer2_outputs[10094]);
    assign outputs[9359] = ~(layer2_outputs[3337]);
    assign outputs[9360] = layer2_outputs[2632];
    assign outputs[9361] = ~((layer2_outputs[3122]) ^ (layer2_outputs[8128]));
    assign outputs[9362] = ~(layer2_outputs[9892]);
    assign outputs[9363] = layer2_outputs[5537];
    assign outputs[9364] = layer2_outputs[2329];
    assign outputs[9365] = ~((layer2_outputs[2073]) ^ (layer2_outputs[6414]));
    assign outputs[9366] = (layer2_outputs[12671]) & ~(layer2_outputs[6414]);
    assign outputs[9367] = layer2_outputs[1756];
    assign outputs[9368] = layer2_outputs[8258];
    assign outputs[9369] = layer2_outputs[297];
    assign outputs[9370] = layer2_outputs[10443];
    assign outputs[9371] = ~(layer2_outputs[4829]) | (layer2_outputs[5622]);
    assign outputs[9372] = layer2_outputs[1652];
    assign outputs[9373] = layer2_outputs[6264];
    assign outputs[9374] = layer2_outputs[6105];
    assign outputs[9375] = (layer2_outputs[3654]) & ~(layer2_outputs[3465]);
    assign outputs[9376] = ~(layer2_outputs[6688]);
    assign outputs[9377] = (layer2_outputs[11355]) ^ (layer2_outputs[9065]);
    assign outputs[9378] = (layer2_outputs[7521]) ^ (layer2_outputs[2296]);
    assign outputs[9379] = ~(layer2_outputs[3761]);
    assign outputs[9380] = ~(layer2_outputs[4418]);
    assign outputs[9381] = layer2_outputs[2639];
    assign outputs[9382] = layer2_outputs[1342];
    assign outputs[9383] = ~(layer2_outputs[8931]);
    assign outputs[9384] = ~((layer2_outputs[8115]) ^ (layer2_outputs[2683]));
    assign outputs[9385] = ~((layer2_outputs[8137]) ^ (layer2_outputs[3309]));
    assign outputs[9386] = ~((layer2_outputs[6553]) | (layer2_outputs[12096]));
    assign outputs[9387] = ~((layer2_outputs[12429]) | (layer2_outputs[6382]));
    assign outputs[9388] = ~(layer2_outputs[11027]);
    assign outputs[9389] = layer2_outputs[6634];
    assign outputs[9390] = ~((layer2_outputs[12293]) ^ (layer2_outputs[2863]));
    assign outputs[9391] = (layer2_outputs[4723]) ^ (layer2_outputs[7939]);
    assign outputs[9392] = layer2_outputs[2475];
    assign outputs[9393] = ~((layer2_outputs[9010]) | (layer2_outputs[12395]));
    assign outputs[9394] = (layer2_outputs[2653]) & (layer2_outputs[5222]);
    assign outputs[9395] = layer2_outputs[798];
    assign outputs[9396] = layer2_outputs[10119];
    assign outputs[9397] = (layer2_outputs[11652]) ^ (layer2_outputs[4629]);
    assign outputs[9398] = ~(layer2_outputs[2111]);
    assign outputs[9399] = ~(layer2_outputs[6649]);
    assign outputs[9400] = (layer2_outputs[2558]) ^ (layer2_outputs[2661]);
    assign outputs[9401] = ~((layer2_outputs[11979]) ^ (layer2_outputs[3746]));
    assign outputs[9402] = ~((layer2_outputs[4283]) ^ (layer2_outputs[3247]));
    assign outputs[9403] = (layer2_outputs[6971]) | (layer2_outputs[7528]);
    assign outputs[9404] = ~((layer2_outputs[5496]) ^ (layer2_outputs[10617]));
    assign outputs[9405] = ~(layer2_outputs[1831]);
    assign outputs[9406] = (layer2_outputs[6084]) ^ (layer2_outputs[3583]);
    assign outputs[9407] = ~((layer2_outputs[174]) | (layer2_outputs[2192]));
    assign outputs[9408] = layer2_outputs[7222];
    assign outputs[9409] = ~((layer2_outputs[11657]) | (layer2_outputs[764]));
    assign outputs[9410] = layer2_outputs[6024];
    assign outputs[9411] = (layer2_outputs[3954]) & ~(layer2_outputs[9900]);
    assign outputs[9412] = (layer2_outputs[2636]) ^ (layer2_outputs[1475]);
    assign outputs[9413] = ~((layer2_outputs[11809]) ^ (layer2_outputs[3561]));
    assign outputs[9414] = ~(layer2_outputs[9552]);
    assign outputs[9415] = ~((layer2_outputs[972]) | (layer2_outputs[3703]));
    assign outputs[9416] = ~((layer2_outputs[138]) ^ (layer2_outputs[9207]));
    assign outputs[9417] = layer2_outputs[10700];
    assign outputs[9418] = layer2_outputs[10909];
    assign outputs[9419] = ~(layer2_outputs[5045]);
    assign outputs[9420] = layer2_outputs[11941];
    assign outputs[9421] = layer2_outputs[12424];
    assign outputs[9422] = ~((layer2_outputs[786]) ^ (layer2_outputs[8910]));
    assign outputs[9423] = (layer2_outputs[5026]) | (layer2_outputs[12330]);
    assign outputs[9424] = ~(layer2_outputs[3512]);
    assign outputs[9425] = ~((layer2_outputs[1336]) ^ (layer2_outputs[1802]));
    assign outputs[9426] = (layer2_outputs[7600]) ^ (layer2_outputs[872]);
    assign outputs[9427] = layer2_outputs[11351];
    assign outputs[9428] = ~(layer2_outputs[5143]);
    assign outputs[9429] = ~(layer2_outputs[1539]);
    assign outputs[9430] = ~((layer2_outputs[1342]) ^ (layer2_outputs[757]));
    assign outputs[9431] = ~(layer2_outputs[1640]);
    assign outputs[9432] = (layer2_outputs[7468]) & ~(layer2_outputs[5817]);
    assign outputs[9433] = ~(layer2_outputs[11946]);
    assign outputs[9434] = (layer2_outputs[2268]) & ~(layer2_outputs[7461]);
    assign outputs[9435] = ~(layer2_outputs[9929]);
    assign outputs[9436] = layer2_outputs[6570];
    assign outputs[9437] = (layer2_outputs[9940]) ^ (layer2_outputs[5997]);
    assign outputs[9438] = layer2_outputs[5666];
    assign outputs[9439] = (layer2_outputs[3154]) & ~(layer2_outputs[9475]);
    assign outputs[9440] = layer2_outputs[12499];
    assign outputs[9441] = ~(layer2_outputs[9737]);
    assign outputs[9442] = (layer2_outputs[10039]) & (layer2_outputs[2804]);
    assign outputs[9443] = layer2_outputs[2082];
    assign outputs[9444] = ~(layer2_outputs[9673]);
    assign outputs[9445] = layer2_outputs[2007];
    assign outputs[9446] = ~(layer2_outputs[10616]);
    assign outputs[9447] = (layer2_outputs[1642]) | (layer2_outputs[5247]);
    assign outputs[9448] = ~((layer2_outputs[8982]) ^ (layer2_outputs[609]));
    assign outputs[9449] = (layer2_outputs[3914]) & ~(layer2_outputs[4760]);
    assign outputs[9450] = ~((layer2_outputs[1398]) ^ (layer2_outputs[11974]));
    assign outputs[9451] = layer2_outputs[12282];
    assign outputs[9452] = ~(layer2_outputs[6596]);
    assign outputs[9453] = (layer2_outputs[901]) | (layer2_outputs[11515]);
    assign outputs[9454] = ~(layer2_outputs[11474]);
    assign outputs[9455] = ~(layer2_outputs[1867]);
    assign outputs[9456] = ~(layer2_outputs[12690]);
    assign outputs[9457] = layer2_outputs[4625];
    assign outputs[9458] = ~(layer2_outputs[11656]);
    assign outputs[9459] = ~(layer2_outputs[7284]);
    assign outputs[9460] = ~(layer2_outputs[11501]);
    assign outputs[9461] = ~(layer2_outputs[6918]);
    assign outputs[9462] = ~(layer2_outputs[1137]);
    assign outputs[9463] = ~((layer2_outputs[9291]) ^ (layer2_outputs[3783]));
    assign outputs[9464] = layer2_outputs[2307];
    assign outputs[9465] = layer2_outputs[182];
    assign outputs[9466] = layer2_outputs[4819];
    assign outputs[9467] = ~(layer2_outputs[2537]);
    assign outputs[9468] = ~((layer2_outputs[1931]) ^ (layer2_outputs[5349]));
    assign outputs[9469] = (layer2_outputs[8114]) ^ (layer2_outputs[3918]);
    assign outputs[9470] = (layer2_outputs[1572]) & (layer2_outputs[6358]);
    assign outputs[9471] = (layer2_outputs[3174]) ^ (layer2_outputs[8854]);
    assign outputs[9472] = layer2_outputs[7139];
    assign outputs[9473] = (layer2_outputs[2846]) & (layer2_outputs[1179]);
    assign outputs[9474] = ~(layer2_outputs[3903]);
    assign outputs[9475] = ~(layer2_outputs[11940]);
    assign outputs[9476] = ~(layer2_outputs[12141]);
    assign outputs[9477] = layer2_outputs[11453];
    assign outputs[9478] = layer2_outputs[8802];
    assign outputs[9479] = ~(layer2_outputs[1791]);
    assign outputs[9480] = layer2_outputs[6468];
    assign outputs[9481] = layer2_outputs[2198];
    assign outputs[9482] = layer2_outputs[1748];
    assign outputs[9483] = (layer2_outputs[4799]) & ~(layer2_outputs[8561]);
    assign outputs[9484] = (layer2_outputs[6562]) ^ (layer2_outputs[5460]);
    assign outputs[9485] = ~(layer2_outputs[1137]);
    assign outputs[9486] = layer2_outputs[3493];
    assign outputs[9487] = ~((layer2_outputs[1946]) | (layer2_outputs[6287]));
    assign outputs[9488] = layer2_outputs[10372];
    assign outputs[9489] = (layer2_outputs[2218]) | (layer2_outputs[7762]);
    assign outputs[9490] = (layer2_outputs[12119]) ^ (layer2_outputs[10848]);
    assign outputs[9491] = ~(layer2_outputs[9931]);
    assign outputs[9492] = layer2_outputs[5089];
    assign outputs[9493] = ~(layer2_outputs[4171]);
    assign outputs[9494] = (layer2_outputs[4083]) ^ (layer2_outputs[10131]);
    assign outputs[9495] = layer2_outputs[8162];
    assign outputs[9496] = layer2_outputs[12109];
    assign outputs[9497] = ~(layer2_outputs[12114]) | (layer2_outputs[7230]);
    assign outputs[9498] = ~(layer2_outputs[3143]);
    assign outputs[9499] = ~(layer2_outputs[1278]);
    assign outputs[9500] = ~((layer2_outputs[2997]) ^ (layer2_outputs[6339]));
    assign outputs[9501] = ~((layer2_outputs[8938]) & (layer2_outputs[7363]));
    assign outputs[9502] = ~(layer2_outputs[8754]);
    assign outputs[9503] = ~(layer2_outputs[2674]);
    assign outputs[9504] = (layer2_outputs[8045]) & ~(layer2_outputs[11854]);
    assign outputs[9505] = ~(layer2_outputs[7023]);
    assign outputs[9506] = ~((layer2_outputs[9870]) & (layer2_outputs[2831]));
    assign outputs[9507] = layer2_outputs[8567];
    assign outputs[9508] = ~(layer2_outputs[1521]);
    assign outputs[9509] = layer2_outputs[3462];
    assign outputs[9510] = (layer2_outputs[10637]) ^ (layer2_outputs[224]);
    assign outputs[9511] = layer2_outputs[4032];
    assign outputs[9512] = layer2_outputs[9983];
    assign outputs[9513] = ~(layer2_outputs[7530]);
    assign outputs[9514] = layer2_outputs[4018];
    assign outputs[9515] = ~(layer2_outputs[10613]);
    assign outputs[9516] = layer2_outputs[2118];
    assign outputs[9517] = ~(layer2_outputs[4175]);
    assign outputs[9518] = ~(layer2_outputs[3670]);
    assign outputs[9519] = layer2_outputs[8297];
    assign outputs[9520] = (layer2_outputs[2216]) ^ (layer2_outputs[12069]);
    assign outputs[9521] = ~(layer2_outputs[7394]) | (layer2_outputs[12619]);
    assign outputs[9522] = ~((layer2_outputs[10393]) | (layer2_outputs[1638]));
    assign outputs[9523] = layer2_outputs[4583];
    assign outputs[9524] = ~(layer2_outputs[6350]);
    assign outputs[9525] = (layer2_outputs[12553]) ^ (layer2_outputs[8806]);
    assign outputs[9526] = ~((layer2_outputs[5484]) ^ (layer2_outputs[7409]));
    assign outputs[9527] = layer2_outputs[6996];
    assign outputs[9528] = ~(layer2_outputs[8553]);
    assign outputs[9529] = ~(layer2_outputs[9667]);
    assign outputs[9530] = layer2_outputs[766];
    assign outputs[9531] = ~(layer2_outputs[11450]);
    assign outputs[9532] = layer2_outputs[412];
    assign outputs[9533] = ~((layer2_outputs[8573]) ^ (layer2_outputs[5870]));
    assign outputs[9534] = layer2_outputs[9792];
    assign outputs[9535] = ~((layer2_outputs[10467]) ^ (layer2_outputs[8314]));
    assign outputs[9536] = ~(layer2_outputs[6245]);
    assign outputs[9537] = ~(layer2_outputs[4515]);
    assign outputs[9538] = ~(layer2_outputs[8373]);
    assign outputs[9539] = ~(layer2_outputs[1555]);
    assign outputs[9540] = layer2_outputs[12167];
    assign outputs[9541] = ~(layer2_outputs[3256]);
    assign outputs[9542] = ~(layer2_outputs[9838]);
    assign outputs[9543] = ~(layer2_outputs[7779]);
    assign outputs[9544] = ~(layer2_outputs[10588]);
    assign outputs[9545] = layer2_outputs[10097];
    assign outputs[9546] = ~((layer2_outputs[6946]) ^ (layer2_outputs[2066]));
    assign outputs[9547] = ~(layer2_outputs[10565]);
    assign outputs[9548] = ~(layer2_outputs[5646]);
    assign outputs[9549] = ~(layer2_outputs[11147]);
    assign outputs[9550] = ~(layer2_outputs[10916]);
    assign outputs[9551] = (layer2_outputs[8369]) & ~(layer2_outputs[2203]);
    assign outputs[9552] = ~(layer2_outputs[4702]);
    assign outputs[9553] = ~(layer2_outputs[7954]);
    assign outputs[9554] = (layer2_outputs[6743]) & ~(layer2_outputs[10741]);
    assign outputs[9555] = ~(layer2_outputs[10880]);
    assign outputs[9556] = ~(layer2_outputs[4016]) | (layer2_outputs[10304]);
    assign outputs[9557] = ~((layer2_outputs[5860]) ^ (layer2_outputs[6597]));
    assign outputs[9558] = layer2_outputs[10838];
    assign outputs[9559] = ~((layer2_outputs[344]) ^ (layer2_outputs[3957]));
    assign outputs[9560] = ~(layer2_outputs[6490]) | (layer2_outputs[8298]);
    assign outputs[9561] = (layer2_outputs[4661]) ^ (layer2_outputs[1107]);
    assign outputs[9562] = ~(layer2_outputs[4777]);
    assign outputs[9563] = (layer2_outputs[6566]) | (layer2_outputs[10914]);
    assign outputs[9564] = ~(layer2_outputs[2621]);
    assign outputs[9565] = layer2_outputs[3780];
    assign outputs[9566] = layer2_outputs[4421];
    assign outputs[9567] = (layer2_outputs[4679]) ^ (layer2_outputs[9577]);
    assign outputs[9568] = layer2_outputs[7197];
    assign outputs[9569] = (layer2_outputs[2554]) ^ (layer2_outputs[3157]);
    assign outputs[9570] = layer2_outputs[10133];
    assign outputs[9571] = ~(layer2_outputs[131]);
    assign outputs[9572] = ~(layer2_outputs[6039]);
    assign outputs[9573] = layer2_outputs[11415];
    assign outputs[9574] = layer2_outputs[7913];
    assign outputs[9575] = (layer2_outputs[2351]) & ~(layer2_outputs[12301]);
    assign outputs[9576] = layer2_outputs[5836];
    assign outputs[9577] = (layer2_outputs[10830]) ^ (layer2_outputs[5142]);
    assign outputs[9578] = layer2_outputs[2880];
    assign outputs[9579] = (layer2_outputs[6668]) & (layer2_outputs[6483]);
    assign outputs[9580] = ~(layer2_outputs[151]);
    assign outputs[9581] = layer2_outputs[11901];
    assign outputs[9582] = ~(layer2_outputs[3163]) | (layer2_outputs[3706]);
    assign outputs[9583] = (layer2_outputs[5946]) & ~(layer2_outputs[6321]);
    assign outputs[9584] = layer2_outputs[6307];
    assign outputs[9585] = ~((layer2_outputs[12783]) | (layer2_outputs[12761]));
    assign outputs[9586] = layer2_outputs[11085];
    assign outputs[9587] = ~(layer2_outputs[7302]) | (layer2_outputs[12492]);
    assign outputs[9588] = ~(layer2_outputs[9378]);
    assign outputs[9589] = layer2_outputs[7376];
    assign outputs[9590] = layer2_outputs[4114];
    assign outputs[9591] = layer2_outputs[8818];
    assign outputs[9592] = layer2_outputs[10800];
    assign outputs[9593] = (layer2_outputs[930]) ^ (layer2_outputs[7126]);
    assign outputs[9594] = ~((layer2_outputs[9985]) | (layer2_outputs[10622]));
    assign outputs[9595] = layer2_outputs[9716];
    assign outputs[9596] = layer2_outputs[4997];
    assign outputs[9597] = ~((layer2_outputs[4860]) ^ (layer2_outputs[9017]));
    assign outputs[9598] = layer2_outputs[8308];
    assign outputs[9599] = layer2_outputs[7516];
    assign outputs[9600] = layer2_outputs[5545];
    assign outputs[9601] = layer2_outputs[5478];
    assign outputs[9602] = (layer2_outputs[1128]) ^ (layer2_outputs[6131]);
    assign outputs[9603] = ~((layer2_outputs[9434]) ^ (layer2_outputs[721]));
    assign outputs[9604] = ~(layer2_outputs[4155]);
    assign outputs[9605] = layer2_outputs[4875];
    assign outputs[9606] = (layer2_outputs[4790]) ^ (layer2_outputs[10150]);
    assign outputs[9607] = ~(layer2_outputs[6972]);
    assign outputs[9608] = layer2_outputs[11695];
    assign outputs[9609] = ~(layer2_outputs[4801]);
    assign outputs[9610] = layer2_outputs[10871];
    assign outputs[9611] = ~(layer2_outputs[1867]);
    assign outputs[9612] = layer2_outputs[1220];
    assign outputs[9613] = layer2_outputs[12451];
    assign outputs[9614] = layer2_outputs[3606];
    assign outputs[9615] = ~(layer2_outputs[5119]);
    assign outputs[9616] = ~(layer2_outputs[5512]);
    assign outputs[9617] = (layer2_outputs[897]) ^ (layer2_outputs[1875]);
    assign outputs[9618] = ~(layer2_outputs[7829]);
    assign outputs[9619] = (layer2_outputs[6816]) ^ (layer2_outputs[8979]);
    assign outputs[9620] = ~((layer2_outputs[5892]) | (layer2_outputs[5978]));
    assign outputs[9621] = ~(layer2_outputs[8809]);
    assign outputs[9622] = ~(layer2_outputs[4810]);
    assign outputs[9623] = (layer2_outputs[4347]) ^ (layer2_outputs[2561]);
    assign outputs[9624] = ~(layer2_outputs[11961]);
    assign outputs[9625] = layer2_outputs[1739];
    assign outputs[9626] = layer2_outputs[10444];
    assign outputs[9627] = (layer2_outputs[2537]) ^ (layer2_outputs[2174]);
    assign outputs[9628] = (layer2_outputs[996]) ^ (layer2_outputs[3388]);
    assign outputs[9629] = layer2_outputs[6478];
    assign outputs[9630] = (layer2_outputs[12233]) & (layer2_outputs[6292]);
    assign outputs[9631] = ~(layer2_outputs[9893]);
    assign outputs[9632] = layer2_outputs[9962];
    assign outputs[9633] = (layer2_outputs[2572]) ^ (layer2_outputs[1884]);
    assign outputs[9634] = (layer2_outputs[6529]) | (layer2_outputs[12529]);
    assign outputs[9635] = ~(layer2_outputs[2752]);
    assign outputs[9636] = ~(layer2_outputs[2796]);
    assign outputs[9637] = layer2_outputs[6513];
    assign outputs[9638] = layer2_outputs[3542];
    assign outputs[9639] = ~(layer2_outputs[5573]);
    assign outputs[9640] = (layer2_outputs[2093]) ^ (layer2_outputs[5987]);
    assign outputs[9641] = layer2_outputs[12547];
    assign outputs[9642] = layer2_outputs[9422];
    assign outputs[9643] = layer2_outputs[10645];
    assign outputs[9644] = layer2_outputs[2133];
    assign outputs[9645] = ~(layer2_outputs[7078]);
    assign outputs[9646] = layer2_outputs[9163];
    assign outputs[9647] = layer2_outputs[9277];
    assign outputs[9648] = layer2_outputs[12414];
    assign outputs[9649] = (layer2_outputs[7206]) ^ (layer2_outputs[244]);
    assign outputs[9650] = ~(layer2_outputs[8826]);
    assign outputs[9651] = ~(layer2_outputs[2953]);
    assign outputs[9652] = ~(layer2_outputs[1831]);
    assign outputs[9653] = layer2_outputs[2081];
    assign outputs[9654] = (layer2_outputs[489]) & (layer2_outputs[2371]);
    assign outputs[9655] = (layer2_outputs[4467]) ^ (layer2_outputs[4325]);
    assign outputs[9656] = layer2_outputs[5096];
    assign outputs[9657] = layer2_outputs[12596];
    assign outputs[9658] = ~(layer2_outputs[7490]);
    assign outputs[9659] = layer2_outputs[4568];
    assign outputs[9660] = (layer2_outputs[9157]) ^ (layer2_outputs[11325]);
    assign outputs[9661] = ~((layer2_outputs[9734]) ^ (layer2_outputs[6634]));
    assign outputs[9662] = ~(layer2_outputs[8826]);
    assign outputs[9663] = layer2_outputs[9594];
    assign outputs[9664] = ~(layer2_outputs[1811]);
    assign outputs[9665] = ~(layer2_outputs[12690]);
    assign outputs[9666] = ~(layer2_outputs[938]);
    assign outputs[9667] = (layer2_outputs[75]) ^ (layer2_outputs[8447]);
    assign outputs[9668] = ~(layer2_outputs[4772]);
    assign outputs[9669] = (layer2_outputs[6017]) ^ (layer2_outputs[10403]);
    assign outputs[9670] = ~(layer2_outputs[5417]);
    assign outputs[9671] = ~((layer2_outputs[10699]) | (layer2_outputs[11305]));
    assign outputs[9672] = ~(layer2_outputs[4463]);
    assign outputs[9673] = layer2_outputs[304];
    assign outputs[9674] = ~((layer2_outputs[1479]) ^ (layer2_outputs[3812]));
    assign outputs[9675] = (layer2_outputs[6532]) ^ (layer2_outputs[7497]);
    assign outputs[9676] = (layer2_outputs[2656]) ^ (layer2_outputs[7398]);
    assign outputs[9677] = ~((layer2_outputs[2145]) ^ (layer2_outputs[3486]));
    assign outputs[9678] = ~((layer2_outputs[1632]) & (layer2_outputs[1332]));
    assign outputs[9679] = (layer2_outputs[7993]) & ~(layer2_outputs[6854]);
    assign outputs[9680] = (layer2_outputs[1801]) ^ (layer2_outputs[2413]);
    assign outputs[9681] = ~(layer2_outputs[8999]);
    assign outputs[9682] = ~(layer2_outputs[916]);
    assign outputs[9683] = ~(layer2_outputs[2496]) | (layer2_outputs[10822]);
    assign outputs[9684] = (layer2_outputs[2526]) ^ (layer2_outputs[3202]);
    assign outputs[9685] = layer2_outputs[9661];
    assign outputs[9686] = ~((layer2_outputs[217]) ^ (layer2_outputs[4550]));
    assign outputs[9687] = layer2_outputs[139];
    assign outputs[9688] = layer2_outputs[10722];
    assign outputs[9689] = ~(layer2_outputs[7246]) | (layer2_outputs[624]);
    assign outputs[9690] = ~(layer2_outputs[12620]);
    assign outputs[9691] = ~(layer2_outputs[10784]);
    assign outputs[9692] = (layer2_outputs[12715]) ^ (layer2_outputs[2260]);
    assign outputs[9693] = (layer2_outputs[7069]) & ~(layer2_outputs[8587]);
    assign outputs[9694] = ~((layer2_outputs[11634]) ^ (layer2_outputs[1094]));
    assign outputs[9695] = layer2_outputs[12055];
    assign outputs[9696] = layer2_outputs[5228];
    assign outputs[9697] = layer2_outputs[2072];
    assign outputs[9698] = ~(layer2_outputs[10448]);
    assign outputs[9699] = layer2_outputs[3250];
    assign outputs[9700] = (layer2_outputs[4253]) ^ (layer2_outputs[2726]);
    assign outputs[9701] = ~(layer2_outputs[3699]);
    assign outputs[9702] = ~(layer2_outputs[1650]) | (layer2_outputs[10909]);
    assign outputs[9703] = ~((layer2_outputs[3535]) | (layer2_outputs[6795]));
    assign outputs[9704] = (layer2_outputs[11069]) ^ (layer2_outputs[6824]);
    assign outputs[9705] = layer2_outputs[8290];
    assign outputs[9706] = ~((layer2_outputs[5514]) ^ (layer2_outputs[9980]));
    assign outputs[9707] = ~((layer2_outputs[9639]) ^ (layer2_outputs[7177]));
    assign outputs[9708] = ~(layer2_outputs[12717]);
    assign outputs[9709] = (layer2_outputs[8522]) ^ (layer2_outputs[10789]);
    assign outputs[9710] = ~(layer2_outputs[1667]);
    assign outputs[9711] = (layer2_outputs[10728]) & ~(layer2_outputs[1707]);
    assign outputs[9712] = ~((layer2_outputs[9352]) | (layer2_outputs[1699]));
    assign outputs[9713] = ~((layer2_outputs[5956]) ^ (layer2_outputs[4633]));
    assign outputs[9714] = layer2_outputs[4545];
    assign outputs[9715] = layer2_outputs[9004];
    assign outputs[9716] = ~(layer2_outputs[4320]);
    assign outputs[9717] = ~(layer2_outputs[11656]);
    assign outputs[9718] = (layer2_outputs[8491]) & ~(layer2_outputs[8766]);
    assign outputs[9719] = (layer2_outputs[2101]) & ~(layer2_outputs[2314]);
    assign outputs[9720] = ~((layer2_outputs[4941]) | (layer2_outputs[7507]));
    assign outputs[9721] = layer2_outputs[9857];
    assign outputs[9722] = layer2_outputs[12593];
    assign outputs[9723] = ~((layer2_outputs[1974]) & (layer2_outputs[8681]));
    assign outputs[9724] = layer2_outputs[8775];
    assign outputs[9725] = ~(layer2_outputs[11139]) | (layer2_outputs[7700]);
    assign outputs[9726] = ~(layer2_outputs[5290]);
    assign outputs[9727] = layer2_outputs[9358];
    assign outputs[9728] = (layer2_outputs[8577]) & ~(layer2_outputs[6763]);
    assign outputs[9729] = layer2_outputs[452];
    assign outputs[9730] = ~((layer2_outputs[8122]) | (layer2_outputs[12442]));
    assign outputs[9731] = layer2_outputs[1580];
    assign outputs[9732] = layer2_outputs[98];
    assign outputs[9733] = (layer2_outputs[12379]) | (layer2_outputs[6157]);
    assign outputs[9734] = (layer2_outputs[4486]) ^ (layer2_outputs[11369]);
    assign outputs[9735] = ~((layer2_outputs[6241]) | (layer2_outputs[8554]));
    assign outputs[9736] = layer2_outputs[3323];
    assign outputs[9737] = (layer2_outputs[2007]) & (layer2_outputs[9955]);
    assign outputs[9738] = (layer2_outputs[934]) & ~(layer2_outputs[2191]);
    assign outputs[9739] = ~(layer2_outputs[10110]);
    assign outputs[9740] = ~((layer2_outputs[5898]) ^ (layer2_outputs[3665]));
    assign outputs[9741] = layer2_outputs[11093];
    assign outputs[9742] = layer2_outputs[3089];
    assign outputs[9743] = ~(layer2_outputs[9580]);
    assign outputs[9744] = ~(layer2_outputs[6362]);
    assign outputs[9745] = layer2_outputs[11651];
    assign outputs[9746] = layer2_outputs[7063];
    assign outputs[9747] = ~(layer2_outputs[9338]);
    assign outputs[9748] = ~(layer2_outputs[6753]);
    assign outputs[9749] = ~((layer2_outputs[4554]) | (layer2_outputs[11064]));
    assign outputs[9750] = layer2_outputs[7607];
    assign outputs[9751] = layer2_outputs[10195];
    assign outputs[9752] = layer2_outputs[9102];
    assign outputs[9753] = layer2_outputs[4967];
    assign outputs[9754] = ~(layer2_outputs[7082]);
    assign outputs[9755] = ~(layer2_outputs[12253]);
    assign outputs[9756] = ~(layer2_outputs[7589]) | (layer2_outputs[293]);
    assign outputs[9757] = ~(layer2_outputs[2116]);
    assign outputs[9758] = ~((layer2_outputs[7841]) | (layer2_outputs[8887]));
    assign outputs[9759] = (layer2_outputs[104]) ^ (layer2_outputs[4506]);
    assign outputs[9760] = ~((layer2_outputs[5627]) | (layer2_outputs[3742]));
    assign outputs[9761] = ~(layer2_outputs[10920]);
    assign outputs[9762] = ~((layer2_outputs[9901]) | (layer2_outputs[6939]));
    assign outputs[9763] = (layer2_outputs[5360]) ^ (layer2_outputs[3794]);
    assign outputs[9764] = (layer2_outputs[5357]) ^ (layer2_outputs[11770]);
    assign outputs[9765] = ~((layer2_outputs[4364]) | (layer2_outputs[91]));
    assign outputs[9766] = (layer2_outputs[3223]) & ~(layer2_outputs[5033]);
    assign outputs[9767] = (layer2_outputs[9396]) ^ (layer2_outputs[12727]);
    assign outputs[9768] = layer2_outputs[2288];
    assign outputs[9769] = (layer2_outputs[2158]) ^ (layer2_outputs[11155]);
    assign outputs[9770] = ~(layer2_outputs[8047]);
    assign outputs[9771] = ~(layer2_outputs[1889]);
    assign outputs[9772] = ~(layer2_outputs[1895]);
    assign outputs[9773] = ~(layer2_outputs[8804]);
    assign outputs[9774] = layer2_outputs[4179];
    assign outputs[9775] = ~((layer2_outputs[8894]) ^ (layer2_outputs[191]));
    assign outputs[9776] = ~((layer2_outputs[2214]) ^ (layer2_outputs[8977]));
    assign outputs[9777] = ~(layer2_outputs[9522]);
    assign outputs[9778] = (layer2_outputs[550]) ^ (layer2_outputs[8214]);
    assign outputs[9779] = layer2_outputs[8018];
    assign outputs[9780] = layer2_outputs[6291];
    assign outputs[9781] = (layer2_outputs[3124]) | (layer2_outputs[7194]);
    assign outputs[9782] = ~(layer2_outputs[10424]);
    assign outputs[9783] = (layer2_outputs[6645]) & (layer2_outputs[4563]);
    assign outputs[9784] = ~(layer2_outputs[1539]);
    assign outputs[9785] = (layer2_outputs[11299]) & ~(layer2_outputs[6055]);
    assign outputs[9786] = ~(layer2_outputs[9807]);
    assign outputs[9787] = layer2_outputs[61];
    assign outputs[9788] = ~(layer2_outputs[3328]);
    assign outputs[9789] = ~(layer2_outputs[1390]);
    assign outputs[9790] = ~(layer2_outputs[971]);
    assign outputs[9791] = (layer2_outputs[843]) & ~(layer2_outputs[7491]);
    assign outputs[9792] = (layer2_outputs[10552]) & ~(layer2_outputs[7859]);
    assign outputs[9793] = layer2_outputs[1565];
    assign outputs[9794] = ~(layer2_outputs[7783]);
    assign outputs[9795] = ~((layer2_outputs[5907]) ^ (layer2_outputs[12437]));
    assign outputs[9796] = ~(layer2_outputs[6643]);
    assign outputs[9797] = (layer2_outputs[6023]) & (layer2_outputs[3158]);
    assign outputs[9798] = layer2_outputs[9322];
    assign outputs[9799] = ~((layer2_outputs[9428]) ^ (layer2_outputs[5630]));
    assign outputs[9800] = (layer2_outputs[7496]) ^ (layer2_outputs[7146]);
    assign outputs[9801] = layer2_outputs[2803];
    assign outputs[9802] = ~(layer2_outputs[3521]) | (layer2_outputs[7612]);
    assign outputs[9803] = ~(layer2_outputs[1979]);
    assign outputs[9804] = (layer2_outputs[7769]) & ~(layer2_outputs[7973]);
    assign outputs[9805] = layer2_outputs[3297];
    assign outputs[9806] = ~(layer2_outputs[78]);
    assign outputs[9807] = (layer2_outputs[12152]) | (layer2_outputs[3970]);
    assign outputs[9808] = ~(layer2_outputs[1984]);
    assign outputs[9809] = layer2_outputs[4638];
    assign outputs[9810] = (layer2_outputs[10668]) ^ (layer2_outputs[6858]);
    assign outputs[9811] = layer2_outputs[7843];
    assign outputs[9812] = layer2_outputs[10382];
    assign outputs[9813] = layer2_outputs[3891];
    assign outputs[9814] = layer2_outputs[9744];
    assign outputs[9815] = ~(layer2_outputs[7176]) | (layer2_outputs[11653]);
    assign outputs[9816] = (layer2_outputs[10327]) | (layer2_outputs[8873]);
    assign outputs[9817] = (layer2_outputs[10059]) & (layer2_outputs[12742]);
    assign outputs[9818] = ~((layer2_outputs[4343]) | (layer2_outputs[7381]));
    assign outputs[9819] = ~(layer2_outputs[5226]);
    assign outputs[9820] = (layer2_outputs[4046]) & ~(layer2_outputs[6191]);
    assign outputs[9821] = ~(layer2_outputs[6351]);
    assign outputs[9822] = ~(layer2_outputs[1009]);
    assign outputs[9823] = layer2_outputs[8274];
    assign outputs[9824] = layer2_outputs[6963];
    assign outputs[9825] = ~(layer2_outputs[5392]);
    assign outputs[9826] = ~(layer2_outputs[5889]);
    assign outputs[9827] = layer2_outputs[11612];
    assign outputs[9828] = layer2_outputs[12089];
    assign outputs[9829] = ~((layer2_outputs[10092]) | (layer2_outputs[5826]));
    assign outputs[9830] = ~((layer2_outputs[3634]) & (layer2_outputs[8078]));
    assign outputs[9831] = layer2_outputs[11945];
    assign outputs[9832] = ~(layer2_outputs[3310]);
    assign outputs[9833] = layer2_outputs[11518];
    assign outputs[9834] = layer2_outputs[173];
    assign outputs[9835] = ~(layer2_outputs[8289]);
    assign outputs[9836] = layer2_outputs[5212];
    assign outputs[9837] = ~((layer2_outputs[7904]) ^ (layer2_outputs[9410]));
    assign outputs[9838] = ~(layer2_outputs[2703]);
    assign outputs[9839] = (layer2_outputs[1089]) & (layer2_outputs[3149]);
    assign outputs[9840] = ~(layer2_outputs[351]);
    assign outputs[9841] = ~(layer2_outputs[9800]);
    assign outputs[9842] = (layer2_outputs[3449]) ^ (layer2_outputs[1963]);
    assign outputs[9843] = (layer2_outputs[1522]) ^ (layer2_outputs[3727]);
    assign outputs[9844] = (layer2_outputs[9505]) ^ (layer2_outputs[5166]);
    assign outputs[9845] = (layer2_outputs[8142]) & ~(layer2_outputs[5850]);
    assign outputs[9846] = (layer2_outputs[8729]) & ~(layer2_outputs[10328]);
    assign outputs[9847] = (layer2_outputs[8717]) & ~(layer2_outputs[4037]);
    assign outputs[9848] = layer2_outputs[8973];
    assign outputs[9849] = (layer2_outputs[11672]) & ~(layer2_outputs[6937]);
    assign outputs[9850] = ~(layer2_outputs[12483]);
    assign outputs[9851] = layer2_outputs[785];
    assign outputs[9852] = ~((layer2_outputs[3207]) | (layer2_outputs[7875]));
    assign outputs[9853] = layer2_outputs[3429];
    assign outputs[9854] = ~(layer2_outputs[8254]) | (layer2_outputs[8343]);
    assign outputs[9855] = ~(layer2_outputs[3858]);
    assign outputs[9856] = ~(layer2_outputs[11323]);
    assign outputs[9857] = layer2_outputs[1455];
    assign outputs[9858] = ~(layer2_outputs[9722]);
    assign outputs[9859] = ~(layer2_outputs[1509]);
    assign outputs[9860] = ~(layer2_outputs[5512]);
    assign outputs[9861] = (layer2_outputs[6164]) & (layer2_outputs[5152]);
    assign outputs[9862] = ~(layer2_outputs[8659]) | (layer2_outputs[12798]);
    assign outputs[9863] = ~((layer2_outputs[5465]) & (layer2_outputs[4873]));
    assign outputs[9864] = ~(layer2_outputs[9999]);
    assign outputs[9865] = ~(layer2_outputs[10734]);
    assign outputs[9866] = (layer2_outputs[1894]) & (layer2_outputs[10581]);
    assign outputs[9867] = ~(layer2_outputs[2697]) | (layer2_outputs[8940]);
    assign outputs[9868] = layer2_outputs[5844];
    assign outputs[9869] = layer2_outputs[5024];
    assign outputs[9870] = ~((layer2_outputs[7985]) ^ (layer2_outputs[7925]));
    assign outputs[9871] = ~(layer2_outputs[7357]);
    assign outputs[9872] = ~((layer2_outputs[1446]) ^ (layer2_outputs[11416]));
    assign outputs[9873] = layer2_outputs[7727];
    assign outputs[9874] = ~((layer2_outputs[9543]) ^ (layer2_outputs[172]));
    assign outputs[9875] = (layer2_outputs[2452]) ^ (layer2_outputs[79]);
    assign outputs[9876] = ~(layer2_outputs[7895]);
    assign outputs[9877] = ~((layer2_outputs[2909]) & (layer2_outputs[3138]));
    assign outputs[9878] = ~((layer2_outputs[2225]) ^ (layer2_outputs[5775]));
    assign outputs[9879] = (layer2_outputs[560]) ^ (layer2_outputs[9063]);
    assign outputs[9880] = (layer2_outputs[7951]) & ~(layer2_outputs[7628]);
    assign outputs[9881] = ~(layer2_outputs[7613]);
    assign outputs[9882] = layer2_outputs[6083];
    assign outputs[9883] = ~(layer2_outputs[828]);
    assign outputs[9884] = ~(layer2_outputs[5683]);
    assign outputs[9885] = layer2_outputs[4324];
    assign outputs[9886] = layer2_outputs[5105];
    assign outputs[9887] = ~((layer2_outputs[714]) ^ (layer2_outputs[10237]));
    assign outputs[9888] = layer2_outputs[3686];
    assign outputs[9889] = (layer2_outputs[5064]) ^ (layer2_outputs[1567]);
    assign outputs[9890] = ~(layer2_outputs[2783]);
    assign outputs[9891] = layer2_outputs[10234];
    assign outputs[9892] = (layer2_outputs[2429]) ^ (layer2_outputs[9133]);
    assign outputs[9893] = layer2_outputs[2120];
    assign outputs[9894] = (layer2_outputs[11669]) ^ (layer2_outputs[12203]);
    assign outputs[9895] = layer2_outputs[7526];
    assign outputs[9896] = ~(layer2_outputs[8595]);
    assign outputs[9897] = layer2_outputs[6517];
    assign outputs[9898] = layer2_outputs[108];
    assign outputs[9899] = layer2_outputs[1504];
    assign outputs[9900] = (layer2_outputs[12185]) ^ (layer2_outputs[10831]);
    assign outputs[9901] = ~(layer2_outputs[6360]) | (layer2_outputs[10672]);
    assign outputs[9902] = ~((layer2_outputs[9843]) ^ (layer2_outputs[12073]));
    assign outputs[9903] = layer2_outputs[8886];
    assign outputs[9904] = (layer2_outputs[7114]) | (layer2_outputs[7421]);
    assign outputs[9905] = (layer2_outputs[11701]) ^ (layer2_outputs[7452]);
    assign outputs[9906] = (layer2_outputs[7910]) & ~(layer2_outputs[7106]);
    assign outputs[9907] = ~(layer2_outputs[5581]);
    assign outputs[9908] = (layer2_outputs[619]) ^ (layer2_outputs[9685]);
    assign outputs[9909] = ~((layer2_outputs[4117]) ^ (layer2_outputs[3162]));
    assign outputs[9910] = layer2_outputs[3974];
    assign outputs[9911] = layer2_outputs[11704];
    assign outputs[9912] = ~(layer2_outputs[7255]);
    assign outputs[9913] = layer2_outputs[11257];
    assign outputs[9914] = ~(layer2_outputs[4752]);
    assign outputs[9915] = ~((layer2_outputs[469]) ^ (layer2_outputs[929]));
    assign outputs[9916] = (layer2_outputs[1953]) & (layer2_outputs[7402]);
    assign outputs[9917] = layer2_outputs[7258];
    assign outputs[9918] = ~((layer2_outputs[6202]) ^ (layer2_outputs[12463]));
    assign outputs[9919] = ~(layer2_outputs[4512]);
    assign outputs[9920] = (layer2_outputs[7975]) | (layer2_outputs[4625]);
    assign outputs[9921] = ~(layer2_outputs[8753]);
    assign outputs[9922] = ~(layer2_outputs[8773]);
    assign outputs[9923] = ~(layer2_outputs[9911]);
    assign outputs[9924] = ~(layer2_outputs[7530]);
    assign outputs[9925] = layer2_outputs[9587];
    assign outputs[9926] = layer2_outputs[2741];
    assign outputs[9927] = layer2_outputs[11964];
    assign outputs[9928] = ~(layer2_outputs[6686]);
    assign outputs[9929] = (layer2_outputs[10594]) ^ (layer2_outputs[8778]);
    assign outputs[9930] = ~((layer2_outputs[4439]) | (layer2_outputs[2838]));
    assign outputs[9931] = layer2_outputs[9829];
    assign outputs[9932] = layer2_outputs[7607];
    assign outputs[9933] = layer2_outputs[11400];
    assign outputs[9934] = ~(layer2_outputs[2181]);
    assign outputs[9935] = ~(layer2_outputs[2947]);
    assign outputs[9936] = layer2_outputs[1111];
    assign outputs[9937] = ~((layer2_outputs[9011]) ^ (layer2_outputs[10987]));
    assign outputs[9938] = (layer2_outputs[5868]) ^ (layer2_outputs[10617]);
    assign outputs[9939] = ~((layer2_outputs[1096]) & (layer2_outputs[9408]));
    assign outputs[9940] = ~((layer2_outputs[5409]) ^ (layer2_outputs[7144]));
    assign outputs[9941] = ~(layer2_outputs[6706]) | (layer2_outputs[1844]);
    assign outputs[9942] = (layer2_outputs[11045]) ^ (layer2_outputs[8744]);
    assign outputs[9943] = layer2_outputs[8148];
    assign outputs[9944] = layer2_outputs[9048];
    assign outputs[9945] = layer2_outputs[4032];
    assign outputs[9946] = layer2_outputs[10519];
    assign outputs[9947] = ~(layer2_outputs[3917]);
    assign outputs[9948] = (layer2_outputs[12093]) & (layer2_outputs[10412]);
    assign outputs[9949] = ~((layer2_outputs[5405]) & (layer2_outputs[8900]));
    assign outputs[9950] = ~((layer2_outputs[12730]) ^ (layer2_outputs[3617]));
    assign outputs[9951] = layer2_outputs[8302];
    assign outputs[9952] = ~(layer2_outputs[386]);
    assign outputs[9953] = ~(layer2_outputs[2912]);
    assign outputs[9954] = layer2_outputs[8729];
    assign outputs[9955] = layer2_outputs[12257];
    assign outputs[9956] = ~(layer2_outputs[2300]);
    assign outputs[9957] = layer2_outputs[1074];
    assign outputs[9958] = (layer2_outputs[11523]) ^ (layer2_outputs[261]);
    assign outputs[9959] = layer2_outputs[3188];
    assign outputs[9960] = (layer2_outputs[6393]) & ~(layer2_outputs[2186]);
    assign outputs[9961] = ~((layer2_outputs[7945]) & (layer2_outputs[5884]));
    assign outputs[9962] = ~(layer2_outputs[4601]) | (layer2_outputs[4507]);
    assign outputs[9963] = (layer2_outputs[10266]) ^ (layer2_outputs[6648]);
    assign outputs[9964] = (layer2_outputs[8548]) & ~(layer2_outputs[322]);
    assign outputs[9965] = layer2_outputs[5158];
    assign outputs[9966] = ~(layer2_outputs[12213]);
    assign outputs[9967] = ~(layer2_outputs[7022]);
    assign outputs[9968] = ~((layer2_outputs[10872]) ^ (layer2_outputs[5461]));
    assign outputs[9969] = (layer2_outputs[2289]) & ~(layer2_outputs[8725]);
    assign outputs[9970] = ~(layer2_outputs[8029]);
    assign outputs[9971] = ~((layer2_outputs[11847]) ^ (layer2_outputs[6986]));
    assign outputs[9972] = ~(layer2_outputs[6591]);
    assign outputs[9973] = ~(layer2_outputs[10453]) | (layer2_outputs[12225]);
    assign outputs[9974] = layer2_outputs[10767];
    assign outputs[9975] = layer2_outputs[7588];
    assign outputs[9976] = ~(layer2_outputs[4458]);
    assign outputs[9977] = layer2_outputs[8534];
    assign outputs[9978] = layer2_outputs[5447];
    assign outputs[9979] = ~(layer2_outputs[10815]);
    assign outputs[9980] = ~((layer2_outputs[11360]) ^ (layer2_outputs[9841]));
    assign outputs[9981] = layer2_outputs[275];
    assign outputs[9982] = ~((layer2_outputs[9789]) ^ (layer2_outputs[5776]));
    assign outputs[9983] = (layer2_outputs[5441]) & ~(layer2_outputs[427]);
    assign outputs[9984] = (layer2_outputs[3348]) ^ (layer2_outputs[7270]);
    assign outputs[9985] = ~(layer2_outputs[12030]);
    assign outputs[9986] = ~(layer2_outputs[4727]);
    assign outputs[9987] = ~(layer2_outputs[1879]);
    assign outputs[9988] = ~((layer2_outputs[1592]) ^ (layer2_outputs[11477]));
    assign outputs[9989] = (layer2_outputs[5716]) ^ (layer2_outputs[4091]);
    assign outputs[9990] = layer2_outputs[3197];
    assign outputs[9991] = ~(layer2_outputs[10859]) | (layer2_outputs[11377]);
    assign outputs[9992] = ~((layer2_outputs[10423]) ^ (layer2_outputs[10325]));
    assign outputs[9993] = ~((layer2_outputs[5271]) ^ (layer2_outputs[9878]));
    assign outputs[9994] = layer2_outputs[3095];
    assign outputs[9995] = ~((layer2_outputs[3152]) ^ (layer2_outputs[2574]));
    assign outputs[9996] = ~(layer2_outputs[185]);
    assign outputs[9997] = ~(layer2_outputs[10997]);
    assign outputs[9998] = layer2_outputs[4798];
    assign outputs[9999] = ~(layer2_outputs[8004]);
    assign outputs[10000] = layer2_outputs[8127];
    assign outputs[10001] = (layer2_outputs[772]) ^ (layer2_outputs[4094]);
    assign outputs[10002] = (layer2_outputs[10153]) ^ (layer2_outputs[10856]);
    assign outputs[10003] = ~((layer2_outputs[6530]) ^ (layer2_outputs[11836]));
    assign outputs[10004] = ~(layer2_outputs[4394]);
    assign outputs[10005] = layer2_outputs[7773];
    assign outputs[10006] = ~(layer2_outputs[5730]);
    assign outputs[10007] = (layer2_outputs[5918]) ^ (layer2_outputs[11839]);
    assign outputs[10008] = ~(layer2_outputs[7119]);
    assign outputs[10009] = (layer2_outputs[12110]) & ~(layer2_outputs[3518]);
    assign outputs[10010] = layer2_outputs[10647];
    assign outputs[10011] = ~(layer2_outputs[12027]);
    assign outputs[10012] = (layer2_outputs[11673]) & ~(layer2_outputs[10904]);
    assign outputs[10013] = (layer2_outputs[10041]) ^ (layer2_outputs[5217]);
    assign outputs[10014] = ~(layer2_outputs[7728]);
    assign outputs[10015] = (layer2_outputs[1757]) ^ (layer2_outputs[9330]);
    assign outputs[10016] = layer2_outputs[5694];
    assign outputs[10017] = layer2_outputs[6289];
    assign outputs[10018] = layer2_outputs[4696];
    assign outputs[10019] = ~(layer2_outputs[7572]);
    assign outputs[10020] = ~((layer2_outputs[4883]) ^ (layer2_outputs[9098]));
    assign outputs[10021] = (layer2_outputs[12653]) ^ (layer2_outputs[11618]);
    assign outputs[10022] = ~(layer2_outputs[9918]);
    assign outputs[10023] = ~(layer2_outputs[9086]);
    assign outputs[10024] = ~(layer2_outputs[4418]);
    assign outputs[10025] = ~(layer2_outputs[11789]);
    assign outputs[10026] = ~((layer2_outputs[9323]) ^ (layer2_outputs[6462]));
    assign outputs[10027] = (layer2_outputs[9989]) ^ (layer2_outputs[6550]);
    assign outputs[10028] = ~(layer2_outputs[2935]);
    assign outputs[10029] = (layer2_outputs[4385]) & ~(layer2_outputs[4805]);
    assign outputs[10030] = (layer2_outputs[9001]) | (layer2_outputs[12229]);
    assign outputs[10031] = (layer2_outputs[8692]) ^ (layer2_outputs[4344]);
    assign outputs[10032] = layer2_outputs[7830];
    assign outputs[10033] = ~(layer2_outputs[10249]);
    assign outputs[10034] = ~(layer2_outputs[9188]);
    assign outputs[10035] = (layer2_outputs[5781]) ^ (layer2_outputs[8689]);
    assign outputs[10036] = ~((layer2_outputs[1987]) ^ (layer2_outputs[2701]));
    assign outputs[10037] = ~(layer2_outputs[4267]) | (layer2_outputs[4255]);
    assign outputs[10038] = ~((layer2_outputs[8593]) ^ (layer2_outputs[2835]));
    assign outputs[10039] = ~(layer2_outputs[4656]);
    assign outputs[10040] = ~(layer2_outputs[2723]);
    assign outputs[10041] = ~(layer2_outputs[5088]);
    assign outputs[10042] = layer2_outputs[11083];
    assign outputs[10043] = layer2_outputs[9164];
    assign outputs[10044] = ~((layer2_outputs[12334]) ^ (layer2_outputs[6159]));
    assign outputs[10045] = ~((layer2_outputs[2618]) ^ (layer2_outputs[9799]));
    assign outputs[10046] = ~((layer2_outputs[12076]) ^ (layer2_outputs[2740]));
    assign outputs[10047] = ~((layer2_outputs[6868]) | (layer2_outputs[6813]));
    assign outputs[10048] = ~(layer2_outputs[3416]);
    assign outputs[10049] = ~((layer2_outputs[11582]) ^ (layer2_outputs[466]));
    assign outputs[10050] = ~(layer2_outputs[87]);
    assign outputs[10051] = layer2_outputs[6254];
    assign outputs[10052] = layer2_outputs[1205];
    assign outputs[10053] = layer2_outputs[8653];
    assign outputs[10054] = (layer2_outputs[12538]) ^ (layer2_outputs[8225]);
    assign outputs[10055] = (layer2_outputs[6906]) & ~(layer2_outputs[10459]);
    assign outputs[10056] = layer2_outputs[7757];
    assign outputs[10057] = layer2_outputs[3915];
    assign outputs[10058] = ~(layer2_outputs[4527]);
    assign outputs[10059] = layer2_outputs[572];
    assign outputs[10060] = (layer2_outputs[292]) & ~(layer2_outputs[10177]);
    assign outputs[10061] = ~(layer2_outputs[5743]);
    assign outputs[10062] = layer2_outputs[6434];
    assign outputs[10063] = (layer2_outputs[8150]) & ~(layer2_outputs[6600]);
    assign outputs[10064] = ~((layer2_outputs[1696]) | (layer2_outputs[10435]));
    assign outputs[10065] = ~((layer2_outputs[11374]) & (layer2_outputs[750]));
    assign outputs[10066] = ~(layer2_outputs[6839]) | (layer2_outputs[1111]);
    assign outputs[10067] = (layer2_outputs[5272]) ^ (layer2_outputs[6433]);
    assign outputs[10068] = layer2_outputs[424];
    assign outputs[10069] = layer2_outputs[10035];
    assign outputs[10070] = ~((layer2_outputs[7603]) | (layer2_outputs[11492]));
    assign outputs[10071] = layer2_outputs[791];
    assign outputs[10072] = layer2_outputs[4369];
    assign outputs[10073] = ~(layer2_outputs[5445]);
    assign outputs[10074] = ~(layer2_outputs[4712]);
    assign outputs[10075] = layer2_outputs[4788];
    assign outputs[10076] = (layer2_outputs[1465]) & (layer2_outputs[9204]);
    assign outputs[10077] = ~(layer2_outputs[9652]);
    assign outputs[10078] = ~((layer2_outputs[1289]) ^ (layer2_outputs[5223]));
    assign outputs[10079] = layer2_outputs[4197];
    assign outputs[10080] = ~(layer2_outputs[6519]);
    assign outputs[10081] = layer2_outputs[9245];
    assign outputs[10082] = layer2_outputs[8439];
    assign outputs[10083] = layer2_outputs[12101];
    assign outputs[10084] = layer2_outputs[4041];
    assign outputs[10085] = ~(layer2_outputs[9548]);
    assign outputs[10086] = (layer2_outputs[12523]) & ~(layer2_outputs[119]);
    assign outputs[10087] = ~((layer2_outputs[2534]) ^ (layer2_outputs[11580]));
    assign outputs[10088] = ~(layer2_outputs[8325]);
    assign outputs[10089] = (layer2_outputs[9685]) ^ (layer2_outputs[6130]);
    assign outputs[10090] = layer2_outputs[6311];
    assign outputs[10091] = (layer2_outputs[8521]) & ~(layer2_outputs[5311]);
    assign outputs[10092] = ~((layer2_outputs[10126]) ^ (layer2_outputs[8247]));
    assign outputs[10093] = (layer2_outputs[290]) ^ (layer2_outputs[357]);
    assign outputs[10094] = ~(layer2_outputs[1530]);
    assign outputs[10095] = ~(layer2_outputs[10702]);
    assign outputs[10096] = ~(layer2_outputs[6905]);
    assign outputs[10097] = (layer2_outputs[9448]) ^ (layer2_outputs[1749]);
    assign outputs[10098] = ~(layer2_outputs[5389]);
    assign outputs[10099] = layer2_outputs[10645];
    assign outputs[10100] = ~((layer2_outputs[3953]) ^ (layer2_outputs[1910]));
    assign outputs[10101] = ~(layer2_outputs[1381]);
    assign outputs[10102] = ~(layer2_outputs[5593]);
    assign outputs[10103] = (layer2_outputs[12517]) & ~(layer2_outputs[8152]);
    assign outputs[10104] = layer2_outputs[1097];
    assign outputs[10105] = layer2_outputs[12140];
    assign outputs[10106] = ~(layer2_outputs[9271]) | (layer2_outputs[4618]);
    assign outputs[10107] = (layer2_outputs[7584]) & (layer2_outputs[10354]);
    assign outputs[10108] = layer2_outputs[9342];
    assign outputs[10109] = layer2_outputs[2937];
    assign outputs[10110] = (layer2_outputs[7680]) ^ (layer2_outputs[10333]);
    assign outputs[10111] = ~(layer2_outputs[1531]);
    assign outputs[10112] = layer2_outputs[4009];
    assign outputs[10113] = ~(layer2_outputs[5387]);
    assign outputs[10114] = ~(layer2_outputs[5549]);
    assign outputs[10115] = ~(layer2_outputs[9573]);
    assign outputs[10116] = ~(layer2_outputs[7387]);
    assign outputs[10117] = ~(layer2_outputs[10198]);
    assign outputs[10118] = layer2_outputs[11774];
    assign outputs[10119] = layer2_outputs[7998];
    assign outputs[10120] = layer2_outputs[6066];
    assign outputs[10121] = (layer2_outputs[5303]) & ~(layer2_outputs[6582]);
    assign outputs[10122] = ~(layer2_outputs[5128]);
    assign outputs[10123] = (layer2_outputs[8801]) | (layer2_outputs[9477]);
    assign outputs[10124] = ~((layer2_outputs[8246]) & (layer2_outputs[12591]));
    assign outputs[10125] = layer2_outputs[9324];
    assign outputs[10126] = (layer2_outputs[3214]) ^ (layer2_outputs[9734]);
    assign outputs[10127] = layer2_outputs[642];
    assign outputs[10128] = ~((layer2_outputs[1774]) ^ (layer2_outputs[10502]));
    assign outputs[10129] = ~(layer2_outputs[12335]);
    assign outputs[10130] = ~(layer2_outputs[6026]);
    assign outputs[10131] = ~((layer2_outputs[9867]) | (layer2_outputs[3]));
    assign outputs[10132] = (layer2_outputs[2363]) & ~(layer2_outputs[1365]);
    assign outputs[10133] = (layer2_outputs[8127]) ^ (layer2_outputs[1423]);
    assign outputs[10134] = layer2_outputs[5641];
    assign outputs[10135] = ~(layer2_outputs[10625]) | (layer2_outputs[11519]);
    assign outputs[10136] = (layer2_outputs[10573]) ^ (layer2_outputs[11219]);
    assign outputs[10137] = (layer2_outputs[10544]) ^ (layer2_outputs[10016]);
    assign outputs[10138] = ~(layer2_outputs[5908]);
    assign outputs[10139] = layer2_outputs[8440];
    assign outputs[10140] = ~(layer2_outputs[12290]);
    assign outputs[10141] = ~((layer2_outputs[10914]) ^ (layer2_outputs[1775]));
    assign outputs[10142] = ~(layer2_outputs[460]);
    assign outputs[10143] = layer2_outputs[11207];
    assign outputs[10144] = (layer2_outputs[9939]) ^ (layer2_outputs[1789]);
    assign outputs[10145] = ~(layer2_outputs[8884]);
    assign outputs[10146] = (layer2_outputs[8544]) ^ (layer2_outputs[12071]);
    assign outputs[10147] = (layer2_outputs[10620]) & ~(layer2_outputs[528]);
    assign outputs[10148] = ~(layer2_outputs[4501]) | (layer2_outputs[331]);
    assign outputs[10149] = ~(layer2_outputs[11824]);
    assign outputs[10150] = ~((layer2_outputs[11496]) ^ (layer2_outputs[7088]));
    assign outputs[10151] = layer2_outputs[2511];
    assign outputs[10152] = layer2_outputs[2833];
    assign outputs[10153] = ~(layer2_outputs[941]);
    assign outputs[10154] = ~(layer2_outputs[8724]);
    assign outputs[10155] = (layer2_outputs[2787]) ^ (layer2_outputs[9641]);
    assign outputs[10156] = ~((layer2_outputs[9037]) ^ (layer2_outputs[7565]));
    assign outputs[10157] = ~((layer2_outputs[9415]) ^ (layer2_outputs[9783]));
    assign outputs[10158] = ~((layer2_outputs[3623]) ^ (layer2_outputs[4834]));
    assign outputs[10159] = ~((layer2_outputs[4928]) & (layer2_outputs[7717]));
    assign outputs[10160] = layer2_outputs[4385];
    assign outputs[10161] = (layer2_outputs[3802]) & (layer2_outputs[5542]);
    assign outputs[10162] = layer2_outputs[11631];
    assign outputs[10163] = ~(layer2_outputs[9561]);
    assign outputs[10164] = ~((layer2_outputs[5167]) ^ (layer2_outputs[10294]));
    assign outputs[10165] = ~((layer2_outputs[1665]) | (layer2_outputs[6323]));
    assign outputs[10166] = layer2_outputs[1227];
    assign outputs[10167] = (layer2_outputs[11957]) & (layer2_outputs[469]);
    assign outputs[10168] = ~(layer2_outputs[5981]);
    assign outputs[10169] = ~((layer2_outputs[1922]) ^ (layer2_outputs[3300]));
    assign outputs[10170] = (layer2_outputs[5903]) ^ (layer2_outputs[2097]);
    assign outputs[10171] = ~(layer2_outputs[7598]);
    assign outputs[10172] = layer2_outputs[4488];
    assign outputs[10173] = layer2_outputs[3533];
    assign outputs[10174] = layer2_outputs[1095];
    assign outputs[10175] = layer2_outputs[6602];
    assign outputs[10176] = ~(layer2_outputs[151]);
    assign outputs[10177] = layer2_outputs[3973];
    assign outputs[10178] = ~((layer2_outputs[1277]) | (layer2_outputs[9015]));
    assign outputs[10179] = (layer2_outputs[1916]) & (layer2_outputs[5711]);
    assign outputs[10180] = ~(layer2_outputs[3410]) | (layer2_outputs[4636]);
    assign outputs[10181] = layer2_outputs[12718];
    assign outputs[10182] = layer2_outputs[8159];
    assign outputs[10183] = ~((layer2_outputs[10973]) ^ (layer2_outputs[8536]));
    assign outputs[10184] = layer2_outputs[7024];
    assign outputs[10185] = ~(layer2_outputs[1578]);
    assign outputs[10186] = ~(layer2_outputs[4389]);
    assign outputs[10187] = layer2_outputs[1169];
    assign outputs[10188] = layer2_outputs[1227];
    assign outputs[10189] = layer2_outputs[11330];
    assign outputs[10190] = layer2_outputs[4208];
    assign outputs[10191] = layer2_outputs[9769];
    assign outputs[10192] = layer2_outputs[11798];
    assign outputs[10193] = layer2_outputs[8414];
    assign outputs[10194] = ~(layer2_outputs[12622]);
    assign outputs[10195] = ~(layer2_outputs[2031]);
    assign outputs[10196] = ~((layer2_outputs[10490]) | (layer2_outputs[6607]));
    assign outputs[10197] = ~(layer2_outputs[2771]);
    assign outputs[10198] = ~((layer2_outputs[9928]) ^ (layer2_outputs[8690]));
    assign outputs[10199] = ~(layer2_outputs[1614]);
    assign outputs[10200] = ~(layer2_outputs[9433]);
    assign outputs[10201] = (layer2_outputs[12409]) ^ (layer2_outputs[12687]);
    assign outputs[10202] = layer2_outputs[3637];
    assign outputs[10203] = layer2_outputs[2836];
    assign outputs[10204] = ~(layer2_outputs[2539]) | (layer2_outputs[2348]);
    assign outputs[10205] = layer2_outputs[9246];
    assign outputs[10206] = ~(layer2_outputs[763]);
    assign outputs[10207] = ~(layer2_outputs[9338]);
    assign outputs[10208] = layer2_outputs[7564];
    assign outputs[10209] = (layer2_outputs[10442]) & ~(layer2_outputs[7701]);
    assign outputs[10210] = (layer2_outputs[11897]) | (layer2_outputs[2448]);
    assign outputs[10211] = layer2_outputs[8726];
    assign outputs[10212] = ~(layer2_outputs[5740]);
    assign outputs[10213] = layer2_outputs[8363];
    assign outputs[10214] = layer2_outputs[2477];
    assign outputs[10215] = ~((layer2_outputs[11358]) | (layer2_outputs[8221]));
    assign outputs[10216] = (layer2_outputs[8593]) ^ (layer2_outputs[9023]);
    assign outputs[10217] = (layer2_outputs[10356]) & (layer2_outputs[11398]);
    assign outputs[10218] = (layer2_outputs[9743]) & ~(layer2_outputs[1685]);
    assign outputs[10219] = ~(layer2_outputs[314]);
    assign outputs[10220] = ~(layer2_outputs[2117]);
    assign outputs[10221] = ~(layer2_outputs[3874]);
    assign outputs[10222] = (layer2_outputs[10390]) & ~(layer2_outputs[7423]);
    assign outputs[10223] = ~(layer2_outputs[8583]);
    assign outputs[10224] = ~((layer2_outputs[8781]) ^ (layer2_outputs[6855]));
    assign outputs[10225] = (layer2_outputs[1105]) ^ (layer2_outputs[3406]);
    assign outputs[10226] = (layer2_outputs[3794]) ^ (layer2_outputs[2388]);
    assign outputs[10227] = ~((layer2_outputs[6244]) ^ (layer2_outputs[5979]));
    assign outputs[10228] = layer2_outputs[7062];
    assign outputs[10229] = layer2_outputs[81];
    assign outputs[10230] = ~(layer2_outputs[5353]);
    assign outputs[10231] = ~(layer2_outputs[3642]);
    assign outputs[10232] = (layer2_outputs[902]) ^ (layer2_outputs[1395]);
    assign outputs[10233] = layer2_outputs[8082];
    assign outputs[10234] = ~(layer2_outputs[2911]);
    assign outputs[10235] = ~((layer2_outputs[4176]) ^ (layer2_outputs[7743]));
    assign outputs[10236] = layer2_outputs[5070];
    assign outputs[10237] = ~(layer2_outputs[3198]);
    assign outputs[10238] = (layer2_outputs[11575]) ^ (layer2_outputs[793]);
    assign outputs[10239] = ~(layer2_outputs[4129]);
    assign outputs[10240] = layer2_outputs[9755];
    assign outputs[10241] = (layer2_outputs[6815]) | (layer2_outputs[10147]);
    assign outputs[10242] = layer2_outputs[10117];
    assign outputs[10243] = ~((layer2_outputs[11370]) ^ (layer2_outputs[11391]));
    assign outputs[10244] = layer2_outputs[10540];
    assign outputs[10245] = layer2_outputs[10614];
    assign outputs[10246] = ~(layer2_outputs[7147]);
    assign outputs[10247] = ~(layer2_outputs[4701]) | (layer2_outputs[10353]);
    assign outputs[10248] = ~(layer2_outputs[11030]);
    assign outputs[10249] = (layer2_outputs[4163]) & (layer2_outputs[9006]);
    assign outputs[10250] = ~(layer2_outputs[682]);
    assign outputs[10251] = (layer2_outputs[3700]) ^ (layer2_outputs[12230]);
    assign outputs[10252] = layer2_outputs[522];
    assign outputs[10253] = ~(layer2_outputs[12239]) | (layer2_outputs[10725]);
    assign outputs[10254] = ~((layer2_outputs[1404]) ^ (layer2_outputs[6135]));
    assign outputs[10255] = ~(layer2_outputs[6769]);
    assign outputs[10256] = (layer2_outputs[10819]) ^ (layer2_outputs[1700]);
    assign outputs[10257] = ~((layer2_outputs[3911]) ^ (layer2_outputs[3098]));
    assign outputs[10258] = ~(layer2_outputs[1353]);
    assign outputs[10259] = ~(layer2_outputs[8658]);
    assign outputs[10260] = (layer2_outputs[6506]) ^ (layer2_outputs[6770]);
    assign outputs[10261] = (layer2_outputs[1609]) ^ (layer2_outputs[3364]);
    assign outputs[10262] = layer2_outputs[8992];
    assign outputs[10263] = (layer2_outputs[947]) | (layer2_outputs[1309]);
    assign outputs[10264] = (layer2_outputs[9682]) ^ (layer2_outputs[2058]);
    assign outputs[10265] = ~(layer2_outputs[1005]);
    assign outputs[10266] = layer2_outputs[11243];
    assign outputs[10267] = layer2_outputs[4153];
    assign outputs[10268] = ~(layer2_outputs[4456]);
    assign outputs[10269] = ~(layer2_outputs[1568]);
    assign outputs[10270] = (layer2_outputs[3857]) & (layer2_outputs[7095]);
    assign outputs[10271] = layer2_outputs[12314];
    assign outputs[10272] = ~(layer2_outputs[5080]) | (layer2_outputs[10631]);
    assign outputs[10273] = ~(layer2_outputs[3694]) | (layer2_outputs[527]);
    assign outputs[10274] = (layer2_outputs[9570]) ^ (layer2_outputs[9811]);
    assign outputs[10275] = (layer2_outputs[2362]) ^ (layer2_outputs[4584]);
    assign outputs[10276] = layer2_outputs[9223];
    assign outputs[10277] = ~(layer2_outputs[7690]);
    assign outputs[10278] = (layer2_outputs[4889]) ^ (layer2_outputs[12793]);
    assign outputs[10279] = ~((layer2_outputs[487]) ^ (layer2_outputs[8606]));
    assign outputs[10280] = layer2_outputs[10374];
    assign outputs[10281] = ~(layer2_outputs[3191]);
    assign outputs[10282] = ~((layer2_outputs[12129]) ^ (layer2_outputs[4488]));
    assign outputs[10283] = ~(layer2_outputs[11177]);
    assign outputs[10284] = layer2_outputs[9187];
    assign outputs[10285] = (layer2_outputs[2949]) & ~(layer2_outputs[8964]);
    assign outputs[10286] = ~((layer2_outputs[377]) ^ (layer2_outputs[2178]));
    assign outputs[10287] = ~(layer2_outputs[3737]);
    assign outputs[10288] = (layer2_outputs[5716]) ^ (layer2_outputs[2100]);
    assign outputs[10289] = ~(layer2_outputs[4606]);
    assign outputs[10290] = layer2_outputs[7507];
    assign outputs[10291] = layer2_outputs[3248];
    assign outputs[10292] = layer2_outputs[11001];
    assign outputs[10293] = ~((layer2_outputs[10305]) ^ (layer2_outputs[10509]));
    assign outputs[10294] = (layer2_outputs[9292]) ^ (layer2_outputs[12116]);
    assign outputs[10295] = (layer2_outputs[3340]) ^ (layer2_outputs[8655]);
    assign outputs[10296] = (layer2_outputs[4422]) ^ (layer2_outputs[7228]);
    assign outputs[10297] = layer2_outputs[12625];
    assign outputs[10298] = ~(layer2_outputs[11553]);
    assign outputs[10299] = layer2_outputs[1779];
    assign outputs[10300] = ~((layer2_outputs[12345]) ^ (layer2_outputs[8792]));
    assign outputs[10301] = layer2_outputs[5817];
    assign outputs[10302] = layer2_outputs[6283];
    assign outputs[10303] = ~(layer2_outputs[1014]);
    assign outputs[10304] = ~(layer2_outputs[9845]);
    assign outputs[10305] = ~(layer2_outputs[7419]);
    assign outputs[10306] = (layer2_outputs[11604]) ^ (layer2_outputs[1132]);
    assign outputs[10307] = ~(layer2_outputs[5535]);
    assign outputs[10308] = layer2_outputs[12788];
    assign outputs[10309] = ~((layer2_outputs[168]) ^ (layer2_outputs[10303]));
    assign outputs[10310] = ~(layer2_outputs[3147]);
    assign outputs[10311] = ~(layer2_outputs[5836]);
    assign outputs[10312] = layer2_outputs[9747];
    assign outputs[10313] = layer2_outputs[195];
    assign outputs[10314] = ~(layer2_outputs[5362]);
    assign outputs[10315] = ~(layer2_outputs[5131]);
    assign outputs[10316] = ~(layer2_outputs[10255]);
    assign outputs[10317] = layer2_outputs[12215];
    assign outputs[10318] = ~((layer2_outputs[4862]) | (layer2_outputs[4696]));
    assign outputs[10319] = layer2_outputs[1436];
    assign outputs[10320] = (layer2_outputs[10449]) | (layer2_outputs[434]);
    assign outputs[10321] = ~(layer2_outputs[8964]) | (layer2_outputs[5400]);
    assign outputs[10322] = ~((layer2_outputs[8064]) ^ (layer2_outputs[1951]));
    assign outputs[10323] = ~(layer2_outputs[919]);
    assign outputs[10324] = (layer2_outputs[6044]) ^ (layer2_outputs[11319]);
    assign outputs[10325] = ~((layer2_outputs[11772]) ^ (layer2_outputs[10854]));
    assign outputs[10326] = ~((layer2_outputs[8109]) ^ (layer2_outputs[1496]));
    assign outputs[10327] = ~((layer2_outputs[12432]) ^ (layer2_outputs[7233]));
    assign outputs[10328] = (layer2_outputs[8128]) ^ (layer2_outputs[9243]);
    assign outputs[10329] = ~(layer2_outputs[2433]) | (layer2_outputs[6120]);
    assign outputs[10330] = (layer2_outputs[12601]) ^ (layer2_outputs[5088]);
    assign outputs[10331] = ~(layer2_outputs[8708]);
    assign outputs[10332] = ~(layer2_outputs[8631]) | (layer2_outputs[468]);
    assign outputs[10333] = (layer2_outputs[4352]) ^ (layer2_outputs[10243]);
    assign outputs[10334] = layer2_outputs[6359];
    assign outputs[10335] = layer2_outputs[12728];
    assign outputs[10336] = ~((layer2_outputs[3465]) ^ (layer2_outputs[10411]));
    assign outputs[10337] = (layer2_outputs[173]) & ~(layer2_outputs[9447]);
    assign outputs[10338] = (layer2_outputs[1836]) ^ (layer2_outputs[5287]);
    assign outputs[10339] = layer2_outputs[10351];
    assign outputs[10340] = ~(layer2_outputs[11293]);
    assign outputs[10341] = layer2_outputs[1669];
    assign outputs[10342] = ~(layer2_outputs[11690]) | (layer2_outputs[5976]);
    assign outputs[10343] = ~(layer2_outputs[6313]);
    assign outputs[10344] = layer2_outputs[2008];
    assign outputs[10345] = ~(layer2_outputs[10511]);
    assign outputs[10346] = layer2_outputs[4128];
    assign outputs[10347] = ~((layer2_outputs[1326]) ^ (layer2_outputs[4471]));
    assign outputs[10348] = ~(layer2_outputs[5138]);
    assign outputs[10349] = (layer2_outputs[10245]) ^ (layer2_outputs[9146]);
    assign outputs[10350] = ~((layer2_outputs[3044]) & (layer2_outputs[7903]));
    assign outputs[10351] = ~((layer2_outputs[8744]) ^ (layer2_outputs[12366]));
    assign outputs[10352] = ~(layer2_outputs[8438]);
    assign outputs[10353] = ~(layer2_outputs[6585]) | (layer2_outputs[10898]);
    assign outputs[10354] = ~(layer2_outputs[10313]) | (layer2_outputs[686]);
    assign outputs[10355] = ~(layer2_outputs[5481]);
    assign outputs[10356] = ~((layer2_outputs[4892]) ^ (layer2_outputs[10628]));
    assign outputs[10357] = ~(layer2_outputs[4645]);
    assign outputs[10358] = layer2_outputs[9550];
    assign outputs[10359] = layer2_outputs[12193];
    assign outputs[10360] = ~((layer2_outputs[1348]) ^ (layer2_outputs[2008]));
    assign outputs[10361] = ~(layer2_outputs[4331]);
    assign outputs[10362] = ~(layer2_outputs[6954]);
    assign outputs[10363] = layer2_outputs[2748];
    assign outputs[10364] = ~(layer2_outputs[2109]);
    assign outputs[10365] = (layer2_outputs[8634]) ^ (layer2_outputs[11352]);
    assign outputs[10366] = layer2_outputs[8552];
    assign outputs[10367] = layer2_outputs[280];
    assign outputs[10368] = ~((layer2_outputs[4022]) ^ (layer2_outputs[10417]));
    assign outputs[10369] = ~(layer2_outputs[9134]) | (layer2_outputs[4634]);
    assign outputs[10370] = (layer2_outputs[8461]) ^ (layer2_outputs[3299]);
    assign outputs[10371] = (layer2_outputs[9123]) ^ (layer2_outputs[7214]);
    assign outputs[10372] = layer2_outputs[4442];
    assign outputs[10373] = layer2_outputs[2196];
    assign outputs[10374] = ~(layer2_outputs[11681]);
    assign outputs[10375] = ~(layer2_outputs[3066]) | (layer2_outputs[10776]);
    assign outputs[10376] = ~(layer2_outputs[2904]);
    assign outputs[10377] = layer2_outputs[11877];
    assign outputs[10378] = ~((layer2_outputs[9433]) ^ (layer2_outputs[10790]));
    assign outputs[10379] = layer2_outputs[4277];
    assign outputs[10380] = ~(layer2_outputs[12065]);
    assign outputs[10381] = ~(layer2_outputs[7966]);
    assign outputs[10382] = (layer2_outputs[7176]) ^ (layer2_outputs[11504]);
    assign outputs[10383] = ~((layer2_outputs[5301]) | (layer2_outputs[5875]));
    assign outputs[10384] = ~(layer2_outputs[6525]);
    assign outputs[10385] = layer2_outputs[8901];
    assign outputs[10386] = ~((layer2_outputs[9143]) ^ (layer2_outputs[6699]));
    assign outputs[10387] = ~((layer2_outputs[4734]) ^ (layer2_outputs[210]));
    assign outputs[10388] = (layer2_outputs[2549]) ^ (layer2_outputs[1827]);
    assign outputs[10389] = ~(layer2_outputs[9214]) | (layer2_outputs[10510]);
    assign outputs[10390] = (layer2_outputs[4659]) & ~(layer2_outputs[11551]);
    assign outputs[10391] = ~(layer2_outputs[433]);
    assign outputs[10392] = (layer2_outputs[2030]) ^ (layer2_outputs[2772]);
    assign outputs[10393] = (layer2_outputs[1389]) & ~(layer2_outputs[1284]);
    assign outputs[10394] = layer2_outputs[9228];
    assign outputs[10395] = ~((layer2_outputs[10179]) ^ (layer2_outputs[9445]));
    assign outputs[10396] = ~(layer2_outputs[1155]);
    assign outputs[10397] = ~((layer2_outputs[6117]) | (layer2_outputs[8522]));
    assign outputs[10398] = ~(layer2_outputs[4468]) | (layer2_outputs[5724]);
    assign outputs[10399] = ~(layer2_outputs[8515]);
    assign outputs[10400] = ~(layer2_outputs[6422]);
    assign outputs[10401] = layer2_outputs[6076];
    assign outputs[10402] = (layer2_outputs[12735]) | (layer2_outputs[3034]);
    assign outputs[10403] = ~(layer2_outputs[6004]) | (layer2_outputs[12034]);
    assign outputs[10404] = (layer2_outputs[10281]) | (layer2_outputs[12575]);
    assign outputs[10405] = layer2_outputs[6229];
    assign outputs[10406] = ~(layer2_outputs[585]);
    assign outputs[10407] = (layer2_outputs[4189]) & (layer2_outputs[9854]);
    assign outputs[10408] = ~((layer2_outputs[10194]) ^ (layer2_outputs[7406]));
    assign outputs[10409] = ~(layer2_outputs[1963]);
    assign outputs[10410] = ~(layer2_outputs[6846]);
    assign outputs[10411] = ~(layer2_outputs[10149]) | (layer2_outputs[10607]);
    assign outputs[10412] = (layer2_outputs[8340]) ^ (layer2_outputs[3329]);
    assign outputs[10413] = layer2_outputs[10056];
    assign outputs[10414] = layer2_outputs[2640];
    assign outputs[10415] = (layer2_outputs[7657]) ^ (layer2_outputs[2817]);
    assign outputs[10416] = (layer2_outputs[1656]) | (layer2_outputs[4908]);
    assign outputs[10417] = ~((layer2_outputs[12709]) ^ (layer2_outputs[11407]));
    assign outputs[10418] = ~(layer2_outputs[8797]) | (layer2_outputs[12601]);
    assign outputs[10419] = ~(layer2_outputs[12433]);
    assign outputs[10420] = ~(layer2_outputs[10709]);
    assign outputs[10421] = layer2_outputs[1547];
    assign outputs[10422] = ~(layer2_outputs[1118]) | (layer2_outputs[7208]);
    assign outputs[10423] = ~((layer2_outputs[4158]) ^ (layer2_outputs[8031]));
    assign outputs[10424] = (layer2_outputs[462]) ^ (layer2_outputs[8559]);
    assign outputs[10425] = layer2_outputs[3316];
    assign outputs[10426] = (layer2_outputs[4922]) | (layer2_outputs[6929]);
    assign outputs[10427] = layer2_outputs[7085];
    assign outputs[10428] = layer2_outputs[3981];
    assign outputs[10429] = layer2_outputs[10508];
    assign outputs[10430] = (layer2_outputs[12441]) ^ (layer2_outputs[10214]);
    assign outputs[10431] = ~((layer2_outputs[12557]) ^ (layer2_outputs[11337]));
    assign outputs[10432] = (layer2_outputs[9089]) | (layer2_outputs[10850]);
    assign outputs[10433] = ~(layer2_outputs[5050]);
    assign outputs[10434] = (layer2_outputs[7730]) ^ (layer2_outputs[753]);
    assign outputs[10435] = layer2_outputs[1710];
    assign outputs[10436] = ~(layer2_outputs[9008]) | (layer2_outputs[1329]);
    assign outputs[10437] = ~(layer2_outputs[177]);
    assign outputs[10438] = layer2_outputs[6258];
    assign outputs[10439] = (layer2_outputs[9328]) ^ (layer2_outputs[6740]);
    assign outputs[10440] = (layer2_outputs[1999]) ^ (layer2_outputs[12778]);
    assign outputs[10441] = (layer2_outputs[3825]) ^ (layer2_outputs[2999]);
    assign outputs[10442] = ~((layer2_outputs[8277]) ^ (layer2_outputs[960]));
    assign outputs[10443] = (layer2_outputs[8561]) ^ (layer2_outputs[3926]);
    assign outputs[10444] = (layer2_outputs[1980]) ^ (layer2_outputs[4008]);
    assign outputs[10445] = ~((layer2_outputs[2868]) ^ (layer2_outputs[5051]));
    assign outputs[10446] = layer2_outputs[13];
    assign outputs[10447] = ~(layer2_outputs[8874]) | (layer2_outputs[5285]);
    assign outputs[10448] = ~(layer2_outputs[11883]) | (layer2_outputs[597]);
    assign outputs[10449] = (layer2_outputs[4733]) ^ (layer2_outputs[10275]);
    assign outputs[10450] = (layer2_outputs[4408]) ^ (layer2_outputs[1765]);
    assign outputs[10451] = (layer2_outputs[3811]) ^ (layer2_outputs[4142]);
    assign outputs[10452] = ~(layer2_outputs[12283]) | (layer2_outputs[6061]);
    assign outputs[10453] = (layer2_outputs[11449]) & ~(layer2_outputs[8513]);
    assign outputs[10454] = (layer2_outputs[4290]) ^ (layer2_outputs[8028]);
    assign outputs[10455] = (layer2_outputs[11387]) ^ (layer2_outputs[7931]);
    assign outputs[10456] = ~(layer2_outputs[6474]);
    assign outputs[10457] = ~((layer2_outputs[7732]) ^ (layer2_outputs[10083]));
    assign outputs[10458] = layer2_outputs[9250];
    assign outputs[10459] = layer2_outputs[510];
    assign outputs[10460] = ~((layer2_outputs[3983]) ^ (layer2_outputs[11497]));
    assign outputs[10461] = layer2_outputs[9871];
    assign outputs[10462] = (layer2_outputs[3874]) ^ (layer2_outputs[8012]);
    assign outputs[10463] = ~(layer2_outputs[9751]) | (layer2_outputs[2990]);
    assign outputs[10464] = ~((layer2_outputs[3046]) ^ (layer2_outputs[1777]));
    assign outputs[10465] = (layer2_outputs[3940]) ^ (layer2_outputs[873]);
    assign outputs[10466] = ~(layer2_outputs[8164]);
    assign outputs[10467] = (layer2_outputs[7743]) ^ (layer2_outputs[10085]);
    assign outputs[10468] = ~(layer2_outputs[11682]);
    assign outputs[10469] = (layer2_outputs[238]) & ~(layer2_outputs[1026]);
    assign outputs[10470] = layer2_outputs[2604];
    assign outputs[10471] = ~(layer2_outputs[6006]) | (layer2_outputs[7348]);
    assign outputs[10472] = layer2_outputs[11803];
    assign outputs[10473] = (layer2_outputs[3914]) ^ (layer2_outputs[10512]);
    assign outputs[10474] = layer2_outputs[10576];
    assign outputs[10475] = (layer2_outputs[2276]) ^ (layer2_outputs[2592]);
    assign outputs[10476] = ~((layer2_outputs[4634]) ^ (layer2_outputs[11323]));
    assign outputs[10477] = ~((layer2_outputs[7051]) & (layer2_outputs[11845]));
    assign outputs[10478] = layer2_outputs[11487];
    assign outputs[10479] = layer2_outputs[5713];
    assign outputs[10480] = (layer2_outputs[1163]) ^ (layer2_outputs[10281]);
    assign outputs[10481] = layer2_outputs[477];
    assign outputs[10482] = layer2_outputs[9031];
    assign outputs[10483] = ~(layer2_outputs[7961]) | (layer2_outputs[7110]);
    assign outputs[10484] = layer2_outputs[1557];
    assign outputs[10485] = ~(layer2_outputs[1008]);
    assign outputs[10486] = ~(layer2_outputs[9199]);
    assign outputs[10487] = ~((layer2_outputs[12214]) ^ (layer2_outputs[3142]));
    assign outputs[10488] = layer2_outputs[2900];
    assign outputs[10489] = ~(layer2_outputs[2536]);
    assign outputs[10490] = (layer2_outputs[1114]) ^ (layer2_outputs[12251]);
    assign outputs[10491] = (layer2_outputs[4809]) ^ (layer2_outputs[8436]);
    assign outputs[10492] = ~((layer2_outputs[3820]) & (layer2_outputs[2993]));
    assign outputs[10493] = ~((layer2_outputs[744]) ^ (layer2_outputs[2584]));
    assign outputs[10494] = layer2_outputs[12299];
    assign outputs[10495] = ~((layer2_outputs[11539]) ^ (layer2_outputs[6515]));
    assign outputs[10496] = ~((layer2_outputs[113]) ^ (layer2_outputs[6552]));
    assign outputs[10497] = (layer2_outputs[5577]) & ~(layer2_outputs[7558]);
    assign outputs[10498] = (layer2_outputs[2646]) | (layer2_outputs[3053]);
    assign outputs[10499] = layer2_outputs[2335];
    assign outputs[10500] = ~(layer2_outputs[8285]);
    assign outputs[10501] = layer2_outputs[10239];
    assign outputs[10502] = ~(layer2_outputs[8602]);
    assign outputs[10503] = layer2_outputs[11674];
    assign outputs[10504] = ~((layer2_outputs[7431]) ^ (layer2_outputs[11182]));
    assign outputs[10505] = ~((layer2_outputs[8520]) & (layer2_outputs[9555]));
    assign outputs[10506] = ~((layer2_outputs[8296]) ^ (layer2_outputs[2099]));
    assign outputs[10507] = ~(layer2_outputs[8479]);
    assign outputs[10508] = ~((layer2_outputs[6993]) ^ (layer2_outputs[8472]));
    assign outputs[10509] = layer2_outputs[2886];
    assign outputs[10510] = ~(layer2_outputs[7535]);
    assign outputs[10511] = ~(layer2_outputs[2083]);
    assign outputs[10512] = ~(layer2_outputs[3988]) | (layer2_outputs[9691]);
    assign outputs[10513] = layer2_outputs[5448];
    assign outputs[10514] = (layer2_outputs[8199]) ^ (layer2_outputs[2603]);
    assign outputs[10515] = ~((layer2_outputs[5446]) ^ (layer2_outputs[5752]));
    assign outputs[10516] = ~((layer2_outputs[3463]) & (layer2_outputs[6198]));
    assign outputs[10517] = layer2_outputs[10115];
    assign outputs[10518] = (layer2_outputs[1348]) ^ (layer2_outputs[6046]);
    assign outputs[10519] = ~(layer2_outputs[4236]) | (layer2_outputs[10557]);
    assign outputs[10520] = ~(layer2_outputs[2090]);
    assign outputs[10521] = (layer2_outputs[8760]) ^ (layer2_outputs[11719]);
    assign outputs[10522] = (layer2_outputs[11831]) ^ (layer2_outputs[4119]);
    assign outputs[10523] = layer2_outputs[11859];
    assign outputs[10524] = layer2_outputs[2914];
    assign outputs[10525] = layer2_outputs[4559];
    assign outputs[10526] = ~(layer2_outputs[4170]);
    assign outputs[10527] = ~((layer2_outputs[8549]) ^ (layer2_outputs[4145]));
    assign outputs[10528] = (layer2_outputs[5141]) ^ (layer2_outputs[10137]);
    assign outputs[10529] = ~(layer2_outputs[11392]);
    assign outputs[10530] = ~(layer2_outputs[3302]);
    assign outputs[10531] = (layer2_outputs[4438]) ^ (layer2_outputs[4505]);
    assign outputs[10532] = ~(layer2_outputs[10406]);
    assign outputs[10533] = layer2_outputs[565];
    assign outputs[10534] = layer2_outputs[9755];
    assign outputs[10535] = ~(layer2_outputs[4870]);
    assign outputs[10536] = ~(layer2_outputs[11891]);
    assign outputs[10537] = ~(layer2_outputs[4209]);
    assign outputs[10538] = ~(layer2_outputs[536]);
    assign outputs[10539] = ~(layer2_outputs[4216]);
    assign outputs[10540] = layer2_outputs[9088];
    assign outputs[10541] = ~(layer2_outputs[11878]);
    assign outputs[10542] = ~(layer2_outputs[12049]) | (layer2_outputs[2092]);
    assign outputs[10543] = ~(layer2_outputs[9891]);
    assign outputs[10544] = ~((layer2_outputs[6304]) ^ (layer2_outputs[3042]));
    assign outputs[10545] = ~((layer2_outputs[8096]) ^ (layer2_outputs[4467]));
    assign outputs[10546] = (layer2_outputs[6485]) ^ (layer2_outputs[7036]);
    assign outputs[10547] = ~(layer2_outputs[5135]) | (layer2_outputs[7138]);
    assign outputs[10548] = layer2_outputs[4973];
    assign outputs[10549] = ~((layer2_outputs[12451]) | (layer2_outputs[10669]));
    assign outputs[10550] = ~((layer2_outputs[1690]) & (layer2_outputs[5147]));
    assign outputs[10551] = ~((layer2_outputs[2208]) ^ (layer2_outputs[3355]));
    assign outputs[10552] = layer2_outputs[3111];
    assign outputs[10553] = ~(layer2_outputs[47]);
    assign outputs[10554] = ~(layer2_outputs[3079]);
    assign outputs[10555] = ~(layer2_outputs[4663]);
    assign outputs[10556] = ~((layer2_outputs[11757]) ^ (layer2_outputs[8101]));
    assign outputs[10557] = (layer2_outputs[10537]) & (layer2_outputs[11748]);
    assign outputs[10558] = ~(layer2_outputs[9151]) | (layer2_outputs[10941]);
    assign outputs[10559] = ~((layer2_outputs[12264]) ^ (layer2_outputs[214]));
    assign outputs[10560] = (layer2_outputs[10825]) ^ (layer2_outputs[6404]);
    assign outputs[10561] = layer2_outputs[6292];
    assign outputs[10562] = ~(layer2_outputs[6965]);
    assign outputs[10563] = layer2_outputs[9373];
    assign outputs[10564] = (layer2_outputs[6884]) & (layer2_outputs[2546]);
    assign outputs[10565] = (layer2_outputs[2509]) ^ (layer2_outputs[4106]);
    assign outputs[10566] = ~((layer2_outputs[4610]) ^ (layer2_outputs[3022]));
    assign outputs[10567] = ~((layer2_outputs[398]) & (layer2_outputs[8658]));
    assign outputs[10568] = (layer2_outputs[7018]) ^ (layer2_outputs[9322]);
    assign outputs[10569] = (layer2_outputs[11359]) & (layer2_outputs[9704]);
    assign outputs[10570] = ~(layer2_outputs[3464]);
    assign outputs[10571] = ~(layer2_outputs[9833]);
    assign outputs[10572] = ~((layer2_outputs[11668]) ^ (layer2_outputs[4701]));
    assign outputs[10573] = layer2_outputs[6897];
    assign outputs[10574] = ~(layer2_outputs[9273]);
    assign outputs[10575] = ~((layer2_outputs[7413]) ^ (layer2_outputs[6343]));
    assign outputs[10576] = (layer2_outputs[4152]) ^ (layer2_outputs[8342]);
    assign outputs[10577] = ~((layer2_outputs[1043]) ^ (layer2_outputs[12757]));
    assign outputs[10578] = ~(layer2_outputs[2267]);
    assign outputs[10579] = ~((layer2_outputs[8622]) ^ (layer2_outputs[12411]));
    assign outputs[10580] = ~((layer2_outputs[1853]) ^ (layer2_outputs[4336]));
    assign outputs[10581] = ~(layer2_outputs[6540]);
    assign outputs[10582] = ~(layer2_outputs[11793]);
    assign outputs[10583] = (layer2_outputs[11582]) ^ (layer2_outputs[997]);
    assign outputs[10584] = ~((layer2_outputs[1931]) & (layer2_outputs[5079]));
    assign outputs[10585] = layer2_outputs[365];
    assign outputs[10586] = layer2_outputs[6274];
    assign outputs[10587] = layer2_outputs[8793];
    assign outputs[10588] = layer2_outputs[1989];
    assign outputs[10589] = ~((layer2_outputs[9374]) & (layer2_outputs[11699]));
    assign outputs[10590] = ~((layer2_outputs[4747]) ^ (layer2_outputs[11006]));
    assign outputs[10591] = ~(layer2_outputs[5799]) | (layer2_outputs[7100]);
    assign outputs[10592] = ~(layer2_outputs[9833]);
    assign outputs[10593] = layer2_outputs[8165];
    assign outputs[10594] = layer2_outputs[317];
    assign outputs[10595] = ~(layer2_outputs[9493]);
    assign outputs[10596] = ~(layer2_outputs[9607]) | (layer2_outputs[10019]);
    assign outputs[10597] = ~((layer2_outputs[1267]) ^ (layer2_outputs[3866]));
    assign outputs[10598] = (layer2_outputs[11533]) ^ (layer2_outputs[3346]);
    assign outputs[10599] = (layer2_outputs[2269]) & ~(layer2_outputs[2561]);
    assign outputs[10600] = layer2_outputs[4931];
    assign outputs[10601] = layer2_outputs[10434];
    assign outputs[10602] = ~((layer2_outputs[8939]) ^ (layer2_outputs[5761]));
    assign outputs[10603] = layer2_outputs[5401];
    assign outputs[10604] = ~((layer2_outputs[9445]) & (layer2_outputs[959]));
    assign outputs[10605] = layer2_outputs[282];
    assign outputs[10606] = ~(layer2_outputs[2959]) | (layer2_outputs[10811]);
    assign outputs[10607] = (layer2_outputs[9379]) ^ (layer2_outputs[12550]);
    assign outputs[10608] = (layer2_outputs[6492]) | (layer2_outputs[4255]);
    assign outputs[10609] = layer2_outputs[7462];
    assign outputs[10610] = layer2_outputs[3722];
    assign outputs[10611] = ~((layer2_outputs[5066]) ^ (layer2_outputs[9261]));
    assign outputs[10612] = (layer2_outputs[7529]) ^ (layer2_outputs[10572]);
    assign outputs[10613] = layer2_outputs[9591];
    assign outputs[10614] = (layer2_outputs[4105]) ^ (layer2_outputs[8956]);
    assign outputs[10615] = layer2_outputs[12729];
    assign outputs[10616] = (layer2_outputs[11199]) ^ (layer2_outputs[599]);
    assign outputs[10617] = ~(layer2_outputs[6048]) | (layer2_outputs[1855]);
    assign outputs[10618] = (layer2_outputs[1709]) ^ (layer2_outputs[12599]);
    assign outputs[10619] = (layer2_outputs[6992]) ^ (layer2_outputs[1144]);
    assign outputs[10620] = layer2_outputs[8094];
    assign outputs[10621] = layer2_outputs[1529];
    assign outputs[10622] = (layer2_outputs[3242]) ^ (layer2_outputs[8862]);
    assign outputs[10623] = layer2_outputs[4192];
    assign outputs[10624] = ~((layer2_outputs[981]) ^ (layer2_outputs[11994]));
    assign outputs[10625] = ~(layer2_outputs[3046]) | (layer2_outputs[6075]);
    assign outputs[10626] = ~((layer2_outputs[2866]) ^ (layer2_outputs[9590]));
    assign outputs[10627] = layer2_outputs[391];
    assign outputs[10628] = (layer2_outputs[4322]) & ~(layer2_outputs[4979]);
    assign outputs[10629] = ~(layer2_outputs[5590]);
    assign outputs[10630] = (layer2_outputs[11225]) ^ (layer2_outputs[11888]);
    assign outputs[10631] = ~(layer2_outputs[2852]);
    assign outputs[10632] = (layer2_outputs[11099]) | (layer2_outputs[5731]);
    assign outputs[10633] = ~((layer2_outputs[7017]) ^ (layer2_outputs[5957]));
    assign outputs[10634] = ~((layer2_outputs[4901]) & (layer2_outputs[742]));
    assign outputs[10635] = layer2_outputs[8860];
    assign outputs[10636] = ~((layer2_outputs[8292]) ^ (layer2_outputs[6653]));
    assign outputs[10637] = ~(layer2_outputs[9185]) | (layer2_outputs[4551]);
    assign outputs[10638] = layer2_outputs[3613];
    assign outputs[10639] = ~(layer2_outputs[3622]);
    assign outputs[10640] = (layer2_outputs[3580]) & ~(layer2_outputs[5239]);
    assign outputs[10641] = ~((layer2_outputs[9702]) | (layer2_outputs[2730]));
    assign outputs[10642] = ~(layer2_outputs[10313]) | (layer2_outputs[9109]);
    assign outputs[10643] = (layer2_outputs[12635]) ^ (layer2_outputs[5019]);
    assign outputs[10644] = layer2_outputs[1174];
    assign outputs[10645] = ~(layer2_outputs[8616]);
    assign outputs[10646] = ~((layer2_outputs[7494]) ^ (layer2_outputs[7398]));
    assign outputs[10647] = ~((layer2_outputs[5652]) ^ (layer2_outputs[529]));
    assign outputs[10648] = ~(layer2_outputs[7894]);
    assign outputs[10649] = ~(layer2_outputs[9385]);
    assign outputs[10650] = layer2_outputs[11433];
    assign outputs[10651] = ~(layer2_outputs[8697]) | (layer2_outputs[2782]);
    assign outputs[10652] = layer2_outputs[350];
    assign outputs[10653] = (layer2_outputs[5078]) ^ (layer2_outputs[2672]);
    assign outputs[10654] = (layer2_outputs[858]) & ~(layer2_outputs[8982]);
    assign outputs[10655] = ~(layer2_outputs[1731]) | (layer2_outputs[1790]);
    assign outputs[10656] = ~(layer2_outputs[9311]);
    assign outputs[10657] = ~((layer2_outputs[7940]) ^ (layer2_outputs[12128]));
    assign outputs[10658] = (layer2_outputs[8950]) & ~(layer2_outputs[11355]);
    assign outputs[10659] = ~(layer2_outputs[5534]) | (layer2_outputs[7364]);
    assign outputs[10660] = ~(layer2_outputs[3648]);
    assign outputs[10661] = ~((layer2_outputs[9100]) ^ (layer2_outputs[2864]));
    assign outputs[10662] = (layer2_outputs[9340]) & ~(layer2_outputs[1648]);
    assign outputs[10663] = (layer2_outputs[11028]) ^ (layer2_outputs[3975]);
    assign outputs[10664] = ~((layer2_outputs[184]) & (layer2_outputs[8173]));
    assign outputs[10665] = (layer2_outputs[5057]) ^ (layer2_outputs[347]);
    assign outputs[10666] = ~(layer2_outputs[1608]) | (layer2_outputs[7307]);
    assign outputs[10667] = ~((layer2_outputs[11495]) ^ (layer2_outputs[5954]));
    assign outputs[10668] = ~((layer2_outputs[4560]) ^ (layer2_outputs[8719]));
    assign outputs[10669] = ~(layer2_outputs[12437]);
    assign outputs[10670] = layer2_outputs[4727];
    assign outputs[10671] = ~((layer2_outputs[12672]) | (layer2_outputs[3871]));
    assign outputs[10672] = (layer2_outputs[5446]) ^ (layer2_outputs[11571]);
    assign outputs[10673] = ~((layer2_outputs[4232]) ^ (layer2_outputs[7196]));
    assign outputs[10674] = layer2_outputs[8510];
    assign outputs[10675] = ~((layer2_outputs[10359]) ^ (layer2_outputs[7150]));
    assign outputs[10676] = (layer2_outputs[12020]) ^ (layer2_outputs[4270]);
    assign outputs[10677] = layer2_outputs[7696];
    assign outputs[10678] = ~(layer2_outputs[5186]);
    assign outputs[10679] = (layer2_outputs[9556]) ^ (layer2_outputs[3253]);
    assign outputs[10680] = ~(layer2_outputs[11215]);
    assign outputs[10681] = layer2_outputs[3143];
    assign outputs[10682] = (layer2_outputs[8261]) | (layer2_outputs[6576]);
    assign outputs[10683] = (layer2_outputs[3721]) ^ (layer2_outputs[129]);
    assign outputs[10684] = ~(layer2_outputs[1414]);
    assign outputs[10685] = ~(layer2_outputs[10595]) | (layer2_outputs[4]);
    assign outputs[10686] = ~(layer2_outputs[572]);
    assign outputs[10687] = ~((layer2_outputs[2518]) ^ (layer2_outputs[1703]));
    assign outputs[10688] = ~((layer2_outputs[11182]) ^ (layer2_outputs[7404]));
    assign outputs[10689] = layer2_outputs[1351];
    assign outputs[10690] = (layer2_outputs[6694]) & ~(layer2_outputs[6601]);
    assign outputs[10691] = (layer2_outputs[153]) | (layer2_outputs[3809]);
    assign outputs[10692] = ~((layer2_outputs[6972]) | (layer2_outputs[504]));
    assign outputs[10693] = (layer2_outputs[11676]) ^ (layer2_outputs[5299]);
    assign outputs[10694] = ~(layer2_outputs[3760]);
    assign outputs[10695] = ~((layer2_outputs[8443]) & (layer2_outputs[5433]));
    assign outputs[10696] = (layer2_outputs[341]) ^ (layer2_outputs[3449]);
    assign outputs[10697] = (layer2_outputs[2372]) ^ (layer2_outputs[6249]);
    assign outputs[10698] = ~((layer2_outputs[9914]) ^ (layer2_outputs[2890]));
    assign outputs[10699] = layer2_outputs[11153];
    assign outputs[10700] = (layer2_outputs[2582]) ^ (layer2_outputs[3012]);
    assign outputs[10701] = ~(layer2_outputs[10070]) | (layer2_outputs[9574]);
    assign outputs[10702] = layer2_outputs[6250];
    assign outputs[10703] = (layer2_outputs[9354]) & ~(layer2_outputs[10867]);
    assign outputs[10704] = ~(layer2_outputs[4875]);
    assign outputs[10705] = ~(layer2_outputs[10256]) | (layer2_outputs[7764]);
    assign outputs[10706] = (layer2_outputs[11770]) & (layer2_outputs[2127]);
    assign outputs[10707] = ~((layer2_outputs[11317]) ^ (layer2_outputs[4528]));
    assign outputs[10708] = (layer2_outputs[1881]) ^ (layer2_outputs[6127]);
    assign outputs[10709] = (layer2_outputs[869]) ^ (layer2_outputs[4472]);
    assign outputs[10710] = layer2_outputs[431];
    assign outputs[10711] = layer2_outputs[11686];
    assign outputs[10712] = layer2_outputs[10272];
    assign outputs[10713] = ~(layer2_outputs[4854]);
    assign outputs[10714] = layer2_outputs[8933];
    assign outputs[10715] = ~((layer2_outputs[10717]) ^ (layer2_outputs[8059]));
    assign outputs[10716] = layer2_outputs[11438];
    assign outputs[10717] = layer2_outputs[12473];
    assign outputs[10718] = ~((layer2_outputs[1068]) & (layer2_outputs[5840]));
    assign outputs[10719] = layer2_outputs[9818];
    assign outputs[10720] = layer2_outputs[1411];
    assign outputs[10721] = ~(layer2_outputs[9483]);
    assign outputs[10722] = ~(layer2_outputs[4366]);
    assign outputs[10723] = (layer2_outputs[12196]) & ~(layer2_outputs[9478]);
    assign outputs[10724] = layer2_outputs[934];
    assign outputs[10725] = ~(layer2_outputs[3514]);
    assign outputs[10726] = layer2_outputs[11623];
    assign outputs[10727] = layer2_outputs[558];
    assign outputs[10728] = ~(layer2_outputs[3843]);
    assign outputs[10729] = ~((layer2_outputs[10856]) ^ (layer2_outputs[8379]));
    assign outputs[10730] = (layer2_outputs[10480]) & (layer2_outputs[9324]);
    assign outputs[10731] = (layer2_outputs[8908]) ^ (layer2_outputs[8233]);
    assign outputs[10732] = ~(layer2_outputs[3105]) | (layer2_outputs[1327]);
    assign outputs[10733] = ~(layer2_outputs[4524]);
    assign outputs[10734] = ~(layer2_outputs[9600]);
    assign outputs[10735] = ~(layer2_outputs[6830]);
    assign outputs[10736] = layer2_outputs[2271];
    assign outputs[10737] = ~((layer2_outputs[488]) ^ (layer2_outputs[2180]));
    assign outputs[10738] = ~(layer2_outputs[11520]);
    assign outputs[10739] = ~((layer2_outputs[12648]) | (layer2_outputs[4258]));
    assign outputs[10740] = layer2_outputs[12098];
    assign outputs[10741] = ~((layer2_outputs[395]) & (layer2_outputs[5127]));
    assign outputs[10742] = ~(layer2_outputs[3939]);
    assign outputs[10743] = layer2_outputs[12402];
    assign outputs[10744] = ~(layer2_outputs[7400]);
    assign outputs[10745] = ~(layer2_outputs[7108]);
    assign outputs[10746] = ~((layer2_outputs[8016]) ^ (layer2_outputs[1605]));
    assign outputs[10747] = (layer2_outputs[11166]) ^ (layer2_outputs[2601]);
    assign outputs[10748] = (layer2_outputs[10843]) ^ (layer2_outputs[3823]);
    assign outputs[10749] = layer2_outputs[9154];
    assign outputs[10750] = layer2_outputs[1639];
    assign outputs[10751] = ~((layer2_outputs[4058]) & (layer2_outputs[3475]));
    assign outputs[10752] = ~((layer2_outputs[5097]) & (layer2_outputs[1046]));
    assign outputs[10753] = ~((layer2_outputs[10808]) & (layer2_outputs[12577]));
    assign outputs[10754] = ~(layer2_outputs[6885]);
    assign outputs[10755] = ~(layer2_outputs[10779]);
    assign outputs[10756] = ~((layer2_outputs[10511]) ^ (layer2_outputs[4064]));
    assign outputs[10757] = ~((layer2_outputs[12027]) ^ (layer2_outputs[1204]));
    assign outputs[10758] = ~(layer2_outputs[10400]) | (layer2_outputs[413]);
    assign outputs[10759] = ~(layer2_outputs[10752]);
    assign outputs[10760] = layer2_outputs[4304];
    assign outputs[10761] = (layer2_outputs[6167]) ^ (layer2_outputs[1188]);
    assign outputs[10762] = ~(layer2_outputs[10962]);
    assign outputs[10763] = ~(layer2_outputs[12055]) | (layer2_outputs[2063]);
    assign outputs[10764] = ~(layer2_outputs[394]) | (layer2_outputs[1540]);
    assign outputs[10765] = layer2_outputs[4185];
    assign outputs[10766] = ~(layer2_outputs[3596]) | (layer2_outputs[2185]);
    assign outputs[10767] = ~((layer2_outputs[2878]) ^ (layer2_outputs[1474]));
    assign outputs[10768] = (layer2_outputs[6058]) ^ (layer2_outputs[8999]);
    assign outputs[10769] = layer2_outputs[12084];
    assign outputs[10770] = layer2_outputs[3525];
    assign outputs[10771] = layer2_outputs[9513];
    assign outputs[10772] = ~((layer2_outputs[6366]) ^ (layer2_outputs[9033]));
    assign outputs[10773] = (layer2_outputs[9546]) & ~(layer2_outputs[12284]);
    assign outputs[10774] = ~((layer2_outputs[9403]) ^ (layer2_outputs[2075]));
    assign outputs[10775] = ~(layer2_outputs[8605]);
    assign outputs[10776] = ~(layer2_outputs[9478]);
    assign outputs[10777] = layer2_outputs[11258];
    assign outputs[10778] = layer2_outputs[11587];
    assign outputs[10779] = ~((layer2_outputs[12798]) | (layer2_outputs[5766]));
    assign outputs[10780] = ~((layer2_outputs[12486]) & (layer2_outputs[6177]));
    assign outputs[10781] = layer2_outputs[2493];
    assign outputs[10782] = layer2_outputs[9192];
    assign outputs[10783] = ~((layer2_outputs[6460]) ^ (layer2_outputs[11977]));
    assign outputs[10784] = ~((layer2_outputs[10262]) ^ (layer2_outputs[422]));
    assign outputs[10785] = ~(layer2_outputs[8758]) | (layer2_outputs[8156]);
    assign outputs[10786] = ~((layer2_outputs[10356]) ^ (layer2_outputs[3260]));
    assign outputs[10787] = (layer2_outputs[10258]) & ~(layer2_outputs[7475]);
    assign outputs[10788] = ~(layer2_outputs[10038]) | (layer2_outputs[6850]);
    assign outputs[10789] = ~(layer2_outputs[8584]);
    assign outputs[10790] = ~(layer2_outputs[1499]);
    assign outputs[10791] = ~((layer2_outputs[399]) ^ (layer2_outputs[4719]));
    assign outputs[10792] = layer2_outputs[1705];
    assign outputs[10793] = (layer2_outputs[9843]) | (layer2_outputs[5527]);
    assign outputs[10794] = ~(layer2_outputs[9817]);
    assign outputs[10795] = ~(layer2_outputs[11178]) | (layer2_outputs[2417]);
    assign outputs[10796] = layer2_outputs[6258];
    assign outputs[10797] = layer2_outputs[3752];
    assign outputs[10798] = ~((layer2_outputs[4597]) & (layer2_outputs[9073]));
    assign outputs[10799] = ~(layer2_outputs[9509]);
    assign outputs[10800] = (layer2_outputs[1842]) ^ (layer2_outputs[3660]);
    assign outputs[10801] = layer2_outputs[10306];
    assign outputs[10802] = layer2_outputs[7787];
    assign outputs[10803] = ~(layer2_outputs[1675]);
    assign outputs[10804] = ~((layer2_outputs[2285]) ^ (layer2_outputs[7098]));
    assign outputs[10805] = ~(layer2_outputs[8861]) | (layer2_outputs[3706]);
    assign outputs[10806] = ~((layer2_outputs[4755]) ^ (layer2_outputs[150]));
    assign outputs[10807] = layer2_outputs[12723];
    assign outputs[10808] = (layer2_outputs[10633]) ^ (layer2_outputs[12551]);
    assign outputs[10809] = (layer2_outputs[12759]) ^ (layer2_outputs[5156]);
    assign outputs[10810] = ~((layer2_outputs[3426]) ^ (layer2_outputs[6410]));
    assign outputs[10811] = ~(layer2_outputs[1446]);
    assign outputs[10812] = ~(layer2_outputs[3418]);
    assign outputs[10813] = layer2_outputs[2168];
    assign outputs[10814] = (layer2_outputs[12117]) & (layer2_outputs[7904]);
    assign outputs[10815] = layer2_outputs[5894];
    assign outputs[10816] = ~((layer2_outputs[3368]) ^ (layer2_outputs[4598]));
    assign outputs[10817] = (layer2_outputs[11380]) ^ (layer2_outputs[10809]);
    assign outputs[10818] = ~(layer2_outputs[4731]);
    assign outputs[10819] = layer2_outputs[12091];
    assign outputs[10820] = ~((layer2_outputs[505]) ^ (layer2_outputs[7728]));
    assign outputs[10821] = layer2_outputs[11621];
    assign outputs[10822] = ~((layer2_outputs[10536]) ^ (layer2_outputs[10787]));
    assign outputs[10823] = ~(layer2_outputs[12436]);
    assign outputs[10824] = (layer2_outputs[7551]) | (layer2_outputs[12783]);
    assign outputs[10825] = (layer2_outputs[9252]) & (layer2_outputs[7213]);
    assign outputs[10826] = ~(layer2_outputs[760]);
    assign outputs[10827] = layer2_outputs[6897];
    assign outputs[10828] = ~(layer2_outputs[5481]);
    assign outputs[10829] = ~(layer2_outputs[12796]);
    assign outputs[10830] = ~((layer2_outputs[6834]) & (layer2_outputs[7539]));
    assign outputs[10831] = layer2_outputs[11378];
    assign outputs[10832] = layer2_outputs[12089];
    assign outputs[10833] = ~(layer2_outputs[2441]);
    assign outputs[10834] = ~(layer2_outputs[8231]);
    assign outputs[10835] = layer2_outputs[2321];
    assign outputs[10836] = layer2_outputs[1900];
    assign outputs[10837] = ~((layer2_outputs[11424]) ^ (layer2_outputs[375]));
    assign outputs[10838] = ~(layer2_outputs[6677]);
    assign outputs[10839] = layer2_outputs[11007];
    assign outputs[10840] = ~(layer2_outputs[4225]);
    assign outputs[10841] = (layer2_outputs[8769]) & (layer2_outputs[6808]);
    assign outputs[10842] = ~(layer2_outputs[992]);
    assign outputs[10843] = ~(layer2_outputs[300]);
    assign outputs[10844] = ~(layer2_outputs[11241]);
    assign outputs[10845] = ~(layer2_outputs[2055]) | (layer2_outputs[2678]);
    assign outputs[10846] = layer2_outputs[4016];
    assign outputs[10847] = ~(layer2_outputs[6254]);
    assign outputs[10848] = ~(layer2_outputs[11412]);
    assign outputs[10849] = layer2_outputs[8224];
    assign outputs[10850] = layer2_outputs[10883];
    assign outputs[10851] = layer2_outputs[6033];
    assign outputs[10852] = (layer2_outputs[12698]) ^ (layer2_outputs[2491]);
    assign outputs[10853] = ~((layer2_outputs[11622]) ^ (layer2_outputs[4375]));
    assign outputs[10854] = (layer2_outputs[11207]) ^ (layer2_outputs[3512]);
    assign outputs[10855] = (layer2_outputs[8870]) & ~(layer2_outputs[12231]);
    assign outputs[10856] = ~((layer2_outputs[5509]) ^ (layer2_outputs[3572]));
    assign outputs[10857] = (layer2_outputs[5211]) & (layer2_outputs[11734]);
    assign outputs[10858] = ~(layer2_outputs[2931]) | (layer2_outputs[7764]);
    assign outputs[10859] = ~((layer2_outputs[11310]) ^ (layer2_outputs[319]));
    assign outputs[10860] = ~((layer2_outputs[11266]) ^ (layer2_outputs[7334]));
    assign outputs[10861] = (layer2_outputs[5174]) ^ (layer2_outputs[7882]);
    assign outputs[10862] = (layer2_outputs[5189]) ^ (layer2_outputs[8030]);
    assign outputs[10863] = layer2_outputs[4239];
    assign outputs[10864] = (layer2_outputs[11575]) | (layer2_outputs[8898]);
    assign outputs[10865] = (layer2_outputs[9190]) ^ (layer2_outputs[9529]);
    assign outputs[10866] = (layer2_outputs[3759]) ^ (layer2_outputs[7101]);
    assign outputs[10867] = layer2_outputs[3701];
    assign outputs[10868] = layer2_outputs[7096];
    assign outputs[10869] = layer2_outputs[10827];
    assign outputs[10870] = (layer2_outputs[5307]) | (layer2_outputs[2273]);
    assign outputs[10871] = ~(layer2_outputs[4045]);
    assign outputs[10872] = (layer2_outputs[9967]) ^ (layer2_outputs[196]);
    assign outputs[10873] = ~(layer2_outputs[12518]) | (layer2_outputs[3628]);
    assign outputs[10874] = ~((layer2_outputs[8743]) & (layer2_outputs[1054]));
    assign outputs[10875] = (layer2_outputs[2177]) ^ (layer2_outputs[2359]);
    assign outputs[10876] = layer2_outputs[1314];
    assign outputs[10877] = ~(layer2_outputs[10849]);
    assign outputs[10878] = ~(layer2_outputs[12796]);
    assign outputs[10879] = (layer2_outputs[10548]) ^ (layer2_outputs[1907]);
    assign outputs[10880] = layer2_outputs[12715];
    assign outputs[10881] = ~((layer2_outputs[11788]) & (layer2_outputs[6140]));
    assign outputs[10882] = (layer2_outputs[4181]) ^ (layer2_outputs[9263]);
    assign outputs[10883] = layer2_outputs[9640];
    assign outputs[10884] = layer2_outputs[9475];
    assign outputs[10885] = ~(layer2_outputs[4446]);
    assign outputs[10886] = layer2_outputs[8227];
    assign outputs[10887] = ~(layer2_outputs[8290]);
    assign outputs[10888] = ~(layer2_outputs[11868]);
    assign outputs[10889] = ~(layer2_outputs[12307]) | (layer2_outputs[1781]);
    assign outputs[10890] = ~((layer2_outputs[5873]) ^ (layer2_outputs[8845]));
    assign outputs[10891] = layer2_outputs[4168];
    assign outputs[10892] = ~((layer2_outputs[6894]) ^ (layer2_outputs[1889]));
    assign outputs[10893] = ~((layer2_outputs[9328]) & (layer2_outputs[12792]));
    assign outputs[10894] = (layer2_outputs[542]) | (layer2_outputs[1460]);
    assign outputs[10895] = layer2_outputs[2265];
    assign outputs[10896] = layer2_outputs[11571];
    assign outputs[10897] = (layer2_outputs[3920]) | (layer2_outputs[2629]);
    assign outputs[10898] = (layer2_outputs[6096]) ^ (layer2_outputs[4604]);
    assign outputs[10899] = layer2_outputs[924];
    assign outputs[10900] = layer2_outputs[8383];
    assign outputs[10901] = layer2_outputs[3903];
    assign outputs[10902] = layer2_outputs[11342];
    assign outputs[10903] = layer2_outputs[2676];
    assign outputs[10904] = ~((layer2_outputs[2455]) ^ (layer2_outputs[10452]));
    assign outputs[10905] = ~((layer2_outputs[335]) ^ (layer2_outputs[1788]));
    assign outputs[10906] = layer2_outputs[10405];
    assign outputs[10907] = layer2_outputs[675];
    assign outputs[10908] = ~(layer2_outputs[2474]);
    assign outputs[10909] = (layer2_outputs[12282]) & (layer2_outputs[4262]);
    assign outputs[10910] = ~(layer2_outputs[3800]) | (layer2_outputs[4056]);
    assign outputs[10911] = ~(layer2_outputs[4135]);
    assign outputs[10912] = ~(layer2_outputs[11025]);
    assign outputs[10913] = layer2_outputs[12559];
    assign outputs[10914] = (layer2_outputs[2129]) ^ (layer2_outputs[4881]);
    assign outputs[10915] = (layer2_outputs[3252]) ^ (layer2_outputs[11717]);
    assign outputs[10916] = (layer2_outputs[11142]) ^ (layer2_outputs[9496]);
    assign outputs[10917] = ~(layer2_outputs[2372]);
    assign outputs[10918] = ~((layer2_outputs[5515]) ^ (layer2_outputs[8259]));
    assign outputs[10919] = layer2_outputs[6921];
    assign outputs[10920] = ~(layer2_outputs[5274]);
    assign outputs[10921] = (layer2_outputs[3209]) ^ (layer2_outputs[9346]);
    assign outputs[10922] = (layer2_outputs[3128]) ^ (layer2_outputs[712]);
    assign outputs[10923] = (layer2_outputs[1352]) | (layer2_outputs[10089]);
    assign outputs[10924] = layer2_outputs[9876];
    assign outputs[10925] = ~((layer2_outputs[3954]) ^ (layer2_outputs[3791]));
    assign outputs[10926] = layer2_outputs[1389];
    assign outputs[10927] = ~((layer2_outputs[3271]) ^ (layer2_outputs[11921]));
    assign outputs[10928] = (layer2_outputs[11722]) & (layer2_outputs[2727]);
    assign outputs[10929] = ~(layer2_outputs[3617]);
    assign outputs[10930] = layer2_outputs[2379];
    assign outputs[10931] = layer2_outputs[391];
    assign outputs[10932] = ~((layer2_outputs[6609]) ^ (layer2_outputs[2410]));
    assign outputs[10933] = layer2_outputs[1828];
    assign outputs[10934] = layer2_outputs[5176];
    assign outputs[10935] = ~(layer2_outputs[1550]);
    assign outputs[10936] = ~(layer2_outputs[9700]) | (layer2_outputs[2364]);
    assign outputs[10937] = ~((layer2_outputs[1840]) ^ (layer2_outputs[6493]));
    assign outputs[10938] = (layer2_outputs[5181]) ^ (layer2_outputs[7553]);
    assign outputs[10939] = ~(layer2_outputs[1580]);
    assign outputs[10940] = ~(layer2_outputs[11649]);
    assign outputs[10941] = (layer2_outputs[2498]) ^ (layer2_outputs[4664]);
    assign outputs[10942] = ~((layer2_outputs[184]) & (layer2_outputs[1008]));
    assign outputs[10943] = (layer2_outputs[2851]) & (layer2_outputs[9586]);
    assign outputs[10944] = ~(layer2_outputs[12615]);
    assign outputs[10945] = (layer2_outputs[6671]) | (layer2_outputs[8282]);
    assign outputs[10946] = ~((layer2_outputs[5874]) ^ (layer2_outputs[2223]));
    assign outputs[10947] = ~(layer2_outputs[7327]);
    assign outputs[10948] = (layer2_outputs[1645]) ^ (layer2_outputs[1958]);
    assign outputs[10949] = ~((layer2_outputs[2347]) ^ (layer2_outputs[7130]));
    assign outputs[10950] = layer2_outputs[10748];
    assign outputs[10951] = ~((layer2_outputs[1217]) ^ (layer2_outputs[3478]));
    assign outputs[10952] = layer2_outputs[11804];
    assign outputs[10953] = ~(layer2_outputs[4588]) | (layer2_outputs[5054]);
    assign outputs[10954] = (layer2_outputs[387]) | (layer2_outputs[2464]);
    assign outputs[10955] = layer2_outputs[7110];
    assign outputs[10956] = layer2_outputs[1066];
    assign outputs[10957] = layer2_outputs[2665];
    assign outputs[10958] = ~((layer2_outputs[7142]) ^ (layer2_outputs[3828]));
    assign outputs[10959] = ~((layer2_outputs[11899]) ^ (layer2_outputs[6853]));
    assign outputs[10960] = (layer2_outputs[11670]) ^ (layer2_outputs[9055]);
    assign outputs[10961] = ~(layer2_outputs[10588]) | (layer2_outputs[3615]);
    assign outputs[10962] = ~(layer2_outputs[1719]);
    assign outputs[10963] = ~(layer2_outputs[11291]);
    assign outputs[10964] = (layer2_outputs[9229]) ^ (layer2_outputs[6023]);
    assign outputs[10965] = (layer2_outputs[6505]) ^ (layer2_outputs[788]);
    assign outputs[10966] = ~((layer2_outputs[2545]) & (layer2_outputs[6298]));
    assign outputs[10967] = ~(layer2_outputs[6372]) | (layer2_outputs[4715]);
    assign outputs[10968] = ~((layer2_outputs[6472]) ^ (layer2_outputs[7022]));
    assign outputs[10969] = layer2_outputs[7081];
    assign outputs[10970] = ~(layer2_outputs[453]);
    assign outputs[10971] = layer2_outputs[11660];
    assign outputs[10972] = (layer2_outputs[312]) & (layer2_outputs[6908]);
    assign outputs[10973] = (layer2_outputs[6120]) ^ (layer2_outputs[3084]);
    assign outputs[10974] = layer2_outputs[8423];
    assign outputs[10975] = ~((layer2_outputs[4713]) & (layer2_outputs[4392]));
    assign outputs[10976] = (layer2_outputs[89]) ^ (layer2_outputs[697]);
    assign outputs[10977] = ~(layer2_outputs[4423]);
    assign outputs[10978] = layer2_outputs[2912];
    assign outputs[10979] = ~((layer2_outputs[1974]) ^ (layer2_outputs[170]));
    assign outputs[10980] = layer2_outputs[2194];
    assign outputs[10981] = ~(layer2_outputs[8357]) | (layer2_outputs[7752]);
    assign outputs[10982] = layer2_outputs[3671];
    assign outputs[10983] = ~(layer2_outputs[11513]) | (layer2_outputs[3119]);
    assign outputs[10984] = ~((layer2_outputs[10907]) ^ (layer2_outputs[3055]));
    assign outputs[10985] = ~(layer2_outputs[10535]);
    assign outputs[10986] = ~(layer2_outputs[9509]);
    assign outputs[10987] = (layer2_outputs[6413]) ^ (layer2_outputs[2929]);
    assign outputs[10988] = ~((layer2_outputs[7760]) ^ (layer2_outputs[8281]));
    assign outputs[10989] = (layer2_outputs[3131]) ^ (layer2_outputs[1740]);
    assign outputs[10990] = ~((layer2_outputs[6368]) & (layer2_outputs[7736]));
    assign outputs[10991] = (layer2_outputs[4253]) & ~(layer2_outputs[2651]);
    assign outputs[10992] = ~(layer2_outputs[12629]);
    assign outputs[10993] = ~(layer2_outputs[12687]);
    assign outputs[10994] = (layer2_outputs[4685]) | (layer2_outputs[10323]);
    assign outputs[10995] = ~((layer2_outputs[3856]) & (layer2_outputs[9937]));
    assign outputs[10996] = ~(layer2_outputs[10587]);
    assign outputs[10997] = ~(layer2_outputs[4125]);
    assign outputs[10998] = ~(layer2_outputs[7392]);
    assign outputs[10999] = 1'b1;
    assign outputs[11000] = ~(layer2_outputs[5557]);
    assign outputs[11001] = layer2_outputs[3247];
    assign outputs[11002] = ~(layer2_outputs[7560]);
    assign outputs[11003] = ~((layer2_outputs[12097]) ^ (layer2_outputs[10842]));
    assign outputs[11004] = ~((layer2_outputs[5470]) ^ (layer2_outputs[9121]));
    assign outputs[11005] = ~(layer2_outputs[12775]);
    assign outputs[11006] = ~((layer2_outputs[6049]) ^ (layer2_outputs[6319]));
    assign outputs[11007] = (layer2_outputs[11165]) ^ (layer2_outputs[3750]);
    assign outputs[11008] = ~(layer2_outputs[7770]);
    assign outputs[11009] = (layer2_outputs[11386]) ^ (layer2_outputs[7478]);
    assign outputs[11010] = ~(layer2_outputs[3725]);
    assign outputs[11011] = ~((layer2_outputs[2091]) ^ (layer2_outputs[3360]));
    assign outputs[11012] = (layer2_outputs[7389]) ^ (layer2_outputs[2746]);
    assign outputs[11013] = (layer2_outputs[12240]) ^ (layer2_outputs[8382]);
    assign outputs[11014] = ~(layer2_outputs[10028]) | (layer2_outputs[5193]);
    assign outputs[11015] = layer2_outputs[1411];
    assign outputs[11016] = ~(layer2_outputs[9312]);
    assign outputs[11017] = ~((layer2_outputs[6944]) ^ (layer2_outputs[5921]));
    assign outputs[11018] = ~(layer2_outputs[12618]);
    assign outputs[11019] = ~(layer2_outputs[11364]);
    assign outputs[11020] = layer2_outputs[12032];
    assign outputs[11021] = ~(layer2_outputs[5177]);
    assign outputs[11022] = (layer2_outputs[11227]) & (layer2_outputs[10979]);
    assign outputs[11023] = ~((layer2_outputs[11251]) ^ (layer2_outputs[3492]));
    assign outputs[11024] = layer2_outputs[9029];
    assign outputs[11025] = ~(layer2_outputs[5784]);
    assign outputs[11026] = (layer2_outputs[4994]) ^ (layer2_outputs[11841]);
    assign outputs[11027] = layer2_outputs[7251];
    assign outputs[11028] = (layer2_outputs[136]) & ~(layer2_outputs[8845]);
    assign outputs[11029] = (layer2_outputs[11851]) ^ (layer2_outputs[10161]);
    assign outputs[11030] = ~((layer2_outputs[7460]) ^ (layer2_outputs[531]));
    assign outputs[11031] = ~(layer2_outputs[3461]);
    assign outputs[11032] = ~(layer2_outputs[9608]);
    assign outputs[11033] = (layer2_outputs[10598]) ^ (layer2_outputs[4890]);
    assign outputs[11034] = (layer2_outputs[4716]) ^ (layer2_outputs[12746]);
    assign outputs[11035] = ~(layer2_outputs[1878]);
    assign outputs[11036] = ~((layer2_outputs[10589]) ^ (layer2_outputs[4992]));
    assign outputs[11037] = layer2_outputs[7787];
    assign outputs[11038] = layer2_outputs[6291];
    assign outputs[11039] = ~((layer2_outputs[1628]) & (layer2_outputs[12699]));
    assign outputs[11040] = (layer2_outputs[4348]) & (layer2_outputs[6446]);
    assign outputs[11041] = (layer2_outputs[11546]) | (layer2_outputs[4540]);
    assign outputs[11042] = (layer2_outputs[1896]) | (layer2_outputs[12371]);
    assign outputs[11043] = layer2_outputs[8878];
    assign outputs[11044] = (layer2_outputs[10175]) & ~(layer2_outputs[2425]);
    assign outputs[11045] = ~(layer2_outputs[11998]);
    assign outputs[11046] = ~(layer2_outputs[9957]) | (layer2_outputs[2219]);
    assign outputs[11047] = layer2_outputs[617];
    assign outputs[11048] = (layer2_outputs[6997]) ^ (layer2_outputs[251]);
    assign outputs[11049] = ~(layer2_outputs[3805]);
    assign outputs[11050] = ~((layer2_outputs[6479]) | (layer2_outputs[6072]));
    assign outputs[11051] = layer2_outputs[11621];
    assign outputs[11052] = layer2_outputs[238];
    assign outputs[11053] = ~(layer2_outputs[3464]) | (layer2_outputs[2492]);
    assign outputs[11054] = (layer2_outputs[3448]) ^ (layer2_outputs[11806]);
    assign outputs[11055] = ~(layer2_outputs[9861]);
    assign outputs[11056] = layer2_outputs[282];
    assign outputs[11057] = ~((layer2_outputs[4926]) & (layer2_outputs[1341]));
    assign outputs[11058] = (layer2_outputs[4697]) ^ (layer2_outputs[2309]);
    assign outputs[11059] = ~(layer2_outputs[7892]);
    assign outputs[11060] = (layer2_outputs[1953]) ^ (layer2_outputs[4837]);
    assign outputs[11061] = ~(layer2_outputs[9495]);
    assign outputs[11062] = layer2_outputs[8232];
    assign outputs[11063] = layer2_outputs[3841];
    assign outputs[11064] = layer2_outputs[12221];
    assign outputs[11065] = ~((layer2_outputs[2559]) ^ (layer2_outputs[3243]));
    assign outputs[11066] = (layer2_outputs[9326]) | (layer2_outputs[41]);
    assign outputs[11067] = ~(layer2_outputs[1006]);
    assign outputs[11068] = layer2_outputs[4941];
    assign outputs[11069] = ~(layer2_outputs[6990]);
    assign outputs[11070] = layer2_outputs[10351];
    assign outputs[11071] = ~(layer2_outputs[65]);
    assign outputs[11072] = ~(layer2_outputs[7426]);
    assign outputs[11073] = (layer2_outputs[4043]) ^ (layer2_outputs[11059]);
    assign outputs[11074] = layer2_outputs[9301];
    assign outputs[11075] = (layer2_outputs[5649]) ^ (layer2_outputs[3018]);
    assign outputs[11076] = ~(layer2_outputs[12512]);
    assign outputs[11077] = layer2_outputs[4612];
    assign outputs[11078] = layer2_outputs[4490];
    assign outputs[11079] = (layer2_outputs[2966]) & ~(layer2_outputs[9661]);
    assign outputs[11080] = layer2_outputs[1984];
    assign outputs[11081] = ~(layer2_outputs[6786]) | (layer2_outputs[10221]);
    assign outputs[11082] = ~(layer2_outputs[7211]);
    assign outputs[11083] = ~(layer2_outputs[10340]);
    assign outputs[11084] = ~(layer2_outputs[5741]);
    assign outputs[11085] = ~(layer2_outputs[5681]);
    assign outputs[11086] = ~(layer2_outputs[11338]);
    assign outputs[11087] = (layer2_outputs[7841]) | (layer2_outputs[2419]);
    assign outputs[11088] = ~(layer2_outputs[12395]) | (layer2_outputs[4604]);
    assign outputs[11089] = ~(layer2_outputs[724]);
    assign outputs[11090] = layer2_outputs[3223];
    assign outputs[11091] = layer2_outputs[5618];
    assign outputs[11092] = (layer2_outputs[426]) ^ (layer2_outputs[1091]);
    assign outputs[11093] = (layer2_outputs[7947]) ^ (layer2_outputs[5266]);
    assign outputs[11094] = (layer2_outputs[5200]) ^ (layer2_outputs[10355]);
    assign outputs[11095] = ~(layer2_outputs[76]);
    assign outputs[11096] = ~((layer2_outputs[9039]) ^ (layer2_outputs[4570]));
    assign outputs[11097] = layer2_outputs[3009];
    assign outputs[11098] = (layer2_outputs[12508]) | (layer2_outputs[4523]);
    assign outputs[11099] = layer2_outputs[3187];
    assign outputs[11100] = (layer2_outputs[2187]) | (layer2_outputs[3133]);
    assign outputs[11101] = layer2_outputs[2467];
    assign outputs[11102] = ~((layer2_outputs[7692]) ^ (layer2_outputs[9319]));
    assign outputs[11103] = ~((layer2_outputs[9186]) ^ (layer2_outputs[11394]));
    assign outputs[11104] = ~(layer2_outputs[4020]);
    assign outputs[11105] = ~(layer2_outputs[11681]);
    assign outputs[11106] = ~(layer2_outputs[5751]) | (layer2_outputs[8073]);
    assign outputs[11107] = ~(layer2_outputs[4761]) | (layer2_outputs[5495]);
    assign outputs[11108] = (layer2_outputs[11105]) ^ (layer2_outputs[7844]);
    assign outputs[11109] = layer2_outputs[1363];
    assign outputs[11110] = ~(layer2_outputs[10370]);
    assign outputs[11111] = layer2_outputs[2469];
    assign outputs[11112] = ~(layer2_outputs[4433]);
    assign outputs[11113] = ~((layer2_outputs[439]) ^ (layer2_outputs[2658]));
    assign outputs[11114] = layer2_outputs[2780];
    assign outputs[11115] = layer2_outputs[6958];
    assign outputs[11116] = ~(layer2_outputs[390]) | (layer2_outputs[12209]);
    assign outputs[11117] = ~(layer2_outputs[3445]) | (layer2_outputs[8025]);
    assign outputs[11118] = (layer2_outputs[10354]) ^ (layer2_outputs[11675]);
    assign outputs[11119] = ~(layer2_outputs[603]) | (layer2_outputs[1509]);
    assign outputs[11120] = layer2_outputs[10405];
    assign outputs[11121] = (layer2_outputs[11371]) ^ (layer2_outputs[12460]);
    assign outputs[11122] = layer2_outputs[1412];
    assign outputs[11123] = ~(layer2_outputs[6195]);
    assign outputs[11124] = layer2_outputs[2753];
    assign outputs[11125] = ~((layer2_outputs[11632]) ^ (layer2_outputs[1749]));
    assign outputs[11126] = ~(layer2_outputs[6699]) | (layer2_outputs[148]);
    assign outputs[11127] = layer2_outputs[4464];
    assign outputs[11128] = ~((layer2_outputs[388]) & (layer2_outputs[8141]));
    assign outputs[11129] = layer2_outputs[2264];
    assign outputs[11130] = (layer2_outputs[10227]) ^ (layer2_outputs[12149]);
    assign outputs[11131] = layer2_outputs[2694];
    assign outputs[11132] = ~(layer2_outputs[9312]);
    assign outputs[11133] = ~((layer2_outputs[808]) ^ (layer2_outputs[11790]));
    assign outputs[11134] = layer2_outputs[8795];
    assign outputs[11135] = (layer2_outputs[9933]) | (layer2_outputs[8458]);
    assign outputs[11136] = (layer2_outputs[1338]) | (layer2_outputs[7109]);
    assign outputs[11137] = ~(layer2_outputs[3990]) | (layer2_outputs[4794]);
    assign outputs[11138] = (layer2_outputs[2440]) ^ (layer2_outputs[5491]);
    assign outputs[11139] = ~((layer2_outputs[7941]) ^ (layer2_outputs[4611]));
    assign outputs[11140] = ~(layer2_outputs[10468]);
    assign outputs[11141] = ~(layer2_outputs[10826]) | (layer2_outputs[3686]);
    assign outputs[11142] = layer2_outputs[2697];
    assign outputs[11143] = (layer2_outputs[6973]) & (layer2_outputs[2947]);
    assign outputs[11144] = layer2_outputs[2155];
    assign outputs[11145] = layer2_outputs[7953];
    assign outputs[11146] = ~((layer2_outputs[1141]) ^ (layer2_outputs[12389]));
    assign outputs[11147] = ~((layer2_outputs[4382]) | (layer2_outputs[7442]));
    assign outputs[11148] = layer2_outputs[8869];
    assign outputs[11149] = layer2_outputs[12195];
    assign outputs[11150] = ~(layer2_outputs[5999]);
    assign outputs[11151] = layer2_outputs[8163];
    assign outputs[11152] = (layer2_outputs[114]) | (layer2_outputs[4121]);
    assign outputs[11153] = ~(layer2_outputs[735]);
    assign outputs[11154] = ~(layer2_outputs[4250]) | (layer2_outputs[1970]);
    assign outputs[11155] = ~(layer2_outputs[4988]);
    assign outputs[11156] = ~((layer2_outputs[11912]) | (layer2_outputs[3571]));
    assign outputs[11157] = (layer2_outputs[10864]) ^ (layer2_outputs[4287]);
    assign outputs[11158] = layer2_outputs[493];
    assign outputs[11159] = (layer2_outputs[2556]) & ~(layer2_outputs[10861]);
    assign outputs[11160] = layer2_outputs[7077];
    assign outputs[11161] = (layer2_outputs[9437]) ^ (layer2_outputs[8871]);
    assign outputs[11162] = layer2_outputs[13];
    assign outputs[11163] = layer2_outputs[10739];
    assign outputs[11164] = (layer2_outputs[8851]) ^ (layer2_outputs[1700]);
    assign outputs[11165] = ~((layer2_outputs[4374]) & (layer2_outputs[10288]));
    assign outputs[11166] = layer2_outputs[1420];
    assign outputs[11167] = (layer2_outputs[12319]) & ~(layer2_outputs[143]);
    assign outputs[11168] = ~((layer2_outputs[2945]) ^ (layer2_outputs[7540]));
    assign outputs[11169] = ~(layer2_outputs[8106]);
    assign outputs[11170] = layer2_outputs[2153];
    assign outputs[11171] = ~(layer2_outputs[7294]);
    assign outputs[11172] = layer2_outputs[10720];
    assign outputs[11173] = (layer2_outputs[4494]) | (layer2_outputs[6560]);
    assign outputs[11174] = ~(layer2_outputs[3399]);
    assign outputs[11175] = layer2_outputs[10466];
    assign outputs[11176] = (layer2_outputs[3757]) ^ (layer2_outputs[3260]);
    assign outputs[11177] = ~((layer2_outputs[938]) ^ (layer2_outputs[11163]));
    assign outputs[11178] = (layer2_outputs[5043]) ^ (layer2_outputs[5947]);
    assign outputs[11179] = layer2_outputs[5865];
    assign outputs[11180] = layer2_outputs[4380];
    assign outputs[11181] = (layer2_outputs[8431]) ^ (layer2_outputs[6128]);
    assign outputs[11182] = ~(layer2_outputs[12285]);
    assign outputs[11183] = (layer2_outputs[7497]) & ~(layer2_outputs[11672]);
    assign outputs[11184] = (layer2_outputs[1670]) & ~(layer2_outputs[5815]);
    assign outputs[11185] = (layer2_outputs[5968]) | (layer2_outputs[9521]);
    assign outputs[11186] = ~((layer2_outputs[8693]) ^ (layer2_outputs[12563]));
    assign outputs[11187] = ~((layer2_outputs[3806]) | (layer2_outputs[2240]));
    assign outputs[11188] = ~((layer2_outputs[118]) | (layer2_outputs[4791]));
    assign outputs[11189] = ~(layer2_outputs[11046]);
    assign outputs[11190] = ~(layer2_outputs[7221]) | (layer2_outputs[2597]);
    assign outputs[11191] = layer2_outputs[7693];
    assign outputs[11192] = (layer2_outputs[10793]) ^ (layer2_outputs[6376]);
    assign outputs[11193] = (layer2_outputs[6738]) & ~(layer2_outputs[12239]);
    assign outputs[11194] = ~(layer2_outputs[807]) | (layer2_outputs[11555]);
    assign outputs[11195] = (layer2_outputs[7578]) & (layer2_outputs[2717]);
    assign outputs[11196] = ~(layer2_outputs[4275]);
    assign outputs[11197] = (layer2_outputs[6459]) | (layer2_outputs[7145]);
    assign outputs[11198] = ~(layer2_outputs[666]);
    assign outputs[11199] = layer2_outputs[3647];
    assign outputs[11200] = (layer2_outputs[1321]) | (layer2_outputs[2785]);
    assign outputs[11201] = ~(layer2_outputs[11576]) | (layer2_outputs[12308]);
    assign outputs[11202] = ~((layer2_outputs[8441]) ^ (layer2_outputs[4165]));
    assign outputs[11203] = (layer2_outputs[7313]) ^ (layer2_outputs[6087]);
    assign outputs[11204] = ~((layer2_outputs[1498]) & (layer2_outputs[8085]));
    assign outputs[11205] = ~((layer2_outputs[10794]) ^ (layer2_outputs[2705]));
    assign outputs[11206] = (layer2_outputs[4247]) ^ (layer2_outputs[12295]);
    assign outputs[11207] = ~(layer2_outputs[249]);
    assign outputs[11208] = ~((layer2_outputs[12423]) ^ (layer2_outputs[1199]));
    assign outputs[11209] = layer2_outputs[1524];
    assign outputs[11210] = ~(layer2_outputs[8787]);
    assign outputs[11211] = ~((layer2_outputs[8429]) | (layer2_outputs[3352]));
    assign outputs[11212] = ~((layer2_outputs[11268]) ^ (layer2_outputs[258]));
    assign outputs[11213] = layer2_outputs[2151];
    assign outputs[11214] = ~(layer2_outputs[1322]);
    assign outputs[11215] = ~(layer2_outputs[6227]);
    assign outputs[11216] = ~((layer2_outputs[9882]) ^ (layer2_outputs[9221]));
    assign outputs[11217] = ~(layer2_outputs[384]);
    assign outputs[11218] = ~((layer2_outputs[12246]) | (layer2_outputs[12699]));
    assign outputs[11219] = ~(layer2_outputs[656]);
    assign outputs[11220] = ~(layer2_outputs[10597]);
    assign outputs[11221] = ~((layer2_outputs[5685]) ^ (layer2_outputs[12118]));
    assign outputs[11222] = 1'b1;
    assign outputs[11223] = ~(layer2_outputs[12173]);
    assign outputs[11224] = (layer2_outputs[7248]) | (layer2_outputs[663]);
    assign outputs[11225] = ~(layer2_outputs[10445]) | (layer2_outputs[37]);
    assign outputs[11226] = ~((layer2_outputs[2028]) & (layer2_outputs[5937]));
    assign outputs[11227] = ~((layer2_outputs[544]) ^ (layer2_outputs[7611]));
    assign outputs[11228] = layer2_outputs[1003];
    assign outputs[11229] = layer2_outputs[10940];
    assign outputs[11230] = ~((layer2_outputs[4073]) ^ (layer2_outputs[703]));
    assign outputs[11231] = (layer2_outputs[12535]) ^ (layer2_outputs[1595]);
    assign outputs[11232] = ~(layer2_outputs[9376]);
    assign outputs[11233] = (layer2_outputs[7122]) ^ (layer2_outputs[3011]);
    assign outputs[11234] = layer2_outputs[5930];
    assign outputs[11235] = ~(layer2_outputs[3784]);
    assign outputs[11236] = (layer2_outputs[6055]) ^ (layer2_outputs[4569]);
    assign outputs[11237] = layer2_outputs[1708];
    assign outputs[11238] = layer2_outputs[10654];
    assign outputs[11239] = ~((layer2_outputs[848]) & (layer2_outputs[11669]));
    assign outputs[11240] = ~((layer2_outputs[6430]) & (layer2_outputs[8198]));
    assign outputs[11241] = layer2_outputs[7165];
    assign outputs[11242] = layer2_outputs[12417];
    assign outputs[11243] = ~((layer2_outputs[9276]) | (layer2_outputs[2940]));
    assign outputs[11244] = ~((layer2_outputs[12700]) | (layer2_outputs[1888]));
    assign outputs[11245] = (layer2_outputs[12401]) ^ (layer2_outputs[3167]);
    assign outputs[11246] = ~(layer2_outputs[5757]);
    assign outputs[11247] = (layer2_outputs[3836]) ^ (layer2_outputs[4316]);
    assign outputs[11248] = (layer2_outputs[4859]) ^ (layer2_outputs[4648]);
    assign outputs[11249] = layer2_outputs[9867];
    assign outputs[11250] = (layer2_outputs[4168]) & ~(layer2_outputs[1769]);
    assign outputs[11251] = (layer2_outputs[11885]) | (layer2_outputs[10743]);
    assign outputs[11252] = layer2_outputs[9404];
    assign outputs[11253] = ~(layer2_outputs[2805]) | (layer2_outputs[3591]);
    assign outputs[11254] = ~((layer2_outputs[10456]) ^ (layer2_outputs[9486]));
    assign outputs[11255] = layer2_outputs[2682];
    assign outputs[11256] = ~(layer2_outputs[4680]);
    assign outputs[11257] = ~(layer2_outputs[7722]);
    assign outputs[11258] = (layer2_outputs[6908]) & (layer2_outputs[12534]);
    assign outputs[11259] = 1'b0;
    assign outputs[11260] = layer2_outputs[2882];
    assign outputs[11261] = ~((layer2_outputs[9487]) ^ (layer2_outputs[12558]));
    assign outputs[11262] = ~(layer2_outputs[1192]);
    assign outputs[11263] = (layer2_outputs[1433]) | (layer2_outputs[110]);
    assign outputs[11264] = layer2_outputs[6012];
    assign outputs[11265] = ~(layer2_outputs[3030]);
    assign outputs[11266] = (layer2_outputs[7677]) & ~(layer2_outputs[680]);
    assign outputs[11267] = ~((layer2_outputs[9748]) ^ (layer2_outputs[6896]));
    assign outputs[11268] = ~(layer2_outputs[12499]);
    assign outputs[11269] = ~((layer2_outputs[1235]) ^ (layer2_outputs[7440]));
    assign outputs[11270] = ~(layer2_outputs[10671]);
    assign outputs[11271] = ~((layer2_outputs[4956]) ^ (layer2_outputs[11874]));
    assign outputs[11272] = ~((layer2_outputs[11353]) ^ (layer2_outputs[12303]));
    assign outputs[11273] = layer2_outputs[9353];
    assign outputs[11274] = (layer2_outputs[11701]) ^ (layer2_outputs[10058]);
    assign outputs[11275] = (layer2_outputs[4362]) & ~(layer2_outputs[6368]);
    assign outputs[11276] = layer2_outputs[6592];
    assign outputs[11277] = (layer2_outputs[8105]) ^ (layer2_outputs[9720]);
    assign outputs[11278] = layer2_outputs[4609];
    assign outputs[11279] = ~(layer2_outputs[9519]) | (layer2_outputs[12324]);
    assign outputs[11280] = (layer2_outputs[6992]) & (layer2_outputs[4055]);
    assign outputs[11281] = ~((layer2_outputs[4565]) ^ (layer2_outputs[8755]));
    assign outputs[11282] = (layer2_outputs[8581]) ^ (layer2_outputs[5066]);
    assign outputs[11283] = ~(layer2_outputs[10261]);
    assign outputs[11284] = ~(layer2_outputs[294]);
    assign outputs[11285] = ~((layer2_outputs[7699]) & (layer2_outputs[4776]));
    assign outputs[11286] = ~(layer2_outputs[12679]);
    assign outputs[11287] = layer2_outputs[4922];
    assign outputs[11288] = ~(layer2_outputs[11058]);
    assign outputs[11289] = ~((layer2_outputs[9782]) ^ (layer2_outputs[10478]));
    assign outputs[11290] = ~(layer2_outputs[10807]);
    assign outputs[11291] = ~((layer2_outputs[12029]) ^ (layer2_outputs[903]));
    assign outputs[11292] = ~((layer2_outputs[1714]) ^ (layer2_outputs[11128]));
    assign outputs[11293] = ~(layer2_outputs[9401]);
    assign outputs[11294] = layer2_outputs[6772];
    assign outputs[11295] = layer2_outputs[4730];
    assign outputs[11296] = ~(layer2_outputs[4036]);
    assign outputs[11297] = (layer2_outputs[4102]) ^ (layer2_outputs[231]);
    assign outputs[11298] = layer2_outputs[389];
    assign outputs[11299] = layer2_outputs[11597];
    assign outputs[11300] = layer2_outputs[6092];
    assign outputs[11301] = ~((layer2_outputs[5031]) ^ (layer2_outputs[9005]));
    assign outputs[11302] = layer2_outputs[7798];
    assign outputs[11303] = ~((layer2_outputs[10418]) & (layer2_outputs[4011]));
    assign outputs[11304] = layer2_outputs[3455];
    assign outputs[11305] = (layer2_outputs[11409]) ^ (layer2_outputs[2281]);
    assign outputs[11306] = (layer2_outputs[1902]) ^ (layer2_outputs[2177]);
    assign outputs[11307] = (layer2_outputs[10612]) ^ (layer2_outputs[5546]);
    assign outputs[11308] = (layer2_outputs[3456]) ^ (layer2_outputs[2349]);
    assign outputs[11309] = ~((layer2_outputs[12603]) | (layer2_outputs[902]));
    assign outputs[11310] = ~((layer2_outputs[5064]) | (layer2_outputs[7817]));
    assign outputs[11311] = ~((layer2_outputs[6433]) | (layer2_outputs[11393]));
    assign outputs[11312] = (layer2_outputs[1224]) ^ (layer2_outputs[5294]);
    assign outputs[11313] = ~((layer2_outputs[9517]) ^ (layer2_outputs[252]));
    assign outputs[11314] = ~(layer2_outputs[6059]);
    assign outputs[11315] = layer2_outputs[5920];
    assign outputs[11316] = layer2_outputs[11966];
    assign outputs[11317] = ~(layer2_outputs[1225]) | (layer2_outputs[9941]);
    assign outputs[11318] = layer2_outputs[2321];
    assign outputs[11319] = ~(layer2_outputs[7164]);
    assign outputs[11320] = (layer2_outputs[11663]) ^ (layer2_outputs[10080]);
    assign outputs[11321] = ~(layer2_outputs[906]);
    assign outputs[11322] = layer2_outputs[12631];
    assign outputs[11323] = ~(layer2_outputs[2037]);
    assign outputs[11324] = ~((layer2_outputs[11898]) & (layer2_outputs[5370]));
    assign outputs[11325] = layer2_outputs[1242];
    assign outputs[11326] = (layer2_outputs[10562]) ^ (layer2_outputs[1897]);
    assign outputs[11327] = (layer2_outputs[2041]) ^ (layer2_outputs[7343]);
    assign outputs[11328] = ~((layer2_outputs[2739]) ^ (layer2_outputs[6363]));
    assign outputs[11329] = ~((layer2_outputs[10959]) & (layer2_outputs[7688]));
    assign outputs[11330] = layer2_outputs[4916];
    assign outputs[11331] = ~((layer2_outputs[5542]) ^ (layer2_outputs[6088]));
    assign outputs[11332] = (layer2_outputs[4507]) ^ (layer2_outputs[5306]);
    assign outputs[11333] = layer2_outputs[12031];
    assign outputs[11334] = layer2_outputs[6893];
    assign outputs[11335] = (layer2_outputs[3133]) & (layer2_outputs[1587]);
    assign outputs[11336] = (layer2_outputs[8452]) ^ (layer2_outputs[3661]);
    assign outputs[11337] = (layer2_outputs[9505]) | (layer2_outputs[4509]);
    assign outputs[11338] = ~((layer2_outputs[4575]) | (layer2_outputs[5612]));
    assign outputs[11339] = layer2_outputs[12113];
    assign outputs[11340] = layer2_outputs[970];
    assign outputs[11341] = ~((layer2_outputs[4226]) ^ (layer2_outputs[12156]));
    assign outputs[11342] = layer2_outputs[10732];
    assign outputs[11343] = ~((layer2_outputs[12785]) & (layer2_outputs[631]));
    assign outputs[11344] = ~((layer2_outputs[256]) ^ (layer2_outputs[5700]));
    assign outputs[11345] = layer2_outputs[9468];
    assign outputs[11346] = ~(layer2_outputs[167]);
    assign outputs[11347] = ~(layer2_outputs[8741]);
    assign outputs[11348] = ~((layer2_outputs[6054]) ^ (layer2_outputs[10613]));
    assign outputs[11349] = (layer2_outputs[6747]) & (layer2_outputs[8747]);
    assign outputs[11350] = (layer2_outputs[11481]) ^ (layer2_outputs[6652]);
    assign outputs[11351] = layer2_outputs[7684];
    assign outputs[11352] = layer2_outputs[11987];
    assign outputs[11353] = ~(layer2_outputs[2175]);
    assign outputs[11354] = (layer2_outputs[9715]) ^ (layer2_outputs[5004]);
    assign outputs[11355] = layer2_outputs[10985];
    assign outputs[11356] = ~((layer2_outputs[12370]) ^ (layer2_outputs[11994]));
    assign outputs[11357] = layer2_outputs[8150];
    assign outputs[11358] = layer2_outputs[7474];
    assign outputs[11359] = ~((layer2_outputs[9138]) & (layer2_outputs[8812]));
    assign outputs[11360] = ~((layer2_outputs[7156]) ^ (layer2_outputs[4519]));
    assign outputs[11361] = ~(layer2_outputs[7434]) | (layer2_outputs[2832]);
    assign outputs[11362] = layer2_outputs[7010];
    assign outputs[11363] = (layer2_outputs[4044]) ^ (layer2_outputs[4285]);
    assign outputs[11364] = layer2_outputs[12430];
    assign outputs[11365] = layer2_outputs[4857];
    assign outputs[11366] = ~(layer2_outputs[11268]);
    assign outputs[11367] = layer2_outputs[5627];
    assign outputs[11368] = (layer2_outputs[7722]) ^ (layer2_outputs[9182]);
    assign outputs[11369] = ~(layer2_outputs[9783]);
    assign outputs[11370] = (layer2_outputs[10132]) ^ (layer2_outputs[10130]);
    assign outputs[11371] = (layer2_outputs[1473]) | (layer2_outputs[7066]);
    assign outputs[11372] = ~((layer2_outputs[6232]) & (layer2_outputs[2775]));
    assign outputs[11373] = (layer2_outputs[9902]) ^ (layer2_outputs[5698]);
    assign outputs[11374] = (layer2_outputs[2428]) & ~(layer2_outputs[7128]);
    assign outputs[11375] = ~(layer2_outputs[11646]);
    assign outputs[11376] = ~((layer2_outputs[2330]) ^ (layer2_outputs[10638]));
    assign outputs[11377] = layer2_outputs[11115];
    assign outputs[11378] = ~(layer2_outputs[6175]);
    assign outputs[11379] = ~(layer2_outputs[2759]);
    assign outputs[11380] = (layer2_outputs[2631]) ^ (layer2_outputs[7044]);
    assign outputs[11381] = layer2_outputs[681];
    assign outputs[11382] = ~((layer2_outputs[9508]) ^ (layer2_outputs[9285]));
    assign outputs[11383] = layer2_outputs[3646];
    assign outputs[11384] = ~((layer2_outputs[12596]) ^ (layer2_outputs[6255]));
    assign outputs[11385] = ~((layer2_outputs[11256]) ^ (layer2_outputs[593]));
    assign outputs[11386] = layer2_outputs[9598];
    assign outputs[11387] = ~((layer2_outputs[1844]) ^ (layer2_outputs[12292]));
    assign outputs[11388] = (layer2_outputs[6479]) ^ (layer2_outputs[6272]);
    assign outputs[11389] = ~(layer2_outputs[11649]);
    assign outputs[11390] = (layer2_outputs[12227]) | (layer2_outputs[6899]);
    assign outputs[11391] = ~(layer2_outputs[10284]);
    assign outputs[11392] = ~(layer2_outputs[8186]);
    assign outputs[11393] = ~(layer2_outputs[4632]);
    assign outputs[11394] = ~(layer2_outputs[8928]) | (layer2_outputs[11852]);
    assign outputs[11395] = layer2_outputs[6261];
    assign outputs[11396] = layer2_outputs[5371];
    assign outputs[11397] = ~(layer2_outputs[11548]);
    assign outputs[11398] = (layer2_outputs[6221]) ^ (layer2_outputs[8709]);
    assign outputs[11399] = ~((layer2_outputs[8099]) & (layer2_outputs[12641]));
    assign outputs[11400] = ~(layer2_outputs[5239]) | (layer2_outputs[7472]);
    assign outputs[11401] = ~(layer2_outputs[12115]);
    assign outputs[11402] = ~(layer2_outputs[2070]);
    assign outputs[11403] = ~(layer2_outputs[1468]);
    assign outputs[11404] = ~(layer2_outputs[284]);
    assign outputs[11405] = layer2_outputs[1798];
    assign outputs[11406] = (layer2_outputs[6301]) ^ (layer2_outputs[11163]);
    assign outputs[11407] = (layer2_outputs[11089]) | (layer2_outputs[7190]);
    assign outputs[11408] = ~((layer2_outputs[2636]) ^ (layer2_outputs[11318]));
    assign outputs[11409] = (layer2_outputs[9350]) | (layer2_outputs[5464]);
    assign outputs[11410] = layer2_outputs[9854];
    assign outputs[11411] = ~((layer2_outputs[5419]) ^ (layer2_outputs[2499]));
    assign outputs[11412] = (layer2_outputs[5825]) ^ (layer2_outputs[5443]);
    assign outputs[11413] = ~(layer2_outputs[7478]) | (layer2_outputs[2053]);
    assign outputs[11414] = (layer2_outputs[2015]) & (layer2_outputs[3345]);
    assign outputs[11415] = layer2_outputs[4043];
    assign outputs[11416] = ~(layer2_outputs[9096]);
    assign outputs[11417] = layer2_outputs[7349];
    assign outputs[11418] = layer2_outputs[1254];
    assign outputs[11419] = ~(layer2_outputs[10790]) | (layer2_outputs[5841]);
    assign outputs[11420] = ~((layer2_outputs[10025]) ^ (layer2_outputs[11579]));
    assign outputs[11421] = layer2_outputs[2330];
    assign outputs[11422] = ~(layer2_outputs[1854]);
    assign outputs[11423] = ~((layer2_outputs[6114]) & (layer2_outputs[4037]));
    assign outputs[11424] = layer2_outputs[10718];
    assign outputs[11425] = ~((layer2_outputs[6126]) ^ (layer2_outputs[6689]));
    assign outputs[11426] = ~(layer2_outputs[9924]) | (layer2_outputs[9]);
    assign outputs[11427] = layer2_outputs[11327];
    assign outputs[11428] = ~((layer2_outputs[3991]) ^ (layer2_outputs[6543]));
    assign outputs[11429] = ~((layer2_outputs[8799]) & (layer2_outputs[1732]));
    assign outputs[11430] = ~((layer2_outputs[6545]) ^ (layer2_outputs[10900]));
    assign outputs[11431] = ~(layer2_outputs[7831]) | (layer2_outputs[6115]);
    assign outputs[11432] = ~((layer2_outputs[10465]) ^ (layer2_outputs[10492]));
    assign outputs[11433] = layer2_outputs[7828];
    assign outputs[11434] = ~((layer2_outputs[1988]) ^ (layer2_outputs[11534]));
    assign outputs[11435] = ~(layer2_outputs[2474]);
    assign outputs[11436] = (layer2_outputs[12358]) & (layer2_outputs[6730]);
    assign outputs[11437] = ~(layer2_outputs[5179]);
    assign outputs[11438] = (layer2_outputs[11274]) ^ (layer2_outputs[3090]);
    assign outputs[11439] = layer2_outputs[2076];
    assign outputs[11440] = ~(layer2_outputs[3081]) | (layer2_outputs[4726]);
    assign outputs[11441] = layer2_outputs[9923];
    assign outputs[11442] = ~(layer2_outputs[7617]) | (layer2_outputs[2828]);
    assign outputs[11443] = (layer2_outputs[7966]) ^ (layer2_outputs[3470]);
    assign outputs[11444] = layer2_outputs[2808];
    assign outputs[11445] = ~(layer2_outputs[6129]);
    assign outputs[11446] = ~((layer2_outputs[9679]) ^ (layer2_outputs[4213]));
    assign outputs[11447] = (layer2_outputs[2085]) | (layer2_outputs[11423]);
    assign outputs[11448] = ~(layer2_outputs[2161]);
    assign outputs[11449] = layer2_outputs[6436];
    assign outputs[11450] = (layer2_outputs[264]) ^ (layer2_outputs[8923]);
    assign outputs[11451] = (layer2_outputs[7347]) & (layer2_outputs[6636]);
    assign outputs[11452] = ~((layer2_outputs[1203]) ^ (layer2_outputs[7889]));
    assign outputs[11453] = ~(layer2_outputs[10233]);
    assign outputs[11454] = ~((layer2_outputs[128]) ^ (layer2_outputs[8909]));
    assign outputs[11455] = ~((layer2_outputs[12493]) ^ (layer2_outputs[2732]));
    assign outputs[11456] = ~(layer2_outputs[12094]);
    assign outputs[11457] = (layer2_outputs[3773]) ^ (layer2_outputs[767]);
    assign outputs[11458] = ~((layer2_outputs[9925]) ^ (layer2_outputs[1037]));
    assign outputs[11459] = ~((layer2_outputs[1671]) & (layer2_outputs[9511]));
    assign outputs[11460] = layer2_outputs[8323];
    assign outputs[11461] = ~(layer2_outputs[2394]) | (layer2_outputs[1471]);
    assign outputs[11462] = ~((layer2_outputs[5118]) ^ (layer2_outputs[10178]));
    assign outputs[11463] = ~(layer2_outputs[12367]) | (layer2_outputs[1859]);
    assign outputs[11464] = ~(layer2_outputs[11849]) | (layer2_outputs[2873]);
    assign outputs[11465] = (layer2_outputs[4751]) ^ (layer2_outputs[6678]);
    assign outputs[11466] = layer2_outputs[8856];
    assign outputs[11467] = ~((layer2_outputs[12718]) | (layer2_outputs[3498]));
    assign outputs[11468] = ~((layer2_outputs[7661]) ^ (layer2_outputs[2249]));
    assign outputs[11469] = (layer2_outputs[42]) ^ (layer2_outputs[2820]);
    assign outputs[11470] = ~(layer2_outputs[6412]);
    assign outputs[11471] = (layer2_outputs[11206]) ^ (layer2_outputs[2431]);
    assign outputs[11472] = (layer2_outputs[5450]) | (layer2_outputs[11662]);
    assign outputs[11473] = (layer2_outputs[11532]) ^ (layer2_outputs[12070]);
    assign outputs[11474] = ~((layer2_outputs[11882]) ^ (layer2_outputs[1393]));
    assign outputs[11475] = (layer2_outputs[7843]) ^ (layer2_outputs[3663]);
    assign outputs[11476] = (layer2_outputs[16]) ^ (layer2_outputs[5453]);
    assign outputs[11477] = (layer2_outputs[1161]) | (layer2_outputs[9010]);
    assign outputs[11478] = (layer2_outputs[12343]) ^ (layer2_outputs[8263]);
    assign outputs[11479] = layer2_outputs[6956];
    assign outputs[11480] = (layer2_outputs[10306]) ^ (layer2_outputs[2324]);
    assign outputs[11481] = (layer2_outputs[2418]) ^ (layer2_outputs[8181]);
    assign outputs[11482] = ~(layer2_outputs[8579]);
    assign outputs[11483] = layer2_outputs[7372];
    assign outputs[11484] = ~(layer2_outputs[4894]);
    assign outputs[11485] = layer2_outputs[3841];
    assign outputs[11486] = layer2_outputs[5308];
    assign outputs[11487] = layer2_outputs[170];
    assign outputs[11488] = (layer2_outputs[9944]) & (layer2_outputs[9124]);
    assign outputs[11489] = ~(layer2_outputs[2907]);
    assign outputs[11490] = ~(layer2_outputs[10493]);
    assign outputs[11491] = ~(layer2_outputs[9430]);
    assign outputs[11492] = (layer2_outputs[11671]) ^ (layer2_outputs[10667]);
    assign outputs[11493] = ~((layer2_outputs[6858]) ^ (layer2_outputs[5175]));
    assign outputs[11494] = ~(layer2_outputs[9269]);
    assign outputs[11495] = layer2_outputs[2935];
    assign outputs[11496] = (layer2_outputs[628]) ^ (layer2_outputs[7070]);
    assign outputs[11497] = (layer2_outputs[12321]) ^ (layer2_outputs[12538]);
    assign outputs[11498] = layer2_outputs[8449];
    assign outputs[11499] = ~(layer2_outputs[2803]);
    assign outputs[11500] = layer2_outputs[5015];
    assign outputs[11501] = ~(layer2_outputs[11741]);
    assign outputs[11502] = layer2_outputs[4834];
    assign outputs[11503] = ~(layer2_outputs[8902]);
    assign outputs[11504] = ~(layer2_outputs[3095]);
    assign outputs[11505] = ~((layer2_outputs[416]) ^ (layer2_outputs[376]));
    assign outputs[11506] = ~(layer2_outputs[6186]);
    assign outputs[11507] = ~(layer2_outputs[4522]);
    assign outputs[11508] = ~(layer2_outputs[8791]) | (layer2_outputs[3176]);
    assign outputs[11509] = (layer2_outputs[2719]) ^ (layer2_outputs[2915]);
    assign outputs[11510] = ~(layer2_outputs[1078]) | (layer2_outputs[6577]);
    assign outputs[11511] = (layer2_outputs[1131]) & ~(layer2_outputs[5146]);
    assign outputs[11512] = ~(layer2_outputs[9534]) | (layer2_outputs[4081]);
    assign outputs[11513] = ~(layer2_outputs[9927]) | (layer2_outputs[11125]);
    assign outputs[11514] = layer2_outputs[11590];
    assign outputs[11515] = ~(layer2_outputs[6932]);
    assign outputs[11516] = ~(layer2_outputs[1715]);
    assign outputs[11517] = ~((layer2_outputs[10691]) | (layer2_outputs[1767]));
    assign outputs[11518] = layer2_outputs[1852];
    assign outputs[11519] = (layer2_outputs[11541]) ^ (layer2_outputs[2042]);
    assign outputs[11520] = layer2_outputs[6806];
    assign outputs[11521] = layer2_outputs[12021];
    assign outputs[11522] = ~((layer2_outputs[5126]) ^ (layer2_outputs[5861]));
    assign outputs[11523] = (layer2_outputs[8478]) ^ (layer2_outputs[6598]);
    assign outputs[11524] = (layer2_outputs[12462]) & ~(layer2_outputs[6424]);
    assign outputs[11525] = (layer2_outputs[7384]) ^ (layer2_outputs[2038]);
    assign outputs[11526] = layer2_outputs[10903];
    assign outputs[11527] = ~(layer2_outputs[12396]);
    assign outputs[11528] = (layer2_outputs[3590]) & (layer2_outputs[12198]);
    assign outputs[11529] = ~(layer2_outputs[2035]);
    assign outputs[11530] = (layer2_outputs[4596]) | (layer2_outputs[11545]);
    assign outputs[11531] = ~((layer2_outputs[9489]) ^ (layer2_outputs[4178]));
    assign outputs[11532] = ~(layer2_outputs[6424]);
    assign outputs[11533] = layer2_outputs[5383];
    assign outputs[11534] = (layer2_outputs[1869]) ^ (layer2_outputs[12632]);
    assign outputs[11535] = ~(layer2_outputs[5198]);
    assign outputs[11536] = ~((layer2_outputs[642]) ^ (layer2_outputs[12075]));
    assign outputs[11537] = ~((layer2_outputs[8258]) ^ (layer2_outputs[4228]));
    assign outputs[11538] = ~(layer2_outputs[10151]);
    assign outputs[11539] = ~(layer2_outputs[6109]) | (layer2_outputs[6600]);
    assign outputs[11540] = (layer2_outputs[3589]) & ~(layer2_outputs[1401]);
    assign outputs[11541] = layer2_outputs[1900];
    assign outputs[11542] = layer2_outputs[895];
    assign outputs[11543] = layer2_outputs[936];
    assign outputs[11544] = ~((layer2_outputs[12485]) ^ (layer2_outputs[4149]));
    assign outputs[11545] = ~(layer2_outputs[380]);
    assign outputs[11546] = layer2_outputs[5220];
    assign outputs[11547] = (layer2_outputs[1374]) ^ (layer2_outputs[8545]);
    assign outputs[11548] = ~(layer2_outputs[190]);
    assign outputs[11549] = ~((layer2_outputs[7331]) | (layer2_outputs[4270]));
    assign outputs[11550] = ~(layer2_outputs[11492]);
    assign outputs[11551] = ~(layer2_outputs[8655]);
    assign outputs[11552] = layer2_outputs[10682];
    assign outputs[11553] = ~(layer2_outputs[12276]);
    assign outputs[11554] = ~(layer2_outputs[3717]);
    assign outputs[11555] = layer2_outputs[7778];
    assign outputs[11556] = ~(layer2_outputs[10378]);
    assign outputs[11557] = (layer2_outputs[8418]) & ~(layer2_outputs[2137]);
    assign outputs[11558] = ~(layer2_outputs[3035]);
    assign outputs[11559] = ~(layer2_outputs[6693]);
    assign outputs[11560] = layer2_outputs[12514];
    assign outputs[11561] = ~(layer2_outputs[10799]);
    assign outputs[11562] = ~((layer2_outputs[3454]) ^ (layer2_outputs[4021]));
    assign outputs[11563] = ~(layer2_outputs[10253]);
    assign outputs[11564] = layer2_outputs[3127];
    assign outputs[11565] = ~(layer2_outputs[12784]);
    assign outputs[11566] = (layer2_outputs[1345]) ^ (layer2_outputs[9985]);
    assign outputs[11567] = ~(layer2_outputs[4243]);
    assign outputs[11568] = ~((layer2_outputs[5337]) ^ (layer2_outputs[8987]));
    assign outputs[11569] = layer2_outputs[4370];
    assign outputs[11570] = layer2_outputs[387];
    assign outputs[11571] = layer2_outputs[9468];
    assign outputs[11572] = layer2_outputs[7485];
    assign outputs[11573] = ~((layer2_outputs[11457]) & (layer2_outputs[4140]));
    assign outputs[11574] = layer2_outputs[4263];
    assign outputs[11575] = (layer2_outputs[350]) & ~(layer2_outputs[5879]);
    assign outputs[11576] = ~(layer2_outputs[3630]);
    assign outputs[11577] = layer2_outputs[5622];
    assign outputs[11578] = layer2_outputs[568];
    assign outputs[11579] = layer2_outputs[3801];
    assign outputs[11580] = ~(layer2_outputs[3782]);
    assign outputs[11581] = (layer2_outputs[9248]) ^ (layer2_outputs[12608]);
    assign outputs[11582] = ~(layer2_outputs[12025]) | (layer2_outputs[10579]);
    assign outputs[11583] = layer2_outputs[3772];
    assign outputs[11584] = (layer2_outputs[6243]) ^ (layer2_outputs[324]);
    assign outputs[11585] = ~(layer2_outputs[2737]);
    assign outputs[11586] = ~(layer2_outputs[984]);
    assign outputs[11587] = ~(layer2_outputs[11445]);
    assign outputs[11588] = ~(layer2_outputs[4406]);
    assign outputs[11589] = ~(layer2_outputs[3422]);
    assign outputs[11590] = ~((layer2_outputs[5373]) & (layer2_outputs[11375]));
    assign outputs[11591] = ~(layer2_outputs[1057]);
    assign outputs[11592] = (layer2_outputs[6710]) ^ (layer2_outputs[2955]);
    assign outputs[11593] = ~((layer2_outputs[24]) ^ (layer2_outputs[9081]));
    assign outputs[11594] = ~(layer2_outputs[12611]);
    assign outputs[11595] = (layer2_outputs[11794]) | (layer2_outputs[12277]);
    assign outputs[11596] = ~(layer2_outputs[3200]) | (layer2_outputs[6136]);
    assign outputs[11597] = ~(layer2_outputs[9869]);
    assign outputs[11598] = layer2_outputs[12254];
    assign outputs[11599] = layer2_outputs[10414];
    assign outputs[11600] = (layer2_outputs[202]) & (layer2_outputs[4182]);
    assign outputs[11601] = layer2_outputs[776];
    assign outputs[11602] = ~(layer2_outputs[7968]);
    assign outputs[11603] = layer2_outputs[8777];
    assign outputs[11604] = layer2_outputs[7231];
    assign outputs[11605] = ~((layer2_outputs[4441]) & (layer2_outputs[3320]));
    assign outputs[11606] = (layer2_outputs[8715]) ^ (layer2_outputs[2877]);
    assign outputs[11607] = layer2_outputs[7965];
    assign outputs[11608] = (layer2_outputs[447]) ^ (layer2_outputs[5607]);
    assign outputs[11609] = ~(layer2_outputs[11841]) | (layer2_outputs[7032]);
    assign outputs[11610] = ~((layer2_outputs[2336]) | (layer2_outputs[11177]));
    assign outputs[11611] = ~(layer2_outputs[2078]) | (layer2_outputs[8617]);
    assign outputs[11612] = layer2_outputs[260];
    assign outputs[11613] = layer2_outputs[2456];
    assign outputs[11614] = ~(layer2_outputs[2846]);
    assign outputs[11615] = layer2_outputs[3325];
    assign outputs[11616] = ~(layer2_outputs[972]);
    assign outputs[11617] = (layer2_outputs[2655]) & ~(layer2_outputs[1753]);
    assign outputs[11618] = (layer2_outputs[12610]) ^ (layer2_outputs[1136]);
    assign outputs[11619] = (layer2_outputs[4307]) ^ (layer2_outputs[11417]);
    assign outputs[11620] = ~(layer2_outputs[6903]);
    assign outputs[11621] = layer2_outputs[1812];
    assign outputs[11622] = (layer2_outputs[9417]) & ~(layer2_outputs[7443]);
    assign outputs[11623] = (layer2_outputs[4420]) & ~(layer2_outputs[8778]);
    assign outputs[11624] = (layer2_outputs[5271]) ^ (layer2_outputs[6927]);
    assign outputs[11625] = ~((layer2_outputs[8696]) ^ (layer2_outputs[5492]));
    assign outputs[11626] = ~((layer2_outputs[10456]) ^ (layer2_outputs[9692]));
    assign outputs[11627] = ~((layer2_outputs[4061]) | (layer2_outputs[7417]));
    assign outputs[11628] = ~(layer2_outputs[6467]) | (layer2_outputs[3375]);
    assign outputs[11629] = (layer2_outputs[1011]) & (layer2_outputs[5872]);
    assign outputs[11630] = ~(layer2_outputs[12181]) | (layer2_outputs[5620]);
    assign outputs[11631] = ~(layer2_outputs[8550]);
    assign outputs[11632] = layer2_outputs[6814];
    assign outputs[11633] = ~((layer2_outputs[12633]) ^ (layer2_outputs[5116]));
    assign outputs[11634] = ~(layer2_outputs[8892]);
    assign outputs[11635] = (layer2_outputs[3557]) & ~(layer2_outputs[12664]);
    assign outputs[11636] = ~((layer2_outputs[5139]) ^ (layer2_outputs[7739]));
    assign outputs[11637] = (layer2_outputs[1218]) ^ (layer2_outputs[3379]);
    assign outputs[11638] = ~((layer2_outputs[2346]) ^ (layer2_outputs[4469]));
    assign outputs[11639] = ~(layer2_outputs[5566]);
    assign outputs[11640] = layer2_outputs[6429];
    assign outputs[11641] = (layer2_outputs[12155]) ^ (layer2_outputs[4196]);
    assign outputs[11642] = ~((layer2_outputs[8205]) ^ (layer2_outputs[971]));
    assign outputs[11643] = ~(layer2_outputs[9215]);
    assign outputs[11644] = ~((layer2_outputs[6410]) ^ (layer2_outputs[4286]));
    assign outputs[11645] = ~(layer2_outputs[754]) | (layer2_outputs[7223]);
    assign outputs[11646] = (layer2_outputs[11389]) & ~(layer2_outputs[10879]);
    assign outputs[11647] = (layer2_outputs[3835]) & (layer2_outputs[8669]);
    assign outputs[11648] = layer2_outputs[9620];
    assign outputs[11649] = layer2_outputs[1723];
    assign outputs[11650] = ~(layer2_outputs[2940]);
    assign outputs[11651] = layer2_outputs[2985];
    assign outputs[11652] = ~(layer2_outputs[8647]);
    assign outputs[11653] = ~(layer2_outputs[2001]);
    assign outputs[11654] = ~((layer2_outputs[915]) ^ (layer2_outputs[2579]));
    assign outputs[11655] = ~((layer2_outputs[6138]) | (layer2_outputs[2475]));
    assign outputs[11656] = ~(layer2_outputs[9576]);
    assign outputs[11657] = ~(layer2_outputs[11860]) | (layer2_outputs[11819]);
    assign outputs[11658] = (layer2_outputs[2080]) ^ (layer2_outputs[11517]);
    assign outputs[11659] = ~(layer2_outputs[4918]);
    assign outputs[11660] = ~(layer2_outputs[11499]);
    assign outputs[11661] = layer2_outputs[10234];
    assign outputs[11662] = layer2_outputs[4204];
    assign outputs[11663] = (layer2_outputs[4206]) ^ (layer2_outputs[7638]);
    assign outputs[11664] = layer2_outputs[5460];
    assign outputs[11665] = ~(layer2_outputs[4078]) | (layer2_outputs[5153]);
    assign outputs[11666] = ~(layer2_outputs[7053]);
    assign outputs[11667] = ~(layer2_outputs[12190]);
    assign outputs[11668] = ~((layer2_outputs[11221]) ^ (layer2_outputs[11077]));
    assign outputs[11669] = ~((layer2_outputs[4477]) ^ (layer2_outputs[10998]));
    assign outputs[11670] = layer2_outputs[7767];
    assign outputs[11671] = ~((layer2_outputs[1397]) ^ (layer2_outputs[6171]));
    assign outputs[11672] = ~(layer2_outputs[1234]);
    assign outputs[11673] = layer2_outputs[10246];
    assign outputs[11674] = layer2_outputs[3431];
    assign outputs[11675] = ~(layer2_outputs[4048]);
    assign outputs[11676] = layer2_outputs[5383];
    assign outputs[11677] = (layer2_outputs[8834]) & (layer2_outputs[3409]);
    assign outputs[11678] = layer2_outputs[12081];
    assign outputs[11679] = (layer2_outputs[3608]) ^ (layer2_outputs[998]);
    assign outputs[11680] = ~(layer2_outputs[9132]);
    assign outputs[11681] = ~((layer2_outputs[8650]) ^ (layer2_outputs[3764]));
    assign outputs[11682] = layer2_outputs[4998];
    assign outputs[11683] = ~(layer2_outputs[11689]);
    assign outputs[11684] = (layer2_outputs[6160]) | (layer2_outputs[4718]);
    assign outputs[11685] = layer2_outputs[10724];
    assign outputs[11686] = ~((layer2_outputs[3386]) ^ (layer2_outputs[148]));
    assign outputs[11687] = ~(layer2_outputs[5677]);
    assign outputs[11688] = ~((layer2_outputs[4414]) & (layer2_outputs[2286]));
    assign outputs[11689] = layer2_outputs[2173];
    assign outputs[11690] = (layer2_outputs[2926]) | (layer2_outputs[7512]);
    assign outputs[11691] = layer2_outputs[9518];
    assign outputs[11692] = ~(layer2_outputs[73]);
    assign outputs[11693] = (layer2_outputs[7803]) & ~(layer2_outputs[11766]);
    assign outputs[11694] = layer2_outputs[7540];
    assign outputs[11695] = layer2_outputs[7936];
    assign outputs[11696] = ~((layer2_outputs[10868]) & (layer2_outputs[6152]));
    assign outputs[11697] = ~(layer2_outputs[4553]);
    assign outputs[11698] = layer2_outputs[1240];
    assign outputs[11699] = ~(layer2_outputs[3109]);
    assign outputs[11700] = (layer2_outputs[6200]) ^ (layer2_outputs[8480]);
    assign outputs[11701] = ~((layer2_outputs[2819]) ^ (layer2_outputs[8277]));
    assign outputs[11702] = ~(layer2_outputs[10181]);
    assign outputs[11703] = layer2_outputs[12043];
    assign outputs[11704] = layer2_outputs[3003];
    assign outputs[11705] = ~(layer2_outputs[5531]);
    assign outputs[11706] = ~(layer2_outputs[9873]);
    assign outputs[11707] = ~(layer2_outputs[1925]);
    assign outputs[11708] = (layer2_outputs[6720]) | (layer2_outputs[813]);
    assign outputs[11709] = (layer2_outputs[5180]) & (layer2_outputs[7767]);
    assign outputs[11710] = ~(layer2_outputs[10254]);
    assign outputs[11711] = ~(layer2_outputs[5961]);
    assign outputs[11712] = (layer2_outputs[1463]) ^ (layer2_outputs[5904]);
    assign outputs[11713] = layer2_outputs[11783];
    assign outputs[11714] = (layer2_outputs[10747]) & ~(layer2_outputs[3338]);
    assign outputs[11715] = ~((layer2_outputs[8574]) ^ (layer2_outputs[8855]));
    assign outputs[11716] = layer2_outputs[4775];
    assign outputs[11717] = layer2_outputs[533];
    assign outputs[11718] = ~(layer2_outputs[8294]);
    assign outputs[11719] = layer2_outputs[7707];
    assign outputs[11720] = layer2_outputs[12794];
    assign outputs[11721] = ~(layer2_outputs[473]);
    assign outputs[11722] = (layer2_outputs[9617]) & ~(layer2_outputs[12154]);
    assign outputs[11723] = ~(layer2_outputs[7711]);
    assign outputs[11724] = ~(layer2_outputs[8415]);
    assign outputs[11725] = layer2_outputs[2961];
    assign outputs[11726] = (layer2_outputs[3567]) ^ (layer2_outputs[6079]);
    assign outputs[11727] = ~(layer2_outputs[9252]);
    assign outputs[11728] = ~((layer2_outputs[3584]) | (layer2_outputs[1548]));
    assign outputs[11729] = (layer2_outputs[8654]) ^ (layer2_outputs[2881]);
    assign outputs[11730] = ~((layer2_outputs[4893]) | (layer2_outputs[10542]));
    assign outputs[11731] = (layer2_outputs[8090]) ^ (layer2_outputs[1826]);
    assign outputs[11732] = ~(layer2_outputs[3423]);
    assign outputs[11733] = layer2_outputs[3995];
    assign outputs[11734] = ~((layer2_outputs[3813]) & (layer2_outputs[9149]));
    assign outputs[11735] = ~((layer2_outputs[11489]) & (layer2_outputs[8571]));
    assign outputs[11736] = (layer2_outputs[10963]) ^ (layer2_outputs[5332]);
    assign outputs[11737] = ~(layer2_outputs[6155]);
    assign outputs[11738] = layer2_outputs[1170];
    assign outputs[11739] = (layer2_outputs[6288]) & ~(layer2_outputs[923]);
    assign outputs[11740] = ~(layer2_outputs[11440]);
    assign outputs[11741] = (layer2_outputs[8328]) ^ (layer2_outputs[6651]);
    assign outputs[11742] = ~((layer2_outputs[9210]) & (layer2_outputs[6340]));
    assign outputs[11743] = layer2_outputs[6045];
    assign outputs[11744] = layer2_outputs[7576];
    assign outputs[11745] = ~(layer2_outputs[3946]);
    assign outputs[11746] = ~(layer2_outputs[9932]);
    assign outputs[11747] = (layer2_outputs[5514]) ^ (layer2_outputs[4328]);
    assign outputs[11748] = (layer2_outputs[9628]) ^ (layer2_outputs[7459]);
    assign outputs[11749] = ~((layer2_outputs[6841]) ^ (layer2_outputs[2287]));
    assign outputs[11750] = ~(layer2_outputs[10671]);
    assign outputs[11751] = (layer2_outputs[7729]) & ~(layer2_outputs[8504]);
    assign outputs[11752] = ~(layer2_outputs[11430]) | (layer2_outputs[4571]);
    assign outputs[11753] = ~(layer2_outputs[322]);
    assign outputs[11754] = ~(layer2_outputs[55]);
    assign outputs[11755] = ~(layer2_outputs[573]);
    assign outputs[11756] = ~(layer2_outputs[6903]);
    assign outputs[11757] = layer2_outputs[7013];
    assign outputs[11758] = (layer2_outputs[10668]) ^ (layer2_outputs[9956]);
    assign outputs[11759] = layer2_outputs[6453];
    assign outputs[11760] = (layer2_outputs[1899]) ^ (layer2_outputs[1851]);
    assign outputs[11761] = ~(layer2_outputs[6558]);
    assign outputs[11762] = layer2_outputs[6099];
    assign outputs[11763] = ~(layer2_outputs[10205]);
    assign outputs[11764] = ~((layer2_outputs[8283]) ^ (layer2_outputs[3310]));
    assign outputs[11765] = layer2_outputs[179];
    assign outputs[11766] = layer2_outputs[6690];
    assign outputs[11767] = ~(layer2_outputs[9079]) | (layer2_outputs[3641]);
    assign outputs[11768] = ~((layer2_outputs[10194]) & (layer2_outputs[1351]));
    assign outputs[11769] = ~(layer2_outputs[1022]);
    assign outputs[11770] = ~(layer2_outputs[5806]) | (layer2_outputs[10922]);
    assign outputs[11771] = layer2_outputs[676];
    assign outputs[11772] = (layer2_outputs[7642]) ^ (layer2_outputs[11611]);
    assign outputs[11773] = (layer2_outputs[7618]) ^ (layer2_outputs[1582]);
    assign outputs[11774] = layer2_outputs[7187];
    assign outputs[11775] = (layer2_outputs[4994]) & (layer2_outputs[3408]);
    assign outputs[11776] = ~((layer2_outputs[9429]) ^ (layer2_outputs[2297]));
    assign outputs[11777] = (layer2_outputs[1795]) & (layer2_outputs[10414]);
    assign outputs[11778] = ~(layer2_outputs[1766]);
    assign outputs[11779] = (layer2_outputs[1640]) ^ (layer2_outputs[3281]);
    assign outputs[11780] = (layer2_outputs[10529]) ^ (layer2_outputs[12536]);
    assign outputs[11781] = layer2_outputs[8610];
    assign outputs[11782] = layer2_outputs[4272];
    assign outputs[11783] = ~((layer2_outputs[7676]) ^ (layer2_outputs[1634]));
    assign outputs[11784] = layer2_outputs[7360];
    assign outputs[11785] = (layer2_outputs[3196]) ^ (layer2_outputs[4640]);
    assign outputs[11786] = ~(layer2_outputs[5488]) | (layer2_outputs[9994]);
    assign outputs[11787] = (layer2_outputs[862]) ^ (layer2_outputs[5837]);
    assign outputs[11788] = ~(layer2_outputs[10054]) | (layer2_outputs[7659]);
    assign outputs[11789] = ~(layer2_outputs[492]);
    assign outputs[11790] = (layer2_outputs[11910]) & ~(layer2_outputs[6427]);
    assign outputs[11791] = (layer2_outputs[8079]) ^ (layer2_outputs[8975]);
    assign outputs[11792] = layer2_outputs[11730];
    assign outputs[11793] = (layer2_outputs[6499]) ^ (layer2_outputs[1374]);
    assign outputs[11794] = ~(layer2_outputs[6826]);
    assign outputs[11795] = ~(layer2_outputs[5283]);
    assign outputs[11796] = ~(layer2_outputs[7348]) | (layer2_outputs[9267]);
    assign outputs[11797] = ~(layer2_outputs[4462]);
    assign outputs[11798] = ~(layer2_outputs[9000]);
    assign outputs[11799] = ~(layer2_outputs[7851]);
    assign outputs[11800] = ~((layer2_outputs[3796]) ^ (layer2_outputs[11854]));
    assign outputs[11801] = ~(layer2_outputs[629]);
    assign outputs[11802] = layer2_outputs[3680];
    assign outputs[11803] = layer2_outputs[846];
    assign outputs[11804] = layer2_outputs[6736];
    assign outputs[11805] = ~((layer2_outputs[2644]) ^ (layer2_outputs[2176]));
    assign outputs[11806] = ~(layer2_outputs[1378]) | (layer2_outputs[7656]);
    assign outputs[11807] = ~(layer2_outputs[1578]);
    assign outputs[11808] = (layer2_outputs[2353]) & (layer2_outputs[2224]);
    assign outputs[11809] = ~((layer2_outputs[3696]) ^ (layer2_outputs[6295]));
    assign outputs[11810] = ~(layer2_outputs[3160]);
    assign outputs[11811] = layer2_outputs[11782];
    assign outputs[11812] = ~((layer2_outputs[1301]) ^ (layer2_outputs[11573]));
    assign outputs[11813] = (layer2_outputs[11739]) & (layer2_outputs[9131]);
    assign outputs[11814] = (layer2_outputs[11425]) & ~(layer2_outputs[684]);
    assign outputs[11815] = layer2_outputs[7884];
    assign outputs[11816] = layer2_outputs[2662];
    assign outputs[11817] = layer2_outputs[11022];
    assign outputs[11818] = ~((layer2_outputs[6476]) | (layer2_outputs[4059]));
    assign outputs[11819] = ~(layer2_outputs[9699]);
    assign outputs[11820] = ~(layer2_outputs[573]);
    assign outputs[11821] = ~((layer2_outputs[6629]) ^ (layer2_outputs[1375]));
    assign outputs[11822] = ~(layer2_outputs[9898]);
    assign outputs[11823] = (layer2_outputs[252]) ^ (layer2_outputs[11768]);
    assign outputs[11824] = ~((layer2_outputs[12265]) ^ (layer2_outputs[2365]));
    assign outputs[11825] = ~((layer2_outputs[5966]) ^ (layer2_outputs[3793]));
    assign outputs[11826] = ~(layer2_outputs[12371]) | (layer2_outputs[11]);
    assign outputs[11827] = ~(layer2_outputs[3994]);
    assign outputs[11828] = layer2_outputs[10307];
    assign outputs[11829] = layer2_outputs[12636];
    assign outputs[11830] = layer2_outputs[6438];
    assign outputs[11831] = ~(layer2_outputs[4943]);
    assign outputs[11832] = layer2_outputs[9917];
    assign outputs[11833] = ~((layer2_outputs[989]) ^ (layer2_outputs[10641]));
    assign outputs[11834] = ~(layer2_outputs[11135]);
    assign outputs[11835] = layer2_outputs[6077];
    assign outputs[11836] = (layer2_outputs[7052]) ^ (layer2_outputs[45]);
    assign outputs[11837] = ~(layer2_outputs[3940]) | (layer2_outputs[3849]);
    assign outputs[11838] = layer2_outputs[621];
    assign outputs[11839] = layer2_outputs[6618];
    assign outputs[11840] = layer2_outputs[11564];
    assign outputs[11841] = ~(layer2_outputs[2086]);
    assign outputs[11842] = layer2_outputs[9173];
    assign outputs[11843] = (layer2_outputs[5104]) & ~(layer2_outputs[2848]);
    assign outputs[11844] = (layer2_outputs[2523]) ^ (layer2_outputs[4938]);
    assign outputs[11845] = (layer2_outputs[8986]) & ~(layer2_outputs[6419]);
    assign outputs[11846] = ~(layer2_outputs[12695]);
    assign outputs[11847] = (layer2_outputs[10535]) & (layer2_outputs[6761]);
    assign outputs[11848] = ~(layer2_outputs[1143]);
    assign outputs[11849] = ~((layer2_outputs[9791]) ^ (layer2_outputs[7391]));
    assign outputs[11850] = layer2_outputs[2690];
    assign outputs[11851] = ~(layer2_outputs[8104]);
    assign outputs[11852] = layer2_outputs[925];
    assign outputs[11853] = (layer2_outputs[6786]) ^ (layer2_outputs[5898]);
    assign outputs[11854] = ~(layer2_outputs[7546]);
    assign outputs[11855] = ~((layer2_outputs[12665]) ^ (layer2_outputs[7250]));
    assign outputs[11856] = (layer2_outputs[3372]) ^ (layer2_outputs[836]);
    assign outputs[11857] = ~((layer2_outputs[1406]) ^ (layer2_outputs[1047]));
    assign outputs[11858] = layer2_outputs[5399];
    assign outputs[11859] = ~(layer2_outputs[5969]);
    assign outputs[11860] = (layer2_outputs[511]) & ~(layer2_outputs[7328]);
    assign outputs[11861] = ~((layer2_outputs[4624]) ^ (layer2_outputs[12286]));
    assign outputs[11862] = ~(layer2_outputs[6123]);
    assign outputs[11863] = layer2_outputs[6563];
    assign outputs[11864] = (layer2_outputs[4841]) & ~(layer2_outputs[2756]);
    assign outputs[11865] = layer2_outputs[6056];
    assign outputs[11866] = layer2_outputs[10461];
    assign outputs[11867] = ~(layer2_outputs[10192]);
    assign outputs[11868] = layer2_outputs[12206];
    assign outputs[11869] = layer2_outputs[4095];
    assign outputs[11870] = layer2_outputs[11887];
    assign outputs[11871] = ~((layer2_outputs[3397]) ^ (layer2_outputs[7056]));
    assign outputs[11872] = (layer2_outputs[8607]) ^ (layer2_outputs[705]);
    assign outputs[11873] = layer2_outputs[7772];
    assign outputs[11874] = layer2_outputs[4117];
    assign outputs[11875] = ~(layer2_outputs[1442]);
    assign outputs[11876] = ~(layer2_outputs[12382]);
    assign outputs[11877] = ~((layer2_outputs[8569]) ^ (layer2_outputs[5367]));
    assign outputs[11878] = layer2_outputs[5453];
    assign outputs[11879] = ~(layer2_outputs[5693]);
    assign outputs[11880] = ~((layer2_outputs[5570]) & (layer2_outputs[4303]));
    assign outputs[11881] = layer2_outputs[1725];
    assign outputs[11882] = (layer2_outputs[11986]) ^ (layer2_outputs[10118]);
    assign outputs[11883] = ~(layer2_outputs[5139]);
    assign outputs[11884] = ~((layer2_outputs[12406]) ^ (layer2_outputs[1190]));
    assign outputs[11885] = (layer2_outputs[9706]) & (layer2_outputs[8984]);
    assign outputs[11886] = ~((layer2_outputs[3991]) ^ (layer2_outputs[3734]));
    assign outputs[11887] = ~(layer2_outputs[12758]);
    assign outputs[11888] = ~(layer2_outputs[4054]);
    assign outputs[11889] = ~(layer2_outputs[6207]);
    assign outputs[11890] = layer2_outputs[10222];
    assign outputs[11891] = ~(layer2_outputs[10300]);
    assign outputs[11892] = (layer2_outputs[7344]) & ~(layer2_outputs[5309]);
    assign outputs[11893] = layer2_outputs[12416];
    assign outputs[11894] = ~((layer2_outputs[1499]) & (layer2_outputs[8042]));
    assign outputs[11895] = ~((layer2_outputs[12524]) ^ (layer2_outputs[8280]));
    assign outputs[11896] = ~(layer2_outputs[9800]);
    assign outputs[11897] = layer2_outputs[6658];
    assign outputs[11898] = ~(layer2_outputs[11180]);
    assign outputs[11899] = (layer2_outputs[11068]) ^ (layer2_outputs[3036]);
    assign outputs[11900] = (layer2_outputs[9649]) & ~(layer2_outputs[7364]);
    assign outputs[11901] = ~(layer2_outputs[8211]);
    assign outputs[11902] = layer2_outputs[4066];
    assign outputs[11903] = layer2_outputs[8926];
    assign outputs[11904] = ~((layer2_outputs[3936]) ^ (layer2_outputs[10392]));
    assign outputs[11905] = (layer2_outputs[10045]) ^ (layer2_outputs[9151]);
    assign outputs[11906] = layer2_outputs[11734];
    assign outputs[11907] = (layer2_outputs[3279]) & (layer2_outputs[3705]);
    assign outputs[11908] = (layer2_outputs[10923]) ^ (layer2_outputs[11363]);
    assign outputs[11909] = ~(layer2_outputs[3182]);
    assign outputs[11910] = layer2_outputs[7035];
    assign outputs[11911] = ~((layer2_outputs[1636]) ^ (layer2_outputs[876]));
    assign outputs[11912] = layer2_outputs[11494];
    assign outputs[11913] = ~(layer2_outputs[3452]);
    assign outputs[11914] = ~(layer2_outputs[8445]);
    assign outputs[11915] = layer2_outputs[7092];
    assign outputs[11916] = layer2_outputs[4714];
    assign outputs[11917] = (layer2_outputs[905]) ^ (layer2_outputs[12793]);
    assign outputs[11918] = ~(layer2_outputs[2022]);
    assign outputs[11919] = (layer2_outputs[5569]) ^ (layer2_outputs[10438]);
    assign outputs[11920] = layer2_outputs[5114];
    assign outputs[11921] = ~((layer2_outputs[9740]) ^ (layer2_outputs[2895]));
    assign outputs[11922] = ~((layer2_outputs[1050]) & (layer2_outputs[7164]));
    assign outputs[11923] = (layer2_outputs[11875]) | (layer2_outputs[8879]);
    assign outputs[11924] = ~(layer2_outputs[7199]);
    assign outputs[11925] = layer2_outputs[6602];
    assign outputs[11926] = (layer2_outputs[2453]) & (layer2_outputs[2750]);
    assign outputs[11927] = layer2_outputs[8946];
    assign outputs[11928] = ~(layer2_outputs[7240]);
    assign outputs[11929] = ~(layer2_outputs[121]);
    assign outputs[11930] = ~((layer2_outputs[273]) | (layer2_outputs[1190]));
    assign outputs[11931] = ~(layer2_outputs[5797]);
    assign outputs[11932] = ~(layer2_outputs[8660]) | (layer2_outputs[8121]);
    assign outputs[11933] = layer2_outputs[7997];
    assign outputs[11934] = ~((layer2_outputs[7802]) | (layer2_outputs[3246]));
    assign outputs[11935] = ~(layer2_outputs[995]);
    assign outputs[11936] = ~((layer2_outputs[4413]) ^ (layer2_outputs[2979]));
    assign outputs[11937] = (layer2_outputs[9030]) & ~(layer2_outputs[1034]);
    assign outputs[11938] = layer2_outputs[4981];
    assign outputs[11939] = ~(layer2_outputs[10336]);
    assign outputs[11940] = layer2_outputs[3137];
    assign outputs[11941] = (layer2_outputs[8954]) & ~(layer2_outputs[1163]);
    assign outputs[11942] = ~(layer2_outputs[3588]);
    assign outputs[11943] = (layer2_outputs[3273]) & ~(layer2_outputs[2516]);
    assign outputs[11944] = ~(layer2_outputs[7379]);
    assign outputs[11945] = layer2_outputs[9135];
    assign outputs[11946] = (layer2_outputs[123]) | (layer2_outputs[9336]);
    assign outputs[11947] = ~((layer2_outputs[9305]) ^ (layer2_outputs[6489]));
    assign outputs[11948] = ~((layer2_outputs[10098]) ^ (layer2_outputs[12031]));
    assign outputs[11949] = ~(layer2_outputs[10090]);
    assign outputs[11950] = ~(layer2_outputs[1410]) | (layer2_outputs[6456]);
    assign outputs[11951] = ~(layer2_outputs[4202]);
    assign outputs[11952] = ~((layer2_outputs[2819]) & (layer2_outputs[10828]));
    assign outputs[11953] = layer2_outputs[6539];
    assign outputs[11954] = (layer2_outputs[10950]) & ~(layer2_outputs[10902]);
    assign outputs[11955] = ~(layer2_outputs[10026]);
    assign outputs[11956] = layer2_outputs[1995];
    assign outputs[11957] = ~(layer2_outputs[624]) | (layer2_outputs[2251]);
    assign outputs[11958] = ~(layer2_outputs[7499]) | (layer2_outputs[2634]);
    assign outputs[11959] = (layer2_outputs[7314]) ^ (layer2_outputs[3934]);
    assign outputs[11960] = (layer2_outputs[4738]) & (layer2_outputs[12267]);
    assign outputs[11961] = layer2_outputs[3570];
    assign outputs[11962] = ~(layer2_outputs[12095]);
    assign outputs[11963] = layer2_outputs[785];
    assign outputs[11964] = layer2_outputs[11541];
    assign outputs[11965] = ~(layer2_outputs[10705]);
    assign outputs[11966] = ~((layer2_outputs[7504]) ^ (layer2_outputs[11614]));
    assign outputs[11967] = ~(layer2_outputs[3414]) | (layer2_outputs[8236]);
    assign outputs[11968] = ~(layer2_outputs[5583]);
    assign outputs[11969] = ~((layer2_outputs[4846]) ^ (layer2_outputs[3818]));
    assign outputs[11970] = (layer2_outputs[5267]) & ~(layer2_outputs[11653]);
    assign outputs[11971] = ~(layer2_outputs[10504]);
    assign outputs[11972] = ~(layer2_outputs[65]);
    assign outputs[11973] = layer2_outputs[12189];
    assign outputs[11974] = ~(layer2_outputs[5493]);
    assign outputs[11975] = ~((layer2_outputs[5834]) | (layer2_outputs[5404]));
    assign outputs[11976] = ~(layer2_outputs[6604]) | (layer2_outputs[11558]);
    assign outputs[11977] = ~((layer2_outputs[7201]) ^ (layer2_outputs[1113]));
    assign outputs[11978] = ~((layer2_outputs[660]) & (layer2_outputs[6198]));
    assign outputs[11979] = ~(layer2_outputs[1996]);
    assign outputs[11980] = (layer2_outputs[11604]) ^ (layer2_outputs[2513]);
    assign outputs[11981] = layer2_outputs[6010];
    assign outputs[11982] = ~(layer2_outputs[7759]) | (layer2_outputs[2769]);
    assign outputs[11983] = layer2_outputs[5448];
    assign outputs[11984] = (layer2_outputs[11048]) & (layer2_outputs[6336]);
    assign outputs[11985] = (layer2_outputs[12]) & ~(layer2_outputs[8458]);
    assign outputs[11986] = layer2_outputs[2189];
    assign outputs[11987] = ~(layer2_outputs[1875]);
    assign outputs[11988] = layer2_outputs[884];
    assign outputs[11989] = ~((layer2_outputs[4226]) | (layer2_outputs[12008]));
    assign outputs[11990] = (layer2_outputs[4562]) | (layer2_outputs[1714]);
    assign outputs[11991] = ~(layer2_outputs[2975]);
    assign outputs[11992] = layer2_outputs[12374];
    assign outputs[11993] = (layer2_outputs[9390]) ^ (layer2_outputs[9856]);
    assign outputs[11994] = ~(layer2_outputs[7008]);
    assign outputs[11995] = (layer2_outputs[11813]) ^ (layer2_outputs[5169]);
    assign outputs[11996] = (layer2_outputs[4242]) ^ (layer2_outputs[5046]);
    assign outputs[11997] = ~(layer2_outputs[5145]);
    assign outputs[11998] = (layer2_outputs[12102]) ^ (layer2_outputs[5687]);
    assign outputs[11999] = ~(layer2_outputs[9839]);
    assign outputs[12000] = ~(layer2_outputs[5656]);
    assign outputs[12001] = (layer2_outputs[1830]) ^ (layer2_outputs[5123]);
    assign outputs[12002] = (layer2_outputs[6960]) ^ (layer2_outputs[6991]);
    assign outputs[12003] = (layer2_outputs[8951]) & (layer2_outputs[659]);
    assign outputs[12004] = (layer2_outputs[3244]) | (layer2_outputs[3577]);
    assign outputs[12005] = layer2_outputs[5756];
    assign outputs[12006] = ~(layer2_outputs[8516]);
    assign outputs[12007] = (layer2_outputs[1075]) | (layer2_outputs[5827]);
    assign outputs[12008] = ~(layer2_outputs[4065]);
    assign outputs[12009] = layer2_outputs[11421];
    assign outputs[12010] = layer2_outputs[10672];
    assign outputs[12011] = layer2_outputs[8493];
    assign outputs[12012] = ~(layer2_outputs[11500]);
    assign outputs[12013] = layer2_outputs[8591];
    assign outputs[12014] = ~(layer2_outputs[1691]);
    assign outputs[12015] = ~((layer2_outputs[6622]) ^ (layer2_outputs[3662]));
    assign outputs[12016] = layer2_outputs[5539];
    assign outputs[12017] = ~(layer2_outputs[11693]);
    assign outputs[12018] = (layer2_outputs[11797]) ^ (layer2_outputs[372]);
    assign outputs[12019] = ~((layer2_outputs[64]) | (layer2_outputs[6657]));
    assign outputs[12020] = ~((layer2_outputs[8494]) ^ (layer2_outputs[9960]));
    assign outputs[12021] = ~(layer2_outputs[6016]);
    assign outputs[12022] = (layer2_outputs[6377]) ^ (layer2_outputs[627]);
    assign outputs[12023] = ~(layer2_outputs[10241]);
    assign outputs[12024] = ~(layer2_outputs[2114]);
    assign outputs[12025] = ~(layer2_outputs[9903]) | (layer2_outputs[4508]);
    assign outputs[12026] = ~(layer2_outputs[4345]);
    assign outputs[12027] = layer2_outputs[12202];
    assign outputs[12028] = ~(layer2_outputs[6712]);
    assign outputs[12029] = ~((layer2_outputs[8133]) | (layer2_outputs[4384]));
    assign outputs[12030] = ~(layer2_outputs[7849]);
    assign outputs[12031] = ~((layer2_outputs[2356]) | (layer2_outputs[12682]));
    assign outputs[12032] = (layer2_outputs[1125]) ^ (layer2_outputs[1618]);
    assign outputs[12033] = ~(layer2_outputs[3907]);
    assign outputs[12034] = (layer2_outputs[3258]) ^ (layer2_outputs[298]);
    assign outputs[12035] = ~(layer2_outputs[4586]);
    assign outputs[12036] = ~(layer2_outputs[940]);
    assign outputs[12037] = layer2_outputs[8426];
    assign outputs[12038] = layer2_outputs[4888];
    assign outputs[12039] = ~((layer2_outputs[7143]) ^ (layer2_outputs[3344]));
    assign outputs[12040] = ~((layer2_outputs[643]) ^ (layer2_outputs[1796]));
    assign outputs[12041] = ~(layer2_outputs[7516]);
    assign outputs[12042] = layer2_outputs[9193];
    assign outputs[12043] = ~((layer2_outputs[5430]) ^ (layer2_outputs[3762]));
    assign outputs[12044] = ~(layer2_outputs[8766]);
    assign outputs[12045] = layer2_outputs[8981];
    assign outputs[12046] = layer2_outputs[878];
    assign outputs[12047] = ~(layer2_outputs[2439]);
    assign outputs[12048] = (layer2_outputs[6949]) ^ (layer2_outputs[5783]);
    assign outputs[12049] = layer2_outputs[2360];
    assign outputs[12050] = ~((layer2_outputs[11138]) & (layer2_outputs[2551]));
    assign outputs[12051] = (layer2_outputs[6270]) & (layer2_outputs[8692]);
    assign outputs[12052] = layer2_outputs[6620];
    assign outputs[12053] = (layer2_outputs[9826]) ^ (layer2_outputs[4019]);
    assign outputs[12054] = ~(layer2_outputs[12302]);
    assign outputs[12055] = ~(layer2_outputs[10297]);
    assign outputs[12056] = layer2_outputs[10347];
    assign outputs[12057] = ~((layer2_outputs[8645]) ^ (layer2_outputs[888]));
    assign outputs[12058] = ~(layer2_outputs[2367]);
    assign outputs[12059] = (layer2_outputs[6337]) ^ (layer2_outputs[8089]);
    assign outputs[12060] = ~(layer2_outputs[3755]);
    assign outputs[12061] = layer2_outputs[6976];
    assign outputs[12062] = ~((layer2_outputs[7850]) & (layer2_outputs[2165]));
    assign outputs[12063] = layer2_outputs[1312];
    assign outputs[12064] = (layer2_outputs[2801]) | (layer2_outputs[3361]);
    assign outputs[12065] = layer2_outputs[2422];
    assign outputs[12066] = layer2_outputs[12773];
    assign outputs[12067] = (layer2_outputs[1940]) ^ (layer2_outputs[9607]);
    assign outputs[12068] = layer2_outputs[5261];
    assign outputs[12069] = layer2_outputs[8527];
    assign outputs[12070] = (layer2_outputs[12244]) ^ (layer2_outputs[4259]);
    assign outputs[12071] = ~((layer2_outputs[736]) | (layer2_outputs[11087]));
    assign outputs[12072] = ~(layer2_outputs[11648]);
    assign outputs[12073] = ~(layer2_outputs[7644]);
    assign outputs[12074] = layer2_outputs[452];
    assign outputs[12075] = ~(layer2_outputs[5272]);
    assign outputs[12076] = ~((layer2_outputs[3513]) ^ (layer2_outputs[3581]));
    assign outputs[12077] = (layer2_outputs[1156]) & (layer2_outputs[2968]);
    assign outputs[12078] = layer2_outputs[9107];
    assign outputs[12079] = (layer2_outputs[2997]) & (layer2_outputs[8462]);
    assign outputs[12080] = ~(layer2_outputs[12025]);
    assign outputs[12081] = ~(layer2_outputs[6820]);
    assign outputs[12082] = (layer2_outputs[4097]) ^ (layer2_outputs[11818]);
    assign outputs[12083] = (layer2_outputs[9731]) & (layer2_outputs[4916]);
    assign outputs[12084] = ~((layer2_outputs[12777]) ^ (layer2_outputs[5292]));
    assign outputs[12085] = ~(layer2_outputs[11185]);
    assign outputs[12086] = (layer2_outputs[8121]) & ~(layer2_outputs[6118]);
    assign outputs[12087] = ~(layer2_outputs[5530]);
    assign outputs[12088] = layer2_outputs[936];
    assign outputs[12089] = ~(layer2_outputs[638]) | (layer2_outputs[1437]);
    assign outputs[12090] = ~((layer2_outputs[2262]) & (layer2_outputs[8281]));
    assign outputs[12091] = (layer2_outputs[5320]) ^ (layer2_outputs[9526]);
    assign outputs[12092] = ~(layer2_outputs[6743]) | (layer2_outputs[2461]);
    assign outputs[12093] = layer2_outputs[7318];
    assign outputs[12094] = (layer2_outputs[2540]) & ~(layer2_outputs[7483]);
    assign outputs[12095] = (layer2_outputs[5344]) ^ (layer2_outputs[2743]);
    assign outputs[12096] = (layer2_outputs[8496]) ^ (layer2_outputs[12546]);
    assign outputs[12097] = ~(layer2_outputs[7216]);
    assign outputs[12098] = ~((layer2_outputs[10055]) ^ (layer2_outputs[8241]));
    assign outputs[12099] = ~((layer2_outputs[9014]) ^ (layer2_outputs[755]));
    assign outputs[12100] = ~((layer2_outputs[10240]) ^ (layer2_outputs[4675]));
    assign outputs[12101] = ~(layer2_outputs[1824]);
    assign outputs[12102] = (layer2_outputs[728]) & ~(layer2_outputs[247]);
    assign outputs[12103] = ~(layer2_outputs[3614]);
    assign outputs[12104] = layer2_outputs[8260];
    assign outputs[12105] = layer2_outputs[5434];
    assign outputs[12106] = layer2_outputs[9069];
    assign outputs[12107] = layer2_outputs[4371];
    assign outputs[12108] = (layer2_outputs[9425]) ^ (layer2_outputs[8492]);
    assign outputs[12109] = ~((layer2_outputs[6546]) ^ (layer2_outputs[5934]));
    assign outputs[12110] = layer2_outputs[12565];
    assign outputs[12111] = ~(layer2_outputs[5182]) | (layer2_outputs[2662]);
    assign outputs[12112] = layer2_outputs[5444];
    assign outputs[12113] = ~(layer2_outputs[6098]);
    assign outputs[12114] = (layer2_outputs[8834]) & ~(layer2_outputs[11985]);
    assign outputs[12115] = (layer2_outputs[15]) ^ (layer2_outputs[7396]);
    assign outputs[12116] = layer2_outputs[1177];
    assign outputs[12117] = layer2_outputs[8343];
    assign outputs[12118] = ~(layer2_outputs[11095]) | (layer2_outputs[455]);
    assign outputs[12119] = layer2_outputs[8483];
    assign outputs[12120] = ~(layer2_outputs[12484]);
    assign outputs[12121] = layer2_outputs[2963];
    assign outputs[12122] = (layer2_outputs[2009]) & (layer2_outputs[12186]);
    assign outputs[12123] = (layer2_outputs[4173]) ^ (layer2_outputs[10285]);
    assign outputs[12124] = layer2_outputs[7351];
    assign outputs[12125] = ~(layer2_outputs[5046]) | (layer2_outputs[11015]);
    assign outputs[12126] = ~(layer2_outputs[9548]);
    assign outputs[12127] = ~((layer2_outputs[7220]) ^ (layer2_outputs[3922]));
    assign outputs[12128] = ~((layer2_outputs[2734]) & (layer2_outputs[12356]));
    assign outputs[12129] = (layer2_outputs[10764]) & (layer2_outputs[9013]);
    assign outputs[12130] = ~(layer2_outputs[1308]);
    assign outputs[12131] = (layer2_outputs[12412]) ^ (layer2_outputs[4786]);
    assign outputs[12132] = (layer2_outputs[2108]) ^ (layer2_outputs[928]);
    assign outputs[12133] = layer2_outputs[6804];
    assign outputs[12134] = ~((layer2_outputs[7679]) & (layer2_outputs[6988]));
    assign outputs[12135] = (layer2_outputs[82]) ^ (layer2_outputs[7891]);
    assign outputs[12136] = ~((layer2_outputs[5501]) | (layer2_outputs[6582]));
    assign outputs[12137] = layer2_outputs[8735];
    assign outputs[12138] = layer2_outputs[4602];
    assign outputs[12139] = ~(layer2_outputs[9571]);
    assign outputs[12140] = ~(layer2_outputs[10974]);
    assign outputs[12141] = ~(layer2_outputs[976]);
    assign outputs[12142] = (layer2_outputs[10078]) ^ (layer2_outputs[7988]);
    assign outputs[12143] = layer2_outputs[11837];
    assign outputs[12144] = (layer2_outputs[11210]) & ~(layer2_outputs[12182]);
    assign outputs[12145] = (layer2_outputs[9660]) ^ (layer2_outputs[8896]);
    assign outputs[12146] = layer2_outputs[680];
    assign outputs[12147] = layer2_outputs[6751];
    assign outputs[12148] = ~(layer2_outputs[1145]);
    assign outputs[12149] = ~((layer2_outputs[7939]) ^ (layer2_outputs[4511]));
    assign outputs[12150] = ~((layer2_outputs[9052]) ^ (layer2_outputs[11717]));
    assign outputs[12151] = layer2_outputs[3153];
    assign outputs[12152] = ~(layer2_outputs[7942]);
    assign outputs[12153] = ~(layer2_outputs[11500]);
    assign outputs[12154] = layer2_outputs[7502];
    assign outputs[12155] = ~(layer2_outputs[4115]);
    assign outputs[12156] = ~(layer2_outputs[8233]);
    assign outputs[12157] = ~(layer2_outputs[5084]);
    assign outputs[12158] = ~(layer2_outputs[9356]);
    assign outputs[12159] = layer2_outputs[3277];
    assign outputs[12160] = ~((layer2_outputs[8832]) ^ (layer2_outputs[10432]));
    assign outputs[12161] = (layer2_outputs[3543]) ^ (layer2_outputs[8366]);
    assign outputs[12162] = layer2_outputs[7230];
    assign outputs[12163] = ~(layer2_outputs[9584]);
    assign outputs[12164] = (layer2_outputs[11760]) & (layer2_outputs[3239]);
    assign outputs[12165] = ~(layer2_outputs[2073]);
    assign outputs[12166] = ~(layer2_outputs[6516]);
    assign outputs[12167] = (layer2_outputs[6399]) ^ (layer2_outputs[123]);
    assign outputs[12168] = (layer2_outputs[5171]) ^ (layer2_outputs[12115]);
    assign outputs[12169] = ~(layer2_outputs[5801]);
    assign outputs[12170] = ~((layer2_outputs[6402]) ^ (layer2_outputs[475]));
    assign outputs[12171] = (layer2_outputs[1092]) ^ (layer2_outputs[7801]);
    assign outputs[12172] = layer2_outputs[10801];
    assign outputs[12173] = ~(layer2_outputs[4386]);
    assign outputs[12174] = layer2_outputs[2609];
    assign outputs[12175] = (layer2_outputs[880]) & ~(layer2_outputs[10510]);
    assign outputs[12176] = layer2_outputs[3059];
    assign outputs[12177] = ~((layer2_outputs[5829]) ^ (layer2_outputs[5342]));
    assign outputs[12178] = layer2_outputs[5959];
    assign outputs[12179] = ~(layer2_outputs[6541]);
    assign outputs[12180] = ~(layer2_outputs[3529]);
    assign outputs[12181] = layer2_outputs[1073];
    assign outputs[12182] = (layer2_outputs[6993]) & ~(layer2_outputs[6799]);
    assign outputs[12183] = ~(layer2_outputs[4660]);
    assign outputs[12184] = 1'b1;
    assign outputs[12185] = layer2_outputs[4775];
    assign outputs[12186] = (layer2_outputs[11494]) & (layer2_outputs[3923]);
    assign outputs[12187] = layer2_outputs[1874];
    assign outputs[12188] = layer2_outputs[5597];
    assign outputs[12189] = ~(layer2_outputs[294]);
    assign outputs[12190] = ~((layer2_outputs[3952]) | (layer2_outputs[3219]));
    assign outputs[12191] = layer2_outputs[3287];
    assign outputs[12192] = ~(layer2_outputs[9644]);
    assign outputs[12193] = ~(layer2_outputs[4637]);
    assign outputs[12194] = (layer2_outputs[3972]) | (layer2_outputs[10099]);
    assign outputs[12195] = ~((layer2_outputs[10895]) | (layer2_outputs[1130]));
    assign outputs[12196] = ~((layer2_outputs[1203]) ^ (layer2_outputs[218]));
    assign outputs[12197] = ~((layer2_outputs[5347]) ^ (layer2_outputs[10055]));
    assign outputs[12198] = ~((layer2_outputs[6856]) ^ (layer2_outputs[5376]));
    assign outputs[12199] = ~((layer2_outputs[5009]) ^ (layer2_outputs[8543]));
    assign outputs[12200] = (layer2_outputs[7705]) ^ (layer2_outputs[7572]);
    assign outputs[12201] = ~((layer2_outputs[11846]) | (layer2_outputs[10615]));
    assign outputs[12202] = ~((layer2_outputs[7980]) & (layer2_outputs[11925]));
    assign outputs[12203] = ~(layer2_outputs[6817]);
    assign outputs[12204] = ~(layer2_outputs[10711]);
    assign outputs[12205] = layer2_outputs[10371];
    assign outputs[12206] = ~((layer2_outputs[10268]) ^ (layer2_outputs[6561]));
    assign outputs[12207] = layer2_outputs[2270];
    assign outputs[12208] = (layer2_outputs[7960]) & ~(layer2_outputs[4499]);
    assign outputs[12209] = (layer2_outputs[1812]) ^ (layer2_outputs[144]);
    assign outputs[12210] = ~(layer2_outputs[10388]);
    assign outputs[12211] = ~(layer2_outputs[9095]);
    assign outputs[12212] = (layer2_outputs[9568]) ^ (layer2_outputs[12274]);
    assign outputs[12213] = layer2_outputs[7605];
    assign outputs[12214] = ~(layer2_outputs[12180]);
    assign outputs[12215] = ~(layer2_outputs[5003]) | (layer2_outputs[535]);
    assign outputs[12216] = layer2_outputs[3919];
    assign outputs[12217] = ~(layer2_outputs[5451]) | (layer2_outputs[4101]);
    assign outputs[12218] = ~((layer2_outputs[1683]) ^ (layer2_outputs[7669]));
    assign outputs[12219] = ~((layer2_outputs[8803]) ^ (layer2_outputs[10799]));
    assign outputs[12220] = ~(layer2_outputs[6420]) | (layer2_outputs[10285]);
    assign outputs[12221] = layer2_outputs[6312];
    assign outputs[12222] = (layer2_outputs[3130]) & ~(layer2_outputs[9110]);
    assign outputs[12223] = ~(layer2_outputs[6896]);
    assign outputs[12224] = ~(layer2_outputs[1463]);
    assign outputs[12225] = (layer2_outputs[8242]) & ~(layer2_outputs[7099]);
    assign outputs[12226] = layer2_outputs[1289];
    assign outputs[12227] = layer2_outputs[10264];
    assign outputs[12228] = (layer2_outputs[4954]) & ~(layer2_outputs[860]);
    assign outputs[12229] = ~(layer2_outputs[2020]);
    assign outputs[12230] = layer2_outputs[12414];
    assign outputs[12231] = (layer2_outputs[9431]) & (layer2_outputs[7814]);
    assign outputs[12232] = ~(layer2_outputs[6604]) | (layer2_outputs[8096]);
    assign outputs[12233] = (layer2_outputs[3826]) & ~(layer2_outputs[1196]);
    assign outputs[12234] = ~(layer2_outputs[6667]);
    assign outputs[12235] = ~(layer2_outputs[6351]);
    assign outputs[12236] = ~((layer2_outputs[7023]) | (layer2_outputs[10173]));
    assign outputs[12237] = (layer2_outputs[11567]) ^ (layer2_outputs[2075]);
    assign outputs[12238] = ~((layer2_outputs[6855]) ^ (layer2_outputs[4476]));
    assign outputs[12239] = ~((layer2_outputs[9980]) & (layer2_outputs[3635]));
    assign outputs[12240] = ~(layer2_outputs[5573]);
    assign outputs[12241] = ~(layer2_outputs[11583]);
    assign outputs[12242] = ~(layer2_outputs[10935]);
    assign outputs[12243] = ~(layer2_outputs[10168]);
    assign outputs[12244] = (layer2_outputs[11535]) ^ (layer2_outputs[1226]);
    assign outputs[12245] = (layer2_outputs[10279]) & ~(layer2_outputs[2146]);
    assign outputs[12246] = layer2_outputs[9645];
    assign outputs[12247] = (layer2_outputs[9205]) & ~(layer2_outputs[1162]);
    assign outputs[12248] = ~(layer2_outputs[2913]);
    assign outputs[12249] = layer2_outputs[9717];
    assign outputs[12250] = ~(layer2_outputs[7914]);
    assign outputs[12251] = ~(layer2_outputs[11307]);
    assign outputs[12252] = layer2_outputs[4773];
    assign outputs[12253] = ~(layer2_outputs[9862]);
    assign outputs[12254] = layer2_outputs[7029];
    assign outputs[12255] = layer2_outputs[4265];
    assign outputs[12256] = (layer2_outputs[975]) ^ (layer2_outputs[5670]);
    assign outputs[12257] = (layer2_outputs[5335]) ^ (layer2_outputs[4280]);
    assign outputs[12258] = layer2_outputs[4];
    assign outputs[12259] = layer2_outputs[4587];
    assign outputs[12260] = layer2_outputs[5614];
    assign outputs[12261] = ~(layer2_outputs[1038]);
    assign outputs[12262] = ~(layer2_outputs[10913]);
    assign outputs[12263] = ~(layer2_outputs[2401]);
    assign outputs[12264] = ~(layer2_outputs[2960]);
    assign outputs[12265] = (layer2_outputs[4361]) ^ (layer2_outputs[6713]);
    assign outputs[12266] = ~(layer2_outputs[10967]);
    assign outputs[12267] = ~(layer2_outputs[5285]);
    assign outputs[12268] = (layer2_outputs[12413]) & ~(layer2_outputs[12419]);
    assign outputs[12269] = ~(layer2_outputs[5762]);
    assign outputs[12270] = layer2_outputs[4790];
    assign outputs[12271] = layer2_outputs[4923];
    assign outputs[12272] = (layer2_outputs[9662]) ^ (layer2_outputs[3123]);
    assign outputs[12273] = layer2_outputs[10137];
    assign outputs[12274] = layer2_outputs[386];
    assign outputs[12275] = layer2_outputs[979];
    assign outputs[12276] = layer2_outputs[8476];
    assign outputs[12277] = (layer2_outputs[4827]) ^ (layer2_outputs[1728]);
    assign outputs[12278] = ~(layer2_outputs[3502]);
    assign outputs[12279] = layer2_outputs[3408];
    assign outputs[12280] = ~(layer2_outputs[2250]);
    assign outputs[12281] = ~((layer2_outputs[11332]) ^ (layer2_outputs[11708]));
    assign outputs[12282] = layer2_outputs[4799];
    assign outputs[12283] = ~(layer2_outputs[1890]);
    assign outputs[12284] = ~((layer2_outputs[3330]) | (layer2_outputs[6869]));
    assign outputs[12285] = (layer2_outputs[3013]) ^ (layer2_outputs[11617]);
    assign outputs[12286] = ~(layer2_outputs[10192]);
    assign outputs[12287] = layer2_outputs[3509];
    assign outputs[12288] = ~(layer2_outputs[9191]);
    assign outputs[12289] = (layer2_outputs[956]) ^ (layer2_outputs[10551]);
    assign outputs[12290] = ~((layer2_outputs[8651]) ^ (layer2_outputs[1434]));
    assign outputs[12291] = layer2_outputs[8243];
    assign outputs[12292] = (layer2_outputs[5643]) ^ (layer2_outputs[7698]);
    assign outputs[12293] = ~((layer2_outputs[10197]) ^ (layer2_outputs[7844]));
    assign outputs[12294] = layer2_outputs[11415];
    assign outputs[12295] = ~(layer2_outputs[11017]);
    assign outputs[12296] = layer2_outputs[4141];
    assign outputs[12297] = ~(layer2_outputs[10468]);
    assign outputs[12298] = ~(layer2_outputs[5743]);
    assign outputs[12299] = layer2_outputs[9289];
    assign outputs[12300] = ~((layer2_outputs[2079]) | (layer2_outputs[10141]));
    assign outputs[12301] = layer2_outputs[403];
    assign outputs[12302] = ~(layer2_outputs[10864]);
    assign outputs[12303] = (layer2_outputs[7120]) ^ (layer2_outputs[3004]);
    assign outputs[12304] = layer2_outputs[10186];
    assign outputs[12305] = ~(layer2_outputs[917]);
    assign outputs[12306] = (layer2_outputs[11265]) ^ (layer2_outputs[7866]);
    assign outputs[12307] = (layer2_outputs[3920]) ^ (layer2_outputs[11460]);
    assign outputs[12308] = (layer2_outputs[8223]) & ~(layer2_outputs[9171]);
    assign outputs[12309] = ~(layer2_outputs[3985]);
    assign outputs[12310] = (layer2_outputs[2766]) ^ (layer2_outputs[9072]);
    assign outputs[12311] = layer2_outputs[5304];
    assign outputs[12312] = (layer2_outputs[11791]) ^ (layer2_outputs[12177]);
    assign outputs[12313] = ~((layer2_outputs[1110]) ^ (layer2_outputs[2977]));
    assign outputs[12314] = ~((layer2_outputs[2895]) ^ (layer2_outputs[1453]));
    assign outputs[12315] = (layer2_outputs[9604]) & ~(layer2_outputs[6973]);
    assign outputs[12316] = ~((layer2_outputs[3659]) ^ (layer2_outputs[1084]));
    assign outputs[12317] = (layer2_outputs[5593]) ^ (layer2_outputs[3708]);
    assign outputs[12318] = layer2_outputs[7457];
    assign outputs[12319] = ~((layer2_outputs[8756]) | (layer2_outputs[10401]));
    assign outputs[12320] = ~((layer2_outputs[9804]) ^ (layer2_outputs[1990]));
    assign outputs[12321] = layer2_outputs[7959];
    assign outputs[12322] = layer2_outputs[12519];
    assign outputs[12323] = (layer2_outputs[8839]) ^ (layer2_outputs[1063]);
    assign outputs[12324] = ~(layer2_outputs[71]);
    assign outputs[12325] = ~(layer2_outputs[6750]);
    assign outputs[12326] = ~(layer2_outputs[12728]) | (layer2_outputs[7737]);
    assign outputs[12327] = ~((layer2_outputs[2283]) ^ (layer2_outputs[154]));
    assign outputs[12328] = ~(layer2_outputs[1755]);
    assign outputs[12329] = layer2_outputs[2655];
    assign outputs[12330] = ~(layer2_outputs[11193]);
    assign outputs[12331] = layer2_outputs[12788];
    assign outputs[12332] = ~((layer2_outputs[6578]) | (layer2_outputs[4741]));
    assign outputs[12333] = ~((layer2_outputs[5071]) ^ (layer2_outputs[9343]));
    assign outputs[12334] = ~(layer2_outputs[8026]);
    assign outputs[12335] = ~(layer2_outputs[3336]) | (layer2_outputs[6395]);
    assign outputs[12336] = (layer2_outputs[4320]) & (layer2_outputs[6377]);
    assign outputs[12337] = ~(layer2_outputs[11143]) | (layer2_outputs[12479]);
    assign outputs[12338] = layer2_outputs[12756];
    assign outputs[12339] = ~((layer2_outputs[7573]) | (layer2_outputs[6151]));
    assign outputs[12340] = layer2_outputs[6393];
    assign outputs[12341] = (layer2_outputs[11245]) | (layer2_outputs[1261]);
    assign outputs[12342] = layer2_outputs[7664];
    assign outputs[12343] = layer2_outputs[1144];
    assign outputs[12344] = ~(layer2_outputs[6036]);
    assign outputs[12345] = layer2_outputs[2856];
    assign outputs[12346] = layer2_outputs[11424];
    assign outputs[12347] = ~(layer2_outputs[7375]);
    assign outputs[12348] = ~((layer2_outputs[3183]) & (layer2_outputs[882]));
    assign outputs[12349] = (layer2_outputs[8053]) & (layer2_outputs[2109]);
    assign outputs[12350] = (layer2_outputs[9316]) ^ (layer2_outputs[2462]);
    assign outputs[12351] = (layer2_outputs[58]) ^ (layer2_outputs[6158]);
    assign outputs[12352] = layer2_outputs[3127];
    assign outputs[12353] = layer2_outputs[3480];
    assign outputs[12354] = ~(layer2_outputs[7715]);
    assign outputs[12355] = ~((layer2_outputs[10252]) ^ (layer2_outputs[6457]));
    assign outputs[12356] = ~((layer2_outputs[9596]) ^ (layer2_outputs[9304]));
    assign outputs[12357] = layer2_outputs[11780];
    assign outputs[12358] = layer2_outputs[10921];
    assign outputs[12359] = ~(layer2_outputs[482]);
    assign outputs[12360] = ~(layer2_outputs[12611]);
    assign outputs[12361] = layer2_outputs[4070];
    assign outputs[12362] = layer2_outputs[3093];
    assign outputs[12363] = ~(layer2_outputs[1738]);
    assign outputs[12364] = ~(layer2_outputs[10931]);
    assign outputs[12365] = layer2_outputs[139];
    assign outputs[12366] = (layer2_outputs[11053]) ^ (layer2_outputs[3115]);
    assign outputs[12367] = layer2_outputs[6628];
    assign outputs[12368] = ~(layer2_outputs[12158]) | (layer2_outputs[951]);
    assign outputs[12369] = layer2_outputs[4407];
    assign outputs[12370] = ~(layer2_outputs[262]) | (layer2_outputs[5300]);
    assign outputs[12371] = ~((layer2_outputs[4702]) & (layer2_outputs[8538]));
    assign outputs[12372] = layer2_outputs[5942];
    assign outputs[12373] = layer2_outputs[10555];
    assign outputs[12374] = (layer2_outputs[2781]) ^ (layer2_outputs[56]);
    assign outputs[12375] = ~((layer2_outputs[9417]) ^ (layer2_outputs[6917]));
    assign outputs[12376] = (layer2_outputs[5479]) ^ (layer2_outputs[4229]);
    assign outputs[12377] = layer2_outputs[11814];
    assign outputs[12378] = (layer2_outputs[9070]) ^ (layer2_outputs[6268]);
    assign outputs[12379] = layer2_outputs[5100];
    assign outputs[12380] = ~((layer2_outputs[3410]) ^ (layer2_outputs[12187]));
    assign outputs[12381] = ~((layer2_outputs[5318]) & (layer2_outputs[4314]));
    assign outputs[12382] = (layer2_outputs[7472]) & ~(layer2_outputs[10036]);
    assign outputs[12383] = layer2_outputs[4948];
    assign outputs[12384] = ~(layer2_outputs[9601]);
    assign outputs[12385] = ~(layer2_outputs[6464]);
    assign outputs[12386] = layer2_outputs[7108];
    assign outputs[12387] = (layer2_outputs[1239]) ^ (layer2_outputs[1458]);
    assign outputs[12388] = ~(layer2_outputs[328]);
    assign outputs[12389] = layer2_outputs[7725];
    assign outputs[12390] = ~((layer2_outputs[12344]) ^ (layer2_outputs[4669]));
    assign outputs[12391] = (layer2_outputs[11461]) | (layer2_outputs[1035]);
    assign outputs[12392] = ~(layer2_outputs[7406]);
    assign outputs[12393] = ~(layer2_outputs[7203]) | (layer2_outputs[5385]);
    assign outputs[12394] = (layer2_outputs[3039]) ^ (layer2_outputs[12531]);
    assign outputs[12395] = layer2_outputs[12111];
    assign outputs[12396] = ~((layer2_outputs[8932]) ^ (layer2_outputs[2797]));
    assign outputs[12397] = ~(layer2_outputs[7047]);
    assign outputs[12398] = layer2_outputs[7523];
    assign outputs[12399] = ~((layer2_outputs[12209]) ^ (layer2_outputs[11304]));
    assign outputs[12400] = ~(layer2_outputs[1967]);
    assign outputs[12401] = ~((layer2_outputs[1355]) ^ (layer2_outputs[482]));
    assign outputs[12402] = ~(layer2_outputs[7357]);
    assign outputs[12403] = ~((layer2_outputs[12782]) | (layer2_outputs[4115]));
    assign outputs[12404] = ~(layer2_outputs[10410]);
    assign outputs[12405] = ~(layer2_outputs[6069]);
    assign outputs[12406] = layer2_outputs[9054];
    assign outputs[12407] = ~(layer2_outputs[3957]);
    assign outputs[12408] = ~((layer2_outputs[1036]) ^ (layer2_outputs[6184]));
    assign outputs[12409] = (layer2_outputs[4277]) | (layer2_outputs[142]);
    assign outputs[12410] = ~((layer2_outputs[11216]) ^ (layer2_outputs[11616]));
    assign outputs[12411] = ~((layer2_outputs[11504]) ^ (layer2_outputs[10558]));
    assign outputs[12412] = layer2_outputs[6880];
    assign outputs[12413] = ~(layer2_outputs[27]) | (layer2_outputs[11699]);
    assign outputs[12414] = ~((layer2_outputs[6226]) | (layer2_outputs[10538]));
    assign outputs[12415] = ~((layer2_outputs[6974]) ^ (layer2_outputs[5581]));
    assign outputs[12416] = ~((layer2_outputs[6943]) ^ (layer2_outputs[9360]));
    assign outputs[12417] = layer2_outputs[9994];
    assign outputs[12418] = ~(layer2_outputs[6153]);
    assign outputs[12419] = ~(layer2_outputs[9329]);
    assign outputs[12420] = (layer2_outputs[9565]) ^ (layer2_outputs[563]);
    assign outputs[12421] = layer2_outputs[12373];
    assign outputs[12422] = ~(layer2_outputs[513]);
    assign outputs[12423] = layer2_outputs[5315];
    assign outputs[12424] = ~(layer2_outputs[8132]);
    assign outputs[12425] = ~(layer2_outputs[4544]);
    assign outputs[12426] = ~(layer2_outputs[8075]);
    assign outputs[12427] = ~((layer2_outputs[514]) ^ (layer2_outputs[5849]));
    assign outputs[12428] = ~(layer2_outputs[1977]);
    assign outputs[12429] = ~(layer2_outputs[4304]);
    assign outputs[12430] = ~(layer2_outputs[1067]);
    assign outputs[12431] = ~(layer2_outputs[180]) | (layer2_outputs[4735]);
    assign outputs[12432] = (layer2_outputs[10685]) & (layer2_outputs[9949]);
    assign outputs[12433] = (layer2_outputs[7308]) & (layer2_outputs[7317]);
    assign outputs[12434] = ~((layer2_outputs[3177]) | (layer2_outputs[10710]));
    assign outputs[12435] = ~((layer2_outputs[9247]) ^ (layer2_outputs[255]));
    assign outputs[12436] = ~((layer2_outputs[3563]) & (layer2_outputs[2094]));
    assign outputs[12437] = layer2_outputs[3326];
    assign outputs[12438] = layer2_outputs[11875];
    assign outputs[12439] = ~(layer2_outputs[5549]) | (layer2_outputs[11058]);
    assign outputs[12440] = ~(layer2_outputs[2059]);
    assign outputs[12441] = ~(layer2_outputs[12509]);
    assign outputs[12442] = ~(layer2_outputs[10096]) | (layer2_outputs[973]);
    assign outputs[12443] = (layer2_outputs[5439]) ^ (layer2_outputs[8682]);
    assign outputs[12444] = ~(layer2_outputs[4962]);
    assign outputs[12445] = ~((layer2_outputs[10844]) ^ (layer2_outputs[5591]));
    assign outputs[12446] = layer2_outputs[7873];
    assign outputs[12447] = layer2_outputs[7605];
    assign outputs[12448] = ~(layer2_outputs[9299]);
    assign outputs[12449] = ~(layer2_outputs[2573]);
    assign outputs[12450] = layer2_outputs[1764];
    assign outputs[12451] = (layer2_outputs[5962]) & ~(layer2_outputs[2029]);
    assign outputs[12452] = layer2_outputs[7554];
    assign outputs[12453] = ~(layer2_outputs[11329]);
    assign outputs[12454] = layer2_outputs[2241];
    assign outputs[12455] = layer2_outputs[5804];
    assign outputs[12456] = layer2_outputs[12088];
    assign outputs[12457] = layer2_outputs[1520];
    assign outputs[12458] = ~(layer2_outputs[5977]);
    assign outputs[12459] = (layer2_outputs[6347]) | (layer2_outputs[8196]);
    assign outputs[12460] = ~((layer2_outputs[9075]) ^ (layer2_outputs[7888]));
    assign outputs[12461] = ~(layer2_outputs[4724]);
    assign outputs[12462] = ~(layer2_outputs[5049]);
    assign outputs[12463] = (layer2_outputs[8815]) & ~(layer2_outputs[4715]);
    assign outputs[12464] = layer2_outputs[6627];
    assign outputs[12465] = (layer2_outputs[6214]) & ~(layer2_outputs[8883]);
    assign outputs[12466] = (layer2_outputs[3484]) ^ (layer2_outputs[6196]);
    assign outputs[12467] = (layer2_outputs[10908]) ^ (layer2_outputs[6684]);
    assign outputs[12468] = ~(layer2_outputs[5625]);
    assign outputs[12469] = ~(layer2_outputs[10933]);
    assign outputs[12470] = ~(layer2_outputs[8676]);
    assign outputs[12471] = (layer2_outputs[5865]) | (layer2_outputs[1211]);
    assign outputs[12472] = ~(layer2_outputs[3312]);
    assign outputs[12473] = layer2_outputs[3239];
    assign outputs[12474] = ~(layer2_outputs[6465]);
    assign outputs[12475] = ~(layer2_outputs[12169]);
    assign outputs[12476] = ~((layer2_outputs[525]) | (layer2_outputs[12524]));
    assign outputs[12477] = ~(layer2_outputs[9779]);
    assign outputs[12478] = (layer2_outputs[70]) ^ (layer2_outputs[4179]);
    assign outputs[12479] = layer2_outputs[7374];
    assign outputs[12480] = ~((layer2_outputs[8669]) ^ (layer2_outputs[2729]));
    assign outputs[12481] = layer2_outputs[8723];
    assign outputs[12482] = ~(layer2_outputs[601]) | (layer2_outputs[11120]);
    assign outputs[12483] = layer2_outputs[6335];
    assign outputs[12484] = (layer2_outputs[9388]) ^ (layer2_outputs[2152]);
    assign outputs[12485] = (layer2_outputs[8113]) ^ (layer2_outputs[12028]);
    assign outputs[12486] = layer2_outputs[538];
    assign outputs[12487] = ~(layer2_outputs[3479]) | (layer2_outputs[12392]);
    assign outputs[12488] = (layer2_outputs[8175]) ^ (layer2_outputs[423]);
    assign outputs[12489] = ~(layer2_outputs[12096]) | (layer2_outputs[7868]);
    assign outputs[12490] = ~(layer2_outputs[1630]);
    assign outputs[12491] = layer2_outputs[3276];
    assign outputs[12492] = layer2_outputs[10531];
    assign outputs[12493] = ~(layer2_outputs[4724]) | (layer2_outputs[11072]);
    assign outputs[12494] = ~(layer2_outputs[3286]);
    assign outputs[12495] = (layer2_outputs[3551]) & ~(layer2_outputs[10060]);
    assign outputs[12496] = layer2_outputs[4709];
    assign outputs[12497] = (layer2_outputs[2340]) ^ (layer2_outputs[5633]);
    assign outputs[12498] = (layer2_outputs[4640]) ^ (layer2_outputs[7652]);
    assign outputs[12499] = (layer2_outputs[6962]) & ~(layer2_outputs[3934]);
    assign outputs[12500] = ~(layer2_outputs[2282]);
    assign outputs[12501] = ~(layer2_outputs[3049]);
    assign outputs[12502] = layer2_outputs[3509];
    assign outputs[12503] = (layer2_outputs[10893]) & ~(layer2_outputs[4983]);
    assign outputs[12504] = ~(layer2_outputs[7361]);
    assign outputs[12505] = ~(layer2_outputs[11082]);
    assign outputs[12506] = (layer2_outputs[10787]) & (layer2_outputs[12016]);
    assign outputs[12507] = layer2_outputs[9938];
    assign outputs[12508] = ~(layer2_outputs[9987]);
    assign outputs[12509] = (layer2_outputs[8716]) & ~(layer2_outputs[332]);
    assign outputs[12510] = ~(layer2_outputs[1062]);
    assign outputs[12511] = layer2_outputs[4432];
    assign outputs[12512] = ~(layer2_outputs[2552]);
    assign outputs[12513] = layer2_outputs[9064];
    assign outputs[12514] = ~(layer2_outputs[9969]);
    assign outputs[12515] = (layer2_outputs[9831]) ^ (layer2_outputs[2629]);
    assign outputs[12516] = layer2_outputs[10164];
    assign outputs[12517] = ~((layer2_outputs[1091]) ^ (layer2_outputs[5642]));
    assign outputs[12518] = ~(layer2_outputs[7926]) | (layer2_outputs[9625]);
    assign outputs[12519] = ~((layer2_outputs[12063]) & (layer2_outputs[3770]));
    assign outputs[12520] = ~(layer2_outputs[3699]);
    assign outputs[12521] = (layer2_outputs[6369]) & ~(layer2_outputs[9752]);
    assign outputs[12522] = ~(layer2_outputs[1992]) | (layer2_outputs[462]);
    assign outputs[12523] = ~((layer2_outputs[6884]) ^ (layer2_outputs[6724]));
    assign outputs[12524] = (layer2_outputs[4516]) & (layer2_outputs[10210]);
    assign outputs[12525] = ~((layer2_outputs[12328]) | (layer2_outputs[10001]));
    assign outputs[12526] = (layer2_outputs[2845]) ^ (layer2_outputs[6635]);
    assign outputs[12527] = ~(layer2_outputs[1260]);
    assign outputs[12528] = layer2_outputs[1500];
    assign outputs[12529] = ~((layer2_outputs[11385]) ^ (layer2_outputs[11406]));
    assign outputs[12530] = (layer2_outputs[10615]) ^ (layer2_outputs[4365]);
    assign outputs[12531] = layer2_outputs[6300];
    assign outputs[12532] = layer2_outputs[1501];
    assign outputs[12533] = (layer2_outputs[3144]) | (layer2_outputs[309]);
    assign outputs[12534] = (layer2_outputs[11057]) ^ (layer2_outputs[9836]);
    assign outputs[12535] = layer2_outputs[1207];
    assign outputs[12536] = ~((layer2_outputs[299]) ^ (layer2_outputs[6100]));
    assign outputs[12537] = (layer2_outputs[179]) & (layer2_outputs[9346]);
    assign outputs[12538] = ~(layer2_outputs[3469]);
    assign outputs[12539] = (layer2_outputs[2103]) | (layer2_outputs[777]);
    assign outputs[12540] = ~(layer2_outputs[5397]);
    assign outputs[12541] = layer2_outputs[7131];
    assign outputs[12542] = layer2_outputs[1721];
    assign outputs[12543] = ~((layer2_outputs[4581]) ^ (layer2_outputs[5654]));
    assign outputs[12544] = (layer2_outputs[10915]) & (layer2_outputs[5948]);
    assign outputs[12545] = (layer2_outputs[6169]) ^ (layer2_outputs[12212]);
    assign outputs[12546] = layer2_outputs[5436];
    assign outputs[12547] = ~((layer2_outputs[11404]) ^ (layer2_outputs[6219]));
    assign outputs[12548] = (layer2_outputs[692]) & ~(layer2_outputs[10142]);
    assign outputs[12549] = ~((layer2_outputs[1029]) & (layer2_outputs[5278]));
    assign outputs[12550] = ~(layer2_outputs[10139]);
    assign outputs[12551] = ~(layer2_outputs[7239]);
    assign outputs[12552] = layer2_outputs[3290];
    assign outputs[12553] = ~((layer2_outputs[3056]) & (layer2_outputs[4300]));
    assign outputs[12554] = ~(layer2_outputs[716]);
    assign outputs[12555] = ~((layer2_outputs[7555]) ^ (layer2_outputs[12205]));
    assign outputs[12556] = ~((layer2_outputs[620]) ^ (layer2_outputs[9892]));
    assign outputs[12557] = (layer2_outputs[3184]) ^ (layer2_outputs[4630]);
    assign outputs[12558] = ~((layer2_outputs[8248]) ^ (layer2_outputs[8460]));
    assign outputs[12559] = ~(layer2_outputs[2608]);
    assign outputs[12560] = ~((layer2_outputs[2859]) ^ (layer2_outputs[4364]));
    assign outputs[12561] = ~((layer2_outputs[10145]) ^ (layer2_outputs[11263]));
    assign outputs[12562] = ~((layer2_outputs[11636]) ^ (layer2_outputs[2242]));
    assign outputs[12563] = ~(layer2_outputs[11382]);
    assign outputs[12564] = layer2_outputs[7834];
    assign outputs[12565] = layer2_outputs[2406];
    assign outputs[12566] = ~((layer2_outputs[548]) | (layer2_outputs[5843]));
    assign outputs[12567] = (layer2_outputs[2809]) & (layer2_outputs[10207]);
    assign outputs[12568] = ~(layer2_outputs[7281]);
    assign outputs[12569] = (layer2_outputs[8239]) ^ (layer2_outputs[1048]);
    assign outputs[12570] = layer2_outputs[7295];
    assign outputs[12571] = layer2_outputs[7324];
    assign outputs[12572] = ~(layer2_outputs[11753]);
    assign outputs[12573] = (layer2_outputs[1157]) & ~(layer2_outputs[10928]);
    assign outputs[12574] = ~((layer2_outputs[1794]) & (layer2_outputs[404]));
    assign outputs[12575] = ~(layer2_outputs[1843]);
    assign outputs[12576] = ~((layer2_outputs[4071]) ^ (layer2_outputs[8762]));
    assign outputs[12577] = ~(layer2_outputs[10785]);
    assign outputs[12578] = ~(layer2_outputs[408]);
    assign outputs[12579] = layer2_outputs[11021];
    assign outputs[12580] = (layer2_outputs[7141]) ^ (layer2_outputs[12640]);
    assign outputs[12581] = ~(layer2_outputs[2681]);
    assign outputs[12582] = layer2_outputs[3057];
    assign outputs[12583] = ~((layer2_outputs[8608]) ^ (layer2_outputs[6503]));
    assign outputs[12584] = ~((layer2_outputs[7461]) ^ (layer2_outputs[2137]));
    assign outputs[12585] = (layer2_outputs[349]) ^ (layer2_outputs[1734]);
    assign outputs[12586] = (layer2_outputs[3626]) & (layer2_outputs[1721]);
    assign outputs[12587] = ~(layer2_outputs[7117]);
    assign outputs[12588] = (layer2_outputs[7170]) & ~(layer2_outputs[11512]);
    assign outputs[12589] = (layer2_outputs[7387]) | (layer2_outputs[6713]);
    assign outputs[12590] = ~((layer2_outputs[9959]) ^ (layer2_outputs[6426]));
    assign outputs[12591] = layer2_outputs[7524];
    assign outputs[12592] = (layer2_outputs[12553]) & ~(layer2_outputs[9275]);
    assign outputs[12593] = ~((layer2_outputs[5626]) & (layer2_outputs[4064]));
    assign outputs[12594] = ~((layer2_outputs[12632]) ^ (layer2_outputs[3125]));
    assign outputs[12595] = ~(layer2_outputs[7396]);
    assign outputs[12596] = ~(layer2_outputs[8157]);
    assign outputs[12597] = (layer2_outputs[650]) ^ (layer2_outputs[6749]);
    assign outputs[12598] = ~(layer2_outputs[9356]);
    assign outputs[12599] = (layer2_outputs[3531]) ^ (layer2_outputs[10346]);
    assign outputs[12600] = layer2_outputs[8816];
    assign outputs[12601] = (layer2_outputs[5648]) & ~(layer2_outputs[3598]);
    assign outputs[12602] = ~(layer2_outputs[2970]);
    assign outputs[12603] = ~((layer2_outputs[5750]) | (layer2_outputs[4266]));
    assign outputs[12604] = layer2_outputs[4555];
    assign outputs[12605] = ~(layer2_outputs[3672]);
    assign outputs[12606] = ~(layer2_outputs[824]);
    assign outputs[12607] = ~((layer2_outputs[602]) & (layer2_outputs[5075]));
    assign outputs[12608] = (layer2_outputs[1865]) ^ (layer2_outputs[7332]);
    assign outputs[12609] = (layer2_outputs[7885]) ^ (layer2_outputs[780]);
    assign outputs[12610] = layer2_outputs[12241];
    assign outputs[12611] = ~((layer2_outputs[5623]) ^ (layer2_outputs[11301]));
    assign outputs[12612] = layer2_outputs[7848];
    assign outputs[12613] = (layer2_outputs[8056]) & ~(layer2_outputs[5403]);
    assign outputs[12614] = ~(layer2_outputs[8509]);
    assign outputs[12615] = layer2_outputs[4096];
    assign outputs[12616] = (layer2_outputs[1068]) & ~(layer2_outputs[9414]);
    assign outputs[12617] = (layer2_outputs[8240]) ^ (layer2_outputs[5252]);
    assign outputs[12618] = layer2_outputs[402];
    assign outputs[12619] = layer2_outputs[10067];
    assign outputs[12620] = ~((layer2_outputs[8027]) | (layer2_outputs[11498]));
    assign outputs[12621] = (layer2_outputs[12654]) ^ (layer2_outputs[10999]);
    assign outputs[12622] = layer2_outputs[667];
    assign outputs[12623] = ~(layer2_outputs[4042]);
    assign outputs[12624] = ~((layer2_outputs[9966]) ^ (layer2_outputs[6518]));
    assign outputs[12625] = ~(layer2_outputs[401]);
    assign outputs[12626] = ~(layer2_outputs[804]);
    assign outputs[12627] = ~(layer2_outputs[11993]);
    assign outputs[12628] = layer2_outputs[2374];
    assign outputs[12629] = layer2_outputs[6997];
    assign outputs[12630] = (layer2_outputs[2178]) ^ (layer2_outputs[9115]);
    assign outputs[12631] = layer2_outputs[11911];
    assign outputs[12632] = ~((layer2_outputs[1661]) ^ (layer2_outputs[11230]));
    assign outputs[12633] = (layer2_outputs[872]) & ~(layer2_outputs[5683]);
    assign outputs[12634] = (layer2_outputs[8022]) ^ (layer2_outputs[1407]);
    assign outputs[12635] = ~((layer2_outputs[11981]) ^ (layer2_outputs[12054]));
    assign outputs[12636] = (layer2_outputs[9469]) & ~(layer2_outputs[9133]);
    assign outputs[12637] = ~(layer2_outputs[248]) | (layer2_outputs[8996]);
    assign outputs[12638] = (layer2_outputs[7258]) & (layer2_outputs[3417]);
    assign outputs[12639] = layer2_outputs[9380];
    assign outputs[12640] = layer2_outputs[6962];
    assign outputs[12641] = ~(layer2_outputs[7781]) | (layer2_outputs[8053]);
    assign outputs[12642] = ~((layer2_outputs[10658]) ^ (layer2_outputs[3477]));
    assign outputs[12643] = ~((layer2_outputs[8648]) ^ (layer2_outputs[6514]));
    assign outputs[12644] = (layer2_outputs[366]) & ~(layer2_outputs[12391]);
    assign outputs[12645] = ~((layer2_outputs[2547]) | (layer2_outputs[3736]));
    assign outputs[12646] = ~(layer2_outputs[157]);
    assign outputs[12647] = ~(layer2_outputs[2306]);
    assign outputs[12648] = layer2_outputs[8292];
    assign outputs[12649] = (layer2_outputs[3006]) & ~(layer2_outputs[12333]);
    assign outputs[12650] = ~((layer2_outputs[12772]) ^ (layer2_outputs[2427]));
    assign outputs[12651] = ~(layer2_outputs[12310]);
    assign outputs[12652] = ~((layer2_outputs[11908]) ^ (layer2_outputs[5537]));
    assign outputs[12653] = ~(layer2_outputs[2670]);
    assign outputs[12654] = layer2_outputs[10276];
    assign outputs[12655] = ~(layer2_outputs[8183]);
    assign outputs[12656] = (layer2_outputs[7513]) ^ (layer2_outputs[4940]);
    assign outputs[12657] = layer2_outputs[1823];
    assign outputs[12658] = (layer2_outputs[11810]) ^ (layer2_outputs[11214]);
    assign outputs[12659] = (layer2_outputs[3014]) ^ (layer2_outputs[5130]);
    assign outputs[12660] = ~(layer2_outputs[250]);
    assign outputs[12661] = (layer2_outputs[5293]) ^ (layer2_outputs[6524]);
    assign outputs[12662] = layer2_outputs[9036];
    assign outputs[12663] = (layer2_outputs[8470]) | (layer2_outputs[8188]);
    assign outputs[12664] = ~((layer2_outputs[5959]) ^ (layer2_outputs[6100]));
    assign outputs[12665] = ~(layer2_outputs[10757]);
    assign outputs[12666] = layer2_outputs[6645];
    assign outputs[12667] = (layer2_outputs[658]) ^ (layer2_outputs[2728]);
    assign outputs[12668] = layer2_outputs[2985];
    assign outputs[12669] = (layer2_outputs[6998]) & (layer2_outputs[11959]);
    assign outputs[12670] = ~(layer2_outputs[28]);
    assign outputs[12671] = layer2_outputs[9157];
    assign outputs[12672] = ~(layer2_outputs[3501]);
    assign outputs[12673] = layer2_outputs[341];
    assign outputs[12674] = ~(layer2_outputs[12620]);
    assign outputs[12675] = (layer2_outputs[2417]) | (layer2_outputs[488]);
    assign outputs[12676] = ~((layer2_outputs[11145]) ^ (layer2_outputs[1148]));
    assign outputs[12677] = (layer2_outputs[5547]) & (layer2_outputs[11853]);
    assign outputs[12678] = (layer2_outputs[6178]) & ~(layer2_outputs[10600]);
    assign outputs[12679] = (layer2_outputs[11827]) | (layer2_outputs[7941]);
    assign outputs[12680] = (layer2_outputs[5211]) & ~(layer2_outputs[5237]);
    assign outputs[12681] = (layer2_outputs[10633]) ^ (layer2_outputs[10982]);
    assign outputs[12682] = ~(layer2_outputs[5210]);
    assign outputs[12683] = layer2_outputs[8070];
    assign outputs[12684] = layer2_outputs[11036];
    assign outputs[12685] = layer2_outputs[1170];
    assign outputs[12686] = (layer2_outputs[6119]) & ~(layer2_outputs[11720]);
    assign outputs[12687] = ~(layer2_outputs[7254]);
    assign outputs[12688] = (layer2_outputs[1174]) ^ (layer2_outputs[10093]);
    assign outputs[12689] = ~((layer2_outputs[5640]) ^ (layer2_outputs[12478]));
    assign outputs[12690] = ~(layer2_outputs[253]);
    assign outputs[12691] = ~(layer2_outputs[4946]);
    assign outputs[12692] = layer2_outputs[1898];
    assign outputs[12693] = ~((layer2_outputs[3687]) ^ (layer2_outputs[409]));
    assign outputs[12694] = ~(layer2_outputs[11061]);
    assign outputs[12695] = ~((layer2_outputs[1582]) ^ (layer2_outputs[9162]));
    assign outputs[12696] = (layer2_outputs[5375]) | (layer2_outputs[6917]);
    assign outputs[12697] = ~(layer2_outputs[9494]) | (layer2_outputs[268]);
    assign outputs[12698] = (layer2_outputs[3607]) & ~(layer2_outputs[8374]);
    assign outputs[12699] = (layer2_outputs[5318]) ^ (layer2_outputs[1589]);
    assign outputs[12700] = ~((layer2_outputs[152]) ^ (layer2_outputs[6348]));
    assign outputs[12701] = ~((layer2_outputs[372]) ^ (layer2_outputs[7986]));
    assign outputs[12702] = (layer2_outputs[7782]) & (layer2_outputs[2751]);
    assign outputs[12703] = ~((layer2_outputs[722]) ^ (layer2_outputs[6800]));
    assign outputs[12704] = ~(layer2_outputs[10945]);
    assign outputs[12705] = ~((layer2_outputs[1074]) ^ (layer2_outputs[8305]));
    assign outputs[12706] = layer2_outputs[11271];
    assign outputs[12707] = layer2_outputs[8885];
    assign outputs[12708] = layer2_outputs[8293];
    assign outputs[12709] = (layer2_outputs[1552]) & (layer2_outputs[4520]);
    assign outputs[12710] = ~((layer2_outputs[1928]) ^ (layer2_outputs[2084]));
    assign outputs[12711] = layer2_outputs[1437];
    assign outputs[12712] = layer2_outputs[11051];
    assign outputs[12713] = ~(layer2_outputs[5186]);
    assign outputs[12714] = ~((layer2_outputs[9630]) ^ (layer2_outputs[3188]));
    assign outputs[12715] = ~(layer2_outputs[3064]);
    assign outputs[12716] = ~((layer2_outputs[11855]) ^ (layer2_outputs[9804]));
    assign outputs[12717] = (layer2_outputs[1271]) & (layer2_outputs[5680]);
    assign outputs[12718] = layer2_outputs[5942];
    assign outputs[12719] = layer2_outputs[1177];
    assign outputs[12720] = layer2_outputs[10366];
    assign outputs[12721] = (layer2_outputs[9002]) ^ (layer2_outputs[2807]);
    assign outputs[12722] = (layer2_outputs[10979]) ^ (layer2_outputs[11248]);
    assign outputs[12723] = ~(layer2_outputs[7104]);
    assign outputs[12724] = ~((layer2_outputs[7339]) ^ (layer2_outputs[6378]));
    assign outputs[12725] = (layer2_outputs[11940]) & ~(layer2_outputs[2429]);
    assign outputs[12726] = layer2_outputs[8564];
    assign outputs[12727] = layer2_outputs[11936];
    assign outputs[12728] = (layer2_outputs[9821]) ^ (layer2_outputs[9683]);
    assign outputs[12729] = ~(layer2_outputs[4003]);
    assign outputs[12730] = (layer2_outputs[11309]) ^ (layer2_outputs[5604]);
    assign outputs[12731] = (layer2_outputs[1591]) | (layer2_outputs[10159]);
    assign outputs[12732] = layer2_outputs[5434];
    assign outputs[12733] = ~(layer2_outputs[526]);
    assign outputs[12734] = ~(layer2_outputs[9026]) | (layer2_outputs[1970]);
    assign outputs[12735] = ~(layer2_outputs[8506]);
    assign outputs[12736] = (layer2_outputs[12418]) | (layer2_outputs[9821]);
    assign outputs[12737] = (layer2_outputs[2107]) | (layer2_outputs[8376]);
    assign outputs[12738] = (layer2_outputs[4182]) & (layer2_outputs[1408]);
    assign outputs[12739] = ~((layer2_outputs[864]) ^ (layer2_outputs[8747]));
    assign outputs[12740] = layer2_outputs[4688];
    assign outputs[12741] = ~((layer2_outputs[2465]) ^ (layer2_outputs[3272]));
    assign outputs[12742] = (layer2_outputs[3202]) ^ (layer2_outputs[3015]);
    assign outputs[12743] = layer2_outputs[5047];
    assign outputs[12744] = ~(layer2_outputs[10381]);
    assign outputs[12745] = (layer2_outputs[11232]) ^ (layer2_outputs[11253]);
    assign outputs[12746] = layer2_outputs[10350];
    assign outputs[12747] = ~(layer2_outputs[4454]);
    assign outputs[12748] = layer2_outputs[10177];
    assign outputs[12749] = layer2_outputs[10486];
    assign outputs[12750] = layer2_outputs[11748];
    assign outputs[12751] = layer2_outputs[529];
    assign outputs[12752] = ~(layer2_outputs[6508]) | (layer2_outputs[1832]);
    assign outputs[12753] = ~(layer2_outputs[3585]);
    assign outputs[12754] = layer2_outputs[6755];
    assign outputs[12755] = (layer2_outputs[106]) ^ (layer2_outputs[7280]);
    assign outputs[12756] = layer2_outputs[8998];
    assign outputs[12757] = ~(layer2_outputs[6009]);
    assign outputs[12758] = ~(layer2_outputs[8675]);
    assign outputs[12759] = ~((layer2_outputs[12556]) & (layer2_outputs[6665]));
    assign outputs[12760] = ~((layer2_outputs[10189]) ^ (layer2_outputs[6253]));
    assign outputs[12761] = ~(layer2_outputs[1505]);
    assign outputs[12762] = (layer2_outputs[11700]) & ~(layer2_outputs[7826]);
    assign outputs[12763] = layer2_outputs[1295];
    assign outputs[12764] = ~(layer2_outputs[10036]);
    assign outputs[12765] = ~((layer2_outputs[7543]) ^ (layer2_outputs[3012]));
    assign outputs[12766] = ~(layer2_outputs[10601]) | (layer2_outputs[7718]);
    assign outputs[12767] = ~(layer2_outputs[8848]);
    assign outputs[12768] = ~(layer2_outputs[6401]);
    assign outputs[12769] = layer2_outputs[8570];
    assign outputs[12770] = ~(layer2_outputs[7111]);
    assign outputs[12771] = ~(layer2_outputs[78]);
    assign outputs[12772] = ~(layer2_outputs[7161]);
    assign outputs[12773] = ~(layer2_outputs[1136]) | (layer2_outputs[2395]);
    assign outputs[12774] = layer2_outputs[9053];
    assign outputs[12775] = ~(layer2_outputs[765]);
    assign outputs[12776] = ~((layer2_outputs[3462]) ^ (layer2_outputs[6319]));
    assign outputs[12777] = ~((layer2_outputs[1031]) ^ (layer2_outputs[5863]));
    assign outputs[12778] = (layer2_outputs[11173]) & ~(layer2_outputs[9325]);
    assign outputs[12779] = layer2_outputs[2847];
    assign outputs[12780] = ~(layer2_outputs[2918]);
    assign outputs[12781] = ~((layer2_outputs[6666]) & (layer2_outputs[8356]));
    assign outputs[12782] = (layer2_outputs[5951]) ^ (layer2_outputs[3941]);
    assign outputs[12783] = ~(layer2_outputs[11811]);
    assign outputs[12784] = layer2_outputs[8869];
    assign outputs[12785] = ~(layer2_outputs[8124]);
    assign outputs[12786] = (layer2_outputs[12380]) ^ (layer2_outputs[10074]);
    assign outputs[12787] = ~(layer2_outputs[8102]);
    assign outputs[12788] = (layer2_outputs[360]) & ~(layer2_outputs[90]);
    assign outputs[12789] = (layer2_outputs[4435]) ^ (layer2_outputs[11019]);
    assign outputs[12790] = layer2_outputs[2598];
    assign outputs[12791] = (layer2_outputs[5860]) & (layer2_outputs[6752]);
    assign outputs[12792] = ~((layer2_outputs[9664]) ^ (layer2_outputs[45]));
    assign outputs[12793] = layer2_outputs[3027];
    assign outputs[12794] = ~(layer2_outputs[3452]);
    assign outputs[12795] = layer2_outputs[10427];
    assign outputs[12796] = ~(layer2_outputs[11737]);
    assign outputs[12797] = (layer2_outputs[12561]) & ~(layer2_outputs[4439]);
    assign outputs[12798] = layer2_outputs[6690];
    assign outputs[12799] = (layer2_outputs[3714]) ^ (layer2_outputs[7591]);
endmodule
