library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(2559 downto 0);
    signal layer1_outputs : std_logic_vector(2559 downto 0);
    signal layer2_outputs : std_logic_vector(2559 downto 0);
    signal layer3_outputs : std_logic_vector(2559 downto 0);
    signal layer4_outputs : std_logic_vector(2559 downto 0);
    signal layer5_outputs : std_logic_vector(2559 downto 0);
    signal layer6_outputs : std_logic_vector(2559 downto 0);

begin

    layer0_outputs(0) <= (inputs(254)) and (inputs(43));
    layer0_outputs(1) <= (inputs(235)) xor (inputs(140));
    layer0_outputs(2) <= not(inputs(24)) or (inputs(27));
    layer0_outputs(3) <= '0';
    layer0_outputs(4) <= not(inputs(43));
    layer0_outputs(5) <= inputs(146);
    layer0_outputs(6) <= not((inputs(143)) xor (inputs(174)));
    layer0_outputs(7) <= not(inputs(255)) or (inputs(0));
    layer0_outputs(8) <= '1';
    layer0_outputs(9) <= '1';
    layer0_outputs(10) <= not(inputs(111));
    layer0_outputs(11) <= (inputs(58)) or (inputs(126));
    layer0_outputs(12) <= (inputs(221)) or (inputs(1));
    layer0_outputs(13) <= (inputs(216)) or (inputs(224));
    layer0_outputs(14) <= inputs(30);
    layer0_outputs(15) <= '1';
    layer0_outputs(16) <= not(inputs(69)) or (inputs(3));
    layer0_outputs(17) <= (inputs(86)) and not (inputs(30));
    layer0_outputs(18) <= not(inputs(124));
    layer0_outputs(19) <= not((inputs(193)) or (inputs(224)));
    layer0_outputs(20) <= not(inputs(179));
    layer0_outputs(21) <= '1';
    layer0_outputs(22) <= (inputs(75)) xor (inputs(46));
    layer0_outputs(23) <= (inputs(55)) or (inputs(113));
    layer0_outputs(24) <= '0';
    layer0_outputs(25) <= not(inputs(223));
    layer0_outputs(26) <= not(inputs(252)) or (inputs(42));
    layer0_outputs(27) <= (inputs(121)) and not (inputs(242));
    layer0_outputs(28) <= not(inputs(210));
    layer0_outputs(29) <= '0';
    layer0_outputs(30) <= inputs(135);
    layer0_outputs(31) <= '1';
    layer0_outputs(32) <= (inputs(255)) xor (inputs(75));
    layer0_outputs(33) <= inputs(133);
    layer0_outputs(34) <= (inputs(220)) xor (inputs(173));
    layer0_outputs(35) <= '1';
    layer0_outputs(36) <= '1';
    layer0_outputs(37) <= (inputs(236)) and not (inputs(202));
    layer0_outputs(38) <= not(inputs(221));
    layer0_outputs(39) <= not((inputs(207)) or (inputs(193)));
    layer0_outputs(40) <= not(inputs(222));
    layer0_outputs(41) <= '0';
    layer0_outputs(42) <= inputs(102);
    layer0_outputs(43) <= (inputs(38)) or (inputs(101));
    layer0_outputs(44) <= (inputs(187)) or (inputs(189));
    layer0_outputs(45) <= '0';
    layer0_outputs(46) <= (inputs(218)) or (inputs(208));
    layer0_outputs(47) <= '0';
    layer0_outputs(48) <= '0';
    layer0_outputs(49) <= '0';
    layer0_outputs(50) <= not(inputs(205));
    layer0_outputs(51) <= (inputs(109)) or (inputs(159));
    layer0_outputs(52) <= not((inputs(33)) and (inputs(46)));
    layer0_outputs(53) <= not(inputs(167));
    layer0_outputs(54) <= (inputs(190)) or (inputs(141));
    layer0_outputs(55) <= inputs(60);
    layer0_outputs(56) <= inputs(151);
    layer0_outputs(57) <= '1';
    layer0_outputs(58) <= inputs(153);
    layer0_outputs(59) <= (inputs(157)) and (inputs(32));
    layer0_outputs(60) <= (inputs(207)) and not (inputs(97));
    layer0_outputs(61) <= not(inputs(119));
    layer0_outputs(62) <= not((inputs(145)) and (inputs(166)));
    layer0_outputs(63) <= '1';
    layer0_outputs(64) <= '0';
    layer0_outputs(65) <= (inputs(200)) and not (inputs(46));
    layer0_outputs(66) <= not(inputs(115)) or (inputs(152));
    layer0_outputs(67) <= (inputs(120)) or (inputs(105));
    layer0_outputs(68) <= inputs(149);
    layer0_outputs(69) <= (inputs(173)) or (inputs(210));
    layer0_outputs(70) <= not(inputs(44)) or (inputs(137));
    layer0_outputs(71) <= '0';
    layer0_outputs(72) <= inputs(167);
    layer0_outputs(73) <= (inputs(176)) xor (inputs(82));
    layer0_outputs(74) <= not(inputs(134));
    layer0_outputs(75) <= not((inputs(109)) and (inputs(5)));
    layer0_outputs(76) <= (inputs(185)) and not (inputs(64));
    layer0_outputs(77) <= (inputs(99)) or (inputs(107));
    layer0_outputs(78) <= '1';
    layer0_outputs(79) <= '1';
    layer0_outputs(80) <= not(inputs(1)) or (inputs(22));
    layer0_outputs(81) <= '0';
    layer0_outputs(82) <= '1';
    layer0_outputs(83) <= (inputs(207)) and not (inputs(17));
    layer0_outputs(84) <= '1';
    layer0_outputs(85) <= '1';
    layer0_outputs(86) <= (inputs(133)) and (inputs(12));
    layer0_outputs(87) <= inputs(111);
    layer0_outputs(88) <= not(inputs(79));
    layer0_outputs(89) <= not((inputs(240)) and (inputs(244)));
    layer0_outputs(90) <= (inputs(196)) or (inputs(213));
    layer0_outputs(91) <= '0';
    layer0_outputs(92) <= (inputs(142)) or (inputs(217));
    layer0_outputs(93) <= (inputs(43)) or (inputs(58));
    layer0_outputs(94) <= (inputs(203)) and (inputs(152));
    layer0_outputs(95) <= (inputs(221)) and not (inputs(94));
    layer0_outputs(96) <= inputs(195);
    layer0_outputs(97) <= (inputs(154)) or (inputs(204));
    layer0_outputs(98) <= not(inputs(136));
    layer0_outputs(99) <= (inputs(90)) and (inputs(135));
    layer0_outputs(100) <= not(inputs(62));
    layer0_outputs(101) <= '1';
    layer0_outputs(102) <= (inputs(58)) and (inputs(138));
    layer0_outputs(103) <= (inputs(244)) and not (inputs(29));
    layer0_outputs(104) <= '1';
    layer0_outputs(105) <= not((inputs(111)) or (inputs(43)));
    layer0_outputs(106) <= '1';
    layer0_outputs(107) <= not((inputs(166)) or (inputs(102)));
    layer0_outputs(108) <= '0';
    layer0_outputs(109) <= (inputs(246)) and not (inputs(151));
    layer0_outputs(110) <= (inputs(180)) and not (inputs(98));
    layer0_outputs(111) <= not(inputs(165));
    layer0_outputs(112) <= not(inputs(179)) or (inputs(213));
    layer0_outputs(113) <= (inputs(164)) or (inputs(88));
    layer0_outputs(114) <= not((inputs(2)) or (inputs(140)));
    layer0_outputs(115) <= not((inputs(209)) or (inputs(31)));
    layer0_outputs(116) <= not(inputs(115)) or (inputs(106));
    layer0_outputs(117) <= '1';
    layer0_outputs(118) <= '1';
    layer0_outputs(119) <= inputs(249);
    layer0_outputs(120) <= not(inputs(59)) or (inputs(62));
    layer0_outputs(121) <= inputs(192);
    layer0_outputs(122) <= not((inputs(146)) or (inputs(235)));
    layer0_outputs(123) <= not(inputs(6));
    layer0_outputs(124) <= (inputs(107)) or (inputs(29));
    layer0_outputs(125) <= '1';
    layer0_outputs(126) <= '1';
    layer0_outputs(127) <= not(inputs(33)) or (inputs(132));
    layer0_outputs(128) <= not((inputs(98)) or (inputs(192)));
    layer0_outputs(129) <= not(inputs(71)) or (inputs(50));
    layer0_outputs(130) <= not((inputs(47)) or (inputs(252)));
    layer0_outputs(131) <= (inputs(78)) or (inputs(61));
    layer0_outputs(132) <= not((inputs(246)) or (inputs(160)));
    layer0_outputs(133) <= not((inputs(203)) or (inputs(160)));
    layer0_outputs(134) <= inputs(142);
    layer0_outputs(135) <= not(inputs(86)) or (inputs(74));
    layer0_outputs(136) <= inputs(126);
    layer0_outputs(137) <= '1';
    layer0_outputs(138) <= (inputs(97)) and (inputs(31));
    layer0_outputs(139) <= '0';
    layer0_outputs(140) <= not(inputs(118));
    layer0_outputs(141) <= (inputs(148)) and (inputs(219));
    layer0_outputs(142) <= not(inputs(209));
    layer0_outputs(143) <= not(inputs(55));
    layer0_outputs(144) <= (inputs(2)) or (inputs(234));
    layer0_outputs(145) <= '1';
    layer0_outputs(146) <= inputs(31);
    layer0_outputs(147) <= not(inputs(7)) or (inputs(13));
    layer0_outputs(148) <= not(inputs(143));
    layer0_outputs(149) <= not((inputs(215)) and (inputs(156)));
    layer0_outputs(150) <= (inputs(114)) or (inputs(201));
    layer0_outputs(151) <= not(inputs(162));
    layer0_outputs(152) <= '0';
    layer0_outputs(153) <= not(inputs(22));
    layer0_outputs(154) <= (inputs(116)) or (inputs(52));
    layer0_outputs(155) <= inputs(113);
    layer0_outputs(156) <= (inputs(25)) and not (inputs(85));
    layer0_outputs(157) <= inputs(24);
    layer0_outputs(158) <= '0';
    layer0_outputs(159) <= (inputs(34)) and not (inputs(158));
    layer0_outputs(160) <= not((inputs(206)) or (inputs(147)));
    layer0_outputs(161) <= not(inputs(11)) or (inputs(73));
    layer0_outputs(162) <= not(inputs(77));
    layer0_outputs(163) <= (inputs(121)) and not (inputs(87));
    layer0_outputs(164) <= not((inputs(169)) and (inputs(230)));
    layer0_outputs(165) <= inputs(110);
    layer0_outputs(166) <= (inputs(193)) and (inputs(4));
    layer0_outputs(167) <= not(inputs(96)) or (inputs(205));
    layer0_outputs(168) <= inputs(132);
    layer0_outputs(169) <= not(inputs(236)) or (inputs(238));
    layer0_outputs(170) <= '1';
    layer0_outputs(171) <= not(inputs(150));
    layer0_outputs(172) <= not(inputs(34)) or (inputs(115));
    layer0_outputs(173) <= not(inputs(233)) or (inputs(238));
    layer0_outputs(174) <= (inputs(22)) xor (inputs(133));
    layer0_outputs(175) <= (inputs(159)) and (inputs(183));
    layer0_outputs(176) <= '1';
    layer0_outputs(177) <= inputs(211);
    layer0_outputs(178) <= '1';
    layer0_outputs(179) <= inputs(161);
    layer0_outputs(180) <= not((inputs(226)) and (inputs(28)));
    layer0_outputs(181) <= not(inputs(212));
    layer0_outputs(182) <= '1';
    layer0_outputs(183) <= not(inputs(130)) or (inputs(136));
    layer0_outputs(184) <= (inputs(94)) and not (inputs(70));
    layer0_outputs(185) <= not((inputs(75)) or (inputs(92)));
    layer0_outputs(186) <= not(inputs(141));
    layer0_outputs(187) <= not(inputs(255)) or (inputs(159));
    layer0_outputs(188) <= inputs(85);
    layer0_outputs(189) <= not(inputs(164)) or (inputs(125));
    layer0_outputs(190) <= inputs(191);
    layer0_outputs(191) <= not(inputs(148)) or (inputs(39));
    layer0_outputs(192) <= not(inputs(100));
    layer0_outputs(193) <= '0';
    layer0_outputs(194) <= (inputs(81)) and (inputs(104));
    layer0_outputs(195) <= (inputs(32)) and not (inputs(153));
    layer0_outputs(196) <= '0';
    layer0_outputs(197) <= (inputs(170)) and (inputs(142));
    layer0_outputs(198) <= (inputs(253)) or (inputs(226));
    layer0_outputs(199) <= not((inputs(238)) or (inputs(135)));
    layer0_outputs(200) <= (inputs(227)) or (inputs(153));
    layer0_outputs(201) <= '0';
    layer0_outputs(202) <= (inputs(94)) xor (inputs(61));
    layer0_outputs(203) <= (inputs(144)) and not (inputs(33));
    layer0_outputs(204) <= not((inputs(189)) and (inputs(163)));
    layer0_outputs(205) <= not(inputs(196));
    layer0_outputs(206) <= not(inputs(32)) or (inputs(220));
    layer0_outputs(207) <= not((inputs(90)) or (inputs(225)));
    layer0_outputs(208) <= (inputs(140)) and not (inputs(118));
    layer0_outputs(209) <= (inputs(187)) or (inputs(130));
    layer0_outputs(210) <= '0';
    layer0_outputs(211) <= '1';
    layer0_outputs(212) <= (inputs(156)) and (inputs(101));
    layer0_outputs(213) <= not(inputs(93));
    layer0_outputs(214) <= '1';
    layer0_outputs(215) <= (inputs(149)) and (inputs(150));
    layer0_outputs(216) <= inputs(2);
    layer0_outputs(217) <= '1';
    layer0_outputs(218) <= not(inputs(104));
    layer0_outputs(219) <= not((inputs(137)) or (inputs(251)));
    layer0_outputs(220) <= inputs(16);
    layer0_outputs(221) <= (inputs(35)) and not (inputs(10));
    layer0_outputs(222) <= '0';
    layer0_outputs(223) <= not(inputs(198)) or (inputs(231));
    layer0_outputs(224) <= inputs(45);
    layer0_outputs(225) <= '1';
    layer0_outputs(226) <= (inputs(173)) and not (inputs(12));
    layer0_outputs(227) <= not(inputs(157));
    layer0_outputs(228) <= not((inputs(28)) and (inputs(75)));
    layer0_outputs(229) <= not(inputs(21)) or (inputs(65));
    layer0_outputs(230) <= not(inputs(228));
    layer0_outputs(231) <= (inputs(35)) and not (inputs(126));
    layer0_outputs(232) <= not((inputs(34)) or (inputs(145)));
    layer0_outputs(233) <= (inputs(67)) and not (inputs(235));
    layer0_outputs(234) <= not((inputs(35)) xor (inputs(11)));
    layer0_outputs(235) <= not(inputs(188)) or (inputs(184));
    layer0_outputs(236) <= (inputs(154)) and (inputs(102));
    layer0_outputs(237) <= not(inputs(214));
    layer0_outputs(238) <= not((inputs(223)) or (inputs(106)));
    layer0_outputs(239) <= (inputs(103)) and not (inputs(175));
    layer0_outputs(240) <= not(inputs(12)) or (inputs(130));
    layer0_outputs(241) <= '0';
    layer0_outputs(242) <= not(inputs(231));
    layer0_outputs(243) <= (inputs(128)) and not (inputs(236));
    layer0_outputs(244) <= '1';
    layer0_outputs(245) <= (inputs(143)) xor (inputs(101));
    layer0_outputs(246) <= not(inputs(191));
    layer0_outputs(247) <= not((inputs(134)) or (inputs(137)));
    layer0_outputs(248) <= (inputs(14)) and not (inputs(131));
    layer0_outputs(249) <= '0';
    layer0_outputs(250) <= not(inputs(154));
    layer0_outputs(251) <= inputs(105);
    layer0_outputs(252) <= not((inputs(144)) or (inputs(185)));
    layer0_outputs(253) <= not(inputs(190));
    layer0_outputs(254) <= '1';
    layer0_outputs(255) <= not((inputs(111)) or (inputs(122)));
    layer0_outputs(256) <= inputs(228);
    layer0_outputs(257) <= not(inputs(63)) or (inputs(2));
    layer0_outputs(258) <= '0';
    layer0_outputs(259) <= (inputs(99)) or (inputs(129));
    layer0_outputs(260) <= not(inputs(6)) or (inputs(247));
    layer0_outputs(261) <= (inputs(230)) and (inputs(231));
    layer0_outputs(262) <= inputs(105);
    layer0_outputs(263) <= not((inputs(232)) and (inputs(45)));
    layer0_outputs(264) <= '0';
    layer0_outputs(265) <= '1';
    layer0_outputs(266) <= inputs(167);
    layer0_outputs(267) <= (inputs(179)) and not (inputs(44));
    layer0_outputs(268) <= '0';
    layer0_outputs(269) <= (inputs(88)) and not (inputs(238));
    layer0_outputs(270) <= (inputs(13)) or (inputs(104));
    layer0_outputs(271) <= not(inputs(165));
    layer0_outputs(272) <= (inputs(108)) or (inputs(161));
    layer0_outputs(273) <= inputs(228);
    layer0_outputs(274) <= not(inputs(221)) or (inputs(66));
    layer0_outputs(275) <= inputs(19);
    layer0_outputs(276) <= inputs(180);
    layer0_outputs(277) <= not((inputs(168)) or (inputs(152)));
    layer0_outputs(278) <= (inputs(241)) and not (inputs(112));
    layer0_outputs(279) <= '1';
    layer0_outputs(280) <= not((inputs(159)) and (inputs(225)));
    layer0_outputs(281) <= inputs(131);
    layer0_outputs(282) <= '0';
    layer0_outputs(283) <= not(inputs(21)) or (inputs(144));
    layer0_outputs(284) <= '0';
    layer0_outputs(285) <= inputs(115);
    layer0_outputs(286) <= not((inputs(126)) and (inputs(10)));
    layer0_outputs(287) <= not(inputs(23)) or (inputs(45));
    layer0_outputs(288) <= '0';
    layer0_outputs(289) <= inputs(3);
    layer0_outputs(290) <= not(inputs(71));
    layer0_outputs(291) <= '0';
    layer0_outputs(292) <= not((inputs(218)) or (inputs(177)));
    layer0_outputs(293) <= (inputs(122)) and (inputs(89));
    layer0_outputs(294) <= inputs(92);
    layer0_outputs(295) <= not(inputs(209)) or (inputs(60));
    layer0_outputs(296) <= inputs(247);
    layer0_outputs(297) <= not((inputs(177)) or (inputs(171)));
    layer0_outputs(298) <= '1';
    layer0_outputs(299) <= '1';
    layer0_outputs(300) <= '0';
    layer0_outputs(301) <= not(inputs(62)) or (inputs(171));
    layer0_outputs(302) <= not(inputs(92));
    layer0_outputs(303) <= not(inputs(16));
    layer0_outputs(304) <= (inputs(95)) or (inputs(209));
    layer0_outputs(305) <= (inputs(228)) and not (inputs(95));
    layer0_outputs(306) <= not(inputs(221)) or (inputs(241));
    layer0_outputs(307) <= (inputs(163)) or (inputs(178));
    layer0_outputs(308) <= not(inputs(232));
    layer0_outputs(309) <= not(inputs(163));
    layer0_outputs(310) <= not(inputs(218)) or (inputs(124));
    layer0_outputs(311) <= (inputs(83)) and not (inputs(62));
    layer0_outputs(312) <= not((inputs(69)) or (inputs(39)));
    layer0_outputs(313) <= '0';
    layer0_outputs(314) <= (inputs(50)) and not (inputs(253));
    layer0_outputs(315) <= not(inputs(114));
    layer0_outputs(316) <= '0';
    layer0_outputs(317) <= '0';
    layer0_outputs(318) <= inputs(20);
    layer0_outputs(319) <= inputs(61);
    layer0_outputs(320) <= inputs(146);
    layer0_outputs(321) <= inputs(107);
    layer0_outputs(322) <= (inputs(191)) and not (inputs(73));
    layer0_outputs(323) <= '0';
    layer0_outputs(324) <= not((inputs(181)) xor (inputs(191)));
    layer0_outputs(325) <= (inputs(199)) and not (inputs(127));
    layer0_outputs(326) <= (inputs(123)) or (inputs(137));
    layer0_outputs(327) <= '0';
    layer0_outputs(328) <= inputs(113);
    layer0_outputs(329) <= (inputs(178)) and (inputs(141));
    layer0_outputs(330) <= not(inputs(72));
    layer0_outputs(331) <= (inputs(112)) and not (inputs(151));
    layer0_outputs(332) <= (inputs(227)) or (inputs(143));
    layer0_outputs(333) <= '1';
    layer0_outputs(334) <= '1';
    layer0_outputs(335) <= not(inputs(22));
    layer0_outputs(336) <= (inputs(254)) and not (inputs(50));
    layer0_outputs(337) <= '0';
    layer0_outputs(338) <= not((inputs(175)) or (inputs(221)));
    layer0_outputs(339) <= '1';
    layer0_outputs(340) <= not(inputs(110));
    layer0_outputs(341) <= not((inputs(205)) xor (inputs(76)));
    layer0_outputs(342) <= not((inputs(29)) and (inputs(37)));
    layer0_outputs(343) <= not((inputs(162)) and (inputs(124)));
    layer0_outputs(344) <= '0';
    layer0_outputs(345) <= (inputs(82)) or (inputs(99));
    layer0_outputs(346) <= inputs(145);
    layer0_outputs(347) <= (inputs(37)) or (inputs(253));
    layer0_outputs(348) <= not(inputs(145));
    layer0_outputs(349) <= '1';
    layer0_outputs(350) <= not((inputs(215)) and (inputs(159)));
    layer0_outputs(351) <= (inputs(148)) or (inputs(63));
    layer0_outputs(352) <= (inputs(187)) and not (inputs(154));
    layer0_outputs(353) <= (inputs(113)) or (inputs(185));
    layer0_outputs(354) <= inputs(131);
    layer0_outputs(355) <= '0';
    layer0_outputs(356) <= not(inputs(101)) or (inputs(105));
    layer0_outputs(357) <= (inputs(211)) or (inputs(179));
    layer0_outputs(358) <= '0';
    layer0_outputs(359) <= not((inputs(144)) or (inputs(244)));
    layer0_outputs(360) <= not(inputs(106));
    layer0_outputs(361) <= not(inputs(12)) or (inputs(33));
    layer0_outputs(362) <= (inputs(73)) or (inputs(237));
    layer0_outputs(363) <= not((inputs(113)) xor (inputs(166)));
    layer0_outputs(364) <= '1';
    layer0_outputs(365) <= not((inputs(57)) or (inputs(12)));
    layer0_outputs(366) <= not(inputs(84)) or (inputs(122));
    layer0_outputs(367) <= not(inputs(58)) or (inputs(214));
    layer0_outputs(368) <= not((inputs(49)) and (inputs(131)));
    layer0_outputs(369) <= '1';
    layer0_outputs(370) <= inputs(91);
    layer0_outputs(371) <= not(inputs(159)) or (inputs(30));
    layer0_outputs(372) <= inputs(243);
    layer0_outputs(373) <= (inputs(91)) and not (inputs(204));
    layer0_outputs(374) <= '1';
    layer0_outputs(375) <= not(inputs(117));
    layer0_outputs(376) <= '0';
    layer0_outputs(377) <= not(inputs(106)) or (inputs(207));
    layer0_outputs(378) <= not(inputs(227)) or (inputs(31));
    layer0_outputs(379) <= not(inputs(3)) or (inputs(217));
    layer0_outputs(380) <= inputs(124);
    layer0_outputs(381) <= (inputs(113)) xor (inputs(100));
    layer0_outputs(382) <= '0';
    layer0_outputs(383) <= not((inputs(197)) or (inputs(149)));
    layer0_outputs(384) <= '0';
    layer0_outputs(385) <= (inputs(159)) xor (inputs(23));
    layer0_outputs(386) <= not(inputs(12)) or (inputs(97));
    layer0_outputs(387) <= not(inputs(190));
    layer0_outputs(388) <= (inputs(15)) and not (inputs(118));
    layer0_outputs(389) <= '0';
    layer0_outputs(390) <= inputs(150);
    layer0_outputs(391) <= (inputs(249)) or (inputs(202));
    layer0_outputs(392) <= '1';
    layer0_outputs(393) <= not((inputs(217)) and (inputs(252)));
    layer0_outputs(394) <= not(inputs(38)) or (inputs(135));
    layer0_outputs(395) <= not((inputs(46)) and (inputs(109)));
    layer0_outputs(396) <= not(inputs(63));
    layer0_outputs(397) <= '0';
    layer0_outputs(398) <= '0';
    layer0_outputs(399) <= not(inputs(217));
    layer0_outputs(400) <= (inputs(203)) and not (inputs(58));
    layer0_outputs(401) <= '0';
    layer0_outputs(402) <= not(inputs(13)) or (inputs(193));
    layer0_outputs(403) <= '0';
    layer0_outputs(404) <= (inputs(150)) or (inputs(102));
    layer0_outputs(405) <= inputs(173);
    layer0_outputs(406) <= inputs(60);
    layer0_outputs(407) <= '1';
    layer0_outputs(408) <= (inputs(90)) and not (inputs(236));
    layer0_outputs(409) <= inputs(34);
    layer0_outputs(410) <= not(inputs(121));
    layer0_outputs(411) <= (inputs(207)) or (inputs(138));
    layer0_outputs(412) <= not(inputs(85));
    layer0_outputs(413) <= '0';
    layer0_outputs(414) <= not(inputs(144));
    layer0_outputs(415) <= inputs(88);
    layer0_outputs(416) <= inputs(141);
    layer0_outputs(417) <= '0';
    layer0_outputs(418) <= not(inputs(219)) or (inputs(222));
    layer0_outputs(419) <= (inputs(169)) and not (inputs(20));
    layer0_outputs(420) <= not(inputs(55));
    layer0_outputs(421) <= not(inputs(126));
    layer0_outputs(422) <= '0';
    layer0_outputs(423) <= '1';
    layer0_outputs(424) <= inputs(32);
    layer0_outputs(425) <= not(inputs(94));
    layer0_outputs(426) <= not(inputs(226));
    layer0_outputs(427) <= '0';
    layer0_outputs(428) <= '1';
    layer0_outputs(429) <= '1';
    layer0_outputs(430) <= not((inputs(224)) or (inputs(110)));
    layer0_outputs(431) <= (inputs(142)) and not (inputs(148));
    layer0_outputs(432) <= inputs(34);
    layer0_outputs(433) <= not(inputs(229)) or (inputs(2));
    layer0_outputs(434) <= '1';
    layer0_outputs(435) <= (inputs(44)) or (inputs(49));
    layer0_outputs(436) <= inputs(215);
    layer0_outputs(437) <= '1';
    layer0_outputs(438) <= (inputs(50)) or (inputs(188));
    layer0_outputs(439) <= '1';
    layer0_outputs(440) <= (inputs(80)) and (inputs(162));
    layer0_outputs(441) <= not((inputs(166)) and (inputs(153)));
    layer0_outputs(442) <= not(inputs(91));
    layer0_outputs(443) <= (inputs(26)) and not (inputs(211));
    layer0_outputs(444) <= inputs(85);
    layer0_outputs(445) <= inputs(116);
    layer0_outputs(446) <= (inputs(128)) or (inputs(104));
    layer0_outputs(447) <= not((inputs(234)) or (inputs(26)));
    layer0_outputs(448) <= '1';
    layer0_outputs(449) <= not(inputs(99));
    layer0_outputs(450) <= inputs(132);
    layer0_outputs(451) <= (inputs(197)) and (inputs(108));
    layer0_outputs(452) <= not(inputs(161)) or (inputs(77));
    layer0_outputs(453) <= (inputs(23)) or (inputs(180));
    layer0_outputs(454) <= '1';
    layer0_outputs(455) <= not((inputs(202)) and (inputs(192)));
    layer0_outputs(456) <= '1';
    layer0_outputs(457) <= not((inputs(23)) and (inputs(34)));
    layer0_outputs(458) <= '1';
    layer0_outputs(459) <= not(inputs(130)) or (inputs(151));
    layer0_outputs(460) <= inputs(111);
    layer0_outputs(461) <= (inputs(120)) and not (inputs(208));
    layer0_outputs(462) <= not(inputs(174)) or (inputs(40));
    layer0_outputs(463) <= not(inputs(96));
    layer0_outputs(464) <= (inputs(194)) xor (inputs(204));
    layer0_outputs(465) <= not(inputs(183));
    layer0_outputs(466) <= not(inputs(234));
    layer0_outputs(467) <= (inputs(176)) and (inputs(222));
    layer0_outputs(468) <= inputs(65);
    layer0_outputs(469) <= not(inputs(94));
    layer0_outputs(470) <= inputs(100);
    layer0_outputs(471) <= '1';
    layer0_outputs(472) <= not(inputs(167)) or (inputs(208));
    layer0_outputs(473) <= '0';
    layer0_outputs(474) <= not((inputs(57)) and (inputs(236)));
    layer0_outputs(475) <= inputs(126);
    layer0_outputs(476) <= not(inputs(234));
    layer0_outputs(477) <= inputs(199);
    layer0_outputs(478) <= not((inputs(181)) or (inputs(164)));
    layer0_outputs(479) <= inputs(135);
    layer0_outputs(480) <= not(inputs(166));
    layer0_outputs(481) <= not((inputs(132)) or (inputs(161)));
    layer0_outputs(482) <= '1';
    layer0_outputs(483) <= inputs(150);
    layer0_outputs(484) <= not(inputs(91));
    layer0_outputs(485) <= not(inputs(141)) or (inputs(3));
    layer0_outputs(486) <= (inputs(215)) and (inputs(171));
    layer0_outputs(487) <= inputs(42);
    layer0_outputs(488) <= '1';
    layer0_outputs(489) <= (inputs(32)) xor (inputs(1));
    layer0_outputs(490) <= (inputs(20)) and not (inputs(107));
    layer0_outputs(491) <= '0';
    layer0_outputs(492) <= (inputs(235)) and not (inputs(93));
    layer0_outputs(493) <= '0';
    layer0_outputs(494) <= inputs(99);
    layer0_outputs(495) <= not((inputs(67)) and (inputs(0)));
    layer0_outputs(496) <= (inputs(122)) or (inputs(207));
    layer0_outputs(497) <= (inputs(231)) or (inputs(207));
    layer0_outputs(498) <= not((inputs(154)) or (inputs(101)));
    layer0_outputs(499) <= (inputs(242)) and not (inputs(22));
    layer0_outputs(500) <= not((inputs(184)) and (inputs(82)));
    layer0_outputs(501) <= '1';
    layer0_outputs(502) <= inputs(1);
    layer0_outputs(503) <= '0';
    layer0_outputs(504) <= not(inputs(95));
    layer0_outputs(505) <= not((inputs(36)) or (inputs(65)));
    layer0_outputs(506) <= not((inputs(79)) or (inputs(160)));
    layer0_outputs(507) <= (inputs(88)) xor (inputs(96));
    layer0_outputs(508) <= not(inputs(93)) or (inputs(119));
    layer0_outputs(509) <= '0';
    layer0_outputs(510) <= not(inputs(77));
    layer0_outputs(511) <= (inputs(108)) and not (inputs(24));
    layer0_outputs(512) <= (inputs(74)) and (inputs(77));
    layer0_outputs(513) <= not((inputs(219)) or (inputs(1)));
    layer0_outputs(514) <= (inputs(145)) or (inputs(4));
    layer0_outputs(515) <= not(inputs(115)) or (inputs(26));
    layer0_outputs(516) <= not(inputs(102));
    layer0_outputs(517) <= not(inputs(44));
    layer0_outputs(518) <= inputs(120);
    layer0_outputs(519) <= not((inputs(141)) or (inputs(39)));
    layer0_outputs(520) <= (inputs(238)) and not (inputs(99));
    layer0_outputs(521) <= '0';
    layer0_outputs(522) <= (inputs(101)) or (inputs(247));
    layer0_outputs(523) <= not(inputs(50)) or (inputs(15));
    layer0_outputs(524) <= not(inputs(202)) or (inputs(52));
    layer0_outputs(525) <= not(inputs(198));
    layer0_outputs(526) <= (inputs(65)) xor (inputs(65));
    layer0_outputs(527) <= '0';
    layer0_outputs(528) <= not(inputs(0)) or (inputs(150));
    layer0_outputs(529) <= not(inputs(150));
    layer0_outputs(530) <= '1';
    layer0_outputs(531) <= '1';
    layer0_outputs(532) <= not(inputs(249));
    layer0_outputs(533) <= (inputs(72)) and not (inputs(227));
    layer0_outputs(534) <= inputs(46);
    layer0_outputs(535) <= (inputs(242)) and not (inputs(148));
    layer0_outputs(536) <= (inputs(174)) or (inputs(181));
    layer0_outputs(537) <= not((inputs(55)) or (inputs(167)));
    layer0_outputs(538) <= not(inputs(107));
    layer0_outputs(539) <= not((inputs(255)) and (inputs(114)));
    layer0_outputs(540) <= not(inputs(239)) or (inputs(250));
    layer0_outputs(541) <= '1';
    layer0_outputs(542) <= (inputs(71)) and not (inputs(126));
    layer0_outputs(543) <= inputs(119);
    layer0_outputs(544) <= '0';
    layer0_outputs(545) <= not(inputs(240)) or (inputs(206));
    layer0_outputs(546) <= (inputs(81)) and not (inputs(169));
    layer0_outputs(547) <= not((inputs(10)) and (inputs(76)));
    layer0_outputs(548) <= inputs(165);
    layer0_outputs(549) <= not(inputs(247));
    layer0_outputs(550) <= '1';
    layer0_outputs(551) <= (inputs(99)) or (inputs(37));
    layer0_outputs(552) <= (inputs(187)) xor (inputs(83));
    layer0_outputs(553) <= '0';
    layer0_outputs(554) <= not(inputs(252));
    layer0_outputs(555) <= not((inputs(171)) and (inputs(241)));
    layer0_outputs(556) <= not(inputs(109));
    layer0_outputs(557) <= inputs(182);
    layer0_outputs(558) <= '0';
    layer0_outputs(559) <= not(inputs(126)) or (inputs(164));
    layer0_outputs(560) <= not(inputs(239));
    layer0_outputs(561) <= '1';
    layer0_outputs(562) <= not(inputs(170)) or (inputs(67));
    layer0_outputs(563) <= (inputs(57)) and not (inputs(26));
    layer0_outputs(564) <= not((inputs(104)) xor (inputs(178)));
    layer0_outputs(565) <= (inputs(205)) and not (inputs(160));
    layer0_outputs(566) <= (inputs(42)) and not (inputs(21));
    layer0_outputs(567) <= '0';
    layer0_outputs(568) <= not(inputs(97));
    layer0_outputs(569) <= (inputs(6)) or (inputs(71));
    layer0_outputs(570) <= not(inputs(68));
    layer0_outputs(571) <= (inputs(5)) and (inputs(59));
    layer0_outputs(572) <= inputs(145);
    layer0_outputs(573) <= inputs(120);
    layer0_outputs(574) <= inputs(80);
    layer0_outputs(575) <= not(inputs(114)) or (inputs(72));
    layer0_outputs(576) <= '1';
    layer0_outputs(577) <= not(inputs(23));
    layer0_outputs(578) <= (inputs(150)) and not (inputs(134));
    layer0_outputs(579) <= '0';
    layer0_outputs(580) <= '1';
    layer0_outputs(581) <= not(inputs(146));
    layer0_outputs(582) <= '0';
    layer0_outputs(583) <= (inputs(167)) and not (inputs(188));
    layer0_outputs(584) <= not(inputs(208)) or (inputs(254));
    layer0_outputs(585) <= not((inputs(216)) or (inputs(189)));
    layer0_outputs(586) <= (inputs(192)) or (inputs(227));
    layer0_outputs(587) <= (inputs(210)) and not (inputs(62));
    layer0_outputs(588) <= inputs(196);
    layer0_outputs(589) <= not(inputs(96)) or (inputs(18));
    layer0_outputs(590) <= inputs(252);
    layer0_outputs(591) <= not((inputs(197)) or (inputs(217)));
    layer0_outputs(592) <= not(inputs(156));
    layer0_outputs(593) <= '1';
    layer0_outputs(594) <= inputs(194);
    layer0_outputs(595) <= '0';
    layer0_outputs(596) <= (inputs(162)) and (inputs(139));
    layer0_outputs(597) <= not(inputs(19));
    layer0_outputs(598) <= inputs(5);
    layer0_outputs(599) <= not(inputs(164));
    layer0_outputs(600) <= '0';
    layer0_outputs(601) <= not(inputs(151)) or (inputs(18));
    layer0_outputs(602) <= not(inputs(213));
    layer0_outputs(603) <= not(inputs(21)) or (inputs(212));
    layer0_outputs(604) <= (inputs(158)) and not (inputs(182));
    layer0_outputs(605) <= not((inputs(253)) xor (inputs(22)));
    layer0_outputs(606) <= (inputs(129)) or (inputs(77));
    layer0_outputs(607) <= '1';
    layer0_outputs(608) <= (inputs(239)) and not (inputs(254));
    layer0_outputs(609) <= '1';
    layer0_outputs(610) <= (inputs(251)) or (inputs(137));
    layer0_outputs(611) <= not(inputs(199)) or (inputs(202));
    layer0_outputs(612) <= not(inputs(61));
    layer0_outputs(613) <= (inputs(74)) or (inputs(179));
    layer0_outputs(614) <= not(inputs(51)) or (inputs(105));
    layer0_outputs(615) <= (inputs(64)) and (inputs(77));
    layer0_outputs(616) <= '1';
    layer0_outputs(617) <= inputs(75);
    layer0_outputs(618) <= (inputs(89)) and not (inputs(127));
    layer0_outputs(619) <= (inputs(253)) and not (inputs(74));
    layer0_outputs(620) <= (inputs(209)) and (inputs(180));
    layer0_outputs(621) <= '0';
    layer0_outputs(622) <= not((inputs(156)) and (inputs(110)));
    layer0_outputs(623) <= '1';
    layer0_outputs(624) <= inputs(135);
    layer0_outputs(625) <= (inputs(144)) and not (inputs(199));
    layer0_outputs(626) <= inputs(178);
    layer0_outputs(627) <= not(inputs(86)) or (inputs(249));
    layer0_outputs(628) <= (inputs(157)) xor (inputs(175));
    layer0_outputs(629) <= inputs(238);
    layer0_outputs(630) <= not(inputs(82)) or (inputs(167));
    layer0_outputs(631) <= '1';
    layer0_outputs(632) <= (inputs(62)) and (inputs(251));
    layer0_outputs(633) <= inputs(117);
    layer0_outputs(634) <= not((inputs(219)) and (inputs(182)));
    layer0_outputs(635) <= (inputs(195)) or (inputs(143));
    layer0_outputs(636) <= (inputs(43)) and not (inputs(229));
    layer0_outputs(637) <= '1';
    layer0_outputs(638) <= (inputs(237)) and (inputs(15));
    layer0_outputs(639) <= not(inputs(41));
    layer0_outputs(640) <= (inputs(4)) and not (inputs(221));
    layer0_outputs(641) <= not(inputs(89)) or (inputs(212));
    layer0_outputs(642) <= not((inputs(86)) or (inputs(248)));
    layer0_outputs(643) <= (inputs(68)) xor (inputs(194));
    layer0_outputs(644) <= not(inputs(136)) or (inputs(146));
    layer0_outputs(645) <= not(inputs(216));
    layer0_outputs(646) <= inputs(196);
    layer0_outputs(647) <= inputs(129);
    layer0_outputs(648) <= (inputs(223)) or (inputs(33));
    layer0_outputs(649) <= not(inputs(176)) or (inputs(224));
    layer0_outputs(650) <= (inputs(194)) and (inputs(109));
    layer0_outputs(651) <= not(inputs(198)) or (inputs(58));
    layer0_outputs(652) <= not((inputs(154)) and (inputs(57)));
    layer0_outputs(653) <= not(inputs(20));
    layer0_outputs(654) <= not(inputs(43));
    layer0_outputs(655) <= not(inputs(105)) or (inputs(2));
    layer0_outputs(656) <= not((inputs(11)) and (inputs(50)));
    layer0_outputs(657) <= not(inputs(200)) or (inputs(210));
    layer0_outputs(658) <= (inputs(82)) and not (inputs(253));
    layer0_outputs(659) <= (inputs(203)) or (inputs(80));
    layer0_outputs(660) <= not(inputs(233));
    layer0_outputs(661) <= not(inputs(205));
    layer0_outputs(662) <= (inputs(64)) and not (inputs(65));
    layer0_outputs(663) <= not(inputs(162));
    layer0_outputs(664) <= (inputs(103)) or (inputs(46));
    layer0_outputs(665) <= (inputs(103)) or (inputs(212));
    layer0_outputs(666) <= (inputs(13)) xor (inputs(137));
    layer0_outputs(667) <= not(inputs(208));
    layer0_outputs(668) <= '0';
    layer0_outputs(669) <= '1';
    layer0_outputs(670) <= not((inputs(19)) or (inputs(253)));
    layer0_outputs(671) <= not((inputs(79)) and (inputs(136)));
    layer0_outputs(672) <= not((inputs(114)) xor (inputs(178)));
    layer0_outputs(673) <= inputs(80);
    layer0_outputs(674) <= inputs(87);
    layer0_outputs(675) <= (inputs(17)) and not (inputs(157));
    layer0_outputs(676) <= inputs(32);
    layer0_outputs(677) <= inputs(135);
    layer0_outputs(678) <= inputs(227);
    layer0_outputs(679) <= '1';
    layer0_outputs(680) <= inputs(105);
    layer0_outputs(681) <= '0';
    layer0_outputs(682) <= '1';
    layer0_outputs(683) <= '1';
    layer0_outputs(684) <= '0';
    layer0_outputs(685) <= (inputs(215)) and not (inputs(166));
    layer0_outputs(686) <= (inputs(233)) and not (inputs(23));
    layer0_outputs(687) <= '1';
    layer0_outputs(688) <= not((inputs(132)) or (inputs(243)));
    layer0_outputs(689) <= '1';
    layer0_outputs(690) <= '1';
    layer0_outputs(691) <= '0';
    layer0_outputs(692) <= not(inputs(160));
    layer0_outputs(693) <= '0';
    layer0_outputs(694) <= not((inputs(62)) or (inputs(232)));
    layer0_outputs(695) <= not(inputs(9));
    layer0_outputs(696) <= (inputs(98)) and not (inputs(10));
    layer0_outputs(697) <= '1';
    layer0_outputs(698) <= (inputs(181)) and (inputs(65));
    layer0_outputs(699) <= not(inputs(124));
    layer0_outputs(700) <= inputs(142);
    layer0_outputs(701) <= not((inputs(39)) and (inputs(82)));
    layer0_outputs(702) <= not((inputs(73)) xor (inputs(150)));
    layer0_outputs(703) <= '0';
    layer0_outputs(704) <= inputs(20);
    layer0_outputs(705) <= inputs(113);
    layer0_outputs(706) <= '1';
    layer0_outputs(707) <= not(inputs(127));
    layer0_outputs(708) <= '1';
    layer0_outputs(709) <= '1';
    layer0_outputs(710) <= (inputs(204)) or (inputs(188));
    layer0_outputs(711) <= not(inputs(143));
    layer0_outputs(712) <= '1';
    layer0_outputs(713) <= (inputs(76)) and not (inputs(194));
    layer0_outputs(714) <= inputs(129);
    layer0_outputs(715) <= (inputs(0)) and not (inputs(97));
    layer0_outputs(716) <= inputs(125);
    layer0_outputs(717) <= inputs(82);
    layer0_outputs(718) <= (inputs(31)) and (inputs(202));
    layer0_outputs(719) <= (inputs(204)) or (inputs(51));
    layer0_outputs(720) <= not((inputs(227)) xor (inputs(93)));
    layer0_outputs(721) <= inputs(65);
    layer0_outputs(722) <= not((inputs(155)) or (inputs(27)));
    layer0_outputs(723) <= not(inputs(97));
    layer0_outputs(724) <= (inputs(63)) or (inputs(37));
    layer0_outputs(725) <= not((inputs(86)) xor (inputs(206)));
    layer0_outputs(726) <= not(inputs(12)) or (inputs(166));
    layer0_outputs(727) <= not((inputs(177)) xor (inputs(251)));
    layer0_outputs(728) <= '1';
    layer0_outputs(729) <= inputs(66);
    layer0_outputs(730) <= '0';
    layer0_outputs(731) <= inputs(24);
    layer0_outputs(732) <= (inputs(235)) and not (inputs(237));
    layer0_outputs(733) <= not((inputs(47)) or (inputs(61)));
    layer0_outputs(734) <= not(inputs(100)) or (inputs(210));
    layer0_outputs(735) <= inputs(229);
    layer0_outputs(736) <= inputs(127);
    layer0_outputs(737) <= not(inputs(238));
    layer0_outputs(738) <= not((inputs(69)) or (inputs(246)));
    layer0_outputs(739) <= '0';
    layer0_outputs(740) <= (inputs(121)) and not (inputs(100));
    layer0_outputs(741) <= (inputs(135)) xor (inputs(235));
    layer0_outputs(742) <= inputs(230);
    layer0_outputs(743) <= not((inputs(102)) or (inputs(172)));
    layer0_outputs(744) <= (inputs(166)) and not (inputs(254));
    layer0_outputs(745) <= not((inputs(206)) or (inputs(43)));
    layer0_outputs(746) <= inputs(92);
    layer0_outputs(747) <= not((inputs(249)) or (inputs(237)));
    layer0_outputs(748) <= inputs(2);
    layer0_outputs(749) <= (inputs(77)) and not (inputs(237));
    layer0_outputs(750) <= not(inputs(120));
    layer0_outputs(751) <= not(inputs(76)) or (inputs(212));
    layer0_outputs(752) <= (inputs(254)) or (inputs(90));
    layer0_outputs(753) <= (inputs(21)) and (inputs(245));
    layer0_outputs(754) <= inputs(94);
    layer0_outputs(755) <= (inputs(224)) and (inputs(252));
    layer0_outputs(756) <= '1';
    layer0_outputs(757) <= '0';
    layer0_outputs(758) <= '0';
    layer0_outputs(759) <= (inputs(155)) and not (inputs(15));
    layer0_outputs(760) <= not((inputs(141)) and (inputs(9)));
    layer0_outputs(761) <= (inputs(116)) and (inputs(67));
    layer0_outputs(762) <= '1';
    layer0_outputs(763) <= not(inputs(166)) or (inputs(56));
    layer0_outputs(764) <= '0';
    layer0_outputs(765) <= (inputs(172)) and not (inputs(72));
    layer0_outputs(766) <= not((inputs(53)) or (inputs(142)));
    layer0_outputs(767) <= not((inputs(140)) and (inputs(192)));
    layer0_outputs(768) <= inputs(70);
    layer0_outputs(769) <= not((inputs(245)) xor (inputs(231)));
    layer0_outputs(770) <= not((inputs(210)) xor (inputs(101)));
    layer0_outputs(771) <= inputs(78);
    layer0_outputs(772) <= (inputs(70)) and not (inputs(79));
    layer0_outputs(773) <= (inputs(153)) and (inputs(234));
    layer0_outputs(774) <= (inputs(103)) and not (inputs(127));
    layer0_outputs(775) <= '0';
    layer0_outputs(776) <= not((inputs(129)) or (inputs(127)));
    layer0_outputs(777) <= not(inputs(7)) or (inputs(34));
    layer0_outputs(778) <= inputs(69);
    layer0_outputs(779) <= '1';
    layer0_outputs(780) <= (inputs(99)) and (inputs(126));
    layer0_outputs(781) <= not(inputs(146)) or (inputs(206));
    layer0_outputs(782) <= (inputs(236)) and not (inputs(113));
    layer0_outputs(783) <= '1';
    layer0_outputs(784) <= (inputs(131)) and not (inputs(14));
    layer0_outputs(785) <= not(inputs(207));
    layer0_outputs(786) <= not(inputs(161));
    layer0_outputs(787) <= inputs(180);
    layer0_outputs(788) <= (inputs(0)) or (inputs(252));
    layer0_outputs(789) <= not((inputs(183)) or (inputs(120)));
    layer0_outputs(790) <= '1';
    layer0_outputs(791) <= not((inputs(167)) xor (inputs(48)));
    layer0_outputs(792) <= not(inputs(55));
    layer0_outputs(793) <= not((inputs(208)) and (inputs(250)));
    layer0_outputs(794) <= inputs(134);
    layer0_outputs(795) <= not((inputs(30)) or (inputs(168)));
    layer0_outputs(796) <= '1';
    layer0_outputs(797) <= '1';
    layer0_outputs(798) <= not(inputs(63));
    layer0_outputs(799) <= '0';
    layer0_outputs(800) <= (inputs(9)) or (inputs(24));
    layer0_outputs(801) <= (inputs(168)) and not (inputs(9));
    layer0_outputs(802) <= inputs(164);
    layer0_outputs(803) <= inputs(3);
    layer0_outputs(804) <= (inputs(245)) and not (inputs(62));
    layer0_outputs(805) <= not(inputs(201)) or (inputs(13));
    layer0_outputs(806) <= '1';
    layer0_outputs(807) <= not((inputs(177)) xor (inputs(196)));
    layer0_outputs(808) <= '0';
    layer0_outputs(809) <= inputs(125);
    layer0_outputs(810) <= '0';
    layer0_outputs(811) <= '0';
    layer0_outputs(812) <= not(inputs(230));
    layer0_outputs(813) <= not(inputs(15));
    layer0_outputs(814) <= not((inputs(213)) or (inputs(225)));
    layer0_outputs(815) <= not(inputs(54)) or (inputs(56));
    layer0_outputs(816) <= not(inputs(176));
    layer0_outputs(817) <= '0';
    layer0_outputs(818) <= (inputs(163)) xor (inputs(84));
    layer0_outputs(819) <= (inputs(41)) and (inputs(22));
    layer0_outputs(820) <= '1';
    layer0_outputs(821) <= (inputs(250)) and not (inputs(173));
    layer0_outputs(822) <= inputs(228);
    layer0_outputs(823) <= (inputs(235)) and not (inputs(126));
    layer0_outputs(824) <= not((inputs(121)) or (inputs(151)));
    layer0_outputs(825) <= '1';
    layer0_outputs(826) <= (inputs(5)) and (inputs(123));
    layer0_outputs(827) <= not((inputs(171)) xor (inputs(221)));
    layer0_outputs(828) <= '1';
    layer0_outputs(829) <= not(inputs(38));
    layer0_outputs(830) <= '1';
    layer0_outputs(831) <= (inputs(228)) and not (inputs(43));
    layer0_outputs(832) <= not((inputs(84)) and (inputs(121)));
    layer0_outputs(833) <= inputs(151);
    layer0_outputs(834) <= '1';
    layer0_outputs(835) <= '0';
    layer0_outputs(836) <= not((inputs(176)) and (inputs(18)));
    layer0_outputs(837) <= not((inputs(67)) and (inputs(106)));
    layer0_outputs(838) <= not((inputs(78)) or (inputs(30)));
    layer0_outputs(839) <= not(inputs(172)) or (inputs(79));
    layer0_outputs(840) <= (inputs(168)) and not (inputs(92));
    layer0_outputs(841) <= (inputs(138)) and not (inputs(69));
    layer0_outputs(842) <= (inputs(112)) and not (inputs(11));
    layer0_outputs(843) <= (inputs(220)) and not (inputs(92));
    layer0_outputs(844) <= not(inputs(27)) or (inputs(25));
    layer0_outputs(845) <= (inputs(157)) and (inputs(9));
    layer0_outputs(846) <= '1';
    layer0_outputs(847) <= (inputs(93)) and (inputs(48));
    layer0_outputs(848) <= not(inputs(75));
    layer0_outputs(849) <= not((inputs(222)) or (inputs(3)));
    layer0_outputs(850) <= not(inputs(213)) or (inputs(109));
    layer0_outputs(851) <= (inputs(128)) and not (inputs(254));
    layer0_outputs(852) <= not((inputs(152)) and (inputs(62)));
    layer0_outputs(853) <= '0';
    layer0_outputs(854) <= not(inputs(221)) or (inputs(54));
    layer0_outputs(855) <= '1';
    layer0_outputs(856) <= not((inputs(249)) and (inputs(80)));
    layer0_outputs(857) <= not((inputs(82)) or (inputs(133)));
    layer0_outputs(858) <= '1';
    layer0_outputs(859) <= '0';
    layer0_outputs(860) <= '1';
    layer0_outputs(861) <= not((inputs(236)) or (inputs(209)));
    layer0_outputs(862) <= (inputs(86)) and not (inputs(100));
    layer0_outputs(863) <= not(inputs(171)) or (inputs(166));
    layer0_outputs(864) <= (inputs(153)) and not (inputs(172));
    layer0_outputs(865) <= inputs(161);
    layer0_outputs(866) <= not(inputs(28));
    layer0_outputs(867) <= (inputs(20)) and not (inputs(160));
    layer0_outputs(868) <= '1';
    layer0_outputs(869) <= not(inputs(230));
    layer0_outputs(870) <= (inputs(180)) and (inputs(86));
    layer0_outputs(871) <= not((inputs(191)) or (inputs(180)));
    layer0_outputs(872) <= inputs(228);
    layer0_outputs(873) <= '0';
    layer0_outputs(874) <= not((inputs(168)) or (inputs(201)));
    layer0_outputs(875) <= inputs(203);
    layer0_outputs(876) <= not((inputs(204)) or (inputs(44)));
    layer0_outputs(877) <= not(inputs(137)) or (inputs(123));
    layer0_outputs(878) <= (inputs(130)) or (inputs(211));
    layer0_outputs(879) <= inputs(101);
    layer0_outputs(880) <= not(inputs(96)) or (inputs(214));
    layer0_outputs(881) <= not(inputs(228));
    layer0_outputs(882) <= '0';
    layer0_outputs(883) <= (inputs(137)) and (inputs(73));
    layer0_outputs(884) <= not((inputs(30)) or (inputs(20)));
    layer0_outputs(885) <= not(inputs(102)) or (inputs(183));
    layer0_outputs(886) <= not(inputs(52));
    layer0_outputs(887) <= not(inputs(30));
    layer0_outputs(888) <= inputs(46);
    layer0_outputs(889) <= (inputs(7)) xor (inputs(177));
    layer0_outputs(890) <= '0';
    layer0_outputs(891) <= '1';
    layer0_outputs(892) <= not(inputs(64));
    layer0_outputs(893) <= not(inputs(65)) or (inputs(155));
    layer0_outputs(894) <= not((inputs(142)) or (inputs(142)));
    layer0_outputs(895) <= not(inputs(242)) or (inputs(26));
    layer0_outputs(896) <= (inputs(251)) and not (inputs(181));
    layer0_outputs(897) <= inputs(98);
    layer0_outputs(898) <= inputs(227);
    layer0_outputs(899) <= inputs(104);
    layer0_outputs(900) <= (inputs(116)) and not (inputs(179));
    layer0_outputs(901) <= (inputs(158)) and (inputs(227));
    layer0_outputs(902) <= '0';
    layer0_outputs(903) <= inputs(37);
    layer0_outputs(904) <= not(inputs(224)) or (inputs(58));
    layer0_outputs(905) <= '0';
    layer0_outputs(906) <= not(inputs(218)) or (inputs(107));
    layer0_outputs(907) <= not((inputs(84)) and (inputs(81)));
    layer0_outputs(908) <= (inputs(185)) and (inputs(141));
    layer0_outputs(909) <= inputs(147);
    layer0_outputs(910) <= inputs(119);
    layer0_outputs(911) <= not(inputs(36)) or (inputs(110));
    layer0_outputs(912) <= '1';
    layer0_outputs(913) <= '0';
    layer0_outputs(914) <= (inputs(119)) or (inputs(83));
    layer0_outputs(915) <= (inputs(53)) and not (inputs(190));
    layer0_outputs(916) <= '1';
    layer0_outputs(917) <= not(inputs(23)) or (inputs(39));
    layer0_outputs(918) <= inputs(82);
    layer0_outputs(919) <= inputs(232);
    layer0_outputs(920) <= '1';
    layer0_outputs(921) <= not(inputs(254)) or (inputs(27));
    layer0_outputs(922) <= inputs(168);
    layer0_outputs(923) <= (inputs(37)) and not (inputs(160));
    layer0_outputs(924) <= not(inputs(226)) or (inputs(145));
    layer0_outputs(925) <= inputs(251);
    layer0_outputs(926) <= not((inputs(103)) or (inputs(177)));
    layer0_outputs(927) <= inputs(47);
    layer0_outputs(928) <= '1';
    layer0_outputs(929) <= not((inputs(65)) or (inputs(83)));
    layer0_outputs(930) <= not(inputs(77)) or (inputs(224));
    layer0_outputs(931) <= inputs(144);
    layer0_outputs(932) <= (inputs(223)) or (inputs(182));
    layer0_outputs(933) <= not((inputs(240)) and (inputs(104)));
    layer0_outputs(934) <= '1';
    layer0_outputs(935) <= (inputs(8)) or (inputs(69));
    layer0_outputs(936) <= inputs(188);
    layer0_outputs(937) <= inputs(226);
    layer0_outputs(938) <= not(inputs(24));
    layer0_outputs(939) <= (inputs(119)) and (inputs(140));
    layer0_outputs(940) <= not(inputs(91));
    layer0_outputs(941) <= inputs(84);
    layer0_outputs(942) <= '0';
    layer0_outputs(943) <= (inputs(67)) and (inputs(239));
    layer0_outputs(944) <= not(inputs(80)) or (inputs(173));
    layer0_outputs(945) <= '1';
    layer0_outputs(946) <= not(inputs(125)) or (inputs(116));
    layer0_outputs(947) <= not(inputs(125)) or (inputs(49));
    layer0_outputs(948) <= not((inputs(36)) and (inputs(192)));
    layer0_outputs(949) <= not(inputs(5));
    layer0_outputs(950) <= '0';
    layer0_outputs(951) <= (inputs(84)) and not (inputs(230));
    layer0_outputs(952) <= '0';
    layer0_outputs(953) <= not(inputs(181)) or (inputs(225));
    layer0_outputs(954) <= '0';
    layer0_outputs(955) <= '1';
    layer0_outputs(956) <= not(inputs(19));
    layer0_outputs(957) <= not((inputs(75)) and (inputs(101)));
    layer0_outputs(958) <= (inputs(204)) and not (inputs(163));
    layer0_outputs(959) <= not(inputs(50)) or (inputs(212));
    layer0_outputs(960) <= not(inputs(118)) or (inputs(78));
    layer0_outputs(961) <= inputs(132);
    layer0_outputs(962) <= inputs(214);
    layer0_outputs(963) <= (inputs(28)) or (inputs(125));
    layer0_outputs(964) <= (inputs(60)) or (inputs(75));
    layer0_outputs(965) <= '0';
    layer0_outputs(966) <= (inputs(77)) or (inputs(32));
    layer0_outputs(967) <= not(inputs(25));
    layer0_outputs(968) <= not(inputs(129)) or (inputs(0));
    layer0_outputs(969) <= inputs(102);
    layer0_outputs(970) <= inputs(36);
    layer0_outputs(971) <= not(inputs(145)) or (inputs(121));
    layer0_outputs(972) <= not(inputs(165));
    layer0_outputs(973) <= (inputs(174)) and not (inputs(15));
    layer0_outputs(974) <= '0';
    layer0_outputs(975) <= '1';
    layer0_outputs(976) <= '1';
    layer0_outputs(977) <= not(inputs(110));
    layer0_outputs(978) <= not(inputs(242));
    layer0_outputs(979) <= inputs(99);
    layer0_outputs(980) <= not(inputs(117));
    layer0_outputs(981) <= not((inputs(82)) or (inputs(144)));
    layer0_outputs(982) <= '0';
    layer0_outputs(983) <= not(inputs(133));
    layer0_outputs(984) <= '0';
    layer0_outputs(985) <= (inputs(83)) or (inputs(204));
    layer0_outputs(986) <= not((inputs(120)) and (inputs(25)));
    layer0_outputs(987) <= (inputs(234)) or (inputs(171));
    layer0_outputs(988) <= '1';
    layer0_outputs(989) <= not(inputs(255));
    layer0_outputs(990) <= not((inputs(21)) or (inputs(234)));
    layer0_outputs(991) <= (inputs(93)) or (inputs(146));
    layer0_outputs(992) <= '1';
    layer0_outputs(993) <= '1';
    layer0_outputs(994) <= inputs(47);
    layer0_outputs(995) <= '0';
    layer0_outputs(996) <= inputs(23);
    layer0_outputs(997) <= inputs(141);
    layer0_outputs(998) <= (inputs(135)) or (inputs(63));
    layer0_outputs(999) <= not(inputs(26));
    layer0_outputs(1000) <= '1';
    layer0_outputs(1001) <= (inputs(226)) or (inputs(44));
    layer0_outputs(1002) <= not((inputs(254)) and (inputs(1)));
    layer0_outputs(1003) <= (inputs(45)) and (inputs(41));
    layer0_outputs(1004) <= not(inputs(186));
    layer0_outputs(1005) <= '1';
    layer0_outputs(1006) <= '0';
    layer0_outputs(1007) <= not(inputs(230));
    layer0_outputs(1008) <= (inputs(10)) and not (inputs(146));
    layer0_outputs(1009) <= '1';
    layer0_outputs(1010) <= inputs(145);
    layer0_outputs(1011) <= '1';
    layer0_outputs(1012) <= '0';
    layer0_outputs(1013) <= inputs(27);
    layer0_outputs(1014) <= (inputs(32)) and (inputs(186));
    layer0_outputs(1015) <= '0';
    layer0_outputs(1016) <= '1';
    layer0_outputs(1017) <= inputs(119);
    layer0_outputs(1018) <= not(inputs(66));
    layer0_outputs(1019) <= (inputs(121)) and (inputs(101));
    layer0_outputs(1020) <= '1';
    layer0_outputs(1021) <= inputs(61);
    layer0_outputs(1022) <= not(inputs(74));
    layer0_outputs(1023) <= (inputs(81)) and not (inputs(60));
    layer0_outputs(1024) <= not((inputs(228)) and (inputs(39)));
    layer0_outputs(1025) <= (inputs(146)) and not (inputs(1));
    layer0_outputs(1026) <= (inputs(72)) or (inputs(236));
    layer0_outputs(1027) <= not((inputs(25)) or (inputs(57)));
    layer0_outputs(1028) <= '0';
    layer0_outputs(1029) <= inputs(200);
    layer0_outputs(1030) <= not(inputs(167));
    layer0_outputs(1031) <= not(inputs(182)) or (inputs(138));
    layer0_outputs(1032) <= not(inputs(215)) or (inputs(183));
    layer0_outputs(1033) <= '1';
    layer0_outputs(1034) <= '1';
    layer0_outputs(1035) <= (inputs(134)) and not (inputs(191));
    layer0_outputs(1036) <= inputs(31);
    layer0_outputs(1037) <= not((inputs(199)) and (inputs(57)));
    layer0_outputs(1038) <= (inputs(74)) xor (inputs(80));
    layer0_outputs(1039) <= not(inputs(13)) or (inputs(70));
    layer0_outputs(1040) <= '1';
    layer0_outputs(1041) <= (inputs(66)) and (inputs(113));
    layer0_outputs(1042) <= inputs(179);
    layer0_outputs(1043) <= not((inputs(167)) and (inputs(171)));
    layer0_outputs(1044) <= not((inputs(64)) or (inputs(64)));
    layer0_outputs(1045) <= inputs(100);
    layer0_outputs(1046) <= '1';
    layer0_outputs(1047) <= not(inputs(245));
    layer0_outputs(1048) <= '1';
    layer0_outputs(1049) <= '1';
    layer0_outputs(1050) <= '0';
    layer0_outputs(1051) <= (inputs(106)) and (inputs(78));
    layer0_outputs(1052) <= not(inputs(83));
    layer0_outputs(1053) <= not(inputs(143));
    layer0_outputs(1054) <= not(inputs(249));
    layer0_outputs(1055) <= inputs(227);
    layer0_outputs(1056) <= inputs(197);
    layer0_outputs(1057) <= (inputs(137)) and not (inputs(214));
    layer0_outputs(1058) <= not(inputs(11));
    layer0_outputs(1059) <= (inputs(10)) and not (inputs(54));
    layer0_outputs(1060) <= '0';
    layer0_outputs(1061) <= not(inputs(52));
    layer0_outputs(1062) <= inputs(129);
    layer0_outputs(1063) <= inputs(175);
    layer0_outputs(1064) <= inputs(22);
    layer0_outputs(1065) <= not(inputs(34));
    layer0_outputs(1066) <= not((inputs(131)) or (inputs(34)));
    layer0_outputs(1067) <= not(inputs(133)) or (inputs(7));
    layer0_outputs(1068) <= (inputs(30)) or (inputs(186));
    layer0_outputs(1069) <= (inputs(106)) and not (inputs(80));
    layer0_outputs(1070) <= inputs(109);
    layer0_outputs(1071) <= inputs(253);
    layer0_outputs(1072) <= (inputs(19)) or (inputs(237));
    layer0_outputs(1073) <= inputs(159);
    layer0_outputs(1074) <= not(inputs(107)) or (inputs(128));
    layer0_outputs(1075) <= inputs(18);
    layer0_outputs(1076) <= not(inputs(36)) or (inputs(154));
    layer0_outputs(1077) <= '0';
    layer0_outputs(1078) <= (inputs(247)) and not (inputs(59));
    layer0_outputs(1079) <= inputs(248);
    layer0_outputs(1080) <= '1';
    layer0_outputs(1081) <= not(inputs(105));
    layer0_outputs(1082) <= not(inputs(246));
    layer0_outputs(1083) <= inputs(83);
    layer0_outputs(1084) <= '0';
    layer0_outputs(1085) <= inputs(93);
    layer0_outputs(1086) <= '0';
    layer0_outputs(1087) <= (inputs(115)) and not (inputs(223));
    layer0_outputs(1088) <= not((inputs(117)) xor (inputs(35)));
    layer0_outputs(1089) <= not(inputs(207));
    layer0_outputs(1090) <= '0';
    layer0_outputs(1091) <= (inputs(136)) and not (inputs(245));
    layer0_outputs(1092) <= (inputs(148)) and (inputs(95));
    layer0_outputs(1093) <= (inputs(78)) or (inputs(16));
    layer0_outputs(1094) <= inputs(136);
    layer0_outputs(1095) <= inputs(4);
    layer0_outputs(1096) <= not((inputs(141)) or (inputs(158)));
    layer0_outputs(1097) <= (inputs(216)) or (inputs(232));
    layer0_outputs(1098) <= '0';
    layer0_outputs(1099) <= not((inputs(157)) or (inputs(84)));
    layer0_outputs(1100) <= (inputs(63)) xor (inputs(50));
    layer0_outputs(1101) <= not(inputs(8));
    layer0_outputs(1102) <= '1';
    layer0_outputs(1103) <= '0';
    layer0_outputs(1104) <= '0';
    layer0_outputs(1105) <= (inputs(55)) and not (inputs(90));
    layer0_outputs(1106) <= '1';
    layer0_outputs(1107) <= '1';
    layer0_outputs(1108) <= '0';
    layer0_outputs(1109) <= not(inputs(190)) or (inputs(192));
    layer0_outputs(1110) <= not((inputs(184)) or (inputs(196)));
    layer0_outputs(1111) <= '0';
    layer0_outputs(1112) <= not(inputs(122));
    layer0_outputs(1113) <= not(inputs(149)) or (inputs(141));
    layer0_outputs(1114) <= not(inputs(31)) or (inputs(244));
    layer0_outputs(1115) <= not(inputs(224));
    layer0_outputs(1116) <= not((inputs(67)) or (inputs(225)));
    layer0_outputs(1117) <= not((inputs(203)) or (inputs(96)));
    layer0_outputs(1118) <= (inputs(54)) and not (inputs(87));
    layer0_outputs(1119) <= not(inputs(25));
    layer0_outputs(1120) <= (inputs(140)) or (inputs(157));
    layer0_outputs(1121) <= (inputs(147)) and not (inputs(119));
    layer0_outputs(1122) <= '0';
    layer0_outputs(1123) <= inputs(107);
    layer0_outputs(1124) <= inputs(20);
    layer0_outputs(1125) <= '0';
    layer0_outputs(1126) <= not(inputs(178));
    layer0_outputs(1127) <= not(inputs(100));
    layer0_outputs(1128) <= not((inputs(36)) xor (inputs(19)));
    layer0_outputs(1129) <= (inputs(146)) or (inputs(52));
    layer0_outputs(1130) <= (inputs(225)) or (inputs(241));
    layer0_outputs(1131) <= inputs(130);
    layer0_outputs(1132) <= (inputs(97)) and not (inputs(161));
    layer0_outputs(1133) <= (inputs(159)) or (inputs(103));
    layer0_outputs(1134) <= '1';
    layer0_outputs(1135) <= (inputs(138)) or (inputs(175));
    layer0_outputs(1136) <= '1';
    layer0_outputs(1137) <= not((inputs(244)) or (inputs(246)));
    layer0_outputs(1138) <= inputs(67);
    layer0_outputs(1139) <= '0';
    layer0_outputs(1140) <= '1';
    layer0_outputs(1141) <= not(inputs(20));
    layer0_outputs(1142) <= '0';
    layer0_outputs(1143) <= (inputs(158)) and not (inputs(210));
    layer0_outputs(1144) <= not((inputs(53)) xor (inputs(160)));
    layer0_outputs(1145) <= not(inputs(36)) or (inputs(132));
    layer0_outputs(1146) <= not((inputs(116)) and (inputs(174)));
    layer0_outputs(1147) <= '1';
    layer0_outputs(1148) <= (inputs(118)) and not (inputs(207));
    layer0_outputs(1149) <= not(inputs(114));
    layer0_outputs(1150) <= '1';
    layer0_outputs(1151) <= not(inputs(96));
    layer0_outputs(1152) <= inputs(212);
    layer0_outputs(1153) <= '1';
    layer0_outputs(1154) <= inputs(9);
    layer0_outputs(1155) <= not(inputs(201)) or (inputs(152));
    layer0_outputs(1156) <= not(inputs(138));
    layer0_outputs(1157) <= '0';
    layer0_outputs(1158) <= inputs(76);
    layer0_outputs(1159) <= (inputs(23)) and not (inputs(159));
    layer0_outputs(1160) <= (inputs(138)) and not (inputs(76));
    layer0_outputs(1161) <= not(inputs(255));
    layer0_outputs(1162) <= inputs(63);
    layer0_outputs(1163) <= not(inputs(155)) or (inputs(49));
    layer0_outputs(1164) <= inputs(239);
    layer0_outputs(1165) <= (inputs(121)) xor (inputs(176));
    layer0_outputs(1166) <= inputs(109);
    layer0_outputs(1167) <= not(inputs(118)) or (inputs(99));
    layer0_outputs(1168) <= not((inputs(120)) and (inputs(2)));
    layer0_outputs(1169) <= not((inputs(137)) and (inputs(41)));
    layer0_outputs(1170) <= not(inputs(251)) or (inputs(249));
    layer0_outputs(1171) <= (inputs(16)) and not (inputs(233));
    layer0_outputs(1172) <= not((inputs(170)) and (inputs(143)));
    layer0_outputs(1173) <= '0';
    layer0_outputs(1174) <= not(inputs(153)) or (inputs(18));
    layer0_outputs(1175) <= '1';
    layer0_outputs(1176) <= inputs(233);
    layer0_outputs(1177) <= not(inputs(120)) or (inputs(163));
    layer0_outputs(1178) <= inputs(135);
    layer0_outputs(1179) <= inputs(163);
    layer0_outputs(1180) <= not(inputs(92)) or (inputs(191));
    layer0_outputs(1181) <= inputs(119);
    layer0_outputs(1182) <= (inputs(241)) and (inputs(21));
    layer0_outputs(1183) <= inputs(56);
    layer0_outputs(1184) <= not((inputs(232)) and (inputs(23)));
    layer0_outputs(1185) <= not(inputs(178)) or (inputs(199));
    layer0_outputs(1186) <= not(inputs(100)) or (inputs(39));
    layer0_outputs(1187) <= (inputs(140)) xor (inputs(128));
    layer0_outputs(1188) <= '1';
    layer0_outputs(1189) <= not(inputs(90));
    layer0_outputs(1190) <= not((inputs(75)) or (inputs(183)));
    layer0_outputs(1191) <= not(inputs(70));
    layer0_outputs(1192) <= (inputs(124)) or (inputs(155));
    layer0_outputs(1193) <= '1';
    layer0_outputs(1194) <= not(inputs(118));
    layer0_outputs(1195) <= inputs(243);
    layer0_outputs(1196) <= not((inputs(223)) or (inputs(170)));
    layer0_outputs(1197) <= (inputs(25)) and not (inputs(57));
    layer0_outputs(1198) <= '1';
    layer0_outputs(1199) <= '1';
    layer0_outputs(1200) <= not(inputs(155)) or (inputs(156));
    layer0_outputs(1201) <= '1';
    layer0_outputs(1202) <= not(inputs(147));
    layer0_outputs(1203) <= not((inputs(223)) or (inputs(195)));
    layer0_outputs(1204) <= (inputs(88)) and not (inputs(94));
    layer0_outputs(1205) <= '1';
    layer0_outputs(1206) <= '0';
    layer0_outputs(1207) <= not(inputs(212)) or (inputs(33));
    layer0_outputs(1208) <= (inputs(164)) and (inputs(42));
    layer0_outputs(1209) <= inputs(86);
    layer0_outputs(1210) <= not(inputs(209));
    layer0_outputs(1211) <= '0';
    layer0_outputs(1212) <= inputs(129);
    layer0_outputs(1213) <= not(inputs(24));
    layer0_outputs(1214) <= '0';
    layer0_outputs(1215) <= inputs(254);
    layer0_outputs(1216) <= (inputs(100)) or (inputs(219));
    layer0_outputs(1217) <= '0';
    layer0_outputs(1218) <= not(inputs(16));
    layer0_outputs(1219) <= (inputs(220)) or (inputs(108));
    layer0_outputs(1220) <= inputs(76);
    layer0_outputs(1221) <= not((inputs(12)) and (inputs(57)));
    layer0_outputs(1222) <= inputs(49);
    layer0_outputs(1223) <= (inputs(66)) or (inputs(115));
    layer0_outputs(1224) <= not((inputs(199)) or (inputs(223)));
    layer0_outputs(1225) <= not((inputs(26)) or (inputs(16)));
    layer0_outputs(1226) <= not(inputs(178));
    layer0_outputs(1227) <= not(inputs(246));
    layer0_outputs(1228) <= not((inputs(180)) xor (inputs(198)));
    layer0_outputs(1229) <= not(inputs(130));
    layer0_outputs(1230) <= inputs(183);
    layer0_outputs(1231) <= (inputs(10)) or (inputs(36));
    layer0_outputs(1232) <= '1';
    layer0_outputs(1233) <= (inputs(249)) xor (inputs(35));
    layer0_outputs(1234) <= (inputs(254)) xor (inputs(189));
    layer0_outputs(1235) <= inputs(1);
    layer0_outputs(1236) <= (inputs(36)) and not (inputs(25));
    layer0_outputs(1237) <= (inputs(145)) and (inputs(8));
    layer0_outputs(1238) <= not(inputs(28)) or (inputs(190));
    layer0_outputs(1239) <= (inputs(88)) and not (inputs(112));
    layer0_outputs(1240) <= (inputs(255)) or (inputs(121));
    layer0_outputs(1241) <= '1';
    layer0_outputs(1242) <= inputs(218);
    layer0_outputs(1243) <= '1';
    layer0_outputs(1244) <= (inputs(111)) and not (inputs(3));
    layer0_outputs(1245) <= '1';
    layer0_outputs(1246) <= inputs(211);
    layer0_outputs(1247) <= inputs(208);
    layer0_outputs(1248) <= '1';
    layer0_outputs(1249) <= (inputs(95)) or (inputs(230));
    layer0_outputs(1250) <= inputs(174);
    layer0_outputs(1251) <= '0';
    layer0_outputs(1252) <= inputs(68);
    layer0_outputs(1253) <= not(inputs(59)) or (inputs(236));
    layer0_outputs(1254) <= not((inputs(215)) and (inputs(208)));
    layer0_outputs(1255) <= not((inputs(190)) or (inputs(53)));
    layer0_outputs(1256) <= '0';
    layer0_outputs(1257) <= not((inputs(157)) and (inputs(31)));
    layer0_outputs(1258) <= not((inputs(38)) or (inputs(14)));
    layer0_outputs(1259) <= not(inputs(127)) or (inputs(31));
    layer0_outputs(1260) <= (inputs(186)) or (inputs(85));
    layer0_outputs(1261) <= (inputs(8)) xor (inputs(216));
    layer0_outputs(1262) <= inputs(125);
    layer0_outputs(1263) <= (inputs(140)) or (inputs(31));
    layer0_outputs(1264) <= not(inputs(228));
    layer0_outputs(1265) <= not((inputs(236)) or (inputs(22)));
    layer0_outputs(1266) <= not(inputs(116));
    layer0_outputs(1267) <= inputs(245);
    layer0_outputs(1268) <= '0';
    layer0_outputs(1269) <= (inputs(201)) and (inputs(210));
    layer0_outputs(1270) <= (inputs(147)) and not (inputs(72));
    layer0_outputs(1271) <= not(inputs(221)) or (inputs(159));
    layer0_outputs(1272) <= (inputs(193)) and not (inputs(218));
    layer0_outputs(1273) <= not((inputs(119)) and (inputs(209)));
    layer0_outputs(1274) <= inputs(113);
    layer0_outputs(1275) <= (inputs(179)) and not (inputs(174));
    layer0_outputs(1276) <= '1';
    layer0_outputs(1277) <= not(inputs(61));
    layer0_outputs(1278) <= inputs(59);
    layer0_outputs(1279) <= inputs(197);
    layer0_outputs(1280) <= not((inputs(172)) or (inputs(205)));
    layer0_outputs(1281) <= '1';
    layer0_outputs(1282) <= not((inputs(229)) and (inputs(242)));
    layer0_outputs(1283) <= '1';
    layer0_outputs(1284) <= not(inputs(24)) or (inputs(208));
    layer0_outputs(1285) <= not(inputs(78));
    layer0_outputs(1286) <= inputs(123);
    layer0_outputs(1287) <= inputs(106);
    layer0_outputs(1288) <= not((inputs(190)) or (inputs(157)));
    layer0_outputs(1289) <= not(inputs(157));
    layer0_outputs(1290) <= (inputs(161)) and not (inputs(61));
    layer0_outputs(1291) <= not((inputs(44)) and (inputs(54)));
    layer0_outputs(1292) <= (inputs(224)) or (inputs(209));
    layer0_outputs(1293) <= not(inputs(224));
    layer0_outputs(1294) <= (inputs(131)) and (inputs(108));
    layer0_outputs(1295) <= '0';
    layer0_outputs(1296) <= not(inputs(109)) or (inputs(105));
    layer0_outputs(1297) <= not((inputs(34)) or (inputs(146)));
    layer0_outputs(1298) <= not(inputs(71)) or (inputs(152));
    layer0_outputs(1299) <= (inputs(18)) and not (inputs(129));
    layer0_outputs(1300) <= '1';
    layer0_outputs(1301) <= (inputs(212)) or (inputs(232));
    layer0_outputs(1302) <= '0';
    layer0_outputs(1303) <= (inputs(112)) and not (inputs(78));
    layer0_outputs(1304) <= not(inputs(125)) or (inputs(187));
    layer0_outputs(1305) <= '1';
    layer0_outputs(1306) <= (inputs(86)) and not (inputs(48));
    layer0_outputs(1307) <= '1';
    layer0_outputs(1308) <= (inputs(172)) and (inputs(112));
    layer0_outputs(1309) <= not(inputs(16));
    layer0_outputs(1310) <= (inputs(98)) and not (inputs(153));
    layer0_outputs(1311) <= inputs(84);
    layer0_outputs(1312) <= not(inputs(216));
    layer0_outputs(1313) <= inputs(200);
    layer0_outputs(1314) <= '0';
    layer0_outputs(1315) <= not(inputs(22));
    layer0_outputs(1316) <= (inputs(207)) and (inputs(47));
    layer0_outputs(1317) <= '1';
    layer0_outputs(1318) <= '0';
    layer0_outputs(1319) <= '0';
    layer0_outputs(1320) <= (inputs(114)) and not (inputs(91));
    layer0_outputs(1321) <= inputs(45);
    layer0_outputs(1322) <= (inputs(140)) or (inputs(66));
    layer0_outputs(1323) <= not(inputs(153));
    layer0_outputs(1324) <= not(inputs(129));
    layer0_outputs(1325) <= not(inputs(223));
    layer0_outputs(1326) <= (inputs(182)) and (inputs(42));
    layer0_outputs(1327) <= (inputs(17)) or (inputs(43));
    layer0_outputs(1328) <= not(inputs(26)) or (inputs(4));
    layer0_outputs(1329) <= (inputs(132)) and not (inputs(167));
    layer0_outputs(1330) <= '0';
    layer0_outputs(1331) <= not(inputs(157));
    layer0_outputs(1332) <= not(inputs(27));
    layer0_outputs(1333) <= (inputs(71)) and (inputs(67));
    layer0_outputs(1334) <= '0';
    layer0_outputs(1335) <= (inputs(137)) and not (inputs(80));
    layer0_outputs(1336) <= (inputs(103)) and not (inputs(14));
    layer0_outputs(1337) <= not(inputs(176)) or (inputs(115));
    layer0_outputs(1338) <= not(inputs(112));
    layer0_outputs(1339) <= (inputs(206)) or (inputs(64));
    layer0_outputs(1340) <= not(inputs(88)) or (inputs(130));
    layer0_outputs(1341) <= not(inputs(193)) or (inputs(154));
    layer0_outputs(1342) <= '1';
    layer0_outputs(1343) <= not((inputs(151)) and (inputs(202)));
    layer0_outputs(1344) <= (inputs(192)) or (inputs(94));
    layer0_outputs(1345) <= (inputs(232)) xor (inputs(3));
    layer0_outputs(1346) <= inputs(229);
    layer0_outputs(1347) <= not(inputs(243));
    layer0_outputs(1348) <= not(inputs(27));
    layer0_outputs(1349) <= (inputs(28)) and not (inputs(225));
    layer0_outputs(1350) <= (inputs(95)) and not (inputs(8));
    layer0_outputs(1351) <= not((inputs(56)) or (inputs(245)));
    layer0_outputs(1352) <= not((inputs(75)) or (inputs(95)));
    layer0_outputs(1353) <= not((inputs(45)) or (inputs(59)));
    layer0_outputs(1354) <= not(inputs(21));
    layer0_outputs(1355) <= (inputs(24)) and not (inputs(230));
    layer0_outputs(1356) <= inputs(98);
    layer0_outputs(1357) <= (inputs(249)) and not (inputs(12));
    layer0_outputs(1358) <= inputs(142);
    layer0_outputs(1359) <= not(inputs(149));
    layer0_outputs(1360) <= not(inputs(38));
    layer0_outputs(1361) <= not(inputs(60));
    layer0_outputs(1362) <= (inputs(243)) and not (inputs(137));
    layer0_outputs(1363) <= '1';
    layer0_outputs(1364) <= not(inputs(219));
    layer0_outputs(1365) <= (inputs(165)) or (inputs(219));
    layer0_outputs(1366) <= (inputs(69)) and not (inputs(211));
    layer0_outputs(1367) <= not((inputs(254)) or (inputs(43)));
    layer0_outputs(1368) <= (inputs(79)) and (inputs(225));
    layer0_outputs(1369) <= not(inputs(213));
    layer0_outputs(1370) <= not(inputs(242)) or (inputs(122));
    layer0_outputs(1371) <= (inputs(255)) and not (inputs(92));
    layer0_outputs(1372) <= not(inputs(162));
    layer0_outputs(1373) <= not((inputs(235)) or (inputs(85)));
    layer0_outputs(1374) <= not(inputs(133)) or (inputs(253));
    layer0_outputs(1375) <= not((inputs(23)) or (inputs(194)));
    layer0_outputs(1376) <= not((inputs(108)) xor (inputs(111)));
    layer0_outputs(1377) <= '1';
    layer0_outputs(1378) <= (inputs(41)) and not (inputs(103));
    layer0_outputs(1379) <= not((inputs(250)) and (inputs(150)));
    layer0_outputs(1380) <= inputs(28);
    layer0_outputs(1381) <= not((inputs(251)) and (inputs(197)));
    layer0_outputs(1382) <= not((inputs(236)) and (inputs(131)));
    layer0_outputs(1383) <= not(inputs(8));
    layer0_outputs(1384) <= not(inputs(30)) or (inputs(153));
    layer0_outputs(1385) <= not(inputs(16)) or (inputs(80));
    layer0_outputs(1386) <= (inputs(209)) or (inputs(128));
    layer0_outputs(1387) <= '0';
    layer0_outputs(1388) <= not(inputs(24));
    layer0_outputs(1389) <= not(inputs(166));
    layer0_outputs(1390) <= '0';
    layer0_outputs(1391) <= (inputs(153)) or (inputs(66));
    layer0_outputs(1392) <= not(inputs(86)) or (inputs(81));
    layer0_outputs(1393) <= (inputs(41)) or (inputs(71));
    layer0_outputs(1394) <= '1';
    layer0_outputs(1395) <= '0';
    layer0_outputs(1396) <= '1';
    layer0_outputs(1397) <= '0';
    layer0_outputs(1398) <= not((inputs(171)) and (inputs(174)));
    layer0_outputs(1399) <= inputs(90);
    layer0_outputs(1400) <= inputs(104);
    layer0_outputs(1401) <= not(inputs(220)) or (inputs(92));
    layer0_outputs(1402) <= (inputs(223)) and not (inputs(235));
    layer0_outputs(1403) <= (inputs(168)) and not (inputs(16));
    layer0_outputs(1404) <= (inputs(224)) or (inputs(201));
    layer0_outputs(1405) <= not((inputs(66)) xor (inputs(81)));
    layer0_outputs(1406) <= not(inputs(38));
    layer0_outputs(1407) <= (inputs(12)) and not (inputs(25));
    layer0_outputs(1408) <= not((inputs(248)) or (inputs(93)));
    layer0_outputs(1409) <= (inputs(22)) and not (inputs(129));
    layer0_outputs(1410) <= (inputs(255)) or (inputs(208));
    layer0_outputs(1411) <= not(inputs(135)) or (inputs(143));
    layer0_outputs(1412) <= '1';
    layer0_outputs(1413) <= not(inputs(200)) or (inputs(139));
    layer0_outputs(1414) <= not((inputs(250)) or (inputs(198)));
    layer0_outputs(1415) <= not((inputs(144)) or (inputs(30)));
    layer0_outputs(1416) <= (inputs(223)) and not (inputs(46));
    layer0_outputs(1417) <= not((inputs(48)) xor (inputs(90)));
    layer0_outputs(1418) <= not(inputs(123));
    layer0_outputs(1419) <= not((inputs(149)) or (inputs(198)));
    layer0_outputs(1420) <= (inputs(80)) or (inputs(149));
    layer0_outputs(1421) <= not((inputs(78)) or (inputs(186)));
    layer0_outputs(1422) <= '0';
    layer0_outputs(1423) <= not((inputs(81)) and (inputs(130)));
    layer0_outputs(1424) <= '1';
    layer0_outputs(1425) <= '1';
    layer0_outputs(1426) <= (inputs(1)) and (inputs(200));
    layer0_outputs(1427) <= (inputs(103)) and not (inputs(98));
    layer0_outputs(1428) <= not(inputs(123)) or (inputs(192));
    layer0_outputs(1429) <= not((inputs(3)) or (inputs(104)));
    layer0_outputs(1430) <= (inputs(4)) xor (inputs(59));
    layer0_outputs(1431) <= not(inputs(160));
    layer0_outputs(1432) <= not(inputs(118));
    layer0_outputs(1433) <= not((inputs(19)) or (inputs(212)));
    layer0_outputs(1434) <= '1';
    layer0_outputs(1435) <= inputs(169);
    layer0_outputs(1436) <= not(inputs(245));
    layer0_outputs(1437) <= (inputs(176)) or (inputs(32));
    layer0_outputs(1438) <= (inputs(68)) or (inputs(114));
    layer0_outputs(1439) <= not(inputs(202));
    layer0_outputs(1440) <= '1';
    layer0_outputs(1441) <= (inputs(97)) or (inputs(93));
    layer0_outputs(1442) <= not((inputs(207)) and (inputs(104)));
    layer0_outputs(1443) <= not(inputs(196));
    layer0_outputs(1444) <= (inputs(35)) and (inputs(103));
    layer0_outputs(1445) <= not(inputs(116)) or (inputs(239));
    layer0_outputs(1446) <= (inputs(117)) and (inputs(147));
    layer0_outputs(1447) <= (inputs(242)) or (inputs(161));
    layer0_outputs(1448) <= (inputs(94)) and not (inputs(92));
    layer0_outputs(1449) <= '1';
    layer0_outputs(1450) <= inputs(32);
    layer0_outputs(1451) <= inputs(116);
    layer0_outputs(1452) <= not(inputs(195));
    layer0_outputs(1453) <= not(inputs(118));
    layer0_outputs(1454) <= '0';
    layer0_outputs(1455) <= '1';
    layer0_outputs(1456) <= '0';
    layer0_outputs(1457) <= '1';
    layer0_outputs(1458) <= inputs(120);
    layer0_outputs(1459) <= (inputs(175)) or (inputs(120));
    layer0_outputs(1460) <= '1';
    layer0_outputs(1461) <= '1';
    layer0_outputs(1462) <= not(inputs(76));
    layer0_outputs(1463) <= inputs(103);
    layer0_outputs(1464) <= not(inputs(169));
    layer0_outputs(1465) <= not((inputs(202)) and (inputs(67)));
    layer0_outputs(1466) <= not((inputs(31)) and (inputs(184)));
    layer0_outputs(1467) <= '0';
    layer0_outputs(1468) <= not((inputs(51)) and (inputs(89)));
    layer0_outputs(1469) <= not(inputs(163));
    layer0_outputs(1470) <= '1';
    layer0_outputs(1471) <= not(inputs(47)) or (inputs(191));
    layer0_outputs(1472) <= '1';
    layer0_outputs(1473) <= '0';
    layer0_outputs(1474) <= not((inputs(109)) or (inputs(174)));
    layer0_outputs(1475) <= not(inputs(9));
    layer0_outputs(1476) <= (inputs(42)) or (inputs(34));
    layer0_outputs(1477) <= (inputs(20)) and not (inputs(203));
    layer0_outputs(1478) <= not((inputs(229)) and (inputs(28)));
    layer0_outputs(1479) <= inputs(73);
    layer0_outputs(1480) <= not(inputs(194));
    layer0_outputs(1481) <= inputs(206);
    layer0_outputs(1482) <= (inputs(68)) and not (inputs(154));
    layer0_outputs(1483) <= not((inputs(165)) or (inputs(190)));
    layer0_outputs(1484) <= not(inputs(239)) or (inputs(176));
    layer0_outputs(1485) <= not((inputs(181)) or (inputs(168)));
    layer0_outputs(1486) <= '0';
    layer0_outputs(1487) <= not((inputs(178)) or (inputs(174)));
    layer0_outputs(1488) <= (inputs(68)) and not (inputs(236));
    layer0_outputs(1489) <= not(inputs(0));
    layer0_outputs(1490) <= not((inputs(100)) and (inputs(128)));
    layer0_outputs(1491) <= (inputs(19)) and (inputs(73));
    layer0_outputs(1492) <= not((inputs(240)) and (inputs(204)));
    layer0_outputs(1493) <= (inputs(121)) and (inputs(47));
    layer0_outputs(1494) <= not(inputs(200));
    layer0_outputs(1495) <= not(inputs(71));
    layer0_outputs(1496) <= '0';
    layer0_outputs(1497) <= '1';
    layer0_outputs(1498) <= (inputs(247)) and not (inputs(17));
    layer0_outputs(1499) <= inputs(155);
    layer0_outputs(1500) <= '0';
    layer0_outputs(1501) <= '1';
    layer0_outputs(1502) <= inputs(158);
    layer0_outputs(1503) <= not((inputs(48)) or (inputs(96)));
    layer0_outputs(1504) <= (inputs(220)) and (inputs(72));
    layer0_outputs(1505) <= not(inputs(229));
    layer0_outputs(1506) <= '1';
    layer0_outputs(1507) <= not((inputs(220)) and (inputs(74)));
    layer0_outputs(1508) <= not((inputs(50)) xor (inputs(140)));
    layer0_outputs(1509) <= inputs(76);
    layer0_outputs(1510) <= (inputs(177)) and not (inputs(52));
    layer0_outputs(1511) <= (inputs(121)) and not (inputs(127));
    layer0_outputs(1512) <= '1';
    layer0_outputs(1513) <= not((inputs(255)) or (inputs(2)));
    layer0_outputs(1514) <= (inputs(204)) and (inputs(192));
    layer0_outputs(1515) <= inputs(179);
    layer0_outputs(1516) <= (inputs(195)) and not (inputs(62));
    layer0_outputs(1517) <= '0';
    layer0_outputs(1518) <= not(inputs(83)) or (inputs(56));
    layer0_outputs(1519) <= not((inputs(245)) and (inputs(187)));
    layer0_outputs(1520) <= (inputs(193)) and not (inputs(4));
    layer0_outputs(1521) <= not(inputs(28)) or (inputs(149));
    layer0_outputs(1522) <= not(inputs(25));
    layer0_outputs(1523) <= not(inputs(40));
    layer0_outputs(1524) <= not(inputs(38)) or (inputs(152));
    layer0_outputs(1525) <= not(inputs(162));
    layer0_outputs(1526) <= not(inputs(209)) or (inputs(240));
    layer0_outputs(1527) <= (inputs(76)) or (inputs(13));
    layer0_outputs(1528) <= (inputs(253)) and (inputs(141));
    layer0_outputs(1529) <= not((inputs(164)) or (inputs(165)));
    layer0_outputs(1530) <= not(inputs(247));
    layer0_outputs(1531) <= '0';
    layer0_outputs(1532) <= not((inputs(64)) or (inputs(37)));
    layer0_outputs(1533) <= (inputs(111)) and not (inputs(57));
    layer0_outputs(1534) <= '1';
    layer0_outputs(1535) <= not(inputs(104)) or (inputs(221));
    layer0_outputs(1536) <= '0';
    layer0_outputs(1537) <= '0';
    layer0_outputs(1538) <= inputs(91);
    layer0_outputs(1539) <= (inputs(116)) and not (inputs(5));
    layer0_outputs(1540) <= '1';
    layer0_outputs(1541) <= (inputs(164)) and not (inputs(239));
    layer0_outputs(1542) <= not(inputs(82)) or (inputs(227));
    layer0_outputs(1543) <= '0';
    layer0_outputs(1544) <= inputs(173);
    layer0_outputs(1545) <= inputs(31);
    layer0_outputs(1546) <= '1';
    layer0_outputs(1547) <= not((inputs(155)) or (inputs(107)));
    layer0_outputs(1548) <= inputs(34);
    layer0_outputs(1549) <= not(inputs(45));
    layer0_outputs(1550) <= not((inputs(156)) or (inputs(122)));
    layer0_outputs(1551) <= '0';
    layer0_outputs(1552) <= inputs(182);
    layer0_outputs(1553) <= not(inputs(91)) or (inputs(136));
    layer0_outputs(1554) <= (inputs(81)) and not (inputs(235));
    layer0_outputs(1555) <= not(inputs(46));
    layer0_outputs(1556) <= '0';
    layer0_outputs(1557) <= not(inputs(92)) or (inputs(0));
    layer0_outputs(1558) <= '0';
    layer0_outputs(1559) <= inputs(224);
    layer0_outputs(1560) <= not(inputs(27));
    layer0_outputs(1561) <= not(inputs(211));
    layer0_outputs(1562) <= not(inputs(132)) or (inputs(197));
    layer0_outputs(1563) <= '0';
    layer0_outputs(1564) <= inputs(25);
    layer0_outputs(1565) <= not(inputs(15));
    layer0_outputs(1566) <= not((inputs(39)) or (inputs(11)));
    layer0_outputs(1567) <= not(inputs(40)) or (inputs(89));
    layer0_outputs(1568) <= '1';
    layer0_outputs(1569) <= not(inputs(52));
    layer0_outputs(1570) <= not(inputs(201));
    layer0_outputs(1571) <= not(inputs(111));
    layer0_outputs(1572) <= (inputs(20)) and (inputs(72));
    layer0_outputs(1573) <= not(inputs(41));
    layer0_outputs(1574) <= inputs(47);
    layer0_outputs(1575) <= (inputs(74)) and not (inputs(54));
    layer0_outputs(1576) <= not(inputs(118)) or (inputs(25));
    layer0_outputs(1577) <= '0';
    layer0_outputs(1578) <= not((inputs(233)) and (inputs(105)));
    layer0_outputs(1579) <= not(inputs(154));
    layer0_outputs(1580) <= not(inputs(56)) or (inputs(136));
    layer0_outputs(1581) <= inputs(182);
    layer0_outputs(1582) <= not(inputs(205)) or (inputs(108));
    layer0_outputs(1583) <= not(inputs(89)) or (inputs(38));
    layer0_outputs(1584) <= not(inputs(67));
    layer0_outputs(1585) <= (inputs(218)) and not (inputs(198));
    layer0_outputs(1586) <= inputs(93);
    layer0_outputs(1587) <= (inputs(75)) and not (inputs(176));
    layer0_outputs(1588) <= not(inputs(229));
    layer0_outputs(1589) <= (inputs(176)) and not (inputs(166));
    layer0_outputs(1590) <= (inputs(104)) or (inputs(239));
    layer0_outputs(1591) <= '1';
    layer0_outputs(1592) <= inputs(151);
    layer0_outputs(1593) <= not(inputs(224)) or (inputs(100));
    layer0_outputs(1594) <= not(inputs(241)) or (inputs(145));
    layer0_outputs(1595) <= (inputs(101)) and not (inputs(95));
    layer0_outputs(1596) <= '1';
    layer0_outputs(1597) <= (inputs(91)) or (inputs(157));
    layer0_outputs(1598) <= not(inputs(178));
    layer0_outputs(1599) <= not(inputs(45)) or (inputs(103));
    layer0_outputs(1600) <= '0';
    layer0_outputs(1601) <= not(inputs(63)) or (inputs(222));
    layer0_outputs(1602) <= (inputs(3)) or (inputs(195));
    layer0_outputs(1603) <= not(inputs(23)) or (inputs(124));
    layer0_outputs(1604) <= inputs(164);
    layer0_outputs(1605) <= not(inputs(68));
    layer0_outputs(1606) <= (inputs(56)) and (inputs(39));
    layer0_outputs(1607) <= (inputs(48)) and not (inputs(29));
    layer0_outputs(1608) <= inputs(68);
    layer0_outputs(1609) <= '0';
    layer0_outputs(1610) <= not(inputs(7)) or (inputs(239));
    layer0_outputs(1611) <= inputs(19);
    layer0_outputs(1612) <= not(inputs(234)) or (inputs(29));
    layer0_outputs(1613) <= not((inputs(134)) and (inputs(189)));
    layer0_outputs(1614) <= '0';
    layer0_outputs(1615) <= '0';
    layer0_outputs(1616) <= not(inputs(222)) or (inputs(219));
    layer0_outputs(1617) <= not(inputs(70));
    layer0_outputs(1618) <= not(inputs(184));
    layer0_outputs(1619) <= (inputs(1)) xor (inputs(227));
    layer0_outputs(1620) <= not(inputs(152));
    layer0_outputs(1621) <= inputs(63);
    layer0_outputs(1622) <= not(inputs(197)) or (inputs(28));
    layer0_outputs(1623) <= inputs(166);
    layer0_outputs(1624) <= not(inputs(50)) or (inputs(35));
    layer0_outputs(1625) <= not(inputs(227)) or (inputs(157));
    layer0_outputs(1626) <= '0';
    layer0_outputs(1627) <= '1';
    layer0_outputs(1628) <= (inputs(123)) and (inputs(55));
    layer0_outputs(1629) <= not(inputs(226));
    layer0_outputs(1630) <= not((inputs(177)) or (inputs(205)));
    layer0_outputs(1631) <= not((inputs(247)) and (inputs(199)));
    layer0_outputs(1632) <= (inputs(230)) and not (inputs(165));
    layer0_outputs(1633) <= (inputs(243)) and (inputs(240));
    layer0_outputs(1634) <= not(inputs(13)) or (inputs(163));
    layer0_outputs(1635) <= inputs(105);
    layer0_outputs(1636) <= '0';
    layer0_outputs(1637) <= inputs(114);
    layer0_outputs(1638) <= not(inputs(12)) or (inputs(146));
    layer0_outputs(1639) <= not((inputs(108)) or (inputs(171)));
    layer0_outputs(1640) <= not(inputs(52)) or (inputs(18));
    layer0_outputs(1641) <= (inputs(196)) or (inputs(149));
    layer0_outputs(1642) <= not((inputs(169)) or (inputs(4)));
    layer0_outputs(1643) <= not(inputs(8));
    layer0_outputs(1644) <= not(inputs(49));
    layer0_outputs(1645) <= not(inputs(187)) or (inputs(15));
    layer0_outputs(1646) <= (inputs(71)) xor (inputs(79));
    layer0_outputs(1647) <= '0';
    layer0_outputs(1648) <= not(inputs(7)) or (inputs(104));
    layer0_outputs(1649) <= (inputs(176)) xor (inputs(121));
    layer0_outputs(1650) <= (inputs(163)) or (inputs(195));
    layer0_outputs(1651) <= inputs(59);
    layer0_outputs(1652) <= '1';
    layer0_outputs(1653) <= not(inputs(139));
    layer0_outputs(1654) <= (inputs(173)) and (inputs(220));
    layer0_outputs(1655) <= inputs(153);
    layer0_outputs(1656) <= not(inputs(230)) or (inputs(207));
    layer0_outputs(1657) <= not(inputs(204)) or (inputs(30));
    layer0_outputs(1658) <= '0';
    layer0_outputs(1659) <= '0';
    layer0_outputs(1660) <= (inputs(239)) or (inputs(195));
    layer0_outputs(1661) <= not((inputs(95)) or (inputs(139)));
    layer0_outputs(1662) <= not(inputs(35)) or (inputs(154));
    layer0_outputs(1663) <= (inputs(101)) or (inputs(177));
    layer0_outputs(1664) <= '1';
    layer0_outputs(1665) <= not((inputs(92)) xor (inputs(222)));
    layer0_outputs(1666) <= (inputs(202)) and not (inputs(139));
    layer0_outputs(1667) <= not(inputs(156));
    layer0_outputs(1668) <= not(inputs(8)) or (inputs(13));
    layer0_outputs(1669) <= '0';
    layer0_outputs(1670) <= inputs(197);
    layer0_outputs(1671) <= not(inputs(88));
    layer0_outputs(1672) <= (inputs(139)) xor (inputs(80));
    layer0_outputs(1673) <= '0';
    layer0_outputs(1674) <= (inputs(51)) or (inputs(185));
    layer0_outputs(1675) <= inputs(182);
    layer0_outputs(1676) <= (inputs(226)) and (inputs(245));
    layer0_outputs(1677) <= inputs(100);
    layer0_outputs(1678) <= not(inputs(165));
    layer0_outputs(1679) <= not(inputs(189)) or (inputs(18));
    layer0_outputs(1680) <= '1';
    layer0_outputs(1681) <= not((inputs(231)) or (inputs(54)));
    layer0_outputs(1682) <= not(inputs(184));
    layer0_outputs(1683) <= '0';
    layer0_outputs(1684) <= (inputs(189)) and not (inputs(115));
    layer0_outputs(1685) <= not(inputs(3)) or (inputs(232));
    layer0_outputs(1686) <= '0';
    layer0_outputs(1687) <= not(inputs(165)) or (inputs(14));
    layer0_outputs(1688) <= not(inputs(85)) or (inputs(112));
    layer0_outputs(1689) <= not((inputs(108)) and (inputs(44)));
    layer0_outputs(1690) <= '1';
    layer0_outputs(1691) <= inputs(137);
    layer0_outputs(1692) <= (inputs(162)) or (inputs(160));
    layer0_outputs(1693) <= not(inputs(245));
    layer0_outputs(1694) <= not(inputs(132)) or (inputs(1));
    layer0_outputs(1695) <= not(inputs(217));
    layer0_outputs(1696) <= '0';
    layer0_outputs(1697) <= inputs(119);
    layer0_outputs(1698) <= not(inputs(244));
    layer0_outputs(1699) <= (inputs(146)) and (inputs(231));
    layer0_outputs(1700) <= '1';
    layer0_outputs(1701) <= not(inputs(71)) or (inputs(31));
    layer0_outputs(1702) <= not(inputs(129));
    layer0_outputs(1703) <= (inputs(210)) or (inputs(230));
    layer0_outputs(1704) <= inputs(94);
    layer0_outputs(1705) <= (inputs(63)) and (inputs(13));
    layer0_outputs(1706) <= inputs(126);
    layer0_outputs(1707) <= '0';
    layer0_outputs(1708) <= inputs(98);
    layer0_outputs(1709) <= not(inputs(112));
    layer0_outputs(1710) <= not(inputs(236)) or (inputs(84));
    layer0_outputs(1711) <= '1';
    layer0_outputs(1712) <= (inputs(99)) or (inputs(172));
    layer0_outputs(1713) <= (inputs(186)) and not (inputs(197));
    layer0_outputs(1714) <= not(inputs(83));
    layer0_outputs(1715) <= (inputs(48)) and (inputs(25));
    layer0_outputs(1716) <= not((inputs(84)) or (inputs(103)));
    layer0_outputs(1717) <= not(inputs(188));
    layer0_outputs(1718) <= '0';
    layer0_outputs(1719) <= inputs(83);
    layer0_outputs(1720) <= (inputs(173)) and not (inputs(230));
    layer0_outputs(1721) <= (inputs(34)) or (inputs(196));
    layer0_outputs(1722) <= inputs(42);
    layer0_outputs(1723) <= not((inputs(142)) or (inputs(233)));
    layer0_outputs(1724) <= (inputs(26)) or (inputs(175));
    layer0_outputs(1725) <= not(inputs(2));
    layer0_outputs(1726) <= not(inputs(20)) or (inputs(162));
    layer0_outputs(1727) <= not(inputs(132));
    layer0_outputs(1728) <= not((inputs(118)) xor (inputs(1)));
    layer0_outputs(1729) <= inputs(140);
    layer0_outputs(1730) <= not(inputs(162));
    layer0_outputs(1731) <= (inputs(228)) and not (inputs(84));
    layer0_outputs(1732) <= '0';
    layer0_outputs(1733) <= not(inputs(151)) or (inputs(222));
    layer0_outputs(1734) <= '1';
    layer0_outputs(1735) <= '1';
    layer0_outputs(1736) <= not(inputs(238));
    layer0_outputs(1737) <= not(inputs(162)) or (inputs(159));
    layer0_outputs(1738) <= inputs(151);
    layer0_outputs(1739) <= '0';
    layer0_outputs(1740) <= not((inputs(200)) xor (inputs(158)));
    layer0_outputs(1741) <= '0';
    layer0_outputs(1742) <= '0';
    layer0_outputs(1743) <= '0';
    layer0_outputs(1744) <= (inputs(27)) or (inputs(47));
    layer0_outputs(1745) <= '1';
    layer0_outputs(1746) <= not((inputs(99)) or (inputs(97)));
    layer0_outputs(1747) <= '1';
    layer0_outputs(1748) <= (inputs(31)) and not (inputs(37));
    layer0_outputs(1749) <= (inputs(95)) xor (inputs(47));
    layer0_outputs(1750) <= not(inputs(156)) or (inputs(215));
    layer0_outputs(1751) <= '0';
    layer0_outputs(1752) <= not((inputs(76)) and (inputs(26)));
    layer0_outputs(1753) <= not(inputs(61));
    layer0_outputs(1754) <= '1';
    layer0_outputs(1755) <= not(inputs(233));
    layer0_outputs(1756) <= inputs(210);
    layer0_outputs(1757) <= '1';
    layer0_outputs(1758) <= not(inputs(5));
    layer0_outputs(1759) <= not(inputs(148)) or (inputs(18));
    layer0_outputs(1760) <= not(inputs(214)) or (inputs(135));
    layer0_outputs(1761) <= not(inputs(150));
    layer0_outputs(1762) <= inputs(213);
    layer0_outputs(1763) <= inputs(236);
    layer0_outputs(1764) <= '0';
    layer0_outputs(1765) <= not(inputs(77)) or (inputs(182));
    layer0_outputs(1766) <= inputs(118);
    layer0_outputs(1767) <= not(inputs(0)) or (inputs(81));
    layer0_outputs(1768) <= (inputs(83)) and not (inputs(209));
    layer0_outputs(1769) <= inputs(175);
    layer0_outputs(1770) <= (inputs(3)) and (inputs(44));
    layer0_outputs(1771) <= (inputs(222)) or (inputs(33));
    layer0_outputs(1772) <= (inputs(251)) or (inputs(234));
    layer0_outputs(1773) <= (inputs(179)) or (inputs(204));
    layer0_outputs(1774) <= inputs(138);
    layer0_outputs(1775) <= not(inputs(134));
    layer0_outputs(1776) <= '0';
    layer0_outputs(1777) <= '0';
    layer0_outputs(1778) <= (inputs(37)) and not (inputs(144));
    layer0_outputs(1779) <= not((inputs(216)) and (inputs(174)));
    layer0_outputs(1780) <= not(inputs(96));
    layer0_outputs(1781) <= not(inputs(116));
    layer0_outputs(1782) <= (inputs(96)) and not (inputs(6));
    layer0_outputs(1783) <= (inputs(5)) and not (inputs(252));
    layer0_outputs(1784) <= inputs(107);
    layer0_outputs(1785) <= (inputs(215)) and not (inputs(203));
    layer0_outputs(1786) <= '0';
    layer0_outputs(1787) <= inputs(158);
    layer0_outputs(1788) <= inputs(194);
    layer0_outputs(1789) <= not(inputs(162));
    layer0_outputs(1790) <= (inputs(6)) and (inputs(31));
    layer0_outputs(1791) <= (inputs(197)) or (inputs(53));
    layer0_outputs(1792) <= '0';
    layer0_outputs(1793) <= not(inputs(93));
    layer0_outputs(1794) <= (inputs(138)) xor (inputs(160));
    layer0_outputs(1795) <= not((inputs(161)) xor (inputs(218)));
    layer0_outputs(1796) <= (inputs(44)) or (inputs(109));
    layer0_outputs(1797) <= (inputs(94)) and (inputs(42));
    layer0_outputs(1798) <= '0';
    layer0_outputs(1799) <= (inputs(87)) or (inputs(149));
    layer0_outputs(1800) <= inputs(241);
    layer0_outputs(1801) <= not(inputs(165)) or (inputs(50));
    layer0_outputs(1802) <= not(inputs(168));
    layer0_outputs(1803) <= inputs(143);
    layer0_outputs(1804) <= not((inputs(172)) and (inputs(250)));
    layer0_outputs(1805) <= not(inputs(255)) or (inputs(252));
    layer0_outputs(1806) <= (inputs(89)) and (inputs(243));
    layer0_outputs(1807) <= not((inputs(98)) and (inputs(128)));
    layer0_outputs(1808) <= (inputs(160)) and not (inputs(129));
    layer0_outputs(1809) <= (inputs(21)) or (inputs(166));
    layer0_outputs(1810) <= not((inputs(160)) xor (inputs(46)));
    layer0_outputs(1811) <= (inputs(36)) or (inputs(70));
    layer0_outputs(1812) <= not(inputs(18));
    layer0_outputs(1813) <= (inputs(64)) and not (inputs(181));
    layer0_outputs(1814) <= (inputs(133)) and (inputs(68));
    layer0_outputs(1815) <= not(inputs(74));
    layer0_outputs(1816) <= not(inputs(28)) or (inputs(173));
    layer0_outputs(1817) <= (inputs(187)) or (inputs(218));
    layer0_outputs(1818) <= not(inputs(19));
    layer0_outputs(1819) <= (inputs(229)) and not (inputs(151));
    layer0_outputs(1820) <= not(inputs(156));
    layer0_outputs(1821) <= '1';
    layer0_outputs(1822) <= '1';
    layer0_outputs(1823) <= not(inputs(211));
    layer0_outputs(1824) <= not((inputs(77)) or (inputs(107)));
    layer0_outputs(1825) <= '0';
    layer0_outputs(1826) <= inputs(225);
    layer0_outputs(1827) <= '0';
    layer0_outputs(1828) <= not(inputs(240)) or (inputs(133));
    layer0_outputs(1829) <= (inputs(147)) and not (inputs(248));
    layer0_outputs(1830) <= not((inputs(59)) and (inputs(18)));
    layer0_outputs(1831) <= not(inputs(217));
    layer0_outputs(1832) <= not(inputs(255)) or (inputs(43));
    layer0_outputs(1833) <= '0';
    layer0_outputs(1834) <= '0';
    layer0_outputs(1835) <= inputs(254);
    layer0_outputs(1836) <= inputs(58);
    layer0_outputs(1837) <= not((inputs(111)) or (inputs(196)));
    layer0_outputs(1838) <= '1';
    layer0_outputs(1839) <= not((inputs(238)) xor (inputs(238)));
    layer0_outputs(1840) <= not((inputs(179)) and (inputs(145)));
    layer0_outputs(1841) <= not(inputs(213));
    layer0_outputs(1842) <= '0';
    layer0_outputs(1843) <= (inputs(128)) or (inputs(155));
    layer0_outputs(1844) <= inputs(46);
    layer0_outputs(1845) <= not(inputs(91)) or (inputs(88));
    layer0_outputs(1846) <= (inputs(149)) or (inputs(126));
    layer0_outputs(1847) <= not((inputs(232)) and (inputs(92)));
    layer0_outputs(1848) <= '1';
    layer0_outputs(1849) <= not(inputs(171)) or (inputs(98));
    layer0_outputs(1850) <= not((inputs(250)) and (inputs(253)));
    layer0_outputs(1851) <= (inputs(151)) or (inputs(123));
    layer0_outputs(1852) <= '1';
    layer0_outputs(1853) <= not((inputs(61)) or (inputs(163)));
    layer0_outputs(1854) <= not((inputs(206)) or (inputs(66)));
    layer0_outputs(1855) <= '0';
    layer0_outputs(1856) <= inputs(106);
    layer0_outputs(1857) <= '0';
    layer0_outputs(1858) <= '0';
    layer0_outputs(1859) <= (inputs(161)) and not (inputs(87));
    layer0_outputs(1860) <= (inputs(117)) and not (inputs(2));
    layer0_outputs(1861) <= (inputs(35)) or (inputs(153));
    layer0_outputs(1862) <= not(inputs(213));
    layer0_outputs(1863) <= not(inputs(164));
    layer0_outputs(1864) <= not(inputs(44)) or (inputs(230));
    layer0_outputs(1865) <= not((inputs(163)) or (inputs(250)));
    layer0_outputs(1866) <= not((inputs(8)) and (inputs(59)));
    layer0_outputs(1867) <= (inputs(165)) and not (inputs(30));
    layer0_outputs(1868) <= not((inputs(147)) and (inputs(108)));
    layer0_outputs(1869) <= '1';
    layer0_outputs(1870) <= '1';
    layer0_outputs(1871) <= not(inputs(14));
    layer0_outputs(1872) <= inputs(155);
    layer0_outputs(1873) <= inputs(121);
    layer0_outputs(1874) <= (inputs(206)) and not (inputs(122));
    layer0_outputs(1875) <= '0';
    layer0_outputs(1876) <= (inputs(229)) or (inputs(157));
    layer0_outputs(1877) <= '1';
    layer0_outputs(1878) <= (inputs(221)) xor (inputs(173));
    layer0_outputs(1879) <= not((inputs(198)) and (inputs(39)));
    layer0_outputs(1880) <= not(inputs(194));
    layer0_outputs(1881) <= (inputs(191)) or (inputs(232));
    layer0_outputs(1882) <= not(inputs(115));
    layer0_outputs(1883) <= not(inputs(183));
    layer0_outputs(1884) <= '0';
    layer0_outputs(1885) <= not(inputs(222));
    layer0_outputs(1886) <= (inputs(231)) or (inputs(192));
    layer0_outputs(1887) <= inputs(202);
    layer0_outputs(1888) <= inputs(183);
    layer0_outputs(1889) <= inputs(58);
    layer0_outputs(1890) <= (inputs(0)) xor (inputs(0));
    layer0_outputs(1891) <= inputs(100);
    layer0_outputs(1892) <= not(inputs(39)) or (inputs(219));
    layer0_outputs(1893) <= (inputs(197)) or (inputs(185));
    layer0_outputs(1894) <= not(inputs(76)) or (inputs(29));
    layer0_outputs(1895) <= inputs(223);
    layer0_outputs(1896) <= not(inputs(61)) or (inputs(86));
    layer0_outputs(1897) <= (inputs(183)) and (inputs(108));
    layer0_outputs(1898) <= not((inputs(76)) or (inputs(31)));
    layer0_outputs(1899) <= not(inputs(94)) or (inputs(136));
    layer0_outputs(1900) <= (inputs(69)) and (inputs(205));
    layer0_outputs(1901) <= '0';
    layer0_outputs(1902) <= (inputs(85)) and not (inputs(177));
    layer0_outputs(1903) <= '1';
    layer0_outputs(1904) <= not(inputs(84));
    layer0_outputs(1905) <= not(inputs(117));
    layer0_outputs(1906) <= (inputs(246)) or (inputs(111));
    layer0_outputs(1907) <= not(inputs(175));
    layer0_outputs(1908) <= not(inputs(203));
    layer0_outputs(1909) <= not((inputs(124)) or (inputs(92)));
    layer0_outputs(1910) <= (inputs(253)) and not (inputs(232));
    layer0_outputs(1911) <= (inputs(133)) and not (inputs(187));
    layer0_outputs(1912) <= (inputs(6)) or (inputs(69));
    layer0_outputs(1913) <= not(inputs(142)) or (inputs(240));
    layer0_outputs(1914) <= '1';
    layer0_outputs(1915) <= (inputs(240)) and not (inputs(45));
    layer0_outputs(1916) <= (inputs(218)) or (inputs(160));
    layer0_outputs(1917) <= inputs(56);
    layer0_outputs(1918) <= not(inputs(163));
    layer0_outputs(1919) <= not(inputs(245));
    layer0_outputs(1920) <= not(inputs(48));
    layer0_outputs(1921) <= not((inputs(15)) xor (inputs(51)));
    layer0_outputs(1922) <= not(inputs(156)) or (inputs(232));
    layer0_outputs(1923) <= '0';
    layer0_outputs(1924) <= not(inputs(151)) or (inputs(176));
    layer0_outputs(1925) <= not((inputs(79)) and (inputs(35)));
    layer0_outputs(1926) <= '1';
    layer0_outputs(1927) <= not(inputs(13));
    layer0_outputs(1928) <= inputs(89);
    layer0_outputs(1929) <= inputs(240);
    layer0_outputs(1930) <= '1';
    layer0_outputs(1931) <= not((inputs(42)) or (inputs(208)));
    layer0_outputs(1932) <= (inputs(136)) and not (inputs(233));
    layer0_outputs(1933) <= not(inputs(184));
    layer0_outputs(1934) <= not(inputs(25)) or (inputs(232));
    layer0_outputs(1935) <= '1';
    layer0_outputs(1936) <= (inputs(190)) xor (inputs(179));
    layer0_outputs(1937) <= '0';
    layer0_outputs(1938) <= not(inputs(122));
    layer0_outputs(1939) <= inputs(183);
    layer0_outputs(1940) <= not((inputs(140)) and (inputs(212)));
    layer0_outputs(1941) <= inputs(8);
    layer0_outputs(1942) <= not(inputs(106));
    layer0_outputs(1943) <= not(inputs(94));
    layer0_outputs(1944) <= not(inputs(58));
    layer0_outputs(1945) <= not((inputs(103)) or (inputs(118)));
    layer0_outputs(1946) <= inputs(253);
    layer0_outputs(1947) <= not(inputs(145));
    layer0_outputs(1948) <= (inputs(108)) and not (inputs(193));
    layer0_outputs(1949) <= inputs(177);
    layer0_outputs(1950) <= not((inputs(132)) and (inputs(252)));
    layer0_outputs(1951) <= '1';
    layer0_outputs(1952) <= '1';
    layer0_outputs(1953) <= (inputs(235)) and not (inputs(78));
    layer0_outputs(1954) <= '0';
    layer0_outputs(1955) <= inputs(112);
    layer0_outputs(1956) <= '1';
    layer0_outputs(1957) <= not((inputs(214)) or (inputs(11)));
    layer0_outputs(1958) <= not((inputs(163)) and (inputs(48)));
    layer0_outputs(1959) <= (inputs(218)) or (inputs(173));
    layer0_outputs(1960) <= inputs(61);
    layer0_outputs(1961) <= not(inputs(180));
    layer0_outputs(1962) <= '0';
    layer0_outputs(1963) <= '0';
    layer0_outputs(1964) <= '0';
    layer0_outputs(1965) <= not(inputs(139));
    layer0_outputs(1966) <= '0';
    layer0_outputs(1967) <= not(inputs(195));
    layer0_outputs(1968) <= (inputs(151)) and not (inputs(179));
    layer0_outputs(1969) <= not(inputs(101));
    layer0_outputs(1970) <= inputs(168);
    layer0_outputs(1971) <= inputs(202);
    layer0_outputs(1972) <= not((inputs(60)) and (inputs(186)));
    layer0_outputs(1973) <= not((inputs(148)) or (inputs(98)));
    layer0_outputs(1974) <= not((inputs(128)) or (inputs(76)));
    layer0_outputs(1975) <= not(inputs(98)) or (inputs(171));
    layer0_outputs(1976) <= (inputs(231)) and not (inputs(110));
    layer0_outputs(1977) <= (inputs(204)) or (inputs(102));
    layer0_outputs(1978) <= not(inputs(252)) or (inputs(173));
    layer0_outputs(1979) <= (inputs(9)) and not (inputs(24));
    layer0_outputs(1980) <= not(inputs(136)) or (inputs(242));
    layer0_outputs(1981) <= inputs(224);
    layer0_outputs(1982) <= (inputs(179)) and not (inputs(107));
    layer0_outputs(1983) <= (inputs(89)) and not (inputs(16));
    layer0_outputs(1984) <= not(inputs(24)) or (inputs(226));
    layer0_outputs(1985) <= '1';
    layer0_outputs(1986) <= not((inputs(219)) xor (inputs(179)));
    layer0_outputs(1987) <= not((inputs(8)) or (inputs(212)));
    layer0_outputs(1988) <= not((inputs(101)) and (inputs(97)));
    layer0_outputs(1989) <= inputs(77);
    layer0_outputs(1990) <= (inputs(138)) and not (inputs(195));
    layer0_outputs(1991) <= inputs(27);
    layer0_outputs(1992) <= (inputs(122)) and not (inputs(122));
    layer0_outputs(1993) <= (inputs(190)) and (inputs(92));
    layer0_outputs(1994) <= not((inputs(108)) or (inputs(222)));
    layer0_outputs(1995) <= not((inputs(250)) and (inputs(180)));
    layer0_outputs(1996) <= (inputs(213)) and (inputs(60));
    layer0_outputs(1997) <= inputs(117);
    layer0_outputs(1998) <= not((inputs(209)) or (inputs(96)));
    layer0_outputs(1999) <= inputs(106);
    layer0_outputs(2000) <= (inputs(53)) and not (inputs(204));
    layer0_outputs(2001) <= (inputs(135)) xor (inputs(153));
    layer0_outputs(2002) <= not(inputs(235));
    layer0_outputs(2003) <= (inputs(52)) xor (inputs(179));
    layer0_outputs(2004) <= '0';
    layer0_outputs(2005) <= (inputs(209)) and (inputs(26));
    layer0_outputs(2006) <= (inputs(173)) xor (inputs(7));
    layer0_outputs(2007) <= not((inputs(148)) or (inputs(54)));
    layer0_outputs(2008) <= not(inputs(152));
    layer0_outputs(2009) <= (inputs(148)) and not (inputs(241));
    layer0_outputs(2010) <= not((inputs(212)) and (inputs(217)));
    layer0_outputs(2011) <= '0';
    layer0_outputs(2012) <= not(inputs(51)) or (inputs(90));
    layer0_outputs(2013) <= '1';
    layer0_outputs(2014) <= not((inputs(133)) and (inputs(205)));
    layer0_outputs(2015) <= (inputs(134)) or (inputs(235));
    layer0_outputs(2016) <= (inputs(194)) and not (inputs(129));
    layer0_outputs(2017) <= '1';
    layer0_outputs(2018) <= inputs(59);
    layer0_outputs(2019) <= (inputs(8)) and not (inputs(15));
    layer0_outputs(2020) <= not(inputs(16));
    layer0_outputs(2021) <= (inputs(255)) and not (inputs(97));
    layer0_outputs(2022) <= not(inputs(197)) or (inputs(112));
    layer0_outputs(2023) <= (inputs(85)) or (inputs(198));
    layer0_outputs(2024) <= not((inputs(90)) and (inputs(53)));
    layer0_outputs(2025) <= not(inputs(50)) or (inputs(248));
    layer0_outputs(2026) <= not(inputs(212));
    layer0_outputs(2027) <= inputs(181);
    layer0_outputs(2028) <= (inputs(177)) and not (inputs(248));
    layer0_outputs(2029) <= not((inputs(113)) and (inputs(2)));
    layer0_outputs(2030) <= '1';
    layer0_outputs(2031) <= (inputs(45)) or (inputs(145));
    layer0_outputs(2032) <= not(inputs(159));
    layer0_outputs(2033) <= not(inputs(8)) or (inputs(18));
    layer0_outputs(2034) <= not((inputs(180)) or (inputs(174)));
    layer0_outputs(2035) <= (inputs(95)) or (inputs(218));
    layer0_outputs(2036) <= inputs(138);
    layer0_outputs(2037) <= not(inputs(119));
    layer0_outputs(2038) <= inputs(151);
    layer0_outputs(2039) <= not((inputs(90)) and (inputs(229)));
    layer0_outputs(2040) <= '1';
    layer0_outputs(2041) <= not(inputs(68)) or (inputs(191));
    layer0_outputs(2042) <= not(inputs(247));
    layer0_outputs(2043) <= inputs(222);
    layer0_outputs(2044) <= (inputs(106)) and not (inputs(194));
    layer0_outputs(2045) <= (inputs(58)) and not (inputs(86));
    layer0_outputs(2046) <= not(inputs(82));
    layer0_outputs(2047) <= '1';
    layer0_outputs(2048) <= (inputs(147)) and not (inputs(133));
    layer0_outputs(2049) <= not(inputs(143));
    layer0_outputs(2050) <= '1';
    layer0_outputs(2051) <= '0';
    layer0_outputs(2052) <= '0';
    layer0_outputs(2053) <= '1';
    layer0_outputs(2054) <= not((inputs(183)) or (inputs(13)));
    layer0_outputs(2055) <= not(inputs(155));
    layer0_outputs(2056) <= (inputs(35)) and (inputs(247));
    layer0_outputs(2057) <= not(inputs(80)) or (inputs(83));
    layer0_outputs(2058) <= inputs(110);
    layer0_outputs(2059) <= inputs(50);
    layer0_outputs(2060) <= (inputs(73)) and not (inputs(43));
    layer0_outputs(2061) <= inputs(121);
    layer0_outputs(2062) <= (inputs(57)) and not (inputs(252));
    layer0_outputs(2063) <= not(inputs(135));
    layer0_outputs(2064) <= not((inputs(36)) or (inputs(10)));
    layer0_outputs(2065) <= not(inputs(131));
    layer0_outputs(2066) <= not(inputs(232));
    layer0_outputs(2067) <= not(inputs(221));
    layer0_outputs(2068) <= inputs(122);
    layer0_outputs(2069) <= not((inputs(5)) and (inputs(145)));
    layer0_outputs(2070) <= inputs(148);
    layer0_outputs(2071) <= not((inputs(189)) and (inputs(111)));
    layer0_outputs(2072) <= not(inputs(5)) or (inputs(89));
    layer0_outputs(2073) <= not(inputs(186)) or (inputs(21));
    layer0_outputs(2074) <= not(inputs(214));
    layer0_outputs(2075) <= '1';
    layer0_outputs(2076) <= not((inputs(97)) xor (inputs(69)));
    layer0_outputs(2077) <= inputs(85);
    layer0_outputs(2078) <= '0';
    layer0_outputs(2079) <= '1';
    layer0_outputs(2080) <= '0';
    layer0_outputs(2081) <= not((inputs(95)) or (inputs(33)));
    layer0_outputs(2082) <= '0';
    layer0_outputs(2083) <= '1';
    layer0_outputs(2084) <= (inputs(11)) and (inputs(220));
    layer0_outputs(2085) <= (inputs(189)) or (inputs(238));
    layer0_outputs(2086) <= (inputs(180)) xor (inputs(13));
    layer0_outputs(2087) <= not((inputs(152)) or (inputs(15)));
    layer0_outputs(2088) <= '1';
    layer0_outputs(2089) <= inputs(181);
    layer0_outputs(2090) <= not(inputs(224));
    layer0_outputs(2091) <= inputs(19);
    layer0_outputs(2092) <= inputs(88);
    layer0_outputs(2093) <= '1';
    layer0_outputs(2094) <= inputs(117);
    layer0_outputs(2095) <= not(inputs(18)) or (inputs(82));
    layer0_outputs(2096) <= not(inputs(165));
    layer0_outputs(2097) <= not(inputs(136)) or (inputs(216));
    layer0_outputs(2098) <= '1';
    layer0_outputs(2099) <= not(inputs(215)) or (inputs(123));
    layer0_outputs(2100) <= (inputs(210)) or (inputs(14));
    layer0_outputs(2101) <= inputs(233);
    layer0_outputs(2102) <= inputs(166);
    layer0_outputs(2103) <= (inputs(244)) or (inputs(246));
    layer0_outputs(2104) <= inputs(106);
    layer0_outputs(2105) <= not(inputs(202));
    layer0_outputs(2106) <= '0';
    layer0_outputs(2107) <= (inputs(158)) and not (inputs(36));
    layer0_outputs(2108) <= (inputs(65)) or (inputs(21));
    layer0_outputs(2109) <= (inputs(49)) or (inputs(53));
    layer0_outputs(2110) <= (inputs(181)) or (inputs(37));
    layer0_outputs(2111) <= not(inputs(55)) or (inputs(105));
    layer0_outputs(2112) <= '0';
    layer0_outputs(2113) <= '1';
    layer0_outputs(2114) <= (inputs(53)) and not (inputs(158));
    layer0_outputs(2115) <= not((inputs(245)) and (inputs(231)));
    layer0_outputs(2116) <= not((inputs(185)) and (inputs(32)));
    layer0_outputs(2117) <= (inputs(162)) or (inputs(202));
    layer0_outputs(2118) <= (inputs(130)) or (inputs(112));
    layer0_outputs(2119) <= not(inputs(20)) or (inputs(205));
    layer0_outputs(2120) <= inputs(16);
    layer0_outputs(2121) <= inputs(69);
    layer0_outputs(2122) <= not(inputs(240));
    layer0_outputs(2123) <= (inputs(202)) or (inputs(248));
    layer0_outputs(2124) <= inputs(93);
    layer0_outputs(2125) <= '0';
    layer0_outputs(2126) <= (inputs(7)) or (inputs(69));
    layer0_outputs(2127) <= '1';
    layer0_outputs(2128) <= (inputs(24)) and not (inputs(71));
    layer0_outputs(2129) <= not(inputs(163)) or (inputs(179));
    layer0_outputs(2130) <= inputs(240);
    layer0_outputs(2131) <= '0';
    layer0_outputs(2132) <= (inputs(208)) or (inputs(72));
    layer0_outputs(2133) <= (inputs(108)) and not (inputs(42));
    layer0_outputs(2134) <= (inputs(26)) or (inputs(51));
    layer0_outputs(2135) <= not(inputs(113));
    layer0_outputs(2136) <= '1';
    layer0_outputs(2137) <= inputs(17);
    layer0_outputs(2138) <= not(inputs(20)) or (inputs(210));
    layer0_outputs(2139) <= not(inputs(217)) or (inputs(63));
    layer0_outputs(2140) <= inputs(147);
    layer0_outputs(2141) <= inputs(248);
    layer0_outputs(2142) <= (inputs(238)) or (inputs(195));
    layer0_outputs(2143) <= '1';
    layer0_outputs(2144) <= '1';
    layer0_outputs(2145) <= '0';
    layer0_outputs(2146) <= not(inputs(134));
    layer0_outputs(2147) <= not(inputs(188)) or (inputs(12));
    layer0_outputs(2148) <= (inputs(124)) or (inputs(2));
    layer0_outputs(2149) <= inputs(185);
    layer0_outputs(2150) <= '0';
    layer0_outputs(2151) <= not((inputs(56)) and (inputs(170)));
    layer0_outputs(2152) <= (inputs(138)) and not (inputs(80));
    layer0_outputs(2153) <= (inputs(166)) or (inputs(59));
    layer0_outputs(2154) <= '1';
    layer0_outputs(2155) <= (inputs(81)) and (inputs(213));
    layer0_outputs(2156) <= '1';
    layer0_outputs(2157) <= '0';
    layer0_outputs(2158) <= not((inputs(87)) and (inputs(53)));
    layer0_outputs(2159) <= not(inputs(177));
    layer0_outputs(2160) <= '1';
    layer0_outputs(2161) <= not(inputs(131));
    layer0_outputs(2162) <= inputs(126);
    layer0_outputs(2163) <= '1';
    layer0_outputs(2164) <= not(inputs(246)) or (inputs(102));
    layer0_outputs(2165) <= inputs(47);
    layer0_outputs(2166) <= not(inputs(83));
    layer0_outputs(2167) <= inputs(130);
    layer0_outputs(2168) <= not(inputs(254));
    layer0_outputs(2169) <= not(inputs(208));
    layer0_outputs(2170) <= not(inputs(4)) or (inputs(221));
    layer0_outputs(2171) <= (inputs(198)) or (inputs(225));
    layer0_outputs(2172) <= not((inputs(198)) or (inputs(201)));
    layer0_outputs(2173) <= not(inputs(127)) or (inputs(154));
    layer0_outputs(2174) <= not(inputs(29));
    layer0_outputs(2175) <= not((inputs(200)) and (inputs(235)));
    layer0_outputs(2176) <= not((inputs(66)) or (inputs(76)));
    layer0_outputs(2177) <= (inputs(158)) and not (inputs(137));
    layer0_outputs(2178) <= not(inputs(229));
    layer0_outputs(2179) <= (inputs(191)) and not (inputs(7));
    layer0_outputs(2180) <= '0';
    layer0_outputs(2181) <= not(inputs(126));
    layer0_outputs(2182) <= not((inputs(196)) and (inputs(241)));
    layer0_outputs(2183) <= (inputs(24)) and not (inputs(86));
    layer0_outputs(2184) <= '0';
    layer0_outputs(2185) <= (inputs(188)) or (inputs(157));
    layer0_outputs(2186) <= (inputs(154)) and not (inputs(17));
    layer0_outputs(2187) <= not(inputs(246));
    layer0_outputs(2188) <= not((inputs(60)) and (inputs(237)));
    layer0_outputs(2189) <= not(inputs(133));
    layer0_outputs(2190) <= (inputs(15)) xor (inputs(88));
    layer0_outputs(2191) <= inputs(102);
    layer0_outputs(2192) <= not(inputs(7));
    layer0_outputs(2193) <= not(inputs(195));
    layer0_outputs(2194) <= (inputs(189)) and not (inputs(240));
    layer0_outputs(2195) <= inputs(2);
    layer0_outputs(2196) <= not((inputs(188)) or (inputs(11)));
    layer0_outputs(2197) <= not(inputs(193)) or (inputs(57));
    layer0_outputs(2198) <= inputs(243);
    layer0_outputs(2199) <= not(inputs(187)) or (inputs(59));
    layer0_outputs(2200) <= not((inputs(246)) and (inputs(125)));
    layer0_outputs(2201) <= (inputs(87)) and not (inputs(136));
    layer0_outputs(2202) <= '1';
    layer0_outputs(2203) <= not((inputs(64)) or (inputs(181)));
    layer0_outputs(2204) <= not((inputs(179)) or (inputs(11)));
    layer0_outputs(2205) <= not(inputs(9));
    layer0_outputs(2206) <= inputs(131);
    layer0_outputs(2207) <= not(inputs(69));
    layer0_outputs(2208) <= not(inputs(139));
    layer0_outputs(2209) <= '0';
    layer0_outputs(2210) <= (inputs(17)) and not (inputs(149));
    layer0_outputs(2211) <= not(inputs(57)) or (inputs(117));
    layer0_outputs(2212) <= (inputs(73)) and (inputs(130));
    layer0_outputs(2213) <= inputs(193);
    layer0_outputs(2214) <= inputs(168);
    layer0_outputs(2215) <= not(inputs(86));
    layer0_outputs(2216) <= not(inputs(164));
    layer0_outputs(2217) <= '1';
    layer0_outputs(2218) <= (inputs(60)) and (inputs(177));
    layer0_outputs(2219) <= '1';
    layer0_outputs(2220) <= not(inputs(37)) or (inputs(127));
    layer0_outputs(2221) <= not(inputs(80));
    layer0_outputs(2222) <= inputs(48);
    layer0_outputs(2223) <= (inputs(141)) or (inputs(3));
    layer0_outputs(2224) <= (inputs(234)) and (inputs(14));
    layer0_outputs(2225) <= (inputs(89)) and not (inputs(144));
    layer0_outputs(2226) <= (inputs(217)) and not (inputs(152));
    layer0_outputs(2227) <= not((inputs(99)) or (inputs(130)));
    layer0_outputs(2228) <= not((inputs(189)) and (inputs(162)));
    layer0_outputs(2229) <= not(inputs(136));
    layer0_outputs(2230) <= inputs(114);
    layer0_outputs(2231) <= (inputs(40)) or (inputs(113));
    layer0_outputs(2232) <= '0';
    layer0_outputs(2233) <= not((inputs(164)) or (inputs(154)));
    layer0_outputs(2234) <= (inputs(212)) or (inputs(197));
    layer0_outputs(2235) <= (inputs(64)) and (inputs(248));
    layer0_outputs(2236) <= inputs(106);
    layer0_outputs(2237) <= inputs(73);
    layer0_outputs(2238) <= not(inputs(199));
    layer0_outputs(2239) <= not(inputs(125));
    layer0_outputs(2240) <= (inputs(60)) and not (inputs(219));
    layer0_outputs(2241) <= (inputs(104)) or (inputs(192));
    layer0_outputs(2242) <= '1';
    layer0_outputs(2243) <= '1';
    layer0_outputs(2244) <= (inputs(77)) xor (inputs(134));
    layer0_outputs(2245) <= '1';
    layer0_outputs(2246) <= not(inputs(37)) or (inputs(251));
    layer0_outputs(2247) <= (inputs(237)) and not (inputs(14));
    layer0_outputs(2248) <= '0';
    layer0_outputs(2249) <= not(inputs(203));
    layer0_outputs(2250) <= (inputs(48)) and not (inputs(51));
    layer0_outputs(2251) <= '1';
    layer0_outputs(2252) <= inputs(255);
    layer0_outputs(2253) <= (inputs(189)) and not (inputs(125));
    layer0_outputs(2254) <= not(inputs(0));
    layer0_outputs(2255) <= not(inputs(132));
    layer0_outputs(2256) <= '0';
    layer0_outputs(2257) <= inputs(224);
    layer0_outputs(2258) <= (inputs(33)) or (inputs(214));
    layer0_outputs(2259) <= inputs(76);
    layer0_outputs(2260) <= not(inputs(181));
    layer0_outputs(2261) <= inputs(171);
    layer0_outputs(2262) <= not(inputs(106)) or (inputs(230));
    layer0_outputs(2263) <= (inputs(253)) and (inputs(18));
    layer0_outputs(2264) <= (inputs(238)) or (inputs(49));
    layer0_outputs(2265) <= not(inputs(145)) or (inputs(143));
    layer0_outputs(2266) <= not((inputs(17)) and (inputs(222)));
    layer0_outputs(2267) <= '1';
    layer0_outputs(2268) <= not((inputs(222)) and (inputs(107)));
    layer0_outputs(2269) <= not(inputs(212));
    layer0_outputs(2270) <= not((inputs(163)) xor (inputs(177)));
    layer0_outputs(2271) <= '1';
    layer0_outputs(2272) <= not(inputs(183));
    layer0_outputs(2273) <= '0';
    layer0_outputs(2274) <= not(inputs(7)) or (inputs(190));
    layer0_outputs(2275) <= (inputs(139)) and not (inputs(116));
    layer0_outputs(2276) <= (inputs(209)) and not (inputs(219));
    layer0_outputs(2277) <= not(inputs(31));
    layer0_outputs(2278) <= not(inputs(132)) or (inputs(48));
    layer0_outputs(2279) <= (inputs(223)) and (inputs(115));
    layer0_outputs(2280) <= (inputs(218)) and (inputs(229));
    layer0_outputs(2281) <= not(inputs(143)) or (inputs(251));
    layer0_outputs(2282) <= inputs(231);
    layer0_outputs(2283) <= (inputs(133)) and not (inputs(252));
    layer0_outputs(2284) <= not(inputs(176));
    layer0_outputs(2285) <= not(inputs(53));
    layer0_outputs(2286) <= not((inputs(230)) or (inputs(155)));
    layer0_outputs(2287) <= (inputs(34)) and (inputs(240));
    layer0_outputs(2288) <= not(inputs(206));
    layer0_outputs(2289) <= (inputs(91)) or (inputs(142));
    layer0_outputs(2290) <= (inputs(15)) xor (inputs(144));
    layer0_outputs(2291) <= (inputs(63)) and not (inputs(201));
    layer0_outputs(2292) <= not((inputs(113)) and (inputs(169)));
    layer0_outputs(2293) <= '0';
    layer0_outputs(2294) <= (inputs(165)) and not (inputs(243));
    layer0_outputs(2295) <= '1';
    layer0_outputs(2296) <= (inputs(4)) and not (inputs(49));
    layer0_outputs(2297) <= not(inputs(196));
    layer0_outputs(2298) <= (inputs(109)) or (inputs(188));
    layer0_outputs(2299) <= not(inputs(110));
    layer0_outputs(2300) <= not((inputs(72)) and (inputs(149)));
    layer0_outputs(2301) <= not(inputs(2));
    layer0_outputs(2302) <= (inputs(220)) or (inputs(97));
    layer0_outputs(2303) <= '1';
    layer0_outputs(2304) <= not((inputs(14)) or (inputs(174)));
    layer0_outputs(2305) <= not((inputs(87)) and (inputs(146)));
    layer0_outputs(2306) <= not((inputs(239)) or (inputs(131)));
    layer0_outputs(2307) <= not((inputs(247)) or (inputs(162)));
    layer0_outputs(2308) <= not(inputs(61));
    layer0_outputs(2309) <= not((inputs(84)) or (inputs(86)));
    layer0_outputs(2310) <= inputs(230);
    layer0_outputs(2311) <= '0';
    layer0_outputs(2312) <= not(inputs(130));
    layer0_outputs(2313) <= not(inputs(44)) or (inputs(239));
    layer0_outputs(2314) <= inputs(104);
    layer0_outputs(2315) <= (inputs(244)) xor (inputs(44));
    layer0_outputs(2316) <= inputs(243);
    layer0_outputs(2317) <= '0';
    layer0_outputs(2318) <= not(inputs(167));
    layer0_outputs(2319) <= (inputs(56)) and (inputs(21));
    layer0_outputs(2320) <= not(inputs(120)) or (inputs(161));
    layer0_outputs(2321) <= not((inputs(251)) and (inputs(22)));
    layer0_outputs(2322) <= (inputs(111)) or (inputs(210));
    layer0_outputs(2323) <= not((inputs(206)) or (inputs(18)));
    layer0_outputs(2324) <= (inputs(65)) and not (inputs(236));
    layer0_outputs(2325) <= not(inputs(229));
    layer0_outputs(2326) <= (inputs(90)) and not (inputs(116));
    layer0_outputs(2327) <= (inputs(160)) or (inputs(79));
    layer0_outputs(2328) <= not(inputs(125));
    layer0_outputs(2329) <= inputs(182);
    layer0_outputs(2330) <= inputs(207);
    layer0_outputs(2331) <= (inputs(83)) and (inputs(204));
    layer0_outputs(2332) <= not((inputs(7)) and (inputs(112)));
    layer0_outputs(2333) <= '1';
    layer0_outputs(2334) <= '1';
    layer0_outputs(2335) <= not(inputs(93));
    layer0_outputs(2336) <= inputs(85);
    layer0_outputs(2337) <= not(inputs(77));
    layer0_outputs(2338) <= not((inputs(115)) and (inputs(52)));
    layer0_outputs(2339) <= (inputs(254)) and (inputs(34));
    layer0_outputs(2340) <= '1';
    layer0_outputs(2341) <= '0';
    layer0_outputs(2342) <= not(inputs(248)) or (inputs(17));
    layer0_outputs(2343) <= not((inputs(134)) or (inputs(68)));
    layer0_outputs(2344) <= (inputs(43)) and (inputs(54));
    layer0_outputs(2345) <= (inputs(10)) and (inputs(7));
    layer0_outputs(2346) <= not(inputs(239));
    layer0_outputs(2347) <= inputs(149);
    layer0_outputs(2348) <= not((inputs(183)) and (inputs(94)));
    layer0_outputs(2349) <= '1';
    layer0_outputs(2350) <= '1';
    layer0_outputs(2351) <= not((inputs(192)) and (inputs(112)));
    layer0_outputs(2352) <= not((inputs(79)) or (inputs(1)));
    layer0_outputs(2353) <= (inputs(22)) and not (inputs(248));
    layer0_outputs(2354) <= (inputs(201)) and (inputs(178));
    layer0_outputs(2355) <= not(inputs(41)) or (inputs(68));
    layer0_outputs(2356) <= (inputs(53)) or (inputs(24));
    layer0_outputs(2357) <= not(inputs(168));
    layer0_outputs(2358) <= not((inputs(110)) or (inputs(219)));
    layer0_outputs(2359) <= '0';
    layer0_outputs(2360) <= inputs(113);
    layer0_outputs(2361) <= '0';
    layer0_outputs(2362) <= not(inputs(112));
    layer0_outputs(2363) <= inputs(72);
    layer0_outputs(2364) <= inputs(105);
    layer0_outputs(2365) <= not((inputs(174)) or (inputs(97)));
    layer0_outputs(2366) <= (inputs(189)) and not (inputs(17));
    layer0_outputs(2367) <= not(inputs(193));
    layer0_outputs(2368) <= '0';
    layer0_outputs(2369) <= inputs(43);
    layer0_outputs(2370) <= (inputs(227)) and not (inputs(233));
    layer0_outputs(2371) <= not(inputs(13)) or (inputs(243));
    layer0_outputs(2372) <= (inputs(50)) or (inputs(7));
    layer0_outputs(2373) <= '1';
    layer0_outputs(2374) <= (inputs(119)) and (inputs(192));
    layer0_outputs(2375) <= (inputs(8)) and not (inputs(98));
    layer0_outputs(2376) <= (inputs(107)) and not (inputs(153));
    layer0_outputs(2377) <= not(inputs(46));
    layer0_outputs(2378) <= inputs(139);
    layer0_outputs(2379) <= (inputs(158)) or (inputs(146));
    layer0_outputs(2380) <= not(inputs(156)) or (inputs(68));
    layer0_outputs(2381) <= (inputs(168)) and not (inputs(96));
    layer0_outputs(2382) <= inputs(196);
    layer0_outputs(2383) <= (inputs(74)) and (inputs(111));
    layer0_outputs(2384) <= (inputs(205)) or (inputs(24));
    layer0_outputs(2385) <= not(inputs(38));
    layer0_outputs(2386) <= '0';
    layer0_outputs(2387) <= '1';
    layer0_outputs(2388) <= not(inputs(159)) or (inputs(104));
    layer0_outputs(2389) <= inputs(99);
    layer0_outputs(2390) <= (inputs(26)) and not (inputs(4));
    layer0_outputs(2391) <= (inputs(100)) and not (inputs(2));
    layer0_outputs(2392) <= '0';
    layer0_outputs(2393) <= '1';
    layer0_outputs(2394) <= '1';
    layer0_outputs(2395) <= (inputs(100)) or (inputs(115));
    layer0_outputs(2396) <= inputs(170);
    layer0_outputs(2397) <= not(inputs(131)) or (inputs(40));
    layer0_outputs(2398) <= (inputs(119)) or (inputs(100));
    layer0_outputs(2399) <= not(inputs(12)) or (inputs(213));
    layer0_outputs(2400) <= not(inputs(148));
    layer0_outputs(2401) <= not((inputs(54)) or (inputs(20)));
    layer0_outputs(2402) <= not(inputs(42));
    layer0_outputs(2403) <= '1';
    layer0_outputs(2404) <= not((inputs(69)) or (inputs(101)));
    layer0_outputs(2405) <= (inputs(98)) and (inputs(172));
    layer0_outputs(2406) <= (inputs(64)) and not (inputs(217));
    layer0_outputs(2407) <= not(inputs(150)) or (inputs(92));
    layer0_outputs(2408) <= (inputs(232)) or (inputs(61));
    layer0_outputs(2409) <= not((inputs(233)) and (inputs(189)));
    layer0_outputs(2410) <= not(inputs(90));
    layer0_outputs(2411) <= not(inputs(156));
    layer0_outputs(2412) <= not((inputs(163)) or (inputs(100)));
    layer0_outputs(2413) <= not(inputs(167));
    layer0_outputs(2414) <= (inputs(2)) and (inputs(47));
    layer0_outputs(2415) <= (inputs(40)) or (inputs(79));
    layer0_outputs(2416) <= '0';
    layer0_outputs(2417) <= '1';
    layer0_outputs(2418) <= (inputs(79)) and not (inputs(147));
    layer0_outputs(2419) <= inputs(115);
    layer0_outputs(2420) <= '1';
    layer0_outputs(2421) <= (inputs(7)) and not (inputs(29));
    layer0_outputs(2422) <= not((inputs(221)) and (inputs(33)));
    layer0_outputs(2423) <= not(inputs(84)) or (inputs(32));
    layer0_outputs(2424) <= '1';
    layer0_outputs(2425) <= inputs(203);
    layer0_outputs(2426) <= '0';
    layer0_outputs(2427) <= '0';
    layer0_outputs(2428) <= not((inputs(150)) or (inputs(198)));
    layer0_outputs(2429) <= not(inputs(128));
    layer0_outputs(2430) <= '0';
    layer0_outputs(2431) <= not(inputs(162)) or (inputs(153));
    layer0_outputs(2432) <= not(inputs(226));
    layer0_outputs(2433) <= '1';
    layer0_outputs(2434) <= (inputs(159)) and (inputs(219));
    layer0_outputs(2435) <= (inputs(192)) or (inputs(146));
    layer0_outputs(2436) <= not((inputs(223)) or (inputs(38)));
    layer0_outputs(2437) <= not((inputs(62)) and (inputs(59)));
    layer0_outputs(2438) <= '1';
    layer0_outputs(2439) <= '0';
    layer0_outputs(2440) <= inputs(136);
    layer0_outputs(2441) <= not(inputs(74)) or (inputs(118));
    layer0_outputs(2442) <= inputs(136);
    layer0_outputs(2443) <= inputs(255);
    layer0_outputs(2444) <= not(inputs(211)) or (inputs(199));
    layer0_outputs(2445) <= not(inputs(88));
    layer0_outputs(2446) <= (inputs(139)) or (inputs(249));
    layer0_outputs(2447) <= not(inputs(110));
    layer0_outputs(2448) <= '0';
    layer0_outputs(2449) <= not(inputs(138));
    layer0_outputs(2450) <= inputs(217);
    layer0_outputs(2451) <= not(inputs(71));
    layer0_outputs(2452) <= not(inputs(97));
    layer0_outputs(2453) <= '0';
    layer0_outputs(2454) <= not((inputs(19)) and (inputs(87)));
    layer0_outputs(2455) <= '1';
    layer0_outputs(2456) <= not((inputs(211)) or (inputs(175)));
    layer0_outputs(2457) <= (inputs(238)) and (inputs(231));
    layer0_outputs(2458) <= not(inputs(21)) or (inputs(194));
    layer0_outputs(2459) <= not(inputs(5)) or (inputs(188));
    layer0_outputs(2460) <= '1';
    layer0_outputs(2461) <= not(inputs(121)) or (inputs(111));
    layer0_outputs(2462) <= inputs(226);
    layer0_outputs(2463) <= (inputs(180)) and (inputs(150));
    layer0_outputs(2464) <= '0';
    layer0_outputs(2465) <= not(inputs(152));
    layer0_outputs(2466) <= not((inputs(33)) xor (inputs(144)));
    layer0_outputs(2467) <= not(inputs(57));
    layer0_outputs(2468) <= (inputs(141)) or (inputs(144));
    layer0_outputs(2469) <= not((inputs(72)) and (inputs(48)));
    layer0_outputs(2470) <= not(inputs(228));
    layer0_outputs(2471) <= (inputs(29)) or (inputs(132));
    layer0_outputs(2472) <= '0';
    layer0_outputs(2473) <= (inputs(135)) and not (inputs(188));
    layer0_outputs(2474) <= '1';
    layer0_outputs(2475) <= not(inputs(74)) or (inputs(148));
    layer0_outputs(2476) <= (inputs(73)) and (inputs(37));
    layer0_outputs(2477) <= '1';
    layer0_outputs(2478) <= '0';
    layer0_outputs(2479) <= not((inputs(105)) and (inputs(226)));
    layer0_outputs(2480) <= '1';
    layer0_outputs(2481) <= inputs(232);
    layer0_outputs(2482) <= not(inputs(147));
    layer0_outputs(2483) <= '0';
    layer0_outputs(2484) <= not(inputs(176));
    layer0_outputs(2485) <= (inputs(102)) xor (inputs(132));
    layer0_outputs(2486) <= not((inputs(126)) and (inputs(20)));
    layer0_outputs(2487) <= (inputs(94)) and not (inputs(139));
    layer0_outputs(2488) <= not((inputs(38)) and (inputs(11)));
    layer0_outputs(2489) <= '0';
    layer0_outputs(2490) <= not((inputs(73)) and (inputs(248)));
    layer0_outputs(2491) <= (inputs(52)) and (inputs(112));
    layer0_outputs(2492) <= not(inputs(169)) or (inputs(157));
    layer0_outputs(2493) <= '0';
    layer0_outputs(2494) <= not((inputs(71)) and (inputs(45)));
    layer0_outputs(2495) <= (inputs(6)) and (inputs(238));
    layer0_outputs(2496) <= not(inputs(36));
    layer0_outputs(2497) <= '0';
    layer0_outputs(2498) <= not(inputs(108)) or (inputs(178));
    layer0_outputs(2499) <= '0';
    layer0_outputs(2500) <= inputs(25);
    layer0_outputs(2501) <= not(inputs(156)) or (inputs(206));
    layer0_outputs(2502) <= inputs(176);
    layer0_outputs(2503) <= not((inputs(126)) or (inputs(164)));
    layer0_outputs(2504) <= '0';
    layer0_outputs(2505) <= (inputs(28)) and not (inputs(102));
    layer0_outputs(2506) <= not(inputs(116)) or (inputs(5));
    layer0_outputs(2507) <= inputs(99);
    layer0_outputs(2508) <= (inputs(162)) or (inputs(219));
    layer0_outputs(2509) <= (inputs(51)) and not (inputs(108));
    layer0_outputs(2510) <= (inputs(45)) and not (inputs(16));
    layer0_outputs(2511) <= (inputs(160)) and not (inputs(10));
    layer0_outputs(2512) <= (inputs(45)) or (inputs(26));
    layer0_outputs(2513) <= inputs(123);
    layer0_outputs(2514) <= '1';
    layer0_outputs(2515) <= not(inputs(184)) or (inputs(172));
    layer0_outputs(2516) <= not((inputs(76)) or (inputs(60)));
    layer0_outputs(2517) <= not(inputs(100));
    layer0_outputs(2518) <= (inputs(195)) or (inputs(178));
    layer0_outputs(2519) <= '1';
    layer0_outputs(2520) <= (inputs(193)) and not (inputs(255));
    layer0_outputs(2521) <= (inputs(181)) and not (inputs(236));
    layer0_outputs(2522) <= (inputs(20)) or (inputs(247));
    layer0_outputs(2523) <= not((inputs(117)) xor (inputs(48)));
    layer0_outputs(2524) <= not((inputs(5)) or (inputs(156)));
    layer0_outputs(2525) <= not(inputs(42)) or (inputs(67));
    layer0_outputs(2526) <= (inputs(228)) and not (inputs(180));
    layer0_outputs(2527) <= inputs(99);
    layer0_outputs(2528) <= (inputs(39)) and not (inputs(118));
    layer0_outputs(2529) <= not((inputs(83)) and (inputs(25)));
    layer0_outputs(2530) <= inputs(85);
    layer0_outputs(2531) <= inputs(7);
    layer0_outputs(2532) <= '0';
    layer0_outputs(2533) <= not((inputs(236)) and (inputs(161)));
    layer0_outputs(2534) <= not((inputs(61)) or (inputs(123)));
    layer0_outputs(2535) <= (inputs(9)) and not (inputs(17));
    layer0_outputs(2536) <= (inputs(116)) xor (inputs(104));
    layer0_outputs(2537) <= (inputs(66)) xor (inputs(193));
    layer0_outputs(2538) <= not(inputs(205));
    layer0_outputs(2539) <= not(inputs(113)) or (inputs(74));
    layer0_outputs(2540) <= not(inputs(242)) or (inputs(89));
    layer0_outputs(2541) <= inputs(255);
    layer0_outputs(2542) <= not(inputs(13));
    layer0_outputs(2543) <= (inputs(47)) or (inputs(247));
    layer0_outputs(2544) <= not(inputs(21));
    layer0_outputs(2545) <= inputs(137);
    layer0_outputs(2546) <= '1';
    layer0_outputs(2547) <= inputs(156);
    layer0_outputs(2548) <= not((inputs(225)) or (inputs(189)));
    layer0_outputs(2549) <= not(inputs(27));
    layer0_outputs(2550) <= not((inputs(193)) or (inputs(148)));
    layer0_outputs(2551) <= not(inputs(36));
    layer0_outputs(2552) <= inputs(96);
    layer0_outputs(2553) <= (inputs(79)) and (inputs(12));
    layer0_outputs(2554) <= not((inputs(52)) or (inputs(115)));
    layer0_outputs(2555) <= '1';
    layer0_outputs(2556) <= '0';
    layer0_outputs(2557) <= not(inputs(60));
    layer0_outputs(2558) <= (inputs(41)) or (inputs(226));
    layer0_outputs(2559) <= (inputs(96)) and not (inputs(210));
    layer1_outputs(0) <= not(layer0_outputs(752));
    layer1_outputs(1) <= '1';
    layer1_outputs(2) <= not(layer0_outputs(559));
    layer1_outputs(3) <= (layer0_outputs(468)) and (layer0_outputs(123));
    layer1_outputs(4) <= '0';
    layer1_outputs(5) <= (layer0_outputs(1503)) and not (layer0_outputs(1867));
    layer1_outputs(6) <= layer0_outputs(1215);
    layer1_outputs(7) <= (layer0_outputs(1478)) and not (layer0_outputs(1111));
    layer1_outputs(8) <= layer0_outputs(426);
    layer1_outputs(9) <= '0';
    layer1_outputs(10) <= '0';
    layer1_outputs(11) <= '0';
    layer1_outputs(12) <= not(layer0_outputs(1236)) or (layer0_outputs(1791));
    layer1_outputs(13) <= layer0_outputs(1916);
    layer1_outputs(14) <= not(layer0_outputs(1007));
    layer1_outputs(15) <= not((layer0_outputs(1848)) or (layer0_outputs(1557)));
    layer1_outputs(16) <= not((layer0_outputs(2051)) and (layer0_outputs(1227)));
    layer1_outputs(17) <= not((layer0_outputs(816)) xor (layer0_outputs(194)));
    layer1_outputs(18) <= '1';
    layer1_outputs(19) <= not((layer0_outputs(2024)) or (layer0_outputs(1674)));
    layer1_outputs(20) <= layer0_outputs(1282);
    layer1_outputs(21) <= '1';
    layer1_outputs(22) <= '0';
    layer1_outputs(23) <= layer0_outputs(2447);
    layer1_outputs(24) <= '1';
    layer1_outputs(25) <= (layer0_outputs(2043)) and (layer0_outputs(291));
    layer1_outputs(26) <= layer0_outputs(1724);
    layer1_outputs(27) <= not((layer0_outputs(674)) or (layer0_outputs(1252)));
    layer1_outputs(28) <= not(layer0_outputs(898));
    layer1_outputs(29) <= not(layer0_outputs(1314)) or (layer0_outputs(854));
    layer1_outputs(30) <= not((layer0_outputs(514)) or (layer0_outputs(190)));
    layer1_outputs(31) <= not(layer0_outputs(2132));
    layer1_outputs(32) <= (layer0_outputs(683)) and (layer0_outputs(45));
    layer1_outputs(33) <= layer0_outputs(1352);
    layer1_outputs(34) <= '0';
    layer1_outputs(35) <= (layer0_outputs(489)) and not (layer0_outputs(1074));
    layer1_outputs(36) <= '1';
    layer1_outputs(37) <= not((layer0_outputs(294)) or (layer0_outputs(2218)));
    layer1_outputs(38) <= '1';
    layer1_outputs(39) <= not(layer0_outputs(951));
    layer1_outputs(40) <= not((layer0_outputs(2530)) and (layer0_outputs(926)));
    layer1_outputs(41) <= '0';
    layer1_outputs(42) <= layer0_outputs(165);
    layer1_outputs(43) <= layer0_outputs(505);
    layer1_outputs(44) <= not(layer0_outputs(1865)) or (layer0_outputs(1917));
    layer1_outputs(45) <= not(layer0_outputs(160));
    layer1_outputs(46) <= (layer0_outputs(1665)) and not (layer0_outputs(2058));
    layer1_outputs(47) <= not(layer0_outputs(188));
    layer1_outputs(48) <= not(layer0_outputs(1360));
    layer1_outputs(49) <= not((layer0_outputs(2530)) and (layer0_outputs(2481)));
    layer1_outputs(50) <= not(layer0_outputs(71));
    layer1_outputs(51) <= (layer0_outputs(1058)) and not (layer0_outputs(1083));
    layer1_outputs(52) <= not((layer0_outputs(2087)) or (layer0_outputs(2476)));
    layer1_outputs(53) <= (layer0_outputs(2503)) and (layer0_outputs(2070));
    layer1_outputs(54) <= '0';
    layer1_outputs(55) <= not(layer0_outputs(1561));
    layer1_outputs(56) <= layer0_outputs(851);
    layer1_outputs(57) <= (layer0_outputs(1211)) and not (layer0_outputs(1040));
    layer1_outputs(58) <= '1';
    layer1_outputs(59) <= not(layer0_outputs(1756));
    layer1_outputs(60) <= (layer0_outputs(628)) and not (layer0_outputs(954));
    layer1_outputs(61) <= not(layer0_outputs(661));
    layer1_outputs(62) <= not(layer0_outputs(2313));
    layer1_outputs(63) <= not(layer0_outputs(1127)) or (layer0_outputs(970));
    layer1_outputs(64) <= (layer0_outputs(1284)) and not (layer0_outputs(1886));
    layer1_outputs(65) <= not(layer0_outputs(1797)) or (layer0_outputs(1014));
    layer1_outputs(66) <= '1';
    layer1_outputs(67) <= layer0_outputs(1047);
    layer1_outputs(68) <= '1';
    layer1_outputs(69) <= not((layer0_outputs(2179)) or (layer0_outputs(1165)));
    layer1_outputs(70) <= (layer0_outputs(920)) or (layer0_outputs(21));
    layer1_outputs(71) <= not(layer0_outputs(621));
    layer1_outputs(72) <= '0';
    layer1_outputs(73) <= (layer0_outputs(1105)) and not (layer0_outputs(2264));
    layer1_outputs(74) <= (layer0_outputs(182)) and not (layer0_outputs(1996));
    layer1_outputs(75) <= (layer0_outputs(786)) and (layer0_outputs(1115));
    layer1_outputs(76) <= (layer0_outputs(511)) and not (layer0_outputs(1604));
    layer1_outputs(77) <= not((layer0_outputs(590)) and (layer0_outputs(1532)));
    layer1_outputs(78) <= (layer0_outputs(131)) or (layer0_outputs(347));
    layer1_outputs(79) <= not(layer0_outputs(2353)) or (layer0_outputs(1542));
    layer1_outputs(80) <= (layer0_outputs(1790)) and not (layer0_outputs(799));
    layer1_outputs(81) <= not(layer0_outputs(1949)) or (layer0_outputs(1631));
    layer1_outputs(82) <= '1';
    layer1_outputs(83) <= (layer0_outputs(2310)) and not (layer0_outputs(2243));
    layer1_outputs(84) <= not((layer0_outputs(847)) and (layer0_outputs(2392)));
    layer1_outputs(85) <= layer0_outputs(2428);
    layer1_outputs(86) <= not(layer0_outputs(2076)) or (layer0_outputs(512));
    layer1_outputs(87) <= not(layer0_outputs(1918));
    layer1_outputs(88) <= not(layer0_outputs(168));
    layer1_outputs(89) <= not((layer0_outputs(1849)) or (layer0_outputs(1814)));
    layer1_outputs(90) <= not(layer0_outputs(2404)) or (layer0_outputs(508));
    layer1_outputs(91) <= (layer0_outputs(882)) and not (layer0_outputs(1969));
    layer1_outputs(92) <= not(layer0_outputs(810));
    layer1_outputs(93) <= layer0_outputs(494);
    layer1_outputs(94) <= (layer0_outputs(2383)) and (layer0_outputs(2018));
    layer1_outputs(95) <= not(layer0_outputs(915));
    layer1_outputs(96) <= (layer0_outputs(1499)) and not (layer0_outputs(1430));
    layer1_outputs(97) <= (layer0_outputs(1800)) and (layer0_outputs(1479));
    layer1_outputs(98) <= layer0_outputs(2354);
    layer1_outputs(99) <= '1';
    layer1_outputs(100) <= '0';
    layer1_outputs(101) <= layer0_outputs(538);
    layer1_outputs(102) <= '0';
    layer1_outputs(103) <= (layer0_outputs(253)) and (layer0_outputs(1126));
    layer1_outputs(104) <= '0';
    layer1_outputs(105) <= (layer0_outputs(1691)) and (layer0_outputs(975));
    layer1_outputs(106) <= '0';
    layer1_outputs(107) <= (layer0_outputs(2033)) and not (layer0_outputs(1649));
    layer1_outputs(108) <= layer0_outputs(1963);
    layer1_outputs(109) <= '0';
    layer1_outputs(110) <= not(layer0_outputs(875)) or (layer0_outputs(1861));
    layer1_outputs(111) <= (layer0_outputs(1389)) and (layer0_outputs(1195));
    layer1_outputs(112) <= (layer0_outputs(1816)) or (layer0_outputs(1686));
    layer1_outputs(113) <= not(layer0_outputs(1938));
    layer1_outputs(114) <= '0';
    layer1_outputs(115) <= '1';
    layer1_outputs(116) <= not((layer0_outputs(1039)) and (layer0_outputs(2509)));
    layer1_outputs(117) <= not((layer0_outputs(2382)) or (layer0_outputs(304)));
    layer1_outputs(118) <= (layer0_outputs(2296)) and not (layer0_outputs(1271));
    layer1_outputs(119) <= layer0_outputs(266);
    layer1_outputs(120) <= (layer0_outputs(2341)) and (layer0_outputs(109));
    layer1_outputs(121) <= (layer0_outputs(633)) and not (layer0_outputs(630));
    layer1_outputs(122) <= layer0_outputs(1366);
    layer1_outputs(123) <= not(layer0_outputs(460)) or (layer0_outputs(336));
    layer1_outputs(124) <= not(layer0_outputs(610)) or (layer0_outputs(1197));
    layer1_outputs(125) <= not((layer0_outputs(245)) or (layer0_outputs(2168)));
    layer1_outputs(126) <= (layer0_outputs(142)) and not (layer0_outputs(2035));
    layer1_outputs(127) <= '1';
    layer1_outputs(128) <= (layer0_outputs(2449)) and not (layer0_outputs(1544));
    layer1_outputs(129) <= not(layer0_outputs(1849)) or (layer0_outputs(1583));
    layer1_outputs(130) <= (layer0_outputs(2054)) and not (layer0_outputs(1094));
    layer1_outputs(131) <= '0';
    layer1_outputs(132) <= '0';
    layer1_outputs(133) <= '1';
    layer1_outputs(134) <= (layer0_outputs(1382)) or (layer0_outputs(975));
    layer1_outputs(135) <= '1';
    layer1_outputs(136) <= not(layer0_outputs(184)) or (layer0_outputs(1734));
    layer1_outputs(137) <= not((layer0_outputs(1473)) and (layer0_outputs(1521)));
    layer1_outputs(138) <= (layer0_outputs(2284)) or (layer0_outputs(326));
    layer1_outputs(139) <= '0';
    layer1_outputs(140) <= layer0_outputs(829);
    layer1_outputs(141) <= not((layer0_outputs(2301)) and (layer0_outputs(2225)));
    layer1_outputs(142) <= not((layer0_outputs(820)) or (layer0_outputs(1031)));
    layer1_outputs(143) <= layer0_outputs(218);
    layer1_outputs(144) <= '1';
    layer1_outputs(145) <= layer0_outputs(1349);
    layer1_outputs(146) <= '0';
    layer1_outputs(147) <= layer0_outputs(2034);
    layer1_outputs(148) <= not(layer0_outputs(331)) or (layer0_outputs(701));
    layer1_outputs(149) <= not(layer0_outputs(1348)) or (layer0_outputs(2520));
    layer1_outputs(150) <= (layer0_outputs(605)) and not (layer0_outputs(220));
    layer1_outputs(151) <= '1';
    layer1_outputs(152) <= (layer0_outputs(959)) and not (layer0_outputs(2373));
    layer1_outputs(153) <= not(layer0_outputs(2225));
    layer1_outputs(154) <= '1';
    layer1_outputs(155) <= not(layer0_outputs(824));
    layer1_outputs(156) <= (layer0_outputs(2509)) and (layer0_outputs(2167));
    layer1_outputs(157) <= layer0_outputs(397);
    layer1_outputs(158) <= layer0_outputs(2148);
    layer1_outputs(159) <= not(layer0_outputs(1520));
    layer1_outputs(160) <= not(layer0_outputs(1296));
    layer1_outputs(161) <= not(layer0_outputs(808)) or (layer0_outputs(1735));
    layer1_outputs(162) <= layer0_outputs(104);
    layer1_outputs(163) <= (layer0_outputs(1515)) and not (layer0_outputs(966));
    layer1_outputs(164) <= '0';
    layer1_outputs(165) <= not(layer0_outputs(2226));
    layer1_outputs(166) <= layer0_outputs(2258);
    layer1_outputs(167) <= (layer0_outputs(1201)) or (layer0_outputs(2075));
    layer1_outputs(168) <= not((layer0_outputs(2384)) and (layer0_outputs(1400)));
    layer1_outputs(169) <= (layer0_outputs(1853)) xor (layer0_outputs(222));
    layer1_outputs(170) <= (layer0_outputs(1035)) and not (layer0_outputs(912));
    layer1_outputs(171) <= layer0_outputs(1017);
    layer1_outputs(172) <= not((layer0_outputs(1380)) or (layer0_outputs(1802)));
    layer1_outputs(173) <= not((layer0_outputs(440)) and (layer0_outputs(762)));
    layer1_outputs(174) <= not((layer0_outputs(1813)) and (layer0_outputs(2112)));
    layer1_outputs(175) <= not(layer0_outputs(2374)) or (layer0_outputs(631));
    layer1_outputs(176) <= not((layer0_outputs(1117)) or (layer0_outputs(791)));
    layer1_outputs(177) <= not((layer0_outputs(1405)) and (layer0_outputs(1973)));
    layer1_outputs(178) <= '0';
    layer1_outputs(179) <= '0';
    layer1_outputs(180) <= (layer0_outputs(1365)) or (layer0_outputs(386));
    layer1_outputs(181) <= (layer0_outputs(1208)) and (layer0_outputs(982));
    layer1_outputs(182) <= (layer0_outputs(1710)) and not (layer0_outputs(1436));
    layer1_outputs(183) <= (layer0_outputs(1323)) and not (layer0_outputs(1469));
    layer1_outputs(184) <= '1';
    layer1_outputs(185) <= (layer0_outputs(861)) or (layer0_outputs(2521));
    layer1_outputs(186) <= not(layer0_outputs(2459)) or (layer0_outputs(2104));
    layer1_outputs(187) <= layer0_outputs(1387);
    layer1_outputs(188) <= '0';
    layer1_outputs(189) <= layer0_outputs(1520);
    layer1_outputs(190) <= layer0_outputs(445);
    layer1_outputs(191) <= (layer0_outputs(2010)) or (layer0_outputs(810));
    layer1_outputs(192) <= '0';
    layer1_outputs(193) <= not((layer0_outputs(207)) and (layer0_outputs(130)));
    layer1_outputs(194) <= not(layer0_outputs(1269));
    layer1_outputs(195) <= (layer0_outputs(465)) and not (layer0_outputs(1621));
    layer1_outputs(196) <= layer0_outputs(1540);
    layer1_outputs(197) <= not(layer0_outputs(1277)) or (layer0_outputs(1612));
    layer1_outputs(198) <= (layer0_outputs(998)) and (layer0_outputs(1507));
    layer1_outputs(199) <= layer0_outputs(1945);
    layer1_outputs(200) <= not((layer0_outputs(1792)) or (layer0_outputs(2122)));
    layer1_outputs(201) <= '1';
    layer1_outputs(202) <= not(layer0_outputs(551));
    layer1_outputs(203) <= (layer0_outputs(1699)) and not (layer0_outputs(479));
    layer1_outputs(204) <= (layer0_outputs(2164)) and not (layer0_outputs(798));
    layer1_outputs(205) <= layer0_outputs(470);
    layer1_outputs(206) <= not(layer0_outputs(162));
    layer1_outputs(207) <= not((layer0_outputs(1179)) or (layer0_outputs(269)));
    layer1_outputs(208) <= not((layer0_outputs(722)) and (layer0_outputs(1981)));
    layer1_outputs(209) <= layer0_outputs(2236);
    layer1_outputs(210) <= (layer0_outputs(1490)) and (layer0_outputs(2114));
    layer1_outputs(211) <= '0';
    layer1_outputs(212) <= not(layer0_outputs(982));
    layer1_outputs(213) <= (layer0_outputs(1286)) and not (layer0_outputs(1140));
    layer1_outputs(214) <= (layer0_outputs(909)) xor (layer0_outputs(1766));
    layer1_outputs(215) <= not((layer0_outputs(285)) or (layer0_outputs(2507)));
    layer1_outputs(216) <= not(layer0_outputs(1508));
    layer1_outputs(217) <= (layer0_outputs(478)) and not (layer0_outputs(2153));
    layer1_outputs(218) <= not(layer0_outputs(1024)) or (layer0_outputs(552));
    layer1_outputs(219) <= not((layer0_outputs(1088)) or (layer0_outputs(1956)));
    layer1_outputs(220) <= (layer0_outputs(2180)) and not (layer0_outputs(13));
    layer1_outputs(221) <= '0';
    layer1_outputs(222) <= not(layer0_outputs(2471));
    layer1_outputs(223) <= not((layer0_outputs(608)) and (layer0_outputs(1694)));
    layer1_outputs(224) <= layer0_outputs(1974);
    layer1_outputs(225) <= '1';
    layer1_outputs(226) <= not(layer0_outputs(2319)) or (layer0_outputs(2407));
    layer1_outputs(227) <= not(layer0_outputs(2213));
    layer1_outputs(228) <= not(layer0_outputs(463));
    layer1_outputs(229) <= '0';
    layer1_outputs(230) <= '1';
    layer1_outputs(231) <= '1';
    layer1_outputs(232) <= not((layer0_outputs(2545)) or (layer0_outputs(1725)));
    layer1_outputs(233) <= not((layer0_outputs(173)) or (layer0_outputs(1511)));
    layer1_outputs(234) <= '1';
    layer1_outputs(235) <= not(layer0_outputs(1861)) or (layer0_outputs(653));
    layer1_outputs(236) <= not(layer0_outputs(312));
    layer1_outputs(237) <= '0';
    layer1_outputs(238) <= (layer0_outputs(2226)) and not (layer0_outputs(367));
    layer1_outputs(239) <= '1';
    layer1_outputs(240) <= not((layer0_outputs(95)) and (layer0_outputs(813)));
    layer1_outputs(241) <= not((layer0_outputs(15)) or (layer0_outputs(126)));
    layer1_outputs(242) <= not((layer0_outputs(1032)) or (layer0_outputs(1233)));
    layer1_outputs(243) <= '0';
    layer1_outputs(244) <= '0';
    layer1_outputs(245) <= not((layer0_outputs(557)) and (layer0_outputs(1970)));
    layer1_outputs(246) <= not(layer0_outputs(691));
    layer1_outputs(247) <= not(layer0_outputs(2055)) or (layer0_outputs(1804));
    layer1_outputs(248) <= (layer0_outputs(1739)) and not (layer0_outputs(187));
    layer1_outputs(249) <= not((layer0_outputs(1026)) or (layer0_outputs(2508)));
    layer1_outputs(250) <= (layer0_outputs(1950)) or (layer0_outputs(257));
    layer1_outputs(251) <= not(layer0_outputs(1150)) or (layer0_outputs(2388));
    layer1_outputs(252) <= '0';
    layer1_outputs(253) <= '0';
    layer1_outputs(254) <= not(layer0_outputs(1303)) or (layer0_outputs(2163));
    layer1_outputs(255) <= (layer0_outputs(1884)) and not (layer0_outputs(1304));
    layer1_outputs(256) <= not(layer0_outputs(2401));
    layer1_outputs(257) <= not(layer0_outputs(2398)) or (layer0_outputs(1659));
    layer1_outputs(258) <= (layer0_outputs(2003)) and not (layer0_outputs(2363));
    layer1_outputs(259) <= not(layer0_outputs(123));
    layer1_outputs(260) <= (layer0_outputs(1778)) and not (layer0_outputs(1549));
    layer1_outputs(261) <= '1';
    layer1_outputs(262) <= '1';
    layer1_outputs(263) <= (layer0_outputs(1803)) and (layer0_outputs(595));
    layer1_outputs(264) <= not(layer0_outputs(2256));
    layer1_outputs(265) <= not((layer0_outputs(831)) and (layer0_outputs(1198)));
    layer1_outputs(266) <= not((layer0_outputs(554)) or (layer0_outputs(1992)));
    layer1_outputs(267) <= not(layer0_outputs(332));
    layer1_outputs(268) <= '1';
    layer1_outputs(269) <= '0';
    layer1_outputs(270) <= layer0_outputs(973);
    layer1_outputs(271) <= (layer0_outputs(73)) and not (layer0_outputs(907));
    layer1_outputs(272) <= '1';
    layer1_outputs(273) <= not((layer0_outputs(769)) or (layer0_outputs(391)));
    layer1_outputs(274) <= '0';
    layer1_outputs(275) <= '0';
    layer1_outputs(276) <= '0';
    layer1_outputs(277) <= not(layer0_outputs(1133)) or (layer0_outputs(774));
    layer1_outputs(278) <= not(layer0_outputs(148)) or (layer0_outputs(224));
    layer1_outputs(279) <= (layer0_outputs(396)) or (layer0_outputs(671));
    layer1_outputs(280) <= '1';
    layer1_outputs(281) <= (layer0_outputs(2394)) and not (layer0_outputs(109));
    layer1_outputs(282) <= (layer0_outputs(1528)) and not (layer0_outputs(1807));
    layer1_outputs(283) <= (layer0_outputs(403)) and not (layer0_outputs(2017));
    layer1_outputs(284) <= '0';
    layer1_outputs(285) <= not(layer0_outputs(1342)) or (layer0_outputs(93));
    layer1_outputs(286) <= '1';
    layer1_outputs(287) <= layer0_outputs(1689);
    layer1_outputs(288) <= not(layer0_outputs(61)) or (layer0_outputs(883));
    layer1_outputs(289) <= not(layer0_outputs(2125)) or (layer0_outputs(609));
    layer1_outputs(290) <= not(layer0_outputs(1601));
    layer1_outputs(291) <= not((layer0_outputs(2551)) and (layer0_outputs(584)));
    layer1_outputs(292) <= '1';
    layer1_outputs(293) <= (layer0_outputs(1423)) and (layer0_outputs(1328));
    layer1_outputs(294) <= (layer0_outputs(1986)) or (layer0_outputs(380));
    layer1_outputs(295) <= (layer0_outputs(2306)) and (layer0_outputs(1529));
    layer1_outputs(296) <= not(layer0_outputs(2360)) or (layer0_outputs(2479));
    layer1_outputs(297) <= not(layer0_outputs(501));
    layer1_outputs(298) <= layer0_outputs(843);
    layer1_outputs(299) <= layer0_outputs(1716);
    layer1_outputs(300) <= (layer0_outputs(1005)) and not (layer0_outputs(695));
    layer1_outputs(301) <= '1';
    layer1_outputs(302) <= not(layer0_outputs(1556));
    layer1_outputs(303) <= (layer0_outputs(1646)) and not (layer0_outputs(861));
    layer1_outputs(304) <= (layer0_outputs(758)) and not (layer0_outputs(1823));
    layer1_outputs(305) <= (layer0_outputs(1016)) or (layer0_outputs(1282));
    layer1_outputs(306) <= '1';
    layer1_outputs(307) <= '0';
    layer1_outputs(308) <= layer0_outputs(108);
    layer1_outputs(309) <= not(layer0_outputs(2557)) or (layer0_outputs(224));
    layer1_outputs(310) <= '0';
    layer1_outputs(311) <= not(layer0_outputs(610));
    layer1_outputs(312) <= '0';
    layer1_outputs(313) <= (layer0_outputs(186)) and not (layer0_outputs(2166));
    layer1_outputs(314) <= not((layer0_outputs(258)) and (layer0_outputs(2114)));
    layer1_outputs(315) <= '1';
    layer1_outputs(316) <= layer0_outputs(2544);
    layer1_outputs(317) <= not(layer0_outputs(1802)) or (layer0_outputs(733));
    layer1_outputs(318) <= not(layer0_outputs(879));
    layer1_outputs(319) <= not(layer0_outputs(2032)) or (layer0_outputs(54));
    layer1_outputs(320) <= '1';
    layer1_outputs(321) <= layer0_outputs(1376);
    layer1_outputs(322) <= not(layer0_outputs(951));
    layer1_outputs(323) <= not(layer0_outputs(1364));
    layer1_outputs(324) <= not((layer0_outputs(418)) or (layer0_outputs(369)));
    layer1_outputs(325) <= not(layer0_outputs(1099)) or (layer0_outputs(1793));
    layer1_outputs(326) <= (layer0_outputs(98)) and not (layer0_outputs(2269));
    layer1_outputs(327) <= (layer0_outputs(575)) and (layer0_outputs(445));
    layer1_outputs(328) <= '1';
    layer1_outputs(329) <= (layer0_outputs(2457)) and not (layer0_outputs(244));
    layer1_outputs(330) <= '1';
    layer1_outputs(331) <= not(layer0_outputs(1881));
    layer1_outputs(332) <= layer0_outputs(1184);
    layer1_outputs(333) <= not((layer0_outputs(1160)) or (layer0_outputs(483)));
    layer1_outputs(334) <= '1';
    layer1_outputs(335) <= not(layer0_outputs(825)) or (layer0_outputs(2516));
    layer1_outputs(336) <= not(layer0_outputs(2002));
    layer1_outputs(337) <= not(layer0_outputs(757));
    layer1_outputs(338) <= not((layer0_outputs(1418)) and (layer0_outputs(1292)));
    layer1_outputs(339) <= not(layer0_outputs(1907)) or (layer0_outputs(296));
    layer1_outputs(340) <= (layer0_outputs(482)) and (layer0_outputs(636));
    layer1_outputs(341) <= '0';
    layer1_outputs(342) <= not(layer0_outputs(2408)) or (layer0_outputs(2270));
    layer1_outputs(343) <= layer0_outputs(489);
    layer1_outputs(344) <= '0';
    layer1_outputs(345) <= (layer0_outputs(115)) and not (layer0_outputs(2220));
    layer1_outputs(346) <= (layer0_outputs(2542)) and not (layer0_outputs(1408));
    layer1_outputs(347) <= '0';
    layer1_outputs(348) <= '1';
    layer1_outputs(349) <= (layer0_outputs(919)) and not (layer0_outputs(591));
    layer1_outputs(350) <= not((layer0_outputs(2501)) and (layer0_outputs(502)));
    layer1_outputs(351) <= '0';
    layer1_outputs(352) <= not((layer0_outputs(1153)) or (layer0_outputs(780)));
    layer1_outputs(353) <= layer0_outputs(2288);
    layer1_outputs(354) <= '0';
    layer1_outputs(355) <= layer0_outputs(1727);
    layer1_outputs(356) <= not(layer0_outputs(497));
    layer1_outputs(357) <= layer0_outputs(601);
    layer1_outputs(358) <= '1';
    layer1_outputs(359) <= '1';
    layer1_outputs(360) <= (layer0_outputs(383)) and (layer0_outputs(1799));
    layer1_outputs(361) <= layer0_outputs(932);
    layer1_outputs(362) <= '0';
    layer1_outputs(363) <= '1';
    layer1_outputs(364) <= not((layer0_outputs(542)) and (layer0_outputs(1746)));
    layer1_outputs(365) <= not((layer0_outputs(733)) and (layer0_outputs(341)));
    layer1_outputs(366) <= not(layer0_outputs(313)) or (layer0_outputs(2490));
    layer1_outputs(367) <= '1';
    layer1_outputs(368) <= not(layer0_outputs(1789));
    layer1_outputs(369) <= not(layer0_outputs(572));
    layer1_outputs(370) <= (layer0_outputs(2487)) and not (layer0_outputs(701));
    layer1_outputs(371) <= (layer0_outputs(225)) and not (layer0_outputs(181));
    layer1_outputs(372) <= not(layer0_outputs(787));
    layer1_outputs(373) <= '0';
    layer1_outputs(374) <= '0';
    layer1_outputs(375) <= (layer0_outputs(2063)) and not (layer0_outputs(949));
    layer1_outputs(376) <= (layer0_outputs(1051)) or (layer0_outputs(2543));
    layer1_outputs(377) <= layer0_outputs(2544);
    layer1_outputs(378) <= '1';
    layer1_outputs(379) <= not(layer0_outputs(929));
    layer1_outputs(380) <= not(layer0_outputs(843));
    layer1_outputs(381) <= not(layer0_outputs(1817));
    layer1_outputs(382) <= layer0_outputs(1447);
    layer1_outputs(383) <= not((layer0_outputs(375)) or (layer0_outputs(2223)));
    layer1_outputs(384) <= '0';
    layer1_outputs(385) <= not(layer0_outputs(1157)) or (layer0_outputs(2251));
    layer1_outputs(386) <= layer0_outputs(340);
    layer1_outputs(387) <= (layer0_outputs(1638)) and not (layer0_outputs(1760));
    layer1_outputs(388) <= not((layer0_outputs(1151)) or (layer0_outputs(2402)));
    layer1_outputs(389) <= layer0_outputs(1706);
    layer1_outputs(390) <= not(layer0_outputs(798)) or (layer0_outputs(159));
    layer1_outputs(391) <= (layer0_outputs(2441)) and not (layer0_outputs(1358));
    layer1_outputs(392) <= (layer0_outputs(1775)) or (layer0_outputs(1074));
    layer1_outputs(393) <= not(layer0_outputs(2458)) or (layer0_outputs(1187));
    layer1_outputs(394) <= '0';
    layer1_outputs(395) <= not((layer0_outputs(1468)) and (layer0_outputs(1225)));
    layer1_outputs(396) <= (layer0_outputs(49)) xor (layer0_outputs(383));
    layer1_outputs(397) <= (layer0_outputs(166)) and not (layer0_outputs(2355));
    layer1_outputs(398) <= not(layer0_outputs(311)) or (layer0_outputs(2457));
    layer1_outputs(399) <= not((layer0_outputs(1241)) or (layer0_outputs(1585)));
    layer1_outputs(400) <= (layer0_outputs(2525)) and not (layer0_outputs(74));
    layer1_outputs(401) <= (layer0_outputs(323)) and not (layer0_outputs(2306));
    layer1_outputs(402) <= (layer0_outputs(1968)) and (layer0_outputs(1806));
    layer1_outputs(403) <= (layer0_outputs(1964)) and not (layer0_outputs(815));
    layer1_outputs(404) <= not((layer0_outputs(727)) or (layer0_outputs(1473)));
    layer1_outputs(405) <= layer0_outputs(878);
    layer1_outputs(406) <= (layer0_outputs(2224)) or (layer0_outputs(940));
    layer1_outputs(407) <= not((layer0_outputs(1523)) or (layer0_outputs(2099)));
    layer1_outputs(408) <= '0';
    layer1_outputs(409) <= not(layer0_outputs(748));
    layer1_outputs(410) <= '0';
    layer1_outputs(411) <= not((layer0_outputs(850)) or (layer0_outputs(2093)));
    layer1_outputs(412) <= (layer0_outputs(58)) and (layer0_outputs(2520));
    layer1_outputs(413) <= (layer0_outputs(1886)) and not (layer0_outputs(363));
    layer1_outputs(414) <= '0';
    layer1_outputs(415) <= '1';
    layer1_outputs(416) <= '1';
    layer1_outputs(417) <= not((layer0_outputs(1440)) or (layer0_outputs(776)));
    layer1_outputs(418) <= not(layer0_outputs(1145));
    layer1_outputs(419) <= not(layer0_outputs(2378));
    layer1_outputs(420) <= not((layer0_outputs(1428)) or (layer0_outputs(819)));
    layer1_outputs(421) <= not(layer0_outputs(1110));
    layer1_outputs(422) <= not(layer0_outputs(2367)) or (layer0_outputs(1362));
    layer1_outputs(423) <= (layer0_outputs(1249)) and not (layer0_outputs(1681));
    layer1_outputs(424) <= layer0_outputs(1930);
    layer1_outputs(425) <= not((layer0_outputs(2052)) and (layer0_outputs(1787)));
    layer1_outputs(426) <= not((layer0_outputs(1052)) or (layer0_outputs(1702)));
    layer1_outputs(427) <= '0';
    layer1_outputs(428) <= layer0_outputs(2214);
    layer1_outputs(429) <= not(layer0_outputs(295)) or (layer0_outputs(2094));
    layer1_outputs(430) <= not(layer0_outputs(921)) or (layer0_outputs(692));
    layer1_outputs(431) <= not(layer0_outputs(1967));
    layer1_outputs(432) <= not((layer0_outputs(2129)) and (layer0_outputs(599)));
    layer1_outputs(433) <= (layer0_outputs(66)) and not (layer0_outputs(897));
    layer1_outputs(434) <= (layer0_outputs(373)) and not (layer0_outputs(1900));
    layer1_outputs(435) <= not((layer0_outputs(1810)) xor (layer0_outputs(1156)));
    layer1_outputs(436) <= (layer0_outputs(1426)) and not (layer0_outputs(1214));
    layer1_outputs(437) <= not(layer0_outputs(300)) or (layer0_outputs(441));
    layer1_outputs(438) <= layer0_outputs(1805);
    layer1_outputs(439) <= (layer0_outputs(2080)) and not (layer0_outputs(1469));
    layer1_outputs(440) <= not(layer0_outputs(1920)) or (layer0_outputs(1991));
    layer1_outputs(441) <= not(layer0_outputs(2021));
    layer1_outputs(442) <= not((layer0_outputs(1216)) or (layer0_outputs(1209)));
    layer1_outputs(443) <= layer0_outputs(1873);
    layer1_outputs(444) <= '1';
    layer1_outputs(445) <= not(layer0_outputs(238));
    layer1_outputs(446) <= not(layer0_outputs(1410));
    layer1_outputs(447) <= '1';
    layer1_outputs(448) <= not((layer0_outputs(1081)) or (layer0_outputs(2552)));
    layer1_outputs(449) <= layer0_outputs(1590);
    layer1_outputs(450) <= '1';
    layer1_outputs(451) <= '0';
    layer1_outputs(452) <= not(layer0_outputs(1995)) or (layer0_outputs(2302));
    layer1_outputs(453) <= (layer0_outputs(87)) and not (layer0_outputs(2173));
    layer1_outputs(454) <= layer0_outputs(1427);
    layer1_outputs(455) <= not(layer0_outputs(1368)) or (layer0_outputs(180));
    layer1_outputs(456) <= layer0_outputs(2423);
    layer1_outputs(457) <= '0';
    layer1_outputs(458) <= not(layer0_outputs(2186)) or (layer0_outputs(785));
    layer1_outputs(459) <= layer0_outputs(1983);
    layer1_outputs(460) <= (layer0_outputs(315)) or (layer0_outputs(2280));
    layer1_outputs(461) <= not((layer0_outputs(845)) or (layer0_outputs(486)));
    layer1_outputs(462) <= layer0_outputs(200);
    layer1_outputs(463) <= layer0_outputs(1045);
    layer1_outputs(464) <= '1';
    layer1_outputs(465) <= not((layer0_outputs(1641)) or (layer0_outputs(2413)));
    layer1_outputs(466) <= not((layer0_outputs(1909)) and (layer0_outputs(1297)));
    layer1_outputs(467) <= '1';
    layer1_outputs(468) <= not((layer0_outputs(65)) xor (layer0_outputs(2379)));
    layer1_outputs(469) <= layer0_outputs(2429);
    layer1_outputs(470) <= layer0_outputs(44);
    layer1_outputs(471) <= layer0_outputs(1134);
    layer1_outputs(472) <= (layer0_outputs(960)) and not (layer0_outputs(2339));
    layer1_outputs(473) <= '0';
    layer1_outputs(474) <= layer0_outputs(1256);
    layer1_outputs(475) <= (layer0_outputs(1415)) and (layer0_outputs(1970));
    layer1_outputs(476) <= not(layer0_outputs(668)) or (layer0_outputs(1396));
    layer1_outputs(477) <= (layer0_outputs(76)) and not (layer0_outputs(761));
    layer1_outputs(478) <= not((layer0_outputs(832)) or (layer0_outputs(1936)));
    layer1_outputs(479) <= '0';
    layer1_outputs(480) <= not(layer0_outputs(1351));
    layer1_outputs(481) <= (layer0_outputs(1324)) and not (layer0_outputs(1453));
    layer1_outputs(482) <= (layer0_outputs(18)) or (layer0_outputs(1671));
    layer1_outputs(483) <= not(layer0_outputs(2559)) or (layer0_outputs(1429));
    layer1_outputs(484) <= (layer0_outputs(1248)) or (layer0_outputs(1553));
    layer1_outputs(485) <= (layer0_outputs(1634)) or (layer0_outputs(1036));
    layer1_outputs(486) <= (layer0_outputs(284)) and (layer0_outputs(1196));
    layer1_outputs(487) <= not(layer0_outputs(1706));
    layer1_outputs(488) <= not((layer0_outputs(2157)) and (layer0_outputs(2385)));
    layer1_outputs(489) <= layer0_outputs(292);
    layer1_outputs(490) <= not(layer0_outputs(1070));
    layer1_outputs(491) <= layer0_outputs(1801);
    layer1_outputs(492) <= not((layer0_outputs(373)) and (layer0_outputs(862)));
    layer1_outputs(493) <= layer0_outputs(2364);
    layer1_outputs(494) <= layer0_outputs(2309);
    layer1_outputs(495) <= layer0_outputs(1156);
    layer1_outputs(496) <= layer0_outputs(2065);
    layer1_outputs(497) <= (layer0_outputs(366)) or (layer0_outputs(2334));
    layer1_outputs(498) <= '0';
    layer1_outputs(499) <= not(layer0_outputs(1227)) or (layer0_outputs(1867));
    layer1_outputs(500) <= layer0_outputs(204);
    layer1_outputs(501) <= not((layer0_outputs(1221)) xor (layer0_outputs(266)));
    layer1_outputs(502) <= '1';
    layer1_outputs(503) <= '0';
    layer1_outputs(504) <= not(layer0_outputs(736));
    layer1_outputs(505) <= not(layer0_outputs(2079)) or (layer0_outputs(641));
    layer1_outputs(506) <= not((layer0_outputs(2527)) or (layer0_outputs(477)));
    layer1_outputs(507) <= not(layer0_outputs(598)) or (layer0_outputs(168));
    layer1_outputs(508) <= not((layer0_outputs(1580)) or (layer0_outputs(2074)));
    layer1_outputs(509) <= not(layer0_outputs(1567)) or (layer0_outputs(1650));
    layer1_outputs(510) <= '1';
    layer1_outputs(511) <= not((layer0_outputs(2052)) or (layer0_outputs(225)));
    layer1_outputs(512) <= not((layer0_outputs(1458)) and (layer0_outputs(2329)));
    layer1_outputs(513) <= not(layer0_outputs(2282));
    layer1_outputs(514) <= not(layer0_outputs(1081)) or (layer0_outputs(41));
    layer1_outputs(515) <= layer0_outputs(1528);
    layer1_outputs(516) <= not((layer0_outputs(319)) or (layer0_outputs(858)));
    layer1_outputs(517) <= (layer0_outputs(1569)) and not (layer0_outputs(73));
    layer1_outputs(518) <= not((layer0_outputs(845)) and (layer0_outputs(1023)));
    layer1_outputs(519) <= (layer0_outputs(318)) and not (layer0_outputs(1838));
    layer1_outputs(520) <= not((layer0_outputs(2055)) or (layer0_outputs(801)));
    layer1_outputs(521) <= '0';
    layer1_outputs(522) <= '0';
    layer1_outputs(523) <= (layer0_outputs(11)) and (layer0_outputs(2465));
    layer1_outputs(524) <= (layer0_outputs(1092)) and not (layer0_outputs(1118));
    layer1_outputs(525) <= (layer0_outputs(426)) or (layer0_outputs(2412));
    layer1_outputs(526) <= not(layer0_outputs(1568));
    layer1_outputs(527) <= (layer0_outputs(1855)) and (layer0_outputs(1244));
    layer1_outputs(528) <= not(layer0_outputs(1194));
    layer1_outputs(529) <= (layer0_outputs(848)) and (layer0_outputs(2310));
    layer1_outputs(530) <= not(layer0_outputs(288)) or (layer0_outputs(1664));
    layer1_outputs(531) <= '0';
    layer1_outputs(532) <= layer0_outputs(869);
    layer1_outputs(533) <= not(layer0_outputs(57)) or (layer0_outputs(171));
    layer1_outputs(534) <= not((layer0_outputs(1389)) and (layer0_outputs(2138)));
    layer1_outputs(535) <= layer0_outputs(272);
    layer1_outputs(536) <= (layer0_outputs(1666)) or (layer0_outputs(1898));
    layer1_outputs(537) <= not(layer0_outputs(1525));
    layer1_outputs(538) <= not((layer0_outputs(697)) or (layer0_outputs(233)));
    layer1_outputs(539) <= (layer0_outputs(1491)) and not (layer0_outputs(1837));
    layer1_outputs(540) <= not((layer0_outputs(252)) or (layer0_outputs(796)));
    layer1_outputs(541) <= not((layer0_outputs(2141)) or (layer0_outputs(2208)));
    layer1_outputs(542) <= (layer0_outputs(1262)) and not (layer0_outputs(2491));
    layer1_outputs(543) <= layer0_outputs(68);
    layer1_outputs(544) <= '0';
    layer1_outputs(545) <= (layer0_outputs(936)) and not (layer0_outputs(2040));
    layer1_outputs(546) <= layer0_outputs(644);
    layer1_outputs(547) <= (layer0_outputs(1870)) and not (layer0_outputs(783));
    layer1_outputs(548) <= '1';
    layer1_outputs(549) <= not(layer0_outputs(2128));
    layer1_outputs(550) <= not(layer0_outputs(2262));
    layer1_outputs(551) <= layer0_outputs(465);
    layer1_outputs(552) <= (layer0_outputs(2175)) xor (layer0_outputs(934));
    layer1_outputs(553) <= '1';
    layer1_outputs(554) <= not(layer0_outputs(1677));
    layer1_outputs(555) <= not(layer0_outputs(1529));
    layer1_outputs(556) <= not((layer0_outputs(721)) xor (layer0_outputs(16)));
    layer1_outputs(557) <= layer0_outputs(2518);
    layer1_outputs(558) <= not(layer0_outputs(335));
    layer1_outputs(559) <= '0';
    layer1_outputs(560) <= '1';
    layer1_outputs(561) <= layer0_outputs(1668);
    layer1_outputs(562) <= '0';
    layer1_outputs(563) <= (layer0_outputs(746)) and not (layer0_outputs(1135));
    layer1_outputs(564) <= '1';
    layer1_outputs(565) <= (layer0_outputs(740)) and not (layer0_outputs(523));
    layer1_outputs(566) <= (layer0_outputs(1953)) or (layer0_outputs(1267));
    layer1_outputs(567) <= not((layer0_outputs(1238)) or (layer0_outputs(1088)));
    layer1_outputs(568) <= (layer0_outputs(834)) or (layer0_outputs(1747));
    layer1_outputs(569) <= '1';
    layer1_outputs(570) <= not((layer0_outputs(192)) or (layer0_outputs(1783)));
    layer1_outputs(571) <= layer0_outputs(983);
    layer1_outputs(572) <= not(layer0_outputs(549)) or (layer0_outputs(1501));
    layer1_outputs(573) <= not(layer0_outputs(921)) or (layer0_outputs(128));
    layer1_outputs(574) <= '0';
    layer1_outputs(575) <= not(layer0_outputs(2117));
    layer1_outputs(576) <= not(layer0_outputs(1749)) or (layer0_outputs(119));
    layer1_outputs(577) <= not((layer0_outputs(1689)) or (layer0_outputs(1205)));
    layer1_outputs(578) <= '1';
    layer1_outputs(579) <= '0';
    layer1_outputs(580) <= (layer0_outputs(1922)) or (layer0_outputs(665));
    layer1_outputs(581) <= not(layer0_outputs(778));
    layer1_outputs(582) <= not(layer0_outputs(888));
    layer1_outputs(583) <= (layer0_outputs(1075)) and not (layer0_outputs(729));
    layer1_outputs(584) <= not(layer0_outputs(528)) or (layer0_outputs(1645));
    layer1_outputs(585) <= not(layer0_outputs(817)) or (layer0_outputs(2053));
    layer1_outputs(586) <= not(layer0_outputs(1101)) or (layer0_outputs(574));
    layer1_outputs(587) <= '1';
    layer1_outputs(588) <= not((layer0_outputs(2025)) or (layer0_outputs(1172)));
    layer1_outputs(589) <= not(layer0_outputs(937));
    layer1_outputs(590) <= not((layer0_outputs(1625)) xor (layer0_outputs(992)));
    layer1_outputs(591) <= not(layer0_outputs(1284));
    layer1_outputs(592) <= (layer0_outputs(1463)) and not (layer0_outputs(1142));
    layer1_outputs(593) <= not(layer0_outputs(1180));
    layer1_outputs(594) <= not(layer0_outputs(326));
    layer1_outputs(595) <= not(layer0_outputs(2082)) or (layer0_outputs(1598));
    layer1_outputs(596) <= not(layer0_outputs(1944));
    layer1_outputs(597) <= not(layer0_outputs(231));
    layer1_outputs(598) <= (layer0_outputs(906)) and (layer0_outputs(1933));
    layer1_outputs(599) <= (layer0_outputs(1301)) or (layer0_outputs(616));
    layer1_outputs(600) <= (layer0_outputs(237)) and (layer0_outputs(371));
    layer1_outputs(601) <= not(layer0_outputs(2061));
    layer1_outputs(602) <= not(layer0_outputs(585)) or (layer0_outputs(1316));
    layer1_outputs(603) <= not(layer0_outputs(2339)) or (layer0_outputs(1852));
    layer1_outputs(604) <= layer0_outputs(2203);
    layer1_outputs(605) <= '0';
    layer1_outputs(606) <= layer0_outputs(750);
    layer1_outputs(607) <= '0';
    layer1_outputs(608) <= (layer0_outputs(1154)) and not (layer0_outputs(787));
    layer1_outputs(609) <= (layer0_outputs(1191)) or (layer0_outputs(90));
    layer1_outputs(610) <= not(layer0_outputs(2020)) or (layer0_outputs(170));
    layer1_outputs(611) <= not((layer0_outputs(1485)) and (layer0_outputs(1855)));
    layer1_outputs(612) <= (layer0_outputs(1977)) or (layer0_outputs(150));
    layer1_outputs(613) <= layer0_outputs(1687);
    layer1_outputs(614) <= not(layer0_outputs(574)) or (layer0_outputs(541));
    layer1_outputs(615) <= '1';
    layer1_outputs(616) <= '1';
    layer1_outputs(617) <= '1';
    layer1_outputs(618) <= '0';
    layer1_outputs(619) <= not(layer0_outputs(1623));
    layer1_outputs(620) <= layer0_outputs(677);
    layer1_outputs(621) <= not(layer0_outputs(2496));
    layer1_outputs(622) <= not(layer0_outputs(2335));
    layer1_outputs(623) <= '1';
    layer1_outputs(624) <= not((layer0_outputs(2469)) or (layer0_outputs(1737)));
    layer1_outputs(625) <= (layer0_outputs(112)) and (layer0_outputs(2276));
    layer1_outputs(626) <= (layer0_outputs(2440)) and not (layer0_outputs(690));
    layer1_outputs(627) <= (layer0_outputs(2340)) and (layer0_outputs(2344));
    layer1_outputs(628) <= (layer0_outputs(2314)) and (layer0_outputs(935));
    layer1_outputs(629) <= '1';
    layer1_outputs(630) <= not(layer0_outputs(2131)) or (layer0_outputs(550));
    layer1_outputs(631) <= not(layer0_outputs(425));
    layer1_outputs(632) <= (layer0_outputs(2303)) or (layer0_outputs(2295));
    layer1_outputs(633) <= (layer0_outputs(1290)) and (layer0_outputs(2248));
    layer1_outputs(634) <= not((layer0_outputs(1574)) or (layer0_outputs(404)));
    layer1_outputs(635) <= layer0_outputs(2486);
    layer1_outputs(636) <= (layer0_outputs(2064)) or (layer0_outputs(655));
    layer1_outputs(637) <= not(layer0_outputs(1301)) or (layer0_outputs(867));
    layer1_outputs(638) <= not(layer0_outputs(273));
    layer1_outputs(639) <= not(layer0_outputs(803));
    layer1_outputs(640) <= '0';
    layer1_outputs(641) <= not(layer0_outputs(2183));
    layer1_outputs(642) <= '1';
    layer1_outputs(643) <= not(layer0_outputs(2329));
    layer1_outputs(644) <= layer0_outputs(584);
    layer1_outputs(645) <= layer0_outputs(2216);
    layer1_outputs(646) <= (layer0_outputs(1462)) and not (layer0_outputs(349));
    layer1_outputs(647) <= '1';
    layer1_outputs(648) <= (layer0_outputs(318)) and not (layer0_outputs(1339));
    layer1_outputs(649) <= (layer0_outputs(1797)) or (layer0_outputs(190));
    layer1_outputs(650) <= not(layer0_outputs(1561));
    layer1_outputs(651) <= not(layer0_outputs(361)) or (layer0_outputs(637));
    layer1_outputs(652) <= layer0_outputs(840);
    layer1_outputs(653) <= layer0_outputs(136);
    layer1_outputs(654) <= not((layer0_outputs(593)) xor (layer0_outputs(1434)));
    layer1_outputs(655) <= '0';
    layer1_outputs(656) <= not(layer0_outputs(2169)) or (layer0_outputs(2185));
    layer1_outputs(657) <= (layer0_outputs(1452)) and not (layer0_outputs(735));
    layer1_outputs(658) <= (layer0_outputs(177)) and not (layer0_outputs(2442));
    layer1_outputs(659) <= '1';
    layer1_outputs(660) <= '1';
    layer1_outputs(661) <= '0';
    layer1_outputs(662) <= not(layer0_outputs(1758));
    layer1_outputs(663) <= (layer0_outputs(2377)) xor (layer0_outputs(1381));
    layer1_outputs(664) <= not(layer0_outputs(197)) or (layer0_outputs(749));
    layer1_outputs(665) <= (layer0_outputs(1699)) and not (layer0_outputs(1291));
    layer1_outputs(666) <= not(layer0_outputs(2274)) or (layer0_outputs(1251));
    layer1_outputs(667) <= layer0_outputs(827);
    layer1_outputs(668) <= not((layer0_outputs(96)) and (layer0_outputs(348)));
    layer1_outputs(669) <= (layer0_outputs(1700)) and not (layer0_outputs(720));
    layer1_outputs(670) <= (layer0_outputs(2482)) and (layer0_outputs(462));
    layer1_outputs(671) <= (layer0_outputs(49)) xor (layer0_outputs(1635));
    layer1_outputs(672) <= not(layer0_outputs(2247)) or (layer0_outputs(635));
    layer1_outputs(673) <= not(layer0_outputs(2266)) or (layer0_outputs(113));
    layer1_outputs(674) <= (layer0_outputs(937)) and not (layer0_outputs(1288));
    layer1_outputs(675) <= not(layer0_outputs(1972)) or (layer0_outputs(208));
    layer1_outputs(676) <= not((layer0_outputs(2348)) xor (layer0_outputs(467)));
    layer1_outputs(677) <= '0';
    layer1_outputs(678) <= not((layer0_outputs(2116)) and (layer0_outputs(1075)));
    layer1_outputs(679) <= not(layer0_outputs(1989));
    layer1_outputs(680) <= layer0_outputs(791);
    layer1_outputs(681) <= '1';
    layer1_outputs(682) <= layer0_outputs(1369);
    layer1_outputs(683) <= (layer0_outputs(1168)) and not (layer0_outputs(867));
    layer1_outputs(684) <= (layer0_outputs(2484)) and not (layer0_outputs(1040));
    layer1_outputs(685) <= (layer0_outputs(151)) or (layer0_outputs(178));
    layer1_outputs(686) <= not((layer0_outputs(157)) or (layer0_outputs(97)));
    layer1_outputs(687) <= (layer0_outputs(1404)) or (layer0_outputs(1977));
    layer1_outputs(688) <= not(layer0_outputs(1888));
    layer1_outputs(689) <= '1';
    layer1_outputs(690) <= '0';
    layer1_outputs(691) <= (layer0_outputs(81)) xor (layer0_outputs(243));
    layer1_outputs(692) <= (layer0_outputs(267)) and not (layer0_outputs(199));
    layer1_outputs(693) <= (layer0_outputs(659)) or (layer0_outputs(807));
    layer1_outputs(694) <= not((layer0_outputs(2091)) or (layer0_outputs(2045)));
    layer1_outputs(695) <= not((layer0_outputs(303)) and (layer0_outputs(1841)));
    layer1_outputs(696) <= not(layer0_outputs(686)) or (layer0_outputs(737));
    layer1_outputs(697) <= (layer0_outputs(1844)) or (layer0_outputs(1894));
    layer1_outputs(698) <= (layer0_outputs(911)) or (layer0_outputs(1899));
    layer1_outputs(699) <= '0';
    layer1_outputs(700) <= (layer0_outputs(984)) and (layer0_outputs(179));
    layer1_outputs(701) <= (layer0_outputs(2471)) or (layer0_outputs(747));
    layer1_outputs(702) <= '0';
    layer1_outputs(703) <= not(layer0_outputs(670));
    layer1_outputs(704) <= (layer0_outputs(330)) and not (layer0_outputs(2301));
    layer1_outputs(705) <= (layer0_outputs(1162)) and (layer0_outputs(2461));
    layer1_outputs(706) <= (layer0_outputs(176)) and not (layer0_outputs(2308));
    layer1_outputs(707) <= layer0_outputs(2159);
    layer1_outputs(708) <= '1';
    layer1_outputs(709) <= layer0_outputs(1919);
    layer1_outputs(710) <= (layer0_outputs(1242)) and not (layer0_outputs(2466));
    layer1_outputs(711) <= '0';
    layer1_outputs(712) <= not(layer0_outputs(481));
    layer1_outputs(713) <= (layer0_outputs(739)) and not (layer0_outputs(375));
    layer1_outputs(714) <= not((layer0_outputs(2342)) or (layer0_outputs(1087)));
    layer1_outputs(715) <= (layer0_outputs(1697)) and not (layer0_outputs(1359));
    layer1_outputs(716) <= (layer0_outputs(296)) and not (layer0_outputs(2149));
    layer1_outputs(717) <= (layer0_outputs(899)) or (layer0_outputs(704));
    layer1_outputs(718) <= (layer0_outputs(741)) and not (layer0_outputs(1863));
    layer1_outputs(719) <= not(layer0_outputs(2035));
    layer1_outputs(720) <= layer0_outputs(1882);
    layer1_outputs(721) <= layer0_outputs(989);
    layer1_outputs(722) <= not((layer0_outputs(2139)) and (layer0_outputs(1129)));
    layer1_outputs(723) <= not(layer0_outputs(220));
    layer1_outputs(724) <= layer0_outputs(2081);
    layer1_outputs(725) <= not(layer0_outputs(566)) or (layer0_outputs(675));
    layer1_outputs(726) <= (layer0_outputs(1130)) and not (layer0_outputs(2317));
    layer1_outputs(727) <= '1';
    layer1_outputs(728) <= '0';
    layer1_outputs(729) <= not(layer0_outputs(1233));
    layer1_outputs(730) <= not(layer0_outputs(2113)) or (layer0_outputs(994));
    layer1_outputs(731) <= not((layer0_outputs(664)) xor (layer0_outputs(2368)));
    layer1_outputs(732) <= not(layer0_outputs(1017));
    layer1_outputs(733) <= (layer0_outputs(1337)) and not (layer0_outputs(2242));
    layer1_outputs(734) <= (layer0_outputs(188)) or (layer0_outputs(1610));
    layer1_outputs(735) <= (layer0_outputs(169)) and not (layer0_outputs(2466));
    layer1_outputs(736) <= (layer0_outputs(1607)) and (layer0_outputs(1590));
    layer1_outputs(737) <= layer0_outputs(1310);
    layer1_outputs(738) <= '0';
    layer1_outputs(739) <= not(layer0_outputs(2515)) or (layer0_outputs(2336));
    layer1_outputs(740) <= (layer0_outputs(724)) and (layer0_outputs(1962));
    layer1_outputs(741) <= not(layer0_outputs(1468));
    layer1_outputs(742) <= not(layer0_outputs(1852)) or (layer0_outputs(2432));
    layer1_outputs(743) <= (layer0_outputs(1451)) and not (layer0_outputs(682));
    layer1_outputs(744) <= not((layer0_outputs(141)) or (layer0_outputs(1078)));
    layer1_outputs(745) <= (layer0_outputs(1956)) or (layer0_outputs(70));
    layer1_outputs(746) <= (layer0_outputs(1360)) and (layer0_outputs(851));
    layer1_outputs(747) <= (layer0_outputs(1190)) and not (layer0_outputs(1484));
    layer1_outputs(748) <= (layer0_outputs(1554)) and not (layer0_outputs(1136));
    layer1_outputs(749) <= (layer0_outputs(589)) and not (layer0_outputs(597));
    layer1_outputs(750) <= (layer0_outputs(1504)) and not (layer0_outputs(265));
    layer1_outputs(751) <= not(layer0_outputs(737)) or (layer0_outputs(1874));
    layer1_outputs(752) <= '0';
    layer1_outputs(753) <= not((layer0_outputs(1613)) and (layer0_outputs(617)));
    layer1_outputs(754) <= layer0_outputs(1796);
    layer1_outputs(755) <= layer0_outputs(1817);
    layer1_outputs(756) <= '1';
    layer1_outputs(757) <= '1';
    layer1_outputs(758) <= (layer0_outputs(300)) or (layer0_outputs(2227));
    layer1_outputs(759) <= (layer0_outputs(167)) or (layer0_outputs(223));
    layer1_outputs(760) <= not(layer0_outputs(2485)) or (layer0_outputs(1605));
    layer1_outputs(761) <= not((layer0_outputs(2332)) and (layer0_outputs(480)));
    layer1_outputs(762) <= layer0_outputs(2089);
    layer1_outputs(763) <= not(layer0_outputs(770));
    layer1_outputs(764) <= (layer0_outputs(2187)) and (layer0_outputs(927));
    layer1_outputs(765) <= not(layer0_outputs(1578));
    layer1_outputs(766) <= '1';
    layer1_outputs(767) <= '0';
    layer1_outputs(768) <= not(layer0_outputs(678));
    layer1_outputs(769) <= not((layer0_outputs(1060)) and (layer0_outputs(1319)));
    layer1_outputs(770) <= not(layer0_outputs(768)) or (layer0_outputs(1033));
    layer1_outputs(771) <= '0';
    layer1_outputs(772) <= not(layer0_outputs(2110)) or (layer0_outputs(953));
    layer1_outputs(773) <= not(layer0_outputs(570));
    layer1_outputs(774) <= not(layer0_outputs(1509));
    layer1_outputs(775) <= layer0_outputs(635);
    layer1_outputs(776) <= not((layer0_outputs(2143)) and (layer0_outputs(2287)));
    layer1_outputs(777) <= not(layer0_outputs(2163)) or (layer0_outputs(2557));
    layer1_outputs(778) <= not(layer0_outputs(1858)) or (layer0_outputs(1145));
    layer1_outputs(779) <= not(layer0_outputs(338)) or (layer0_outputs(2435));
    layer1_outputs(780) <= not(layer0_outputs(259));
    layer1_outputs(781) <= '0';
    layer1_outputs(782) <= layer0_outputs(2549);
    layer1_outputs(783) <= not(layer0_outputs(755)) or (layer0_outputs(1803));
    layer1_outputs(784) <= not((layer0_outputs(2438)) or (layer0_outputs(1568)));
    layer1_outputs(785) <= '0';
    layer1_outputs(786) <= layer0_outputs(72);
    layer1_outputs(787) <= not(layer0_outputs(446));
    layer1_outputs(788) <= (layer0_outputs(161)) or (layer0_outputs(1637));
    layer1_outputs(789) <= '0';
    layer1_outputs(790) <= not((layer0_outputs(1235)) and (layer0_outputs(682)));
    layer1_outputs(791) <= not(layer0_outputs(1732)) or (layer0_outputs(1985));
    layer1_outputs(792) <= not(layer0_outputs(2099)) or (layer0_outputs(731));
    layer1_outputs(793) <= not((layer0_outputs(1690)) and (layer0_outputs(1167)));
    layer1_outputs(794) <= layer0_outputs(357);
    layer1_outputs(795) <= not(layer0_outputs(512)) or (layer0_outputs(1370));
    layer1_outputs(796) <= layer0_outputs(471);
    layer1_outputs(797) <= not(layer0_outputs(1149)) or (layer0_outputs(586));
    layer1_outputs(798) <= layer0_outputs(333);
    layer1_outputs(799) <= not((layer0_outputs(2375)) or (layer0_outputs(1072)));
    layer1_outputs(800) <= not(layer0_outputs(2444));
    layer1_outputs(801) <= not(layer0_outputs(1883));
    layer1_outputs(802) <= layer0_outputs(114);
    layer1_outputs(803) <= layer0_outputs(1918);
    layer1_outputs(804) <= not((layer0_outputs(563)) and (layer0_outputs(1217)));
    layer1_outputs(805) <= layer0_outputs(1290);
    layer1_outputs(806) <= '0';
    layer1_outputs(807) <= not(layer0_outputs(2550));
    layer1_outputs(808) <= not(layer0_outputs(911)) or (layer0_outputs(2000));
    layer1_outputs(809) <= (layer0_outputs(452)) and not (layer0_outputs(988));
    layer1_outputs(810) <= (layer0_outputs(2100)) and not (layer0_outputs(1667));
    layer1_outputs(811) <= not(layer0_outputs(322)) or (layer0_outputs(928));
    layer1_outputs(812) <= (layer0_outputs(1300)) or (layer0_outputs(1343));
    layer1_outputs(813) <= layer0_outputs(529);
    layer1_outputs(814) <= not(layer0_outputs(1866)) or (layer0_outputs(459));
    layer1_outputs(815) <= (layer0_outputs(1131)) and (layer0_outputs(132));
    layer1_outputs(816) <= (layer0_outputs(2177)) and not (layer0_outputs(236));
    layer1_outputs(817) <= '1';
    layer1_outputs(818) <= '1';
    layer1_outputs(819) <= layer0_outputs(894);
    layer1_outputs(820) <= not(layer0_outputs(2281)) or (layer0_outputs(1302));
    layer1_outputs(821) <= '1';
    layer1_outputs(822) <= '0';
    layer1_outputs(823) <= not(layer0_outputs(2524)) or (layer0_outputs(1371));
    layer1_outputs(824) <= layer0_outputs(2257);
    layer1_outputs(825) <= (layer0_outputs(667)) and not (layer0_outputs(923));
    layer1_outputs(826) <= not((layer0_outputs(1565)) and (layer0_outputs(490)));
    layer1_outputs(827) <= (layer0_outputs(1171)) and not (layer0_outputs(2265));
    layer1_outputs(828) <= not(layer0_outputs(2318));
    layer1_outputs(829) <= not(layer0_outputs(2342));
    layer1_outputs(830) <= not(layer0_outputs(987)) or (layer0_outputs(1844));
    layer1_outputs(831) <= (layer0_outputs(514)) or (layer0_outputs(1187));
    layer1_outputs(832) <= layer0_outputs(2450);
    layer1_outputs(833) <= layer0_outputs(309);
    layer1_outputs(834) <= not(layer0_outputs(564));
    layer1_outputs(835) <= (layer0_outputs(1399)) and not (layer0_outputs(1599));
    layer1_outputs(836) <= '1';
    layer1_outputs(837) <= (layer0_outputs(2359)) and not (layer0_outputs(2298));
    layer1_outputs(838) <= '0';
    layer1_outputs(839) <= layer0_outputs(2134);
    layer1_outputs(840) <= not((layer0_outputs(387)) and (layer0_outputs(1392)));
    layer1_outputs(841) <= '1';
    layer1_outputs(842) <= (layer0_outputs(342)) and (layer0_outputs(870));
    layer1_outputs(843) <= not((layer0_outputs(935)) and (layer0_outputs(274)));
    layer1_outputs(844) <= (layer0_outputs(1876)) and (layer0_outputs(395));
    layer1_outputs(845) <= not(layer0_outputs(707));
    layer1_outputs(846) <= (layer0_outputs(2273)) or (layer0_outputs(2501));
    layer1_outputs(847) <= not((layer0_outputs(2222)) and (layer0_outputs(1336)));
    layer1_outputs(848) <= not(layer0_outputs(792)) or (layer0_outputs(2246));
    layer1_outputs(849) <= layer0_outputs(1593);
    layer1_outputs(850) <= '1';
    layer1_outputs(851) <= (layer0_outputs(1069)) and (layer0_outputs(1441));
    layer1_outputs(852) <= '0';
    layer1_outputs(853) <= (layer0_outputs(549)) or (layer0_outputs(2510));
    layer1_outputs(854) <= '1';
    layer1_outputs(855) <= (layer0_outputs(1273)) or (layer0_outputs(1877));
    layer1_outputs(856) <= not(layer0_outputs(1986)) or (layer0_outputs(228));
    layer1_outputs(857) <= not(layer0_outputs(1251)) or (layer0_outputs(1489));
    layer1_outputs(858) <= (layer0_outputs(2084)) and not (layer0_outputs(1398));
    layer1_outputs(859) <= layer0_outputs(2027);
    layer1_outputs(860) <= not((layer0_outputs(2258)) or (layer0_outputs(1644)));
    layer1_outputs(861) <= '1';
    layer1_outputs(862) <= not((layer0_outputs(627)) or (layer0_outputs(602)));
    layer1_outputs(863) <= (layer0_outputs(1151)) or (layer0_outputs(2388));
    layer1_outputs(864) <= '1';
    layer1_outputs(865) <= (layer0_outputs(638)) and not (layer0_outputs(85));
    layer1_outputs(866) <= not((layer0_outputs(1343)) or (layer0_outputs(1875)));
    layer1_outputs(867) <= layer0_outputs(871);
    layer1_outputs(868) <= '1';
    layer1_outputs(869) <= not((layer0_outputs(1585)) and (layer0_outputs(890)));
    layer1_outputs(870) <= not((layer0_outputs(226)) xor (layer0_outputs(907)));
    layer1_outputs(871) <= not(layer0_outputs(1712));
    layer1_outputs(872) <= layer0_outputs(1639);
    layer1_outputs(873) <= '0';
    layer1_outputs(874) <= layer0_outputs(255);
    layer1_outputs(875) <= layer0_outputs(1964);
    layer1_outputs(876) <= '1';
    layer1_outputs(877) <= '0';
    layer1_outputs(878) <= (layer0_outputs(2498)) or (layer0_outputs(1715));
    layer1_outputs(879) <= not(layer0_outputs(1341)) or (layer0_outputs(543));
    layer1_outputs(880) <= '0';
    layer1_outputs(881) <= (layer0_outputs(1319)) and not (layer0_outputs(1068));
    layer1_outputs(882) <= not((layer0_outputs(107)) or (layer0_outputs(2261)));
    layer1_outputs(883) <= (layer0_outputs(1222)) and not (layer0_outputs(321));
    layer1_outputs(884) <= not(layer0_outputs(177)) or (layer0_outputs(653));
    layer1_outputs(885) <= '1';
    layer1_outputs(886) <= not(layer0_outputs(1183));
    layer1_outputs(887) <= not((layer0_outputs(1811)) xor (layer0_outputs(1783)));
    layer1_outputs(888) <= '1';
    layer1_outputs(889) <= not(layer0_outputs(1472)) or (layer0_outputs(2177));
    layer1_outputs(890) <= '1';
    layer1_outputs(891) <= '1';
    layer1_outputs(892) <= (layer0_outputs(407)) and (layer0_outputs(2085));
    layer1_outputs(893) <= not(layer0_outputs(1452));
    layer1_outputs(894) <= not((layer0_outputs(2348)) or (layer0_outputs(1630)));
    layer1_outputs(895) <= (layer0_outputs(1618)) and (layer0_outputs(1486));
    layer1_outputs(896) <= (layer0_outputs(37)) and (layer0_outputs(1062));
    layer1_outputs(897) <= not(layer0_outputs(2064));
    layer1_outputs(898) <= layer0_outputs(2413);
    layer1_outputs(899) <= '1';
    layer1_outputs(900) <= not(layer0_outputs(453)) or (layer0_outputs(2336));
    layer1_outputs(901) <= (layer0_outputs(1503)) or (layer0_outputs(1477));
    layer1_outputs(902) <= not((layer0_outputs(170)) or (layer0_outputs(550)));
    layer1_outputs(903) <= not((layer0_outputs(496)) or (layer0_outputs(2165)));
    layer1_outputs(904) <= not(layer0_outputs(2230));
    layer1_outputs(905) <= not(layer0_outputs(516)) or (layer0_outputs(617));
    layer1_outputs(906) <= '0';
    layer1_outputs(907) <= '0';
    layer1_outputs(908) <= '1';
    layer1_outputs(909) <= '0';
    layer1_outputs(910) <= (layer0_outputs(1144)) and not (layer0_outputs(643));
    layer1_outputs(911) <= (layer0_outputs(644)) and (layer0_outputs(80));
    layer1_outputs(912) <= '0';
    layer1_outputs(913) <= '1';
    layer1_outputs(914) <= '0';
    layer1_outputs(915) <= not(layer0_outputs(2077));
    layer1_outputs(916) <= layer0_outputs(412);
    layer1_outputs(917) <= (layer0_outputs(1908)) and not (layer0_outputs(1763));
    layer1_outputs(918) <= layer0_outputs(1238);
    layer1_outputs(919) <= (layer0_outputs(1541)) or (layer0_outputs(1878));
    layer1_outputs(920) <= not(layer0_outputs(1435)) or (layer0_outputs(256));
    layer1_outputs(921) <= not(layer0_outputs(1309)) or (layer0_outputs(213));
    layer1_outputs(922) <= layer0_outputs(2046);
    layer1_outputs(923) <= not(layer0_outputs(1837));
    layer1_outputs(924) <= not((layer0_outputs(1565)) or (layer0_outputs(2531)));
    layer1_outputs(925) <= not(layer0_outputs(2105));
    layer1_outputs(926) <= layer0_outputs(1417);
    layer1_outputs(927) <= layer0_outputs(2435);
    layer1_outputs(928) <= not(layer0_outputs(1289));
    layer1_outputs(929) <= (layer0_outputs(1213)) and (layer0_outputs(1723));
    layer1_outputs(930) <= (layer0_outputs(2332)) and not (layer0_outputs(404));
    layer1_outputs(931) <= not(layer0_outputs(1190)) or (layer0_outputs(2207));
    layer1_outputs(932) <= '0';
    layer1_outputs(933) <= '0';
    layer1_outputs(934) <= not((layer0_outputs(500)) or (layer0_outputs(652)));
    layer1_outputs(935) <= not(layer0_outputs(1175));
    layer1_outputs(936) <= not(layer0_outputs(517));
    layer1_outputs(937) <= not(layer0_outputs(957));
    layer1_outputs(938) <= not(layer0_outputs(2117));
    layer1_outputs(939) <= '0';
    layer1_outputs(940) <= not(layer0_outputs(1831)) or (layer0_outputs(2376));
    layer1_outputs(941) <= (layer0_outputs(2198)) or (layer0_outputs(2267));
    layer1_outputs(942) <= not((layer0_outputs(611)) and (layer0_outputs(772)));
    layer1_outputs(943) <= not(layer0_outputs(1794)) or (layer0_outputs(1204));
    layer1_outputs(944) <= (layer0_outputs(775)) and not (layer0_outputs(2049));
    layer1_outputs(945) <= layer0_outputs(1694);
    layer1_outputs(946) <= not(layer0_outputs(699)) or (layer0_outputs(277));
    layer1_outputs(947) <= (layer0_outputs(1371)) and not (layer0_outputs(943));
    layer1_outputs(948) <= layer0_outputs(2436);
    layer1_outputs(949) <= layer0_outputs(2016);
    layer1_outputs(950) <= not((layer0_outputs(752)) or (layer0_outputs(419)));
    layer1_outputs(951) <= (layer0_outputs(873)) and not (layer0_outputs(1245));
    layer1_outputs(952) <= layer0_outputs(410);
    layer1_outputs(953) <= (layer0_outputs(1793)) and not (layer0_outputs(1589));
    layer1_outputs(954) <= '1';
    layer1_outputs(955) <= (layer0_outputs(1089)) or (layer0_outputs(1804));
    layer1_outputs(956) <= not(layer0_outputs(833)) or (layer0_outputs(1959));
    layer1_outputs(957) <= '1';
    layer1_outputs(958) <= (layer0_outputs(1253)) and (layer0_outputs(641));
    layer1_outputs(959) <= (layer0_outputs(406)) and not (layer0_outputs(1207));
    layer1_outputs(960) <= not(layer0_outputs(466)) or (layer0_outputs(1984));
    layer1_outputs(961) <= '1';
    layer1_outputs(962) <= not(layer0_outputs(55));
    layer1_outputs(963) <= layer0_outputs(894);
    layer1_outputs(964) <= (layer0_outputs(2472)) and not (layer0_outputs(415));
    layer1_outputs(965) <= not((layer0_outputs(456)) or (layer0_outputs(1594)));
    layer1_outputs(966) <= '1';
    layer1_outputs(967) <= (layer0_outputs(713)) or (layer0_outputs(1810));
    layer1_outputs(968) <= (layer0_outputs(1217)) and (layer0_outputs(1721));
    layer1_outputs(969) <= layer0_outputs(1064);
    layer1_outputs(970) <= '1';
    layer1_outputs(971) <= not(layer0_outputs(10));
    layer1_outputs(972) <= not(layer0_outputs(588));
    layer1_outputs(973) <= not(layer0_outputs(972));
    layer1_outputs(974) <= '0';
    layer1_outputs(975) <= '1';
    layer1_outputs(976) <= not((layer0_outputs(263)) xor (layer0_outputs(1272)));
    layer1_outputs(977) <= layer0_outputs(1588);
    layer1_outputs(978) <= not(layer0_outputs(1982)) or (layer0_outputs(1497));
    layer1_outputs(979) <= not(layer0_outputs(1526));
    layer1_outputs(980) <= (layer0_outputs(61)) or (layer0_outputs(1044));
    layer1_outputs(981) <= layer0_outputs(1208);
    layer1_outputs(982) <= layer0_outputs(2178);
    layer1_outputs(983) <= '0';
    layer1_outputs(984) <= not((layer0_outputs(136)) and (layer0_outputs(626)));
    layer1_outputs(985) <= '1';
    layer1_outputs(986) <= (layer0_outputs(122)) and (layer0_outputs(886));
    layer1_outputs(987) <= layer0_outputs(2381);
    layer1_outputs(988) <= layer0_outputs(67);
    layer1_outputs(989) <= '0';
    layer1_outputs(990) <= not((layer0_outputs(1633)) or (layer0_outputs(449)));
    layer1_outputs(991) <= (layer0_outputs(1972)) and not (layer0_outputs(545));
    layer1_outputs(992) <= (layer0_outputs(859)) and (layer0_outputs(622));
    layer1_outputs(993) <= (layer0_outputs(751)) and (layer0_outputs(1085));
    layer1_outputs(994) <= '1';
    layer1_outputs(995) <= not((layer0_outputs(925)) and (layer0_outputs(2345)));
    layer1_outputs(996) <= not(layer0_outputs(620)) or (layer0_outputs(2116));
    layer1_outputs(997) <= layer0_outputs(1945);
    layer1_outputs(998) <= '0';
    layer1_outputs(999) <= not((layer0_outputs(503)) and (layer0_outputs(2291)));
    layer1_outputs(1000) <= (layer0_outputs(2463)) and (layer0_outputs(1431));
    layer1_outputs(1001) <= not(layer0_outputs(1085));
    layer1_outputs(1002) <= layer0_outputs(1273);
    layer1_outputs(1003) <= not(layer0_outputs(411));
    layer1_outputs(1004) <= '1';
    layer1_outputs(1005) <= (layer0_outputs(2429)) and not (layer0_outputs(2270));
    layer1_outputs(1006) <= not(layer0_outputs(849)) or (layer0_outputs(2445));
    layer1_outputs(1007) <= (layer0_outputs(1736)) and not (layer0_outputs(2145));
    layer1_outputs(1008) <= not((layer0_outputs(931)) and (layer0_outputs(2211)));
    layer1_outputs(1009) <= not(layer0_outputs(1167));
    layer1_outputs(1010) <= not(layer0_outputs(1655)) or (layer0_outputs(474));
    layer1_outputs(1011) <= '0';
    layer1_outputs(1012) <= not(layer0_outputs(1505));
    layer1_outputs(1013) <= (layer0_outputs(818)) and not (layer0_outputs(1654));
    layer1_outputs(1014) <= not(layer0_outputs(929));
    layer1_outputs(1015) <= layer0_outputs(1313);
    layer1_outputs(1016) <= not((layer0_outputs(1731)) and (layer0_outputs(293)));
    layer1_outputs(1017) <= '1';
    layer1_outputs(1018) <= not((layer0_outputs(40)) and (layer0_outputs(1657)));
    layer1_outputs(1019) <= (layer0_outputs(607)) and not (layer0_outputs(2323));
    layer1_outputs(1020) <= '0';
    layer1_outputs(1021) <= (layer0_outputs(1976)) and not (layer0_outputs(1355));
    layer1_outputs(1022) <= (layer0_outputs(2277)) or (layer0_outputs(758));
    layer1_outputs(1023) <= '1';
    layer1_outputs(1024) <= (layer0_outputs(836)) and not (layer0_outputs(2333));
    layer1_outputs(1025) <= not(layer0_outputs(2431)) or (layer0_outputs(431));
    layer1_outputs(1026) <= (layer0_outputs(1443)) and not (layer0_outputs(392));
    layer1_outputs(1027) <= layer0_outputs(874);
    layer1_outputs(1028) <= not(layer0_outputs(2460)) or (layer0_outputs(1678));
    layer1_outputs(1029) <= '1';
    layer1_outputs(1030) <= '0';
    layer1_outputs(1031) <= not(layer0_outputs(2098)) or (layer0_outputs(2042));
    layer1_outputs(1032) <= '0';
    layer1_outputs(1033) <= not(layer0_outputs(2077));
    layer1_outputs(1034) <= layer0_outputs(1859);
    layer1_outputs(1035) <= (layer0_outputs(567)) and not (layer0_outputs(602));
    layer1_outputs(1036) <= '0';
    layer1_outputs(1037) <= (layer0_outputs(960)) and not (layer0_outputs(350));
    layer1_outputs(1038) <= (layer0_outputs(2153)) or (layer0_outputs(1091));
    layer1_outputs(1039) <= not(layer0_outputs(2050));
    layer1_outputs(1040) <= layer0_outputs(2307);
    layer1_outputs(1041) <= not((layer0_outputs(1216)) or (layer0_outputs(1413)));
    layer1_outputs(1042) <= not((layer0_outputs(700)) or (layer0_outputs(685)));
    layer1_outputs(1043) <= (layer0_outputs(1611)) and not (layer0_outputs(2496));
    layer1_outputs(1044) <= '0';
    layer1_outputs(1045) <= not(layer0_outputs(2028)) or (layer0_outputs(2543));
    layer1_outputs(1046) <= not(layer0_outputs(241));
    layer1_outputs(1047) <= not(layer0_outputs(1962)) or (layer0_outputs(2090));
    layer1_outputs(1048) <= (layer0_outputs(347)) or (layer0_outputs(1049));
    layer1_outputs(1049) <= not((layer0_outputs(1615)) and (layer0_outputs(1467)));
    layer1_outputs(1050) <= not(layer0_outputs(1738)) or (layer0_outputs(2094));
    layer1_outputs(1051) <= not(layer0_outputs(2096));
    layer1_outputs(1052) <= layer0_outputs(2118);
    layer1_outputs(1053) <= not(layer0_outputs(398)) or (layer0_outputs(1752));
    layer1_outputs(1054) <= not(layer0_outputs(2174)) or (layer0_outputs(235));
    layer1_outputs(1055) <= (layer0_outputs(368)) and not (layer0_outputs(1049));
    layer1_outputs(1056) <= not((layer0_outputs(1828)) and (layer0_outputs(2038)));
    layer1_outputs(1057) <= not(layer0_outputs(142)) or (layer0_outputs(1773));
    layer1_outputs(1058) <= not((layer0_outputs(148)) and (layer0_outputs(1542)));
    layer1_outputs(1059) <= (layer0_outputs(232)) and not (layer0_outputs(351));
    layer1_outputs(1060) <= '0';
    layer1_outputs(1061) <= '1';
    layer1_outputs(1062) <= not(layer0_outputs(1084));
    layer1_outputs(1063) <= not((layer0_outputs(78)) or (layer0_outputs(904)));
    layer1_outputs(1064) <= not(layer0_outputs(1416)) or (layer0_outputs(1472));
    layer1_outputs(1065) <= (layer0_outputs(2548)) xor (layer0_outputs(195));
    layer1_outputs(1066) <= '0';
    layer1_outputs(1067) <= (layer0_outputs(121)) and not (layer0_outputs(2474));
    layer1_outputs(1068) <= (layer0_outputs(1547)) and not (layer0_outputs(1733));
    layer1_outputs(1069) <= not((layer0_outputs(1952)) or (layer0_outputs(2522)));
    layer1_outputs(1070) <= '1';
    layer1_outputs(1071) <= not((layer0_outputs(1798)) or (layer0_outputs(1027)));
    layer1_outputs(1072) <= not((layer0_outputs(1185)) xor (layer0_outputs(2400)));
    layer1_outputs(1073) <= (layer0_outputs(28)) and not (layer0_outputs(559));
    layer1_outputs(1074) <= layer0_outputs(155);
    layer1_outputs(1075) <= not(layer0_outputs(732)) or (layer0_outputs(1801));
    layer1_outputs(1076) <= '0';
    layer1_outputs(1077) <= not(layer0_outputs(800));
    layer1_outputs(1078) <= '1';
    layer1_outputs(1079) <= not(layer0_outputs(1293)) or (layer0_outputs(1653));
    layer1_outputs(1080) <= (layer0_outputs(2370)) or (layer0_outputs(1018));
    layer1_outputs(1081) <= '0';
    layer1_outputs(1082) <= not(layer0_outputs(1)) or (layer0_outputs(2205));
    layer1_outputs(1083) <= layer0_outputs(2244);
    layer1_outputs(1084) <= '0';
    layer1_outputs(1085) <= '1';
    layer1_outputs(1086) <= (layer0_outputs(273)) or (layer0_outputs(865));
    layer1_outputs(1087) <= (layer0_outputs(1875)) and not (layer0_outputs(872));
    layer1_outputs(1088) <= not(layer0_outputs(251));
    layer1_outputs(1089) <= (layer0_outputs(1275)) and not (layer0_outputs(402));
    layer1_outputs(1090) <= (layer0_outputs(2195)) and (layer0_outputs(837));
    layer1_outputs(1091) <= (layer0_outputs(26)) and not (layer0_outputs(680));
    layer1_outputs(1092) <= (layer0_outputs(316)) and not (layer0_outputs(1305));
    layer1_outputs(1093) <= '1';
    layer1_outputs(1094) <= (layer0_outputs(930)) and (layer0_outputs(876));
    layer1_outputs(1095) <= '1';
    layer1_outputs(1096) <= (layer0_outputs(1882)) and (layer0_outputs(1537));
    layer1_outputs(1097) <= '1';
    layer1_outputs(1098) <= not((layer0_outputs(1682)) or (layer0_outputs(705)));
    layer1_outputs(1099) <= '0';
    layer1_outputs(1100) <= '1';
    layer1_outputs(1101) <= not((layer0_outputs(1232)) or (layer0_outputs(980)));
    layer1_outputs(1102) <= (layer0_outputs(1012)) and not (layer0_outputs(1587));
    layer1_outputs(1103) <= (layer0_outputs(1942)) and not (layer0_outputs(1784));
    layer1_outputs(1104) <= not((layer0_outputs(676)) and (layer0_outputs(1884)));
    layer1_outputs(1105) <= not(layer0_outputs(1606)) or (layer0_outputs(1868));
    layer1_outputs(1106) <= (layer0_outputs(792)) and not (layer0_outputs(185));
    layer1_outputs(1107) <= not(layer0_outputs(1123));
    layer1_outputs(1108) <= '0';
    layer1_outputs(1109) <= layer0_outputs(1553);
    layer1_outputs(1110) <= layer0_outputs(1398);
    layer1_outputs(1111) <= layer0_outputs(124);
    layer1_outputs(1112) <= not(layer0_outputs(1416));
    layer1_outputs(1113) <= (layer0_outputs(1055)) or (layer0_outputs(424));
    layer1_outputs(1114) <= layer0_outputs(346);
    layer1_outputs(1115) <= (layer0_outputs(1911)) and not (layer0_outputs(1730));
    layer1_outputs(1116) <= (layer0_outputs(573)) xor (layer0_outputs(7));
    layer1_outputs(1117) <= (layer0_outputs(1640)) and not (layer0_outputs(1310));
    layer1_outputs(1118) <= (layer0_outputs(1330)) and not (layer0_outputs(2221));
    layer1_outputs(1119) <= '1';
    layer1_outputs(1120) <= '0';
    layer1_outputs(1121) <= '1';
    layer1_outputs(1122) <= '1';
    layer1_outputs(1123) <= layer0_outputs(1048);
    layer1_outputs(1124) <= (layer0_outputs(1560)) and not (layer0_outputs(690));
    layer1_outputs(1125) <= (layer0_outputs(2320)) and (layer0_outputs(837));
    layer1_outputs(1126) <= not((layer0_outputs(2442)) and (layer0_outputs(2190)));
    layer1_outputs(1127) <= not(layer0_outputs(1315));
    layer1_outputs(1128) <= (layer0_outputs(767)) and (layer0_outputs(986));
    layer1_outputs(1129) <= (layer0_outputs(2281)) and (layer0_outputs(102));
    layer1_outputs(1130) <= layer0_outputs(1598);
    layer1_outputs(1131) <= '1';
    layer1_outputs(1132) <= '1';
    layer1_outputs(1133) <= not((layer0_outputs(1070)) and (layer0_outputs(1580)));
    layer1_outputs(1134) <= not(layer0_outputs(2503)) or (layer0_outputs(200));
    layer1_outputs(1135) <= layer0_outputs(2519);
    layer1_outputs(1136) <= (layer0_outputs(1660)) or (layer0_outputs(1734));
    layer1_outputs(1137) <= '1';
    layer1_outputs(1138) <= '1';
    layer1_outputs(1139) <= '1';
    layer1_outputs(1140) <= '0';
    layer1_outputs(1141) <= not((layer0_outputs(507)) and (layer0_outputs(115)));
    layer1_outputs(1142) <= (layer0_outputs(1174)) and not (layer0_outputs(1782));
    layer1_outputs(1143) <= not((layer0_outputs(294)) or (layer0_outputs(615)));
    layer1_outputs(1144) <= not((layer0_outputs(36)) or (layer0_outputs(2243)));
    layer1_outputs(1145) <= '0';
    layer1_outputs(1146) <= (layer0_outputs(131)) or (layer0_outputs(1634));
    layer1_outputs(1147) <= layer0_outputs(833);
    layer1_outputs(1148) <= layer0_outputs(1424);
    layer1_outputs(1149) <= '0';
    layer1_outputs(1150) <= not((layer0_outputs(1304)) and (layer0_outputs(146)));
    layer1_outputs(1151) <= not(layer0_outputs(216)) or (layer0_outputs(565));
    layer1_outputs(1152) <= not((layer0_outputs(206)) xor (layer0_outputs(153)));
    layer1_outputs(1153) <= '0';
    layer1_outputs(1154) <= (layer0_outputs(64)) and not (layer0_outputs(774));
    layer1_outputs(1155) <= (layer0_outputs(182)) and not (layer0_outputs(2192));
    layer1_outputs(1156) <= not(layer0_outputs(2425)) or (layer0_outputs(1307));
    layer1_outputs(1157) <= (layer0_outputs(1679)) and (layer0_outputs(157));
    layer1_outputs(1158) <= '0';
    layer1_outputs(1159) <= not((layer0_outputs(1005)) or (layer0_outputs(1424)));
    layer1_outputs(1160) <= not(layer0_outputs(1267));
    layer1_outputs(1161) <= (layer0_outputs(399)) or (layer0_outputs(589));
    layer1_outputs(1162) <= not(layer0_outputs(2556)) or (layer0_outputs(1745));
    layer1_outputs(1163) <= '0';
    layer1_outputs(1164) <= not(layer0_outputs(1231)) or (layer0_outputs(906));
    layer1_outputs(1165) <= not(layer0_outputs(1329)) or (layer0_outputs(4));
    layer1_outputs(1166) <= not((layer0_outputs(1024)) or (layer0_outputs(234)));
    layer1_outputs(1167) <= (layer0_outputs(1858)) and (layer0_outputs(1707));
    layer1_outputs(1168) <= (layer0_outputs(2194)) and not (layer0_outputs(1892));
    layer1_outputs(1169) <= not(layer0_outputs(1660)) or (layer0_outputs(1369));
    layer1_outputs(1170) <= layer0_outputs(2322);
    layer1_outputs(1171) <= '0';
    layer1_outputs(1172) <= layer0_outputs(1260);
    layer1_outputs(1173) <= layer0_outputs(686);
    layer1_outputs(1174) <= not(layer0_outputs(2204)) or (layer0_outputs(1488));
    layer1_outputs(1175) <= (layer0_outputs(1407)) and not (layer0_outputs(967));
    layer1_outputs(1176) <= '1';
    layer1_outputs(1177) <= (layer0_outputs(2245)) and not (layer0_outputs(2529));
    layer1_outputs(1178) <= not(layer0_outputs(1100));
    layer1_outputs(1179) <= '0';
    layer1_outputs(1180) <= layer0_outputs(1412);
    layer1_outputs(1181) <= (layer0_outputs(280)) or (layer0_outputs(616));
    layer1_outputs(1182) <= layer0_outputs(842);
    layer1_outputs(1183) <= (layer0_outputs(2119)) and (layer0_outputs(1114));
    layer1_outputs(1184) <= not(layer0_outputs(156)) or (layer0_outputs(374));
    layer1_outputs(1185) <= not(layer0_outputs(2004));
    layer1_outputs(1186) <= (layer0_outputs(1746)) and not (layer0_outputs(50));
    layer1_outputs(1187) <= layer0_outputs(1965);
    layer1_outputs(1188) <= '0';
    layer1_outputs(1189) <= layer0_outputs(742);
    layer1_outputs(1190) <= '1';
    layer1_outputs(1191) <= not(layer0_outputs(309)) or (layer0_outputs(759));
    layer1_outputs(1192) <= not(layer0_outputs(886));
    layer1_outputs(1193) <= (layer0_outputs(328)) or (layer0_outputs(923));
    layer1_outputs(1194) <= layer0_outputs(278);
    layer1_outputs(1195) <= '0';
    layer1_outputs(1196) <= not(layer0_outputs(601)) or (layer0_outputs(2431));
    layer1_outputs(1197) <= '1';
    layer1_outputs(1198) <= (layer0_outputs(1413)) and not (layer0_outputs(1410));
    layer1_outputs(1199) <= not(layer0_outputs(270));
    layer1_outputs(1200) <= not((layer0_outputs(378)) or (layer0_outputs(378)));
    layer1_outputs(1201) <= layer0_outputs(569);
    layer1_outputs(1202) <= not(layer0_outputs(673)) or (layer0_outputs(391));
    layer1_outputs(1203) <= '1';
    layer1_outputs(1204) <= not((layer0_outputs(1138)) and (layer0_outputs(2086)));
    layer1_outputs(1205) <= (layer0_outputs(706)) and (layer0_outputs(811));
    layer1_outputs(1206) <= not((layer0_outputs(1066)) and (layer0_outputs(1043)));
    layer1_outputs(1207) <= (layer0_outputs(1000)) or (layer0_outputs(133));
    layer1_outputs(1208) <= layer0_outputs(2096);
    layer1_outputs(1209) <= not(layer0_outputs(1976)) or (layer0_outputs(372));
    layer1_outputs(1210) <= (layer0_outputs(1943)) and not (layer0_outputs(1220));
    layer1_outputs(1211) <= layer0_outputs(2369);
    layer1_outputs(1212) <= '0';
    layer1_outputs(1213) <= layer0_outputs(1815);
    layer1_outputs(1214) <= not((layer0_outputs(636)) or (layer0_outputs(1678)));
    layer1_outputs(1215) <= (layer0_outputs(893)) and (layer0_outputs(557));
    layer1_outputs(1216) <= not(layer0_outputs(20));
    layer1_outputs(1217) <= (layer0_outputs(320)) and (layer0_outputs(1109));
    layer1_outputs(1218) <= '1';
    layer1_outputs(1219) <= layer0_outputs(191);
    layer1_outputs(1220) <= not(layer0_outputs(1444));
    layer1_outputs(1221) <= (layer0_outputs(1052)) and (layer0_outputs(1786));
    layer1_outputs(1222) <= (layer0_outputs(0)) and not (layer0_outputs(106));
    layer1_outputs(1223) <= not(layer0_outputs(183));
    layer1_outputs(1224) <= (layer0_outputs(2013)) or (layer0_outputs(2072));
    layer1_outputs(1225) <= not(layer0_outputs(1458));
    layer1_outputs(1226) <= not((layer0_outputs(1658)) and (layer0_outputs(1732)));
    layer1_outputs(1227) <= '0';
    layer1_outputs(1228) <= '1';
    layer1_outputs(1229) <= not(layer0_outputs(978));
    layer1_outputs(1230) <= layer0_outputs(968);
    layer1_outputs(1231) <= not((layer0_outputs(394)) and (layer0_outputs(930)));
    layer1_outputs(1232) <= '0';
    layer1_outputs(1233) <= '1';
    layer1_outputs(1234) <= '0';
    layer1_outputs(1235) <= layer0_outputs(1719);
    layer1_outputs(1236) <= not(layer0_outputs(1445));
    layer1_outputs(1237) <= not((layer0_outputs(2137)) and (layer0_outputs(1691)));
    layer1_outputs(1238) <= layer0_outputs(371);
    layer1_outputs(1239) <= '1';
    layer1_outputs(1240) <= not(layer0_outputs(1771));
    layer1_outputs(1241) <= (layer0_outputs(952)) and not (layer0_outputs(2536));
    layer1_outputs(1242) <= '0';
    layer1_outputs(1243) <= (layer0_outputs(2380)) and not (layer0_outputs(1018));
    layer1_outputs(1244) <= not(layer0_outputs(1720)) or (layer0_outputs(414));
    layer1_outputs(1245) <= not(layer0_outputs(2488)) or (layer0_outputs(1594));
    layer1_outputs(1246) <= layer0_outputs(1350);
    layer1_outputs(1247) <= not(layer0_outputs(872));
    layer1_outputs(1248) <= layer0_outputs(1983);
    layer1_outputs(1249) <= not((layer0_outputs(1125)) and (layer0_outputs(317)));
    layer1_outputs(1250) <= (layer0_outputs(1143)) or (layer0_outputs(556));
    layer1_outputs(1251) <= '1';
    layer1_outputs(1252) <= not((layer0_outputs(2113)) and (layer0_outputs(2473)));
    layer1_outputs(1253) <= not((layer0_outputs(1193)) or (layer0_outputs(1995)));
    layer1_outputs(1254) <= '0';
    layer1_outputs(1255) <= not(layer0_outputs(1059)) or (layer0_outputs(2272));
    layer1_outputs(1256) <= '1';
    layer1_outputs(1257) <= not(layer0_outputs(405)) or (layer0_outputs(498));
    layer1_outputs(1258) <= (layer0_outputs(1832)) or (layer0_outputs(2436));
    layer1_outputs(1259) <= not((layer0_outputs(2188)) xor (layer0_outputs(841)));
    layer1_outputs(1260) <= not((layer0_outputs(2512)) and (layer0_outputs(634)));
    layer1_outputs(1261) <= (layer0_outputs(2090)) and not (layer0_outputs(1025));
    layer1_outputs(1262) <= not(layer0_outputs(1677)) or (layer0_outputs(415));
    layer1_outputs(1263) <= layer0_outputs(786);
    layer1_outputs(1264) <= (layer0_outputs(1543)) and (layer0_outputs(1511));
    layer1_outputs(1265) <= '0';
    layer1_outputs(1266) <= layer0_outputs(2537);
    layer1_outputs(1267) <= not((layer0_outputs(2519)) or (layer0_outputs(1136)));
    layer1_outputs(1268) <= (layer0_outputs(2091)) xor (layer0_outputs(2249));
    layer1_outputs(1269) <= (layer0_outputs(1215)) or (layer0_outputs(2322));
    layer1_outputs(1270) <= layer0_outputs(2008);
    layer1_outputs(1271) <= layer0_outputs(2060);
    layer1_outputs(1272) <= (layer0_outputs(2472)) and (layer0_outputs(571));
    layer1_outputs(1273) <= '0';
    layer1_outputs(1274) <= not(layer0_outputs(734)) or (layer0_outputs(1712));
    layer1_outputs(1275) <= not(layer0_outputs(698)) or (layer0_outputs(1146));
    layer1_outputs(1276) <= layer0_outputs(1054);
    layer1_outputs(1277) <= not(layer0_outputs(1120));
    layer1_outputs(1278) <= not(layer0_outputs(2020)) or (layer0_outputs(1517));
    layer1_outputs(1279) <= not(layer0_outputs(2386)) or (layer0_outputs(325));
    layer1_outputs(1280) <= (layer0_outputs(552)) and (layer0_outputs(1722));
    layer1_outputs(1281) <= layer0_outputs(2452);
    layer1_outputs(1282) <= '1';
    layer1_outputs(1283) <= '0';
    layer1_outputs(1284) <= not(layer0_outputs(1131));
    layer1_outputs(1285) <= (layer0_outputs(2196)) and (layer0_outputs(698));
    layer1_outputs(1286) <= '0';
    layer1_outputs(1287) <= (layer0_outputs(262)) and not (layer0_outputs(1997));
    layer1_outputs(1288) <= not(layer0_outputs(2286));
    layer1_outputs(1289) <= not(layer0_outputs(2554)) or (layer0_outputs(36));
    layer1_outputs(1290) <= (layer0_outputs(646)) or (layer0_outputs(121));
    layer1_outputs(1291) <= (layer0_outputs(1228)) or (layer0_outputs(1755));
    layer1_outputs(1292) <= '1';
    layer1_outputs(1293) <= (layer0_outputs(1789)) xor (layer0_outputs(1113));
    layer1_outputs(1294) <= layer0_outputs(417);
    layer1_outputs(1295) <= not(layer0_outputs(1036));
    layer1_outputs(1296) <= not((layer0_outputs(1189)) or (layer0_outputs(875)));
    layer1_outputs(1297) <= (layer0_outputs(922)) or (layer0_outputs(256));
    layer1_outputs(1298) <= '0';
    layer1_outputs(1299) <= (layer0_outputs(2019)) and not (layer0_outputs(781));
    layer1_outputs(1300) <= (layer0_outputs(1771)) and not (layer0_outputs(803));
    layer1_outputs(1301) <= (layer0_outputs(163)) or (layer0_outputs(1656));
    layer1_outputs(1302) <= '0';
    layer1_outputs(1303) <= (layer0_outputs(1698)) xor (layer0_outputs(1381));
    layer1_outputs(1304) <= not((layer0_outputs(1941)) and (layer0_outputs(1960)));
    layer1_outputs(1305) <= not(layer0_outputs(58));
    layer1_outputs(1306) <= not(layer0_outputs(1862));
    layer1_outputs(1307) <= not((layer0_outputs(198)) or (layer0_outputs(1170)));
    layer1_outputs(1308) <= not(layer0_outputs(1518));
    layer1_outputs(1309) <= (layer0_outputs(708)) or (layer0_outputs(1880));
    layer1_outputs(1310) <= not(layer0_outputs(2558));
    layer1_outputs(1311) <= layer0_outputs(2309);
    layer1_outputs(1312) <= '1';
    layer1_outputs(1313) <= layer0_outputs(2135);
    layer1_outputs(1314) <= (layer0_outputs(464)) and not (layer0_outputs(2298));
    layer1_outputs(1315) <= (layer0_outputs(1893)) and not (layer0_outputs(879));
    layer1_outputs(1316) <= '1';
    layer1_outputs(1317) <= (layer0_outputs(1538)) or (layer0_outputs(1340));
    layer1_outputs(1318) <= not(layer0_outputs(540)) or (layer0_outputs(663));
    layer1_outputs(1319) <= '1';
    layer1_outputs(1320) <= not(layer0_outputs(219));
    layer1_outputs(1321) <= '1';
    layer1_outputs(1322) <= layer0_outputs(2475);
    layer1_outputs(1323) <= not((layer0_outputs(1536)) and (layer0_outputs(201)));
    layer1_outputs(1324) <= not(layer0_outputs(384)) or (layer0_outputs(1379));
    layer1_outputs(1325) <= '0';
    layer1_outputs(1326) <= not(layer0_outputs(536));
    layer1_outputs(1327) <= not(layer0_outputs(1110));
    layer1_outputs(1328) <= (layer0_outputs(684)) and not (layer0_outputs(2546));
    layer1_outputs(1329) <= not(layer0_outputs(2418));
    layer1_outputs(1330) <= (layer0_outputs(853)) or (layer0_outputs(488));
    layer1_outputs(1331) <= '1';
    layer1_outputs(1332) <= not(layer0_outputs(2335));
    layer1_outputs(1333) <= not((layer0_outputs(1346)) xor (layer0_outputs(2082)));
    layer1_outputs(1334) <= (layer0_outputs(1742)) and not (layer0_outputs(1652));
    layer1_outputs(1335) <= (layer0_outputs(1785)) or (layer0_outputs(614));
    layer1_outputs(1336) <= '1';
    layer1_outputs(1337) <= (layer0_outputs(1194)) and (layer0_outputs(499));
    layer1_outputs(1338) <= layer0_outputs(1846);
    layer1_outputs(1339) <= not(layer0_outputs(702)) or (layer0_outputs(522));
    layer1_outputs(1340) <= not(layer0_outputs(2067));
    layer1_outputs(1341) <= not((layer0_outputs(1806)) and (layer0_outputs(0)));
    layer1_outputs(1342) <= not(layer0_outputs(852)) or (layer0_outputs(1461));
    layer1_outputs(1343) <= not(layer0_outputs(2511)) or (layer0_outputs(1295));
    layer1_outputs(1344) <= not(layer0_outputs(1763));
    layer1_outputs(1345) <= not(layer0_outputs(2423)) or (layer0_outputs(647));
    layer1_outputs(1346) <= '1';
    layer1_outputs(1347) <= (layer0_outputs(718)) and (layer0_outputs(327));
    layer1_outputs(1348) <= layer0_outputs(2167);
    layer1_outputs(1349) <= layer0_outputs(2146);
    layer1_outputs(1350) <= '1';
    layer1_outputs(1351) <= not(layer0_outputs(1119));
    layer1_outputs(1352) <= (layer0_outputs(1937)) and (layer0_outputs(1395));
    layer1_outputs(1353) <= '1';
    layer1_outputs(1354) <= (layer0_outputs(1253)) xor (layer0_outputs(1303));
    layer1_outputs(1355) <= not(layer0_outputs(1695)) or (layer0_outputs(1570));
    layer1_outputs(1356) <= '1';
    layer1_outputs(1357) <= not(layer0_outputs(657)) or (layer0_outputs(10));
    layer1_outputs(1358) <= not(layer0_outputs(1446));
    layer1_outputs(1359) <= not(layer0_outputs(662)) or (layer0_outputs(1020));
    layer1_outputs(1360) <= not((layer0_outputs(185)) and (layer0_outputs(271)));
    layer1_outputs(1361) <= '1';
    layer1_outputs(1362) <= (layer0_outputs(2184)) and (layer0_outputs(2283));
    layer1_outputs(1363) <= (layer0_outputs(1927)) and not (layer0_outputs(2523));
    layer1_outputs(1364) <= layer0_outputs(1285);
    layer1_outputs(1365) <= (layer0_outputs(2375)) and not (layer0_outputs(1608));
    layer1_outputs(1366) <= '0';
    layer1_outputs(1367) <= not(layer0_outputs(227));
    layer1_outputs(1368) <= '1';
    layer1_outputs(1369) <= '0';
    layer1_outputs(1370) <= (layer0_outputs(2444)) or (layer0_outputs(16));
    layer1_outputs(1371) <= '0';
    layer1_outputs(1372) <= not(layer0_outputs(2047)) or (layer0_outputs(134));
    layer1_outputs(1373) <= layer0_outputs(259);
    layer1_outputs(1374) <= not((layer0_outputs(2517)) and (layer0_outputs(623)));
    layer1_outputs(1375) <= not(layer0_outputs(331));
    layer1_outputs(1376) <= not(layer0_outputs(1274));
    layer1_outputs(1377) <= not(layer0_outputs(967));
    layer1_outputs(1378) <= '0';
    layer1_outputs(1379) <= not(layer0_outputs(2389));
    layer1_outputs(1380) <= not(layer0_outputs(1632)) or (layer0_outputs(2036));
    layer1_outputs(1381) <= layer0_outputs(624);
    layer1_outputs(1382) <= layer0_outputs(515);
    layer1_outputs(1383) <= '0';
    layer1_outputs(1384) <= (layer0_outputs(1237)) and not (layer0_outputs(2299));
    layer1_outputs(1385) <= (layer0_outputs(1620)) and not (layer0_outputs(2219));
    layer1_outputs(1386) <= not(layer0_outputs(1670)) or (layer0_outputs(1686));
    layer1_outputs(1387) <= (layer0_outputs(100)) and not (layer0_outputs(433));
    layer1_outputs(1388) <= not(layer0_outputs(1197)) or (layer0_outputs(322));
    layer1_outputs(1389) <= layer0_outputs(1617);
    layer1_outputs(1390) <= '0';
    layer1_outputs(1391) <= not((layer0_outputs(955)) and (layer0_outputs(2331)));
    layer1_outputs(1392) <= not(layer0_outputs(1278)) or (layer0_outputs(2535));
    layer1_outputs(1393) <= (layer0_outputs(1224)) and (layer0_outputs(821));
    layer1_outputs(1394) <= not(layer0_outputs(1152));
    layer1_outputs(1395) <= layer0_outputs(487);
    layer1_outputs(1396) <= not(layer0_outputs(997)) or (layer0_outputs(366));
    layer1_outputs(1397) <= not(layer0_outputs(642));
    layer1_outputs(1398) <= not(layer0_outputs(772));
    layer1_outputs(1399) <= '0';
    layer1_outputs(1400) <= not(layer0_outputs(1611));
    layer1_outputs(1401) <= layer0_outputs(1759);
    layer1_outputs(1402) <= not((layer0_outputs(72)) and (layer0_outputs(1800)));
    layer1_outputs(1403) <= layer0_outputs(525);
    layer1_outputs(1404) <= (layer0_outputs(1148)) and not (layer0_outputs(154));
    layer1_outputs(1405) <= (layer0_outputs(1388)) or (layer0_outputs(209));
    layer1_outputs(1406) <= (layer0_outputs(596)) and not (layer0_outputs(2399));
    layer1_outputs(1407) <= (layer0_outputs(2016)) and not (layer0_outputs(1363));
    layer1_outputs(1408) <= not(layer0_outputs(196)) or (layer0_outputs(21));
    layer1_outputs(1409) <= not(layer0_outputs(1850)) or (layer0_outputs(484));
    layer1_outputs(1410) <= not(layer0_outputs(1326));
    layer1_outputs(1411) <= not(layer0_outputs(990)) or (layer0_outputs(176));
    layer1_outputs(1412) <= (layer0_outputs(2193)) or (layer0_outputs(1338));
    layer1_outputs(1413) <= layer0_outputs(1152);
    layer1_outputs(1414) <= not(layer0_outputs(2494)) or (layer0_outputs(1118));
    layer1_outputs(1415) <= not((layer0_outputs(1577)) xor (layer0_outputs(433)));
    layer1_outputs(1416) <= not(layer0_outputs(778));
    layer1_outputs(1417) <= not(layer0_outputs(370));
    layer1_outputs(1418) <= (layer0_outputs(2142)) or (layer0_outputs(450));
    layer1_outputs(1419) <= '0';
    layer1_outputs(1420) <= layer0_outputs(381);
    layer1_outputs(1421) <= '1';
    layer1_outputs(1422) <= (layer0_outputs(1331)) and not (layer0_outputs(1414));
    layer1_outputs(1423) <= not(layer0_outputs(1819));
    layer1_outputs(1424) <= layer0_outputs(320);
    layer1_outputs(1425) <= not(layer0_outputs(1659)) or (layer0_outputs(728));
    layer1_outputs(1426) <= not((layer0_outputs(1246)) and (layer0_outputs(1485)));
    layer1_outputs(1427) <= not((layer0_outputs(646)) and (layer0_outputs(1871)));
    layer1_outputs(1428) <= '0';
    layer1_outputs(1429) <= (layer0_outputs(65)) and not (layer0_outputs(1401));
    layer1_outputs(1430) <= '0';
    layer1_outputs(1431) <= (layer0_outputs(1449)) or (layer0_outputs(2137));
    layer1_outputs(1432) <= not(layer0_outputs(222)) or (layer0_outputs(85));
    layer1_outputs(1433) <= '0';
    layer1_outputs(1434) <= '1';
    layer1_outputs(1435) <= not(layer0_outputs(963)) or (layer0_outputs(933));
    layer1_outputs(1436) <= not(layer0_outputs(1917));
    layer1_outputs(1437) <= '0';
    layer1_outputs(1438) <= '0';
    layer1_outputs(1439) <= layer0_outputs(941);
    layer1_outputs(1440) <= layer0_outputs(714);
    layer1_outputs(1441) <= not(layer0_outputs(1495));
    layer1_outputs(1442) <= not(layer0_outputs(597)) or (layer0_outputs(251));
    layer1_outputs(1443) <= (layer0_outputs(2060)) or (layer0_outputs(1522));
    layer1_outputs(1444) <= (layer0_outputs(47)) or (layer0_outputs(1377));
    layer1_outputs(1445) <= '1';
    layer1_outputs(1446) <= '0';
    layer1_outputs(1447) <= not(layer0_outputs(1780));
    layer1_outputs(1448) <= layer0_outputs(1762);
    layer1_outputs(1449) <= '0';
    layer1_outputs(1450) <= not((layer0_outputs(1584)) and (layer0_outputs(438)));
    layer1_outputs(1451) <= (layer0_outputs(1139)) and not (layer0_outputs(515));
    layer1_outputs(1452) <= not((layer0_outputs(1328)) and (layer0_outputs(427)));
    layer1_outputs(1453) <= '1';
    layer1_outputs(1454) <= not(layer0_outputs(2454));
    layer1_outputs(1455) <= not(layer0_outputs(2008));
    layer1_outputs(1456) <= (layer0_outputs(917)) and not (layer0_outputs(1768));
    layer1_outputs(1457) <= (layer0_outputs(962)) and (layer0_outputs(120));
    layer1_outputs(1458) <= layer0_outputs(2038);
    layer1_outputs(1459) <= (layer0_outputs(1494)) and not (layer0_outputs(311));
    layer1_outputs(1460) <= not((layer0_outputs(1924)) and (layer0_outputs(338)));
    layer1_outputs(1461) <= (layer0_outputs(359)) or (layer0_outputs(658));
    layer1_outputs(1462) <= '1';
    layer1_outputs(1463) <= layer0_outputs(1202);
    layer1_outputs(1464) <= (layer0_outputs(2446)) or (layer0_outputs(711));
    layer1_outputs(1465) <= not(layer0_outputs(4));
    layer1_outputs(1466) <= '0';
    layer1_outputs(1467) <= (layer0_outputs(1545)) and not (layer0_outputs(1386));
    layer1_outputs(1468) <= '0';
    layer1_outputs(1469) <= not(layer0_outputs(2473));
    layer1_outputs(1470) <= not(layer0_outputs(400));
    layer1_outputs(1471) <= not((layer0_outputs(1552)) and (layer0_outputs(1721)));
    layer1_outputs(1472) <= (layer0_outputs(41)) and not (layer0_outputs(2416));
    layer1_outputs(1473) <= layer0_outputs(1484);
    layer1_outputs(1474) <= not(layer0_outputs(2135));
    layer1_outputs(1475) <= not(layer0_outputs(1739)) or (layer0_outputs(334));
    layer1_outputs(1476) <= not(layer0_outputs(60));
    layer1_outputs(1477) <= layer0_outputs(789);
    layer1_outputs(1478) <= not((layer0_outputs(1184)) or (layer0_outputs(639)));
    layer1_outputs(1479) <= not((layer0_outputs(725)) or (layer0_outputs(753)));
    layer1_outputs(1480) <= (layer0_outputs(1655)) and not (layer0_outputs(1426));
    layer1_outputs(1481) <= not((layer0_outputs(89)) or (layer0_outputs(2347)));
    layer1_outputs(1482) <= not((layer0_outputs(672)) or (layer0_outputs(1320)));
    layer1_outputs(1483) <= not((layer0_outputs(486)) and (layer0_outputs(2172)));
    layer1_outputs(1484) <= (layer0_outputs(518)) and not (layer0_outputs(578));
    layer1_outputs(1485) <= '0';
    layer1_outputs(1486) <= layer0_outputs(1042);
    layer1_outputs(1487) <= (layer0_outputs(1929)) and not (layer0_outputs(2319));
    layer1_outputs(1488) <= not(layer0_outputs(660)) or (layer0_outputs(506));
    layer1_outputs(1489) <= not(layer0_outputs(2230));
    layer1_outputs(1490) <= '0';
    layer1_outputs(1491) <= '0';
    layer1_outputs(1492) <= (layer0_outputs(277)) or (layer0_outputs(1958));
    layer1_outputs(1493) <= not((layer0_outputs(1391)) and (layer0_outputs(1612)));
    layer1_outputs(1494) <= '1';
    layer1_outputs(1495) <= not(layer0_outputs(1938));
    layer1_outputs(1496) <= not(layer0_outputs(1073));
    layer1_outputs(1497) <= not(layer0_outputs(461));
    layer1_outputs(1498) <= layer0_outputs(1836);
    layer1_outputs(1499) <= not(layer0_outputs(393)) or (layer0_outputs(1234));
    layer1_outputs(1500) <= (layer0_outputs(2175)) and not (layer0_outputs(1726));
    layer1_outputs(1501) <= (layer0_outputs(916)) or (layer0_outputs(1820));
    layer1_outputs(1502) <= '0';
    layer1_outputs(1503) <= '0';
    layer1_outputs(1504) <= not(layer0_outputs(1571));
    layer1_outputs(1505) <= '1';
    layer1_outputs(1506) <= (layer0_outputs(1438)) and (layer0_outputs(1318));
    layer1_outputs(1507) <= layer0_outputs(297);
    layer1_outputs(1508) <= (layer0_outputs(1778)) and not (layer0_outputs(1353));
    layer1_outputs(1509) <= (layer0_outputs(1321)) or (layer0_outputs(116));
    layer1_outputs(1510) <= (layer0_outputs(1096)) and (layer0_outputs(1439));
    layer1_outputs(1511) <= (layer0_outputs(2255)) and not (layer0_outputs(1450));
    layer1_outputs(1512) <= (layer0_outputs(2256)) or (layer0_outputs(441));
    layer1_outputs(1513) <= (layer0_outputs(1936)) and not (layer0_outputs(2505));
    layer1_outputs(1514) <= (layer0_outputs(454)) and not (layer0_outputs(1406));
    layer1_outputs(1515) <= not(layer0_outputs(884));
    layer1_outputs(1516) <= not(layer0_outputs(2192)) or (layer0_outputs(1053));
    layer1_outputs(1517) <= not((layer0_outputs(388)) or (layer0_outputs(283)));
    layer1_outputs(1518) <= '0';
    layer1_outputs(1519) <= '0';
    layer1_outputs(1520) <= (layer0_outputs(147)) and not (layer0_outputs(2468));
    layer1_outputs(1521) <= '1';
    layer1_outputs(1522) <= not(layer0_outputs(931));
    layer1_outputs(1523) <= '1';
    layer1_outputs(1524) <= layer0_outputs(1082);
    layer1_outputs(1525) <= (layer0_outputs(69)) and not (layer0_outputs(369));
    layer1_outputs(1526) <= (layer0_outputs(2430)) or (layer0_outputs(26));
    layer1_outputs(1527) <= not((layer0_outputs(1228)) or (layer0_outputs(2025)));
    layer1_outputs(1528) <= (layer0_outputs(2487)) and (layer0_outputs(1619));
    layer1_outputs(1529) <= '1';
    layer1_outputs(1530) <= (layer0_outputs(1872)) or (layer0_outputs(1747));
    layer1_outputs(1531) <= layer0_outputs(132);
    layer1_outputs(1532) <= not(layer0_outputs(1791)) or (layer0_outputs(1237));
    layer1_outputs(1533) <= '0';
    layer1_outputs(1534) <= '1';
    layer1_outputs(1535) <= layer0_outputs(199);
    layer1_outputs(1536) <= not(layer0_outputs(571));
    layer1_outputs(1537) <= (layer0_outputs(90)) and not (layer0_outputs(310));
    layer1_outputs(1538) <= not((layer0_outputs(1130)) or (layer0_outputs(1753)));
    layer1_outputs(1539) <= not(layer0_outputs(22)) or (layer0_outputs(254));
    layer1_outputs(1540) <= (layer0_outputs(2204)) and not (layer0_outputs(2098));
    layer1_outputs(1541) <= not((layer0_outputs(1509)) and (layer0_outputs(916)));
    layer1_outputs(1542) <= (layer0_outputs(775)) and not (layer0_outputs(307));
    layer1_outputs(1543) <= '1';
    layer1_outputs(1544) <= (layer0_outputs(1616)) or (layer0_outputs(626));
    layer1_outputs(1545) <= layer0_outputs(1942);
    layer1_outputs(1546) <= '0';
    layer1_outputs(1547) <= (layer0_outputs(1500)) and not (layer0_outputs(1839));
    layer1_outputs(1548) <= layer0_outputs(2249);
    layer1_outputs(1549) <= layer0_outputs(410);
    layer1_outputs(1550) <= not(layer0_outputs(100)) or (layer0_outputs(1080));
    layer1_outputs(1551) <= not((layer0_outputs(2239)) or (layer0_outputs(1311)));
    layer1_outputs(1552) <= layer0_outputs(717);
    layer1_outputs(1553) <= (layer0_outputs(480)) and not (layer0_outputs(1042));
    layer1_outputs(1554) <= layer0_outputs(940);
    layer1_outputs(1555) <= '1';
    layer1_outputs(1556) <= (layer0_outputs(903)) and not (layer0_outputs(1367));
    layer1_outputs(1557) <= (layer0_outputs(455)) or (layer0_outputs(2172));
    layer1_outputs(1558) <= not((layer0_outputs(2141)) or (layer0_outputs(319)));
    layer1_outputs(1559) <= (layer0_outputs(688)) and (layer0_outputs(2148));
    layer1_outputs(1560) <= (layer0_outputs(716)) xor (layer0_outputs(211));
    layer1_outputs(1561) <= (layer0_outputs(755)) and not (layer0_outputs(2288));
    layer1_outputs(1562) <= (layer0_outputs(744)) xor (layer0_outputs(1206));
    layer1_outputs(1563) <= layer0_outputs(2255);
    layer1_outputs(1564) <= not(layer0_outputs(1781)) or (layer0_outputs(470));
    layer1_outputs(1565) <= not(layer0_outputs(2328)) or (layer0_outputs(1135));
    layer1_outputs(1566) <= not(layer0_outputs(140)) or (layer0_outputs(1193));
    layer1_outputs(1567) <= (layer0_outputs(145)) xor (layer0_outputs(2070));
    layer1_outputs(1568) <= not(layer0_outputs(6));
    layer1_outputs(1569) <= not(layer0_outputs(1071)) or (layer0_outputs(568));
    layer1_outputs(1570) <= '1';
    layer1_outputs(1571) <= '1';
    layer1_outputs(1572) <= not(layer0_outputs(710));
    layer1_outputs(1573) <= not((layer0_outputs(962)) and (layer0_outputs(2402)));
    layer1_outputs(1574) <= not(layer0_outputs(1845));
    layer1_outputs(1575) <= (layer0_outputs(398)) and not (layer0_outputs(428));
    layer1_outputs(1576) <= (layer0_outputs(1482)) and not (layer0_outputs(476));
    layer1_outputs(1577) <= not(layer0_outputs(713)) or (layer0_outputs(2410));
    layer1_outputs(1578) <= (layer0_outputs(1189)) or (layer0_outputs(1128));
    layer1_outputs(1579) <= not(layer0_outputs(1007)) or (layer0_outputs(2221));
    layer1_outputs(1580) <= layer0_outputs(1818);
    layer1_outputs(1581) <= not(layer0_outputs(2538));
    layer1_outputs(1582) <= not(layer0_outputs(1100)) or (layer0_outputs(2449));
    layer1_outputs(1583) <= not(layer0_outputs(1354));
    layer1_outputs(1584) <= '1';
    layer1_outputs(1585) <= '0';
    layer1_outputs(1586) <= layer0_outputs(2218);
    layer1_outputs(1587) <= not(layer0_outputs(1047)) or (layer0_outputs(2420));
    layer1_outputs(1588) <= '0';
    layer1_outputs(1589) <= layer0_outputs(2166);
    layer1_outputs(1590) <= layer0_outputs(308);
    layer1_outputs(1591) <= '1';
    layer1_outputs(1592) <= '0';
    layer1_outputs(1593) <= (layer0_outputs(856)) or (layer0_outputs(1625));
    layer1_outputs(1594) <= not(layer0_outputs(1635));
    layer1_outputs(1595) <= not(layer0_outputs(522));
    layer1_outputs(1596) <= (layer0_outputs(33)) and not (layer0_outputs(826));
    layer1_outputs(1597) <= '1';
    layer1_outputs(1598) <= '1';
    layer1_outputs(1599) <= (layer0_outputs(1332)) and not (layer0_outputs(38));
    layer1_outputs(1600) <= layer0_outputs(1714);
    layer1_outputs(1601) <= not(layer0_outputs(221)) or (layer0_outputs(2277));
    layer1_outputs(1602) <= (layer0_outputs(1947)) and (layer0_outputs(2197));
    layer1_outputs(1603) <= '0';
    layer1_outputs(1604) <= layer0_outputs(1885);
    layer1_outputs(1605) <= not((layer0_outputs(1068)) and (layer0_outputs(2497)));
    layer1_outputs(1606) <= not(layer0_outputs(19)) or (layer0_outputs(518));
    layer1_outputs(1607) <= (layer0_outputs(1765)) and not (layer0_outputs(1192));
    layer1_outputs(1608) <= layer0_outputs(1035);
    layer1_outputs(1609) <= '0';
    layer1_outputs(1610) <= '0';
    layer1_outputs(1611) <= '0';
    layer1_outputs(1612) <= not(layer0_outputs(1531));
    layer1_outputs(1613) <= (layer0_outputs(1280)) and not (layer0_outputs(1807));
    layer1_outputs(1614) <= not(layer0_outputs(1943)) or (layer0_outputs(1043));
    layer1_outputs(1615) <= not(layer0_outputs(1533)) or (layer0_outputs(1460));
    layer1_outputs(1616) <= '0';
    layer1_outputs(1617) <= layer0_outputs(2231);
    layer1_outputs(1618) <= '0';
    layer1_outputs(1619) <= not(layer0_outputs(2291)) or (layer0_outputs(1317));
    layer1_outputs(1620) <= not(layer0_outputs(1913)) or (layer0_outputs(1341));
    layer1_outputs(1621) <= not(layer0_outputs(149)) or (layer0_outputs(2048));
    layer1_outputs(1622) <= not((layer0_outputs(1264)) and (layer0_outputs(1347)));
    layer1_outputs(1623) <= '1';
    layer1_outputs(1624) <= '1';
    layer1_outputs(1625) <= not(layer0_outputs(1592)) or (layer0_outputs(1011));
    layer1_outputs(1626) <= not(layer0_outputs(2349));
    layer1_outputs(1627) <= not(layer0_outputs(51));
    layer1_outputs(1628) <= '0';
    layer1_outputs(1629) <= not(layer0_outputs(868));
    layer1_outputs(1630) <= '0';
    layer1_outputs(1631) <= not((layer0_outputs(1581)) or (layer0_outputs(1497)));
    layer1_outputs(1632) <= layer0_outputs(1603);
    layer1_outputs(1633) <= (layer0_outputs(1948)) or (layer0_outputs(1717));
    layer1_outputs(1634) <= (layer0_outputs(2285)) and not (layer0_outputs(1811));
    layer1_outputs(1635) <= layer0_outputs(996);
    layer1_outputs(1636) <= not(layer0_outputs(1186));
    layer1_outputs(1637) <= not(layer0_outputs(1073));
    layer1_outputs(1638) <= layer0_outputs(1619);
    layer1_outputs(1639) <= (layer0_outputs(1891)) and (layer0_outputs(30));
    layer1_outputs(1640) <= layer0_outputs(39);
    layer1_outputs(1641) <= layer0_outputs(1780);
    layer1_outputs(1642) <= not((layer0_outputs(1027)) or (layer0_outputs(262)));
    layer1_outputs(1643) <= not(layer0_outputs(696)) or (layer0_outputs(2039));
    layer1_outputs(1644) <= not(layer0_outputs(1720)) or (layer0_outputs(1181));
    layer1_outputs(1645) <= not(layer0_outputs(2)) or (layer0_outputs(1486));
    layer1_outputs(1646) <= (layer0_outputs(2238)) or (layer0_outputs(1001));
    layer1_outputs(1647) <= not((layer0_outputs(685)) or (layer0_outputs(1934)));
    layer1_outputs(1648) <= layer0_outputs(1730);
    layer1_outputs(1649) <= '1';
    layer1_outputs(1650) <= not((layer0_outputs(1928)) or (layer0_outputs(2233)));
    layer1_outputs(1651) <= (layer0_outputs(2080)) and (layer0_outputs(2499));
    layer1_outputs(1652) <= layer0_outputs(74);
    layer1_outputs(1653) <= not((layer0_outputs(751)) or (layer0_outputs(117)));
    layer1_outputs(1654) <= not(layer0_outputs(1994));
    layer1_outputs(1655) <= not((layer0_outputs(2456)) and (layer0_outputs(1039)));
    layer1_outputs(1656) <= '1';
    layer1_outputs(1657) <= (layer0_outputs(75)) or (layer0_outputs(2069));
    layer1_outputs(1658) <= (layer0_outputs(1847)) or (layer0_outputs(1547));
    layer1_outputs(1659) <= not(layer0_outputs(1618)) or (layer0_outputs(1177));
    layer1_outputs(1660) <= layer0_outputs(1441);
    layer1_outputs(1661) <= not((layer0_outputs(362)) and (layer0_outputs(283)));
    layer1_outputs(1662) <= not(layer0_outputs(1226));
    layer1_outputs(1663) <= not(layer0_outputs(216)) or (layer0_outputs(2315));
    layer1_outputs(1664) <= layer0_outputs(1279);
    layer1_outputs(1665) <= not(layer0_outputs(2121));
    layer1_outputs(1666) <= (layer0_outputs(1842)) and (layer0_outputs(1683));
    layer1_outputs(1667) <= not((layer0_outputs(2409)) or (layer0_outputs(1474)));
    layer1_outputs(1668) <= (layer0_outputs(94)) and (layer0_outputs(444));
    layer1_outputs(1669) <= not(layer0_outputs(760)) or (layer0_outputs(1502));
    layer1_outputs(1670) <= layer0_outputs(543);
    layer1_outputs(1671) <= (layer0_outputs(1254)) and not (layer0_outputs(1524));
    layer1_outputs(1672) <= not((layer0_outputs(1080)) or (layer0_outputs(364)));
    layer1_outputs(1673) <= not(layer0_outputs(1824)) or (layer0_outputs(1607));
    layer1_outputs(1674) <= not(layer0_outputs(2195)) or (layer0_outputs(2199));
    layer1_outputs(1675) <= not(layer0_outputs(2318));
    layer1_outputs(1676) <= '1';
    layer1_outputs(1677) <= (layer0_outputs(1868)) and not (layer0_outputs(1116));
    layer1_outputs(1678) <= (layer0_outputs(747)) or (layer0_outputs(125));
    layer1_outputs(1679) <= not(layer0_outputs(964));
    layer1_outputs(1680) <= '1';
    layer1_outputs(1681) <= (layer0_outputs(519)) and not (layer0_outputs(2115));
    layer1_outputs(1682) <= '0';
    layer1_outputs(1683) <= '1';
    layer1_outputs(1684) <= '0';
    layer1_outputs(1685) <= '1';
    layer1_outputs(1686) <= not((layer0_outputs(805)) or (layer0_outputs(2139)));
    layer1_outputs(1687) <= not(layer0_outputs(1857)) or (layer0_outputs(2359));
    layer1_outputs(1688) <= '1';
    layer1_outputs(1689) <= not(layer0_outputs(1851)) or (layer0_outputs(1218));
    layer1_outputs(1690) <= (layer0_outputs(839)) and (layer0_outputs(1885));
    layer1_outputs(1691) <= (layer0_outputs(2155)) and not (layer0_outputs(1499));
    layer1_outputs(1692) <= not(layer0_outputs(111));
    layer1_outputs(1693) <= '1';
    layer1_outputs(1694) <= (layer0_outputs(110)) and not (layer0_outputs(740));
    layer1_outputs(1695) <= not(layer0_outputs(2252));
    layer1_outputs(1696) <= not((layer0_outputs(581)) or (layer0_outputs(2357)));
    layer1_outputs(1697) <= (layer0_outputs(429)) and not (layer0_outputs(2066));
    layer1_outputs(1698) <= (layer0_outputs(83)) or (layer0_outputs(715));
    layer1_outputs(1699) <= not(layer0_outputs(1269)) or (layer0_outputs(2292));
    layer1_outputs(1700) <= layer0_outputs(444);
    layer1_outputs(1701) <= '0';
    layer1_outputs(1702) <= '1';
    layer1_outputs(1703) <= layer0_outputs(560);
    layer1_outputs(1704) <= not(layer0_outputs(1056));
    layer1_outputs(1705) <= '1';
    layer1_outputs(1706) <= (layer0_outputs(1239)) and not (layer0_outputs(645));
    layer1_outputs(1707) <= not((layer0_outputs(365)) or (layer0_outputs(1038)));
    layer1_outputs(1708) <= (layer0_outputs(1232)) and not (layer0_outputs(2304));
    layer1_outputs(1709) <= '1';
    layer1_outputs(1710) <= layer0_outputs(2364);
    layer1_outputs(1711) <= layer0_outputs(1437);
    layer1_outputs(1712) <= not((layer0_outputs(1992)) and (layer0_outputs(1919)));
    layer1_outputs(1713) <= not(layer0_outputs(1651)) or (layer0_outputs(1261));
    layer1_outputs(1714) <= not((layer0_outputs(1822)) or (layer0_outputs(1011)));
    layer1_outputs(1715) <= '1';
    layer1_outputs(1716) <= not(layer0_outputs(1082)) or (layer0_outputs(855));
    layer1_outputs(1717) <= '0';
    layer1_outputs(1718) <= '0';
    layer1_outputs(1719) <= (layer0_outputs(1333)) and not (layer0_outputs(2181));
    layer1_outputs(1720) <= not(layer0_outputs(1973));
    layer1_outputs(1721) <= '0';
    layer1_outputs(1722) <= '0';
    layer1_outputs(1723) <= (layer0_outputs(400)) and not (layer0_outputs(2427));
    layer1_outputs(1724) <= '1';
    layer1_outputs(1725) <= (layer0_outputs(1788)) and not (layer0_outputs(92));
    layer1_outputs(1726) <= (layer0_outputs(1555)) and (layer0_outputs(2101));
    layer1_outputs(1727) <= (layer0_outputs(1397)) or (layer0_outputs(2525));
    layer1_outputs(1728) <= (layer0_outputs(2506)) and not (layer0_outputs(1498));
    layer1_outputs(1729) <= layer0_outputs(1437);
    layer1_outputs(1730) <= not(layer0_outputs(324));
    layer1_outputs(1731) <= not(layer0_outputs(1022)) or (layer0_outputs(1708));
    layer1_outputs(1732) <= (layer0_outputs(269)) and not (layer0_outputs(2547));
    layer1_outputs(1733) <= (layer0_outputs(1378)) and not (layer0_outputs(1318));
    layer1_outputs(1734) <= not(layer0_outputs(565)) or (layer0_outputs(1570));
    layer1_outputs(1735) <= '1';
    layer1_outputs(1736) <= not(layer0_outputs(1582));
    layer1_outputs(1737) <= (layer0_outputs(260)) or (layer0_outputs(2110));
    layer1_outputs(1738) <= not(layer0_outputs(1958));
    layer1_outputs(1739) <= not(layer0_outputs(1796)) or (layer0_outputs(77));
    layer1_outputs(1740) <= '0';
    layer1_outputs(1741) <= not((layer0_outputs(1255)) or (layer0_outputs(1808)));
    layer1_outputs(1742) <= layer0_outputs(743);
    layer1_outputs(1743) <= not(layer0_outputs(2085));
    layer1_outputs(1744) <= (layer0_outputs(1404)) or (layer0_outputs(2101));
    layer1_outputs(1745) <= '1';
    layer1_outputs(1746) <= not((layer0_outputs(2222)) and (layer0_outputs(991)));
    layer1_outputs(1747) <= not((layer0_outputs(203)) xor (layer0_outputs(1344)));
    layer1_outputs(1748) <= not((layer0_outputs(1001)) or (layer0_outputs(1333)));
    layer1_outputs(1749) <= not((layer0_outputs(527)) or (layer0_outputs(1022)));
    layer1_outputs(1750) <= not(layer0_outputs(1166)) or (layer0_outputs(2305));
    layer1_outputs(1751) <= (layer0_outputs(1414)) and not (layer0_outputs(1440));
    layer1_outputs(1752) <= not(layer0_outputs(1336));
    layer1_outputs(1753) <= '0';
    layer1_outputs(1754) <= not(layer0_outputs(53));
    layer1_outputs(1755) <= '1';
    layer1_outputs(1756) <= not(layer0_outputs(1629));
    layer1_outputs(1757) <= (layer0_outputs(306)) or (layer0_outputs(434));
    layer1_outputs(1758) <= (layer0_outputs(705)) and not (layer0_outputs(2125));
    layer1_outputs(1759) <= '1';
    layer1_outputs(1760) <= (layer0_outputs(140)) and not (layer0_outputs(2140));
    layer1_outputs(1761) <= not((layer0_outputs(1961)) or (layer0_outputs(1464)));
    layer1_outputs(1762) <= not(layer0_outputs(2411));
    layer1_outputs(1763) <= not(layer0_outputs(1387)) or (layer0_outputs(422));
    layer1_outputs(1764) <= not(layer0_outputs(2357));
    layer1_outputs(1765) <= not(layer0_outputs(1327));
    layer1_outputs(1766) <= not(layer0_outputs(2513)) or (layer0_outputs(24));
    layer1_outputs(1767) <= '0';
    layer1_outputs(1768) <= (layer0_outputs(208)) and (layer0_outputs(946));
    layer1_outputs(1769) <= layer0_outputs(1288);
    layer1_outputs(1770) <= (layer0_outputs(1429)) and (layer0_outputs(1963));
    layer1_outputs(1771) <= '1';
    layer1_outputs(1772) <= (layer0_outputs(129)) or (layer0_outputs(2190));
    layer1_outputs(1773) <= '0';
    layer1_outputs(1774) <= (layer0_outputs(2526)) and not (layer0_outputs(154));
    layer1_outputs(1775) <= (layer0_outputs(892)) or (layer0_outputs(1138));
    layer1_outputs(1776) <= not((layer0_outputs(2324)) or (layer0_outputs(93)));
    layer1_outputs(1777) <= not(layer0_outputs(650));
    layer1_outputs(1778) <= (layer0_outputs(457)) or (layer0_outputs(1417));
    layer1_outputs(1779) <= not(layer0_outputs(1890)) or (layer0_outputs(2483));
    layer1_outputs(1780) <= layer0_outputs(183);
    layer1_outputs(1781) <= not((layer0_outputs(2349)) or (layer0_outputs(240)));
    layer1_outputs(1782) <= (layer0_outputs(1767)) or (layer0_outputs(439));
    layer1_outputs(1783) <= layer0_outputs(1378);
    layer1_outputs(1784) <= not((layer0_outputs(1498)) or (layer0_outputs(2100)));
    layer1_outputs(1785) <= not((layer0_outputs(2518)) or (layer0_outputs(1688)));
    layer1_outputs(1786) <= (layer0_outputs(2405)) and not (layer0_outputs(2147));
    layer1_outputs(1787) <= '0';
    layer1_outputs(1788) <= '0';
    layer1_outputs(1789) <= (layer0_outputs(2324)) and not (layer0_outputs(1820));
    layer1_outputs(1790) <= not((layer0_outputs(554)) or (layer0_outputs(797)));
    layer1_outputs(1791) <= not(layer0_outputs(961)) or (layer0_outputs(850));
    layer1_outputs(1792) <= not(layer0_outputs(124));
    layer1_outputs(1793) <= not(layer0_outputs(193)) or (layer0_outputs(1149));
    layer1_outputs(1794) <= '1';
    layer1_outputs(1795) <= not((layer0_outputs(357)) and (layer0_outputs(1243)));
    layer1_outputs(1796) <= (layer0_outputs(2299)) and not (layer0_outputs(999));
    layer1_outputs(1797) <= layer0_outputs(1178);
    layer1_outputs(1798) <= not((layer0_outputs(1865)) and (layer0_outputs(914)));
    layer1_outputs(1799) <= layer0_outputs(304);
    layer1_outputs(1800) <= layer0_outputs(2241);
    layer1_outputs(1801) <= not(layer0_outputs(1072));
    layer1_outputs(1802) <= not(layer0_outputs(1422)) or (layer0_outputs(1709));
    layer1_outputs(1803) <= (layer0_outputs(1257)) and (layer0_outputs(918));
    layer1_outputs(1804) <= (layer0_outputs(1338)) and (layer0_outputs(1622));
    layer1_outputs(1805) <= '0';
    layer1_outputs(1806) <= '0';
    layer1_outputs(1807) <= (layer0_outputs(1597)) and not (layer0_outputs(1346));
    layer1_outputs(1808) <= (layer0_outputs(2044)) and (layer0_outputs(1915));
    layer1_outputs(1809) <= not((layer0_outputs(5)) or (layer0_outputs(476)));
    layer1_outputs(1810) <= not(layer0_outputs(1582)) or (layer0_outputs(2103));
    layer1_outputs(1811) <= (layer0_outputs(153)) and not (layer0_outputs(1912));
    layer1_outputs(1812) <= not(layer0_outputs(908)) or (layer0_outputs(946));
    layer1_outputs(1813) <= '1';
    layer1_outputs(1814) <= not(layer0_outputs(1139)) or (layer0_outputs(254));
    layer1_outputs(1815) <= not(layer0_outputs(2019));
    layer1_outputs(1816) <= layer0_outputs(640);
    layer1_outputs(1817) <= '0';
    layer1_outputs(1818) <= (layer0_outputs(2372)) and not (layer0_outputs(23));
    layer1_outputs(1819) <= (layer0_outputs(1058)) xor (layer0_outputs(1842));
    layer1_outputs(1820) <= '1';
    layer1_outputs(1821) <= (layer0_outputs(2328)) and not (layer0_outputs(2086));
    layer1_outputs(1822) <= '0';
    layer1_outputs(1823) <= not((layer0_outputs(44)) xor (layer0_outputs(2010)));
    layer1_outputs(1824) <= not(layer0_outputs(2534));
    layer1_outputs(1825) <= not(layer0_outputs(673)) or (layer0_outputs(1425));
    layer1_outputs(1826) <= layer0_outputs(1141);
    layer1_outputs(1827) <= not(layer0_outputs(1900)) or (layer0_outputs(1415));
    layer1_outputs(1828) <= not(layer0_outputs(25));
    layer1_outputs(1829) <= (layer0_outputs(1514)) and (layer0_outputs(2106));
    layer1_outputs(1830) <= layer0_outputs(1693);
    layer1_outputs(1831) <= (layer0_outputs(1496)) and (layer0_outputs(876));
    layer1_outputs(1832) <= not((layer0_outputs(945)) or (layer0_outputs(1978)));
    layer1_outputs(1833) <= layer0_outputs(1399);
    layer1_outputs(1834) <= '0';
    layer1_outputs(1835) <= layer0_outputs(1750);
    layer1_outputs(1836) <= not((layer0_outputs(2391)) and (layer0_outputs(2118)));
    layer1_outputs(1837) <= (layer0_outputs(1483)) and not (layer0_outputs(1340));
    layer1_outputs(1838) <= not(layer0_outputs(1495));
    layer1_outputs(1839) <= '0';
    layer1_outputs(1840) <= not(layer0_outputs(664)) or (layer0_outputs(1623));
    layer1_outputs(1841) <= not((layer0_outputs(1843)) and (layer0_outputs(1365)));
    layer1_outputs(1842) <= '0';
    layer1_outputs(1843) <= not(layer0_outputs(542)) or (layer0_outputs(1788));
    layer1_outputs(1844) <= (layer0_outputs(2488)) or (layer0_outputs(46));
    layer1_outputs(1845) <= (layer0_outputs(2419)) and (layer0_outputs(2437));
    layer1_outputs(1846) <= layer0_outputs(2210);
    layer1_outputs(1847) <= not(layer0_outputs(1372));
    layer1_outputs(1848) <= not(layer0_outputs(651));
    layer1_outputs(1849) <= not(layer0_outputs(1286));
    layer1_outputs(1850) <= not(layer0_outputs(1079));
    layer1_outputs(1851) <= '1';
    layer1_outputs(1852) <= not(layer0_outputs(1003)) or (layer0_outputs(59));
    layer1_outputs(1853) <= layer0_outputs(241);
    layer1_outputs(1854) <= not(layer0_outputs(726));
    layer1_outputs(1855) <= layer0_outputs(2325);
    layer1_outputs(1856) <= not((layer0_outputs(71)) and (layer0_outputs(231)));
    layer1_outputs(1857) <= not((layer0_outputs(1132)) and (layer0_outputs(1393)));
    layer1_outputs(1858) <= (layer0_outputs(732)) and not (layer0_outputs(2482));
    layer1_outputs(1859) <= not(layer0_outputs(1693));
    layer1_outputs(1860) <= not(layer0_outputs(163)) or (layer0_outputs(1250));
    layer1_outputs(1861) <= '1';
    layer1_outputs(1862) <= '0';
    layer1_outputs(1863) <= layer0_outputs(2278);
    layer1_outputs(1864) <= '0';
    layer1_outputs(1865) <= layer0_outputs(2142);
    layer1_outputs(1866) <= (layer0_outputs(1863)) and not (layer0_outputs(773));
    layer1_outputs(1867) <= layer0_outputs(1480);
    layer1_outputs(1868) <= not(layer0_outputs(756)) or (layer0_outputs(2554));
    layer1_outputs(1869) <= '1';
    layer1_outputs(1870) <= '1';
    layer1_outputs(1871) <= not(layer0_outputs(1420));
    layer1_outputs(1872) <= '0';
    layer1_outputs(1873) <= not((layer0_outputs(1397)) or (layer0_outputs(1998)));
    layer1_outputs(1874) <= not(layer0_outputs(1530)) or (layer0_outputs(2182));
    layer1_outputs(1875) <= '1';
    layer1_outputs(1876) <= not((layer0_outputs(1432)) and (layer0_outputs(1931)));
    layer1_outputs(1877) <= layer0_outputs(794);
    layer1_outputs(1878) <= (layer0_outputs(1946)) and not (layer0_outputs(1939));
    layer1_outputs(1879) <= '1';
    layer1_outputs(1880) <= not((layer0_outputs(232)) and (layer0_outputs(484)));
    layer1_outputs(1881) <= layer0_outputs(2058);
    layer1_outputs(1882) <= not(layer0_outputs(1032)) or (layer0_outputs(416));
    layer1_outputs(1883) <= '0';
    layer1_outputs(1884) <= not(layer0_outputs(840));
    layer1_outputs(1885) <= (layer0_outputs(1191)) xor (layer0_outputs(43));
    layer1_outputs(1886) <= layer0_outputs(1182);
    layer1_outputs(1887) <= not((layer0_outputs(1030)) or (layer0_outputs(754)));
    layer1_outputs(1888) <= layer0_outputs(1375);
    layer1_outputs(1889) <= not((layer0_outputs(344)) and (layer0_outputs(2023)));
    layer1_outputs(1890) <= '0';
    layer1_outputs(1891) <= not((layer0_outputs(2386)) and (layer0_outputs(2478)));
    layer1_outputs(1892) <= '0';
    layer1_outputs(1893) <= not(layer0_outputs(438)) or (layer0_outputs(430));
    layer1_outputs(1894) <= not(layer0_outputs(625)) or (layer0_outputs(632));
    layer1_outputs(1895) <= '1';
    layer1_outputs(1896) <= '1';
    layer1_outputs(1897) <= '0';
    layer1_outputs(1898) <= not((layer0_outputs(2371)) and (layer0_outputs(1704)));
    layer1_outputs(1899) <= '1';
    layer1_outputs(1900) <= not(layer0_outputs(290)) or (layer0_outputs(1723));
    layer1_outputs(1901) <= (layer0_outputs(2254)) and (layer0_outputs(1931));
    layer1_outputs(1902) <= not(layer0_outputs(524));
    layer1_outputs(1903) <= not(layer0_outputs(1704));
    layer1_outputs(1904) <= not(layer0_outputs(430));
    layer1_outputs(1905) <= '1';
    layer1_outputs(1906) <= not((layer0_outputs(678)) and (layer0_outputs(596)));
    layer1_outputs(1907) <= not((layer0_outputs(599)) and (layer0_outputs(1823)));
    layer1_outputs(1908) <= not((layer0_outputs(5)) and (layer0_outputs(2476)));
    layer1_outputs(1909) <= layer0_outputs(612);
    layer1_outputs(1910) <= not(layer0_outputs(1835)) or (layer0_outputs(2465));
    layer1_outputs(1911) <= not(layer0_outputs(1263)) or (layer0_outputs(1903));
    layer1_outputs(1912) <= not((layer0_outputs(1818)) and (layer0_outputs(1348)));
    layer1_outputs(1913) <= (layer0_outputs(1370)) and (layer0_outputs(1119));
    layer1_outputs(1914) <= '1';
    layer1_outputs(1915) <= '1';
    layer1_outputs(1916) <= not((layer0_outputs(807)) and (layer0_outputs(1559)));
    layer1_outputs(1917) <= (layer0_outputs(2071)) or (layer0_outputs(1083));
    layer1_outputs(1918) <= layer0_outputs(110);
    layer1_outputs(1919) <= '1';
    layer1_outputs(1920) <= '0';
    layer1_outputs(1921) <= layer0_outputs(794);
    layer1_outputs(1922) <= not((layer0_outputs(857)) and (layer0_outputs(1557)));
    layer1_outputs(1923) <= not(layer0_outputs(2165));
    layer1_outputs(1924) <= not(layer0_outputs(348)) or (layer0_outputs(442));
    layer1_outputs(1925) <= '0';
    layer1_outputs(1926) <= not((layer0_outputs(169)) and (layer0_outputs(1247)));
    layer1_outputs(1927) <= '1';
    layer1_outputs(1928) <= '0';
    layer1_outputs(1929) <= (layer0_outputs(2002)) and (layer0_outputs(1781));
    layer1_outputs(1930) <= '1';
    layer1_outputs(1931) <= (layer0_outputs(1522)) xor (layer0_outputs(1728));
    layer1_outputs(1932) <= (layer0_outputs(245)) or (layer0_outputs(963));
    layer1_outputs(1933) <= (layer0_outputs(2012)) or (layer0_outputs(1259));
    layer1_outputs(1934) <= (layer0_outputs(1669)) and not (layer0_outputs(2188));
    layer1_outputs(1935) <= '0';
    layer1_outputs(1936) <= (layer0_outputs(62)) and not (layer0_outputs(957));
    layer1_outputs(1937) <= not(layer0_outputs(1256)) or (layer0_outputs(1758));
    layer1_outputs(1938) <= not(layer0_outputs(179));
    layer1_outputs(1939) <= layer0_outputs(1860);
    layer1_outputs(1940) <= not((layer0_outputs(2133)) and (layer0_outputs(964)));
    layer1_outputs(1941) <= (layer0_outputs(1826)) and (layer0_outputs(301));
    layer1_outputs(1942) <= not(layer0_outputs(1097));
    layer1_outputs(1943) <= (layer0_outputs(2546)) and not (layer0_outputs(1516));
    layer1_outputs(1944) <= (layer0_outputs(1021)) and not (layer0_outputs(2284));
    layer1_outputs(1945) <= (layer0_outputs(978)) and not (layer0_outputs(1411));
    layer1_outputs(1946) <= not((layer0_outputs(298)) and (layer0_outputs(1841)));
    layer1_outputs(1947) <= not(layer0_outputs(1272));
    layer1_outputs(1948) <= layer0_outputs(2395);
    layer1_outputs(1949) <= not((layer0_outputs(13)) or (layer0_outputs(560)));
    layer1_outputs(1950) <= not(layer0_outputs(1718));
    layer1_outputs(1951) <= (layer0_outputs(2440)) or (layer0_outputs(1455));
    layer1_outputs(1952) <= not(layer0_outputs(2146)) or (layer0_outputs(1519));
    layer1_outputs(1953) <= not((layer0_outputs(1641)) and (layer0_outputs(2207)));
    layer1_outputs(1954) <= not((layer0_outputs(744)) or (layer0_outputs(1213)));
    layer1_outputs(1955) <= layer0_outputs(1748);
    layer1_outputs(1956) <= '1';
    layer1_outputs(1957) <= '0';
    layer1_outputs(1958) <= not(layer0_outputs(2014)) or (layer0_outputs(680));
    layer1_outputs(1959) <= not(layer0_outputs(1643));
    layer1_outputs(1960) <= not(layer0_outputs(801));
    layer1_outputs(1961) <= '1';
    layer1_outputs(1962) <= (layer0_outputs(1434)) or (layer0_outputs(630));
    layer1_outputs(1963) <= not(layer0_outputs(1361));
    layer1_outputs(1964) <= not(layer0_outputs(442));
    layer1_outputs(1965) <= (layer0_outputs(745)) and not (layer0_outputs(314));
    layer1_outputs(1966) <= layer0_outputs(436);
    layer1_outputs(1967) <= (layer0_outputs(2379)) and not (layer0_outputs(1552));
    layer1_outputs(1968) <= '0';
    layer1_outputs(1969) <= not(layer0_outputs(1510)) or (layer0_outputs(1571));
    layer1_outputs(1970) <= not(layer0_outputs(1898)) or (layer0_outputs(1203));
    layer1_outputs(1971) <= layer0_outputs(763);
    layer1_outputs(1972) <= (layer0_outputs(2205)) or (layer0_outputs(146));
    layer1_outputs(1973) <= not(layer0_outputs(1491)) or (layer0_outputs(1767));
    layer1_outputs(1974) <= (layer0_outputs(197)) and not (layer0_outputs(274));
    layer1_outputs(1975) <= (layer0_outputs(1409)) and (layer0_outputs(113));
    layer1_outputs(1976) <= not(layer0_outputs(864)) or (layer0_outputs(1581));
    layer1_outputs(1977) <= layer0_outputs(924);
    layer1_outputs(1978) <= (layer0_outputs(99)) xor (layer0_outputs(2463));
    layer1_outputs(1979) <= not(layer0_outputs(802));
    layer1_outputs(1980) <= (layer0_outputs(1056)) and (layer0_outputs(1178));
    layer1_outputs(1981) <= not(layer0_outputs(742));
    layer1_outputs(1982) <= layer0_outputs(46);
    layer1_outputs(1983) <= not(layer0_outputs(707)) or (layer0_outputs(2260));
    layer1_outputs(1984) <= '0';
    layer1_outputs(1985) <= '0';
    layer1_outputs(1986) <= not((layer0_outputs(2187)) or (layer0_outputs(643)));
    layer1_outputs(1987) <= '0';
    layer1_outputs(1988) <= layer0_outputs(2257);
    layer1_outputs(1989) <= (layer0_outputs(2475)) and not (layer0_outputs(1527));
    layer1_outputs(1990) <= '0';
    layer1_outputs(1991) <= not(layer0_outputs(1987)) or (layer0_outputs(1055));
    layer1_outputs(1992) <= (layer0_outputs(496)) and not (layer0_outputs(2224));
    layer1_outputs(1993) <= not(layer0_outputs(1993));
    layer1_outputs(1994) <= not(layer0_outputs(814));
    layer1_outputs(1995) <= not((layer0_outputs(748)) or (layer0_outputs(645)));
    layer1_outputs(1996) <= not((layer0_outputs(2102)) and (layer0_outputs(356)));
    layer1_outputs(1997) <= (layer0_outputs(1729)) and not (layer0_outputs(782));
    layer1_outputs(1998) <= not(layer0_outputs(1997));
    layer1_outputs(1999) <= not((layer0_outputs(2275)) or (layer0_outputs(1645)));
    layer1_outputs(2000) <= layer0_outputs(2443);
    layer1_outputs(2001) <= layer0_outputs(1824);
    layer1_outputs(2002) <= not(layer0_outputs(981));
    layer1_outputs(2003) <= layer0_outputs(1126);
    layer1_outputs(2004) <= (layer0_outputs(942)) and not (layer0_outputs(1342));
    layer1_outputs(2005) <= not(layer0_outputs(119)) or (layer0_outputs(578));
    layer1_outputs(2006) <= not((layer0_outputs(1291)) and (layer0_outputs(2345)));
    layer1_outputs(2007) <= '0';
    layer1_outputs(2008) <= layer0_outputs(2397);
    layer1_outputs(2009) <= '1';
    layer1_outputs(2010) <= '0';
    layer1_outputs(2011) <= (layer0_outputs(1708)) or (layer0_outputs(1725));
    layer1_outputs(2012) <= not(layer0_outputs(1965));
    layer1_outputs(2013) <= layer0_outputs(239);
    layer1_outputs(2014) <= not(layer0_outputs(928));
    layer1_outputs(2015) <= not(layer0_outputs(491));
    layer1_outputs(2016) <= (layer0_outputs(1183)) or (layer0_outputs(2555));
    layer1_outputs(2017) <= '1';
    layer1_outputs(2018) <= layer0_outputs(1583);
    layer1_outputs(2019) <= (layer0_outputs(2326)) and (layer0_outputs(871));
    layer1_outputs(2020) <= (layer0_outputs(431)) and not (layer0_outputs(866));
    layer1_outputs(2021) <= layer0_outputs(1419);
    layer1_outputs(2022) <= not(layer0_outputs(516)) or (layer0_outputs(495));
    layer1_outputs(2023) <= (layer0_outputs(206)) or (layer0_outputs(437));
    layer1_outputs(2024) <= (layer0_outputs(1280)) and not (layer0_outputs(2510));
    layer1_outputs(2025) <= not(layer0_outputs(2191)) or (layer0_outputs(351));
    layer1_outputs(2026) <= '0';
    layer1_outputs(2027) <= '0';
    layer1_outputs(2028) <= (layer0_outputs(1362)) or (layer0_outputs(759));
    layer1_outputs(2029) <= not(layer0_outputs(2076));
    layer1_outputs(2030) <= layer0_outputs(2434);
    layer1_outputs(2031) <= '1';
    layer1_outputs(2032) <= not(layer0_outputs(2363)) or (layer0_outputs(594));
    layer1_outputs(2033) <= '0';
    layer1_outputs(2034) <= not(layer0_outputs(1895));
    layer1_outputs(2035) <= '1';
    layer1_outputs(2036) <= '1';
    layer1_outputs(2037) <= (layer0_outputs(2217)) and not (layer0_outputs(2425));
    layer1_outputs(2038) <= (layer0_outputs(1464)) and (layer0_outputs(598));
    layer1_outputs(2039) <= not((layer0_outputs(2140)) or (layer0_outputs(155)));
    layer1_outputs(2040) <= (layer0_outputs(434)) or (layer0_outputs(1460));
    layer1_outputs(2041) <= not(layer0_outputs(435));
    layer1_outputs(2042) <= not(layer0_outputs(1098)) or (layer0_outputs(2267));
    layer1_outputs(2043) <= layer0_outputs(657);
    layer1_outputs(2044) <= '1';
    layer1_outputs(2045) <= not(layer0_outputs(1550)) or (layer0_outputs(2031));
    layer1_outputs(2046) <= layer0_outputs(1158);
    layer1_outputs(2047) <= '0';
    layer1_outputs(2048) <= (layer0_outputs(151)) and (layer0_outputs(1757));
    layer1_outputs(2049) <= layer0_outputs(2484);
    layer1_outputs(2050) <= not(layer0_outputs(1383)) or (layer0_outputs(2469));
    layer1_outputs(2051) <= not((layer0_outputs(2259)) and (layer0_outputs(611)));
    layer1_outputs(2052) <= '1';
    layer1_outputs(2053) <= (layer0_outputs(2485)) and not (layer0_outputs(2498));
    layer1_outputs(2054) <= not(layer0_outputs(463));
    layer1_outputs(2055) <= '0';
    layer1_outputs(2056) <= not(layer0_outputs(953));
    layer1_outputs(2057) <= not((layer0_outputs(1164)) or (layer0_outputs(1339)));
    layer1_outputs(2058) <= not(layer0_outputs(1013));
    layer1_outputs(2059) <= not((layer0_outputs(1418)) or (layer0_outputs(2353)));
    layer1_outputs(2060) <= (layer0_outputs(2358)) and not (layer0_outputs(289));
    layer1_outputs(2061) <= layer0_outputs(1957);
    layer1_outputs(2062) <= layer0_outputs(2290);
    layer1_outputs(2063) <= layer0_outputs(2382);
    layer1_outputs(2064) <= '0';
    layer1_outputs(2065) <= not(layer0_outputs(1093));
    layer1_outputs(2066) <= layer0_outputs(815);
    layer1_outputs(2067) <= layer0_outputs(1258);
    layer1_outputs(2068) <= layer0_outputs(658);
    layer1_outputs(2069) <= layer0_outputs(1266);
    layer1_outputs(2070) <= not(layer0_outputs(1960));
    layer1_outputs(2071) <= not(layer0_outputs(493)) or (layer0_outputs(9));
    layer1_outputs(2072) <= (layer0_outputs(816)) and (layer0_outputs(1795));
    layer1_outputs(2073) <= not(layer0_outputs(412)) or (layer0_outputs(2174));
    layer1_outputs(2074) <= (layer0_outputs(2448)) and (layer0_outputs(278));
    layer1_outputs(2075) <= not(layer0_outputs(1910)) or (layer0_outputs(249));
    layer1_outputs(2076) <= not(layer0_outputs(694));
    layer1_outputs(2077) <= not(layer0_outputs(20));
    layer1_outputs(2078) <= '1';
    layer1_outputs(2079) <= not(layer0_outputs(834)) or (layer0_outputs(877));
    layer1_outputs(2080) <= not(layer0_outputs(1564)) or (layer0_outputs(1249));
    layer1_outputs(2081) <= '1';
    layer1_outputs(2082) <= (layer0_outputs(712)) or (layer0_outputs(342));
    layer1_outputs(2083) <= '0';
    layer1_outputs(2084) <= not(layer0_outputs(513)) or (layer0_outputs(1834));
    layer1_outputs(2085) <= layer0_outputs(1266);
    layer1_outputs(2086) <= not(layer0_outputs(1141)) or (layer0_outputs(562));
    layer1_outputs(2087) <= not(layer0_outputs(2505));
    layer1_outputs(2088) <= layer0_outputs(1545);
    layer1_outputs(2089) <= not(layer0_outputs(1650));
    layer1_outputs(2090) <= layer0_outputs(627);
    layer1_outputs(2091) <= not((layer0_outputs(446)) xor (layer0_outputs(1759)));
    layer1_outputs(2092) <= not(layer0_outputs(1539));
    layer1_outputs(2093) <= layer0_outputs(604);
    layer1_outputs(2094) <= (layer0_outputs(1779)) xor (layer0_outputs(1894));
    layer1_outputs(2095) <= (layer0_outputs(1474)) and (layer0_outputs(2260));
    layer1_outputs(2096) <= not((layer0_outputs(948)) or (layer0_outputs(1008)));
    layer1_outputs(2097) <= (layer0_outputs(811)) and (layer0_outputs(1892));
    layer1_outputs(2098) <= (layer0_outputs(2015)) and not (layer0_outputs(788));
    layer1_outputs(2099) <= not((layer0_outputs(1952)) or (layer0_outputs(448)));
    layer1_outputs(2100) <= '1';
    layer1_outputs(2101) <= layer0_outputs(1492);
    layer1_outputs(2102) <= not(layer0_outputs(417)) or (layer0_outputs(1903));
    layer1_outputs(2103) <= not(layer0_outputs(230));
    layer1_outputs(2104) <= (layer0_outputs(708)) xor (layer0_outputs(1949));
    layer1_outputs(2105) <= (layer0_outputs(77)) and not (layer0_outputs(1753));
    layer1_outputs(2106) <= not((layer0_outputs(1856)) and (layer0_outputs(2346)));
    layer1_outputs(2107) <= not(layer0_outputs(2161));
    layer1_outputs(2108) <= not(layer0_outputs(56));
    layer1_outputs(2109) <= '1';
    layer1_outputs(2110) <= '1';
    layer1_outputs(2111) <= (layer0_outputs(2312)) and not (layer0_outputs(2185));
    layer1_outputs(2112) <= not(layer0_outputs(2389));
    layer1_outputs(2113) <= (layer0_outputs(261)) or (layer0_outputs(1165));
    layer1_outputs(2114) <= not(layer0_outputs(2206));
    layer1_outputs(2115) <= not(layer0_outputs(546));
    layer1_outputs(2116) <= (layer0_outputs(1999)) or (layer0_outputs(1095));
    layer1_outputs(2117) <= (layer0_outputs(1535)) or (layer0_outputs(2109));
    layer1_outputs(2118) <= '1';
    layer1_outputs(2119) <= '0';
    layer1_outputs(2120) <= '1';
    layer1_outputs(2121) <= not(layer0_outputs(525));
    layer1_outputs(2122) <= '0';
    layer1_outputs(2123) <= not(layer0_outputs(1578)) or (layer0_outputs(947));
    layer1_outputs(2124) <= not(layer0_outputs(194)) or (layer0_outputs(2333));
    layer1_outputs(2125) <= not((layer0_outputs(1270)) and (layer0_outputs(2297)));
    layer1_outputs(2126) <= '1';
    layer1_outputs(2127) <= not(layer0_outputs(1060)) or (layer0_outputs(667));
    layer1_outputs(2128) <= (layer0_outputs(1104)) and not (layer0_outputs(1200));
    layer1_outputs(2129) <= '0';
    layer1_outputs(2130) <= '0';
    layer1_outputs(2131) <= '1';
    layer1_outputs(2132) <= '1';
    layer1_outputs(2133) <= (layer0_outputs(1335)) xor (layer0_outputs(2105));
    layer1_outputs(2134) <= not(layer0_outputs(2352)) or (layer0_outputs(819));
    layer1_outputs(2135) <= not((layer0_outputs(1808)) and (layer0_outputs(888)));
    layer1_outputs(2136) <= '1';
    layer1_outputs(2137) <= '1';
    layer1_outputs(2138) <= not(layer0_outputs(1502));
    layer1_outputs(2139) <= (layer0_outputs(2037)) and not (layer0_outputs(103));
    layer1_outputs(2140) <= (layer0_outputs(1278)) and not (layer0_outputs(1537));
    layer1_outputs(2141) <= (layer0_outputs(14)) and (layer0_outputs(2134));
    layer1_outputs(2142) <= not((layer0_outputs(555)) and (layer0_outputs(1207)));
    layer1_outputs(2143) <= not(layer0_outputs(2499));
    layer1_outputs(2144) <= '0';
    layer1_outputs(2145) <= (layer0_outputs(2338)) or (layer0_outputs(989));
    layer1_outputs(2146) <= (layer0_outputs(1629)) or (layer0_outputs(1519));
    layer1_outputs(2147) <= (layer0_outputs(1433)) xor (layer0_outputs(1112));
    layer1_outputs(2148) <= not(layer0_outputs(2120));
    layer1_outputs(2149) <= '1';
    layer1_outputs(2150) <= '1';
    layer1_outputs(2151) <= '1';
    layer1_outputs(2152) <= (layer0_outputs(1200)) xor (layer0_outputs(1322));
    layer1_outputs(2153) <= not((layer0_outputs(1762)) and (layer0_outputs(1206)));
    layer1_outputs(2154) <= '0';
    layer1_outputs(2155) <= not((layer0_outputs(548)) or (layer0_outputs(56)));
    layer1_outputs(2156) <= (layer0_outputs(947)) or (layer0_outputs(1567));
    layer1_outputs(2157) <= not(layer0_outputs(2517)) or (layer0_outputs(606));
    layer1_outputs(2158) <= layer0_outputs(1902);
    layer1_outputs(2159) <= layer0_outputs(1476);
    layer1_outputs(2160) <= not((layer0_outputs(1614)) and (layer0_outputs(2540)));
    layer1_outputs(2161) <= layer0_outputs(2366);
    layer1_outputs(2162) <= '1';
    layer1_outputs(2163) <= layer0_outputs(2033);
    layer1_outputs(2164) <= '1';
    layer1_outputs(2165) <= '0';
    layer1_outputs(2166) <= not(layer0_outputs(494));
    layer1_outputs(2167) <= not((layer0_outputs(2164)) or (layer0_outputs(1155)));
    layer1_outputs(2168) <= '0';
    layer1_outputs(2169) <= not(layer0_outputs(1330)) or (layer0_outputs(2115));
    layer1_outputs(2170) <= layer0_outputs(629);
    layer1_outputs(2171) <= not(layer0_outputs(746));
    layer1_outputs(2172) <= (layer0_outputs(1164)) and (layer0_outputs(1558));
    layer1_outputs(2173) <= (layer0_outputs(723)) or (layer0_outputs(2111));
    layer1_outputs(2174) <= (layer0_outputs(874)) and not (layer0_outputs(2438));
    layer1_outputs(2175) <= not((layer0_outputs(32)) or (layer0_outputs(1872)));
    layer1_outputs(2176) <= layer0_outputs(936);
    layer1_outputs(2177) <= not((layer0_outputs(1626)) and (layer0_outputs(2051)));
    layer1_outputs(2178) <= not(layer0_outputs(192));
    layer1_outputs(2179) <= (layer0_outputs(2376)) and not (layer0_outputs(2027));
    layer1_outputs(2180) <= (layer0_outputs(464)) and (layer0_outputs(452));
    layer1_outputs(2181) <= layer0_outputs(2541);
    layer1_outputs(2182) <= (layer0_outputs(765)) and not (layer0_outputs(2539));
    layer1_outputs(2183) <= (layer0_outputs(1092)) and (layer0_outputs(918));
    layer1_outputs(2184) <= (layer0_outputs(977)) and not (layer0_outputs(2419));
    layer1_outputs(2185) <= not(layer0_outputs(2108));
    layer1_outputs(2186) <= '1';
    layer1_outputs(2187) <= (layer0_outputs(1111)) and (layer0_outputs(1270));
    layer1_outputs(2188) <= '1';
    layer1_outputs(2189) <= not((layer0_outputs(6)) or (layer0_outputs(2084)));
    layer1_outputs(2190) <= layer0_outputs(34);
    layer1_outputs(2191) <= not(layer0_outputs(94));
    layer1_outputs(2192) <= not(layer0_outputs(149));
    layer1_outputs(2193) <= not(layer0_outputs(432)) or (layer0_outputs(1642));
    layer1_outputs(2194) <= (layer0_outputs(766)) and not (layer0_outputs(1356));
    layer1_outputs(2195) <= (layer0_outputs(424)) and not (layer0_outputs(396));
    layer1_outputs(2196) <= layer0_outputs(2073);
    layer1_outputs(2197) <= layer0_outputs(53);
    layer1_outputs(2198) <= (layer0_outputs(679)) or (layer0_outputs(2227));
    layer1_outputs(2199) <= '0';
    layer1_outputs(2200) <= '1';
    layer1_outputs(2201) <= '1';
    layer1_outputs(2202) <= not((layer0_outputs(328)) and (layer0_outputs(2072)));
    layer1_outputs(2203) <= (layer0_outputs(2176)) and (layer0_outputs(419));
    layer1_outputs(2204) <= not(layer0_outputs(1713)) or (layer0_outputs(402));
    layer1_outputs(2205) <= layer0_outputs(2432);
    layer1_outputs(2206) <= not(layer0_outputs(2264)) or (layer0_outputs(2136));
    layer1_outputs(2207) <= (layer0_outputs(933)) or (layer0_outputs(2362));
    layer1_outputs(2208) <= (layer0_outputs(1628)) and (layer0_outputs(1439));
    layer1_outputs(2209) <= (layer0_outputs(1373)) and not (layer0_outputs(1816));
    layer1_outputs(2210) <= (layer0_outputs(1067)) and not (layer0_outputs(654));
    layer1_outputs(2211) <= layer0_outputs(1109);
    layer1_outputs(2212) <= '0';
    layer1_outputs(2213) <= not(layer0_outputs(2001));
    layer1_outputs(2214) <= '0';
    layer1_outputs(2215) <= not((layer0_outputs(1671)) or (layer0_outputs(307)));
    layer1_outputs(2216) <= layer0_outputs(1161);
    layer1_outputs(2217) <= '0';
    layer1_outputs(2218) <= (layer0_outputs(483)) and not (layer0_outputs(609));
    layer1_outputs(2219) <= (layer0_outputs(1514)) and not (layer0_outputs(2527));
    layer1_outputs(2220) <= not(layer0_outputs(1526));
    layer1_outputs(2221) <= not((layer0_outputs(1335)) or (layer0_outputs(321)));
    layer1_outputs(2222) <= layer0_outputs(1311);
    layer1_outputs(2223) <= not((layer0_outputs(2540)) or (layer0_outputs(1540)));
    layer1_outputs(2224) <= (layer0_outputs(938)) and (layer0_outputs(1648));
    layer1_outputs(2225) <= layer0_outputs(1490);
    layer1_outputs(2226) <= '0';
    layer1_outputs(2227) <= '0';
    layer1_outputs(2228) <= '0';
    layer1_outputs(2229) <= not((layer0_outputs(1933)) or (layer0_outputs(603)));
    layer1_outputs(2230) <= '1';
    layer1_outputs(2231) <= not((layer0_outputs(1262)) or (layer0_outputs(724)));
    layer1_outputs(2232) <= '0';
    layer1_outputs(2233) <= not((layer0_outputs(2083)) or (layer0_outputs(500)));
    layer1_outputs(2234) <= not(layer0_outputs(1064));
    layer1_outputs(2235) <= (layer0_outputs(1636)) and not (layer0_outputs(1016));
    layer1_outputs(2236) <= (layer0_outputs(1573)) and not (layer0_outputs(2006));
    layer1_outputs(2237) <= '0';
    layer1_outputs(2238) <= '1';
    layer1_outputs(2239) <= '0';
    layer1_outputs(2240) <= not(layer0_outputs(1061));
    layer1_outputs(2241) <= (layer0_outputs(1711)) or (layer0_outputs(1257));
    layer1_outputs(2242) <= not(layer0_outputs(1169)) or (layer0_outputs(776));
    layer1_outputs(2243) <= '0';
    layer1_outputs(2244) <= '1';
    layer1_outputs(2245) <= '0';
    layer1_outputs(2246) <= not(layer0_outputs(848));
    layer1_outputs(2247) <= not((layer0_outputs(897)) or (layer0_outputs(750)));
    layer1_outputs(2248) <= (layer0_outputs(1287)) or (layer0_outputs(1125));
    layer1_outputs(2249) <= not(layer0_outputs(2290));
    layer1_outputs(2250) <= not(layer0_outputs(1297)) or (layer0_outputs(2396));
    layer1_outputs(2251) <= not(layer0_outputs(67)) or (layer0_outputs(2238));
    layer1_outputs(2252) <= '0';
    layer1_outputs(2253) <= (layer0_outputs(1532)) and not (layer0_outputs(1306));
    layer1_outputs(2254) <= not(layer0_outputs(1713)) or (layer0_outputs(689));
    layer1_outputs(2255) <= layer0_outputs(276);
    layer1_outputs(2256) <= (layer0_outputs(2451)) and not (layer0_outputs(2356));
    layer1_outputs(2257) <= (layer0_outputs(1481)) and not (layer0_outputs(2559));
    layer1_outputs(2258) <= not((layer0_outputs(17)) or (layer0_outputs(1192)));
    layer1_outputs(2259) <= '0';
    layer1_outputs(2260) <= layer0_outputs(1815);
    layer1_outputs(2261) <= not((layer0_outputs(577)) xor (layer0_outputs(2362)));
    layer1_outputs(2262) <= not(layer0_outputs(2109));
    layer1_outputs(2263) <= not(layer0_outputs(1876));
    layer1_outputs(2264) <= not(layer0_outputs(524));
    layer1_outputs(2265) <= not(layer0_outputs(1355)) or (layer0_outputs(51));
    layer1_outputs(2266) <= (layer0_outputs(660)) and not (layer0_outputs(1560));
    layer1_outputs(2267) <= not(layer0_outputs(159));
    layer1_outputs(2268) <= '0';
    layer1_outputs(2269) <= layer0_outputs(959);
    layer1_outputs(2270) <= not(layer0_outputs(1443));
    layer1_outputs(2271) <= (layer0_outputs(239)) and not (layer0_outputs(2556));
    layer1_outputs(2272) <= not(layer0_outputs(1981)) or (layer0_outputs(469));
    layer1_outputs(2273) <= not(layer0_outputs(539));
    layer1_outputs(2274) <= (layer0_outputs(887)) or (layer0_outputs(812));
    layer1_outputs(2275) <= not(layer0_outputs(2093)) or (layer0_outputs(1312));
    layer1_outputs(2276) <= '0';
    layer1_outputs(2277) <= not(layer0_outputs(1180));
    layer1_outputs(2278) <= not(layer0_outputs(1400));
    layer1_outputs(2279) <= '1';
    layer1_outputs(2280) <= '0';
    layer1_outputs(2281) <= (layer0_outputs(156)) or (layer0_outputs(1672));
    layer1_outputs(2282) <= '0';
    layer1_outputs(2283) <= layer0_outputs(1603);
    layer1_outputs(2284) <= (layer0_outputs(429)) or (layer0_outputs(213));
    layer1_outputs(2285) <= (layer0_outputs(1530)) and not (layer0_outputs(1729));
    layer1_outputs(2286) <= (layer0_outputs(2292)) or (layer0_outputs(82));
    layer1_outputs(2287) <= (layer0_outputs(533)) and not (layer0_outputs(672));
    layer1_outputs(2288) <= (layer0_outputs(1196)) and (layer0_outputs(2158));
    layer1_outputs(2289) <= not(layer0_outputs(1703));
    layer1_outputs(2290) <= layer0_outputs(980);
    layer1_outputs(2291) <= '1';
    layer1_outputs(2292) <= not(layer0_outputs(228)) or (layer0_outputs(126));
    layer1_outputs(2293) <= not(layer0_outputs(1172)) or (layer0_outputs(310));
    layer1_outputs(2294) <= not((layer0_outputs(317)) and (layer0_outputs(2412)));
    layer1_outputs(2295) <= layer0_outputs(809);
    layer1_outputs(2296) <= not(layer0_outputs(2062));
    layer1_outputs(2297) <= layer0_outputs(1906);
    layer1_outputs(2298) <= '0';
    layer1_outputs(2299) <= (layer0_outputs(1722)) and (layer0_outputs(2439));
    layer1_outputs(2300) <= not(layer0_outputs(1345)) or (layer0_outputs(581));
    layer1_outputs(2301) <= '0';
    layer1_outputs(2302) <= not(layer0_outputs(1120));
    layer1_outputs(2303) <= (layer0_outputs(739)) and (layer0_outputs(1562));
    layer1_outputs(2304) <= (layer0_outputs(1880)) and not (layer0_outputs(1692));
    layer1_outputs(2305) <= not(layer0_outputs(2236));
    layer1_outputs(2306) <= not(layer0_outputs(1));
    layer1_outputs(2307) <= (layer0_outputs(1548)) and not (layer0_outputs(80));
    layer1_outputs(2308) <= layer0_outputs(613);
    layer1_outputs(2309) <= '1';
    layer1_outputs(2310) <= (layer0_outputs(965)) and (layer0_outputs(764));
    layer1_outputs(2311) <= '0';
    layer1_outputs(2312) <= (layer0_outputs(2493)) and (layer0_outputs(1998));
    layer1_outputs(2313) <= '0';
    layer1_outputs(2314) <= layer0_outputs(869);
    layer1_outputs(2315) <= not(layer0_outputs(1230));
    layer1_outputs(2316) <= not(layer0_outputs(353)) or (layer0_outputs(881));
    layer1_outputs(2317) <= not(layer0_outputs(981)) or (layer0_outputs(985));
    layer1_outputs(2318) <= layer0_outputs(1675);
    layer1_outputs(2319) <= layer0_outputs(823);
    layer1_outputs(2320) <= not(layer0_outputs(458)) or (layer0_outputs(854));
    layer1_outputs(2321) <= not((layer0_outputs(1663)) or (layer0_outputs(172)));
    layer1_outputs(2322) <= (layer0_outputs(1359)) and not (layer0_outputs(2289));
    layer1_outputs(2323) <= '1';
    layer1_outputs(2324) <= (layer0_outputs(1021)) and not (layer0_outputs(2209));
    layer1_outputs(2325) <= not((layer0_outputs(1595)) or (layer0_outputs(1121)));
    layer1_outputs(2326) <= (layer0_outputs(2178)) and (layer0_outputs(202));
    layer1_outputs(2327) <= '1';
    layer1_outputs(2328) <= not(layer0_outputs(255));
    layer1_outputs(2329) <= not(layer0_outputs(1045)) or (layer0_outputs(784));
    layer1_outputs(2330) <= '1';
    layer1_outputs(2331) <= layer0_outputs(590);
    layer1_outputs(2332) <= '1';
    layer1_outputs(2333) <= not(layer0_outputs(979));
    layer1_outputs(2334) <= layer0_outputs(302);
    layer1_outputs(2335) <= (layer0_outputs(130)) or (layer0_outputs(1662));
    layer1_outputs(2336) <= '1';
    layer1_outputs(2337) <= not((layer0_outputs(1003)) and (layer0_outputs(2462)));
    layer1_outputs(2338) <= (layer0_outputs(2421)) and (layer0_outputs(813));
    layer1_outputs(2339) <= '0';
    layer1_outputs(2340) <= (layer0_outputs(1718)) and not (layer0_outputs(89));
    layer1_outputs(2341) <= not(layer0_outputs(2315));
    layer1_outputs(2342) <= '0';
    layer1_outputs(2343) <= layer0_outputs(2065);
    layer1_outputs(2344) <= (layer0_outputs(2528)) and not (layer0_outputs(1925));
    layer1_outputs(2345) <= (layer0_outputs(548)) and not (layer0_outputs(2152));
    layer1_outputs(2346) <= (layer0_outputs(838)) and not (layer0_outputs(1176));
    layer1_outputs(2347) <= (layer0_outputs(2313)) and not (layer0_outputs(827));
    layer1_outputs(2348) <= not((layer0_outputs(1244)) and (layer0_outputs(76)));
    layer1_outputs(2349) <= (layer0_outputs(865)) and not (layer0_outputs(2124));
    layer1_outputs(2350) <= (layer0_outputs(788)) or (layer0_outputs(648));
    layer1_outputs(2351) <= layer0_outputs(1069);
    layer1_outputs(2352) <= layer0_outputs(1210);
    layer1_outputs(2353) <= (layer0_outputs(2009)) and not (layer0_outputs(409));
    layer1_outputs(2354) <= not(layer0_outputs(2011)) or (layer0_outputs(2088));
    layer1_outputs(2355) <= not(layer0_outputs(281));
    layer1_outputs(2356) <= '0';
    layer1_outputs(2357) <= not(layer0_outputs(152));
    layer1_outputs(2358) <= layer0_outputs(504);
    layer1_outputs(2359) <= not((layer0_outputs(264)) and (layer0_outputs(1390)));
    layer1_outputs(2360) <= not(layer0_outputs(92));
    layer1_outputs(2361) <= (layer0_outputs(315)) and not (layer0_outputs(1680));
    layer1_outputs(2362) <= '1';
    layer1_outputs(2363) <= not(layer0_outputs(922));
    layer1_outputs(2364) <= not(layer0_outputs(1159));
    layer1_outputs(2365) <= (layer0_outputs(361)) and not (layer0_outputs(718));
    layer1_outputs(2366) <= not(layer0_outputs(754)) or (layer0_outputs(2533));
    layer1_outputs(2367) <= not((layer0_outputs(2532)) and (layer0_outputs(1090)));
    layer1_outputs(2368) <= not(layer0_outputs(286));
    layer1_outputs(2369) <= layer0_outputs(1023);
    layer1_outputs(2370) <= (layer0_outputs(624)) and not (layer0_outputs(1241));
    layer1_outputs(2371) <= '1';
    layer1_outputs(2372) <= layer0_outputs(1772);
    layer1_outputs(2373) <= not((layer0_outputs(956)) and (layer0_outputs(2095)));
    layer1_outputs(2374) <= layer0_outputs(731);
    layer1_outputs(2375) <= not(layer0_outputs(2392)) or (layer0_outputs(271));
    layer1_outputs(2376) <= layer0_outputs(2063);
    layer1_outputs(2377) <= '1';
    layer1_outputs(2378) <= not(layer0_outputs(2535)) or (layer0_outputs(1512));
    layer1_outputs(2379) <= '0';
    layer1_outputs(2380) <= '0';
    layer1_outputs(2381) <= not(layer0_outputs(2393)) or (layer0_outputs(2189));
    layer1_outputs(2382) <= not(layer0_outputs(390));
    layer1_outputs(2383) <= not(layer0_outputs(2410));
    layer1_outputs(2384) <= not(layer0_outputs(2390));
    layer1_outputs(2385) <= not((layer0_outputs(2454)) or (layer0_outputs(1604)));
    layer1_outputs(2386) <= not((layer0_outputs(519)) and (layer0_outputs(285)));
    layer1_outputs(2387) <= not(layer0_outputs(954));
    layer1_outputs(2388) <= not(layer0_outputs(2223));
    layer1_outputs(2389) <= not(layer0_outputs(1924)) or (layer0_outputs(2308));
    layer1_outputs(2390) <= layer0_outputs(1124);
    layer1_outputs(2391) <= (layer0_outputs(345)) and (layer0_outputs(1930));
    layer1_outputs(2392) <= not((layer0_outputs(242)) or (layer0_outputs(675)));
    layer1_outputs(2393) <= not(layer0_outputs(1353));
    layer1_outputs(2394) <= (layer0_outputs(1480)) and not (layer0_outputs(1357));
    layer1_outputs(2395) <= '0';
    layer1_outputs(2396) <= not(layer0_outputs(1247)) or (layer0_outputs(1034));
    layer1_outputs(2397) <= (layer0_outputs(2358)) and not (layer0_outputs(1123));
    layer1_outputs(2398) <= not(layer0_outputs(198));
    layer1_outputs(2399) <= '0';
    layer1_outputs(2400) <= not(layer0_outputs(2502)) or (layer0_outputs(1385));
    layer1_outputs(2401) <= '1';
    layer1_outputs(2402) <= '1';
    layer1_outputs(2403) <= '0';
    layer1_outputs(2404) <= (layer0_outputs(1427)) and (layer0_outputs(764));
    layer1_outputs(2405) <= '1';
    layer1_outputs(2406) <= layer0_outputs(1263);
    layer1_outputs(2407) <= layer0_outputs(1420);
    layer1_outputs(2408) <= not(layer0_outputs(2373)) or (layer0_outputs(1287));
    layer1_outputs(2409) <= (layer0_outputs(2327)) or (layer0_outputs(2507));
    layer1_outputs(2410) <= (layer0_outputs(2550)) and not (layer0_outputs(2387));
    layer1_outputs(2411) <= not((layer0_outputs(455)) or (layer0_outputs(1407)));
    layer1_outputs(2412) <= not(layer0_outputs(2159));
    layer1_outputs(2413) <= not((layer0_outputs(2446)) or (layer0_outputs(1525)));
    layer1_outputs(2414) <= not(layer0_outputs(958));
    layer1_outputs(2415) <= (layer0_outputs(143)) and not (layer0_outputs(535));
    layer1_outputs(2416) <= not(layer0_outputs(1258)) or (layer0_outputs(2046));
    layer1_outputs(2417) <= not((layer0_outputs(1222)) xor (layer0_outputs(704)));
    layer1_outputs(2418) <= (layer0_outputs(1829)) or (layer0_outputs(1223));
    layer1_outputs(2419) <= not(layer0_outputs(2426)) or (layer0_outputs(971));
    layer1_outputs(2420) <= (layer0_outputs(504)) and (layer0_outputs(1854));
    layer1_outputs(2421) <= layer0_outputs(969);
    layer1_outputs(2422) <= layer0_outputs(510);
    layer1_outputs(2423) <= (layer0_outputs(1518)) or (layer0_outputs(1562));
    layer1_outputs(2424) <= not(layer0_outputs(2039));
    layer1_outputs(2425) <= '0';
    layer1_outputs(2426) <= not(layer0_outputs(2126)) or (layer0_outputs(2211));
    layer1_outputs(2427) <= not(layer0_outputs(1087));
    layer1_outputs(2428) <= not((layer0_outputs(910)) or (layer0_outputs(78)));
    layer1_outputs(2429) <= layer0_outputs(2023);
    layer1_outputs(2430) <= not((layer0_outputs(2161)) or (layer0_outputs(799)));
    layer1_outputs(2431) <= not((layer0_outputs(1661)) and (layer0_outputs(229)));
    layer1_outputs(2432) <= not((layer0_outputs(139)) and (layer0_outputs(1705)));
    layer1_outputs(2433) <= (layer0_outputs(379)) and not (layer0_outputs(1990));
    layer1_outputs(2434) <= layer0_outputs(1662);
    layer1_outputs(2435) <= (layer0_outputs(1630)) and (layer0_outputs(893));
    layer1_outputs(2436) <= (layer0_outputs(721)) and (layer0_outputs(2417));
    layer1_outputs(2437) <= layer0_outputs(230);
    layer1_outputs(2438) <= '1';
    layer1_outputs(2439) <= '0';
    layer1_outputs(2440) <= layer0_outputs(1089);
    layer1_outputs(2441) <= (layer0_outputs(1657)) and (layer0_outputs(356));
    layer1_outputs(2442) <= (layer0_outputs(292)) xor (layer0_outputs(846));
    layer1_outputs(2443) <= (layer0_outputs(785)) or (layer0_outputs(1773));
    layer1_outputs(2444) <= (layer0_outputs(1579)) and (layer0_outputs(43));
    layer1_outputs(2445) <= '0';
    layer1_outputs(2446) <= (layer0_outputs(1812)) and (layer0_outputs(716));
    layer1_outputs(2447) <= (layer0_outputs(1899)) and (layer0_outputs(1717));
    layer1_outputs(2448) <= (layer0_outputs(846)) and (layer0_outputs(1004));
    layer1_outputs(2449) <= (layer0_outputs(2170)) and not (layer0_outputs(585));
    layer1_outputs(2450) <= '0';
    layer1_outputs(2451) <= layer0_outputs(532);
    layer1_outputs(2452) <= (layer0_outputs(727)) and (layer0_outputs(450));
    layer1_outputs(2453) <= not((layer0_outputs(814)) or (layer0_outputs(1283)));
    layer1_outputs(2454) <= layer0_outputs(1459);
    layer1_outputs(2455) <= not((layer0_outputs(583)) or (layer0_outputs(656)));
    layer1_outputs(2456) <= '1';
    layer1_outputs(2457) <= '1';
    layer1_outputs(2458) <= layer0_outputs(1231);
    layer1_outputs(2459) <= not((layer0_outputs(1405)) or (layer0_outputs(2)));
    layer1_outputs(2460) <= (layer0_outputs(1321)) and not (layer0_outputs(756));
    layer1_outputs(2461) <= '0';
    layer1_outputs(2462) <= (layer0_outputs(42)) and (layer0_outputs(1447));
    layer1_outputs(2463) <= layer0_outputs(1904);
    layer1_outputs(2464) <= layer0_outputs(771);
    layer1_outputs(2465) <= '0';
    layer1_outputs(2466) <= not((layer0_outputs(1391)) or (layer0_outputs(1009)));
    layer1_outputs(2467) <= not(layer0_outputs(9)) or (layer0_outputs(189));
    layer1_outputs(2468) <= (layer0_outputs(2297)) and not (layer0_outputs(804));
    layer1_outputs(2469) <= (layer0_outputs(25)) xor (layer0_outputs(1179));
    layer1_outputs(2470) <= layer0_outputs(1902);
    layer1_outputs(2471) <= not(layer0_outputs(1065));
    layer1_outputs(2472) <= not(layer0_outputs(881));
    layer1_outputs(2473) <= (layer0_outputs(2352)) and not (layer0_outputs(2253));
    layer1_outputs(2474) <= (layer0_outputs(2385)) and not (layer0_outputs(69));
    layer1_outputs(2475) <= (layer0_outputs(547)) or (layer0_outputs(723));
    layer1_outputs(2476) <= not(layer0_outputs(1279));
    layer1_outputs(2477) <= (layer0_outputs(1835)) or (layer0_outputs(1384));
    layer1_outputs(2478) <= layer0_outputs(958);
    layer1_outputs(2479) <= not(layer0_outputs(1214)) or (layer0_outputs(2071));
    layer1_outputs(2480) <= not(layer0_outputs(1765));
    layer1_outputs(2481) <= not((layer0_outputs(205)) or (layer0_outputs(122)));
    layer1_outputs(2482) <= not(layer0_outputs(1449)) or (layer0_outputs(1166));
    layer1_outputs(2483) <= not((layer0_outputs(2041)) and (layer0_outputs(70)));
    layer1_outputs(2484) <= (layer0_outputs(1969)) and (layer0_outputs(1592));
    layer1_outputs(2485) <= not(layer0_outputs(677));
    layer1_outputs(2486) <= (layer0_outputs(1155)) and not (layer0_outputs(1422));
    layer1_outputs(2487) <= not((layer0_outputs(1595)) or (layer0_outputs(1665)));
    layer1_outputs(2488) <= layer0_outputs(19);
    layer1_outputs(2489) <= not(layer0_outputs(2434));
    layer1_outputs(2490) <= (layer0_outputs(1851)) and (layer0_outputs(2215));
    layer1_outputs(2491) <= not((layer0_outputs(974)) and (layer0_outputs(87)));
    layer1_outputs(2492) <= not(layer0_outputs(620)) or (layer0_outputs(2321));
    layer1_outputs(2493) <= '1';
    layer1_outputs(2494) <= layer0_outputs(218);
    layer1_outputs(2495) <= layer0_outputs(2235);
    layer1_outputs(2496) <= not(layer0_outputs(1549)) or (layer0_outputs(1025));
    layer1_outputs(2497) <= '1';
    layer1_outputs(2498) <= not(layer0_outputs(2122)) or (layer0_outputs(1210));
    layer1_outputs(2499) <= layer0_outputs(1147);
    layer1_outputs(2500) <= '1';
    layer1_outputs(2501) <= (layer0_outputs(1162)) and not (layer0_outputs(2043));
    layer1_outputs(2502) <= (layer0_outputs(2083)) and not (layer0_outputs(330));
    layer1_outputs(2503) <= '0';
    layer1_outputs(2504) <= not(layer0_outputs(479));
    layer1_outputs(2505) <= not((layer0_outputs(403)) and (layer0_outputs(443)));
    layer1_outputs(2506) <= '0';
    layer1_outputs(2507) <= not((layer0_outputs(853)) and (layer0_outputs(648)));
    layer1_outputs(2508) <= (layer0_outputs(908)) and (layer0_outputs(502));
    layer1_outputs(2509) <= layer0_outputs(189);
    layer1_outputs(2510) <= '1';
    layer1_outputs(2511) <= not(layer0_outputs(2316));
    layer1_outputs(2512) <= (layer0_outputs(741)) and not (layer0_outputs(729));
    layer1_outputs(2513) <= '0';
    layer1_outputs(2514) <= (layer0_outputs(830)) and not (layer0_outputs(1701));
    layer1_outputs(2515) <= '1';
    layer1_outputs(2516) <= not(layer0_outputs(2415));
    layer1_outputs(2517) <= '0';
    layer1_outputs(2518) <= not((layer0_outputs(2383)) and (layer0_outputs(821)));
    layer1_outputs(2519) <= '0';
    layer1_outputs(2520) <= not((layer0_outputs(164)) or (layer0_outputs(191)));
    layer1_outputs(2521) <= not(layer0_outputs(481)) or (layer0_outputs(976));
    layer1_outputs(2522) <= '1';
    layer1_outputs(2523) <= not(layer0_outputs(2156)) or (layer0_outputs(2092));
    layer1_outputs(2524) <= not((layer0_outputs(1642)) and (layer0_outputs(885)));
    layer1_outputs(2525) <= not(layer0_outputs(1586));
    layer1_outputs(2526) <= not(layer0_outputs(2524)) or (layer0_outputs(1843));
    layer1_outputs(2527) <= not((layer0_outputs(820)) or (layer0_outputs(1493)));
    layer1_outputs(2528) <= '0';
    layer1_outputs(2529) <= not(layer0_outputs(2391));
    layer1_outputs(2530) <= (layer0_outputs(2029)) xor (layer0_outputs(1299));
    layer1_outputs(2531) <= not(layer0_outputs(903));
    layer1_outputs(2532) <= layer0_outputs(2078);
    layer1_outputs(2533) <= not(layer0_outputs(1264)) or (layer0_outputs(2160));
    layer1_outputs(2534) <= not(layer0_outputs(950));
    layer1_outputs(2535) <= (layer0_outputs(1703)) and not (layer0_outputs(354));
    layer1_outputs(2536) <= (layer0_outputs(2456)) and not (layer0_outputs(1621));
    layer1_outputs(2537) <= not((layer0_outputs(2228)) or (layer0_outputs(1372)));
    layer1_outputs(2538) <= not(layer0_outputs(1265));
    layer1_outputs(2539) <= '1';
    layer1_outputs(2540) <= (layer0_outputs(1218)) and (layer0_outputs(2233));
    layer1_outputs(2541) <= not((layer0_outputs(88)) or (layer0_outputs(105)));
    layer1_outputs(2542) <= not(layer0_outputs(1993)) or (layer0_outputs(2049));
    layer1_outputs(2543) <= not(layer0_outputs(1980));
    layer1_outputs(2544) <= not(layer0_outputs(2151)) or (layer0_outputs(1905));
    layer1_outputs(2545) <= not(layer0_outputs(800));
    layer1_outputs(2546) <= not((layer0_outputs(1430)) or (layer0_outputs(1794)));
    layer1_outputs(2547) <= not(layer0_outputs(1352));
    layer1_outputs(2548) <= layer0_outputs(1181);
    layer1_outputs(2549) <= (layer0_outputs(1421)) and not (layer0_outputs(909));
    layer1_outputs(2550) <= '1';
    layer1_outputs(2551) <= not(layer0_outputs(1593)) or (layer0_outputs(2542));
    layer1_outputs(2552) <= (layer0_outputs(1584)) and (layer0_outputs(358));
    layer1_outputs(2553) <= (layer0_outputs(2470)) and (layer0_outputs(1403));
    layer1_outputs(2554) <= layer0_outputs(1515);
    layer1_outputs(2555) <= '0';
    layer1_outputs(2556) <= (layer0_outputs(1204)) or (layer0_outputs(824));
    layer1_outputs(2557) <= not(layer0_outputs(1419)) or (layer0_outputs(915));
    layer1_outputs(2558) <= '0';
    layer1_outputs(2559) <= not(layer0_outputs(1587)) or (layer0_outputs(2201));
    layer2_outputs(0) <= not((layer1_outputs(105)) or (layer1_outputs(1458)));
    layer2_outputs(1) <= not(layer1_outputs(1019)) or (layer1_outputs(1424));
    layer2_outputs(2) <= (layer1_outputs(1793)) or (layer1_outputs(315));
    layer2_outputs(3) <= (layer1_outputs(603)) or (layer1_outputs(1010));
    layer2_outputs(4) <= (layer1_outputs(2076)) and (layer1_outputs(1876));
    layer2_outputs(5) <= not(layer1_outputs(664));
    layer2_outputs(6) <= not(layer1_outputs(1423)) or (layer1_outputs(1921));
    layer2_outputs(7) <= (layer1_outputs(2519)) and not (layer1_outputs(913));
    layer2_outputs(8) <= '0';
    layer2_outputs(9) <= not(layer1_outputs(1591));
    layer2_outputs(10) <= (layer1_outputs(666)) or (layer1_outputs(1055));
    layer2_outputs(11) <= (layer1_outputs(1394)) and (layer1_outputs(586));
    layer2_outputs(12) <= not((layer1_outputs(526)) and (layer1_outputs(2199)));
    layer2_outputs(13) <= (layer1_outputs(1980)) and not (layer1_outputs(2328));
    layer2_outputs(14) <= not((layer1_outputs(1512)) or (layer1_outputs(725)));
    layer2_outputs(15) <= '0';
    layer2_outputs(16) <= not(layer1_outputs(949));
    layer2_outputs(17) <= (layer1_outputs(2236)) and not (layer1_outputs(1409));
    layer2_outputs(18) <= not((layer1_outputs(596)) and (layer1_outputs(1288)));
    layer2_outputs(19) <= not(layer1_outputs(2536));
    layer2_outputs(20) <= (layer1_outputs(2427)) and not (layer1_outputs(2091));
    layer2_outputs(21) <= not((layer1_outputs(2533)) or (layer1_outputs(2378)));
    layer2_outputs(22) <= (layer1_outputs(372)) and not (layer1_outputs(125));
    layer2_outputs(23) <= not(layer1_outputs(822)) or (layer1_outputs(1588));
    layer2_outputs(24) <= (layer1_outputs(202)) and (layer1_outputs(1354));
    layer2_outputs(25) <= layer1_outputs(2431);
    layer2_outputs(26) <= layer1_outputs(1155);
    layer2_outputs(27) <= not(layer1_outputs(803));
    layer2_outputs(28) <= layer1_outputs(848);
    layer2_outputs(29) <= '1';
    layer2_outputs(30) <= not((layer1_outputs(26)) and (layer1_outputs(2251)));
    layer2_outputs(31) <= not(layer1_outputs(1556));
    layer2_outputs(32) <= not((layer1_outputs(1723)) xor (layer1_outputs(1046)));
    layer2_outputs(33) <= (layer1_outputs(717)) or (layer1_outputs(1763));
    layer2_outputs(34) <= not(layer1_outputs(1340));
    layer2_outputs(35) <= '1';
    layer2_outputs(36) <= not(layer1_outputs(897)) or (layer1_outputs(1655));
    layer2_outputs(37) <= not((layer1_outputs(2257)) and (layer1_outputs(2365)));
    layer2_outputs(38) <= (layer1_outputs(2116)) and not (layer1_outputs(1520));
    layer2_outputs(39) <= not(layer1_outputs(969));
    layer2_outputs(40) <= (layer1_outputs(1921)) and not (layer1_outputs(1443));
    layer2_outputs(41) <= layer1_outputs(1260);
    layer2_outputs(42) <= not((layer1_outputs(1836)) and (layer1_outputs(1183)));
    layer2_outputs(43) <= layer1_outputs(1100);
    layer2_outputs(44) <= layer1_outputs(1424);
    layer2_outputs(45) <= '0';
    layer2_outputs(46) <= not(layer1_outputs(2405)) or (layer1_outputs(948));
    layer2_outputs(47) <= not(layer1_outputs(1143));
    layer2_outputs(48) <= not(layer1_outputs(935)) or (layer1_outputs(1985));
    layer2_outputs(49) <= not(layer1_outputs(383)) or (layer1_outputs(1300));
    layer2_outputs(50) <= layer1_outputs(627);
    layer2_outputs(51) <= not((layer1_outputs(1071)) and (layer1_outputs(1126)));
    layer2_outputs(52) <= not((layer1_outputs(1410)) or (layer1_outputs(1472)));
    layer2_outputs(53) <= (layer1_outputs(1670)) and not (layer1_outputs(542));
    layer2_outputs(54) <= not(layer1_outputs(401)) or (layer1_outputs(1850));
    layer2_outputs(55) <= not(layer1_outputs(2038));
    layer2_outputs(56) <= not(layer1_outputs(341));
    layer2_outputs(57) <= '0';
    layer2_outputs(58) <= layer1_outputs(598);
    layer2_outputs(59) <= not(layer1_outputs(2171));
    layer2_outputs(60) <= (layer1_outputs(365)) and not (layer1_outputs(2168));
    layer2_outputs(61) <= '1';
    layer2_outputs(62) <= not((layer1_outputs(2368)) and (layer1_outputs(388)));
    layer2_outputs(63) <= (layer1_outputs(586)) and not (layer1_outputs(2334));
    layer2_outputs(64) <= layer1_outputs(1687);
    layer2_outputs(65) <= layer1_outputs(2159);
    layer2_outputs(66) <= not((layer1_outputs(1813)) or (layer1_outputs(530)));
    layer2_outputs(67) <= not(layer1_outputs(1707)) or (layer1_outputs(1393));
    layer2_outputs(68) <= layer1_outputs(1012);
    layer2_outputs(69) <= (layer1_outputs(971)) and not (layer1_outputs(259));
    layer2_outputs(70) <= (layer1_outputs(103)) and not (layer1_outputs(925));
    layer2_outputs(71) <= '0';
    layer2_outputs(72) <= '1';
    layer2_outputs(73) <= '0';
    layer2_outputs(74) <= not((layer1_outputs(233)) and (layer1_outputs(2483)));
    layer2_outputs(75) <= layer1_outputs(61);
    layer2_outputs(76) <= not(layer1_outputs(215));
    layer2_outputs(77) <= not((layer1_outputs(2047)) and (layer1_outputs(545)));
    layer2_outputs(78) <= layer1_outputs(2537);
    layer2_outputs(79) <= layer1_outputs(1310);
    layer2_outputs(80) <= not(layer1_outputs(1268)) or (layer1_outputs(845));
    layer2_outputs(81) <= not(layer1_outputs(1373));
    layer2_outputs(82) <= not(layer1_outputs(520)) or (layer1_outputs(139));
    layer2_outputs(83) <= not(layer1_outputs(2197)) or (layer1_outputs(1830));
    layer2_outputs(84) <= not(layer1_outputs(132)) or (layer1_outputs(2492));
    layer2_outputs(85) <= layer1_outputs(1270);
    layer2_outputs(86) <= '1';
    layer2_outputs(87) <= '0';
    layer2_outputs(88) <= not(layer1_outputs(1553));
    layer2_outputs(89) <= layer1_outputs(963);
    layer2_outputs(90) <= (layer1_outputs(932)) and not (layer1_outputs(1185));
    layer2_outputs(91) <= not(layer1_outputs(1105));
    layer2_outputs(92) <= not(layer1_outputs(1257)) or (layer1_outputs(469));
    layer2_outputs(93) <= not((layer1_outputs(149)) or (layer1_outputs(1018)));
    layer2_outputs(94) <= '1';
    layer2_outputs(95) <= not((layer1_outputs(608)) and (layer1_outputs(1795)));
    layer2_outputs(96) <= '1';
    layer2_outputs(97) <= (layer1_outputs(932)) and (layer1_outputs(411));
    layer2_outputs(98) <= not(layer1_outputs(647));
    layer2_outputs(99) <= not(layer1_outputs(2157));
    layer2_outputs(100) <= not(layer1_outputs(2057));
    layer2_outputs(101) <= not((layer1_outputs(601)) xor (layer1_outputs(2113)));
    layer2_outputs(102) <= '1';
    layer2_outputs(103) <= not(layer1_outputs(640));
    layer2_outputs(104) <= not(layer1_outputs(657));
    layer2_outputs(105) <= '0';
    layer2_outputs(106) <= not((layer1_outputs(1489)) or (layer1_outputs(752)));
    layer2_outputs(107) <= not(layer1_outputs(54));
    layer2_outputs(108) <= '0';
    layer2_outputs(109) <= (layer1_outputs(344)) and not (layer1_outputs(1911));
    layer2_outputs(110) <= not((layer1_outputs(570)) or (layer1_outputs(763)));
    layer2_outputs(111) <= layer1_outputs(1434);
    layer2_outputs(112) <= '0';
    layer2_outputs(113) <= not(layer1_outputs(792));
    layer2_outputs(114) <= layer1_outputs(2297);
    layer2_outputs(115) <= not(layer1_outputs(675));
    layer2_outputs(116) <= '0';
    layer2_outputs(117) <= (layer1_outputs(1301)) and not (layer1_outputs(1187));
    layer2_outputs(118) <= not(layer1_outputs(205)) or (layer1_outputs(907));
    layer2_outputs(119) <= layer1_outputs(267);
    layer2_outputs(120) <= (layer1_outputs(1565)) or (layer1_outputs(2526));
    layer2_outputs(121) <= not((layer1_outputs(1630)) or (layer1_outputs(392)));
    layer2_outputs(122) <= not((layer1_outputs(236)) or (layer1_outputs(1054)));
    layer2_outputs(123) <= '0';
    layer2_outputs(124) <= (layer1_outputs(1876)) or (layer1_outputs(2244));
    layer2_outputs(125) <= (layer1_outputs(955)) and not (layer1_outputs(1388));
    layer2_outputs(126) <= (layer1_outputs(13)) and not (layer1_outputs(1532));
    layer2_outputs(127) <= layer1_outputs(673);
    layer2_outputs(128) <= not((layer1_outputs(12)) or (layer1_outputs(415)));
    layer2_outputs(129) <= not(layer1_outputs(1976));
    layer2_outputs(130) <= not(layer1_outputs(311));
    layer2_outputs(131) <= '0';
    layer2_outputs(132) <= (layer1_outputs(811)) and not (layer1_outputs(1122));
    layer2_outputs(133) <= (layer1_outputs(1216)) and (layer1_outputs(817));
    layer2_outputs(134) <= (layer1_outputs(191)) or (layer1_outputs(165));
    layer2_outputs(135) <= '1';
    layer2_outputs(136) <= '0';
    layer2_outputs(137) <= '0';
    layer2_outputs(138) <= not(layer1_outputs(394));
    layer2_outputs(139) <= '0';
    layer2_outputs(140) <= (layer1_outputs(2438)) or (layer1_outputs(2143));
    layer2_outputs(141) <= not(layer1_outputs(2388));
    layer2_outputs(142) <= not(layer1_outputs(157)) or (layer1_outputs(2146));
    layer2_outputs(143) <= not(layer1_outputs(1468)) or (layer1_outputs(1182));
    layer2_outputs(144) <= not((layer1_outputs(1117)) or (layer1_outputs(1656)));
    layer2_outputs(145) <= layer1_outputs(390);
    layer2_outputs(146) <= (layer1_outputs(911)) and (layer1_outputs(1823));
    layer2_outputs(147) <= '1';
    layer2_outputs(148) <= (layer1_outputs(1351)) and not (layer1_outputs(1373));
    layer2_outputs(149) <= not((layer1_outputs(787)) xor (layer1_outputs(854)));
    layer2_outputs(150) <= (layer1_outputs(533)) or (layer1_outputs(240));
    layer2_outputs(151) <= layer1_outputs(799);
    layer2_outputs(152) <= not(layer1_outputs(1081)) or (layer1_outputs(1181));
    layer2_outputs(153) <= not((layer1_outputs(195)) or (layer1_outputs(611)));
    layer2_outputs(154) <= not(layer1_outputs(2398));
    layer2_outputs(155) <= not(layer1_outputs(2485));
    layer2_outputs(156) <= layer1_outputs(1583);
    layer2_outputs(157) <= '1';
    layer2_outputs(158) <= '0';
    layer2_outputs(159) <= not((layer1_outputs(987)) or (layer1_outputs(733)));
    layer2_outputs(160) <= not(layer1_outputs(933)) or (layer1_outputs(1122));
    layer2_outputs(161) <= not(layer1_outputs(1954));
    layer2_outputs(162) <= (layer1_outputs(1453)) xor (layer1_outputs(2101));
    layer2_outputs(163) <= layer1_outputs(1628);
    layer2_outputs(164) <= not(layer1_outputs(2095)) or (layer1_outputs(1367));
    layer2_outputs(165) <= (layer1_outputs(581)) or (layer1_outputs(2223));
    layer2_outputs(166) <= not(layer1_outputs(1294));
    layer2_outputs(167) <= not(layer1_outputs(1360));
    layer2_outputs(168) <= '1';
    layer2_outputs(169) <= not(layer1_outputs(1996));
    layer2_outputs(170) <= not(layer1_outputs(1030)) or (layer1_outputs(1534));
    layer2_outputs(171) <= not((layer1_outputs(1566)) or (layer1_outputs(226)));
    layer2_outputs(172) <= layer1_outputs(825);
    layer2_outputs(173) <= '0';
    layer2_outputs(174) <= not(layer1_outputs(1885)) or (layer1_outputs(1875));
    layer2_outputs(175) <= not((layer1_outputs(254)) and (layer1_outputs(2243)));
    layer2_outputs(176) <= not(layer1_outputs(57)) or (layer1_outputs(1230));
    layer2_outputs(177) <= (layer1_outputs(1004)) or (layer1_outputs(464));
    layer2_outputs(178) <= layer1_outputs(1860);
    layer2_outputs(179) <= (layer1_outputs(239)) and not (layer1_outputs(448));
    layer2_outputs(180) <= '0';
    layer2_outputs(181) <= (layer1_outputs(639)) or (layer1_outputs(975));
    layer2_outputs(182) <= (layer1_outputs(831)) and not (layer1_outputs(2149));
    layer2_outputs(183) <= not(layer1_outputs(714)) or (layer1_outputs(1857));
    layer2_outputs(184) <= not(layer1_outputs(2307)) or (layer1_outputs(2078));
    layer2_outputs(185) <= not(layer1_outputs(601)) or (layer1_outputs(160));
    layer2_outputs(186) <= '1';
    layer2_outputs(187) <= layer1_outputs(1780);
    layer2_outputs(188) <= '1';
    layer2_outputs(189) <= '1';
    layer2_outputs(190) <= not((layer1_outputs(1113)) and (layer1_outputs(1103)));
    layer2_outputs(191) <= not(layer1_outputs(2252)) or (layer1_outputs(2337));
    layer2_outputs(192) <= (layer1_outputs(645)) and not (layer1_outputs(2353));
    layer2_outputs(193) <= layer1_outputs(1800);
    layer2_outputs(194) <= not(layer1_outputs(995));
    layer2_outputs(195) <= not(layer1_outputs(912));
    layer2_outputs(196) <= layer1_outputs(840);
    layer2_outputs(197) <= not((layer1_outputs(1696)) or (layer1_outputs(1746)));
    layer2_outputs(198) <= (layer1_outputs(600)) and not (layer1_outputs(1431));
    layer2_outputs(199) <= '0';
    layer2_outputs(200) <= layer1_outputs(1644);
    layer2_outputs(201) <= layer1_outputs(167);
    layer2_outputs(202) <= layer1_outputs(379);
    layer2_outputs(203) <= not(layer1_outputs(1653));
    layer2_outputs(204) <= (layer1_outputs(1961)) and not (layer1_outputs(2516));
    layer2_outputs(205) <= not(layer1_outputs(653));
    layer2_outputs(206) <= (layer1_outputs(2067)) and (layer1_outputs(755));
    layer2_outputs(207) <= '1';
    layer2_outputs(208) <= not(layer1_outputs(470));
    layer2_outputs(209) <= not((layer1_outputs(2204)) and (layer1_outputs(810)));
    layer2_outputs(210) <= (layer1_outputs(2198)) or (layer1_outputs(315));
    layer2_outputs(211) <= layer1_outputs(2308);
    layer2_outputs(212) <= (layer1_outputs(250)) or (layer1_outputs(1142));
    layer2_outputs(213) <= not(layer1_outputs(1866)) or (layer1_outputs(203));
    layer2_outputs(214) <= not((layer1_outputs(701)) xor (layer1_outputs(1097)));
    layer2_outputs(215) <= (layer1_outputs(1322)) and not (layer1_outputs(2324));
    layer2_outputs(216) <= layer1_outputs(386);
    layer2_outputs(217) <= '0';
    layer2_outputs(218) <= layer1_outputs(2007);
    layer2_outputs(219) <= (layer1_outputs(435)) and not (layer1_outputs(2441));
    layer2_outputs(220) <= layer1_outputs(1676);
    layer2_outputs(221) <= not(layer1_outputs(2481));
    layer2_outputs(222) <= (layer1_outputs(2262)) and not (layer1_outputs(291));
    layer2_outputs(223) <= not(layer1_outputs(164)) or (layer1_outputs(2479));
    layer2_outputs(224) <= not((layer1_outputs(1411)) or (layer1_outputs(1338)));
    layer2_outputs(225) <= not((layer1_outputs(189)) or (layer1_outputs(371)));
    layer2_outputs(226) <= (layer1_outputs(2121)) and not (layer1_outputs(622));
    layer2_outputs(227) <= (layer1_outputs(656)) and not (layer1_outputs(2483));
    layer2_outputs(228) <= not(layer1_outputs(201));
    layer2_outputs(229) <= layer1_outputs(1833);
    layer2_outputs(230) <= not(layer1_outputs(1990)) or (layer1_outputs(578));
    layer2_outputs(231) <= layer1_outputs(2006);
    layer2_outputs(232) <= (layer1_outputs(2391)) or (layer1_outputs(1093));
    layer2_outputs(233) <= not(layer1_outputs(1200));
    layer2_outputs(234) <= (layer1_outputs(830)) and not (layer1_outputs(346));
    layer2_outputs(235) <= (layer1_outputs(465)) and (layer1_outputs(1852));
    layer2_outputs(236) <= not(layer1_outputs(2107));
    layer2_outputs(237) <= layer1_outputs(393);
    layer2_outputs(238) <= not(layer1_outputs(2488));
    layer2_outputs(239) <= not((layer1_outputs(1821)) or (layer1_outputs(1975)));
    layer2_outputs(240) <= (layer1_outputs(616)) and not (layer1_outputs(2382));
    layer2_outputs(241) <= not(layer1_outputs(667)) or (layer1_outputs(2115));
    layer2_outputs(242) <= not(layer1_outputs(1191));
    layer2_outputs(243) <= (layer1_outputs(881)) and (layer1_outputs(1337));
    layer2_outputs(244) <= layer1_outputs(787);
    layer2_outputs(245) <= (layer1_outputs(475)) and (layer1_outputs(820));
    layer2_outputs(246) <= (layer1_outputs(362)) and (layer1_outputs(837));
    layer2_outputs(247) <= '1';
    layer2_outputs(248) <= not(layer1_outputs(2413)) or (layer1_outputs(1699));
    layer2_outputs(249) <= not(layer1_outputs(1339)) or (layer1_outputs(985));
    layer2_outputs(250) <= layer1_outputs(2134);
    layer2_outputs(251) <= not(layer1_outputs(1125));
    layer2_outputs(252) <= not((layer1_outputs(1759)) or (layer1_outputs(2145)));
    layer2_outputs(253) <= (layer1_outputs(507)) and not (layer1_outputs(2424));
    layer2_outputs(254) <= '0';
    layer2_outputs(255) <= not(layer1_outputs(512));
    layer2_outputs(256) <= '1';
    layer2_outputs(257) <= not(layer1_outputs(485));
    layer2_outputs(258) <= (layer1_outputs(112)) and (layer1_outputs(2523));
    layer2_outputs(259) <= '0';
    layer2_outputs(260) <= '1';
    layer2_outputs(261) <= '0';
    layer2_outputs(262) <= (layer1_outputs(1037)) and (layer1_outputs(1516));
    layer2_outputs(263) <= layer1_outputs(2297);
    layer2_outputs(264) <= '1';
    layer2_outputs(265) <= '0';
    layer2_outputs(266) <= not(layer1_outputs(2251));
    layer2_outputs(267) <= not(layer1_outputs(2123));
    layer2_outputs(268) <= not(layer1_outputs(192)) or (layer1_outputs(681));
    layer2_outputs(269) <= (layer1_outputs(2419)) and not (layer1_outputs(2534));
    layer2_outputs(270) <= (layer1_outputs(1065)) and not (layer1_outputs(2543));
    layer2_outputs(271) <= (layer1_outputs(2007)) and (layer1_outputs(2434));
    layer2_outputs(272) <= layer1_outputs(2001);
    layer2_outputs(273) <= '0';
    layer2_outputs(274) <= layer1_outputs(2242);
    layer2_outputs(275) <= '0';
    layer2_outputs(276) <= layer1_outputs(2135);
    layer2_outputs(277) <= '0';
    layer2_outputs(278) <= (layer1_outputs(2232)) and not (layer1_outputs(2177));
    layer2_outputs(279) <= '1';
    layer2_outputs(280) <= '1';
    layer2_outputs(281) <= not(layer1_outputs(773));
    layer2_outputs(282) <= (layer1_outputs(1671)) and not (layer1_outputs(1697));
    layer2_outputs(283) <= (layer1_outputs(2346)) and not (layer1_outputs(1968));
    layer2_outputs(284) <= layer1_outputs(2056);
    layer2_outputs(285) <= not(layer1_outputs(1959)) or (layer1_outputs(2497));
    layer2_outputs(286) <= (layer1_outputs(227)) and not (layer1_outputs(2551));
    layer2_outputs(287) <= (layer1_outputs(981)) and (layer1_outputs(815));
    layer2_outputs(288) <= '1';
    layer2_outputs(289) <= not(layer1_outputs(2372));
    layer2_outputs(290) <= '1';
    layer2_outputs(291) <= (layer1_outputs(2239)) and not (layer1_outputs(901));
    layer2_outputs(292) <= (layer1_outputs(527)) xor (layer1_outputs(209));
    layer2_outputs(293) <= '1';
    layer2_outputs(294) <= (layer1_outputs(953)) and (layer1_outputs(1933));
    layer2_outputs(295) <= '0';
    layer2_outputs(296) <= not(layer1_outputs(1112)) or (layer1_outputs(186));
    layer2_outputs(297) <= not(layer1_outputs(2394));
    layer2_outputs(298) <= (layer1_outputs(552)) xor (layer1_outputs(308));
    layer2_outputs(299) <= (layer1_outputs(1212)) and (layer1_outputs(337));
    layer2_outputs(300) <= not(layer1_outputs(73));
    layer2_outputs(301) <= (layer1_outputs(34)) and not (layer1_outputs(1204));
    layer2_outputs(302) <= '1';
    layer2_outputs(303) <= not(layer1_outputs(2213));
    layer2_outputs(304) <= (layer1_outputs(1372)) and (layer1_outputs(2226));
    layer2_outputs(305) <= not(layer1_outputs(475));
    layer2_outputs(306) <= not(layer1_outputs(1332));
    layer2_outputs(307) <= not(layer1_outputs(300)) or (layer1_outputs(2015));
    layer2_outputs(308) <= '1';
    layer2_outputs(309) <= not((layer1_outputs(1089)) xor (layer1_outputs(6)));
    layer2_outputs(310) <= layer1_outputs(318);
    layer2_outputs(311) <= not(layer1_outputs(1718));
    layer2_outputs(312) <= (layer1_outputs(1283)) and (layer1_outputs(418));
    layer2_outputs(313) <= (layer1_outputs(2042)) or (layer1_outputs(419));
    layer2_outputs(314) <= not(layer1_outputs(1058)) or (layer1_outputs(1259));
    layer2_outputs(315) <= layer1_outputs(1457);
    layer2_outputs(316) <= not(layer1_outputs(2010)) or (layer1_outputs(340));
    layer2_outputs(317) <= (layer1_outputs(1250)) or (layer1_outputs(1794));
    layer2_outputs(318) <= '1';
    layer2_outputs(319) <= '0';
    layer2_outputs(320) <= not(layer1_outputs(1712)) or (layer1_outputs(855));
    layer2_outputs(321) <= (layer1_outputs(2402)) or (layer1_outputs(1435));
    layer2_outputs(322) <= (layer1_outputs(1081)) and not (layer1_outputs(509));
    layer2_outputs(323) <= layer1_outputs(209);
    layer2_outputs(324) <= not((layer1_outputs(354)) and (layer1_outputs(1069)));
    layer2_outputs(325) <= '0';
    layer2_outputs(326) <= not((layer1_outputs(757)) and (layer1_outputs(1302)));
    layer2_outputs(327) <= not(layer1_outputs(1854));
    layer2_outputs(328) <= not((layer1_outputs(2459)) and (layer1_outputs(1186)));
    layer2_outputs(329) <= (layer1_outputs(1860)) and not (layer1_outputs(2143));
    layer2_outputs(330) <= not((layer1_outputs(181)) xor (layer1_outputs(1808)));
    layer2_outputs(331) <= not((layer1_outputs(453)) and (layer1_outputs(99)));
    layer2_outputs(332) <= layer1_outputs(571);
    layer2_outputs(333) <= (layer1_outputs(1343)) or (layer1_outputs(1010));
    layer2_outputs(334) <= not(layer1_outputs(8));
    layer2_outputs(335) <= '0';
    layer2_outputs(336) <= layer1_outputs(1426);
    layer2_outputs(337) <= not((layer1_outputs(408)) and (layer1_outputs(170)));
    layer2_outputs(338) <= (layer1_outputs(872)) and not (layer1_outputs(218));
    layer2_outputs(339) <= '0';
    layer2_outputs(340) <= (layer1_outputs(474)) and (layer1_outputs(1108));
    layer2_outputs(341) <= not((layer1_outputs(2037)) or (layer1_outputs(2242)));
    layer2_outputs(342) <= not(layer1_outputs(27)) or (layer1_outputs(1658));
    layer2_outputs(343) <= (layer1_outputs(1194)) and (layer1_outputs(2339));
    layer2_outputs(344) <= layer1_outputs(1754);
    layer2_outputs(345) <= (layer1_outputs(1733)) or (layer1_outputs(1284));
    layer2_outputs(346) <= not(layer1_outputs(1390)) or (layer1_outputs(31));
    layer2_outputs(347) <= (layer1_outputs(1763)) or (layer1_outputs(1239));
    layer2_outputs(348) <= layer1_outputs(1764);
    layer2_outputs(349) <= layer1_outputs(1000);
    layer2_outputs(350) <= (layer1_outputs(2179)) and not (layer1_outputs(1732));
    layer2_outputs(351) <= (layer1_outputs(1771)) and not (layer1_outputs(1922));
    layer2_outputs(352) <= '1';
    layer2_outputs(353) <= not(layer1_outputs(332));
    layer2_outputs(354) <= '0';
    layer2_outputs(355) <= (layer1_outputs(1084)) and not (layer1_outputs(1057));
    layer2_outputs(356) <= '1';
    layer2_outputs(357) <= (layer1_outputs(804)) or (layer1_outputs(705));
    layer2_outputs(358) <= '1';
    layer2_outputs(359) <= not(layer1_outputs(576)) or (layer1_outputs(1635));
    layer2_outputs(360) <= '1';
    layer2_outputs(361) <= layer1_outputs(445);
    layer2_outputs(362) <= not(layer1_outputs(1981));
    layer2_outputs(363) <= not(layer1_outputs(1646));
    layer2_outputs(364) <= layer1_outputs(2513);
    layer2_outputs(365) <= not(layer1_outputs(1276)) or (layer1_outputs(1074));
    layer2_outputs(366) <= not(layer1_outputs(1726)) or (layer1_outputs(2447));
    layer2_outputs(367) <= (layer1_outputs(153)) and not (layer1_outputs(1878));
    layer2_outputs(368) <= not((layer1_outputs(1659)) and (layer1_outputs(2216)));
    layer2_outputs(369) <= '1';
    layer2_outputs(370) <= (layer1_outputs(1395)) and not (layer1_outputs(347));
    layer2_outputs(371) <= layer1_outputs(810);
    layer2_outputs(372) <= layer1_outputs(183);
    layer2_outputs(373) <= not((layer1_outputs(2039)) xor (layer1_outputs(1047)));
    layer2_outputs(374) <= not((layer1_outputs(784)) and (layer1_outputs(58)));
    layer2_outputs(375) <= (layer1_outputs(23)) and not (layer1_outputs(2316));
    layer2_outputs(376) <= not(layer1_outputs(2018));
    layer2_outputs(377) <= '0';
    layer2_outputs(378) <= not(layer1_outputs(903)) or (layer1_outputs(327));
    layer2_outputs(379) <= not(layer1_outputs(1044)) or (layer1_outputs(1912));
    layer2_outputs(380) <= not(layer1_outputs(903)) or (layer1_outputs(1500));
    layer2_outputs(381) <= not((layer1_outputs(1214)) xor (layer1_outputs(752)));
    layer2_outputs(382) <= not((layer1_outputs(543)) or (layer1_outputs(258)));
    layer2_outputs(383) <= not((layer1_outputs(53)) and (layer1_outputs(889)));
    layer2_outputs(384) <= layer1_outputs(1048);
    layer2_outputs(385) <= layer1_outputs(44);
    layer2_outputs(386) <= '0';
    layer2_outputs(387) <= '0';
    layer2_outputs(388) <= layer1_outputs(321);
    layer2_outputs(389) <= (layer1_outputs(1542)) xor (layer1_outputs(530));
    layer2_outputs(390) <= (layer1_outputs(1034)) and (layer1_outputs(710));
    layer2_outputs(391) <= not((layer1_outputs(2014)) and (layer1_outputs(165)));
    layer2_outputs(392) <= '1';
    layer2_outputs(393) <= '1';
    layer2_outputs(394) <= not(layer1_outputs(373)) or (layer1_outputs(2339));
    layer2_outputs(395) <= not(layer1_outputs(1011)) or (layer1_outputs(1023));
    layer2_outputs(396) <= '1';
    layer2_outputs(397) <= not(layer1_outputs(1269));
    layer2_outputs(398) <= layer1_outputs(1766);
    layer2_outputs(399) <= '0';
    layer2_outputs(400) <= '1';
    layer2_outputs(401) <= not(layer1_outputs(2046));
    layer2_outputs(402) <= not((layer1_outputs(1957)) or (layer1_outputs(1426)));
    layer2_outputs(403) <= layer1_outputs(2530);
    layer2_outputs(404) <= not(layer1_outputs(522)) or (layer1_outputs(1336));
    layer2_outputs(405) <= (layer1_outputs(2064)) and (layer1_outputs(662));
    layer2_outputs(406) <= not(layer1_outputs(2436)) or (layer1_outputs(1769));
    layer2_outputs(407) <= '0';
    layer2_outputs(408) <= not((layer1_outputs(163)) or (layer1_outputs(1187)));
    layer2_outputs(409) <= '0';
    layer2_outputs(410) <= not(layer1_outputs(749));
    layer2_outputs(411) <= layer1_outputs(1951);
    layer2_outputs(412) <= not((layer1_outputs(1935)) and (layer1_outputs(229)));
    layer2_outputs(413) <= (layer1_outputs(626)) and (layer1_outputs(1592));
    layer2_outputs(414) <= '1';
    layer2_outputs(415) <= not(layer1_outputs(177)) or (layer1_outputs(358));
    layer2_outputs(416) <= (layer1_outputs(2290)) or (layer1_outputs(2464));
    layer2_outputs(417) <= '0';
    layer2_outputs(418) <= layer1_outputs(1173);
    layer2_outputs(419) <= '0';
    layer2_outputs(420) <= layer1_outputs(2146);
    layer2_outputs(421) <= '0';
    layer2_outputs(422) <= '1';
    layer2_outputs(423) <= not((layer1_outputs(2181)) and (layer1_outputs(1430)));
    layer2_outputs(424) <= not(layer1_outputs(1262));
    layer2_outputs(425) <= '1';
    layer2_outputs(426) <= '1';
    layer2_outputs(427) <= layer1_outputs(2412);
    layer2_outputs(428) <= not(layer1_outputs(1141));
    layer2_outputs(429) <= (layer1_outputs(1342)) and (layer1_outputs(2321));
    layer2_outputs(430) <= '0';
    layer2_outputs(431) <= layer1_outputs(639);
    layer2_outputs(432) <= layer1_outputs(551);
    layer2_outputs(433) <= '0';
    layer2_outputs(434) <= layer1_outputs(2278);
    layer2_outputs(435) <= not(layer1_outputs(405));
    layer2_outputs(436) <= layer1_outputs(493);
    layer2_outputs(437) <= not(layer1_outputs(1211));
    layer2_outputs(438) <= not(layer1_outputs(1918));
    layer2_outputs(439) <= not((layer1_outputs(1920)) and (layer1_outputs(547)));
    layer2_outputs(440) <= not((layer1_outputs(1268)) and (layer1_outputs(929)));
    layer2_outputs(441) <= (layer1_outputs(2334)) and not (layer1_outputs(2179));
    layer2_outputs(442) <= (layer1_outputs(2079)) and not (layer1_outputs(1958));
    layer2_outputs(443) <= (layer1_outputs(1760)) and (layer1_outputs(290));
    layer2_outputs(444) <= layer1_outputs(148);
    layer2_outputs(445) <= not(layer1_outputs(874));
    layer2_outputs(446) <= (layer1_outputs(1298)) and not (layer1_outputs(1605));
    layer2_outputs(447) <= not(layer1_outputs(977)) or (layer1_outputs(1986));
    layer2_outputs(448) <= '1';
    layer2_outputs(449) <= layer1_outputs(1531);
    layer2_outputs(450) <= layer1_outputs(509);
    layer2_outputs(451) <= not(layer1_outputs(1264)) or (layer1_outputs(2289));
    layer2_outputs(452) <= (layer1_outputs(1917)) or (layer1_outputs(2293));
    layer2_outputs(453) <= '1';
    layer2_outputs(454) <= (layer1_outputs(2211)) and not (layer1_outputs(899));
    layer2_outputs(455) <= (layer1_outputs(1863)) and not (layer1_outputs(501));
    layer2_outputs(456) <= (layer1_outputs(2202)) and not (layer1_outputs(2406));
    layer2_outputs(457) <= not(layer1_outputs(653));
    layer2_outputs(458) <= (layer1_outputs(1115)) and not (layer1_outputs(1002));
    layer2_outputs(459) <= not(layer1_outputs(2138)) or (layer1_outputs(2084));
    layer2_outputs(460) <= not(layer1_outputs(1099)) or (layer1_outputs(1597));
    layer2_outputs(461) <= (layer1_outputs(1936)) and not (layer1_outputs(1392));
    layer2_outputs(462) <= (layer1_outputs(524)) and not (layer1_outputs(484));
    layer2_outputs(463) <= (layer1_outputs(2144)) and (layer1_outputs(806));
    layer2_outputs(464) <= layer1_outputs(742);
    layer2_outputs(465) <= not((layer1_outputs(1121)) or (layer1_outputs(2151)));
    layer2_outputs(466) <= not(layer1_outputs(686));
    layer2_outputs(467) <= not((layer1_outputs(2016)) or (layer1_outputs(629)));
    layer2_outputs(468) <= layer1_outputs(775);
    layer2_outputs(469) <= not(layer1_outputs(898)) or (layer1_outputs(428));
    layer2_outputs(470) <= layer1_outputs(2060);
    layer2_outputs(471) <= (layer1_outputs(891)) and not (layer1_outputs(2293));
    layer2_outputs(472) <= not(layer1_outputs(28)) or (layer1_outputs(1893));
    layer2_outputs(473) <= '1';
    layer2_outputs(474) <= layer1_outputs(2250);
    layer2_outputs(475) <= (layer1_outputs(702)) and (layer1_outputs(2399));
    layer2_outputs(476) <= '1';
    layer2_outputs(477) <= '1';
    layer2_outputs(478) <= '0';
    layer2_outputs(479) <= (layer1_outputs(1578)) or (layer1_outputs(1519));
    layer2_outputs(480) <= layer1_outputs(1681);
    layer2_outputs(481) <= not((layer1_outputs(904)) and (layer1_outputs(2152)));
    layer2_outputs(482) <= not(layer1_outputs(2411));
    layer2_outputs(483) <= layer1_outputs(755);
    layer2_outputs(484) <= layer1_outputs(1574);
    layer2_outputs(485) <= (layer1_outputs(29)) and (layer1_outputs(1320));
    layer2_outputs(486) <= layer1_outputs(2420);
    layer2_outputs(487) <= layer1_outputs(638);
    layer2_outputs(488) <= (layer1_outputs(1968)) or (layer1_outputs(1591));
    layer2_outputs(489) <= (layer1_outputs(401)) and not (layer1_outputs(698));
    layer2_outputs(490) <= (layer1_outputs(879)) or (layer1_outputs(600));
    layer2_outputs(491) <= '1';
    layer2_outputs(492) <= layer1_outputs(316);
    layer2_outputs(493) <= (layer1_outputs(1955)) and not (layer1_outputs(211));
    layer2_outputs(494) <= '0';
    layer2_outputs(495) <= not(layer1_outputs(1380));
    layer2_outputs(496) <= not((layer1_outputs(2217)) or (layer1_outputs(2417)));
    layer2_outputs(497) <= not(layer1_outputs(895)) or (layer1_outputs(2542));
    layer2_outputs(498) <= '0';
    layer2_outputs(499) <= not((layer1_outputs(2344)) and (layer1_outputs(2424)));
    layer2_outputs(500) <= '1';
    layer2_outputs(501) <= (layer1_outputs(1211)) and (layer1_outputs(1032));
    layer2_outputs(502) <= '0';
    layer2_outputs(503) <= layer1_outputs(1423);
    layer2_outputs(504) <= not(layer1_outputs(288)) or (layer1_outputs(1569));
    layer2_outputs(505) <= (layer1_outputs(916)) and (layer1_outputs(2059));
    layer2_outputs(506) <= not((layer1_outputs(382)) and (layer1_outputs(1285)));
    layer2_outputs(507) <= (layer1_outputs(1897)) and not (layer1_outputs(1249));
    layer2_outputs(508) <= (layer1_outputs(1658)) and (layer1_outputs(1772));
    layer2_outputs(509) <= not(layer1_outputs(669));
    layer2_outputs(510) <= layer1_outputs(887);
    layer2_outputs(511) <= '0';
    layer2_outputs(512) <= layer1_outputs(1291);
    layer2_outputs(513) <= (layer1_outputs(122)) xor (layer1_outputs(1262));
    layer2_outputs(514) <= layer1_outputs(1792);
    layer2_outputs(515) <= (layer1_outputs(490)) and not (layer1_outputs(1783));
    layer2_outputs(516) <= not(layer1_outputs(298)) or (layer1_outputs(1505));
    layer2_outputs(517) <= not(layer1_outputs(496));
    layer2_outputs(518) <= '1';
    layer2_outputs(519) <= (layer1_outputs(1276)) or (layer1_outputs(294));
    layer2_outputs(520) <= '1';
    layer2_outputs(521) <= not((layer1_outputs(2269)) or (layer1_outputs(1478)));
    layer2_outputs(522) <= '1';
    layer2_outputs(523) <= (layer1_outputs(326)) or (layer1_outputs(1079));
    layer2_outputs(524) <= '1';
    layer2_outputs(525) <= '1';
    layer2_outputs(526) <= (layer1_outputs(1040)) and (layer1_outputs(2338));
    layer2_outputs(527) <= '0';
    layer2_outputs(528) <= not(layer1_outputs(2065));
    layer2_outputs(529) <= not(layer1_outputs(200)) or (layer1_outputs(409));
    layer2_outputs(530) <= (layer1_outputs(1728)) and not (layer1_outputs(1869));
    layer2_outputs(531) <= not((layer1_outputs(1250)) or (layer1_outputs(1396)));
    layer2_outputs(532) <= (layer1_outputs(263)) and not (layer1_outputs(1421));
    layer2_outputs(533) <= '0';
    layer2_outputs(534) <= not(layer1_outputs(2183)) or (layer1_outputs(1258));
    layer2_outputs(535) <= not(layer1_outputs(1963));
    layer2_outputs(536) <= not(layer1_outputs(2289));
    layer2_outputs(537) <= (layer1_outputs(1784)) or (layer1_outputs(1890));
    layer2_outputs(538) <= not(layer1_outputs(2068));
    layer2_outputs(539) <= '1';
    layer2_outputs(540) <= not(layer1_outputs(2058));
    layer2_outputs(541) <= not(layer1_outputs(930)) or (layer1_outputs(1941));
    layer2_outputs(542) <= layer1_outputs(2520);
    layer2_outputs(543) <= not(layer1_outputs(1406)) or (layer1_outputs(1791));
    layer2_outputs(544) <= not((layer1_outputs(727)) or (layer1_outputs(766)));
    layer2_outputs(545) <= (layer1_outputs(573)) and not (layer1_outputs(1956));
    layer2_outputs(546) <= (layer1_outputs(1482)) and not (layer1_outputs(2475));
    layer2_outputs(547) <= layer1_outputs(856);
    layer2_outputs(548) <= (layer1_outputs(2252)) and not (layer1_outputs(1004));
    layer2_outputs(549) <= '1';
    layer2_outputs(550) <= not(layer1_outputs(874));
    layer2_outputs(551) <= '0';
    layer2_outputs(552) <= '0';
    layer2_outputs(553) <= not(layer1_outputs(2410)) or (layer1_outputs(2232));
    layer2_outputs(554) <= not(layer1_outputs(2175)) or (layer1_outputs(1363));
    layer2_outputs(555) <= not(layer1_outputs(2231));
    layer2_outputs(556) <= not((layer1_outputs(1151)) or (layer1_outputs(1826)));
    layer2_outputs(557) <= '1';
    layer2_outputs(558) <= (layer1_outputs(1012)) and not (layer1_outputs(1209));
    layer2_outputs(559) <= not(layer1_outputs(1640));
    layer2_outputs(560) <= '0';
    layer2_outputs(561) <= not(layer1_outputs(187)) or (layer1_outputs(194));
    layer2_outputs(562) <= '0';
    layer2_outputs(563) <= not((layer1_outputs(1411)) or (layer1_outputs(1309)));
    layer2_outputs(564) <= layer1_outputs(1472);
    layer2_outputs(565) <= (layer1_outputs(1201)) and (layer1_outputs(2125));
    layer2_outputs(566) <= (layer1_outputs(2155)) or (layer1_outputs(531));
    layer2_outputs(567) <= not(layer1_outputs(2249));
    layer2_outputs(568) <= layer1_outputs(2266);
    layer2_outputs(569) <= (layer1_outputs(1181)) and (layer1_outputs(894));
    layer2_outputs(570) <= not((layer1_outputs(1572)) and (layer1_outputs(1476)));
    layer2_outputs(571) <= layer1_outputs(1652);
    layer2_outputs(572) <= not(layer1_outputs(592)) or (layer1_outputs(2267));
    layer2_outputs(573) <= layer1_outputs(1647);
    layer2_outputs(574) <= (layer1_outputs(1675)) and (layer1_outputs(2082));
    layer2_outputs(575) <= '1';
    layer2_outputs(576) <= not((layer1_outputs(112)) and (layer1_outputs(1224)));
    layer2_outputs(577) <= not((layer1_outputs(584)) or (layer1_outputs(7)));
    layer2_outputs(578) <= not(layer1_outputs(1416));
    layer2_outputs(579) <= not(layer1_outputs(323));
    layer2_outputs(580) <= not(layer1_outputs(1013));
    layer2_outputs(581) <= '0';
    layer2_outputs(582) <= not(layer1_outputs(2377));
    layer2_outputs(583) <= layer1_outputs(398);
    layer2_outputs(584) <= not((layer1_outputs(1203)) xor (layer1_outputs(2145)));
    layer2_outputs(585) <= '0';
    layer2_outputs(586) <= '0';
    layer2_outputs(587) <= not((layer1_outputs(1134)) and (layer1_outputs(1738)));
    layer2_outputs(588) <= '0';
    layer2_outputs(589) <= layer1_outputs(1696);
    layer2_outputs(590) <= '1';
    layer2_outputs(591) <= layer1_outputs(1964);
    layer2_outputs(592) <= not(layer1_outputs(886));
    layer2_outputs(593) <= (layer1_outputs(283)) and not (layer1_outputs(683));
    layer2_outputs(594) <= not(layer1_outputs(1056)) or (layer1_outputs(422));
    layer2_outputs(595) <= (layer1_outputs(2205)) and (layer1_outputs(1427));
    layer2_outputs(596) <= '1';
    layer2_outputs(597) <= '1';
    layer2_outputs(598) <= layer1_outputs(1169);
    layer2_outputs(599) <= not(layer1_outputs(1171));
    layer2_outputs(600) <= (layer1_outputs(261)) or (layer1_outputs(2520));
    layer2_outputs(601) <= not(layer1_outputs(1822)) or (layer1_outputs(1432));
    layer2_outputs(602) <= not((layer1_outputs(1853)) and (layer1_outputs(152)));
    layer2_outputs(603) <= (layer1_outputs(2136)) or (layer1_outputs(564));
    layer2_outputs(604) <= not((layer1_outputs(247)) or (layer1_outputs(2100)));
    layer2_outputs(605) <= layer1_outputs(602);
    layer2_outputs(606) <= '1';
    layer2_outputs(607) <= not(layer1_outputs(2168)) or (layer1_outputs(173));
    layer2_outputs(608) <= not(layer1_outputs(2347)) or (layer1_outputs(666));
    layer2_outputs(609) <= not((layer1_outputs(375)) or (layer1_outputs(1389)));
    layer2_outputs(610) <= layer1_outputs(1747);
    layer2_outputs(611) <= '0';
    layer2_outputs(612) <= (layer1_outputs(486)) and not (layer1_outputs(1318));
    layer2_outputs(613) <= layer1_outputs(2275);
    layer2_outputs(614) <= not(layer1_outputs(1525));
    layer2_outputs(615) <= (layer1_outputs(2494)) and (layer1_outputs(1349));
    layer2_outputs(616) <= '1';
    layer2_outputs(617) <= (layer1_outputs(85)) and not (layer1_outputs(2380));
    layer2_outputs(618) <= not((layer1_outputs(1577)) and (layer1_outputs(1116)));
    layer2_outputs(619) <= not((layer1_outputs(298)) or (layer1_outputs(636)));
    layer2_outputs(620) <= not(layer1_outputs(593)) or (layer1_outputs(1722));
    layer2_outputs(621) <= not((layer1_outputs(45)) xor (layer1_outputs(2164)));
    layer2_outputs(622) <= not((layer1_outputs(1715)) or (layer1_outputs(2409)));
    layer2_outputs(623) <= '0';
    layer2_outputs(624) <= '1';
    layer2_outputs(625) <= layer1_outputs(2240);
    layer2_outputs(626) <= (layer1_outputs(1352)) and not (layer1_outputs(184));
    layer2_outputs(627) <= not(layer1_outputs(1203));
    layer2_outputs(628) <= '1';
    layer2_outputs(629) <= not(layer1_outputs(2514));
    layer2_outputs(630) <= layer1_outputs(719);
    layer2_outputs(631) <= not(layer1_outputs(1003));
    layer2_outputs(632) <= not(layer1_outputs(1928)) or (layer1_outputs(573));
    layer2_outputs(633) <= not((layer1_outputs(1939)) and (layer1_outputs(1221)));
    layer2_outputs(634) <= not(layer1_outputs(2428));
    layer2_outputs(635) <= (layer1_outputs(784)) or (layer1_outputs(1033));
    layer2_outputs(636) <= not((layer1_outputs(889)) and (layer1_outputs(920)));
    layer2_outputs(637) <= '1';
    layer2_outputs(638) <= layer1_outputs(631);
    layer2_outputs(639) <= not(layer1_outputs(19));
    layer2_outputs(640) <= layer1_outputs(557);
    layer2_outputs(641) <= (layer1_outputs(705)) and not (layer1_outputs(1275));
    layer2_outputs(642) <= (layer1_outputs(617)) or (layer1_outputs(480));
    layer2_outputs(643) <= layer1_outputs(1320);
    layer2_outputs(644) <= not(layer1_outputs(1888));
    layer2_outputs(645) <= not(layer1_outputs(2152)) or (layer1_outputs(1139));
    layer2_outputs(646) <= not(layer1_outputs(2258)) or (layer1_outputs(1549));
    layer2_outputs(647) <= '0';
    layer2_outputs(648) <= (layer1_outputs(235)) and not (layer1_outputs(2092));
    layer2_outputs(649) <= (layer1_outputs(553)) or (layer1_outputs(1522));
    layer2_outputs(650) <= not((layer1_outputs(783)) or (layer1_outputs(1408)));
    layer2_outputs(651) <= '0';
    layer2_outputs(652) <= (layer1_outputs(80)) and (layer1_outputs(1433));
    layer2_outputs(653) <= '1';
    layer2_outputs(654) <= (layer1_outputs(749)) and (layer1_outputs(1329));
    layer2_outputs(655) <= not(layer1_outputs(1125));
    layer2_outputs(656) <= not((layer1_outputs(867)) and (layer1_outputs(1559)));
    layer2_outputs(657) <= not((layer1_outputs(454)) and (layer1_outputs(47)));
    layer2_outputs(658) <= '1';
    layer2_outputs(659) <= '0';
    layer2_outputs(660) <= layer1_outputs(459);
    layer2_outputs(661) <= not((layer1_outputs(1226)) or (layer1_outputs(2261)));
    layer2_outputs(662) <= (layer1_outputs(433)) and not (layer1_outputs(150));
    layer2_outputs(663) <= not((layer1_outputs(52)) and (layer1_outputs(237)));
    layer2_outputs(664) <= (layer1_outputs(2467)) or (layer1_outputs(1645));
    layer2_outputs(665) <= (layer1_outputs(1761)) and not (layer1_outputs(1002));
    layer2_outputs(666) <= '1';
    layer2_outputs(667) <= not((layer1_outputs(625)) xor (layer1_outputs(1850)));
    layer2_outputs(668) <= not(layer1_outputs(2051)) or (layer1_outputs(972));
    layer2_outputs(669) <= '1';
    layer2_outputs(670) <= layer1_outputs(959);
    layer2_outputs(671) <= (layer1_outputs(2266)) and not (layer1_outputs(1475));
    layer2_outputs(672) <= (layer1_outputs(218)) or (layer1_outputs(893));
    layer2_outputs(673) <= '0';
    layer2_outputs(674) <= layer1_outputs(2159);
    layer2_outputs(675) <= layer1_outputs(1386);
    layer2_outputs(676) <= layer1_outputs(2556);
    layer2_outputs(677) <= (layer1_outputs(1624)) or (layer1_outputs(1061));
    layer2_outputs(678) <= not((layer1_outputs(119)) and (layer1_outputs(49)));
    layer2_outputs(679) <= (layer1_outputs(1595)) and (layer1_outputs(2270));
    layer2_outputs(680) <= '1';
    layer2_outputs(681) <= '0';
    layer2_outputs(682) <= not((layer1_outputs(597)) or (layer1_outputs(747)));
    layer2_outputs(683) <= layer1_outputs(814);
    layer2_outputs(684) <= (layer1_outputs(991)) and not (layer1_outputs(2362));
    layer2_outputs(685) <= not(layer1_outputs(126));
    layer2_outputs(686) <= '1';
    layer2_outputs(687) <= '0';
    layer2_outputs(688) <= not(layer1_outputs(619)) or (layer1_outputs(228));
    layer2_outputs(689) <= '1';
    layer2_outputs(690) <= not((layer1_outputs(1461)) and (layer1_outputs(1111)));
    layer2_outputs(691) <= not((layer1_outputs(375)) and (layer1_outputs(751)));
    layer2_outputs(692) <= '1';
    layer2_outputs(693) <= '1';
    layer2_outputs(694) <= not(layer1_outputs(1288));
    layer2_outputs(695) <= not((layer1_outputs(16)) or (layer1_outputs(264)));
    layer2_outputs(696) <= not((layer1_outputs(343)) and (layer1_outputs(2324)));
    layer2_outputs(697) <= (layer1_outputs(674)) and not (layer1_outputs(568));
    layer2_outputs(698) <= (layer1_outputs(1130)) and not (layer1_outputs(499));
    layer2_outputs(699) <= not(layer1_outputs(843));
    layer2_outputs(700) <= layer1_outputs(2408);
    layer2_outputs(701) <= (layer1_outputs(2517)) and not (layer1_outputs(2330));
    layer2_outputs(702) <= not(layer1_outputs(1600));
    layer2_outputs(703) <= not((layer1_outputs(2397)) and (layer1_outputs(319)));
    layer2_outputs(704) <= '0';
    layer2_outputs(705) <= '0';
    layer2_outputs(706) <= layer1_outputs(1338);
    layer2_outputs(707) <= not((layer1_outputs(368)) or (layer1_outputs(1193)));
    layer2_outputs(708) <= (layer1_outputs(1671)) and not (layer1_outputs(2489));
    layer2_outputs(709) <= '0';
    layer2_outputs(710) <= not((layer1_outputs(1119)) and (layer1_outputs(1321)));
    layer2_outputs(711) <= (layer1_outputs(696)) or (layer1_outputs(1895));
    layer2_outputs(712) <= not(layer1_outputs(2331));
    layer2_outputs(713) <= layer1_outputs(336);
    layer2_outputs(714) <= not(layer1_outputs(737));
    layer2_outputs(715) <= (layer1_outputs(583)) or (layer1_outputs(829));
    layer2_outputs(716) <= not(layer1_outputs(2248)) or (layer1_outputs(2348));
    layer2_outputs(717) <= layer1_outputs(648);
    layer2_outputs(718) <= (layer1_outputs(1843)) and not (layer1_outputs(504));
    layer2_outputs(719) <= (layer1_outputs(440)) and not (layer1_outputs(2087));
    layer2_outputs(720) <= not(layer1_outputs(535));
    layer2_outputs(721) <= (layer1_outputs(162)) and (layer1_outputs(1807));
    layer2_outputs(722) <= (layer1_outputs(1611)) and not (layer1_outputs(2531));
    layer2_outputs(723) <= not(layer1_outputs(1788)) or (layer1_outputs(1676));
    layer2_outputs(724) <= not(layer1_outputs(538)) or (layer1_outputs(1657));
    layer2_outputs(725) <= not((layer1_outputs(169)) and (layer1_outputs(2163)));
    layer2_outputs(726) <= not(layer1_outputs(180)) or (layer1_outputs(988));
    layer2_outputs(727) <= not((layer1_outputs(2420)) xor (layer1_outputs(918)));
    layer2_outputs(728) <= not(layer1_outputs(273)) or (layer1_outputs(1032));
    layer2_outputs(729) <= '0';
    layer2_outputs(730) <= '1';
    layer2_outputs(731) <= '1';
    layer2_outputs(732) <= not((layer1_outputs(106)) and (layer1_outputs(1425)));
    layer2_outputs(733) <= (layer1_outputs(155)) and not (layer1_outputs(120));
    layer2_outputs(734) <= '0';
    layer2_outputs(735) <= not(layer1_outputs(380)) or (layer1_outputs(1859));
    layer2_outputs(736) <= layer1_outputs(1623);
    layer2_outputs(737) <= not((layer1_outputs(1295)) and (layer1_outputs(597)));
    layer2_outputs(738) <= '0';
    layer2_outputs(739) <= '1';
    layer2_outputs(740) <= not(layer1_outputs(569)) or (layer1_outputs(790));
    layer2_outputs(741) <= not(layer1_outputs(0)) or (layer1_outputs(206));
    layer2_outputs(742) <= not(layer1_outputs(1302)) or (layer1_outputs(1256));
    layer2_outputs(743) <= not(layer1_outputs(1632));
    layer2_outputs(744) <= layer1_outputs(2263);
    layer2_outputs(745) <= layer1_outputs(2488);
    layer2_outputs(746) <= not(layer1_outputs(1507)) or (layer1_outputs(2148));
    layer2_outputs(747) <= (layer1_outputs(117)) and (layer1_outputs(503));
    layer2_outputs(748) <= not((layer1_outputs(1509)) and (layer1_outputs(2083)));
    layer2_outputs(749) <= not(layer1_outputs(1261)) or (layer1_outputs(1269));
    layer2_outputs(750) <= '1';
    layer2_outputs(751) <= not(layer1_outputs(833)) or (layer1_outputs(1545));
    layer2_outputs(752) <= '0';
    layer2_outputs(753) <= not(layer1_outputs(304)) or (layer1_outputs(1341));
    layer2_outputs(754) <= '0';
    layer2_outputs(755) <= (layer1_outputs(270)) and (layer1_outputs(1950));
    layer2_outputs(756) <= not(layer1_outputs(1742));
    layer2_outputs(757) <= not(layer1_outputs(1797));
    layer2_outputs(758) <= not(layer1_outputs(1977));
    layer2_outputs(759) <= (layer1_outputs(915)) and not (layer1_outputs(2521));
    layer2_outputs(760) <= not(layer1_outputs(1762));
    layer2_outputs(761) <= layer1_outputs(902);
    layer2_outputs(762) <= layer1_outputs(2112);
    layer2_outputs(763) <= '1';
    layer2_outputs(764) <= (layer1_outputs(866)) and not (layer1_outputs(1874));
    layer2_outputs(765) <= not(layer1_outputs(2227)) or (layer1_outputs(1619));
    layer2_outputs(766) <= (layer1_outputs(528)) and (layer1_outputs(2465));
    layer2_outputs(767) <= not(layer1_outputs(1503)) or (layer1_outputs(2442));
    layer2_outputs(768) <= not((layer1_outputs(281)) and (layer1_outputs(1307)));
    layer2_outputs(769) <= (layer1_outputs(1929)) and not (layer1_outputs(2317));
    layer2_outputs(770) <= layer1_outputs(549);
    layer2_outputs(771) <= (layer1_outputs(299)) and (layer1_outputs(2437));
    layer2_outputs(772) <= not(layer1_outputs(1397));
    layer2_outputs(773) <= not((layer1_outputs(892)) xor (layer1_outputs(951)));
    layer2_outputs(774) <= layer1_outputs(2074);
    layer2_outputs(775) <= not(layer1_outputs(1580));
    layer2_outputs(776) <= not(layer1_outputs(2155)) or (layer1_outputs(479));
    layer2_outputs(777) <= not(layer1_outputs(2052));
    layer2_outputs(778) <= (layer1_outputs(728)) or (layer1_outputs(2545));
    layer2_outputs(779) <= layer1_outputs(1811);
    layer2_outputs(780) <= (layer1_outputs(1439)) and not (layer1_outputs(1846));
    layer2_outputs(781) <= '1';
    layer2_outputs(782) <= not(layer1_outputs(1948));
    layer2_outputs(783) <= '0';
    layer2_outputs(784) <= '1';
    layer2_outputs(785) <= not((layer1_outputs(59)) and (layer1_outputs(942)));
    layer2_outputs(786) <= layer1_outputs(1633);
    layer2_outputs(787) <= not(layer1_outputs(1960)) or (layer1_outputs(207));
    layer2_outputs(788) <= (layer1_outputs(2167)) and not (layer1_outputs(922));
    layer2_outputs(789) <= '0';
    layer2_outputs(790) <= (layer1_outputs(2257)) or (layer1_outputs(1648));
    layer2_outputs(791) <= '1';
    layer2_outputs(792) <= not(layer1_outputs(2078)) or (layer1_outputs(2352));
    layer2_outputs(793) <= layer1_outputs(2301);
    layer2_outputs(794) <= (layer1_outputs(531)) and (layer1_outputs(565));
    layer2_outputs(795) <= not((layer1_outputs(431)) and (layer1_outputs(1099)));
    layer2_outputs(796) <= (layer1_outputs(1711)) and not (layer1_outputs(1172));
    layer2_outputs(797) <= not(layer1_outputs(1290));
    layer2_outputs(798) <= (layer1_outputs(1111)) and (layer1_outputs(2061));
    layer2_outputs(799) <= not((layer1_outputs(1556)) and (layer1_outputs(986)));
    layer2_outputs(800) <= (layer1_outputs(244)) and not (layer1_outputs(1915));
    layer2_outputs(801) <= '1';
    layer2_outputs(802) <= not(layer1_outputs(2));
    layer2_outputs(803) <= (layer1_outputs(2414)) and (layer1_outputs(1385));
    layer2_outputs(804) <= '0';
    layer2_outputs(805) <= not(layer1_outputs(851));
    layer2_outputs(806) <= layer1_outputs(528);
    layer2_outputs(807) <= layer1_outputs(236);
    layer2_outputs(808) <= (layer1_outputs(1471)) and (layer1_outputs(130));
    layer2_outputs(809) <= (layer1_outputs(2024)) and (layer1_outputs(557));
    layer2_outputs(810) <= '1';
    layer2_outputs(811) <= not(layer1_outputs(1765));
    layer2_outputs(812) <= layer1_outputs(2545);
    layer2_outputs(813) <= not(layer1_outputs(1554));
    layer2_outputs(814) <= not(layer1_outputs(968)) or (layer1_outputs(2009));
    layer2_outputs(815) <= layer1_outputs(159);
    layer2_outputs(816) <= (layer1_outputs(2220)) or (layer1_outputs(1448));
    layer2_outputs(817) <= not(layer1_outputs(892)) or (layer1_outputs(145));
    layer2_outputs(818) <= not(layer1_outputs(966));
    layer2_outputs(819) <= not(layer1_outputs(1280));
    layer2_outputs(820) <= layer1_outputs(478);
    layer2_outputs(821) <= not(layer1_outputs(881)) or (layer1_outputs(2316));
    layer2_outputs(822) <= layer1_outputs(1216);
    layer2_outputs(823) <= not(layer1_outputs(513));
    layer2_outputs(824) <= (layer1_outputs(2271)) and not (layer1_outputs(451));
    layer2_outputs(825) <= layer1_outputs(128);
    layer2_outputs(826) <= not(layer1_outputs(549));
    layer2_outputs(827) <= not((layer1_outputs(2040)) and (layer1_outputs(1991)));
    layer2_outputs(828) <= (layer1_outputs(432)) or (layer1_outputs(1418));
    layer2_outputs(829) <= '0';
    layer2_outputs(830) <= '0';
    layer2_outputs(831) <= (layer1_outputs(414)) and not (layer1_outputs(970));
    layer2_outputs(832) <= not((layer1_outputs(1554)) and (layer1_outputs(1871)));
    layer2_outputs(833) <= '0';
    layer2_outputs(834) <= not((layer1_outputs(189)) xor (layer1_outputs(2234)));
    layer2_outputs(835) <= (layer1_outputs(1537)) and not (layer1_outputs(2228));
    layer2_outputs(836) <= '1';
    layer2_outputs(837) <= not(layer1_outputs(546));
    layer2_outputs(838) <= (layer1_outputs(1101)) and (layer1_outputs(1348));
    layer2_outputs(839) <= not(layer1_outputs(2044));
    layer2_outputs(840) <= not(layer1_outputs(224));
    layer2_outputs(841) <= not((layer1_outputs(127)) or (layer1_outputs(66)));
    layer2_outputs(842) <= (layer1_outputs(1007)) and (layer1_outputs(628));
    layer2_outputs(843) <= not(layer1_outputs(1206));
    layer2_outputs(844) <= '1';
    layer2_outputs(845) <= not(layer1_outputs(1180)) or (layer1_outputs(359));
    layer2_outputs(846) <= (layer1_outputs(2555)) and (layer1_outputs(2062));
    layer2_outputs(847) <= (layer1_outputs(1639)) and not (layer1_outputs(1677));
    layer2_outputs(848) <= not((layer1_outputs(2031)) or (layer1_outputs(642)));
    layer2_outputs(849) <= not(layer1_outputs(1736));
    layer2_outputs(850) <= (layer1_outputs(951)) and not (layer1_outputs(1408));
    layer2_outputs(851) <= not(layer1_outputs(865)) or (layer1_outputs(797));
    layer2_outputs(852) <= (layer1_outputs(84)) xor (layer1_outputs(1167));
    layer2_outputs(853) <= layer1_outputs(47);
    layer2_outputs(854) <= layer1_outputs(813);
    layer2_outputs(855) <= not(layer1_outputs(1273)) or (layer1_outputs(1755));
    layer2_outputs(856) <= not(layer1_outputs(443));
    layer2_outputs(857) <= layer1_outputs(571);
    layer2_outputs(858) <= '1';
    layer2_outputs(859) <= not(layer1_outputs(960));
    layer2_outputs(860) <= '1';
    layer2_outputs(861) <= layer1_outputs(1683);
    layer2_outputs(862) <= layer1_outputs(169);
    layer2_outputs(863) <= not(layer1_outputs(1845)) or (layer1_outputs(39));
    layer2_outputs(864) <= (layer1_outputs(453)) or (layer1_outputs(716));
    layer2_outputs(865) <= layer1_outputs(2170);
    layer2_outputs(866) <= (layer1_outputs(676)) and not (layer1_outputs(1593));
    layer2_outputs(867) <= (layer1_outputs(844)) and not (layer1_outputs(1764));
    layer2_outputs(868) <= layer1_outputs(2514);
    layer2_outputs(869) <= layer1_outputs(115);
    layer2_outputs(870) <= not(layer1_outputs(738)) or (layer1_outputs(1927));
    layer2_outputs(871) <= not(layer1_outputs(1235)) or (layer1_outputs(809));
    layer2_outputs(872) <= layer1_outputs(1634);
    layer2_outputs(873) <= not(layer1_outputs(2308));
    layer2_outputs(874) <= not(layer1_outputs(1308));
    layer2_outputs(875) <= (layer1_outputs(46)) and not (layer1_outputs(590));
    layer2_outputs(876) <= not(layer1_outputs(896)) or (layer1_outputs(685));
    layer2_outputs(877) <= not(layer1_outputs(2056)) or (layer1_outputs(2025));
    layer2_outputs(878) <= not(layer1_outputs(2221)) or (layer1_outputs(924));
    layer2_outputs(879) <= (layer1_outputs(176)) and not (layer1_outputs(1201));
    layer2_outputs(880) <= not(layer1_outputs(837)) or (layer1_outputs(1040));
    layer2_outputs(881) <= '0';
    layer2_outputs(882) <= not(layer1_outputs(452));
    layer2_outputs(883) <= layer1_outputs(1519);
    layer2_outputs(884) <= layer1_outputs(1192);
    layer2_outputs(885) <= layer1_outputs(1771);
    layer2_outputs(886) <= not(layer1_outputs(24));
    layer2_outputs(887) <= '1';
    layer2_outputs(888) <= (layer1_outputs(739)) and not (layer1_outputs(1812));
    layer2_outputs(889) <= not(layer1_outputs(544)) or (layer1_outputs(2474));
    layer2_outputs(890) <= layer1_outputs(541);
    layer2_outputs(891) <= not(layer1_outputs(1499)) or (layer1_outputs(1809));
    layer2_outputs(892) <= not((layer1_outputs(2290)) or (layer1_outputs(2255)));
    layer2_outputs(893) <= '1';
    layer2_outputs(894) <= not((layer1_outputs(547)) and (layer1_outputs(2473)));
    layer2_outputs(895) <= not((layer1_outputs(280)) or (layer1_outputs(632)));
    layer2_outputs(896) <= not((layer1_outputs(1609)) and (layer1_outputs(1661)));
    layer2_outputs(897) <= not(layer1_outputs(381));
    layer2_outputs(898) <= not((layer1_outputs(1544)) and (layer1_outputs(2053)));
    layer2_outputs(899) <= layer1_outputs(1488);
    layer2_outputs(900) <= (layer1_outputs(894)) and (layer1_outputs(2047));
    layer2_outputs(901) <= layer1_outputs(1667);
    layer2_outputs(902) <= '0';
    layer2_outputs(903) <= not((layer1_outputs(2080)) or (layer1_outputs(201)));
    layer2_outputs(904) <= layer1_outputs(1748);
    layer2_outputs(905) <= not(layer1_outputs(699)) or (layer1_outputs(1483));
    layer2_outputs(906) <= (layer1_outputs(1085)) or (layer1_outputs(1933));
    layer2_outputs(907) <= not((layer1_outputs(1947)) and (layer1_outputs(331)));
    layer2_outputs(908) <= not(layer1_outputs(322));
    layer2_outputs(909) <= (layer1_outputs(1758)) and not (layer1_outputs(594));
    layer2_outputs(910) <= not((layer1_outputs(61)) and (layer1_outputs(1482)));
    layer2_outputs(911) <= (layer1_outputs(805)) and not (layer1_outputs(990));
    layer2_outputs(912) <= layer1_outputs(602);
    layer2_outputs(913) <= not(layer1_outputs(386)) or (layer1_outputs(206));
    layer2_outputs(914) <= layer1_outputs(2343);
    layer2_outputs(915) <= (layer1_outputs(643)) and (layer1_outputs(2133));
    layer2_outputs(916) <= not(layer1_outputs(1454)) or (layer1_outputs(1720));
    layer2_outputs(917) <= (layer1_outputs(839)) or (layer1_outputs(936));
    layer2_outputs(918) <= (layer1_outputs(1488)) and not (layer1_outputs(73));
    layer2_outputs(919) <= (layer1_outputs(2020)) or (layer1_outputs(687));
    layer2_outputs(920) <= layer1_outputs(2069);
    layer2_outputs(921) <= not(layer1_outputs(2502));
    layer2_outputs(922) <= '1';
    layer2_outputs(923) <= (layer1_outputs(1184)) and not (layer1_outputs(905));
    layer2_outputs(924) <= not((layer1_outputs(1719)) or (layer1_outputs(1029)));
    layer2_outputs(925) <= '1';
    layer2_outputs(926) <= not(layer1_outputs(1664));
    layer2_outputs(927) <= '0';
    layer2_outputs(928) <= '1';
    layer2_outputs(929) <= (layer1_outputs(1750)) xor (layer1_outputs(2134));
    layer2_outputs(930) <= '1';
    layer2_outputs(931) <= layer1_outputs(429);
    layer2_outputs(932) <= not(layer1_outputs(2283));
    layer2_outputs(933) <= '0';
    layer2_outputs(934) <= (layer1_outputs(244)) and not (layer1_outputs(1555));
    layer2_outputs(935) <= not((layer1_outputs(2213)) xor (layer1_outputs(72)));
    layer2_outputs(936) <= not(layer1_outputs(1563)) or (layer1_outputs(1987));
    layer2_outputs(937) <= '1';
    layer2_outputs(938) <= not(layer1_outputs(774)) or (layer1_outputs(333));
    layer2_outputs(939) <= layer1_outputs(2065);
    layer2_outputs(940) <= (layer1_outputs(1132)) or (layer1_outputs(1573));
    layer2_outputs(941) <= not(layer1_outputs(1558)) or (layer1_outputs(685));
    layer2_outputs(942) <= not(layer1_outputs(2002));
    layer2_outputs(943) <= '1';
    layer2_outputs(944) <= not(layer1_outputs(526));
    layer2_outputs(945) <= not(layer1_outputs(474)) or (layer1_outputs(689));
    layer2_outputs(946) <= layer1_outputs(1945);
    layer2_outputs(947) <= layer1_outputs(1801);
    layer2_outputs(948) <= '1';
    layer2_outputs(949) <= (layer1_outputs(252)) and (layer1_outputs(4));
    layer2_outputs(950) <= not((layer1_outputs(282)) and (layer1_outputs(1405)));
    layer2_outputs(951) <= not(layer1_outputs(1504));
    layer2_outputs(952) <= not(layer1_outputs(726));
    layer2_outputs(953) <= not(layer1_outputs(400)) or (layer1_outputs(223));
    layer2_outputs(954) <= '1';
    layer2_outputs(955) <= not(layer1_outputs(32));
    layer2_outputs(956) <= '0';
    layer2_outputs(957) <= not((layer1_outputs(1799)) or (layer1_outputs(1880)));
    layer2_outputs(958) <= layer1_outputs(743);
    layer2_outputs(959) <= not(layer1_outputs(487)) or (layer1_outputs(2408));
    layer2_outputs(960) <= layer1_outputs(715);
    layer2_outputs(961) <= '1';
    layer2_outputs(962) <= layer1_outputs(2166);
    layer2_outputs(963) <= not(layer1_outputs(1729));
    layer2_outputs(964) <= (layer1_outputs(1215)) and not (layer1_outputs(1837));
    layer2_outputs(965) <= not(layer1_outputs(2187)) or (layer1_outputs(2127));
    layer2_outputs(966) <= not(layer1_outputs(420)) or (layer1_outputs(594));
    layer2_outputs(967) <= '0';
    layer2_outputs(968) <= layer1_outputs(2397);
    layer2_outputs(969) <= '0';
    layer2_outputs(970) <= not(layer1_outputs(2304)) or (layer1_outputs(421));
    layer2_outputs(971) <= not((layer1_outputs(158)) and (layer1_outputs(848)));
    layer2_outputs(972) <= not(layer1_outputs(199));
    layer2_outputs(973) <= (layer1_outputs(502)) or (layer1_outputs(777));
    layer2_outputs(974) <= not(layer1_outputs(927));
    layer2_outputs(975) <= not(layer1_outputs(2333));
    layer2_outputs(976) <= (layer1_outputs(1853)) and not (layer1_outputs(1371));
    layer2_outputs(977) <= layer1_outputs(1481);
    layer2_outputs(978) <= not((layer1_outputs(1550)) or (layer1_outputs(175)));
    layer2_outputs(979) <= not((layer1_outputs(864)) and (layer1_outputs(2389)));
    layer2_outputs(980) <= not((layer1_outputs(2426)) or (layer1_outputs(1144)));
    layer2_outputs(981) <= not(layer1_outputs(238)) or (layer1_outputs(246));
    layer2_outputs(982) <= layer1_outputs(2086);
    layer2_outputs(983) <= (layer1_outputs(2178)) and (layer1_outputs(1088));
    layer2_outputs(984) <= not(layer1_outputs(1493));
    layer2_outputs(985) <= not((layer1_outputs(234)) or (layer1_outputs(1196)));
    layer2_outputs(986) <= (layer1_outputs(449)) and not (layer1_outputs(1932));
    layer2_outputs(987) <= (layer1_outputs(562)) and not (layer1_outputs(863));
    layer2_outputs(988) <= '1';
    layer2_outputs(989) <= not((layer1_outputs(1832)) or (layer1_outputs(826)));
    layer2_outputs(990) <= not(layer1_outputs(1672)) or (layer1_outputs(1530));
    layer2_outputs(991) <= layer1_outputs(1784);
    layer2_outputs(992) <= '1';
    layer2_outputs(993) <= '1';
    layer2_outputs(994) <= '1';
    layer2_outputs(995) <= not((layer1_outputs(1667)) and (layer1_outputs(1060)));
    layer2_outputs(996) <= (layer1_outputs(2268)) and not (layer1_outputs(1244));
    layer2_outputs(997) <= not((layer1_outputs(511)) and (layer1_outputs(1547)));
    layer2_outputs(998) <= not((layer1_outputs(1376)) or (layer1_outputs(1297)));
    layer2_outputs(999) <= not((layer1_outputs(1025)) and (layer1_outputs(1400)));
    layer2_outputs(1000) <= (layer1_outputs(1844)) and (layer1_outputs(2508));
    layer2_outputs(1001) <= (layer1_outputs(1221)) and not (layer1_outputs(2118));
    layer2_outputs(1002) <= not(layer1_outputs(2097)) or (layer1_outputs(1170));
    layer2_outputs(1003) <= (layer1_outputs(1311)) xor (layer1_outputs(1767));
    layer2_outputs(1004) <= layer1_outputs(958);
    layer2_outputs(1005) <= (layer1_outputs(772)) or (layer1_outputs(2241));
    layer2_outputs(1006) <= (layer1_outputs(2320)) and (layer1_outputs(1284));
    layer2_outputs(1007) <= not(layer1_outputs(2195)) or (layer1_outputs(2075));
    layer2_outputs(1008) <= not((layer1_outputs(1806)) and (layer1_outputs(20)));
    layer2_outputs(1009) <= not(layer1_outputs(2525));
    layer2_outputs(1010) <= layer1_outputs(2104);
    layer2_outputs(1011) <= not(layer1_outputs(1297)) or (layer1_outputs(2053));
    layer2_outputs(1012) <= (layer1_outputs(782)) and (layer1_outputs(1965));
    layer2_outputs(1013) <= not(layer1_outputs(381));
    layer2_outputs(1014) <= not(layer1_outputs(1098)) or (layer1_outputs(578));
    layer2_outputs(1015) <= layer1_outputs(803);
    layer2_outputs(1016) <= not(layer1_outputs(2103));
    layer2_outputs(1017) <= not(layer1_outputs(771)) or (layer1_outputs(1851));
    layer2_outputs(1018) <= (layer1_outputs(1483)) and not (layer1_outputs(429));
    layer2_outputs(1019) <= layer1_outputs(1943);
    layer2_outputs(1020) <= not((layer1_outputs(2108)) and (layer1_outputs(423)));
    layer2_outputs(1021) <= (layer1_outputs(107)) and not (layer1_outputs(910));
    layer2_outputs(1022) <= (layer1_outputs(931)) or (layer1_outputs(2332));
    layer2_outputs(1023) <= not(layer1_outputs(788));
    layer2_outputs(1024) <= '0';
    layer2_outputs(1025) <= layer1_outputs(396);
    layer2_outputs(1026) <= layer1_outputs(1938);
    layer2_outputs(1027) <= '0';
    layer2_outputs(1028) <= '1';
    layer2_outputs(1029) <= layer1_outputs(1441);
    layer2_outputs(1030) <= layer1_outputs(15);
    layer2_outputs(1031) <= not((layer1_outputs(770)) or (layer1_outputs(2206)));
    layer2_outputs(1032) <= '1';
    layer2_outputs(1033) <= not(layer1_outputs(1345));
    layer2_outputs(1034) <= not(layer1_outputs(828));
    layer2_outputs(1035) <= layer1_outputs(2069);
    layer2_outputs(1036) <= layer1_outputs(1323);
    layer2_outputs(1037) <= not(layer1_outputs(480));
    layer2_outputs(1038) <= not((layer1_outputs(2500)) and (layer1_outputs(1984)));
    layer2_outputs(1039) <= (layer1_outputs(962)) or (layer1_outputs(2345));
    layer2_outputs(1040) <= (layer1_outputs(96)) and not (layer1_outputs(827));
    layer2_outputs(1041) <= layer1_outputs(171);
    layer2_outputs(1042) <= not((layer1_outputs(1904)) and (layer1_outputs(1907)));
    layer2_outputs(1043) <= layer1_outputs(2439);
    layer2_outputs(1044) <= not((layer1_outputs(1531)) or (layer1_outputs(2328)));
    layer2_outputs(1045) <= (layer1_outputs(1980)) and not (layer1_outputs(129));
    layer2_outputs(1046) <= '1';
    layer2_outputs(1047) <= layer1_outputs(87);
    layer2_outputs(1048) <= '0';
    layer2_outputs(1049) <= layer1_outputs(1086);
    layer2_outputs(1050) <= not(layer1_outputs(551));
    layer2_outputs(1051) <= (layer1_outputs(1375)) and (layer1_outputs(1533));
    layer2_outputs(1052) <= not(layer1_outputs(38));
    layer2_outputs(1053) <= '1';
    layer2_outputs(1054) <= not((layer1_outputs(698)) or (layer1_outputs(1962)));
    layer2_outputs(1055) <= layer1_outputs(587);
    layer2_outputs(1056) <= (layer1_outputs(2059)) and (layer1_outputs(1000));
    layer2_outputs(1057) <= layer1_outputs(67);
    layer2_outputs(1058) <= '0';
    layer2_outputs(1059) <= '0';
    layer2_outputs(1060) <= layer1_outputs(1959);
    layer2_outputs(1061) <= '1';
    layer2_outputs(1062) <= layer1_outputs(1977);
    layer2_outputs(1063) <= not((layer1_outputs(1884)) and (layer1_outputs(2556)));
    layer2_outputs(1064) <= not(layer1_outputs(1351));
    layer2_outputs(1065) <= not(layer1_outputs(2262)) or (layer1_outputs(1496));
    layer2_outputs(1066) <= not(layer1_outputs(2050));
    layer2_outputs(1067) <= (layer1_outputs(2329)) and (layer1_outputs(233));
    layer2_outputs(1068) <= (layer1_outputs(1875)) and not (layer1_outputs(1059));
    layer2_outputs(1069) <= not((layer1_outputs(937)) or (layer1_outputs(113)));
    layer2_outputs(1070) <= not(layer1_outputs(2209)) or (layer1_outputs(2147));
    layer2_outputs(1071) <= (layer1_outputs(707)) and not (layer1_outputs(268));
    layer2_outputs(1072) <= layer1_outputs(2385);
    layer2_outputs(1073) <= layer1_outputs(391);
    layer2_outputs(1074) <= '0';
    layer2_outputs(1075) <= layer1_outputs(643);
    layer2_outputs(1076) <= not((layer1_outputs(1756)) or (layer1_outputs(289)));
    layer2_outputs(1077) <= not(layer1_outputs(668));
    layer2_outputs(1078) <= not(layer1_outputs(2429));
    layer2_outputs(1079) <= layer1_outputs(1303);
    layer2_outputs(1080) <= (layer1_outputs(2441)) or (layer1_outputs(1685));
    layer2_outputs(1081) <= not(layer1_outputs(123));
    layer2_outputs(1082) <= layer1_outputs(309);
    layer2_outputs(1083) <= not((layer1_outputs(2532)) and (layer1_outputs(605)));
    layer2_outputs(1084) <= layer1_outputs(2318);
    layer2_outputs(1085) <= '1';
    layer2_outputs(1086) <= not((layer1_outputs(351)) and (layer1_outputs(1923)));
    layer2_outputs(1087) <= not(layer1_outputs(406)) or (layer1_outputs(1305));
    layer2_outputs(1088) <= not((layer1_outputs(542)) or (layer1_outputs(1121)));
    layer2_outputs(1089) <= not(layer1_outputs(1979));
    layer2_outputs(1090) <= layer1_outputs(1896);
    layer2_outputs(1091) <= not(layer1_outputs(460)) or (layer1_outputs(1983));
    layer2_outputs(1092) <= '1';
    layer2_outputs(1093) <= (layer1_outputs(847)) and (layer1_outputs(258));
    layer2_outputs(1094) <= not(layer1_outputs(979));
    layer2_outputs(1095) <= layer1_outputs(143);
    layer2_outputs(1096) <= not(layer1_outputs(1080));
    layer2_outputs(1097) <= layer1_outputs(1687);
    layer2_outputs(1098) <= not(layer1_outputs(1627));
    layer2_outputs(1099) <= '1';
    layer2_outputs(1100) <= '1';
    layer2_outputs(1101) <= '1';
    layer2_outputs(1102) <= not(layer1_outputs(608));
    layer2_outputs(1103) <= not((layer1_outputs(1908)) or (layer1_outputs(1940)));
    layer2_outputs(1104) <= (layer1_outputs(473)) and not (layer1_outputs(1164));
    layer2_outputs(1105) <= not(layer1_outputs(2021)) or (layer1_outputs(1070));
    layer2_outputs(1106) <= (layer1_outputs(1439)) and not (layer1_outputs(2186));
    layer2_outputs(1107) <= '1';
    layer2_outputs(1108) <= not(layer1_outputs(1690));
    layer2_outputs(1109) <= '1';
    layer2_outputs(1110) <= layer1_outputs(2285);
    layer2_outputs(1111) <= '0';
    layer2_outputs(1112) <= '1';
    layer2_outputs(1113) <= not((layer1_outputs(1606)) or (layer1_outputs(2084)));
    layer2_outputs(1114) <= layer1_outputs(1029);
    layer2_outputs(1115) <= (layer1_outputs(290)) and not (layer1_outputs(74));
    layer2_outputs(1116) <= (layer1_outputs(1210)) and (layer1_outputs(1364));
    layer2_outputs(1117) <= '0';
    layer2_outputs(1118) <= layer1_outputs(1544);
    layer2_outputs(1119) <= (layer1_outputs(1660)) and not (layer1_outputs(1381));
    layer2_outputs(1120) <= not((layer1_outputs(17)) xor (layer1_outputs(1102)));
    layer2_outputs(1121) <= not(layer1_outputs(1877)) or (layer1_outputs(410));
    layer2_outputs(1122) <= layer1_outputs(620);
    layer2_outputs(1123) <= '0';
    layer2_outputs(1124) <= not((layer1_outputs(940)) or (layer1_outputs(1213)));
    layer2_outputs(1125) <= '1';
    layer2_outputs(1126) <= layer1_outputs(2278);
    layer2_outputs(1127) <= not((layer1_outputs(1335)) or (layer1_outputs(1938)));
    layer2_outputs(1128) <= not(layer1_outputs(984));
    layer2_outputs(1129) <= '0';
    layer2_outputs(1130) <= (layer1_outputs(1749)) and (layer1_outputs(305));
    layer2_outputs(1131) <= '0';
    layer2_outputs(1132) <= '1';
    layer2_outputs(1133) <= '1';
    layer2_outputs(1134) <= not((layer1_outputs(2196)) or (layer1_outputs(1996)));
    layer2_outputs(1135) <= (layer1_outputs(2386)) or (layer1_outputs(1705));
    layer2_outputs(1136) <= layer1_outputs(2333);
    layer2_outputs(1137) <= not(layer1_outputs(2403)) or (layer1_outputs(812));
    layer2_outputs(1138) <= '0';
    layer2_outputs(1139) <= '1';
    layer2_outputs(1140) <= '0';
    layer2_outputs(1141) <= (layer1_outputs(1123)) and not (layer1_outputs(2509));
    layer2_outputs(1142) <= (layer1_outputs(809)) and not (layer1_outputs(754));
    layer2_outputs(1143) <= not(layer1_outputs(1989)) or (layer1_outputs(1689));
    layer2_outputs(1144) <= layer1_outputs(483);
    layer2_outputs(1145) <= '0';
    layer2_outputs(1146) <= (layer1_outputs(2280)) and not (layer1_outputs(1097));
    layer2_outputs(1147) <= not(layer1_outputs(2342));
    layer2_outputs(1148) <= not((layer1_outputs(94)) and (layer1_outputs(2161)));
    layer2_outputs(1149) <= (layer1_outputs(461)) and (layer1_outputs(1159));
    layer2_outputs(1150) <= (layer1_outputs(1741)) xor (layer1_outputs(2215));
    layer2_outputs(1151) <= layer1_outputs(1397);
    layer2_outputs(1152) <= (layer1_outputs(2117)) and (layer1_outputs(1594));
    layer2_outputs(1153) <= not(layer1_outputs(670));
    layer2_outputs(1154) <= not((layer1_outputs(1775)) or (layer1_outputs(1997)));
    layer2_outputs(1155) <= layer1_outputs(920);
    layer2_outputs(1156) <= '1';
    layer2_outputs(1157) <= layer1_outputs(456);
    layer2_outputs(1158) <= (layer1_outputs(2323)) and not (layer1_outputs(425));
    layer2_outputs(1159) <= (layer1_outputs(2426)) and not (layer1_outputs(622));
    layer2_outputs(1160) <= not(layer1_outputs(88)) or (layer1_outputs(1310));
    layer2_outputs(1161) <= not(layer1_outputs(2026)) or (layer1_outputs(2260));
    layer2_outputs(1162) <= '0';
    layer2_outputs(1163) <= not((layer1_outputs(1109)) and (layer1_outputs(539)));
    layer2_outputs(1164) <= (layer1_outputs(846)) and not (layer1_outputs(667));
    layer2_outputs(1165) <= not(layer1_outputs(473));
    layer2_outputs(1166) <= layer1_outputs(2000);
    layer2_outputs(1167) <= '1';
    layer2_outputs(1168) <= layer1_outputs(982);
    layer2_outputs(1169) <= not(layer1_outputs(168));
    layer2_outputs(1170) <= (layer1_outputs(1994)) and not (layer1_outputs(731));
    layer2_outputs(1171) <= (layer1_outputs(2338)) and not (layer1_outputs(1505));
    layer2_outputs(1172) <= not(layer1_outputs(896)) or (layer1_outputs(975));
    layer2_outputs(1173) <= '1';
    layer2_outputs(1174) <= layer1_outputs(346);
    layer2_outputs(1175) <= layer1_outputs(2541);
    layer2_outputs(1176) <= (layer1_outputs(428)) or (layer1_outputs(2302));
    layer2_outputs(1177) <= (layer1_outputs(2002)) or (layer1_outputs(1245));
    layer2_outputs(1178) <= (layer1_outputs(579)) and not (layer1_outputs(2522));
    layer2_outputs(1179) <= layer1_outputs(1229);
    layer2_outputs(1180) <= layer1_outputs(1345);
    layer2_outputs(1181) <= not((layer1_outputs(1608)) or (layer1_outputs(1573)));
    layer2_outputs(1182) <= not((layer1_outputs(1785)) and (layer1_outputs(2476)));
    layer2_outputs(1183) <= not(layer1_outputs(93));
    layer2_outputs(1184) <= layer1_outputs(1021);
    layer2_outputs(1185) <= not(layer1_outputs(1612)) or (layer1_outputs(921));
    layer2_outputs(1186) <= '1';
    layer2_outputs(1187) <= '0';
    layer2_outputs(1188) <= layer1_outputs(2210);
    layer2_outputs(1189) <= not(layer1_outputs(1197));
    layer2_outputs(1190) <= not(layer1_outputs(1829)) or (layer1_outputs(101));
    layer2_outputs(1191) <= not(layer1_outputs(2418));
    layer2_outputs(1192) <= not((layer1_outputs(2480)) and (layer1_outputs(1528)));
    layer2_outputs(1193) <= (layer1_outputs(1665)) and not (layer1_outputs(2117));
    layer2_outputs(1194) <= layer1_outputs(279);
    layer2_outputs(1195) <= not(layer1_outputs(1157));
    layer2_outputs(1196) <= '0';
    layer2_outputs(1197) <= not((layer1_outputs(780)) and (layer1_outputs(1900)));
    layer2_outputs(1198) <= not(layer1_outputs(1140));
    layer2_outputs(1199) <= not((layer1_outputs(1582)) or (layer1_outputs(1064)));
    layer2_outputs(1200) <= not(layer1_outputs(155)) or (layer1_outputs(663));
    layer2_outputs(1201) <= layer1_outputs(1513);
    layer2_outputs(1202) <= '0';
    layer2_outputs(1203) <= not(layer1_outputs(641));
    layer2_outputs(1204) <= not(layer1_outputs(2548)) or (layer1_outputs(1188));
    layer2_outputs(1205) <= '1';
    layer2_outputs(1206) <= (layer1_outputs(1182)) and not (layer1_outputs(1174));
    layer2_outputs(1207) <= not(layer1_outputs(129));
    layer2_outputs(1208) <= (layer1_outputs(1442)) or (layer1_outputs(946));
    layer2_outputs(1209) <= layer1_outputs(1130);
    layer2_outputs(1210) <= not(layer1_outputs(2049));
    layer2_outputs(1211) <= not((layer1_outputs(2037)) or (layer1_outputs(1688)));
    layer2_outputs(1212) <= not(layer1_outputs(2394)) or (layer1_outputs(1739));
    layer2_outputs(1213) <= not(layer1_outputs(847));
    layer2_outputs(1214) <= (layer1_outputs(1407)) and not (layer1_outputs(2291));
    layer2_outputs(1215) <= layer1_outputs(498);
    layer2_outputs(1216) <= not(layer1_outputs(463));
    layer2_outputs(1217) <= (layer1_outputs(2165)) and not (layer1_outputs(334));
    layer2_outputs(1218) <= (layer1_outputs(1635)) or (layer1_outputs(1649));
    layer2_outputs(1219) <= '0';
    layer2_outputs(1220) <= layer1_outputs(754);
    layer2_outputs(1221) <= not(layer1_outputs(958));
    layer2_outputs(1222) <= '1';
    layer2_outputs(1223) <= not((layer1_outputs(2369)) and (layer1_outputs(1045)));
    layer2_outputs(1224) <= not(layer1_outputs(497));
    layer2_outputs(1225) <= (layer1_outputs(962)) or (layer1_outputs(1495));
    layer2_outputs(1226) <= not((layer1_outputs(781)) or (layer1_outputs(468)));
    layer2_outputs(1227) <= not(layer1_outputs(785)) or (layer1_outputs(1899));
    layer2_outputs(1228) <= layer1_outputs(1532);
    layer2_outputs(1229) <= (layer1_outputs(1675)) or (layer1_outputs(699));
    layer2_outputs(1230) <= not(layer1_outputs(589)) or (layer1_outputs(710));
    layer2_outputs(1231) <= not((layer1_outputs(1152)) or (layer1_outputs(488)));
    layer2_outputs(1232) <= layer1_outputs(2547);
    layer2_outputs(1233) <= '1';
    layer2_outputs(1234) <= not((layer1_outputs(1260)) and (layer1_outputs(1786)));
    layer2_outputs(1235) <= not(layer1_outputs(885)) or (layer1_outputs(980));
    layer2_outputs(1236) <= not(layer1_outputs(1873));
    layer2_outputs(1237) <= '0';
    layer2_outputs(1238) <= not(layer1_outputs(1331));
    layer2_outputs(1239) <= '1';
    layer2_outputs(1240) <= not(layer1_outputs(1273)) or (layer1_outputs(1402));
    layer2_outputs(1241) <= layer1_outputs(2171);
    layer2_outputs(1242) <= '1';
    layer2_outputs(1243) <= '0';
    layer2_outputs(1244) <= not((layer1_outputs(153)) or (layer1_outputs(2340)));
    layer2_outputs(1245) <= '0';
    layer2_outputs(1246) <= not((layer1_outputs(431)) and (layer1_outputs(1447)));
    layer2_outputs(1247) <= not(layer1_outputs(1804));
    layer2_outputs(1248) <= (layer1_outputs(580)) and (layer1_outputs(95));
    layer2_outputs(1249) <= not(layer1_outputs(525));
    layer2_outputs(1250) <= '1';
    layer2_outputs(1251) <= layer1_outputs(1798);
    layer2_outputs(1252) <= (layer1_outputs(1325)) or (layer1_outputs(1384));
    layer2_outputs(1253) <= not((layer1_outputs(1864)) and (layer1_outputs(607)));
    layer2_outputs(1254) <= not(layer1_outputs(741)) or (layer1_outputs(1327));
    layer2_outputs(1255) <= not(layer1_outputs(1247));
    layer2_outputs(1256) <= not(layer1_outputs(588)) or (layer1_outputs(436));
    layer2_outputs(1257) <= (layer1_outputs(2392)) and not (layer1_outputs(271));
    layer2_outputs(1258) <= '1';
    layer2_outputs(1259) <= not(layer1_outputs(580));
    layer2_outputs(1260) <= not(layer1_outputs(1293)) or (layer1_outputs(193));
    layer2_outputs(1261) <= layer1_outputs(126);
    layer2_outputs(1262) <= '0';
    layer2_outputs(1263) <= layer1_outputs(322);
    layer2_outputs(1264) <= layer1_outputs(575);
    layer2_outputs(1265) <= not(layer1_outputs(1818));
    layer2_outputs(1266) <= (layer1_outputs(1031)) and not (layer1_outputs(1966));
    layer2_outputs(1267) <= not((layer1_outputs(22)) and (layer1_outputs(91)));
    layer2_outputs(1268) <= (layer1_outputs(1362)) and not (layer1_outputs(2310));
    layer2_outputs(1269) <= '0';
    layer2_outputs(1270) <= not(layer1_outputs(1400));
    layer2_outputs(1271) <= '0';
    layer2_outputs(1272) <= (layer1_outputs(842)) or (layer1_outputs(546));
    layer2_outputs(1273) <= layer1_outputs(1691);
    layer2_outputs(1274) <= layer1_outputs(1662);
    layer2_outputs(1275) <= not(layer1_outputs(2284));
    layer2_outputs(1276) <= not(layer1_outputs(1146));
    layer2_outputs(1277) <= not(layer1_outputs(823));
    layer2_outputs(1278) <= '0';
    layer2_outputs(1279) <= (layer1_outputs(1651)) xor (layer1_outputs(1975));
    layer2_outputs(1280) <= '0';
    layer2_outputs(1281) <= (layer1_outputs(1575)) and not (layer1_outputs(994));
    layer2_outputs(1282) <= (layer1_outputs(621)) and not (layer1_outputs(2119));
    layer2_outputs(1283) <= not(layer1_outputs(805));
    layer2_outputs(1284) <= not(layer1_outputs(2260)) or (layer1_outputs(1929));
    layer2_outputs(1285) <= not(layer1_outputs(335)) or (layer1_outputs(853));
    layer2_outputs(1286) <= (layer1_outputs(1253)) and not (layer1_outputs(256));
    layer2_outputs(1287) <= '1';
    layer2_outputs(1288) <= not((layer1_outputs(834)) xor (layer1_outputs(2035)));
    layer2_outputs(1289) <= not(layer1_outputs(990));
    layer2_outputs(1290) <= not(layer1_outputs(786));
    layer2_outputs(1291) <= layer1_outputs(2431);
    layer2_outputs(1292) <= (layer1_outputs(1386)) or (layer1_outputs(2354));
    layer2_outputs(1293) <= '1';
    layer2_outputs(1294) <= not((layer1_outputs(566)) and (layer1_outputs(2259)));
    layer2_outputs(1295) <= layer1_outputs(1427);
    layer2_outputs(1296) <= '0';
    layer2_outputs(1297) <= (layer1_outputs(1020)) and not (layer1_outputs(1));
    layer2_outputs(1298) <= not((layer1_outputs(1072)) or (layer1_outputs(2100)));
    layer2_outputs(1299) <= not((layer1_outputs(1490)) xor (layer1_outputs(1722)));
    layer2_outputs(1300) <= layer1_outputs(1992);
    layer2_outputs(1301) <= not(layer1_outputs(2300)) or (layer1_outputs(505));
    layer2_outputs(1302) <= '0';
    layer2_outputs(1303) <= '0';
    layer2_outputs(1304) <= layer1_outputs(1744);
    layer2_outputs(1305) <= (layer1_outputs(890)) or (layer1_outputs(1506));
    layer2_outputs(1306) <= (layer1_outputs(297)) or (layer1_outputs(1061));
    layer2_outputs(1307) <= (layer1_outputs(2098)) and (layer1_outputs(2088));
    layer2_outputs(1308) <= not((layer1_outputs(211)) or (layer1_outputs(1572)));
    layer2_outputs(1309) <= not(layer1_outputs(721)) or (layer1_outputs(1742));
    layer2_outputs(1310) <= not(layer1_outputs(2011));
    layer2_outputs(1311) <= not(layer1_outputs(1441)) or (layer1_outputs(2144));
    layer2_outputs(1312) <= '1';
    layer2_outputs(1313) <= layer1_outputs(1071);
    layer2_outputs(1314) <= (layer1_outputs(1050)) and not (layer1_outputs(1833));
    layer2_outputs(1315) <= (layer1_outputs(66)) xor (layer1_outputs(1999));
    layer2_outputs(1316) <= '0';
    layer2_outputs(1317) <= not(layer1_outputs(1068));
    layer2_outputs(1318) <= not(layer1_outputs(1042)) or (layer1_outputs(1622));
    layer2_outputs(1319) <= not(layer1_outputs(1491)) or (layer1_outputs(2206));
    layer2_outputs(1320) <= not(layer1_outputs(1800)) or (layer1_outputs(1817));
    layer2_outputs(1321) <= '0';
    layer2_outputs(1322) <= not((layer1_outputs(1138)) or (layer1_outputs(41)));
    layer2_outputs(1323) <= not(layer1_outputs(704)) or (layer1_outputs(2330));
    layer2_outputs(1324) <= (layer1_outputs(2074)) and not (layer1_outputs(253));
    layer2_outputs(1325) <= layer1_outputs(349);
    layer2_outputs(1326) <= not(layer1_outputs(1180));
    layer2_outputs(1327) <= '1';
    layer2_outputs(1328) <= layer1_outputs(1047);
    layer2_outputs(1329) <= not(layer1_outputs(247)) or (layer1_outputs(632));
    layer2_outputs(1330) <= '1';
    layer2_outputs(1331) <= (layer1_outputs(1789)) and (layer1_outputs(1599));
    layer2_outputs(1332) <= layer1_outputs(1107);
    layer2_outputs(1333) <= not(layer1_outputs(214)) or (layer1_outputs(2063));
    layer2_outputs(1334) <= '0';
    layer2_outputs(1335) <= (layer1_outputs(1270)) or (layer1_outputs(2367));
    layer2_outputs(1336) <= not(layer1_outputs(1103));
    layer2_outputs(1337) <= not(layer1_outputs(2458));
    layer2_outputs(1338) <= not(layer1_outputs(1455)) or (layer1_outputs(1730));
    layer2_outputs(1339) <= not(layer1_outputs(2032));
    layer2_outputs(1340) <= layer1_outputs(506);
    layer2_outputs(1341) <= layer1_outputs(520);
    layer2_outputs(1342) <= not((layer1_outputs(438)) or (layer1_outputs(1560)));
    layer2_outputs(1343) <= not((layer1_outputs(891)) and (layer1_outputs(64)));
    layer2_outputs(1344) <= '1';
    layer2_outputs(1345) <= layer1_outputs(832);
    layer2_outputs(1346) <= (layer1_outputs(791)) or (layer1_outputs(796));
    layer2_outputs(1347) <= not(layer1_outputs(1437)) or (layer1_outputs(305));
    layer2_outputs(1348) <= not(layer1_outputs(859)) or (layer1_outputs(1389));
    layer2_outputs(1349) <= not(layer1_outputs(2366)) or (layer1_outputs(1851));
    layer2_outputs(1350) <= layer1_outputs(159);
    layer2_outputs(1351) <= (layer1_outputs(2189)) and not (layer1_outputs(2207));
    layer2_outputs(1352) <= not(layer1_outputs(849)) or (layer1_outputs(494));
    layer2_outputs(1353) <= (layer1_outputs(359)) and not (layer1_outputs(973));
    layer2_outputs(1354) <= '0';
    layer2_outputs(1355) <= (layer1_outputs(1602)) and not (layer1_outputs(823));
    layer2_outputs(1356) <= (layer1_outputs(425)) or (layer1_outputs(2186));
    layer2_outputs(1357) <= not(layer1_outputs(505));
    layer2_outputs(1358) <= not((layer1_outputs(2471)) or (layer1_outputs(2343)));
    layer2_outputs(1359) <= not(layer1_outputs(5));
    layer2_outputs(1360) <= not(layer1_outputs(1903));
    layer2_outputs(1361) <= layer1_outputs(1728);
    layer2_outputs(1362) <= not(layer1_outputs(2421));
    layer2_outputs(1363) <= (layer1_outputs(333)) and (layer1_outputs(1144));
    layer2_outputs(1364) <= not((layer1_outputs(471)) xor (layer1_outputs(1372)));
    layer2_outputs(1365) <= not(layer1_outputs(1433)) or (layer1_outputs(506));
    layer2_outputs(1366) <= layer1_outputs(2013);
    layer2_outputs(1367) <= '1';
    layer2_outputs(1368) <= (layer1_outputs(1014)) and not (layer1_outputs(2381));
    layer2_outputs(1369) <= not((layer1_outputs(143)) or (layer1_outputs(1598)));
    layer2_outputs(1370) <= layer1_outputs(1997);
    layer2_outputs(1371) <= '0';
    layer2_outputs(1372) <= not(layer1_outputs(1059));
    layer2_outputs(1373) <= layer1_outputs(1311);
    layer2_outputs(1374) <= layer1_outputs(1881);
    layer2_outputs(1375) <= not(layer1_outputs(377)) or (layer1_outputs(76));
    layer2_outputs(1376) <= (layer1_outputs(691)) and not (layer1_outputs(864));
    layer2_outputs(1377) <= '1';
    layer2_outputs(1378) <= layer1_outputs(1326);
    layer2_outputs(1379) <= layer1_outputs(793);
    layer2_outputs(1380) <= not((layer1_outputs(1393)) and (layer1_outputs(307)));
    layer2_outputs(1381) <= '1';
    layer2_outputs(1382) <= (layer1_outputs(584)) and not (layer1_outputs(212));
    layer2_outputs(1383) <= not(layer1_outputs(2490));
    layer2_outputs(1384) <= '1';
    layer2_outputs(1385) <= layer1_outputs(1231);
    layer2_outputs(1386) <= (layer1_outputs(95)) or (layer1_outputs(172));
    layer2_outputs(1387) <= (layer1_outputs(56)) or (layer1_outputs(2450));
    layer2_outputs(1388) <= '1';
    layer2_outputs(1389) <= not((layer1_outputs(2442)) or (layer1_outputs(548)));
    layer2_outputs(1390) <= layer1_outputs(1462);
    layer2_outputs(1391) <= not(layer1_outputs(790)) or (layer1_outputs(923));
    layer2_outputs(1392) <= not((layer1_outputs(780)) or (layer1_outputs(1467)));
    layer2_outputs(1393) <= (layer1_outputs(1428)) and not (layer1_outputs(1618));
    layer2_outputs(1394) <= '1';
    layer2_outputs(1395) <= '0';
    layer2_outputs(1396) <= '0';
    layer2_outputs(1397) <= (layer1_outputs(511)) and not (layer1_outputs(2522));
    layer2_outputs(1398) <= not(layer1_outputs(446)) or (layer1_outputs(1346));
    layer2_outputs(1399) <= not(layer1_outputs(415));
    layer2_outputs(1400) <= '0';
    layer2_outputs(1401) <= not(layer1_outputs(620));
    layer2_outputs(1402) <= '1';
    layer2_outputs(1403) <= not(layer1_outputs(1796));
    layer2_outputs(1404) <= (layer1_outputs(633)) or (layer1_outputs(430));
    layer2_outputs(1405) <= not(layer1_outputs(2536)) or (layer1_outputs(1186));
    layer2_outputs(1406) <= '0';
    layer2_outputs(1407) <= (layer1_outputs(200)) and not (layer1_outputs(1534));
    layer2_outputs(1408) <= '1';
    layer2_outputs(1409) <= not((layer1_outputs(2140)) or (layer1_outputs(2105)));
    layer2_outputs(1410) <= '0';
    layer2_outputs(1411) <= not((layer1_outputs(1757)) xor (layer1_outputs(928)));
    layer2_outputs(1412) <= '1';
    layer2_outputs(1413) <= not(layer1_outputs(1412));
    layer2_outputs(1414) <= layer1_outputs(1991);
    layer2_outputs(1415) <= layer1_outputs(589);
    layer2_outputs(1416) <= not((layer1_outputs(1219)) and (layer1_outputs(2474)));
    layer2_outputs(1417) <= not(layer1_outputs(2376));
    layer2_outputs(1418) <= not(layer1_outputs(2300));
    layer2_outputs(1419) <= layer1_outputs(78);
    layer2_outputs(1420) <= not((layer1_outputs(2140)) or (layer1_outputs(2501)));
    layer2_outputs(1421) <= not((layer1_outputs(2156)) or (layer1_outputs(2009)));
    layer2_outputs(1422) <= not((layer1_outputs(672)) and (layer1_outputs(1348)));
    layer2_outputs(1423) <= not(layer1_outputs(829)) or (layer1_outputs(1127));
    layer2_outputs(1424) <= not((layer1_outputs(134)) xor (layer1_outputs(2444)));
    layer2_outputs(1425) <= (layer1_outputs(1898)) and not (layer1_outputs(1900));
    layer2_outputs(1426) <= not(layer1_outputs(802));
    layer2_outputs(1427) <= not(layer1_outputs(1617));
    layer2_outputs(1428) <= '0';
    layer2_outputs(1429) <= not(layer1_outputs(725)) or (layer1_outputs(388));
    layer2_outputs(1430) <= (layer1_outputs(1569)) and (layer1_outputs(552));
    layer2_outputs(1431) <= layer1_outputs(604);
    layer2_outputs(1432) <= not((layer1_outputs(1497)) and (layer1_outputs(2477)));
    layer2_outputs(1433) <= '0';
    layer2_outputs(1434) <= (layer1_outputs(2515)) or (layer1_outputs(2279));
    layer2_outputs(1435) <= '0';
    layer2_outputs(1436) <= layer1_outputs(537);
    layer2_outputs(1437) <= (layer1_outputs(1834)) and not (layer1_outputs(2131));
    layer2_outputs(1438) <= not(layer1_outputs(1005));
    layer2_outputs(1439) <= not(layer1_outputs(1972));
    layer2_outputs(1440) <= '1';
    layer2_outputs(1441) <= (layer1_outputs(1469)) xor (layer1_outputs(11));
    layer2_outputs(1442) <= (layer1_outputs(1637)) and (layer1_outputs(283));
    layer2_outputs(1443) <= (layer1_outputs(408)) and not (layer1_outputs(2482));
    layer2_outputs(1444) <= layer1_outputs(849);
    layer2_outputs(1445) <= not(layer1_outputs(2114)) or (layer1_outputs(413));
    layer2_outputs(1446) <= layer1_outputs(2502);
    layer2_outputs(1447) <= not(layer1_outputs(2544)) or (layer1_outputs(2412));
    layer2_outputs(1448) <= layer1_outputs(2415);
    layer2_outputs(1449) <= not(layer1_outputs(1225));
    layer2_outputs(1450) <= (layer1_outputs(1796)) and (layer1_outputs(2189));
    layer2_outputs(1451) <= not((layer1_outputs(432)) or (layer1_outputs(761)));
    layer2_outputs(1452) <= not(layer1_outputs(1476)) or (layer1_outputs(2468));
    layer2_outputs(1453) <= layer1_outputs(2270);
    layer2_outputs(1454) <= (layer1_outputs(1163)) and not (layer1_outputs(963));
    layer2_outputs(1455) <= layer1_outputs(938);
    layer2_outputs(1456) <= not(layer1_outputs(1540)) or (layer1_outputs(1778));
    layer2_outputs(1457) <= (layer1_outputs(1985)) and (layer1_outputs(216));
    layer2_outputs(1458) <= (layer1_outputs(510)) and (layer1_outputs(120));
    layer2_outputs(1459) <= '1';
    layer2_outputs(1460) <= not(layer1_outputs(1590));
    layer2_outputs(1461) <= (layer1_outputs(1252)) or (layer1_outputs(1016));
    layer2_outputs(1462) <= (layer1_outputs(1541)) and not (layer1_outputs(706));
    layer2_outputs(1463) <= layer1_outputs(1998);
    layer2_outputs(1464) <= not(layer1_outputs(489));
    layer2_outputs(1465) <= not(layer1_outputs(565)) or (layer1_outputs(2250));
    layer2_outputs(1466) <= not((layer1_outputs(2531)) or (layer1_outputs(384)));
    layer2_outputs(1467) <= not(layer1_outputs(2003));
    layer2_outputs(1468) <= (layer1_outputs(1805)) and not (layer1_outputs(2215));
    layer2_outputs(1469) <= (layer1_outputs(2461)) and not (layer1_outputs(70));
    layer2_outputs(1470) <= layer1_outputs(919);
    layer2_outputs(1471) <= not(layer1_outputs(1885));
    layer2_outputs(1472) <= layer1_outputs(1692);
    layer2_outputs(1473) <= not((layer1_outputs(1583)) and (layer1_outputs(826)));
    layer2_outputs(1474) <= '0';
    layer2_outputs(1475) <= '1';
    layer2_outputs(1476) <= layer1_outputs(276);
    layer2_outputs(1477) <= not(layer1_outputs(1395));
    layer2_outputs(1478) <= not(layer1_outputs(1246));
    layer2_outputs(1479) <= '0';
    layer2_outputs(1480) <= '1';
    layer2_outputs(1481) <= (layer1_outputs(2435)) and (layer1_outputs(2350));
    layer2_outputs(1482) <= not((layer1_outputs(536)) and (layer1_outputs(2463)));
    layer2_outputs(1483) <= (layer1_outputs(1416)) or (layer1_outputs(1660));
    layer2_outputs(1484) <= not((layer1_outputs(2185)) and (layer1_outputs(2422)));
    layer2_outputs(1485) <= not(layer1_outputs(426)) or (layer1_outputs(396));
    layer2_outputs(1486) <= '0';
    layer2_outputs(1487) <= not(layer1_outputs(1153));
    layer2_outputs(1488) <= not((layer1_outputs(2013)) and (layer1_outputs(693)));
    layer2_outputs(1489) <= (layer1_outputs(1150)) and not (layer1_outputs(525));
    layer2_outputs(1490) <= not(layer1_outputs(582));
    layer2_outputs(1491) <= not((layer1_outputs(407)) and (layer1_outputs(228)));
    layer2_outputs(1492) <= '1';
    layer2_outputs(1493) <= layer1_outputs(2314);
    layer2_outputs(1494) <= (layer1_outputs(1038)) and not (layer1_outputs(293));
    layer2_outputs(1495) <= not(layer1_outputs(321)) or (layer1_outputs(1231));
    layer2_outputs(1496) <= (layer1_outputs(2549)) or (layer1_outputs(2486));
    layer2_outputs(1497) <= (layer1_outputs(16)) or (layer1_outputs(1905));
    layer2_outputs(1498) <= not(layer1_outputs(1015));
    layer2_outputs(1499) <= '0';
    layer2_outputs(1500) <= '0';
    layer2_outputs(1501) <= layer1_outputs(2264);
    layer2_outputs(1502) <= not(layer1_outputs(1502)) or (layer1_outputs(2188));
    layer2_outputs(1503) <= not(layer1_outputs(67));
    layer2_outputs(1504) <= not((layer1_outputs(758)) and (layer1_outputs(1517)));
    layer2_outputs(1505) <= not(layer1_outputs(1473)) or (layer1_outputs(335));
    layer2_outputs(1506) <= not((layer1_outputs(1636)) and (layer1_outputs(2457)));
    layer2_outputs(1507) <= not((layer1_outputs(287)) or (layer1_outputs(1267)));
    layer2_outputs(1508) <= not((layer1_outputs(2498)) or (layer1_outputs(798)));
    layer2_outputs(1509) <= not((layer1_outputs(1880)) or (layer1_outputs(1374)));
    layer2_outputs(1510) <= not(layer1_outputs(1220));
    layer2_outputs(1511) <= not(layer1_outputs(1043)) or (layer1_outputs(2366));
    layer2_outputs(1512) <= (layer1_outputs(327)) and not (layer1_outputs(2469));
    layer2_outputs(1513) <= not(layer1_outputs(1232));
    layer2_outputs(1514) <= '0';
    layer2_outputs(1515) <= not(layer1_outputs(69));
    layer2_outputs(1516) <= '1';
    layer2_outputs(1517) <= not(layer1_outputs(779));
    layer2_outputs(1518) <= (layer1_outputs(1238)) or (layer1_outputs(697));
    layer2_outputs(1519) <= not(layer1_outputs(502));
    layer2_outputs(1520) <= (layer1_outputs(483)) or (layer1_outputs(1138));
    layer2_outputs(1521) <= not(layer1_outputs(90));
    layer2_outputs(1522) <= '1';
    layer2_outputs(1523) <= not(layer1_outputs(2281)) or (layer1_outputs(1659));
    layer2_outputs(1524) <= (layer1_outputs(1378)) and (layer1_outputs(2245));
    layer2_outputs(1525) <= not(layer1_outputs(419)) or (layer1_outputs(2470));
    layer2_outputs(1526) <= '1';
    layer2_outputs(1527) <= layer1_outputs(2351);
    layer2_outputs(1528) <= layer1_outputs(2478);
    layer2_outputs(1529) <= '0';
    layer2_outputs(1530) <= not((layer1_outputs(769)) and (layer1_outputs(735)));
    layer2_outputs(1531) <= not(layer1_outputs(2387));
    layer2_outputs(1532) <= '1';
    layer2_outputs(1533) <= '0';
    layer2_outputs(1534) <= '0';
    layer2_outputs(1535) <= not((layer1_outputs(225)) or (layer1_outputs(630)));
    layer2_outputs(1536) <= (layer1_outputs(2404)) and (layer1_outputs(1192));
    layer2_outputs(1537) <= not((layer1_outputs(532)) or (layer1_outputs(883)));
    layer2_outputs(1538) <= not((layer1_outputs(2080)) or (layer1_outputs(284)));
    layer2_outputs(1539) <= layer1_outputs(119);
    layer2_outputs(1540) <= not((layer1_outputs(272)) or (layer1_outputs(1607)));
    layer2_outputs(1541) <= (layer1_outputs(2319)) or (layer1_outputs(2296));
    layer2_outputs(1542) <= not((layer1_outputs(1105)) or (layer1_outputs(1943)));
    layer2_outputs(1543) <= (layer1_outputs(25)) and (layer1_outputs(1153));
    layer2_outputs(1544) <= layer1_outputs(1147);
    layer2_outputs(1545) <= (layer1_outputs(1321)) and (layer1_outputs(1377));
    layer2_outputs(1546) <= not(layer1_outputs(2085));
    layer2_outputs(1547) <= '0';
    layer2_outputs(1548) <= '1';
    layer2_outputs(1549) <= not(layer1_outputs(1158)) or (layer1_outputs(357));
    layer2_outputs(1550) <= (layer1_outputs(1918)) and (layer1_outputs(2359));
    layer2_outputs(1551) <= not((layer1_outputs(1682)) and (layer1_outputs(1737)));
    layer2_outputs(1552) <= not((layer1_outputs(1939)) or (layer1_outputs(2222)));
    layer2_outputs(1553) <= layer1_outputs(404);
    layer2_outputs(1554) <= (layer1_outputs(1780)) and (layer1_outputs(558));
    layer2_outputs(1555) <= (layer1_outputs(2105)) and not (layer1_outputs(878));
    layer2_outputs(1556) <= (layer1_outputs(517)) or (layer1_outputs(2256));
    layer2_outputs(1557) <= not(layer1_outputs(1744));
    layer2_outputs(1558) <= not((layer1_outputs(1560)) or (layer1_outputs(1165)));
    layer2_outputs(1559) <= not(layer1_outputs(1281)) or (layer1_outputs(60));
    layer2_outputs(1560) <= (layer1_outputs(606)) or (layer1_outputs(2295));
    layer2_outputs(1561) <= layer1_outputs(637);
    layer2_outputs(1562) <= '1';
    layer2_outputs(1563) <= (layer1_outputs(368)) and (layer1_outputs(1989));
    layer2_outputs(1564) <= (layer1_outputs(800)) and not (layer1_outputs(1252));
    layer2_outputs(1565) <= not((layer1_outputs(68)) or (layer1_outputs(1782)));
    layer2_outputs(1566) <= '0';
    layer2_outputs(1567) <= not((layer1_outputs(2224)) or (layer1_outputs(1526)));
    layer2_outputs(1568) <= '1';
    layer2_outputs(1569) <= not(layer1_outputs(684));
    layer2_outputs(1570) <= '1';
    layer2_outputs(1571) <= not((layer1_outputs(1861)) and (layer1_outputs(108)));
    layer2_outputs(1572) <= '1';
    layer2_outputs(1573) <= (layer1_outputs(2471)) and (layer1_outputs(1976));
    layer2_outputs(1574) <= not(layer1_outputs(320)) or (layer1_outputs(1825));
    layer2_outputs(1575) <= '0';
    layer2_outputs(1576) <= not((layer1_outputs(93)) and (layer1_outputs(2551)));
    layer2_outputs(1577) <= '0';
    layer2_outputs(1578) <= layer1_outputs(1558);
    layer2_outputs(1579) <= not(layer1_outputs(2106)) or (layer1_outputs(2012));
    layer2_outputs(1580) <= '0';
    layer2_outputs(1581) <= not(layer1_outputs(1981));
    layer2_outputs(1582) <= not(layer1_outputs(1263)) or (layer1_outputs(583));
    layer2_outputs(1583) <= not(layer1_outputs(1957));
    layer2_outputs(1584) <= (layer1_outputs(2175)) and not (layer1_outputs(982));
    layer2_outputs(1585) <= (layer1_outputs(1892)) and (layer1_outputs(339));
    layer2_outputs(1586) <= '0';
    layer2_outputs(1587) <= not(layer1_outputs(449));
    layer2_outputs(1588) <= layer1_outputs(83);
    layer2_outputs(1589) <= layer1_outputs(2248);
    layer2_outputs(1590) <= '1';
    layer2_outputs(1591) <= not((layer1_outputs(2253)) and (layer1_outputs(986)));
    layer2_outputs(1592) <= not(layer1_outputs(448));
    layer2_outputs(1593) <= (layer1_outputs(1514)) and not (layer1_outputs(462));
    layer2_outputs(1594) <= not(layer1_outputs(2224));
    layer2_outputs(1595) <= not((layer1_outputs(943)) or (layer1_outputs(1684)));
    layer2_outputs(1596) <= not((layer1_outputs(1607)) and (layer1_outputs(1811)));
    layer2_outputs(1597) <= (layer1_outputs(146)) and not (layer1_outputs(2011));
    layer2_outputs(1598) <= layer1_outputs(463);
    layer2_outputs(1599) <= layer1_outputs(1377);
    layer2_outputs(1600) <= layer1_outputs(1734);
    layer2_outputs(1601) <= not(layer1_outputs(138)) or (layer1_outputs(901));
    layer2_outputs(1602) <= layer1_outputs(1710);
    layer2_outputs(1603) <= not(layer1_outputs(1392)) or (layer1_outputs(1643));
    layer2_outputs(1604) <= not(layer1_outputs(1078)) or (layer1_outputs(1695));
    layer2_outputs(1605) <= '0';
    layer2_outputs(1606) <= not(layer1_outputs(1652)) or (layer1_outputs(1707));
    layer2_outputs(1607) <= not(layer1_outputs(188)) or (layer1_outputs(1902));
    layer2_outputs(1608) <= not((layer1_outputs(139)) and (layer1_outputs(2462)));
    layer2_outputs(1609) <= layer1_outputs(1777);
    layer2_outputs(1610) <= layer1_outputs(497);
    layer2_outputs(1611) <= not(layer1_outputs(636));
    layer2_outputs(1612) <= not(layer1_outputs(646)) or (layer1_outputs(379));
    layer2_outputs(1613) <= not(layer1_outputs(334)) or (layer1_outputs(45));
    layer2_outputs(1614) <= (layer1_outputs(1094)) and (layer1_outputs(2341));
    layer2_outputs(1615) <= not(layer1_outputs(1698)) or (layer1_outputs(1923));
    layer2_outputs(1616) <= '0';
    layer2_outputs(1617) <= (layer1_outputs(362)) and not (layer1_outputs(868));
    layer2_outputs(1618) <= not(layer1_outputs(1199)) or (layer1_outputs(1775));
    layer2_outputs(1619) <= (layer1_outputs(1108)) and (layer1_outputs(132));
    layer2_outputs(1620) <= not(layer1_outputs(2107));
    layer2_outputs(1621) <= not(layer1_outputs(2370));
    layer2_outputs(1622) <= layer1_outputs(2208);
    layer2_outputs(1623) <= '0';
    layer2_outputs(1624) <= '0';
    layer2_outputs(1625) <= (layer1_outputs(297)) xor (layer1_outputs(1279));
    layer2_outputs(1626) <= not((layer1_outputs(1328)) or (layer1_outputs(581)));
    layer2_outputs(1627) <= not(layer1_outputs(543));
    layer2_outputs(1628) <= '1';
    layer2_outputs(1629) <= layer1_outputs(172);
    layer2_outputs(1630) <= '0';
    layer2_outputs(1631) <= not(layer1_outputs(1005)) or (layer1_outputs(2279));
    layer2_outputs(1632) <= not(layer1_outputs(2288)) or (layer1_outputs(1528));
    layer2_outputs(1633) <= not(layer1_outputs(1613)) or (layer1_outputs(1145));
    layer2_outputs(1634) <= layer1_outputs(765);
    layer2_outputs(1635) <= not(layer1_outputs(1357)) or (layer1_outputs(1470));
    layer2_outputs(1636) <= not(layer1_outputs(481));
    layer2_outputs(1637) <= '1';
    layer2_outputs(1638) <= not(layer1_outputs(39)) or (layer1_outputs(550));
    layer2_outputs(1639) <= not(layer1_outputs(1719)) or (layer1_outputs(2052));
    layer2_outputs(1640) <= not(layer1_outputs(481));
    layer2_outputs(1641) <= not(layer1_outputs(434));
    layer2_outputs(1642) <= not(layer1_outputs(2360));
    layer2_outputs(1643) <= layer1_outputs(496);
    layer2_outputs(1644) <= not(layer1_outputs(1840));
    layer2_outputs(1645) <= '1';
    layer2_outputs(1646) <= layer1_outputs(150);
    layer2_outputs(1647) <= not(layer1_outputs(2093));
    layer2_outputs(1648) <= (layer1_outputs(997)) and not (layer1_outputs(1874));
    layer2_outputs(1649) <= not(layer1_outputs(2273)) or (layer1_outputs(470));
    layer2_outputs(1650) <= not(layer1_outputs(1428));
    layer2_outputs(1651) <= layer1_outputs(2519);
    layer2_outputs(1652) <= not((layer1_outputs(683)) or (layer1_outputs(2073)));
    layer2_outputs(1653) <= (layer1_outputs(2004)) and (layer1_outputs(385));
    layer2_outputs(1654) <= '1';
    layer2_outputs(1655) <= not((layer1_outputs(2102)) or (layer1_outputs(82)));
    layer2_outputs(1656) <= not((layer1_outputs(1588)) and (layer1_outputs(2120)));
    layer2_outputs(1657) <= '0';
    layer2_outputs(1658) <= not(layer1_outputs(70));
    layer2_outputs(1659) <= not(layer1_outputs(202)) or (layer1_outputs(956));
    layer2_outputs(1660) <= not(layer1_outputs(523));
    layer2_outputs(1661) <= not(layer1_outputs(2373)) or (layer1_outputs(1627));
    layer2_outputs(1662) <= not(layer1_outputs(587));
    layer2_outputs(1663) <= layer1_outputs(987);
    layer2_outputs(1664) <= layer1_outputs(2174);
    layer2_outputs(1665) <= (layer1_outputs(989)) and not (layer1_outputs(1735));
    layer2_outputs(1666) <= '1';
    layer2_outputs(1667) <= layer1_outputs(1564);
    layer2_outputs(1668) <= layer1_outputs(2372);
    layer2_outputs(1669) <= layer1_outputs(2307);
    layer2_outputs(1670) <= (layer1_outputs(1265)) and (layer1_outputs(1686));
    layer2_outputs(1671) <= layer1_outputs(1290);
    layer2_outputs(1672) <= layer1_outputs(717);
    layer2_outputs(1673) <= (layer1_outputs(740)) and not (layer1_outputs(706));
    layer2_outputs(1674) <= (layer1_outputs(1461)) and not (layer1_outputs(418));
    layer2_outputs(1675) <= not((layer1_outputs(1872)) and (layer1_outputs(1548)));
    layer2_outputs(1676) <= not((layer1_outputs(1604)) or (layer1_outputs(1734)));
    layer2_outputs(1677) <= not(layer1_outputs(309));
    layer2_outputs(1678) <= not(layer1_outputs(1415)) or (layer1_outputs(2301));
    layer2_outputs(1679) <= (layer1_outputs(1490)) and (layer1_outputs(529));
    layer2_outputs(1680) <= '1';
    layer2_outputs(1681) <= (layer1_outputs(544)) and (layer1_outputs(880));
    layer2_outputs(1682) <= (layer1_outputs(2165)) and not (layer1_outputs(585));
    layer2_outputs(1683) <= (layer1_outputs(1436)) and not (layer1_outputs(337));
    layer2_outputs(1684) <= not((layer1_outputs(859)) and (layer1_outputs(1475)));
    layer2_outputs(1685) <= (layer1_outputs(1515)) and not (layer1_outputs(2379));
    layer2_outputs(1686) <= (layer1_outputs(1202)) and (layer1_outputs(111));
    layer2_outputs(1687) <= (layer1_outputs(1459)) and not (layer1_outputs(1829));
    layer2_outputs(1688) <= '1';
    layer2_outputs(1689) <= (layer1_outputs(854)) or (layer1_outputs(1864));
    layer2_outputs(1690) <= (layer1_outputs(1589)) and not (layer1_outputs(1552));
    layer2_outputs(1691) <= not(layer1_outputs(1930));
    layer2_outputs(1692) <= not(layer1_outputs(2546));
    layer2_outputs(1693) <= not(layer1_outputs(1248)) or (layer1_outputs(2110));
    layer2_outputs(1694) <= layer1_outputs(556);
    layer2_outputs(1695) <= not(layer1_outputs(482));
    layer2_outputs(1696) <= (layer1_outputs(1232)) and not (layer1_outputs(2320));
    layer2_outputs(1697) <= not(layer1_outputs(1382));
    layer2_outputs(1698) <= '0';
    layer2_outputs(1699) <= not(layer1_outputs(1213)) or (layer1_outputs(1051));
    layer2_outputs(1700) <= not(layer1_outputs(376));
    layer2_outputs(1701) <= not(layer1_outputs(1365)) or (layer1_outputs(650));
    layer2_outputs(1702) <= not(layer1_outputs(48));
    layer2_outputs(1703) <= '1';
    layer2_outputs(1704) <= not((layer1_outputs(1610)) and (layer1_outputs(981)));
    layer2_outputs(1705) <= not(layer1_outputs(915));
    layer2_outputs(1706) <= layer1_outputs(1524);
    layer2_outputs(1707) <= not((layer1_outputs(819)) and (layer1_outputs(123)));
    layer2_outputs(1708) <= '1';
    layer2_outputs(1709) <= not(layer1_outputs(160));
    layer2_outputs(1710) <= not(layer1_outputs(1));
    layer2_outputs(1711) <= not((layer1_outputs(260)) or (layer1_outputs(99)));
    layer2_outputs(1712) <= layer1_outputs(808);
    layer2_outputs(1713) <= not(layer1_outputs(898));
    layer2_outputs(1714) <= not(layer1_outputs(391)) or (layer1_outputs(1513));
    layer2_outputs(1715) <= (layer1_outputs(1788)) and not (layer1_outputs(2438));
    layer2_outputs(1716) <= not(layer1_outputs(2527));
    layer2_outputs(1717) <= '1';
    layer2_outputs(1718) <= not((layer1_outputs(2141)) or (layer1_outputs(570)));
    layer2_outputs(1719) <= not(layer1_outputs(14));
    layer2_outputs(1720) <= not(layer1_outputs(1650));
    layer2_outputs(1721) <= (layer1_outputs(1358)) or (layer1_outputs(1971));
    layer2_outputs(1722) <= (layer1_outputs(21)) or (layer1_outputs(350));
    layer2_outputs(1723) <= not(layer1_outputs(2303));
    layer2_outputs(1724) <= not(layer1_outputs(541));
    layer2_outputs(1725) <= not(layer1_outputs(1057));
    layer2_outputs(1726) <= layer1_outputs(2504);
    layer2_outputs(1727) <= (layer1_outputs(2077)) and not (layer1_outputs(295));
    layer2_outputs(1728) <= layer1_outputs(1340);
    layer2_outputs(1729) <= '1';
    layer2_outputs(1730) <= not(layer1_outputs(834));
    layer2_outputs(1731) <= (layer1_outputs(270)) and (layer1_outputs(2401));
    layer2_outputs(1732) <= layer1_outputs(197);
    layer2_outputs(1733) <= layer1_outputs(2194);
    layer2_outputs(1734) <= not(layer1_outputs(356));
    layer2_outputs(1735) <= layer1_outputs(1306);
    layer2_outputs(1736) <= '0';
    layer2_outputs(1737) <= not(layer1_outputs(1611)) or (layer1_outputs(2456));
    layer2_outputs(1738) <= not((layer1_outputs(2032)) or (layer1_outputs(2139)));
    layer2_outputs(1739) <= (layer1_outputs(1283)) and not (layer1_outputs(2336));
    layer2_outputs(1740) <= not((layer1_outputs(2110)) or (layer1_outputs(50)));
    layer2_outputs(1741) <= not(layer1_outputs(252)) or (layer1_outputs(2136));
    layer2_outputs(1742) <= not(layer1_outputs(1940));
    layer2_outputs(1743) <= not(layer1_outputs(1993)) or (layer1_outputs(614));
    layer2_outputs(1744) <= '1';
    layer2_outputs(1745) <= not(layer1_outputs(203));
    layer2_outputs(1746) <= layer1_outputs(2547);
    layer2_outputs(1747) <= layer1_outputs(1128);
    layer2_outputs(1748) <= (layer1_outputs(26)) and not (layer1_outputs(2000));
    layer2_outputs(1749) <= (layer1_outputs(2319)) and (layer1_outputs(880));
    layer2_outputs(1750) <= layer1_outputs(1375);
    layer2_outputs(1751) <= (layer1_outputs(345)) and not (layer1_outputs(492));
    layer2_outputs(1752) <= layer1_outputs(1193);
    layer2_outputs(1753) <= '1';
    layer2_outputs(1754) <= layer1_outputs(860);
    layer2_outputs(1755) <= not((layer1_outputs(278)) and (layer1_outputs(2046)));
    layer2_outputs(1756) <= (layer1_outputs(1150)) and not (layer1_outputs(495));
    layer2_outputs(1757) <= (layer1_outputs(1503)) and not (layer1_outputs(196));
    layer2_outputs(1758) <= '0';
    layer2_outputs(1759) <= layer1_outputs(2087);
    layer2_outputs(1760) <= (layer1_outputs(938)) or (layer1_outputs(2455));
    layer2_outputs(1761) <= not(layer1_outputs(422));
    layer2_outputs(1762) <= '0';
    layer2_outputs(1763) <= layer1_outputs(113);
    layer2_outputs(1764) <= not(layer1_outputs(590));
    layer2_outputs(1765) <= not(layer1_outputs(2506));
    layer2_outputs(1766) <= (layer1_outputs(1768)) and not (layer1_outputs(1450));
    layer2_outputs(1767) <= not(layer1_outputs(1206));
    layer2_outputs(1768) <= layer1_outputs(1415);
    layer2_outputs(1769) <= not(layer1_outputs(356)) or (layer1_outputs(625));
    layer2_outputs(1770) <= (layer1_outputs(1535)) and not (layer1_outputs(1053));
    layer2_outputs(1771) <= not(layer1_outputs(732));
    layer2_outputs(1772) <= (layer1_outputs(302)) xor (layer1_outputs(1282));
    layer2_outputs(1773) <= (layer1_outputs(344)) and (layer1_outputs(319));
    layer2_outputs(1774) <= layer1_outputs(1228);
    layer2_outputs(1775) <= layer1_outputs(1493);
    layer2_outputs(1776) <= '0';
    layer2_outputs(1777) <= (layer1_outputs(437)) or (layer1_outputs(292));
    layer2_outputs(1778) <= not(layer1_outputs(1787)) or (layer1_outputs(867));
    layer2_outputs(1779) <= not(layer1_outputs(420));
    layer2_outputs(1780) <= (layer1_outputs(2131)) or (layer1_outputs(967));
    layer2_outputs(1781) <= '0';
    layer2_outputs(1782) <= (layer1_outputs(1931)) and not (layer1_outputs(1291));
    layer2_outputs(1783) <= not(layer1_outputs(1236));
    layer2_outputs(1784) <= '0';
    layer2_outputs(1785) <= (layer1_outputs(736)) or (layer1_outputs(1486));
    layer2_outputs(1786) <= not((layer1_outputs(852)) and (layer1_outputs(778)));
    layer2_outputs(1787) <= layer1_outputs(97);
    layer2_outputs(1788) <= '1';
    layer2_outputs(1789) <= not(layer1_outputs(456)) or (layer1_outputs(1479));
    layer2_outputs(1790) <= '1';
    layer2_outputs(1791) <= '0';
    layer2_outputs(1792) <= (layer1_outputs(1700)) or (layer1_outputs(1924));
    layer2_outputs(1793) <= (layer1_outputs(1691)) and not (layer1_outputs(2127));
    layer2_outputs(1794) <= (layer1_outputs(141)) and not (layer1_outputs(1855));
    layer2_outputs(1795) <= '1';
    layer2_outputs(1796) <= not(layer1_outputs(1904)) or (layer1_outputs(349));
    layer2_outputs(1797) <= not(layer1_outputs(1906)) or (layer1_outputs(1820));
    layer2_outputs(1798) <= '1';
    layer2_outputs(1799) <= (layer1_outputs(1746)) xor (layer1_outputs(1614));
    layer2_outputs(1800) <= not((layer1_outputs(1872)) and (layer1_outputs(2223)));
    layer2_outputs(1801) <= (layer1_outputs(25)) or (layer1_outputs(1510));
    layer2_outputs(1802) <= not(layer1_outputs(1315));
    layer2_outputs(1803) <= not(layer1_outputs(1147)) or (layer1_outputs(1456));
    layer2_outputs(1804) <= layer1_outputs(376);
    layer2_outputs(1805) <= (layer1_outputs(1642)) and not (layer1_outputs(2529));
    layer2_outputs(1806) <= '0';
    layer2_outputs(1807) <= layer1_outputs(816);
    layer2_outputs(1808) <= layer1_outputs(2158);
    layer2_outputs(1809) <= not(layer1_outputs(2259)) or (layer1_outputs(135));
    layer2_outputs(1810) <= not(layer1_outputs(1198)) or (layer1_outputs(1815));
    layer2_outputs(1811) <= (layer1_outputs(1786)) and (layer1_outputs(1883));
    layer2_outputs(1812) <= layer1_outputs(2510);
    layer2_outputs(1813) <= '1';
    layer2_outputs(1814) <= not((layer1_outputs(1914)) xor (layer1_outputs(1725)));
    layer2_outputs(1815) <= not(layer1_outputs(974));
    layer2_outputs(1816) <= '1';
    layer2_outputs(1817) <= (layer1_outputs(836)) or (layer1_outputs(970));
    layer2_outputs(1818) <= not(layer1_outputs(131)) or (layer1_outputs(649));
    layer2_outputs(1819) <= layer1_outputs(1849);
    layer2_outputs(1820) <= not(layer1_outputs(907)) or (layer1_outputs(2125));
    layer2_outputs(1821) <= '1';
    layer2_outputs(1822) <= '1';
    layer2_outputs(1823) <= not((layer1_outputs(277)) and (layer1_outputs(1380)));
    layer2_outputs(1824) <= (layer1_outputs(1666)) and (layer1_outputs(1561));
    layer2_outputs(1825) <= (layer1_outputs(1855)) or (layer1_outputs(1073));
    layer2_outputs(1826) <= not(layer1_outputs(771));
    layer2_outputs(1827) <= not((layer1_outputs(1689)) or (layer1_outputs(1341)));
    layer2_outputs(1828) <= not(layer1_outputs(1846)) or (layer1_outputs(2479));
    layer2_outputs(1829) <= layer1_outputs(703);
    layer2_outputs(1830) <= layer1_outputs(652);
    layer2_outputs(1831) <= not(layer1_outputs(1731)) or (layer1_outputs(2374));
    layer2_outputs(1832) <= layer1_outputs(2516);
    layer2_outputs(1833) <= '0';
    layer2_outputs(1834) <= (layer1_outputs(1740)) and (layer1_outputs(2430));
    layer2_outputs(1835) <= '0';
    layer2_outputs(1836) <= '0';
    layer2_outputs(1837) <= not((layer1_outputs(1300)) or (layer1_outputs(367)));
    layer2_outputs(1838) <= not((layer1_outputs(1736)) or (layer1_outputs(1596)));
    layer2_outputs(1839) <= not(layer1_outputs(671)) or (layer1_outputs(1729));
    layer2_outputs(1840) <= (layer1_outputs(694)) and (layer1_outputs(1417));
    layer2_outputs(1841) <= (layer1_outputs(802)) and not (layer1_outputs(77));
    layer2_outputs(1842) <= '1';
    layer2_outputs(1843) <= layer1_outputs(2287);
    layer2_outputs(1844) <= not(layer1_outputs(1009)) or (layer1_outputs(1446));
    layer2_outputs(1845) <= not((layer1_outputs(14)) or (layer1_outputs(686)));
    layer2_outputs(1846) <= '1';
    layer2_outputs(1847) <= layer1_outputs(1594);
    layer2_outputs(1848) <= not((layer1_outputs(1149)) and (layer1_outputs(220)));
    layer2_outputs(1849) <= not((layer1_outputs(2072)) or (layer1_outputs(1992)));
    layer2_outputs(1850) <= not((layer1_outputs(1810)) or (layer1_outputs(1478)));
    layer2_outputs(1851) <= not(layer1_outputs(952));
    layer2_outputs(1852) <= layer1_outputs(2447);
    layer2_outputs(1853) <= not(layer1_outputs(2158));
    layer2_outputs(1854) <= (layer1_outputs(2023)) or (layer1_outputs(1189));
    layer2_outputs(1855) <= layer1_outputs(1773);
    layer2_outputs(1856) <= layer1_outputs(204);
    layer2_outputs(1857) <= not((layer1_outputs(1509)) and (layer1_outputs(1698)));
    layer2_outputs(1858) <= not(layer1_outputs(645)) or (layer1_outputs(2504));
    layer2_outputs(1859) <= not(layer1_outputs(1907));
    layer2_outputs(1860) <= (layer1_outputs(1003)) and not (layer1_outputs(1463));
    layer2_outputs(1861) <= not((layer1_outputs(262)) or (layer1_outputs(798)));
    layer2_outputs(1862) <= (layer1_outputs(588)) and not (layer1_outputs(1184));
    layer2_outputs(1863) <= (layer1_outputs(720)) xor (layer1_outputs(1404));
    layer2_outputs(1864) <= '1';
    layer2_outputs(1865) <= not((layer1_outputs(1662)) or (layer1_outputs(1191)));
    layer2_outputs(1866) <= (layer1_outputs(1616)) and not (layer1_outputs(2496));
    layer2_outputs(1867) <= not(layer1_outputs(2554));
    layer2_outputs(1868) <= layer1_outputs(2231);
    layer2_outputs(1869) <= not(layer1_outputs(43));
    layer2_outputs(1870) <= (layer1_outputs(1496)) or (layer1_outputs(199));
    layer2_outputs(1871) <= not((layer1_outputs(76)) or (layer1_outputs(2249)));
    layer2_outputs(1872) <= not((layer1_outputs(1858)) and (layer1_outputs(2048)));
    layer2_outputs(1873) <= (layer1_outputs(2022)) and not (layer1_outputs(339));
    layer2_outputs(1874) <= (layer1_outputs(1523)) or (layer1_outputs(2477));
    layer2_outputs(1875) <= (layer1_outputs(178)) and not (layer1_outputs(660));
    layer2_outputs(1876) <= '0';
    layer2_outputs(1877) <= layer1_outputs(734);
    layer2_outputs(1878) <= (layer1_outputs(2008)) and not (layer1_outputs(2067));
    layer2_outputs(1879) <= not(layer1_outputs(395)) or (layer1_outputs(1398));
    layer2_outputs(1880) <= (layer1_outputs(789)) and not (layer1_outputs(2539));
    layer2_outputs(1881) <= not((layer1_outputs(1500)) or (layer1_outputs(1467)));
    layer2_outputs(1882) <= layer1_outputs(245);
    layer2_outputs(1883) <= not(layer1_outputs(2363));
    layer2_outputs(1884) <= not(layer1_outputs(1140));
    layer2_outputs(1885) <= (layer1_outputs(1603)) and not (layer1_outputs(1802));
    layer2_outputs(1886) <= layer1_outputs(2476);
    layer2_outputs(1887) <= (layer1_outputs(1129)) and not (layer1_outputs(641));
    layer2_outputs(1888) <= not((layer1_outputs(156)) and (layer1_outputs(929)));
    layer2_outputs(1889) <= (layer1_outputs(762)) and (layer1_outputs(1747));
    layer2_outputs(1890) <= not((layer1_outputs(1440)) and (layer1_outputs(659)));
    layer2_outputs(1891) <= not(layer1_outputs(182)) or (layer1_outputs(2121));
    layer2_outputs(1892) <= not(layer1_outputs(389));
    layer2_outputs(1893) <= '0';
    layer2_outputs(1894) <= (layer1_outputs(1777)) and not (layer1_outputs(1982));
    layer2_outputs(1895) <= (layer1_outputs(799)) and (layer1_outputs(2349));
    layer2_outputs(1896) <= layer1_outputs(945);
    layer2_outputs(1897) <= (layer1_outputs(659)) or (layer1_outputs(1255));
    layer2_outputs(1898) <= not(layer1_outputs(242));
    layer2_outputs(1899) <= '1';
    layer2_outputs(1900) <= '0';
    layer2_outputs(1901) <= not(layer1_outputs(1547));
    layer2_outputs(1902) <= layer1_outputs(1077);
    layer2_outputs(1903) <= not(layer1_outputs(1210)) or (layer1_outputs(1848));
    layer2_outputs(1904) <= '1';
    layer2_outputs(1905) <= layer1_outputs(455);
    layer2_outputs(1906) <= not((layer1_outputs(772)) or (layer1_outputs(2045)));
    layer2_outputs(1907) <= not((layer1_outputs(219)) and (layer1_outputs(1819)));
    layer2_outputs(1908) <= (layer1_outputs(2022)) and not (layer1_outputs(1919));
    layer2_outputs(1909) <= layer1_outputs(1091);
    layer2_outputs(1910) <= not(layer1_outputs(342)) or (layer1_outputs(1816));
    layer2_outputs(1911) <= (layer1_outputs(835)) and not (layer1_outputs(1543));
    layer2_outputs(1912) <= '1';
    layer2_outputs(1913) <= not(layer1_outputs(2513)) or (layer1_outputs(841));
    layer2_outputs(1914) <= layer1_outputs(973);
    layer2_outputs(1915) <= not((layer1_outputs(36)) or (layer1_outputs(1459)));
    layer2_outputs(1916) <= '0';
    layer2_outputs(1917) <= (layer1_outputs(630)) or (layer1_outputs(1350));
    layer2_outputs(1918) <= not((layer1_outputs(851)) and (layer1_outputs(2055)));
    layer2_outputs(1919) <= layer1_outputs(561);
    layer2_outputs(1920) <= (layer1_outputs(1586)) and (layer1_outputs(2274));
    layer2_outputs(1921) <= layer1_outputs(222);
    layer2_outputs(1922) <= not(layer1_outputs(421));
    layer2_outputs(1923) <= not(layer1_outputs(2005)) or (layer1_outputs(2435));
    layer2_outputs(1924) <= '0';
    layer2_outputs(1925) <= '0';
    layer2_outputs(1926) <= (layer1_outputs(1694)) and not (layer1_outputs(556));
    layer2_outputs(1927) <= '0';
    layer2_outputs(1928) <= '1';
    layer2_outputs(1929) <= not(layer1_outputs(2495)) or (layer1_outputs(2363));
    layer2_outputs(1930) <= layer1_outputs(2393);
    layer2_outputs(1931) <= '1';
    layer2_outputs(1932) <= not(layer1_outputs(2481));
    layer2_outputs(1933) <= '1';
    layer2_outputs(1934) <= (layer1_outputs(1480)) and not (layer1_outputs(2209));
    layer2_outputs(1935) <= '0';
    layer2_outputs(1936) <= '1';
    layer2_outputs(1937) <= layer1_outputs(1508);
    layer2_outputs(1938) <= layer1_outputs(4);
    layer2_outputs(1939) <= not((layer1_outputs(232)) and (layer1_outputs(2303)));
    layer2_outputs(1940) <= '0';
    layer2_outputs(1941) <= '1';
    layer2_outputs(1942) <= layer1_outputs(2040);
    layer2_outputs(1943) <= not((layer1_outputs(116)) and (layer1_outputs(37)));
    layer2_outputs(1944) <= not(layer1_outputs(1979));
    layer2_outputs(1945) <= (layer1_outputs(1158)) or (layer1_outputs(1157));
    layer2_outputs(1946) <= not(layer1_outputs(1789)) or (layer1_outputs(2025));
    layer2_outputs(1947) <= not(layer1_outputs(1570)) or (layer1_outputs(759));
    layer2_outputs(1948) <= not(layer1_outputs(1398));
    layer2_outputs(1949) <= (layer1_outputs(1308)) and not (layer1_outputs(1223));
    layer2_outputs(1950) <= not(layer1_outputs(1774));
    layer2_outputs(1951) <= layer1_outputs(555);
    layer2_outputs(1952) <= '0';
    layer2_outputs(1953) <= not(layer1_outputs(1013)) or (layer1_outputs(1838));
    layer2_outputs(1954) <= '0';
    layer2_outputs(1955) <= '1';
    layer2_outputs(1956) <= not(layer1_outputs(2384)) or (layer1_outputs(1970));
    layer2_outputs(1957) <= not(layer1_outputs(1118));
    layer2_outputs(1958) <= not((layer1_outputs(2349)) or (layer1_outputs(911)));
    layer2_outputs(1959) <= not(layer1_outputs(713)) or (layer1_outputs(92));
    layer2_outputs(1960) <= not(layer1_outputs(1487));
    layer2_outputs(1961) <= layer1_outputs(237);
    layer2_outputs(1962) <= '0';
    layer2_outputs(1963) <= not(layer1_outputs(257));
    layer2_outputs(1964) <= not((layer1_outputs(1098)) or (layer1_outputs(1590)));
    layer2_outputs(1965) <= not(layer1_outputs(2405));
    layer2_outputs(1966) <= not(layer1_outputs(276)) or (layer1_outputs(437));
    layer2_outputs(1967) <= not(layer1_outputs(1871));
    layer2_outputs(1968) <= not(layer1_outputs(917));
    layer2_outputs(1969) <= (layer1_outputs(1253)) and (layer1_outputs(694));
    layer2_outputs(1970) <= not(layer1_outputs(1637));
    layer2_outputs(1971) <= (layer1_outputs(2021)) or (layer1_outputs(210));
    layer2_outputs(1972) <= '0';
    layer2_outputs(1973) <= (layer1_outputs(221)) and not (layer1_outputs(2036));
    layer2_outputs(1974) <= not(layer1_outputs(1941)) or (layer1_outputs(2102));
    layer2_outputs(1975) <= not(layer1_outputs(426)) or (layer1_outputs(2521));
    layer2_outputs(1976) <= (layer1_outputs(2017)) and (layer1_outputs(452));
    layer2_outputs(1977) <= (layer1_outputs(873)) and not (layer1_outputs(1183));
    layer2_outputs(1978) <= layer1_outputs(1329);
    layer2_outputs(1979) <= (layer1_outputs(436)) or (layer1_outputs(369));
    layer2_outputs(1980) <= (layer1_outputs(1803)) and not (layer1_outputs(1674));
    layer2_outputs(1981) <= '0';
    layer2_outputs(1982) <= (layer1_outputs(2123)) or (layer1_outputs(899));
    layer2_outputs(1983) <= '0';
    layer2_outputs(1984) <= not(layer1_outputs(2512)) or (layer1_outputs(993));
    layer2_outputs(1985) <= not(layer1_outputs(753));
    layer2_outputs(1986) <= '0';
    layer2_outputs(1987) <= (layer1_outputs(690)) and (layer1_outputs(946));
    layer2_outputs(1988) <= not(layer1_outputs(37));
    layer2_outputs(1989) <= '0';
    layer2_outputs(1990) <= '0';
    layer2_outputs(1991) <= not(layer1_outputs(1518)) or (layer1_outputs(609));
    layer2_outputs(1992) <= not((layer1_outputs(1056)) or (layer1_outputs(1743)));
    layer2_outputs(1993) <= layer1_outputs(1546);
    layer2_outputs(1994) <= '0';
    layer2_outputs(1995) <= '1';
    layer2_outputs(1996) <= layer1_outputs(1028);
    layer2_outputs(1997) <= not(layer1_outputs(1381));
    layer2_outputs(1998) <= '1';
    layer2_outputs(1999) <= not(layer1_outputs(1953));
    layer2_outputs(2000) <= layer1_outputs(2392);
    layer2_outputs(2001) <= (layer1_outputs(253)) and not (layer1_outputs(482));
    layer2_outputs(2002) <= '1';
    layer2_outputs(2003) <= not(layer1_outputs(55));
    layer2_outputs(2004) <= not((layer1_outputs(1512)) or (layer1_outputs(1812)));
    layer2_outputs(2005) <= layer1_outputs(844);
    layer2_outputs(2006) <= '0';
    layer2_outputs(2007) <= not((layer1_outputs(2253)) or (layer1_outputs(875)));
    layer2_outputs(2008) <= not((layer1_outputs(2200)) and (layer1_outputs(1504)));
    layer2_outputs(2009) <= '1';
    layer2_outputs(2010) <= not(layer1_outputs(1499)) or (layer1_outputs(275));
    layer2_outputs(2011) <= '0';
    layer2_outputs(2012) <= (layer1_outputs(2287)) or (layer1_outputs(492));
    layer2_outputs(2013) <= not(layer1_outputs(2436)) or (layer1_outputs(1237));
    layer2_outputs(2014) <= not(layer1_outputs(2060)) or (layer1_outputs(2526));
    layer2_outputs(2015) <= layer1_outputs(136);
    layer2_outputs(2016) <= (layer1_outputs(1663)) and not (layer1_outputs(2364));
    layer2_outputs(2017) <= not(layer1_outputs(1019)) or (layer1_outputs(103));
    layer2_outputs(2018) <= not(layer1_outputs(0));
    layer2_outputs(2019) <= (layer1_outputs(90)) and (layer1_outputs(909));
    layer2_outputs(2020) <= not(layer1_outputs(1882)) or (layer1_outputs(2039));
    layer2_outputs(2021) <= not(layer1_outputs(2192));
    layer2_outputs(2022) <= '0';
    layer2_outputs(2023) <= '1';
    layer2_outputs(2024) <= not(layer1_outputs(2494)) or (layer1_outputs(1248));
    layer2_outputs(2025) <= layer1_outputs(2444);
    layer2_outputs(2026) <= '0';
    layer2_outputs(2027) <= layer1_outputs(1824);
    layer2_outputs(2028) <= (layer1_outputs(266)) or (layer1_outputs(2066));
    layer2_outputs(2029) <= not(layer1_outputs(2305));
    layer2_outputs(2030) <= (layer1_outputs(624)) or (layer1_outputs(1135));
    layer2_outputs(2031) <= '1';
    layer2_outputs(2032) <= not(layer1_outputs(1673)) or (layer1_outputs(1520));
    layer2_outputs(2033) <= layer1_outputs(1301);
    layer2_outputs(2034) <= (layer1_outputs(1655)) and not (layer1_outputs(1772));
    layer2_outputs(2035) <= not(layer1_outputs(807));
    layer2_outputs(2036) <= not(layer1_outputs(650));
    layer2_outputs(2037) <= layer1_outputs(458);
    layer2_outputs(2038) <= (layer1_outputs(427)) and not (layer1_outputs(231));
    layer2_outputs(2039) <= (layer1_outputs(1017)) xor (layer1_outputs(1091));
    layer2_outputs(2040) <= not(layer1_outputs(813));
    layer2_outputs(2041) <= '0';
    layer2_outputs(2042) <= layer1_outputs(33);
    layer2_outputs(2043) <= (layer1_outputs(695)) or (layer1_outputs(2318));
    layer2_outputs(2044) <= (layer1_outputs(1966)) and not (layer1_outputs(2341));
    layer2_outputs(2045) <= '1';
    layer2_outputs(2046) <= (layer1_outputs(1906)) and not (layer1_outputs(361));
    layer2_outputs(2047) <= not((layer1_outputs(1867)) or (layer1_outputs(835)));
    layer2_outputs(2048) <= not(layer1_outputs(80));
    layer2_outputs(2049) <= (layer1_outputs(934)) and not (layer1_outputs(721));
    layer2_outputs(2050) <= (layer1_outputs(1034)) or (layer1_outputs(2185));
    layer2_outputs(2051) <= not((layer1_outputs(2026)) and (layer1_outputs(1217)));
    layer2_outputs(2052) <= not(layer1_outputs(2219)) or (layer1_outputs(1620));
    layer2_outputs(2053) <= not(layer1_outputs(377)) or (layer1_outputs(905));
    layer2_outputs(2054) <= (layer1_outputs(1278)) and not (layer1_outputs(801));
    layer2_outputs(2055) <= '1';
    layer2_outputs(2056) <= not(layer1_outputs(1360));
    layer2_outputs(2057) <= not(layer1_outputs(739));
    layer2_outputs(2058) <= not(layer1_outputs(782)) or (layer1_outputs(2122));
    layer2_outputs(2059) <= not(layer1_outputs(801));
    layer2_outputs(2060) <= layer1_outputs(324);
    layer2_outputs(2061) <= not((layer1_outputs(1178)) and (layer1_outputs(28)));
    layer2_outputs(2062) <= layer1_outputs(1170);
    layer2_outputs(2063) <= not(layer1_outputs(871));
    layer2_outputs(2064) <= (layer1_outputs(281)) and not (layer1_outputs(928));
    layer2_outputs(2065) <= not(layer1_outputs(1837)) or (layer1_outputs(328));
    layer2_outputs(2066) <= (layer1_outputs(1527)) and not (layer1_outputs(1523));
    layer2_outputs(2067) <= not(layer1_outputs(2537));
    layer2_outputs(2068) <= (layer1_outputs(2466)) and (layer1_outputs(1114));
    layer2_outputs(2069) <= (layer1_outputs(730)) and not (layer1_outputs(1049));
    layer2_outputs(2070) <= '0';
    layer2_outputs(2071) <= layer1_outputs(720);
    layer2_outputs(2072) <= not((layer1_outputs(1892)) and (layer1_outputs(1449)));
    layer2_outputs(2073) <= not(layer1_outputs(345));
    layer2_outputs(2074) <= (layer1_outputs(1994)) and not (layer1_outputs(2282));
    layer2_outputs(2075) <= '1';
    layer2_outputs(2076) <= (layer1_outputs(58)) and not (layer1_outputs(1045));
    layer2_outputs(2077) <= '0';
    layer2_outputs(2078) <= layer1_outputs(1263);
    layer2_outputs(2079) <= not(layer1_outputs(988)) or (layer1_outputs(1429));
    layer2_outputs(2080) <= not((layer1_outputs(2553)) or (layer1_outputs(1648)));
    layer2_outputs(2081) <= (layer1_outputs(407)) and not (layer1_outputs(959));
    layer2_outputs(2082) <= (layer1_outputs(1313)) and not (layer1_outputs(819));
    layer2_outputs(2083) <= '1';
    layer2_outputs(2084) <= '0';
    layer2_outputs(2085) <= (layer1_outputs(1159)) and (layer1_outputs(266));
    layer2_outputs(2086) <= (layer1_outputs(2048)) and not (layer1_outputs(1983));
    layer2_outputs(2087) <= not(layer1_outputs(1794)) or (layer1_outputs(2529));
    layer2_outputs(2088) <= not(layer1_outputs(604));
    layer2_outputs(2089) <= '0';
    layer2_outputs(2090) <= (layer1_outputs(708)) and not (layer1_outputs(1128));
    layer2_outputs(2091) <= '0';
    layer2_outputs(2092) <= not((layer1_outputs(2351)) or (layer1_outputs(2548)));
    layer2_outputs(2093) <= not(layer1_outputs(1446)) or (layer1_outputs(746));
    layer2_outputs(2094) <= not(layer1_outputs(862));
    layer2_outputs(2095) <= '0';
    layer2_outputs(2096) <= not(layer1_outputs(1401));
    layer2_outputs(2097) <= (layer1_outputs(2357)) xor (layer1_outputs(2400));
    layer2_outputs(2098) <= not((layer1_outputs(2277)) or (layer1_outputs(1332)));
    layer2_outputs(2099) <= not((layer1_outputs(1602)) and (layer1_outputs(393)));
    layer2_outputs(2100) <= not((layer1_outputs(1773)) and (layer1_outputs(1242)));
    layer2_outputs(2101) <= not((layer1_outputs(1778)) or (layer1_outputs(1188)));
    layer2_outputs(2102) <= not(layer1_outputs(545)) or (layer1_outputs(1361));
    layer2_outputs(2103) <= (layer1_outputs(1214)) and (layer1_outputs(824));
    layer2_outputs(2104) <= not(layer1_outputs(1600));
    layer2_outputs(2105) <= not(layer1_outputs(1222)) or (layer1_outputs(161));
    layer2_outputs(2106) <= (layer1_outputs(2023)) and not (layer1_outputs(1382));
    layer2_outputs(2107) <= not(layer1_outputs(2128)) or (layer1_outputs(857));
    layer2_outputs(2108) <= (layer1_outputs(941)) and (layer1_outputs(1669));
    layer2_outputs(2109) <= not((layer1_outputs(1296)) and (layer1_outputs(1065)));
    layer2_outputs(2110) <= (layer1_outputs(2003)) and (layer1_outputs(1075));
    layer2_outputs(2111) <= not(layer1_outputs(1609)) or (layer1_outputs(1271));
    layer2_outputs(2112) <= '1';
    layer2_outputs(2113) <= '1';
    layer2_outputs(2114) <= (layer1_outputs(2541)) and (layer1_outputs(1727));
    layer2_outputs(2115) <= not(layer1_outputs(2414)) or (layer1_outputs(328));
    layer2_outputs(2116) <= layer1_outputs(665);
    layer2_outputs(2117) <= (layer1_outputs(1580)) xor (layer1_outputs(860));
    layer2_outputs(2118) <= not(layer1_outputs(1903));
    layer2_outputs(2119) <= (layer1_outputs(1390)) and (layer1_outputs(1399));
    layer2_outputs(2120) <= (layer1_outputs(996)) and (layer1_outputs(712));
    layer2_outputs(2121) <= (layer1_outputs(1136)) or (layer1_outputs(681));
    layer2_outputs(2122) <= '0';
    layer2_outputs(2123) <= not(layer1_outputs(1406)) or (layer1_outputs(1218));
    layer2_outputs(2124) <= '0';
    layer2_outputs(2125) <= not(layer1_outputs(1988)) or (layer1_outputs(1704));
    layer2_outputs(2126) <= (layer1_outputs(2448)) and (layer1_outputs(2247));
    layer2_outputs(2127) <= not(layer1_outputs(240));
    layer2_outputs(2128) <= '1';
    layer2_outputs(2129) <= not((layer1_outputs(2517)) and (layer1_outputs(559)));
    layer2_outputs(2130) <= not(layer1_outputs(241)) or (layer1_outputs(469));
    layer2_outputs(2131) <= not(layer1_outputs(1720));
    layer2_outputs(2132) <= not(layer1_outputs(2505));
    layer2_outputs(2133) <= (layer1_outputs(1328)) and not (layer1_outputs(1023));
    layer2_outputs(2134) <= (layer1_outputs(2201)) or (layer1_outputs(1054));
    layer2_outputs(2135) <= '0';
    layer2_outputs(2136) <= (layer1_outputs(1052)) or (layer1_outputs(2472));
    layer2_outputs(2137) <= (layer1_outputs(1149)) or (layer1_outputs(355));
    layer2_outputs(2138) <= not(layer1_outputs(96));
    layer2_outputs(2139) <= not(layer1_outputs(1225));
    layer2_outputs(2140) <= (layer1_outputs(768)) and not (layer1_outputs(1902));
    layer2_outputs(2141) <= (layer1_outputs(173)) or (layer1_outputs(2160));
    layer2_outputs(2142) <= '1';
    layer2_outputs(2143) <= not(layer1_outputs(227)) or (layer1_outputs(2478));
    layer2_outputs(2144) <= (layer1_outputs(1608)) and not (layer1_outputs(1830));
    layer2_outputs(2145) <= layer1_outputs(1653);
    layer2_outputs(2146) <= '1';
    layer2_outputs(2147) <= (layer1_outputs(1581)) and not (layer1_outputs(688));
    layer2_outputs(2148) <= (layer1_outputs(2331)) and not (layer1_outputs(1330));
    layer2_outputs(2149) <= not(layer1_outputs(1247)) or (layer1_outputs(718));
    layer2_outputs(2150) <= layer1_outputs(925);
    layer2_outputs(2151) <= layer1_outputs(1039);
    layer2_outputs(2152) <= (layer1_outputs(2559)) and not (layer1_outputs(2277));
    layer2_outputs(2153) <= not(layer1_outputs(815)) or (layer1_outputs(818));
    layer2_outputs(2154) <= '1';
    layer2_outputs(2155) <= not((layer1_outputs(1835)) and (layer1_outputs(1314)));
    layer2_outputs(2156) <= (layer1_outputs(1643)) and not (layer1_outputs(1930));
    layer2_outputs(2157) <= not(layer1_outputs(1969));
    layer2_outputs(2158) <= (layer1_outputs(1760)) and (layer1_outputs(2299));
    layer2_outputs(2159) <= layer1_outputs(808);
    layer2_outputs(2160) <= (layer1_outputs(1238)) xor (layer1_outputs(1917));
    layer2_outputs(2161) <= '0';
    layer2_outputs(2162) <= (layer1_outputs(1856)) and not (layer1_outputs(1358));
    layer2_outputs(2163) <= layer1_outputs(1208);
    layer2_outputs(2164) <= '0';
    layer2_outputs(2165) <= (layer1_outputs(1014)) and (layer1_outputs(400));
    layer2_outputs(2166) <= layer1_outputs(1567);
    layer2_outputs(2167) <= layer1_outputs(2433);
    layer2_outputs(2168) <= '0';
    layer2_outputs(2169) <= '0';
    layer2_outputs(2170) <= (layer1_outputs(722)) and not (layer1_outputs(532));
    layer2_outputs(2171) <= not(layer1_outputs(1834)) or (layer1_outputs(811));
    layer2_outputs(2172) <= layer1_outputs(613);
    layer2_outputs(2173) <= not((layer1_outputs(760)) or (layer1_outputs(1882)));
    layer2_outputs(2174) <= (layer1_outputs(824)) and not (layer1_outputs(23));
    layer2_outputs(2175) <= layer1_outputs(2114);
    layer2_outputs(2176) <= (layer1_outputs(1678)) or (layer1_outputs(378));
    layer2_outputs(2177) <= not((layer1_outputs(1266)) or (layer1_outputs(177)));
    layer2_outputs(2178) <= not(layer1_outputs(1028)) or (layer1_outputs(1451));
    layer2_outputs(2179) <= '1';
    layer2_outputs(2180) <= not(layer1_outputs(31));
    layer2_outputs(2181) <= not(layer1_outputs(42));
    layer2_outputs(2182) <= (layer1_outputs(2555)) and not (layer1_outputs(226));
    layer2_outputs(2183) <= '0';
    layer2_outputs(2184) <= '0';
    layer2_outputs(2185) <= not((layer1_outputs(1828)) or (layer1_outputs(1581)));
    layer2_outputs(2186) <= layer1_outputs(353);
    layer2_outputs(2187) <= (layer1_outputs(479)) and not (layer1_outputs(2272));
    layer2_outputs(2188) <= '1';
    layer2_outputs(2189) <= '1';
    layer2_outputs(2190) <= '1';
    layer2_outputs(2191) <= (layer1_outputs(2135)) or (layer1_outputs(1757));
    layer2_outputs(2192) <= layer1_outputs(1901);
    layer2_outputs(2193) <= layer1_outputs(1684);
    layer2_outputs(2194) <= (layer1_outputs(1305)) and (layer1_outputs(2315));
    layer2_outputs(2195) <= layer1_outputs(676);
    layer2_outputs(2196) <= not(layer1_outputs(2190)) or (layer1_outputs(2382));
    layer2_outputs(2197) <= not(layer1_outputs(260));
    layer2_outputs(2198) <= (layer1_outputs(1052)) and (layer1_outputs(1468));
    layer2_outputs(2199) <= layer1_outputs(2468);
    layer2_outputs(2200) <= not(layer1_outputs(633)) or (layer1_outputs(1955));
    layer2_outputs(2201) <= not(layer1_outputs(1235));
    layer2_outputs(2202) <= not(layer1_outputs(736)) or (layer1_outputs(900));
    layer2_outputs(2203) <= not(layer1_outputs(2523)) or (layer1_outputs(2407));
    layer2_outputs(2204) <= (layer1_outputs(804)) and not (layer1_outputs(2325));
    layer2_outputs(2205) <= (layer1_outputs(900)) and not (layer1_outputs(1535));
    layer2_outputs(2206) <= layer1_outputs(8);
    layer2_outputs(2207) <= (layer1_outputs(1124)) and not (layer1_outputs(1566));
    layer2_outputs(2208) <= not(layer1_outputs(2018)) or (layer1_outputs(441));
    layer2_outputs(2209) <= layer1_outputs(1510);
    layer2_outputs(2210) <= not(layer1_outputs(1988));
    layer2_outputs(2211) <= '0';
    layer2_outputs(2212) <= not((layer1_outputs(81)) and (layer1_outputs(2064)));
    layer2_outputs(2213) <= (layer1_outputs(1628)) and not (layer1_outputs(1046));
    layer2_outputs(2214) <= '1';
    layer2_outputs(2215) <= not((layer1_outputs(504)) and (layer1_outputs(1367)));
    layer2_outputs(2216) <= layer1_outputs(1114);
    layer2_outputs(2217) <= not((layer1_outputs(2216)) or (layer1_outputs(2276)));
    layer2_outputs(2218) <= not(layer1_outputs(405));
    layer2_outputs(2219) <= not(layer1_outputs(764)) or (layer1_outputs(2304));
    layer2_outputs(2220) <= not(layer1_outputs(1299));
    layer2_outputs(2221) <= (layer1_outputs(2184)) or (layer1_outputs(1142));
    layer2_outputs(2222) <= not(layer1_outputs(2214)) or (layer1_outputs(2015));
    layer2_outputs(2223) <= '1';
    layer2_outputs(2224) <= '1';
    layer2_outputs(2225) <= layer1_outputs(1541);
    layer2_outputs(2226) <= (layer1_outputs(2191)) and (layer1_outputs(147));
    layer2_outputs(2227) <= layer1_outputs(361);
    layer2_outputs(2228) <= not(layer1_outputs(2030));
    layer2_outputs(2229) <= not((layer1_outputs(662)) or (layer1_outputs(2176)));
    layer2_outputs(2230) <= (layer1_outputs(268)) or (layer1_outputs(1470));
    layer2_outputs(2231) <= not(layer1_outputs(33));
    layer2_outputs(2232) <= not(layer1_outputs(744));
    layer2_outputs(2233) <= '1';
    layer2_outputs(2234) <= (layer1_outputs(2097)) and not (layer1_outputs(2456));
    layer2_outputs(2235) <= (layer1_outputs(1849)) and (layer1_outputs(1738));
    layer2_outputs(2236) <= layer1_outputs(955);
    layer2_outputs(2237) <= '1';
    layer2_outputs(2238) <= (layer1_outputs(2421)) and not (layer1_outputs(44));
    layer2_outputs(2239) <= not(layer1_outputs(2045)) or (layer1_outputs(2484));
    layer2_outputs(2240) <= '1';
    layer2_outputs(2241) <= (layer1_outputs(1212)) and not (layer1_outputs(2285));
    layer2_outputs(2242) <= layer1_outputs(634);
    layer2_outputs(2243) <= not((layer1_outputs(1753)) and (layer1_outputs(1854)));
    layer2_outputs(2244) <= not((layer1_outputs(1702)) and (layer1_outputs(1967)));
    layer2_outputs(2245) <= (layer1_outputs(644)) and not (layer1_outputs(709));
    layer2_outputs(2246) <= '1';
    layer2_outputs(2247) <= not((layer1_outputs(2391)) or (layer1_outputs(2317)));
    layer2_outputs(2248) <= layer1_outputs(355);
    layer2_outputs(2249) <= (layer1_outputs(668)) or (layer1_outputs(1721));
    layer2_outputs(2250) <= '0';
    layer2_outputs(2251) <= not((layer1_outputs(2085)) or (layer1_outputs(1146)));
    layer2_outputs(2252) <= layer1_outputs(1484);
    layer2_outputs(2253) <= not((layer1_outputs(718)) or (layer1_outputs(59)));
    layer2_outputs(2254) <= not(layer1_outputs(638));
    layer2_outputs(2255) <= layer1_outputs(1230);
    layer2_outputs(2256) <= '1';
    layer2_outputs(2257) <= '0';
    layer2_outputs(2258) <= not(layer1_outputs(40));
    layer2_outputs(2259) <= (layer1_outputs(2434)) and (layer1_outputs(2387));
    layer2_outputs(2260) <= not(layer1_outputs(20)) or (layer1_outputs(462));
    layer2_outputs(2261) <= (layer1_outputs(374)) and not (layer1_outputs(1176));
    layer2_outputs(2262) <= not((layer1_outputs(1412)) and (layer1_outputs(2373)));
    layer2_outputs(2263) <= (layer1_outputs(357)) or (layer1_outputs(1642));
    layer2_outputs(2264) <= (layer1_outputs(1227)) and (layer1_outputs(1383));
    layer2_outputs(2265) <= not((layer1_outputs(310)) and (layer1_outputs(1599)));
    layer2_outputs(2266) <= layer1_outputs(1543);
    layer2_outputs(2267) <= not(layer1_outputs(329)) or (layer1_outputs(869));
    layer2_outputs(2268) <= not((layer1_outputs(1066)) and (layer1_outputs(41)));
    layer2_outputs(2269) <= layer1_outputs(75);
    layer2_outputs(2270) <= not(layer1_outputs(489));
    layer2_outputs(2271) <= (layer1_outputs(2358)) xor (layer1_outputs(1708));
    layer2_outputs(2272) <= not((layer1_outputs(2525)) and (layer1_outputs(1387)));
    layer2_outputs(2273) <= (layer1_outputs(785)) and not (layer1_outputs(306));
    layer2_outputs(2274) <= '0';
    layer2_outputs(2275) <= layer1_outputs(2089);
    layer2_outputs(2276) <= not((layer1_outputs(1243)) or (layer1_outputs(1017)));
    layer2_outputs(2277) <= (layer1_outputs(2283)) and (layer1_outputs(472));
    layer2_outputs(2278) <= not((layer1_outputs(277)) and (layer1_outputs(2111)));
    layer2_outputs(2279) <= '1';
    layer2_outputs(2280) <= (layer1_outputs(43)) and not (layer1_outputs(2490));
    layer2_outputs(2281) <= not(layer1_outputs(793)) or (layer1_outputs(1716));
    layer2_outputs(2282) <= not(layer1_outputs(2008));
    layer2_outputs(2283) <= (layer1_outputs(142)) and not (layer1_outputs(390));
    layer2_outputs(2284) <= not(layer1_outputs(1173));
    layer2_outputs(2285) <= not((layer1_outputs(807)) or (layer1_outputs(1293)));
    layer2_outputs(2286) <= '1';
    layer2_outputs(2287) <= '1';
    layer2_outputs(2288) <= '0';
    layer2_outputs(2289) <= (layer1_outputs(1964)) and (layer1_outputs(1016));
    layer2_outputs(2290) <= not(layer1_outputs(1365));
    layer2_outputs(2291) <= '1';
    layer2_outputs(2292) <= not(layer1_outputs(692)) or (layer1_outputs(1517));
    layer2_outputs(2293) <= '1';
    layer2_outputs(2294) <= (layer1_outputs(256)) and not (layer1_outputs(314));
    layer2_outputs(2295) <= not(layer1_outputs(2383));
    layer2_outputs(2296) <= not((layer1_outputs(976)) and (layer1_outputs(2344)));
    layer2_outputs(2297) <= layer1_outputs(1840);
    layer2_outputs(2298) <= '1';
    layer2_outputs(2299) <= not(layer1_outputs(735)) or (layer1_outputs(1190));
    layer2_outputs(2300) <= not((layer1_outputs(2161)) and (layer1_outputs(1978)));
    layer2_outputs(2301) <= (layer1_outputs(273)) and not (layer1_outputs(1516));
    layer2_outputs(2302) <= layer1_outputs(13);
    layer2_outputs(2303) <= (layer1_outputs(221)) and (layer1_outputs(655));
    layer2_outputs(2304) <= layer1_outputs(977);
    layer2_outputs(2305) <= layer1_outputs(2066);
    layer2_outputs(2306) <= not((layer1_outputs(161)) or (layer1_outputs(1745)));
    layer2_outputs(2307) <= not(layer1_outputs(2557));
    layer2_outputs(2308) <= layer1_outputs(512);
    layer2_outputs(2309) <= (layer1_outputs(124)) and not (layer1_outputs(2054));
    layer2_outputs(2310) <= layer1_outputs(1797);
    layer2_outputs(2311) <= not(layer1_outputs(695));
    layer2_outputs(2312) <= not(layer1_outputs(2210)) or (layer1_outputs(1112));
    layer2_outputs(2313) <= (layer1_outputs(2172)) and not (layer1_outputs(1694));
    layer2_outputs(2314) <= (layer1_outputs(995)) or (layer1_outputs(841));
    layer2_outputs(2315) <= not(layer1_outputs(953));
    layer2_outputs(2316) <= not(layer1_outputs(382)) or (layer1_outputs(198));
    layer2_outputs(2317) <= layer1_outputs(797);
    layer2_outputs(2318) <= '0';
    layer2_outputs(2319) <= not(layer1_outputs(2463)) or (layer1_outputs(1942));
    layer2_outputs(2320) <= '0';
    layer2_outputs(2321) <= '1';
    layer2_outputs(2322) <= not(layer1_outputs(185)) or (layer1_outputs(592));
    layer2_outputs(2323) <= '1';
    layer2_outputs(2324) <= (layer1_outputs(2221)) and not (layer1_outputs(140));
    layer2_outputs(2325) <= not(layer1_outputs(1998));
    layer2_outputs(2326) <= not((layer1_outputs(1205)) and (layer1_outputs(175)));
    layer2_outputs(2327) <= '0';
    layer2_outputs(2328) <= (layer1_outputs(2282)) and not (layer1_outputs(1870));
    layer2_outputs(2329) <= not(layer1_outputs(2417));
    layer2_outputs(2330) <= (layer1_outputs(2079)) and not (layer1_outputs(566));
    layer2_outputs(2331) <= (layer1_outputs(596)) or (layer1_outputs(1041));
    layer2_outputs(2332) <= '1';
    layer2_outputs(2333) <= not(layer1_outputs(1318));
    layer2_outputs(2334) <= not(layer1_outputs(1704)) or (layer1_outputs(1852));
    layer2_outputs(2335) <= (layer1_outputs(1841)) and not (layer1_outputs(2184));
    layer2_outputs(2336) <= not(layer1_outputs(2306)) or (layer1_outputs(832));
    layer2_outputs(2337) <= (layer1_outputs(34)) and not (layer1_outputs(766));
    layer2_outputs(2338) <= not(layer1_outputs(515));
    layer2_outputs(2339) <= '0';
    layer2_outputs(2340) <= '1';
    layer2_outputs(2341) <= not(layer1_outputs(2469)) or (layer1_outputs(564));
    layer2_outputs(2342) <= layer1_outputs(897);
    layer2_outputs(2343) <= not(layer1_outputs(534));
    layer2_outputs(2344) <= '1';
    layer2_outputs(2345) <= not(layer1_outputs(32)) or (layer1_outputs(286));
    layer2_outputs(2346) <= not(layer1_outputs(147)) or (layer1_outputs(1638));
    layer2_outputs(2347) <= not(layer1_outputs(1205));
    layer2_outputs(2348) <= layer1_outputs(363);
    layer2_outputs(2349) <= (layer1_outputs(1414)) or (layer1_outputs(1847));
    layer2_outputs(2350) <= not(layer1_outputs(514)) or (layer1_outputs(1495));
    layer2_outputs(2351) <= (layer1_outputs(1410)) and not (layer1_outputs(1776));
    layer2_outputs(2352) <= '1';
    layer2_outputs(2353) <= not(layer1_outputs(2299)) or (layer1_outputs(1303));
    layer2_outputs(2354) <= not(layer1_outputs(910));
    layer2_outputs(2355) <= (layer1_outputs(1804)) and not (layer1_outputs(2367));
    layer2_outputs(2356) <= '1';
    layer2_outputs(2357) <= (layer1_outputs(1240)) and (layer1_outputs(495));
    layer2_outputs(2358) <= (layer1_outputs(658)) and not (layer1_outputs(1241));
    layer2_outputs(2359) <= not((layer1_outputs(2440)) and (layer1_outputs(213)));
    layer2_outputs(2360) <= (layer1_outputs(1076)) and not (layer1_outputs(1042));
    layer2_outputs(2361) <= not(layer1_outputs(1116));
    layer2_outputs(2362) <= not(layer1_outputs(966)) or (layer1_outputs(671));
    layer2_outputs(2363) <= '1';
    layer2_outputs(2364) <= layer1_outputs(1626);
    layer2_outputs(2365) <= (layer1_outputs(2208)) and not (layer1_outputs(950));
    layer2_outputs(2366) <= not(layer1_outputs(1274));
    layer2_outputs(2367) <= '0';
    layer2_outputs(2368) <= '0';
    layer2_outputs(2369) <= not((layer1_outputs(2071)) xor (layer1_outputs(1639)));
    layer2_outputs(2370) <= not((layer1_outputs(207)) or (layer1_outputs(741)));
    layer2_outputs(2371) <= layer1_outputs(825);
    layer2_outputs(2372) <= not(layer1_outputs(997));
    layer2_outputs(2373) <= (layer1_outputs(101)) and not (layer1_outputs(2390));
    layer2_outputs(2374) <= not(layer1_outputs(1304)) or (layer1_outputs(627));
    layer2_outputs(2375) <= '1';
    layer2_outputs(2376) <= '0';
    layer2_outputs(2377) <= (layer1_outputs(2311)) and not (layer1_outputs(1174));
    layer2_outputs(2378) <= not(layer1_outputs(1762));
    layer2_outputs(2379) <= (layer1_outputs(2113)) or (layer1_outputs(1884));
    layer2_outputs(2380) <= not(layer1_outputs(336));
    layer2_outputs(2381) <= '0';
    layer2_outputs(2382) <= not(layer1_outputs(1944)) or (layer1_outputs(1025));
    layer2_outputs(2383) <= layer1_outputs(1679);
    layer2_outputs(2384) <= (layer1_outputs(1189)) and not (layer1_outputs(2095));
    layer2_outputs(2385) <= '1';
    layer2_outputs(2386) <= not(layer1_outputs(1455)) or (layer1_outputs(1090));
    layer2_outputs(2387) <= '0';
    layer2_outputs(2388) <= '1';
    layer2_outputs(2389) <= (layer1_outputs(691)) or (layer1_outputs(2475));
    layer2_outputs(2390) <= not(layer1_outputs(1480));
    layer2_outputs(2391) <= not(layer1_outputs(1888));
    layer2_outputs(2392) <= (layer1_outputs(2212)) and not (layer1_outputs(535));
    layer2_outputs(2393) <= '1';
    layer2_outputs(2394) <= layer1_outputs(1498);
    layer2_outputs(2395) <= layer1_outputs(467);
    layer2_outputs(2396) <= layer1_outputs(1177);
    layer2_outputs(2397) <= not((layer1_outputs(1926)) and (layer1_outputs(1261)));
    layer2_outputs(2398) <= (layer1_outputs(2194)) and not (layer1_outputs(487));
    layer2_outputs(2399) <= '0';
    layer2_outputs(2400) <= (layer1_outputs(476)) or (layer1_outputs(291));
    layer2_outputs(2401) <= '1';
    layer2_outputs(2402) <= (layer1_outputs(1335)) and not (layer1_outputs(461));
    layer2_outputs(2403) <= '0';
    layer2_outputs(2404) <= (layer1_outputs(2511)) or (layer1_outputs(1160));
    layer2_outputs(2405) <= not(layer1_outputs(554));
    layer2_outputs(2406) <= '1';
    layer2_outputs(2407) <= '1';
    layer2_outputs(2408) <= not(layer1_outputs(494));
    layer2_outputs(2409) <= not(layer1_outputs(723));
    layer2_outputs(2410) <= not(layer1_outputs(1693));
    layer2_outputs(2411) <= not(layer1_outputs(2462)) or (layer1_outputs(1106));
    layer2_outputs(2412) <= '0';
    layer2_outputs(2413) <= not(layer1_outputs(2167)) or (layer1_outputs(2362));
    layer2_outputs(2414) <= not((layer1_outputs(2268)) and (layer1_outputs(745)));
    layer2_outputs(2415) <= (layer1_outputs(1953)) and not (layer1_outputs(350));
    layer2_outputs(2416) <= layer1_outputs(1622);
    layer2_outputs(2417) <= not(layer1_outputs(1271));
    layer2_outputs(2418) <= not(layer1_outputs(1657));
    layer2_outputs(2419) <= not((layer1_outputs(913)) and (layer1_outputs(1077)));
    layer2_outputs(2420) <= (layer1_outputs(678)) and (layer1_outputs(762));
    layer2_outputs(2421) <= (layer1_outputs(781)) and not (layer1_outputs(133));
    layer2_outputs(2422) <= '1';
    layer2_outputs(2423) <= not(layer1_outputs(1845)) or (layer1_outputs(1501));
    layer2_outputs(2424) <= not(layer1_outputs(398));
    layer2_outputs(2425) <= layer1_outputs(871);
    layer2_outputs(2426) <= '0';
    layer2_outputs(2427) <= not(layer1_outputs(947)) or (layer1_outputs(308));
    layer2_outputs(2428) <= layer1_outputs(423);
    layer2_outputs(2429) <= (layer1_outputs(1151)) or (layer1_outputs(424));
    layer2_outputs(2430) <= not(layer1_outputs(1001));
    layer2_outputs(2431) <= layer1_outputs(2240);
    layer2_outputs(2432) <= not(layer1_outputs(1379));
    layer2_outputs(2433) <= not(layer1_outputs(631));
    layer2_outputs(2434) <= (layer1_outputs(445)) and not (layer1_outputs(195));
    layer2_outputs(2435) <= (layer1_outputs(550)) and not (layer1_outputs(303));
    layer2_outputs(2436) <= not(layer1_outputs(1634)) or (layer1_outputs(2214));
    layer2_outputs(2437) <= '0';
    layer2_outputs(2438) <= '0';
    layer2_outputs(2439) <= not(layer1_outputs(1928)) or (layer1_outputs(1497));
    layer2_outputs(2440) <= not(layer1_outputs(775));
    layer2_outputs(2441) <= not((layer1_outputs(1974)) or (layer1_outputs(2086)));
    layer2_outputs(2442) <= '1';
    layer2_outputs(2443) <= '1';
    layer2_outputs(2444) <= layer1_outputs(2370);
    layer2_outputs(2445) <= '0';
    layer2_outputs(2446) <= (layer1_outputs(249)) and (layer1_outputs(285));
    layer2_outputs(2447) <= (layer1_outputs(1413)) or (layer1_outputs(1323));
    layer2_outputs(2448) <= not((layer1_outputs(2409)) or (layer1_outputs(679)));
    layer2_outputs(2449) <= '0';
    layer2_outputs(2450) <= (layer1_outputs(1601)) and (layer1_outputs(442));
    layer2_outputs(2451) <= not((layer1_outputs(192)) xor (layer1_outputs(1460)));
    layer2_outputs(2452) <= layer1_outputs(1866);
    layer2_outputs(2453) <= not((layer1_outputs(1044)) or (layer1_outputs(1793)));
    layer2_outputs(2454) <= not((layer1_outputs(1137)) or (layer1_outputs(2535)));
    layer2_outputs(2455) <= not(layer1_outputs(1200));
    layer2_outputs(2456) <= not(layer1_outputs(628));
    layer2_outputs(2457) <= not(layer1_outputs(948)) or (layer1_outputs(1593));
    layer2_outputs(2458) <= not((layer1_outputs(2182)) and (layer1_outputs(2273)));
    layer2_outputs(2459) <= not((layer1_outputs(2089)) and (layer1_outputs(1538)));
    layer2_outputs(2460) <= not((layer1_outputs(794)) or (layer1_outputs(1113)));
    layer2_outputs(2461) <= (layer1_outputs(1868)) and (layer1_outputs(1818));
    layer2_outputs(2462) <= not(layer1_outputs(1952));
    layer2_outputs(2463) <= not((layer1_outputs(2239)) or (layer1_outputs(2302)));
    layer2_outputs(2464) <= not(layer1_outputs(1194)) or (layer1_outputs(2070));
    layer2_outputs(2465) <= (layer1_outputs(478)) or (layer1_outputs(712));
    layer2_outputs(2466) <= not(layer1_outputs(1421)) or (layer1_outputs(1670));
    layer2_outputs(2467) <= (layer1_outputs(2265)) and not (layer1_outputs(1177));
    layer2_outputs(2468) <= not((layer1_outputs(870)) or (layer1_outputs(1571)));
    layer2_outputs(2469) <= (layer1_outputs(1664)) and (layer1_outputs(65));
    layer2_outputs(2470) <= not((layer1_outputs(1267)) or (layer1_outputs(1072)));
    layer2_outputs(2471) <= not(layer1_outputs(1647));
    layer2_outputs(2472) <= layer1_outputs(1031);
    layer2_outputs(2473) <= not(layer1_outputs(2452)) or (layer1_outputs(2129));
    layer2_outputs(2474) <= (layer1_outputs(1353)) or (layer1_outputs(1292));
    layer2_outputs(2475) <= '1';
    layer2_outputs(2476) <= not((layer1_outputs(62)) and (layer1_outputs(2350)));
    layer2_outputs(2477) <= (layer1_outputs(1713)) or (layer1_outputs(919));
    layer2_outputs(2478) <= not(layer1_outputs(42));
    layer2_outputs(2479) <= not((layer1_outputs(2389)) or (layer1_outputs(607)));
    layer2_outputs(2480) <= not(layer1_outputs(1879));
    layer2_outputs(2481) <= not((layer1_outputs(1465)) and (layer1_outputs(491)));
    layer2_outputs(2482) <= '1';
    layer2_outputs(2483) <= not(layer1_outputs(1035)) or (layer1_outputs(458));
    layer2_outputs(2484) <= not(layer1_outputs(85));
    layer2_outputs(2485) <= (layer1_outputs(1661)) and (layer1_outputs(1912));
    layer2_outputs(2486) <= not((layer1_outputs(1621)) and (layer1_outputs(338)));
    layer2_outputs(2487) <= not((layer1_outputs(1564)) and (layer1_outputs(2034)));
    layer2_outputs(2488) <= '1';
    layer2_outputs(2489) <= not(layer1_outputs(439)) or (layer1_outputs(2510));
    layer2_outputs(2490) <= not(layer1_outputs(1881));
    layer2_outputs(2491) <= not(layer1_outputs(163));
    layer2_outputs(2492) <= '1';
    layer2_outputs(2493) <= (layer1_outputs(1453)) or (layer1_outputs(1579));
    layer2_outputs(2494) <= (layer1_outputs(2041)) and not (layer1_outputs(682));
    layer2_outputs(2495) <= '0';
    layer2_outputs(2496) <= not(layer1_outputs(2364));
    layer2_outputs(2497) <= layer1_outputs(579);
    layer2_outputs(2498) <= not(layer1_outputs(294)) or (layer1_outputs(2098));
    layer2_outputs(2499) <= '0';
    layer2_outputs(2500) <= (layer1_outputs(1094)) and (layer1_outputs(1474));
    layer2_outputs(2501) <= layer1_outputs(1826);
    layer2_outputs(2502) <= '1';
    layer2_outputs(2503) <= not((layer1_outputs(2326)) and (layer1_outputs(230)));
    layer2_outputs(2504) <= not(layer1_outputs(1859)) or (layer1_outputs(1795));
    layer2_outputs(2505) <= layer1_outputs(2193);
    layer2_outputs(2506) <= (layer1_outputs(1347)) and not (layer1_outputs(2352));
    layer2_outputs(2507) <= (layer1_outputs(1401)) and not (layer1_outputs(1913));
    layer2_outputs(2508) <= (layer1_outputs(1254)) and not (layer1_outputs(468));
    layer2_outputs(2509) <= not(layer1_outputs(303));
    layer2_outputs(2510) <= '0';
    layer2_outputs(2511) <= '0';
    layer2_outputs(2512) <= '0';
    layer2_outputs(2513) <= not(layer1_outputs(743)) or (layer1_outputs(2543));
    layer2_outputs(2514) <= '0';
    layer2_outputs(2515) <= (layer1_outputs(1536)) or (layer1_outputs(1331));
    layer2_outputs(2516) <= not(layer1_outputs(536)) or (layer1_outputs(1087));
    layer2_outputs(2517) <= not((layer1_outputs(2243)) and (layer1_outputs(1454)));
    layer2_outputs(2518) <= not(layer1_outputs(2255));
    layer2_outputs(2519) <= '0';
    layer2_outputs(2520) <= '1';
    layer2_outputs(2521) <= not(layer1_outputs(2403)) or (layer1_outputs(2492));
    layer2_outputs(2522) <= not(layer1_outputs(853));
    layer2_outputs(2523) <= not((layer1_outputs(1403)) or (layer1_outputs(2057)));
    layer2_outputs(2524) <= not(layer1_outputs(275));
    layer2_outputs(2525) <= (layer1_outputs(2137)) and not (layer1_outputs(1402));
    layer2_outputs(2526) <= not((layer1_outputs(446)) xor (layer1_outputs(1048)));
    layer2_outputs(2527) <= '1';
    layer2_outputs(2528) <= (layer1_outputs(2264)) or (layer1_outputs(466));
    layer2_outputs(2529) <= not((layer1_outputs(1835)) or (layer1_outputs(2075)));
    layer2_outputs(2530) <= not(layer1_outputs(1936));
    layer2_outputs(2531) <= layer1_outputs(2128);
    layer2_outputs(2532) <= '1';
    layer2_outputs(2533) <= (layer1_outputs(274)) and not (layer1_outputs(1242));
    layer2_outputs(2534) <= layer1_outputs(1706);
    layer2_outputs(2535) <= (layer1_outputs(30)) and not (layer1_outputs(1006));
    layer2_outputs(2536) <= '1';
    layer2_outputs(2537) <= (layer1_outputs(1287)) and not (layer1_outputs(558));
    layer2_outputs(2538) <= (layer1_outputs(2094)) and not (layer1_outputs(2498));
    layer2_outputs(2539) <= layer1_outputs(2103);
    layer2_outputs(2540) <= not(layer1_outputs(2063));
    layer2_outputs(2541) <= (layer1_outputs(1447)) and (layer1_outputs(1718));
    layer2_outputs(2542) <= layer1_outputs(529);
    layer2_outputs(2543) <= layer1_outputs(2099);
    layer2_outputs(2544) <= not((layer1_outputs(1726)) or (layer1_outputs(1995)));
    layer2_outputs(2545) <= not((layer1_outputs(563)) and (layer1_outputs(539)));
    layer2_outputs(2546) <= '0';
    layer2_outputs(2547) <= (layer1_outputs(740)) and not (layer1_outputs(1916));
    layer2_outputs(2548) <= not(layer1_outputs(248));
    layer2_outputs(2549) <= not(layer1_outputs(1865)) or (layer1_outputs(2196));
    layer2_outputs(2550) <= '1';
    layer2_outputs(2551) <= (layer1_outputs(866)) and not (layer1_outputs(1522));
    layer2_outputs(2552) <= not(layer1_outputs(2495));
    layer2_outputs(2553) <= (layer1_outputs(2116)) or (layer1_outputs(1654));
    layer2_outputs(2554) <= not(layer1_outputs(1511));
    layer2_outputs(2555) <= layer1_outputs(1972);
    layer2_outputs(2556) <= (layer1_outputs(1407)) and not (layer1_outputs(2375));
    layer2_outputs(2557) <= not((layer1_outputs(1498)) and (layer1_outputs(2356)));
    layer2_outputs(2558) <= not((layer1_outputs(1450)) xor (layer1_outputs(1910)));
    layer2_outputs(2559) <= (layer1_outputs(1816)) and (layer1_outputs(351));
    layer3_outputs(0) <= not((layer2_outputs(2432)) or (layer2_outputs(311)));
    layer3_outputs(1) <= not(layer2_outputs(1026)) or (layer2_outputs(756));
    layer3_outputs(2) <= '0';
    layer3_outputs(3) <= not(layer2_outputs(2322)) or (layer2_outputs(103));
    layer3_outputs(4) <= layer2_outputs(103);
    layer3_outputs(5) <= not((layer2_outputs(956)) and (layer2_outputs(312)));
    layer3_outputs(6) <= not(layer2_outputs(1647)) or (layer2_outputs(1642));
    layer3_outputs(7) <= not((layer2_outputs(761)) and (layer2_outputs(996)));
    layer3_outputs(8) <= not(layer2_outputs(269)) or (layer2_outputs(2401));
    layer3_outputs(9) <= not((layer2_outputs(687)) or (layer2_outputs(805)));
    layer3_outputs(10) <= '1';
    layer3_outputs(11) <= not((layer2_outputs(2196)) and (layer2_outputs(2003)));
    layer3_outputs(12) <= '1';
    layer3_outputs(13) <= '1';
    layer3_outputs(14) <= layer2_outputs(670);
    layer3_outputs(15) <= not((layer2_outputs(2480)) and (layer2_outputs(1555)));
    layer3_outputs(16) <= '1';
    layer3_outputs(17) <= (layer2_outputs(682)) and not (layer2_outputs(2104));
    layer3_outputs(18) <= '1';
    layer3_outputs(19) <= not((layer2_outputs(137)) and (layer2_outputs(675)));
    layer3_outputs(20) <= '0';
    layer3_outputs(21) <= (layer2_outputs(1331)) and not (layer2_outputs(326));
    layer3_outputs(22) <= '1';
    layer3_outputs(23) <= not(layer2_outputs(1042)) or (layer2_outputs(834));
    layer3_outputs(24) <= '1';
    layer3_outputs(25) <= not(layer2_outputs(1153));
    layer3_outputs(26) <= layer2_outputs(869);
    layer3_outputs(27) <= not(layer2_outputs(1160));
    layer3_outputs(28) <= not((layer2_outputs(1206)) and (layer2_outputs(1499)));
    layer3_outputs(29) <= layer2_outputs(2165);
    layer3_outputs(30) <= not((layer2_outputs(759)) and (layer2_outputs(471)));
    layer3_outputs(31) <= not((layer2_outputs(91)) xor (layer2_outputs(312)));
    layer3_outputs(32) <= layer2_outputs(137);
    layer3_outputs(33) <= layer2_outputs(2084);
    layer3_outputs(34) <= '0';
    layer3_outputs(35) <= (layer2_outputs(1241)) and not (layer2_outputs(1737));
    layer3_outputs(36) <= layer2_outputs(864);
    layer3_outputs(37) <= (layer2_outputs(1487)) and (layer2_outputs(2126));
    layer3_outputs(38) <= (layer2_outputs(947)) and (layer2_outputs(857));
    layer3_outputs(39) <= '0';
    layer3_outputs(40) <= not(layer2_outputs(919)) or (layer2_outputs(34));
    layer3_outputs(41) <= (layer2_outputs(1941)) and not (layer2_outputs(1389));
    layer3_outputs(42) <= not(layer2_outputs(2374)) or (layer2_outputs(964));
    layer3_outputs(43) <= not((layer2_outputs(1422)) and (layer2_outputs(300)));
    layer3_outputs(44) <= not((layer2_outputs(1883)) and (layer2_outputs(149)));
    layer3_outputs(45) <= '0';
    layer3_outputs(46) <= (layer2_outputs(2373)) or (layer2_outputs(667));
    layer3_outputs(47) <= (layer2_outputs(303)) or (layer2_outputs(206));
    layer3_outputs(48) <= (layer2_outputs(73)) and not (layer2_outputs(748));
    layer3_outputs(49) <= not(layer2_outputs(287)) or (layer2_outputs(2412));
    layer3_outputs(50) <= layer2_outputs(1281);
    layer3_outputs(51) <= layer2_outputs(2215);
    layer3_outputs(52) <= (layer2_outputs(882)) and (layer2_outputs(1733));
    layer3_outputs(53) <= (layer2_outputs(1307)) and not (layer2_outputs(653));
    layer3_outputs(54) <= not((layer2_outputs(1699)) or (layer2_outputs(2533)));
    layer3_outputs(55) <= not((layer2_outputs(1132)) and (layer2_outputs(365)));
    layer3_outputs(56) <= (layer2_outputs(1905)) and (layer2_outputs(796));
    layer3_outputs(57) <= not(layer2_outputs(1339)) or (layer2_outputs(1697));
    layer3_outputs(58) <= not(layer2_outputs(1489)) or (layer2_outputs(814));
    layer3_outputs(59) <= (layer2_outputs(2312)) and not (layer2_outputs(82));
    layer3_outputs(60) <= not((layer2_outputs(1298)) and (layer2_outputs(548)));
    layer3_outputs(61) <= layer2_outputs(180);
    layer3_outputs(62) <= '1';
    layer3_outputs(63) <= '1';
    layer3_outputs(64) <= not(layer2_outputs(513));
    layer3_outputs(65) <= '1';
    layer3_outputs(66) <= not(layer2_outputs(2270)) or (layer2_outputs(883));
    layer3_outputs(67) <= '1';
    layer3_outputs(68) <= not(layer2_outputs(2450));
    layer3_outputs(69) <= not(layer2_outputs(1152));
    layer3_outputs(70) <= not((layer2_outputs(1153)) or (layer2_outputs(770)));
    layer3_outputs(71) <= not((layer2_outputs(577)) or (layer2_outputs(2394)));
    layer3_outputs(72) <= not((layer2_outputs(615)) or (layer2_outputs(679)));
    layer3_outputs(73) <= not(layer2_outputs(1808)) or (layer2_outputs(1995));
    layer3_outputs(74) <= layer2_outputs(1254);
    layer3_outputs(75) <= (layer2_outputs(1795)) or (layer2_outputs(1182));
    layer3_outputs(76) <= '0';
    layer3_outputs(77) <= not(layer2_outputs(401));
    layer3_outputs(78) <= (layer2_outputs(1934)) or (layer2_outputs(2173));
    layer3_outputs(79) <= (layer2_outputs(774)) and (layer2_outputs(1224));
    layer3_outputs(80) <= '0';
    layer3_outputs(81) <= '1';
    layer3_outputs(82) <= not((layer2_outputs(1988)) and (layer2_outputs(2025)));
    layer3_outputs(83) <= (layer2_outputs(2521)) or (layer2_outputs(1109));
    layer3_outputs(84) <= layer2_outputs(2439);
    layer3_outputs(85) <= (layer2_outputs(1637)) or (layer2_outputs(655));
    layer3_outputs(86) <= (layer2_outputs(592)) and (layer2_outputs(1213));
    layer3_outputs(87) <= layer2_outputs(2372);
    layer3_outputs(88) <= not(layer2_outputs(2073));
    layer3_outputs(89) <= (layer2_outputs(843)) and not (layer2_outputs(2462));
    layer3_outputs(90) <= layer2_outputs(1549);
    layer3_outputs(91) <= '1';
    layer3_outputs(92) <= not(layer2_outputs(1442)) or (layer2_outputs(1666));
    layer3_outputs(93) <= not(layer2_outputs(386));
    layer3_outputs(94) <= (layer2_outputs(1165)) and not (layer2_outputs(1768));
    layer3_outputs(95) <= (layer2_outputs(2235)) xor (layer2_outputs(899));
    layer3_outputs(96) <= layer2_outputs(2156);
    layer3_outputs(97) <= layer2_outputs(2559);
    layer3_outputs(98) <= not(layer2_outputs(1859));
    layer3_outputs(99) <= '1';
    layer3_outputs(100) <= not(layer2_outputs(1742)) or (layer2_outputs(1904));
    layer3_outputs(101) <= '1';
    layer3_outputs(102) <= layer2_outputs(2486);
    layer3_outputs(103) <= not(layer2_outputs(1270));
    layer3_outputs(104) <= (layer2_outputs(4)) or (layer2_outputs(1827));
    layer3_outputs(105) <= (layer2_outputs(2362)) and (layer2_outputs(2075));
    layer3_outputs(106) <= not(layer2_outputs(2183)) or (layer2_outputs(1167));
    layer3_outputs(107) <= '1';
    layer3_outputs(108) <= not((layer2_outputs(1357)) and (layer2_outputs(508)));
    layer3_outputs(109) <= not(layer2_outputs(1265)) or (layer2_outputs(528));
    layer3_outputs(110) <= (layer2_outputs(555)) and not (layer2_outputs(2555));
    layer3_outputs(111) <= not((layer2_outputs(2219)) or (layer2_outputs(2495)));
    layer3_outputs(112) <= layer2_outputs(2063);
    layer3_outputs(113) <= not(layer2_outputs(504)) or (layer2_outputs(1463));
    layer3_outputs(114) <= not(layer2_outputs(1077));
    layer3_outputs(115) <= not((layer2_outputs(1958)) or (layer2_outputs(662)));
    layer3_outputs(116) <= not((layer2_outputs(2435)) and (layer2_outputs(1259)));
    layer3_outputs(117) <= layer2_outputs(1709);
    layer3_outputs(118) <= layer2_outputs(2175);
    layer3_outputs(119) <= not(layer2_outputs(435)) or (layer2_outputs(2133));
    layer3_outputs(120) <= not(layer2_outputs(590)) or (layer2_outputs(1719));
    layer3_outputs(121) <= not(layer2_outputs(672)) or (layer2_outputs(296));
    layer3_outputs(122) <= layer2_outputs(250);
    layer3_outputs(123) <= not(layer2_outputs(650)) or (layer2_outputs(929));
    layer3_outputs(124) <= not(layer2_outputs(1130));
    layer3_outputs(125) <= (layer2_outputs(1822)) or (layer2_outputs(2122));
    layer3_outputs(126) <= not((layer2_outputs(1085)) and (layer2_outputs(1193)));
    layer3_outputs(127) <= not(layer2_outputs(2231));
    layer3_outputs(128) <= (layer2_outputs(1855)) and not (layer2_outputs(525));
    layer3_outputs(129) <= not((layer2_outputs(1816)) or (layer2_outputs(714)));
    layer3_outputs(130) <= '0';
    layer3_outputs(131) <= '0';
    layer3_outputs(132) <= not(layer2_outputs(858)) or (layer2_outputs(1755));
    layer3_outputs(133) <= not(layer2_outputs(1278)) or (layer2_outputs(1743));
    layer3_outputs(134) <= layer2_outputs(2541);
    layer3_outputs(135) <= not(layer2_outputs(115));
    layer3_outputs(136) <= not(layer2_outputs(359));
    layer3_outputs(137) <= '0';
    layer3_outputs(138) <= not(layer2_outputs(1819));
    layer3_outputs(139) <= layer2_outputs(2239);
    layer3_outputs(140) <= not(layer2_outputs(1884));
    layer3_outputs(141) <= layer2_outputs(69);
    layer3_outputs(142) <= '0';
    layer3_outputs(143) <= (layer2_outputs(767)) and not (layer2_outputs(1451));
    layer3_outputs(144) <= layer2_outputs(1909);
    layer3_outputs(145) <= not((layer2_outputs(1266)) or (layer2_outputs(1663)));
    layer3_outputs(146) <= not(layer2_outputs(999)) or (layer2_outputs(2099));
    layer3_outputs(147) <= not((layer2_outputs(860)) or (layer2_outputs(1464)));
    layer3_outputs(148) <= not(layer2_outputs(1695));
    layer3_outputs(149) <= not(layer2_outputs(2192));
    layer3_outputs(150) <= not(layer2_outputs(1229));
    layer3_outputs(151) <= not(layer2_outputs(1556)) or (layer2_outputs(156));
    layer3_outputs(152) <= not((layer2_outputs(2145)) and (layer2_outputs(392)));
    layer3_outputs(153) <= (layer2_outputs(593)) and not (layer2_outputs(602));
    layer3_outputs(154) <= layer2_outputs(679);
    layer3_outputs(155) <= not(layer2_outputs(1991)) or (layer2_outputs(2057));
    layer3_outputs(156) <= not((layer2_outputs(827)) xor (layer2_outputs(1528)));
    layer3_outputs(157) <= not((layer2_outputs(297)) and (layer2_outputs(1047)));
    layer3_outputs(158) <= layer2_outputs(932);
    layer3_outputs(159) <= '0';
    layer3_outputs(160) <= '0';
    layer3_outputs(161) <= '0';
    layer3_outputs(162) <= layer2_outputs(2425);
    layer3_outputs(163) <= (layer2_outputs(38)) or (layer2_outputs(1984));
    layer3_outputs(164) <= (layer2_outputs(2521)) or (layer2_outputs(77));
    layer3_outputs(165) <= not(layer2_outputs(1285));
    layer3_outputs(166) <= '0';
    layer3_outputs(167) <= not(layer2_outputs(2328)) or (layer2_outputs(928));
    layer3_outputs(168) <= (layer2_outputs(1044)) and not (layer2_outputs(2046));
    layer3_outputs(169) <= (layer2_outputs(687)) or (layer2_outputs(954));
    layer3_outputs(170) <= not(layer2_outputs(266)) or (layer2_outputs(1625));
    layer3_outputs(171) <= (layer2_outputs(1769)) or (layer2_outputs(834));
    layer3_outputs(172) <= layer2_outputs(1785);
    layer3_outputs(173) <= layer2_outputs(375);
    layer3_outputs(174) <= not((layer2_outputs(2497)) and (layer2_outputs(667)));
    layer3_outputs(175) <= (layer2_outputs(2496)) and not (layer2_outputs(1337));
    layer3_outputs(176) <= '0';
    layer3_outputs(177) <= not(layer2_outputs(1636));
    layer3_outputs(178) <= layer2_outputs(1727);
    layer3_outputs(179) <= (layer2_outputs(2016)) and not (layer2_outputs(2067));
    layer3_outputs(180) <= not(layer2_outputs(959)) or (layer2_outputs(2459));
    layer3_outputs(181) <= layer2_outputs(2015);
    layer3_outputs(182) <= layer2_outputs(2154);
    layer3_outputs(183) <= layer2_outputs(1332);
    layer3_outputs(184) <= not((layer2_outputs(925)) or (layer2_outputs(810)));
    layer3_outputs(185) <= not(layer2_outputs(727));
    layer3_outputs(186) <= not((layer2_outputs(1497)) or (layer2_outputs(543)));
    layer3_outputs(187) <= not((layer2_outputs(2457)) or (layer2_outputs(2111)));
    layer3_outputs(188) <= (layer2_outputs(985)) and not (layer2_outputs(2281));
    layer3_outputs(189) <= layer2_outputs(1069);
    layer3_outputs(190) <= (layer2_outputs(1490)) or (layer2_outputs(1558));
    layer3_outputs(191) <= not(layer2_outputs(1775)) or (layer2_outputs(1725));
    layer3_outputs(192) <= (layer2_outputs(1613)) or (layer2_outputs(1019));
    layer3_outputs(193) <= (layer2_outputs(280)) or (layer2_outputs(930));
    layer3_outputs(194) <= layer2_outputs(253);
    layer3_outputs(195) <= not((layer2_outputs(850)) or (layer2_outputs(449)));
    layer3_outputs(196) <= (layer2_outputs(276)) and not (layer2_outputs(798));
    layer3_outputs(197) <= not(layer2_outputs(1094)) or (layer2_outputs(32));
    layer3_outputs(198) <= not(layer2_outputs(1873));
    layer3_outputs(199) <= (layer2_outputs(201)) or (layer2_outputs(938));
    layer3_outputs(200) <= '0';
    layer3_outputs(201) <= '0';
    layer3_outputs(202) <= not(layer2_outputs(2468));
    layer3_outputs(203) <= (layer2_outputs(1371)) and (layer2_outputs(98));
    layer3_outputs(204) <= (layer2_outputs(138)) or (layer2_outputs(1258));
    layer3_outputs(205) <= layer2_outputs(221);
    layer3_outputs(206) <= not(layer2_outputs(1358));
    layer3_outputs(207) <= not(layer2_outputs(297));
    layer3_outputs(208) <= not(layer2_outputs(1573));
    layer3_outputs(209) <= not(layer2_outputs(565));
    layer3_outputs(210) <= layer2_outputs(2487);
    layer3_outputs(211) <= layer2_outputs(1229);
    layer3_outputs(212) <= not((layer2_outputs(208)) or (layer2_outputs(373)));
    layer3_outputs(213) <= (layer2_outputs(2217)) xor (layer2_outputs(374));
    layer3_outputs(214) <= layer2_outputs(1318);
    layer3_outputs(215) <= not(layer2_outputs(2533)) or (layer2_outputs(1251));
    layer3_outputs(216) <= '0';
    layer3_outputs(217) <= '1';
    layer3_outputs(218) <= not(layer2_outputs(1587));
    layer3_outputs(219) <= not(layer2_outputs(2145)) or (layer2_outputs(2528));
    layer3_outputs(220) <= not(layer2_outputs(2282));
    layer3_outputs(221) <= '1';
    layer3_outputs(222) <= layer2_outputs(336);
    layer3_outputs(223) <= layer2_outputs(2347);
    layer3_outputs(224) <= not(layer2_outputs(362));
    layer3_outputs(225) <= not((layer2_outputs(745)) and (layer2_outputs(1891)));
    layer3_outputs(226) <= layer2_outputs(1360);
    layer3_outputs(227) <= (layer2_outputs(140)) and not (layer2_outputs(1780));
    layer3_outputs(228) <= (layer2_outputs(2359)) and (layer2_outputs(1936));
    layer3_outputs(229) <= (layer2_outputs(2268)) or (layer2_outputs(1312));
    layer3_outputs(230) <= (layer2_outputs(368)) and not (layer2_outputs(217));
    layer3_outputs(231) <= (layer2_outputs(1960)) and (layer2_outputs(1710));
    layer3_outputs(232) <= '0';
    layer3_outputs(233) <= layer2_outputs(447);
    layer3_outputs(234) <= not(layer2_outputs(946)) or (layer2_outputs(2242));
    layer3_outputs(235) <= (layer2_outputs(830)) and (layer2_outputs(2263));
    layer3_outputs(236) <= not((layer2_outputs(631)) and (layer2_outputs(2239)));
    layer3_outputs(237) <= layer2_outputs(571);
    layer3_outputs(238) <= '0';
    layer3_outputs(239) <= not((layer2_outputs(2004)) and (layer2_outputs(600)));
    layer3_outputs(240) <= layer2_outputs(1389);
    layer3_outputs(241) <= not(layer2_outputs(876)) or (layer2_outputs(590));
    layer3_outputs(242) <= (layer2_outputs(495)) and not (layer2_outputs(683));
    layer3_outputs(243) <= layer2_outputs(1643);
    layer3_outputs(244) <= not(layer2_outputs(2379)) or (layer2_outputs(209));
    layer3_outputs(245) <= (layer2_outputs(1839)) or (layer2_outputs(2523));
    layer3_outputs(246) <= layer2_outputs(1727);
    layer3_outputs(247) <= layer2_outputs(2213);
    layer3_outputs(248) <= not(layer2_outputs(2248));
    layer3_outputs(249) <= not(layer2_outputs(66));
    layer3_outputs(250) <= layer2_outputs(214);
    layer3_outputs(251) <= '0';
    layer3_outputs(252) <= layer2_outputs(1677);
    layer3_outputs(253) <= not(layer2_outputs(702)) or (layer2_outputs(2443));
    layer3_outputs(254) <= '0';
    layer3_outputs(255) <= (layer2_outputs(2106)) and not (layer2_outputs(1415));
    layer3_outputs(256) <= (layer2_outputs(1177)) and not (layer2_outputs(1765));
    layer3_outputs(257) <= (layer2_outputs(1029)) or (layer2_outputs(2222));
    layer3_outputs(258) <= '0';
    layer3_outputs(259) <= '0';
    layer3_outputs(260) <= not(layer2_outputs(2543));
    layer3_outputs(261) <= not(layer2_outputs(395));
    layer3_outputs(262) <= not(layer2_outputs(409)) or (layer2_outputs(1853));
    layer3_outputs(263) <= '0';
    layer3_outputs(264) <= not(layer2_outputs(483));
    layer3_outputs(265) <= not(layer2_outputs(2170));
    layer3_outputs(266) <= not(layer2_outputs(1208)) or (layer2_outputs(2280));
    layer3_outputs(267) <= (layer2_outputs(709)) and not (layer2_outputs(1344));
    layer3_outputs(268) <= '1';
    layer3_outputs(269) <= not((layer2_outputs(1656)) xor (layer2_outputs(820)));
    layer3_outputs(270) <= not((layer2_outputs(2498)) and (layer2_outputs(2489)));
    layer3_outputs(271) <= not((layer2_outputs(2182)) or (layer2_outputs(2208)));
    layer3_outputs(272) <= not(layer2_outputs(1366));
    layer3_outputs(273) <= not((layer2_outputs(356)) and (layer2_outputs(142)));
    layer3_outputs(274) <= (layer2_outputs(2241)) and not (layer2_outputs(230));
    layer3_outputs(275) <= '1';
    layer3_outputs(276) <= '1';
    layer3_outputs(277) <= '1';
    layer3_outputs(278) <= not(layer2_outputs(59));
    layer3_outputs(279) <= not(layer2_outputs(1054));
    layer3_outputs(280) <= (layer2_outputs(906)) or (layer2_outputs(1380));
    layer3_outputs(281) <= '0';
    layer3_outputs(282) <= not(layer2_outputs(2317));
    layer3_outputs(283) <= not(layer2_outputs(1123));
    layer3_outputs(284) <= layer2_outputs(281);
    layer3_outputs(285) <= not(layer2_outputs(1410)) or (layer2_outputs(1817));
    layer3_outputs(286) <= layer2_outputs(703);
    layer3_outputs(287) <= not(layer2_outputs(2131));
    layer3_outputs(288) <= (layer2_outputs(2261)) and not (layer2_outputs(2291));
    layer3_outputs(289) <= '0';
    layer3_outputs(290) <= layer2_outputs(225);
    layer3_outputs(291) <= layer2_outputs(389);
    layer3_outputs(292) <= (layer2_outputs(2429)) and (layer2_outputs(1096));
    layer3_outputs(293) <= (layer2_outputs(51)) xor (layer2_outputs(712));
    layer3_outputs(294) <= layer2_outputs(1592);
    layer3_outputs(295) <= '1';
    layer3_outputs(296) <= not(layer2_outputs(750)) or (layer2_outputs(584));
    layer3_outputs(297) <= '1';
    layer3_outputs(298) <= not((layer2_outputs(2264)) and (layer2_outputs(1542)));
    layer3_outputs(299) <= not(layer2_outputs(1886));
    layer3_outputs(300) <= not(layer2_outputs(802)) or (layer2_outputs(370));
    layer3_outputs(301) <= layer2_outputs(913);
    layer3_outputs(302) <= not(layer2_outputs(660)) or (layer2_outputs(2365));
    layer3_outputs(303) <= not(layer2_outputs(2386));
    layer3_outputs(304) <= layer2_outputs(2);
    layer3_outputs(305) <= not((layer2_outputs(1474)) and (layer2_outputs(2183)));
    layer3_outputs(306) <= (layer2_outputs(638)) and not (layer2_outputs(1010));
    layer3_outputs(307) <= (layer2_outputs(1575)) and not (layer2_outputs(426));
    layer3_outputs(308) <= layer2_outputs(1181);
    layer3_outputs(309) <= (layer2_outputs(2556)) and not (layer2_outputs(2166));
    layer3_outputs(310) <= (layer2_outputs(511)) and not (layer2_outputs(634));
    layer3_outputs(311) <= (layer2_outputs(21)) and (layer2_outputs(1206));
    layer3_outputs(312) <= not(layer2_outputs(236));
    layer3_outputs(313) <= not(layer2_outputs(1663));
    layer3_outputs(314) <= not((layer2_outputs(1712)) and (layer2_outputs(630)));
    layer3_outputs(315) <= (layer2_outputs(2117)) or (layer2_outputs(346));
    layer3_outputs(316) <= (layer2_outputs(495)) and not (layer2_outputs(1135));
    layer3_outputs(317) <= '0';
    layer3_outputs(318) <= (layer2_outputs(1626)) and not (layer2_outputs(1953));
    layer3_outputs(319) <= not(layer2_outputs(1945)) or (layer2_outputs(2308));
    layer3_outputs(320) <= '1';
    layer3_outputs(321) <= not(layer2_outputs(1993)) or (layer2_outputs(1882));
    layer3_outputs(322) <= (layer2_outputs(1028)) and not (layer2_outputs(314));
    layer3_outputs(323) <= (layer2_outputs(1894)) and not (layer2_outputs(740));
    layer3_outputs(324) <= not(layer2_outputs(2105)) or (layer2_outputs(1137));
    layer3_outputs(325) <= not(layer2_outputs(2488)) or (layer2_outputs(192));
    layer3_outputs(326) <= layer2_outputs(419);
    layer3_outputs(327) <= (layer2_outputs(688)) and not (layer2_outputs(1473));
    layer3_outputs(328) <= (layer2_outputs(901)) and not (layer2_outputs(663));
    layer3_outputs(329) <= not((layer2_outputs(1545)) and (layer2_outputs(583)));
    layer3_outputs(330) <= (layer2_outputs(1999)) and not (layer2_outputs(1858));
    layer3_outputs(331) <= not((layer2_outputs(705)) or (layer2_outputs(2129)));
    layer3_outputs(332) <= '0';
    layer3_outputs(333) <= '1';
    layer3_outputs(334) <= not((layer2_outputs(417)) or (layer2_outputs(1176)));
    layer3_outputs(335) <= not((layer2_outputs(1072)) or (layer2_outputs(2466)));
    layer3_outputs(336) <= not(layer2_outputs(11));
    layer3_outputs(337) <= not((layer2_outputs(2196)) or (layer2_outputs(1854)));
    layer3_outputs(338) <= '1';
    layer3_outputs(339) <= layer2_outputs(2250);
    layer3_outputs(340) <= (layer2_outputs(512)) or (layer2_outputs(1178));
    layer3_outputs(341) <= layer2_outputs(1184);
    layer3_outputs(342) <= not((layer2_outputs(1217)) and (layer2_outputs(298)));
    layer3_outputs(343) <= (layer2_outputs(1405)) or (layer2_outputs(1829));
    layer3_outputs(344) <= not(layer2_outputs(100));
    layer3_outputs(345) <= not(layer2_outputs(354)) or (layer2_outputs(2266));
    layer3_outputs(346) <= not(layer2_outputs(1726));
    layer3_outputs(347) <= (layer2_outputs(2397)) and (layer2_outputs(701));
    layer3_outputs(348) <= (layer2_outputs(873)) and not (layer2_outputs(1570));
    layer3_outputs(349) <= layer2_outputs(580);
    layer3_outputs(350) <= layer2_outputs(1694);
    layer3_outputs(351) <= (layer2_outputs(1065)) or (layer2_outputs(602));
    layer3_outputs(352) <= '0';
    layer3_outputs(353) <= not((layer2_outputs(473)) or (layer2_outputs(2102)));
    layer3_outputs(354) <= layer2_outputs(2384);
    layer3_outputs(355) <= not((layer2_outputs(1569)) or (layer2_outputs(2179)));
    layer3_outputs(356) <= '1';
    layer3_outputs(357) <= not(layer2_outputs(2041)) or (layer2_outputs(1767));
    layer3_outputs(358) <= (layer2_outputs(951)) or (layer2_outputs(1334));
    layer3_outputs(359) <= layer2_outputs(2310);
    layer3_outputs(360) <= not(layer2_outputs(967));
    layer3_outputs(361) <= not(layer2_outputs(1286)) or (layer2_outputs(1380));
    layer3_outputs(362) <= '1';
    layer3_outputs(363) <= not((layer2_outputs(372)) or (layer2_outputs(2245)));
    layer3_outputs(364) <= layer2_outputs(768);
    layer3_outputs(365) <= (layer2_outputs(1910)) or (layer2_outputs(1425));
    layer3_outputs(366) <= not(layer2_outputs(1565)) or (layer2_outputs(2490));
    layer3_outputs(367) <= not(layer2_outputs(1140)) or (layer2_outputs(1979));
    layer3_outputs(368) <= (layer2_outputs(762)) and (layer2_outputs(2028));
    layer3_outputs(369) <= not((layer2_outputs(1634)) and (layer2_outputs(2194)));
    layer3_outputs(370) <= layer2_outputs(271);
    layer3_outputs(371) <= '0';
    layer3_outputs(372) <= (layer2_outputs(58)) and not (layer2_outputs(819));
    layer3_outputs(373) <= not((layer2_outputs(1657)) and (layer2_outputs(1093)));
    layer3_outputs(374) <= (layer2_outputs(771)) and (layer2_outputs(366));
    layer3_outputs(375) <= (layer2_outputs(509)) and not (layer2_outputs(1784));
    layer3_outputs(376) <= '1';
    layer3_outputs(377) <= not(layer2_outputs(2064));
    layer3_outputs(378) <= not(layer2_outputs(818)) or (layer2_outputs(2229));
    layer3_outputs(379) <= not(layer2_outputs(428)) or (layer2_outputs(1965));
    layer3_outputs(380) <= layer2_outputs(2381);
    layer3_outputs(381) <= '0';
    layer3_outputs(382) <= layer2_outputs(970);
    layer3_outputs(383) <= '0';
    layer3_outputs(384) <= (layer2_outputs(2270)) or (layer2_outputs(1172));
    layer3_outputs(385) <= layer2_outputs(835);
    layer3_outputs(386) <= (layer2_outputs(626)) and not (layer2_outputs(1903));
    layer3_outputs(387) <= '1';
    layer3_outputs(388) <= not(layer2_outputs(16)) or (layer2_outputs(986));
    layer3_outputs(389) <= not((layer2_outputs(1110)) or (layer2_outputs(344)));
    layer3_outputs(390) <= layer2_outputs(2098);
    layer3_outputs(391) <= layer2_outputs(2266);
    layer3_outputs(392) <= not(layer2_outputs(20));
    layer3_outputs(393) <= layer2_outputs(2417);
    layer3_outputs(394) <= (layer2_outputs(1700)) and not (layer2_outputs(2058));
    layer3_outputs(395) <= not((layer2_outputs(305)) and (layer2_outputs(2458)));
    layer3_outputs(396) <= (layer2_outputs(1122)) or (layer2_outputs(2240));
    layer3_outputs(397) <= (layer2_outputs(1058)) or (layer2_outputs(1552));
    layer3_outputs(398) <= not((layer2_outputs(1251)) or (layer2_outputs(1325)));
    layer3_outputs(399) <= not((layer2_outputs(2224)) and (layer2_outputs(939)));
    layer3_outputs(400) <= '0';
    layer3_outputs(401) <= '1';
    layer3_outputs(402) <= not(layer2_outputs(872));
    layer3_outputs(403) <= not(layer2_outputs(93));
    layer3_outputs(404) <= not(layer2_outputs(1357));
    layer3_outputs(405) <= not(layer2_outputs(1894));
    layer3_outputs(406) <= not((layer2_outputs(2382)) or (layer2_outputs(2134)));
    layer3_outputs(407) <= (layer2_outputs(961)) and (layer2_outputs(1277));
    layer3_outputs(408) <= layer2_outputs(1538);
    layer3_outputs(409) <= not(layer2_outputs(1791)) or (layer2_outputs(1846));
    layer3_outputs(410) <= not((layer2_outputs(2142)) and (layer2_outputs(1146)));
    layer3_outputs(411) <= (layer2_outputs(2369)) and not (layer2_outputs(1014));
    layer3_outputs(412) <= (layer2_outputs(790)) or (layer2_outputs(1057));
    layer3_outputs(413) <= (layer2_outputs(1535)) and (layer2_outputs(925));
    layer3_outputs(414) <= '1';
    layer3_outputs(415) <= '0';
    layer3_outputs(416) <= not(layer2_outputs(1891));
    layer3_outputs(417) <= layer2_outputs(2035);
    layer3_outputs(418) <= layer2_outputs(150);
    layer3_outputs(419) <= not(layer2_outputs(95));
    layer3_outputs(420) <= '0';
    layer3_outputs(421) <= (layer2_outputs(1855)) and (layer2_outputs(1751));
    layer3_outputs(422) <= not(layer2_outputs(153)) or (layer2_outputs(1163));
    layer3_outputs(423) <= (layer2_outputs(2301)) and (layer2_outputs(510));
    layer3_outputs(424) <= not((layer2_outputs(993)) and (layer2_outputs(1284)));
    layer3_outputs(425) <= not(layer2_outputs(2403)) or (layer2_outputs(231));
    layer3_outputs(426) <= not(layer2_outputs(1310)) or (layer2_outputs(1022));
    layer3_outputs(427) <= layer2_outputs(363);
    layer3_outputs(428) <= not(layer2_outputs(2366));
    layer3_outputs(429) <= (layer2_outputs(1823)) and not (layer2_outputs(742));
    layer3_outputs(430) <= not(layer2_outputs(1720));
    layer3_outputs(431) <= layer2_outputs(1659);
    layer3_outputs(432) <= '1';
    layer3_outputs(433) <= layer2_outputs(2324);
    layer3_outputs(434) <= not(layer2_outputs(2471)) or (layer2_outputs(1614));
    layer3_outputs(435) <= '0';
    layer3_outputs(436) <= '1';
    layer3_outputs(437) <= not((layer2_outputs(2423)) or (layer2_outputs(3)));
    layer3_outputs(438) <= not(layer2_outputs(1158)) or (layer2_outputs(724));
    layer3_outputs(439) <= not((layer2_outputs(1858)) or (layer2_outputs(2395)));
    layer3_outputs(440) <= layer2_outputs(1286);
    layer3_outputs(441) <= not(layer2_outputs(982)) or (layer2_outputs(2477));
    layer3_outputs(442) <= not(layer2_outputs(21));
    layer3_outputs(443) <= layer2_outputs(1735);
    layer3_outputs(444) <= not(layer2_outputs(2109));
    layer3_outputs(445) <= not(layer2_outputs(1336));
    layer3_outputs(446) <= not(layer2_outputs(1086));
    layer3_outputs(447) <= not((layer2_outputs(1577)) xor (layer2_outputs(462)));
    layer3_outputs(448) <= not(layer2_outputs(1031)) or (layer2_outputs(1620));
    layer3_outputs(449) <= not(layer2_outputs(579));
    layer3_outputs(450) <= not(layer2_outputs(545));
    layer3_outputs(451) <= not(layer2_outputs(566));
    layer3_outputs(452) <= not(layer2_outputs(1379));
    layer3_outputs(453) <= layer2_outputs(427);
    layer3_outputs(454) <= layer2_outputs(1554);
    layer3_outputs(455) <= '0';
    layer3_outputs(456) <= not(layer2_outputs(2456));
    layer3_outputs(457) <= not(layer2_outputs(258));
    layer3_outputs(458) <= not((layer2_outputs(1472)) and (layer2_outputs(1616)));
    layer3_outputs(459) <= (layer2_outputs(2035)) and (layer2_outputs(434));
    layer3_outputs(460) <= (layer2_outputs(577)) or (layer2_outputs(792));
    layer3_outputs(461) <= (layer2_outputs(530)) and (layer2_outputs(2034));
    layer3_outputs(462) <= '0';
    layer3_outputs(463) <= not((layer2_outputs(2244)) or (layer2_outputs(2147)));
    layer3_outputs(464) <= not(layer2_outputs(1048));
    layer3_outputs(465) <= not((layer2_outputs(1135)) and (layer2_outputs(1166)));
    layer3_outputs(466) <= '1';
    layer3_outputs(467) <= '1';
    layer3_outputs(468) <= not((layer2_outputs(1636)) and (layer2_outputs(2087)));
    layer3_outputs(469) <= not(layer2_outputs(1544));
    layer3_outputs(470) <= layer2_outputs(46);
    layer3_outputs(471) <= layer2_outputs(1283);
    layer3_outputs(472) <= not((layer2_outputs(2279)) or (layer2_outputs(1532)));
    layer3_outputs(473) <= layer2_outputs(2478);
    layer3_outputs(474) <= not(layer2_outputs(1426));
    layer3_outputs(475) <= (layer2_outputs(1435)) or (layer2_outputs(1169));
    layer3_outputs(476) <= not(layer2_outputs(724)) or (layer2_outputs(1119));
    layer3_outputs(477) <= '0';
    layer3_outputs(478) <= (layer2_outputs(1810)) and (layer2_outputs(1647));
    layer3_outputs(479) <= layer2_outputs(1556);
    layer3_outputs(480) <= layer2_outputs(124);
    layer3_outputs(481) <= (layer2_outputs(2213)) and not (layer2_outputs(2482));
    layer3_outputs(482) <= layer2_outputs(1837);
    layer3_outputs(483) <= layer2_outputs(1203);
    layer3_outputs(484) <= layer2_outputs(2481);
    layer3_outputs(485) <= layer2_outputs(1902);
    layer3_outputs(486) <= layer2_outputs(541);
    layer3_outputs(487) <= not(layer2_outputs(80));
    layer3_outputs(488) <= not((layer2_outputs(690)) and (layer2_outputs(2371)));
    layer3_outputs(489) <= '0';
    layer3_outputs(490) <= '0';
    layer3_outputs(491) <= '0';
    layer3_outputs(492) <= (layer2_outputs(1037)) and not (layer2_outputs(587));
    layer3_outputs(493) <= '0';
    layer3_outputs(494) <= not(layer2_outputs(465)) or (layer2_outputs(478));
    layer3_outputs(495) <= (layer2_outputs(1525)) and not (layer2_outputs(1998));
    layer3_outputs(496) <= not(layer2_outputs(657));
    layer3_outputs(497) <= (layer2_outputs(1590)) and not (layer2_outputs(1239));
    layer3_outputs(498) <= '1';
    layer3_outputs(499) <= '0';
    layer3_outputs(500) <= (layer2_outputs(1754)) or (layer2_outputs(1314));
    layer3_outputs(501) <= not(layer2_outputs(2408));
    layer3_outputs(502) <= not(layer2_outputs(1594)) or (layer2_outputs(104));
    layer3_outputs(503) <= not((layer2_outputs(1404)) and (layer2_outputs(550)));
    layer3_outputs(504) <= (layer2_outputs(1328)) and not (layer2_outputs(2233));
    layer3_outputs(505) <= (layer2_outputs(132)) and (layer2_outputs(550));
    layer3_outputs(506) <= not(layer2_outputs(1852));
    layer3_outputs(507) <= (layer2_outputs(586)) and not (layer2_outputs(2469));
    layer3_outputs(508) <= layer2_outputs(341);
    layer3_outputs(509) <= layer2_outputs(2029);
    layer3_outputs(510) <= (layer2_outputs(2258)) xor (layer2_outputs(2255));
    layer3_outputs(511) <= not(layer2_outputs(2091)) or (layer2_outputs(1408));
    layer3_outputs(512) <= '1';
    layer3_outputs(513) <= (layer2_outputs(2275)) and not (layer2_outputs(1992));
    layer3_outputs(514) <= not((layer2_outputs(989)) or (layer2_outputs(2048)));
    layer3_outputs(515) <= not((layer2_outputs(597)) or (layer2_outputs(327)));
    layer3_outputs(516) <= not(layer2_outputs(1082));
    layer3_outputs(517) <= '0';
    layer3_outputs(518) <= not(layer2_outputs(1021)) or (layer2_outputs(410));
    layer3_outputs(519) <= not((layer2_outputs(1330)) xor (layer2_outputs(1187)));
    layer3_outputs(520) <= (layer2_outputs(1845)) and (layer2_outputs(1510));
    layer3_outputs(521) <= not(layer2_outputs(1026));
    layer3_outputs(522) <= not((layer2_outputs(982)) or (layer2_outputs(2525)));
    layer3_outputs(523) <= (layer2_outputs(887)) or (layer2_outputs(633));
    layer3_outputs(524) <= not((layer2_outputs(0)) and (layer2_outputs(1316)));
    layer3_outputs(525) <= '0';
    layer3_outputs(526) <= not(layer2_outputs(2159));
    layer3_outputs(527) <= not((layer2_outputs(164)) and (layer2_outputs(1948)));
    layer3_outputs(528) <= not((layer2_outputs(2540)) or (layer2_outputs(1342)));
    layer3_outputs(529) <= (layer2_outputs(1163)) and not (layer2_outputs(854));
    layer3_outputs(530) <= (layer2_outputs(544)) and not (layer2_outputs(258));
    layer3_outputs(531) <= not(layer2_outputs(775)) or (layer2_outputs(804));
    layer3_outputs(532) <= not((layer2_outputs(1937)) and (layer2_outputs(779)));
    layer3_outputs(533) <= '1';
    layer3_outputs(534) <= (layer2_outputs(794)) and not (layer2_outputs(42));
    layer3_outputs(535) <= not(layer2_outputs(1025)) or (layer2_outputs(282));
    layer3_outputs(536) <= not(layer2_outputs(376));
    layer3_outputs(537) <= '0';
    layer3_outputs(538) <= not(layer2_outputs(1466));
    layer3_outputs(539) <= '0';
    layer3_outputs(540) <= (layer2_outputs(2304)) and (layer2_outputs(899));
    layer3_outputs(541) <= (layer2_outputs(2336)) and (layer2_outputs(2499));
    layer3_outputs(542) <= '0';
    layer3_outputs(543) <= layer2_outputs(1872);
    layer3_outputs(544) <= (layer2_outputs(755)) and (layer2_outputs(412));
    layer3_outputs(545) <= not(layer2_outputs(2232));
    layer3_outputs(546) <= not(layer2_outputs(775));
    layer3_outputs(547) <= not((layer2_outputs(2396)) and (layer2_outputs(2037)));
    layer3_outputs(548) <= '0';
    layer3_outputs(549) <= '0';
    layer3_outputs(550) <= not(layer2_outputs(527)) or (layer2_outputs(995));
    layer3_outputs(551) <= not(layer2_outputs(187));
    layer3_outputs(552) <= (layer2_outputs(2420)) and not (layer2_outputs(2011));
    layer3_outputs(553) <= not(layer2_outputs(2231));
    layer3_outputs(554) <= not(layer2_outputs(2351));
    layer3_outputs(555) <= not((layer2_outputs(1395)) and (layer2_outputs(1980)));
    layer3_outputs(556) <= not(layer2_outputs(2500)) or (layer2_outputs(1947));
    layer3_outputs(557) <= (layer2_outputs(2017)) and (layer2_outputs(141));
    layer3_outputs(558) <= (layer2_outputs(1421)) and not (layer2_outputs(725));
    layer3_outputs(559) <= layer2_outputs(1155);
    layer3_outputs(560) <= not((layer2_outputs(2184)) or (layer2_outputs(367)));
    layer3_outputs(561) <= layer2_outputs(1036);
    layer3_outputs(562) <= not(layer2_outputs(2135)) or (layer2_outputs(2447));
    layer3_outputs(563) <= (layer2_outputs(1926)) and not (layer2_outputs(1498));
    layer3_outputs(564) <= not((layer2_outputs(1016)) and (layer2_outputs(1439)));
    layer3_outputs(565) <= '1';
    layer3_outputs(566) <= not((layer2_outputs(1099)) and (layer2_outputs(1214)));
    layer3_outputs(567) <= not((layer2_outputs(1381)) or (layer2_outputs(286)));
    layer3_outputs(568) <= not((layer2_outputs(700)) xor (layer2_outputs(1059)));
    layer3_outputs(569) <= not(layer2_outputs(1221));
    layer3_outputs(570) <= not((layer2_outputs(2211)) and (layer2_outputs(108)));
    layer3_outputs(571) <= layer2_outputs(2539);
    layer3_outputs(572) <= not((layer2_outputs(1576)) and (layer2_outputs(784)));
    layer3_outputs(573) <= (layer2_outputs(818)) xor (layer2_outputs(145));
    layer3_outputs(574) <= layer2_outputs(29);
    layer3_outputs(575) <= (layer2_outputs(167)) or (layer2_outputs(1735));
    layer3_outputs(576) <= not(layer2_outputs(1260)) or (layer2_outputs(2280));
    layer3_outputs(577) <= '1';
    layer3_outputs(578) <= not(layer2_outputs(484));
    layer3_outputs(579) <= not(layer2_outputs(999)) or (layer2_outputs(1257));
    layer3_outputs(580) <= '1';
    layer3_outputs(581) <= (layer2_outputs(127)) and not (layer2_outputs(43));
    layer3_outputs(582) <= not(layer2_outputs(1073));
    layer3_outputs(583) <= not((layer2_outputs(1117)) or (layer2_outputs(754)));
    layer3_outputs(584) <= not(layer2_outputs(235));
    layer3_outputs(585) <= layer2_outputs(2091);
    layer3_outputs(586) <= (layer2_outputs(578)) and (layer2_outputs(173));
    layer3_outputs(587) <= '1';
    layer3_outputs(588) <= not(layer2_outputs(490));
    layer3_outputs(589) <= not((layer2_outputs(1102)) or (layer2_outputs(622)));
    layer3_outputs(590) <= not(layer2_outputs(1843)) or (layer2_outputs(2458));
    layer3_outputs(591) <= '1';
    layer3_outputs(592) <= not((layer2_outputs(2157)) or (layer2_outputs(598)));
    layer3_outputs(593) <= layer2_outputs(1550);
    layer3_outputs(594) <= '0';
    layer3_outputs(595) <= not((layer2_outputs(868)) and (layer2_outputs(1622)));
    layer3_outputs(596) <= not(layer2_outputs(1445)) or (layer2_outputs(1630));
    layer3_outputs(597) <= not(layer2_outputs(1973));
    layer3_outputs(598) <= layer2_outputs(1923);
    layer3_outputs(599) <= not(layer2_outputs(81)) or (layer2_outputs(106));
    layer3_outputs(600) <= (layer2_outputs(1750)) and (layer2_outputs(255));
    layer3_outputs(601) <= not((layer2_outputs(783)) and (layer2_outputs(988)));
    layer3_outputs(602) <= layer2_outputs(1183);
    layer3_outputs(603) <= not(layer2_outputs(1921));
    layer3_outputs(604) <= (layer2_outputs(1882)) and (layer2_outputs(536));
    layer3_outputs(605) <= not(layer2_outputs(1757));
    layer3_outputs(606) <= layer2_outputs(2282);
    layer3_outputs(607) <= not(layer2_outputs(39));
    layer3_outputs(608) <= not(layer2_outputs(1155));
    layer3_outputs(609) <= layer2_outputs(1821);
    layer3_outputs(610) <= (layer2_outputs(992)) and not (layer2_outputs(845));
    layer3_outputs(611) <= '0';
    layer3_outputs(612) <= not(layer2_outputs(1881));
    layer3_outputs(613) <= not((layer2_outputs(1573)) or (layer2_outputs(1527)));
    layer3_outputs(614) <= '1';
    layer3_outputs(615) <= (layer2_outputs(977)) and not (layer2_outputs(324));
    layer3_outputs(616) <= layer2_outputs(1703);
    layer3_outputs(617) <= not((layer2_outputs(652)) or (layer2_outputs(1095)));
    layer3_outputs(618) <= not((layer2_outputs(2209)) and (layer2_outputs(1432)));
    layer3_outputs(619) <= not(layer2_outputs(1560)) or (layer2_outputs(660));
    layer3_outputs(620) <= not((layer2_outputs(1391)) or (layer2_outputs(1338)));
    layer3_outputs(621) <= not(layer2_outputs(556));
    layer3_outputs(622) <= (layer2_outputs(461)) xor (layer2_outputs(1401));
    layer3_outputs(623) <= not(layer2_outputs(638));
    layer3_outputs(624) <= '1';
    layer3_outputs(625) <= layer2_outputs(594);
    layer3_outputs(626) <= '1';
    layer3_outputs(627) <= (layer2_outputs(690)) and not (layer2_outputs(1012));
    layer3_outputs(628) <= not(layer2_outputs(1078)) or (layer2_outputs(1574));
    layer3_outputs(629) <= '0';
    layer3_outputs(630) <= not(layer2_outputs(155));
    layer3_outputs(631) <= layer2_outputs(1460);
    layer3_outputs(632) <= (layer2_outputs(2434)) or (layer2_outputs(1146));
    layer3_outputs(633) <= layer2_outputs(2366);
    layer3_outputs(634) <= not(layer2_outputs(1293));
    layer3_outputs(635) <= not((layer2_outputs(1323)) or (layer2_outputs(2002)));
    layer3_outputs(636) <= '0';
    layer3_outputs(637) <= not(layer2_outputs(1476)) or (layer2_outputs(2106));
    layer3_outputs(638) <= not(layer2_outputs(2514));
    layer3_outputs(639) <= not(layer2_outputs(31));
    layer3_outputs(640) <= not(layer2_outputs(1728));
    layer3_outputs(641) <= (layer2_outputs(2033)) and (layer2_outputs(1149));
    layer3_outputs(642) <= (layer2_outputs(2208)) and (layer2_outputs(1963));
    layer3_outputs(643) <= not(layer2_outputs(193));
    layer3_outputs(644) <= layer2_outputs(2360);
    layer3_outputs(645) <= not(layer2_outputs(1938));
    layer3_outputs(646) <= '0';
    layer3_outputs(647) <= '1';
    layer3_outputs(648) <= layer2_outputs(1952);
    layer3_outputs(649) <= not(layer2_outputs(1610));
    layer3_outputs(650) <= not(layer2_outputs(1274));
    layer3_outputs(651) <= (layer2_outputs(1142)) and (layer2_outputs(1217));
    layer3_outputs(652) <= not(layer2_outputs(1113)) or (layer2_outputs(668));
    layer3_outputs(653) <= not(layer2_outputs(661)) or (layer2_outputs(1817));
    layer3_outputs(654) <= not((layer2_outputs(79)) and (layer2_outputs(1037)));
    layer3_outputs(655) <= not(layer2_outputs(2004));
    layer3_outputs(656) <= not((layer2_outputs(133)) or (layer2_outputs(427)));
    layer3_outputs(657) <= '1';
    layer3_outputs(658) <= (layer2_outputs(122)) or (layer2_outputs(1581));
    layer3_outputs(659) <= not(layer2_outputs(902)) or (layer2_outputs(497));
    layer3_outputs(660) <= not(layer2_outputs(2518));
    layer3_outputs(661) <= not(layer2_outputs(1185)) or (layer2_outputs(2289));
    layer3_outputs(662) <= (layer2_outputs(909)) and (layer2_outputs(582));
    layer3_outputs(663) <= '0';
    layer3_outputs(664) <= not(layer2_outputs(1393));
    layer3_outputs(665) <= not(layer2_outputs(2079));
    layer3_outputs(666) <= not(layer2_outputs(1900));
    layer3_outputs(667) <= not(layer2_outputs(1641));
    layer3_outputs(668) <= not((layer2_outputs(359)) xor (layer2_outputs(1835)));
    layer3_outputs(669) <= (layer2_outputs(345)) or (layer2_outputs(2137));
    layer3_outputs(670) <= '1';
    layer3_outputs(671) <= '0';
    layer3_outputs(672) <= layer2_outputs(445);
    layer3_outputs(673) <= '1';
    layer3_outputs(674) <= not(layer2_outputs(2176));
    layer3_outputs(675) <= not(layer2_outputs(2165));
    layer3_outputs(676) <= not(layer2_outputs(620)) or (layer2_outputs(2380));
    layer3_outputs(677) <= not(layer2_outputs(897));
    layer3_outputs(678) <= not(layer2_outputs(824));
    layer3_outputs(679) <= layer2_outputs(2110);
    layer3_outputs(680) <= '0';
    layer3_outputs(681) <= (layer2_outputs(635)) and not (layer2_outputs(555));
    layer3_outputs(682) <= not((layer2_outputs(592)) or (layer2_outputs(94)));
    layer3_outputs(683) <= (layer2_outputs(800)) and not (layer2_outputs(1008));
    layer3_outputs(684) <= layer2_outputs(1553);
    layer3_outputs(685) <= '0';
    layer3_outputs(686) <= (layer2_outputs(406)) or (layer2_outputs(1087));
    layer3_outputs(687) <= '1';
    layer3_outputs(688) <= layer2_outputs(2317);
    layer3_outputs(689) <= not((layer2_outputs(1933)) xor (layer2_outputs(2389)));
    layer3_outputs(690) <= (layer2_outputs(1939)) or (layer2_outputs(214));
    layer3_outputs(691) <= not(layer2_outputs(66)) or (layer2_outputs(1732));
    layer3_outputs(692) <= not(layer2_outputs(449));
    layer3_outputs(693) <= layer2_outputs(975);
    layer3_outputs(694) <= (layer2_outputs(605)) or (layer2_outputs(2383));
    layer3_outputs(695) <= not((layer2_outputs(1436)) or (layer2_outputs(1062)));
    layer3_outputs(696) <= not(layer2_outputs(161));
    layer3_outputs(697) <= not(layer2_outputs(204));
    layer3_outputs(698) <= not(layer2_outputs(1973)) or (layer2_outputs(1239));
    layer3_outputs(699) <= not((layer2_outputs(281)) and (layer2_outputs(1779)));
    layer3_outputs(700) <= layer2_outputs(820);
    layer3_outputs(701) <= layer2_outputs(639);
    layer3_outputs(702) <= '0';
    layer3_outputs(703) <= not((layer2_outputs(304)) and (layer2_outputs(1302)));
    layer3_outputs(704) <= not(layer2_outputs(1444));
    layer3_outputs(705) <= not(layer2_outputs(421));
    layer3_outputs(706) <= not((layer2_outputs(851)) or (layer2_outputs(1125)));
    layer3_outputs(707) <= layer2_outputs(1996);
    layer3_outputs(708) <= not(layer2_outputs(239));
    layer3_outputs(709) <= not((layer2_outputs(1594)) and (layer2_outputs(919)));
    layer3_outputs(710) <= '1';
    layer3_outputs(711) <= (layer2_outputs(1169)) and not (layer2_outputs(1809));
    layer3_outputs(712) <= layer2_outputs(1416);
    layer3_outputs(713) <= layer2_outputs(1746);
    layer3_outputs(714) <= (layer2_outputs(93)) or (layer2_outputs(1223));
    layer3_outputs(715) <= (layer2_outputs(2156)) and not (layer2_outputs(677));
    layer3_outputs(716) <= layer2_outputs(334);
    layer3_outputs(717) <= not((layer2_outputs(1609)) and (layer2_outputs(1482)));
    layer3_outputs(718) <= not((layer2_outputs(325)) xor (layer2_outputs(405)));
    layer3_outputs(719) <= not(layer2_outputs(2132)) or (layer2_outputs(1250));
    layer3_outputs(720) <= not(layer2_outputs(1326)) or (layer2_outputs(2115));
    layer3_outputs(721) <= not(layer2_outputs(2232));
    layer3_outputs(722) <= (layer2_outputs(1893)) or (layer2_outputs(1688));
    layer3_outputs(723) <= not((layer2_outputs(1016)) and (layer2_outputs(844)));
    layer3_outputs(724) <= not((layer2_outputs(1577)) and (layer2_outputs(2238)));
    layer3_outputs(725) <= layer2_outputs(2127);
    layer3_outputs(726) <= layer2_outputs(1922);
    layer3_outputs(727) <= layer2_outputs(645);
    layer3_outputs(728) <= layer2_outputs(1599);
    layer3_outputs(729) <= not(layer2_outputs(621));
    layer3_outputs(730) <= layer2_outputs(1355);
    layer3_outputs(731) <= layer2_outputs(234);
    layer3_outputs(732) <= not(layer2_outputs(929));
    layer3_outputs(733) <= layer2_outputs(251);
    layer3_outputs(734) <= (layer2_outputs(1671)) and not (layer2_outputs(1617));
    layer3_outputs(735) <= (layer2_outputs(891)) and not (layer2_outputs(2163));
    layer3_outputs(736) <= layer2_outputs(2467);
    layer3_outputs(737) <= '1';
    layer3_outputs(738) <= not(layer2_outputs(299)) or (layer2_outputs(464));
    layer3_outputs(739) <= layer2_outputs(136);
    layer3_outputs(740) <= '0';
    layer3_outputs(741) <= layer2_outputs(890);
    layer3_outputs(742) <= (layer2_outputs(2363)) and not (layer2_outputs(1506));
    layer3_outputs(743) <= '0';
    layer3_outputs(744) <= (layer2_outputs(2025)) and not (layer2_outputs(2039));
    layer3_outputs(745) <= not(layer2_outputs(480)) or (layer2_outputs(1491));
    layer3_outputs(746) <= not(layer2_outputs(2299));
    layer3_outputs(747) <= (layer2_outputs(2454)) and (layer2_outputs(1387));
    layer3_outputs(748) <= not(layer2_outputs(1951)) or (layer2_outputs(1246));
    layer3_outputs(749) <= not((layer2_outputs(2536)) or (layer2_outputs(1628)));
    layer3_outputs(750) <= layer2_outputs(2334);
    layer3_outputs(751) <= not(layer2_outputs(1509));
    layer3_outputs(752) <= (layer2_outputs(1290)) and not (layer2_outputs(1629));
    layer3_outputs(753) <= layer2_outputs(1664);
    layer3_outputs(754) <= not(layer2_outputs(1147));
    layer3_outputs(755) <= layer2_outputs(2216);
    layer3_outputs(756) <= (layer2_outputs(2254)) xor (layer2_outputs(2049));
    layer3_outputs(757) <= not((layer2_outputs(1446)) or (layer2_outputs(808)));
    layer3_outputs(758) <= '0';
    layer3_outputs(759) <= (layer2_outputs(309)) and not (layer2_outputs(1400));
    layer3_outputs(760) <= not(layer2_outputs(720)) or (layer2_outputs(1441));
    layer3_outputs(761) <= (layer2_outputs(797)) or (layer2_outputs(1148));
    layer3_outputs(762) <= not((layer2_outputs(2153)) xor (layer2_outputs(1863)));
    layer3_outputs(763) <= '1';
    layer3_outputs(764) <= not(layer2_outputs(1347));
    layer3_outputs(765) <= (layer2_outputs(1356)) and (layer2_outputs(1120));
    layer3_outputs(766) <= not((layer2_outputs(486)) and (layer2_outputs(2318)));
    layer3_outputs(767) <= (layer2_outputs(553)) and not (layer2_outputs(1196));
    layer3_outputs(768) <= not(layer2_outputs(158)) or (layer2_outputs(2123));
    layer3_outputs(769) <= layer2_outputs(1775);
    layer3_outputs(770) <= '0';
    layer3_outputs(771) <= not(layer2_outputs(1443));
    layer3_outputs(772) <= '1';
    layer3_outputs(773) <= not(layer2_outputs(733));
    layer3_outputs(774) <= (layer2_outputs(1505)) and (layer2_outputs(1671));
    layer3_outputs(775) <= not(layer2_outputs(1769));
    layer3_outputs(776) <= (layer2_outputs(2193)) or (layer2_outputs(231));
    layer3_outputs(777) <= (layer2_outputs(2170)) and (layer2_outputs(1162));
    layer3_outputs(778) <= (layer2_outputs(2479)) and not (layer2_outputs(2427));
    layer3_outputs(779) <= not((layer2_outputs(1495)) xor (layer2_outputs(37)));
    layer3_outputs(780) <= (layer2_outputs(1189)) and not (layer2_outputs(2354));
    layer3_outputs(781) <= (layer2_outputs(2339)) and (layer2_outputs(1546));
    layer3_outputs(782) <= not((layer2_outputs(968)) xor (layer2_outputs(943)));
    layer3_outputs(783) <= not((layer2_outputs(736)) or (layer2_outputs(1329)));
    layer3_outputs(784) <= (layer2_outputs(1182)) or (layer2_outputs(1426));
    layer3_outputs(785) <= layer2_outputs(957);
    layer3_outputs(786) <= '1';
    layer3_outputs(787) <= layer2_outputs(2331);
    layer3_outputs(788) <= not(layer2_outputs(2519)) or (layer2_outputs(965));
    layer3_outputs(789) <= not((layer2_outputs(2461)) or (layer2_outputs(1154)));
    layer3_outputs(790) <= (layer2_outputs(2276)) and (layer2_outputs(2431));
    layer3_outputs(791) <= not(layer2_outputs(2121));
    layer3_outputs(792) <= not(layer2_outputs(2473)) or (layer2_outputs(804));
    layer3_outputs(793) <= layer2_outputs(2234);
    layer3_outputs(794) <= not(layer2_outputs(1869));
    layer3_outputs(795) <= layer2_outputs(1840);
    layer3_outputs(796) <= '0';
    layer3_outputs(797) <= not((layer2_outputs(1041)) or (layer2_outputs(1063)));
    layer3_outputs(798) <= not((layer2_outputs(2256)) or (layer2_outputs(887)));
    layer3_outputs(799) <= layer2_outputs(627);
    layer3_outputs(800) <= layer2_outputs(15);
    layer3_outputs(801) <= (layer2_outputs(1622)) and (layer2_outputs(1788));
    layer3_outputs(802) <= (layer2_outputs(714)) and not (layer2_outputs(1429));
    layer3_outputs(803) <= (layer2_outputs(40)) and not (layer2_outputs(1245));
    layer3_outputs(804) <= not(layer2_outputs(1569));
    layer3_outputs(805) <= layer2_outputs(711);
    layer3_outputs(806) <= (layer2_outputs(2553)) and not (layer2_outputs(1731));
    layer3_outputs(807) <= layer2_outputs(2385);
    layer3_outputs(808) <= '0';
    layer3_outputs(809) <= not((layer2_outputs(1875)) and (layer2_outputs(794)));
    layer3_outputs(810) <= not((layer2_outputs(1979)) or (layer2_outputs(2271)));
    layer3_outputs(811) <= layer2_outputs(1802);
    layer3_outputs(812) <= layer2_outputs(1261);
    layer3_outputs(813) <= (layer2_outputs(147)) and not (layer2_outputs(225));
    layer3_outputs(814) <= (layer2_outputs(1170)) and not (layer2_outputs(572));
    layer3_outputs(815) <= (layer2_outputs(248)) and not (layer2_outputs(2056));
    layer3_outputs(816) <= (layer2_outputs(2520)) or (layer2_outputs(735));
    layer3_outputs(817) <= not(layer2_outputs(1868));
    layer3_outputs(818) <= (layer2_outputs(1385)) and not (layer2_outputs(1713));
    layer3_outputs(819) <= not(layer2_outputs(1771));
    layer3_outputs(820) <= not((layer2_outputs(92)) or (layer2_outputs(651)));
    layer3_outputs(821) <= not((layer2_outputs(1561)) and (layer2_outputs(1240)));
    layer3_outputs(822) <= not(layer2_outputs(1495));
    layer3_outputs(823) <= not(layer2_outputs(26));
    layer3_outputs(824) <= not(layer2_outputs(741));
    layer3_outputs(825) <= not(layer2_outputs(22));
    layer3_outputs(826) <= (layer2_outputs(523)) and not (layer2_outputs(2227));
    layer3_outputs(827) <= not(layer2_outputs(439));
    layer3_outputs(828) <= layer2_outputs(82);
    layer3_outputs(829) <= not(layer2_outputs(1230));
    layer3_outputs(830) <= (layer2_outputs(863)) and not (layer2_outputs(222));
    layer3_outputs(831) <= not(layer2_outputs(2503)) or (layer2_outputs(189));
    layer3_outputs(832) <= '1';
    layer3_outputs(833) <= not(layer2_outputs(252)) or (layer2_outputs(1211));
    layer3_outputs(834) <= layer2_outputs(274);
    layer3_outputs(835) <= not(layer2_outputs(1430)) or (layer2_outputs(47));
    layer3_outputs(836) <= '0';
    layer3_outputs(837) <= (layer2_outputs(1262)) or (layer2_outputs(1257));
    layer3_outputs(838) <= layer2_outputs(1675);
    layer3_outputs(839) <= not(layer2_outputs(482));
    layer3_outputs(840) <= '0';
    layer3_outputs(841) <= layer2_outputs(1345);
    layer3_outputs(842) <= (layer2_outputs(302)) or (layer2_outputs(2406));
    layer3_outputs(843) <= layer2_outputs(2531);
    layer3_outputs(844) <= '1';
    layer3_outputs(845) <= not((layer2_outputs(1431)) or (layer2_outputs(1888)));
    layer3_outputs(846) <= layer2_outputs(1168);
    layer3_outputs(847) <= not(layer2_outputs(1034));
    layer3_outputs(848) <= '0';
    layer3_outputs(849) <= not(layer2_outputs(2481)) or (layer2_outputs(237));
    layer3_outputs(850) <= not(layer2_outputs(1373));
    layer3_outputs(851) <= not(layer2_outputs(2076)) or (layer2_outputs(1684));
    layer3_outputs(852) <= (layer2_outputs(2113)) or (layer2_outputs(861));
    layer3_outputs(853) <= not((layer2_outputs(1043)) and (layer2_outputs(478)));
    layer3_outputs(854) <= layer2_outputs(1126);
    layer3_outputs(855) <= (layer2_outputs(1856)) and (layer2_outputs(1298));
    layer3_outputs(856) <= '1';
    layer3_outputs(857) <= not(layer2_outputs(450)) or (layer2_outputs(348));
    layer3_outputs(858) <= not(layer2_outputs(628));
    layer3_outputs(859) <= not(layer2_outputs(562)) or (layer2_outputs(2349));
    layer3_outputs(860) <= '0';
    layer3_outputs(861) <= '0';
    layer3_outputs(862) <= (layer2_outputs(1449)) and not (layer2_outputs(136));
    layer3_outputs(863) <= (layer2_outputs(2101)) and (layer2_outputs(1000));
    layer3_outputs(864) <= '0';
    layer3_outputs(865) <= not(layer2_outputs(1043)) or (layer2_outputs(1548));
    layer3_outputs(866) <= not(layer2_outputs(139)) or (layer2_outputs(1173));
    layer3_outputs(867) <= not((layer2_outputs(1907)) or (layer2_outputs(941)));
    layer3_outputs(868) <= layer2_outputs(1489);
    layer3_outputs(869) <= layer2_outputs(2556);
    layer3_outputs(870) <= '1';
    layer3_outputs(871) <= not((layer2_outputs(1888)) or (layer2_outputs(210)));
    layer3_outputs(872) <= not((layer2_outputs(858)) and (layer2_outputs(1707)));
    layer3_outputs(873) <= not((layer2_outputs(1680)) xor (layer2_outputs(409)));
    layer3_outputs(874) <= not(layer2_outputs(1353));
    layer3_outputs(875) <= (layer2_outputs(2373)) and (layer2_outputs(1702));
    layer3_outputs(876) <= '1';
    layer3_outputs(877) <= layer2_outputs(1946);
    layer3_outputs(878) <= layer2_outputs(1274);
    layer3_outputs(879) <= '1';
    layer3_outputs(880) <= '0';
    layer3_outputs(881) <= not((layer2_outputs(168)) or (layer2_outputs(2319)));
    layer3_outputs(882) <= not(layer2_outputs(71)) or (layer2_outputs(1730));
    layer3_outputs(883) <= (layer2_outputs(1262)) and not (layer2_outputs(143));
    layer3_outputs(884) <= not((layer2_outputs(569)) and (layer2_outputs(1064)));
    layer3_outputs(885) <= (layer2_outputs(648)) xor (layer2_outputs(521));
    layer3_outputs(886) <= layer2_outputs(152);
    layer3_outputs(887) <= not(layer2_outputs(1914));
    layer3_outputs(888) <= not(layer2_outputs(810)) or (layer2_outputs(2120));
    layer3_outputs(889) <= not((layer2_outputs(294)) or (layer2_outputs(440)));
    layer3_outputs(890) <= (layer2_outputs(921)) and (layer2_outputs(2058));
    layer3_outputs(891) <= layer2_outputs(825);
    layer3_outputs(892) <= '1';
    layer3_outputs(893) <= not(layer2_outputs(205));
    layer3_outputs(894) <= not(layer2_outputs(2119)) or (layer2_outputs(476));
    layer3_outputs(895) <= not((layer2_outputs(699)) and (layer2_outputs(1414)));
    layer3_outputs(896) <= not(layer2_outputs(732));
    layer3_outputs(897) <= not(layer2_outputs(1207)) or (layer2_outputs(2034));
    layer3_outputs(898) <= layer2_outputs(1041);
    layer3_outputs(899) <= (layer2_outputs(322)) and not (layer2_outputs(84));
    layer3_outputs(900) <= not((layer2_outputs(1364)) or (layer2_outputs(2340)));
    layer3_outputs(901) <= not(layer2_outputs(2535));
    layer3_outputs(902) <= not(layer2_outputs(1862));
    layer3_outputs(903) <= not(layer2_outputs(1829)) or (layer2_outputs(1736));
    layer3_outputs(904) <= layer2_outputs(1619);
    layer3_outputs(905) <= layer2_outputs(842);
    layer3_outputs(906) <= not(layer2_outputs(760));
    layer3_outputs(907) <= not(layer2_outputs(1825)) or (layer2_outputs(2189));
    layer3_outputs(908) <= not(layer2_outputs(1219)) or (layer2_outputs(1214));
    layer3_outputs(909) <= '0';
    layer3_outputs(910) <= not((layer2_outputs(1537)) or (layer2_outputs(1969)));
    layer3_outputs(911) <= not(layer2_outputs(81));
    layer3_outputs(912) <= '0';
    layer3_outputs(913) <= layer2_outputs(156);
    layer3_outputs(914) <= not(layer2_outputs(1523));
    layer3_outputs(915) <= '1';
    layer3_outputs(916) <= not(layer2_outputs(2336));
    layer3_outputs(917) <= (layer2_outputs(151)) and not (layer2_outputs(2384));
    layer3_outputs(918) <= not(layer2_outputs(1459)) or (layer2_outputs(6));
    layer3_outputs(919) <= not((layer2_outputs(2368)) and (layer2_outputs(1443)));
    layer3_outputs(920) <= layer2_outputs(2466);
    layer3_outputs(921) <= not(layer2_outputs(1841)) or (layer2_outputs(1148));
    layer3_outputs(922) <= not(layer2_outputs(875)) or (layer2_outputs(905));
    layer3_outputs(923) <= not(layer2_outputs(1366));
    layer3_outputs(924) <= '0';
    layer3_outputs(925) <= (layer2_outputs(1871)) xor (layer2_outputs(96));
    layer3_outputs(926) <= '1';
    layer3_outputs(927) <= (layer2_outputs(2426)) xor (layer2_outputs(1981));
    layer3_outputs(928) <= '0';
    layer3_outputs(929) <= '1';
    layer3_outputs(930) <= not((layer2_outputs(2186)) and (layer2_outputs(2329)));
    layer3_outputs(931) <= not((layer2_outputs(1400)) and (layer2_outputs(2377)));
    layer3_outputs(932) <= not((layer2_outputs(67)) and (layer2_outputs(1831)));
    layer3_outputs(933) <= (layer2_outputs(1584)) and not (layer2_outputs(870));
    layer3_outputs(934) <= layer2_outputs(2204);
    layer3_outputs(935) <= not((layer2_outputs(1530)) xor (layer2_outputs(317)));
    layer3_outputs(936) <= layer2_outputs(1480);
    layer3_outputs(937) <= '1';
    layer3_outputs(938) <= '1';
    layer3_outputs(939) <= not(layer2_outputs(1354)) or (layer2_outputs(170));
    layer3_outputs(940) <= not((layer2_outputs(2516)) and (layer2_outputs(1264)));
    layer3_outputs(941) <= layer2_outputs(1767);
    layer3_outputs(942) <= not((layer2_outputs(658)) xor (layer2_outputs(2248)));
    layer3_outputs(943) <= '0';
    layer3_outputs(944) <= (layer2_outputs(1277)) and not (layer2_outputs(1997));
    layer3_outputs(945) <= (layer2_outputs(1127)) or (layer2_outputs(517));
    layer3_outputs(946) <= not(layer2_outputs(2162));
    layer3_outputs(947) <= not(layer2_outputs(1667));
    layer3_outputs(948) <= not((layer2_outputs(457)) or (layer2_outputs(278)));
    layer3_outputs(949) <= not(layer2_outputs(531));
    layer3_outputs(950) <= not(layer2_outputs(1914)) or (layer2_outputs(1645));
    layer3_outputs(951) <= not((layer2_outputs(673)) and (layer2_outputs(1940)));
    layer3_outputs(952) <= layer2_outputs(1677);
    layer3_outputs(953) <= (layer2_outputs(1001)) and (layer2_outputs(97));
    layer3_outputs(954) <= layer2_outputs(849);
    layer3_outputs(955) <= not((layer2_outputs(1555)) and (layer2_outputs(1793)));
    layer3_outputs(956) <= (layer2_outputs(1923)) and not (layer2_outputs(410));
    layer3_outputs(957) <= not((layer2_outputs(1799)) and (layer2_outputs(917)));
    layer3_outputs(958) <= (layer2_outputs(1598)) or (layer2_outputs(1807));
    layer3_outputs(959) <= (layer2_outputs(717)) or (layer2_outputs(1023));
    layer3_outputs(960) <= (layer2_outputs(337)) and (layer2_outputs(566));
    layer3_outputs(961) <= not(layer2_outputs(2352)) or (layer2_outputs(203));
    layer3_outputs(962) <= (layer2_outputs(542)) or (layer2_outputs(2383));
    layer3_outputs(963) <= (layer2_outputs(1471)) or (layer2_outputs(145));
    layer3_outputs(964) <= not(layer2_outputs(2129));
    layer3_outputs(965) <= '0';
    layer3_outputs(966) <= (layer2_outputs(701)) and not (layer2_outputs(420));
    layer3_outputs(967) <= layer2_outputs(1685);
    layer3_outputs(968) <= not((layer2_outputs(1319)) or (layer2_outputs(1061)));
    layer3_outputs(969) <= layer2_outputs(769);
    layer3_outputs(970) <= not(layer2_outputs(1885)) or (layer2_outputs(1308));
    layer3_outputs(971) <= layer2_outputs(294);
    layer3_outputs(972) <= not(layer2_outputs(1249));
    layer3_outputs(973) <= layer2_outputs(253);
    layer3_outputs(974) <= not((layer2_outputs(129)) and (layer2_outputs(1378)));
    layer3_outputs(975) <= not(layer2_outputs(466));
    layer3_outputs(976) <= '1';
    layer3_outputs(977) <= not(layer2_outputs(986));
    layer3_outputs(978) <= '0';
    layer3_outputs(979) <= (layer2_outputs(64)) and not (layer2_outputs(1718));
    layer3_outputs(980) <= '0';
    layer3_outputs(981) <= not(layer2_outputs(481)) or (layer2_outputs(124));
    layer3_outputs(982) <= not(layer2_outputs(2059));
    layer3_outputs(983) <= layer2_outputs(505);
    layer3_outputs(984) <= not(layer2_outputs(1593)) or (layer2_outputs(1628));
    layer3_outputs(985) <= '0';
    layer3_outputs(986) <= (layer2_outputs(212)) or (layer2_outputs(89));
    layer3_outputs(987) <= not(layer2_outputs(585));
    layer3_outputs(988) <= layer2_outputs(1890);
    layer3_outputs(989) <= '0';
    layer3_outputs(990) <= (layer2_outputs(2299)) and not (layer2_outputs(855));
    layer3_outputs(991) <= '0';
    layer3_outputs(992) <= '0';
    layer3_outputs(993) <= not(layer2_outputs(1530)) or (layer2_outputs(185));
    layer3_outputs(994) <= (layer2_outputs(1482)) or (layer2_outputs(1080));
    layer3_outputs(995) <= not((layer2_outputs(2300)) or (layer2_outputs(1076)));
    layer3_outputs(996) <= not((layer2_outputs(1650)) or (layer2_outputs(220)));
    layer3_outputs(997) <= '0';
    layer3_outputs(998) <= not(layer2_outputs(14));
    layer3_outputs(999) <= not(layer2_outputs(456)) or (layer2_outputs(2062));
    layer3_outputs(1000) <= not((layer2_outputs(5)) or (layer2_outputs(945)));
    layer3_outputs(1001) <= '1';
    layer3_outputs(1002) <= (layer2_outputs(1060)) and not (layer2_outputs(1067));
    layer3_outputs(1003) <= layer2_outputs(117);
    layer3_outputs(1004) <= '0';
    layer3_outputs(1005) <= layer2_outputs(2021);
    layer3_outputs(1006) <= not((layer2_outputs(2316)) or (layer2_outputs(561)));
    layer3_outputs(1007) <= not(layer2_outputs(444));
    layer3_outputs(1008) <= not((layer2_outputs(575)) and (layer2_outputs(1507)));
    layer3_outputs(1009) <= not(layer2_outputs(2306));
    layer3_outputs(1010) <= (layer2_outputs(2493)) or (layer2_outputs(366));
    layer3_outputs(1011) <= layer2_outputs(1620);
    layer3_outputs(1012) <= (layer2_outputs(680)) or (layer2_outputs(23));
    layer3_outputs(1013) <= not(layer2_outputs(603));
    layer3_outputs(1014) <= not(layer2_outputs(1823));
    layer3_outputs(1015) <= '0';
    layer3_outputs(1016) <= not((layer2_outputs(861)) xor (layer2_outputs(90)));
    layer3_outputs(1017) <= not(layer2_outputs(1651)) or (layer2_outputs(1848));
    layer3_outputs(1018) <= not(layer2_outputs(1676));
    layer3_outputs(1019) <= not(layer2_outputs(423)) or (layer2_outputs(744));
    layer3_outputs(1020) <= (layer2_outputs(2505)) or (layer2_outputs(607));
    layer3_outputs(1021) <= '0';
    layer3_outputs(1022) <= layer2_outputs(1060);
    layer3_outputs(1023) <= not((layer2_outputs(73)) and (layer2_outputs(754)));
    layer3_outputs(1024) <= not(layer2_outputs(1811));
    layer3_outputs(1025) <= (layer2_outputs(1578)) or (layer2_outputs(2003));
    layer3_outputs(1026) <= layer2_outputs(1641);
    layer3_outputs(1027) <= not(layer2_outputs(707));
    layer3_outputs(1028) <= not(layer2_outputs(1978));
    layer3_outputs(1029) <= layer2_outputs(2143);
    layer3_outputs(1030) <= not((layer2_outputs(1900)) and (layer2_outputs(399)));
    layer3_outputs(1031) <= layer2_outputs(2066);
    layer3_outputs(1032) <= '1';
    layer3_outputs(1033) <= not(layer2_outputs(1492)) or (layer2_outputs(1601));
    layer3_outputs(1034) <= not(layer2_outputs(432));
    layer3_outputs(1035) <= not((layer2_outputs(483)) and (layer2_outputs(472)));
    layer3_outputs(1036) <= (layer2_outputs(2124)) and (layer2_outputs(1231));
    layer3_outputs(1037) <= not(layer2_outputs(519)) or (layer2_outputs(1265));
    layer3_outputs(1038) <= not(layer2_outputs(961)) or (layer2_outputs(1763));
    layer3_outputs(1039) <= not((layer2_outputs(1887)) xor (layer2_outputs(1420)));
    layer3_outputs(1040) <= not(layer2_outputs(2409));
    layer3_outputs(1041) <= layer2_outputs(871);
    layer3_outputs(1042) <= '0';
    layer3_outputs(1043) <= not(layer2_outputs(2306));
    layer3_outputs(1044) <= not(layer2_outputs(1199));
    layer3_outputs(1045) <= layer2_outputs(1484);
    layer3_outputs(1046) <= (layer2_outputs(2441)) and not (layer2_outputs(892));
    layer3_outputs(1047) <= '0';
    layer3_outputs(1048) <= not((layer2_outputs(296)) or (layer2_outputs(477)));
    layer3_outputs(1049) <= not(layer2_outputs(1470));
    layer3_outputs(1050) <= not(layer2_outputs(395)) or (layer2_outputs(1890));
    layer3_outputs(1051) <= not(layer2_outputs(1698)) or (layer2_outputs(598));
    layer3_outputs(1052) <= not(layer2_outputs(1690));
    layer3_outputs(1053) <= not((layer2_outputs(291)) and (layer2_outputs(567)));
    layer3_outputs(1054) <= '1';
    layer3_outputs(1055) <= (layer2_outputs(715)) xor (layer2_outputs(1597));
    layer3_outputs(1056) <= (layer2_outputs(431)) and (layer2_outputs(2305));
    layer3_outputs(1057) <= not(layer2_outputs(746));
    layer3_outputs(1058) <= '0';
    layer3_outputs(1059) <= not(layer2_outputs(2267)) or (layer2_outputs(167));
    layer3_outputs(1060) <= '0';
    layer3_outputs(1061) <= (layer2_outputs(647)) and not (layer2_outputs(2308));
    layer3_outputs(1062) <= (layer2_outputs(1209)) and not (layer2_outputs(288));
    layer3_outputs(1063) <= not(layer2_outputs(1646));
    layer3_outputs(1064) <= '0';
    layer3_outputs(1065) <= (layer2_outputs(1189)) and not (layer2_outputs(587));
    layer3_outputs(1066) <= not(layer2_outputs(2428)) or (layer2_outputs(2047));
    layer3_outputs(1067) <= layer2_outputs(2189);
    layer3_outputs(1068) <= not(layer2_outputs(2353)) or (layer2_outputs(247));
    layer3_outputs(1069) <= (layer2_outputs(2263)) and not (layer2_outputs(2430));
    layer3_outputs(1070) <= '1';
    layer3_outputs(1071) <= (layer2_outputs(2408)) and not (layer2_outputs(515));
    layer3_outputs(1072) <= '0';
    layer3_outputs(1073) <= layer2_outputs(50);
    layer3_outputs(1074) <= layer2_outputs(536);
    layer3_outputs(1075) <= layer2_outputs(263);
    layer3_outputs(1076) <= not(layer2_outputs(1774));
    layer3_outputs(1077) <= '0';
    layer3_outputs(1078) <= not(layer2_outputs(114)) or (layer2_outputs(1061));
    layer3_outputs(1079) <= (layer2_outputs(1177)) and not (layer2_outputs(1402));
    layer3_outputs(1080) <= '0';
    layer3_outputs(1081) <= (layer2_outputs(1455)) or (layer2_outputs(125));
    layer3_outputs(1082) <= not(layer2_outputs(1291));
    layer3_outputs(1083) <= (layer2_outputs(1684)) or (layer2_outputs(624));
    layer3_outputs(1084) <= not(layer2_outputs(883)) or (layer2_outputs(1205));
    layer3_outputs(1085) <= (layer2_outputs(460)) xor (layer2_outputs(1881));
    layer3_outputs(1086) <= not(layer2_outputs(816));
    layer3_outputs(1087) <= not(layer2_outputs(977)) or (layer2_outputs(2210));
    layer3_outputs(1088) <= layer2_outputs(1644);
    layer3_outputs(1089) <= not(layer2_outputs(1732)) or (layer2_outputs(2537));
    layer3_outputs(1090) <= not(layer2_outputs(2218));
    layer3_outputs(1091) <= not(layer2_outputs(1860)) or (layer2_outputs(333));
    layer3_outputs(1092) <= (layer2_outputs(1689)) or (layer2_outputs(2433));
    layer3_outputs(1093) <= not(layer2_outputs(1445));
    layer3_outputs(1094) <= '0';
    layer3_outputs(1095) <= layer2_outputs(907);
    layer3_outputs(1096) <= not((layer2_outputs(795)) xor (layer2_outputs(2362)));
    layer3_outputs(1097) <= layer2_outputs(332);
    layer3_outputs(1098) <= layer2_outputs(1504);
    layer3_outputs(1099) <= not(layer2_outputs(1311)) or (layer2_outputs(713));
    layer3_outputs(1100) <= (layer2_outputs(1535)) and not (layer2_outputs(1305));
    layer3_outputs(1101) <= not(layer2_outputs(662)) or (layer2_outputs(62));
    layer3_outputs(1102) <= not(layer2_outputs(685));
    layer3_outputs(1103) <= not(layer2_outputs(182)) or (layer2_outputs(1260));
    layer3_outputs(1104) <= layer2_outputs(27);
    layer3_outputs(1105) <= layer2_outputs(676);
    layer3_outputs(1106) <= (layer2_outputs(52)) and not (layer2_outputs(324));
    layer3_outputs(1107) <= (layer2_outputs(2477)) or (layer2_outputs(1656));
    layer3_outputs(1108) <= '1';
    layer3_outputs(1109) <= (layer2_outputs(109)) and not (layer2_outputs(223));
    layer3_outputs(1110) <= (layer2_outputs(726)) and not (layer2_outputs(37));
    layer3_outputs(1111) <= layer2_outputs(70);
    layer3_outputs(1112) <= '0';
    layer3_outputs(1113) <= (layer2_outputs(2217)) and not (layer2_outputs(742));
    layer3_outputs(1114) <= (layer2_outputs(1987)) and (layer2_outputs(262));
    layer3_outputs(1115) <= layer2_outputs(2446);
    layer3_outputs(1116) <= not(layer2_outputs(2368)) or (layer2_outputs(791));
    layer3_outputs(1117) <= (layer2_outputs(1781)) and not (layer2_outputs(490));
    layer3_outputs(1118) <= (layer2_outputs(533)) and not (layer2_outputs(962));
    layer3_outputs(1119) <= not((layer2_outputs(695)) and (layer2_outputs(2199)));
    layer3_outputs(1120) <= not((layer2_outputs(1042)) xor (layer2_outputs(721)));
    layer3_outputs(1121) <= (layer2_outputs(2128)) or (layer2_outputs(1918));
    layer3_outputs(1122) <= layer2_outputs(2042);
    layer3_outputs(1123) <= layer2_outputs(1867);
    layer3_outputs(1124) <= (layer2_outputs(342)) and not (layer2_outputs(2285));
    layer3_outputs(1125) <= (layer2_outputs(749)) or (layer2_outputs(933));
    layer3_outputs(1126) <= '0';
    layer3_outputs(1127) <= (layer2_outputs(1508)) and not (layer2_outputs(491));
    layer3_outputs(1128) <= not(layer2_outputs(1309));
    layer3_outputs(1129) <= not(layer2_outputs(1844));
    layer3_outputs(1130) <= not(layer2_outputs(791)) or (layer2_outputs(308));
    layer3_outputs(1131) <= layer2_outputs(1618);
    layer3_outputs(1132) <= not((layer2_outputs(1462)) or (layer2_outputs(1961)));
    layer3_outputs(1133) <= (layer2_outputs(2197)) and not (layer2_outputs(1188));
    layer3_outputs(1134) <= '1';
    layer3_outputs(1135) <= not(layer2_outputs(812));
    layer3_outputs(1136) <= not((layer2_outputs(2147)) or (layer2_outputs(2167)));
    layer3_outputs(1137) <= not(layer2_outputs(2226));
    layer3_outputs(1138) <= (layer2_outputs(2513)) or (layer2_outputs(1221));
    layer3_outputs(1139) <= '0';
    layer3_outputs(1140) <= (layer2_outputs(2182)) and (layer2_outputs(330));
    layer3_outputs(1141) <= (layer2_outputs(1543)) and (layer2_outputs(2511));
    layer3_outputs(1142) <= '1';
    layer3_outputs(1143) <= not(layer2_outputs(737));
    layer3_outputs(1144) <= layer2_outputs(751);
    layer3_outputs(1145) <= layer2_outputs(60);
    layer3_outputs(1146) <= (layer2_outputs(971)) and not (layer2_outputs(1095));
    layer3_outputs(1147) <= layer2_outputs(1830);
    layer3_outputs(1148) <= not(layer2_outputs(774));
    layer3_outputs(1149) <= '1';
    layer3_outputs(1150) <= layer2_outputs(2342);
    layer3_outputs(1151) <= '1';
    layer3_outputs(1152) <= '0';
    layer3_outputs(1153) <= (layer2_outputs(1720)) and not (layer2_outputs(610));
    layer3_outputs(1154) <= not((layer2_outputs(1692)) or (layer2_outputs(19)));
    layer3_outputs(1155) <= not((layer2_outputs(1563)) or (layer2_outputs(1304)));
    layer3_outputs(1156) <= layer2_outputs(1851);
    layer3_outputs(1157) <= (layer2_outputs(688)) and not (layer2_outputs(817));
    layer3_outputs(1158) <= not(layer2_outputs(1551)) or (layer2_outputs(1185));
    layer3_outputs(1159) <= not(layer2_outputs(787)) or (layer2_outputs(1295));
    layer3_outputs(1160) <= (layer2_outputs(1596)) or (layer2_outputs(1591));
    layer3_outputs(1161) <= not((layer2_outputs(1987)) and (layer2_outputs(2175)));
    layer3_outputs(1162) <= layer2_outputs(1680);
    layer3_outputs(1163) <= layer2_outputs(26);
    layer3_outputs(1164) <= not(layer2_outputs(1225));
    layer3_outputs(1165) <= not(layer2_outputs(288));
    layer3_outputs(1166) <= layer2_outputs(924);
    layer3_outputs(1167) <= (layer2_outputs(1528)) and not (layer2_outputs(2463));
    layer3_outputs(1168) <= (layer2_outputs(101)) or (layer2_outputs(1218));
    layer3_outputs(1169) <= layer2_outputs(2093);
    layer3_outputs(1170) <= not(layer2_outputs(2553));
    layer3_outputs(1171) <= not(layer2_outputs(643)) or (layer2_outputs(2062));
    layer3_outputs(1172) <= layer2_outputs(934);
    layer3_outputs(1173) <= (layer2_outputs(942)) and not (layer2_outputs(1789));
    layer3_outputs(1174) <= '1';
    layer3_outputs(1175) <= layer2_outputs(537);
    layer3_outputs(1176) <= not(layer2_outputs(2449)) or (layer2_outputs(403));
    layer3_outputs(1177) <= not(layer2_outputs(1770)) or (layer2_outputs(753));
    layer3_outputs(1178) <= (layer2_outputs(1716)) or (layer2_outputs(731));
    layer3_outputs(1179) <= not(layer2_outputs(1425)) or (layer2_outputs(1917));
    layer3_outputs(1180) <= not(layer2_outputs(239)) or (layer2_outputs(32));
    layer3_outputs(1181) <= (layer2_outputs(1481)) and not (layer2_outputs(1624));
    layer3_outputs(1182) <= not((layer2_outputs(642)) or (layer2_outputs(1526)));
    layer3_outputs(1183) <= layer2_outputs(361);
    layer3_outputs(1184) <= not((layer2_outputs(233)) or (layer2_outputs(1872)));
    layer3_outputs(1185) <= not((layer2_outputs(623)) or (layer2_outputs(856)));
    layer3_outputs(1186) <= '0';
    layer3_outputs(1187) <= '0';
    layer3_outputs(1188) <= not(layer2_outputs(2346)) or (layer2_outputs(1130));
    layer3_outputs(1189) <= not((layer2_outputs(1597)) and (layer2_outputs(1275)));
    layer3_outputs(1190) <= not((layer2_outputs(785)) and (layer2_outputs(1175)));
    layer3_outputs(1191) <= not(layer2_outputs(778));
    layer3_outputs(1192) <= layer2_outputs(1449);
    layer3_outputs(1193) <= not(layer2_outputs(743));
    layer3_outputs(1194) <= '0';
    layer3_outputs(1195) <= not((layer2_outputs(917)) xor (layer2_outputs(2152)));
    layer3_outputs(1196) <= (layer2_outputs(1395)) and (layer2_outputs(415));
    layer3_outputs(1197) <= not(layer2_outputs(2315));
    layer3_outputs(1198) <= not(layer2_outputs(974)) or (layer2_outputs(2043));
    layer3_outputs(1199) <= not((layer2_outputs(310)) or (layer2_outputs(144)));
    layer3_outputs(1200) <= not(layer2_outputs(768)) or (layer2_outputs(1642));
    layer3_outputs(1201) <= not(layer2_outputs(2206)) or (layer2_outputs(896));
    layer3_outputs(1202) <= not((layer2_outputs(674)) or (layer2_outputs(1378)));
    layer3_outputs(1203) <= not(layer2_outputs(97)) or (layer2_outputs(1348));
    layer3_outputs(1204) <= layer2_outputs(2185);
    layer3_outputs(1205) <= '1';
    layer3_outputs(1206) <= not(layer2_outputs(1033));
    layer3_outputs(1207) <= (layer2_outputs(1658)) xor (layer2_outputs(1932));
    layer3_outputs(1208) <= not(layer2_outputs(2309));
    layer3_outputs(1209) <= (layer2_outputs(2543)) and not (layer2_outputs(1213));
    layer3_outputs(1210) <= (layer2_outputs(2452)) and not (layer2_outputs(806));
    layer3_outputs(1211) <= (layer2_outputs(9)) and not (layer2_outputs(2023));
    layer3_outputs(1212) <= (layer2_outputs(1144)) or (layer2_outputs(1784));
    layer3_outputs(1213) <= (layer2_outputs(1478)) and not (layer2_outputs(904));
    layer3_outputs(1214) <= layer2_outputs(1517);
    layer3_outputs(1215) <= not(layer2_outputs(292));
    layer3_outputs(1216) <= not(layer2_outputs(807)) or (layer2_outputs(369));
    layer3_outputs(1217) <= (layer2_outputs(272)) and (layer2_outputs(18));
    layer3_outputs(1218) <= (layer2_outputs(969)) and (layer2_outputs(1143));
    layer3_outputs(1219) <= not((layer2_outputs(709)) xor (layer2_outputs(1418)));
    layer3_outputs(1220) <= not(layer2_outputs(1838));
    layer3_outputs(1221) <= not(layer2_outputs(1944));
    layer3_outputs(1222) <= layer2_outputs(1516);
    layer3_outputs(1223) <= not(layer2_outputs(760));
    layer3_outputs(1224) <= layer2_outputs(68);
    layer3_outputs(1225) <= not((layer2_outputs(63)) and (layer2_outputs(1199)));
    layer3_outputs(1226) <= (layer2_outputs(1846)) or (layer2_outputs(646));
    layer3_outputs(1227) <= layer2_outputs(1760);
    layer3_outputs(1228) <= (layer2_outputs(2470)) or (layer2_outputs(2401));
    layer3_outputs(1229) <= '1';
    layer3_outputs(1230) <= (layer2_outputs(1685)) and not (layer2_outputs(2551));
    layer3_outputs(1231) <= (layer2_outputs(751)) or (layer2_outputs(1267));
    layer3_outputs(1232) <= not(layer2_outputs(467));
    layer3_outputs(1233) <= not(layer2_outputs(2131));
    layer3_outputs(1234) <= layer2_outputs(615);
    layer3_outputs(1235) <= (layer2_outputs(1311)) and not (layer2_outputs(1234));
    layer3_outputs(1236) <= layer2_outputs(828);
    layer3_outputs(1237) <= (layer2_outputs(458)) or (layer2_outputs(2507));
    layer3_outputs(1238) <= not((layer2_outputs(973)) or (layer2_outputs(1953)));
    layer3_outputs(1239) <= (layer2_outputs(262)) and not (layer2_outputs(2228));
    layer3_outputs(1240) <= '1';
    layer3_outputs(1241) <= (layer2_outputs(2100)) or (layer2_outputs(2030));
    layer3_outputs(1242) <= not(layer2_outputs(1687));
    layer3_outputs(1243) <= '1';
    layer3_outputs(1244) <= layer2_outputs(2434);
    layer3_outputs(1245) <= (layer2_outputs(162)) and (layer2_outputs(2122));
    layer3_outputs(1246) <= (layer2_outputs(459)) xor (layer2_outputs(493));
    layer3_outputs(1247) <= not(layer2_outputs(2074));
    layer3_outputs(1248) <= not((layer2_outputs(397)) and (layer2_outputs(878)));
    layer3_outputs(1249) <= (layer2_outputs(216)) and not (layer2_outputs(2080));
    layer3_outputs(1250) <= not((layer2_outputs(2345)) or (layer2_outputs(1381)));
    layer3_outputs(1251) <= not(layer2_outputs(1172));
    layer3_outputs(1252) <= '1';
    layer3_outputs(1253) <= (layer2_outputs(722)) and not (layer2_outputs(451));
    layer3_outputs(1254) <= (layer2_outputs(943)) xor (layer2_outputs(696));
    layer3_outputs(1255) <= layer2_outputs(2191);
    layer3_outputs(1256) <= not(layer2_outputs(278));
    layer3_outputs(1257) <= '1';
    layer3_outputs(1258) <= layer2_outputs(822);
    layer3_outputs(1259) <= '1';
    layer3_outputs(1260) <= not((layer2_outputs(1368)) or (layer2_outputs(44)));
    layer3_outputs(1261) <= layer2_outputs(257);
    layer3_outputs(1262) <= layer2_outputs(2194);
    layer3_outputs(1263) <= not(layer2_outputs(326));
    layer3_outputs(1264) <= layer2_outputs(2469);
    layer3_outputs(1265) <= not(layer2_outputs(1825));
    layer3_outputs(1266) <= (layer2_outputs(619)) and not (layer2_outputs(24));
    layer3_outputs(1267) <= not(layer2_outputs(1359)) or (layer2_outputs(2424));
    layer3_outputs(1268) <= (layer2_outputs(949)) and (layer2_outputs(1432));
    layer3_outputs(1269) <= layer2_outputs(1771);
    layer3_outputs(1270) <= '0';
    layer3_outputs(1271) <= not((layer2_outputs(2225)) and (layer2_outputs(2425)));
    layer3_outputs(1272) <= (layer2_outputs(2356)) and (layer2_outputs(130));
    layer3_outputs(1273) <= (layer2_outputs(1164)) and (layer2_outputs(378));
    layer3_outputs(1274) <= not((layer2_outputs(2350)) xor (layer2_outputs(564)));
    layer3_outputs(1275) <= (layer2_outputs(1401)) and not (layer2_outputs(551));
    layer3_outputs(1276) <= not(layer2_outputs(831));
    layer3_outputs(1277) <= not(layer2_outputs(2410)) or (layer2_outputs(2114));
    layer3_outputs(1278) <= not(layer2_outputs(847));
    layer3_outputs(1279) <= (layer2_outputs(2489)) and not (layer2_outputs(812));
    layer3_outputs(1280) <= not(layer2_outputs(49)) or (layer2_outputs(2205));
    layer3_outputs(1281) <= not(layer2_outputs(1776)) or (layer2_outputs(2141));
    layer3_outputs(1282) <= not((layer2_outputs(273)) and (layer2_outputs(2294)));
    layer3_outputs(1283) <= (layer2_outputs(309)) and (layer2_outputs(2082));
    layer3_outputs(1284) <= layer2_outputs(202);
    layer3_outputs(1285) <= not(layer2_outputs(1942)) or (layer2_outputs(138));
    layer3_outputs(1286) <= layer2_outputs(2396);
    layer3_outputs(1287) <= not((layer2_outputs(1632)) or (layer2_outputs(1197)));
    layer3_outputs(1288) <= (layer2_outputs(338)) and (layer2_outputs(1819));
    layer3_outputs(1289) <= (layer2_outputs(2018)) and not (layer2_outputs(1925));
    layer3_outputs(1290) <= (layer2_outputs(335)) and not (layer2_outputs(637));
    layer3_outputs(1291) <= '0';
    layer3_outputs(1292) <= not((layer2_outputs(1887)) and (layer2_outputs(1723)));
    layer3_outputs(1293) <= (layer2_outputs(1193)) and not (layer2_outputs(25));
    layer3_outputs(1294) <= layer2_outputs(728);
    layer3_outputs(1295) <= not((layer2_outputs(351)) and (layer2_outputs(51)));
    layer3_outputs(1296) <= layer2_outputs(2253);
    layer3_outputs(1297) <= layer2_outputs(693);
    layer3_outputs(1298) <= not(layer2_outputs(2078));
    layer3_outputs(1299) <= not(layer2_outputs(1557)) or (layer2_outputs(659));
    layer3_outputs(1300) <= (layer2_outputs(291)) and not (layer2_outputs(2219));
    layer3_outputs(1301) <= not(layer2_outputs(1822)) or (layer2_outputs(1896));
    layer3_outputs(1302) <= '0';
    layer3_outputs(1303) <= '0';
    layer3_outputs(1304) <= not((layer2_outputs(39)) xor (layer2_outputs(243)));
    layer3_outputs(1305) <= not((layer2_outputs(1276)) or (layer2_outputs(773)));
    layer3_outputs(1306) <= layer2_outputs(2139);
    layer3_outputs(1307) <= layer2_outputs(956);
    layer3_outputs(1308) <= not(layer2_outputs(2339)) or (layer2_outputs(1014));
    layer3_outputs(1309) <= (layer2_outputs(1865)) and not (layer2_outputs(75));
    layer3_outputs(1310) <= layer2_outputs(2152);
    layer3_outputs(1311) <= (layer2_outputs(1457)) and (layer2_outputs(1407));
    layer3_outputs(1312) <= layer2_outputs(1943);
    layer3_outputs(1313) <= (layer2_outputs(1662)) and (layer2_outputs(1962));
    layer3_outputs(1314) <= (layer2_outputs(382)) or (layer2_outputs(1003));
    layer3_outputs(1315) <= not(layer2_outputs(1128)) or (layer2_outputs(1009));
    layer3_outputs(1316) <= not(layer2_outputs(540));
    layer3_outputs(1317) <= not(layer2_outputs(1168));
    layer3_outputs(1318) <= not(layer2_outputs(284));
    layer3_outputs(1319) <= '0';
    layer3_outputs(1320) <= not((layer2_outputs(473)) and (layer2_outputs(537)));
    layer3_outputs(1321) <= layer2_outputs(2531);
    layer3_outputs(1322) <= '0';
    layer3_outputs(1323) <= not((layer2_outputs(2021)) or (layer2_outputs(2416)));
    layer3_outputs(1324) <= '0';
    layer3_outputs(1325) <= not((layer2_outputs(1079)) xor (layer2_outputs(2228)));
    layer3_outputs(1326) <= not(layer2_outputs(868));
    layer3_outputs(1327) <= layer2_outputs(1852);
    layer3_outputs(1328) <= layer2_outputs(1070);
    layer3_outputs(1329) <= not((layer2_outputs(481)) or (layer2_outputs(1162)));
    layer3_outputs(1330) <= layer2_outputs(2061);
    layer3_outputs(1331) <= (layer2_outputs(1945)) and not (layer2_outputs(2178));
    layer3_outputs(1332) <= not(layer2_outputs(2452)) or (layer2_outputs(2273));
    layer3_outputs(1333) <= '0';
    layer3_outputs(1334) <= layer2_outputs(1930);
    layer3_outputs(1335) <= not(layer2_outputs(2538)) or (layer2_outputs(2344));
    layer3_outputs(1336) <= (layer2_outputs(1504)) or (layer2_outputs(1854));
    layer3_outputs(1337) <= not(layer2_outputs(1365));
    layer3_outputs(1338) <= (layer2_outputs(1818)) or (layer2_outputs(391));
    layer3_outputs(1339) <= layer2_outputs(1336);
    layer3_outputs(1340) <= not((layer2_outputs(350)) or (layer2_outputs(125)));
    layer3_outputs(1341) <= not((layer2_outputs(196)) or (layer2_outputs(1383)));
    layer3_outputs(1342) <= not(layer2_outputs(1989));
    layer3_outputs(1343) <= '1';
    layer3_outputs(1344) <= (layer2_outputs(1943)) or (layer2_outputs(1814));
    layer3_outputs(1345) <= not(layer2_outputs(1372));
    layer3_outputs(1346) <= (layer2_outputs(2214)) xor (layer2_outputs(2268));
    layer3_outputs(1347) <= layer2_outputs(1174);
    layer3_outputs(1348) <= (layer2_outputs(430)) and (layer2_outputs(421));
    layer3_outputs(1349) <= (layer2_outputs(1430)) and (layer2_outputs(2038));
    layer3_outputs(1350) <= (layer2_outputs(276)) and not (layer2_outputs(432));
    layer3_outputs(1351) <= '1';
    layer3_outputs(1352) <= not(layer2_outputs(323));
    layer3_outputs(1353) <= (layer2_outputs(246)) and (layer2_outputs(1849));
    layer3_outputs(1354) <= not(layer2_outputs(1496));
    layer3_outputs(1355) <= (layer2_outputs(881)) and not (layer2_outputs(488));
    layer3_outputs(1356) <= not(layer2_outputs(100)) or (layer2_outputs(518));
    layer3_outputs(1357) <= not(layer2_outputs(877));
    layer3_outputs(1358) <= (layer2_outputs(2295)) xor (layer2_outputs(7));
    layer3_outputs(1359) <= '0';
    layer3_outputs(1360) <= '1';
    layer3_outputs(1361) <= '1';
    layer3_outputs(1362) <= layer2_outputs(131);
    layer3_outputs(1363) <= not(layer2_outputs(908));
    layer3_outputs(1364) <= (layer2_outputs(2508)) and not (layer2_outputs(149));
    layer3_outputs(1365) <= not((layer2_outputs(1974)) xor (layer2_outputs(118)));
    layer3_outputs(1366) <= not((layer2_outputs(1986)) or (layer2_outputs(2501)));
    layer3_outputs(1367) <= not((layer2_outputs(2149)) and (layer2_outputs(1520)));
    layer3_outputs(1368) <= not(layer2_outputs(1427)) or (layer2_outputs(42));
    layer3_outputs(1369) <= (layer2_outputs(2199)) and (layer2_outputs(953));
    layer3_outputs(1370) <= layer2_outputs(2522);
    layer3_outputs(1371) <= '1';
    layer3_outputs(1372) <= not(layer2_outputs(1039)) or (layer2_outputs(1282));
    layer3_outputs(1373) <= not(layer2_outputs(762));
    layer3_outputs(1374) <= '0';
    layer3_outputs(1375) <= '1';
    layer3_outputs(1376) <= '0';
    layer3_outputs(1377) <= not(layer2_outputs(2211));
    layer3_outputs(1378) <= layer2_outputs(779);
    layer3_outputs(1379) <= not((layer2_outputs(371)) and (layer2_outputs(1302)));
    layer3_outputs(1380) <= not(layer2_outputs(1793)) or (layer2_outputs(1256));
    layer3_outputs(1381) <= (layer2_outputs(470)) and not (layer2_outputs(1370));
    layer3_outputs(1382) <= not(layer2_outputs(205)) or (layer2_outputs(2051));
    layer3_outputs(1383) <= '1';
    layer3_outputs(1384) <= not(layer2_outputs(1709));
    layer3_outputs(1385) <= (layer2_outputs(2274)) and not (layer2_outputs(1583));
    layer3_outputs(1386) <= layer2_outputs(777);
    layer3_outputs(1387) <= layer2_outputs(1038);
    layer3_outputs(1388) <= (layer2_outputs(129)) xor (layer2_outputs(448));
    layer3_outputs(1389) <= (layer2_outputs(641)) and not (layer2_outputs(1897));
    layer3_outputs(1390) <= '0';
    layer3_outputs(1391) <= (layer2_outputs(652)) xor (layer2_outputs(2487));
    layer3_outputs(1392) <= not(layer2_outputs(499));
    layer3_outputs(1393) <= layer2_outputs(2474);
    layer3_outputs(1394) <= not(layer2_outputs(1223));
    layer3_outputs(1395) <= not(layer2_outputs(2472));
    layer3_outputs(1396) <= not(layer2_outputs(521)) or (layer2_outputs(1383));
    layer3_outputs(1397) <= (layer2_outputs(2407)) and not (layer2_outputs(2123));
    layer3_outputs(1398) <= layer2_outputs(1284);
    layer3_outputs(1399) <= (layer2_outputs(1446)) and not (layer2_outputs(19));
    layer3_outputs(1400) <= layer2_outputs(918);
    layer3_outputs(1401) <= layer2_outputs(384);
    layer3_outputs(1402) <= (layer2_outputs(1397)) and (layer2_outputs(1186));
    layer3_outputs(1403) <= '0';
    layer3_outputs(1404) <= not((layer2_outputs(1488)) and (layer2_outputs(453)));
    layer3_outputs(1405) <= not(layer2_outputs(1673));
    layer3_outputs(1406) <= (layer2_outputs(2240)) and not (layer2_outputs(1235));
    layer3_outputs(1407) <= not((layer2_outputs(928)) and (layer2_outputs(781)));
    layer3_outputs(1408) <= (layer2_outputs(1952)) and not (layer2_outputs(1714));
    layer3_outputs(1409) <= not(layer2_outputs(769)) or (layer2_outputs(59));
    layer3_outputs(1410) <= not(layer2_outputs(2098));
    layer3_outputs(1411) <= not(layer2_outputs(72)) or (layer2_outputs(1015));
    layer3_outputs(1412) <= not((layer2_outputs(1002)) or (layer2_outputs(952)));
    layer3_outputs(1413) <= not(layer2_outputs(1228)) or (layer2_outputs(1310));
    layer3_outputs(1414) <= not(layer2_outputs(936));
    layer3_outputs(1415) <= layer2_outputs(315);
    layer3_outputs(1416) <= '0';
    layer3_outputs(1417) <= (layer2_outputs(1423)) and not (layer2_outputs(972));
    layer3_outputs(1418) <= '0';
    layer3_outputs(1419) <= (layer2_outputs(1259)) and (layer2_outputs(439));
    layer3_outputs(1420) <= (layer2_outputs(2370)) or (layer2_outputs(196));
    layer3_outputs(1421) <= not((layer2_outputs(765)) or (layer2_outputs(1777)));
    layer3_outputs(1422) <= layer2_outputs(1559);
    layer3_outputs(1423) <= layer2_outputs(1950);
    layer3_outputs(1424) <= not(layer2_outputs(1801));
    layer3_outputs(1425) <= layer2_outputs(1586);
    layer3_outputs(1426) <= not((layer2_outputs(504)) or (layer2_outputs(360)));
    layer3_outputs(1427) <= not((layer2_outputs(2272)) or (layer2_outputs(436)));
    layer3_outputs(1428) <= not(layer2_outputs(1341)) or (layer2_outputs(1493));
    layer3_outputs(1429) <= '1';
    layer3_outputs(1430) <= '1';
    layer3_outputs(1431) <= layer2_outputs(938);
    layer3_outputs(1432) <= '0';
    layer3_outputs(1433) <= '0';
    layer3_outputs(1434) <= not(layer2_outputs(1783)) or (layer2_outputs(1980));
    layer3_outputs(1435) <= layer2_outputs(2394);
    layer3_outputs(1436) <= not(layer2_outputs(2393)) or (layer2_outputs(1838));
    layer3_outputs(1437) <= (layer2_outputs(443)) and not (layer2_outputs(1150));
    layer3_outputs(1438) <= layer2_outputs(1057);
    layer3_outputs(1439) <= (layer2_outputs(1860)) and not (layer2_outputs(2404));
    layer3_outputs(1440) <= (layer2_outputs(387)) and not (layer2_outputs(1329));
    layer3_outputs(1441) <= not(layer2_outputs(2163));
    layer3_outputs(1442) <= (layer2_outputs(1927)) or (layer2_outputs(456));
    layer3_outputs(1443) <= not(layer2_outputs(2265));
    layer3_outputs(1444) <= '0';
    layer3_outputs(1445) <= layer2_outputs(1361);
    layer3_outputs(1446) <= (layer2_outputs(606)) or (layer2_outputs(630));
    layer3_outputs(1447) <= not(layer2_outputs(1025)) or (layer2_outputs(2252));
    layer3_outputs(1448) <= (layer2_outputs(2340)) and (layer2_outputs(670));
    layer3_outputs(1449) <= not(layer2_outputs(2262));
    layer3_outputs(1450) <= (layer2_outputs(2260)) and not (layer2_outputs(445));
    layer3_outputs(1451) <= '0';
    layer3_outputs(1452) <= not((layer2_outputs(479)) and (layer2_outputs(2059)));
    layer3_outputs(1453) <= (layer2_outputs(1490)) or (layer2_outputs(306));
    layer3_outputs(1454) <= '1';
    layer3_outputs(1455) <= not(layer2_outputs(2071)) or (layer2_outputs(1759));
    layer3_outputs(1456) <= layer2_outputs(460);
    layer3_outputs(1457) <= not(layer2_outputs(227));
    layer3_outputs(1458) <= (layer2_outputs(991)) and not (layer2_outputs(1968));
    layer3_outputs(1459) <= not((layer2_outputs(12)) or (layer2_outputs(2464)));
    layer3_outputs(1460) <= not((layer2_outputs(1306)) or (layer2_outputs(1600)));
    layer3_outputs(1461) <= (layer2_outputs(2009)) and (layer2_outputs(1610));
    layer3_outputs(1462) <= layer2_outputs(1957);
    layer3_outputs(1463) <= layer2_outputs(1356);
    layer3_outputs(1464) <= layer2_outputs(2223);
    layer3_outputs(1465) <= (layer2_outputs(2257)) and not (layer2_outputs(2057));
    layer3_outputs(1466) <= (layer2_outputs(2358)) and not (layer2_outputs(1050));
    layer3_outputs(1467) <= layer2_outputs(1602);
    layer3_outputs(1468) <= (layer2_outputs(169)) and not (layer2_outputs(1564));
    layer3_outputs(1469) <= not(layer2_outputs(2118));
    layer3_outputs(1470) <= not((layer2_outputs(43)) or (layer2_outputs(726)));
    layer3_outputs(1471) <= not(layer2_outputs(57));
    layer3_outputs(1472) <= not(layer2_outputs(2390));
    layer3_outputs(1473) <= layer2_outputs(827);
    layer3_outputs(1474) <= not(layer2_outputs(1415));
    layer3_outputs(1475) <= layer2_outputs(1763);
    layer3_outputs(1476) <= layer2_outputs(2431);
    layer3_outputs(1477) <= layer2_outputs(926);
    layer3_outputs(1478) <= not(layer2_outputs(2490));
    layer3_outputs(1479) <= '0';
    layer3_outputs(1480) <= layer2_outputs(1361);
    layer3_outputs(1481) <= (layer2_outputs(1711)) and not (layer2_outputs(1828));
    layer3_outputs(1482) <= not(layer2_outputs(1861));
    layer3_outputs(1483) <= not(layer2_outputs(2471)) or (layer2_outputs(1412));
    layer3_outputs(1484) <= layer2_outputs(89);
    layer3_outputs(1485) <= not(layer2_outputs(493)) or (layer2_outputs(1780));
    layer3_outputs(1486) <= '0';
    layer3_outputs(1487) <= not(layer2_outputs(1640));
    layer3_outputs(1488) <= not(layer2_outputs(442)) or (layer2_outputs(480));
    layer3_outputs(1489) <= layer2_outputs(2014);
    layer3_outputs(1490) <= (layer2_outputs(1092)) or (layer2_outputs(422));
    layer3_outputs(1491) <= '1';
    layer3_outputs(1492) <= '0';
    layer3_outputs(1493) <= not(layer2_outputs(2042)) or (layer2_outputs(1889));
    layer3_outputs(1494) <= not((layer2_outputs(1008)) or (layer2_outputs(2341)));
    layer3_outputs(1495) <= (layer2_outputs(1275)) and not (layer2_outputs(1959));
    layer3_outputs(1496) <= not(layer2_outputs(2119)) or (layer2_outputs(1080));
    layer3_outputs(1497) <= '0';
    layer3_outputs(1498) <= '1';
    layer3_outputs(1499) <= layer2_outputs(1431);
    layer3_outputs(1500) <= not((layer2_outputs(2095)) and (layer2_outputs(1068)));
    layer3_outputs(1501) <= layer2_outputs(76);
    layer3_outputs(1502) <= '1';
    layer3_outputs(1503) <= (layer2_outputs(1180)) or (layer2_outputs(1963));
    layer3_outputs(1504) <= not(layer2_outputs(2484));
    layer3_outputs(1505) <= (layer2_outputs(242)) or (layer2_outputs(719));
    layer3_outputs(1506) <= '0';
    layer3_outputs(1507) <= not((layer2_outputs(2173)) and (layer2_outputs(105)));
    layer3_outputs(1508) <= not(layer2_outputs(755));
    layer3_outputs(1509) <= (layer2_outputs(918)) and not (layer2_outputs(447));
    layer3_outputs(1510) <= layer2_outputs(535);
    layer3_outputs(1511) <= not(layer2_outputs(1340));
    layer3_outputs(1512) <= '1';
    layer3_outputs(1513) <= layer2_outputs(1842);
    layer3_outputs(1514) <= layer2_outputs(1951);
    layer3_outputs(1515) <= (layer2_outputs(1030)) and not (layer2_outputs(941));
    layer3_outputs(1516) <= not(layer2_outputs(40));
    layer3_outputs(1517) <= (layer2_outputs(38)) or (layer2_outputs(1525));
    layer3_outputs(1518) <= (layer2_outputs(109)) and (layer2_outputs(1718));
    layer3_outputs(1519) <= layer2_outputs(1419);
    layer3_outputs(1520) <= layer2_outputs(815);
    layer3_outputs(1521) <= not((layer2_outputs(675)) and (layer2_outputs(487)));
    layer3_outputs(1522) <= not(layer2_outputs(1128)) or (layer2_outputs(1116));
    layer3_outputs(1523) <= not(layer2_outputs(2324)) or (layer2_outputs(1006));
    layer3_outputs(1524) <= layer2_outputs(904);
    layer3_outputs(1525) <= (layer2_outputs(1328)) xor (layer2_outputs(678));
    layer3_outputs(1526) <= (layer2_outputs(277)) or (layer2_outputs(885));
    layer3_outputs(1527) <= layer2_outputs(2269);
    layer3_outputs(1528) <= not(layer2_outputs(916));
    layer3_outputs(1529) <= (layer2_outputs(619)) and not (layer2_outputs(524));
    layer3_outputs(1530) <= not(layer2_outputs(385));
    layer3_outputs(1531) <= not(layer2_outputs(599)) or (layer2_outputs(2298));
    layer3_outputs(1532) <= not(layer2_outputs(972));
    layer3_outputs(1533) <= '0';
    layer3_outputs(1534) <= not(layer2_outputs(438));
    layer3_outputs(1535) <= not(layer2_outputs(1879));
    layer3_outputs(1536) <= not(layer2_outputs(1851));
    layer3_outputs(1537) <= not(layer2_outputs(1256));
    layer3_outputs(1538) <= (layer2_outputs(475)) and (layer2_outputs(1958));
    layer3_outputs(1539) <= (layer2_outputs(581)) and (layer2_outputs(2158));
    layer3_outputs(1540) <= (layer2_outputs(1598)) and not (layer2_outputs(1799));
    layer3_outputs(1541) <= not(layer2_outputs(1204));
    layer3_outputs(1542) <= not(layer2_outputs(272));
    layer3_outputs(1543) <= not(layer2_outputs(407)) or (layer2_outputs(1947));
    layer3_outputs(1544) <= layer2_outputs(898);
    layer3_outputs(1545) <= (layer2_outputs(2100)) and (layer2_outputs(640));
    layer3_outputs(1546) <= (layer2_outputs(546)) and not (layer2_outputs(2116));
    layer3_outputs(1547) <= '1';
    layer3_outputs(1548) <= not(layer2_outputs(113)) or (layer2_outputs(411));
    layer3_outputs(1549) <= '1';
    layer3_outputs(1550) <= layer2_outputs(41);
    layer3_outputs(1551) <= not((layer2_outputs(2451)) and (layer2_outputs(1021)));
    layer3_outputs(1552) <= not((layer2_outputs(1965)) and (layer2_outputs(2169)));
    layer3_outputs(1553) <= (layer2_outputs(1322)) and (layer2_outputs(364));
    layer3_outputs(1554) <= (layer2_outputs(1664)) and not (layer2_outputs(889));
    layer3_outputs(1555) <= (layer2_outputs(2335)) or (layer2_outputs(1723));
    layer3_outputs(1556) <= not(layer2_outputs(1376));
    layer3_outputs(1557) <= layer2_outputs(865);
    layer3_outputs(1558) <= not(layer2_outputs(658)) or (layer2_outputs(782));
    layer3_outputs(1559) <= not(layer2_outputs(1748));
    layer3_outputs(1560) <= '0';
    layer3_outputs(1561) <= (layer2_outputs(413)) and not (layer2_outputs(1503));
    layer3_outputs(1562) <= not(layer2_outputs(1082));
    layer3_outputs(1563) <= '0';
    layer3_outputs(1564) <= not(layer2_outputs(350)) or (layer2_outputs(2212));
    layer3_outputs(1565) <= not(layer2_outputs(2412));
    layer3_outputs(1566) <= '0';
    layer3_outputs(1567) <= layer2_outputs(1668);
    layer3_outputs(1568) <= layer2_outputs(891);
    layer3_outputs(1569) <= (layer2_outputs(417)) and (layer2_outputs(1324));
    layer3_outputs(1570) <= not((layer2_outputs(2200)) or (layer2_outputs(1352)));
    layer3_outputs(1571) <= not(layer2_outputs(2398));
    layer3_outputs(1572) <= not((layer2_outputs(83)) or (layer2_outputs(767)));
    layer3_outputs(1573) <= not(layer2_outputs(1706));
    layer3_outputs(1574) <= layer2_outputs(1089);
    layer3_outputs(1575) <= not(layer2_outputs(1783)) or (layer2_outputs(1377));
    layer3_outputs(1576) <= (layer2_outputs(340)) and not (layer2_outputs(525));
    layer3_outputs(1577) <= not(layer2_outputs(1472)) or (layer2_outputs(2390));
    layer3_outputs(1578) <= (layer2_outputs(261)) and not (layer2_outputs(1892));
    layer3_outputs(1579) <= (layer2_outputs(668)) and not (layer2_outputs(1447));
    layer3_outputs(1580) <= layer2_outputs(676);
    layer3_outputs(1581) <= layer2_outputs(1335);
    layer3_outputs(1582) <= (layer2_outputs(2090)) and not (layer2_outputs(2363));
    layer3_outputs(1583) <= not((layer2_outputs(1667)) xor (layer2_outputs(2421)));
    layer3_outputs(1584) <= layer2_outputs(2507);
    layer3_outputs(1585) <= (layer2_outputs(1893)) and not (layer2_outputs(1388));
    layer3_outputs(1586) <= (layer2_outputs(517)) and (layer2_outputs(1547));
    layer3_outputs(1587) <= not(layer2_outputs(1129));
    layer3_outputs(1588) <= not(layer2_outputs(96));
    layer3_outputs(1589) <= (layer2_outputs(1373)) or (layer2_outputs(213));
    layer3_outputs(1590) <= not(layer2_outputs(1247)) or (layer2_outputs(1810));
    layer3_outputs(1591) <= layer2_outputs(2225);
    layer3_outputs(1592) <= (layer2_outputs(1178)) and not (layer2_outputs(176));
    layer3_outputs(1593) <= (layer2_outputs(2378)) and (layer2_outputs(2018));
    layer3_outputs(1594) <= not((layer2_outputs(1438)) or (layer2_outputs(2424)));
    layer3_outputs(1595) <= not((layer2_outputs(1896)) xor (layer2_outputs(1404)));
    layer3_outputs(1596) <= not(layer2_outputs(1003)) or (layer2_outputs(877));
    layer3_outputs(1597) <= layer2_outputs(1745);
    layer3_outputs(1598) <= '1';
    layer3_outputs(1599) <= not(layer2_outputs(2177)) or (layer2_outputs(2005));
    layer3_outputs(1600) <= '0';
    layer3_outputs(1601) <= (layer2_outputs(90)) and not (layer2_outputs(285));
    layer3_outputs(1602) <= not(layer2_outputs(1612));
    layer3_outputs(1603) <= not(layer2_outputs(2502)) or (layer2_outputs(581));
    layer3_outputs(1604) <= (layer2_outputs(123)) and not (layer2_outputs(2483));
    layer3_outputs(1605) <= not(layer2_outputs(1605)) or (layer2_outputs(1805));
    layer3_outputs(1606) <= (layer2_outputs(2092)) and not (layer2_outputs(1049));
    layer3_outputs(1607) <= not(layer2_outputs(1293));
    layer3_outputs(1608) <= '0';
    layer3_outputs(1609) <= not(layer2_outputs(2285));
    layer3_outputs(1610) <= (layer2_outputs(153)) and not (layer2_outputs(1913));
    layer3_outputs(1611) <= not((layer2_outputs(2532)) or (layer2_outputs(1463)));
    layer3_outputs(1612) <= not(layer2_outputs(540)) or (layer2_outputs(1766));
    layer3_outputs(1613) <= (layer2_outputs(963)) or (layer2_outputs(197));
    layer3_outputs(1614) <= (layer2_outputs(1175)) and not (layer2_outputs(2545));
    layer3_outputs(1615) <= not((layer2_outputs(1862)) and (layer2_outputs(1111)));
    layer3_outputs(1616) <= layer2_outputs(465);
    layer3_outputs(1617) <= layer2_outputs(2000);
    layer3_outputs(1618) <= (layer2_outputs(890)) and (layer2_outputs(430));
    layer3_outputs(1619) <= '1';
    layer3_outputs(1620) <= layer2_outputs(2357);
    layer3_outputs(1621) <= not(layer2_outputs(405)) or (layer2_outputs(1562));
    layer3_outputs(1622) <= (layer2_outputs(1200)) and not (layer2_outputs(1609));
    layer3_outputs(1623) <= layer2_outputs(2417);
    layer3_outputs(1624) <= layer2_outputs(2323);
    layer3_outputs(1625) <= layer2_outputs(515);
    layer3_outputs(1626) <= layer2_outputs(53);
    layer3_outputs(1627) <= layer2_outputs(2348);
    layer3_outputs(1628) <= '1';
    layer3_outputs(1629) <= '1';
    layer3_outputs(1630) <= layer2_outputs(1065);
    layer3_outputs(1631) <= '1';
    layer3_outputs(1632) <= (layer2_outputs(1670)) and (layer2_outputs(586));
    layer3_outputs(1633) <= '0';
    layer3_outputs(1634) <= not(layer2_outputs(570)) or (layer2_outputs(1198));
    layer3_outputs(1635) <= not((layer2_outputs(1253)) and (layer2_outputs(2376)));
    layer3_outputs(1636) <= (layer2_outputs(1837)) and (layer2_outputs(1935));
    layer3_outputs(1637) <= not((layer2_outputs(2198)) or (layer2_outputs(1145)));
    layer3_outputs(1638) <= not((layer2_outputs(1006)) and (layer2_outputs(1119)));
    layer3_outputs(1639) <= '0';
    layer3_outputs(1640) <= not(layer2_outputs(567)) or (layer2_outputs(406));
    layer3_outputs(1641) <= '0';
    layer3_outputs(1642) <= (layer2_outputs(2251)) or (layer2_outputs(1750));
    layer3_outputs(1643) <= layer2_outputs(635);
    layer3_outputs(1644) <= not((layer2_outputs(2081)) xor (layer2_outputs(204)));
    layer3_outputs(1645) <= layer2_outputs(604);
    layer3_outputs(1646) <= (layer2_outputs(1227)) and (layer2_outputs(1865));
    layer3_outputs(1647) <= not((layer2_outputs(218)) and (layer2_outputs(942)));
    layer3_outputs(1648) <= not(layer2_outputs(1578)) or (layer2_outputs(1512));
    layer3_outputs(1649) <= '0';
    layer3_outputs(1650) <= (layer2_outputs(195)) and not (layer2_outputs(1461));
    layer3_outputs(1651) <= (layer2_outputs(1513)) xor (layer2_outputs(1910));
    layer3_outputs(1652) <= not(layer2_outputs(1989)) or (layer2_outputs(1788));
    layer3_outputs(1653) <= '0';
    layer3_outputs(1654) <= layer2_outputs(416);
    layer3_outputs(1655) <= not(layer2_outputs(120));
    layer3_outputs(1656) <= not(layer2_outputs(2504));
    layer3_outputs(1657) <= (layer2_outputs(1593)) and (layer2_outputs(267));
    layer3_outputs(1658) <= not(layer2_outputs(298)) or (layer2_outputs(1864));
    layer3_outputs(1659) <= not(layer2_outputs(1652));
    layer3_outputs(1660) <= not((layer2_outputs(1627)) and (layer2_outputs(649)));
    layer3_outputs(1661) <= not(layer2_outputs(455));
    layer3_outputs(1662) <= layer2_outputs(2024);
    layer3_outputs(1663) <= '0';
    layer3_outputs(1664) <= (layer2_outputs(503)) and (layer2_outputs(1321));
    layer3_outputs(1665) <= not(layer2_outputs(2114)) or (layer2_outputs(862));
    layer3_outputs(1666) <= not(layer2_outputs(969));
    layer3_outputs(1667) <= layer2_outputs(2544);
    layer3_outputs(1668) <= '0';
    layer3_outputs(1669) <= (layer2_outputs(689)) or (layer2_outputs(2375));
    layer3_outputs(1670) <= '0';
    layer3_outputs(1671) <= '0';
    layer3_outputs(1672) <= (layer2_outputs(1289)) and not (layer2_outputs(2343));
    layer3_outputs(1673) <= layer2_outputs(622);
    layer3_outputs(1674) <= layer2_outputs(2325);
    layer3_outputs(1675) <= (layer2_outputs(2013)) and not (layer2_outputs(236));
    layer3_outputs(1676) <= not(layer2_outputs(1219));
    layer3_outputs(1677) <= not(layer2_outputs(1572));
    layer3_outputs(1678) <= not((layer2_outputs(1737)) or (layer2_outputs(1462)));
    layer3_outputs(1679) <= not(layer2_outputs(1078));
    layer3_outputs(1680) <= layer2_outputs(2325);
    layer3_outputs(1681) <= '0';
    layer3_outputs(1682) <= '1';
    layer3_outputs(1683) <= layer2_outputs(164);
    layer3_outputs(1684) <= (layer2_outputs(1024)) and not (layer2_outputs(1110));
    layer3_outputs(1685) <= (layer2_outputs(2496)) or (layer2_outputs(1283));
    layer3_outputs(1686) <= (layer2_outputs(191)) and (layer2_outputs(2443));
    layer3_outputs(1687) <= not(layer2_outputs(2529));
    layer3_outputs(1688) <= not(layer2_outputs(2291));
    layer3_outputs(1689) <= not(layer2_outputs(2148)) or (layer2_outputs(1778));
    layer3_outputs(1690) <= not((layer2_outputs(1194)) or (layer2_outputs(1587)));
    layer3_outputs(1691) <= (layer2_outputs(325)) and not (layer2_outputs(1411));
    layer3_outputs(1692) <= not(layer2_outputs(1116));
    layer3_outputs(1693) <= (layer2_outputs(1762)) and not (layer2_outputs(2215));
    layer3_outputs(1694) <= (layer2_outputs(2467)) and (layer2_outputs(401));
    layer3_outputs(1695) <= (layer2_outputs(2393)) or (layer2_outputs(2139));
    layer3_outputs(1696) <= not(layer2_outputs(1533)) or (layer2_outputs(1144));
    layer3_outputs(1697) <= not(layer2_outputs(1129)) or (layer2_outputs(77));
    layer3_outputs(1698) <= (layer2_outputs(2039)) and (layer2_outputs(1603));
    layer3_outputs(1699) <= not(layer2_outputs(134)) or (layer2_outputs(2278));
    layer3_outputs(1700) <= not(layer2_outputs(2361));
    layer3_outputs(1701) <= not((layer2_outputs(2468)) or (layer2_outputs(1085)));
    layer3_outputs(1702) <= '0';
    layer3_outputs(1703) <= '0';
    layer3_outputs(1704) <= '0';
    layer3_outputs(1705) <= (layer2_outputs(924)) and not (layer2_outputs(597));
    layer3_outputs(1706) <= layer2_outputs(1554);
    layer3_outputs(1707) <= not((layer2_outputs(2404)) and (layer2_outputs(1094)));
    layer3_outputs(1708) <= not((layer2_outputs(1184)) and (layer2_outputs(1485)));
    layer3_outputs(1709) <= layer2_outputs(503);
    layer3_outputs(1710) <= (layer2_outputs(1140)) or (layer2_outputs(2552));
    layer3_outputs(1711) <= '1';
    layer3_outputs(1712) <= (layer2_outputs(2277)) and not (layer2_outputs(522));
    layer3_outputs(1713) <= (layer2_outputs(1849)) or (layer2_outputs(2436));
    layer3_outputs(1714) <= not(layer2_outputs(2097)) or (layer2_outputs(433));
    layer3_outputs(1715) <= layer2_outputs(318);
    layer3_outputs(1716) <= layer2_outputs(1093);
    layer3_outputs(1717) <= (layer2_outputs(435)) and not (layer2_outputs(1920));
    layer3_outputs(1718) <= (layer2_outputs(1880)) and (layer2_outputs(246));
    layer3_outputs(1719) <= not((layer2_outputs(264)) or (layer2_outputs(506)));
    layer3_outputs(1720) <= layer2_outputs(944);
    layer3_outputs(1721) <= '1';
    layer3_outputs(1722) <= not(layer2_outputs(1570));
    layer3_outputs(1723) <= not(layer2_outputs(41));
    layer3_outputs(1724) <= (layer2_outputs(787)) and (layer2_outputs(388));
    layer3_outputs(1725) <= (layer2_outputs(1629)) or (layer2_outputs(2494));
    layer3_outputs(1726) <= layer2_outputs(437);
    layer3_outputs(1727) <= not((layer2_outputs(1222)) and (layer2_outputs(1058)));
    layer3_outputs(1728) <= not(layer2_outputs(1804));
    layer3_outputs(1729) <= not((layer2_outputs(1938)) and (layer2_outputs(2405)));
    layer3_outputs(1730) <= layer2_outputs(1454);
    layer3_outputs(1731) <= not((layer2_outputs(55)) or (layer2_outputs(321)));
    layer3_outputs(1732) <= not((layer2_outputs(1399)) or (layer2_outputs(357)));
    layer3_outputs(1733) <= (layer2_outputs(669)) or (layer2_outputs(730));
    layer3_outputs(1734) <= not(layer2_outputs(2522));
    layer3_outputs(1735) <= '1';
    layer3_outputs(1736) <= '0';
    layer3_outputs(1737) <= '1';
    layer3_outputs(1738) <= not(layer2_outputs(991));
    layer3_outputs(1739) <= not(layer2_outputs(379));
    layer3_outputs(1740) <= not(layer2_outputs(440)) or (layer2_outputs(836));
    layer3_outputs(1741) <= (layer2_outputs(2321)) or (layer2_outputs(948));
    layer3_outputs(1742) <= not(layer2_outputs(900));
    layer3_outputs(1743) <= not((layer2_outputs(2515)) and (layer2_outputs(543)));
    layer3_outputs(1744) <= not(layer2_outputs(1740));
    layer3_outputs(1745) <= layer2_outputs(2292);
    layer3_outputs(1746) <= layer2_outputs(2313);
    layer3_outputs(1747) <= (layer2_outputs(2330)) or (layer2_outputs(1154));
    layer3_outputs(1748) <= not(layer2_outputs(2498));
    layer3_outputs(1749) <= not(layer2_outputs(353));
    layer3_outputs(1750) <= not(layer2_outputs(1734));
    layer3_outputs(1751) <= not(layer2_outputs(831));
    layer3_outputs(1752) <= not((layer2_outputs(937)) or (layer2_outputs(897)));
    layer3_outputs(1753) <= not(layer2_outputs(2279));
    layer3_outputs(1754) <= not(layer2_outputs(363)) or (layer2_outputs(2329));
    layer3_outputs(1755) <= (layer2_outputs(399)) and (layer2_outputs(1075));
    layer3_outputs(1756) <= (layer2_outputs(232)) or (layer2_outputs(1390));
    layer3_outputs(1757) <= (layer2_outputs(1954)) or (layer2_outputs(966));
    layer3_outputs(1758) <= not(layer2_outputs(1067));
    layer3_outputs(1759) <= not(layer2_outputs(2074)) or (layer2_outputs(576));
    layer3_outputs(1760) <= not(layer2_outputs(2438)) or (layer2_outputs(54));
    layer3_outputs(1761) <= not(layer2_outputs(1927));
    layer3_outputs(1762) <= not(layer2_outputs(2295)) or (layer2_outputs(1496));
    layer3_outputs(1763) <= '1';
    layer3_outputs(1764) <= not(layer2_outputs(1832));
    layer3_outputs(1765) <= not(layer2_outputs(1122));
    layer3_outputs(1766) <= not(layer2_outputs(2247)) or (layer2_outputs(931));
    layer3_outputs(1767) <= not((layer2_outputs(1929)) or (layer2_outputs(2517)));
    layer3_outputs(1768) <= (layer2_outputs(1359)) or (layer2_outputs(2436));
    layer3_outputs(1769) <= layer2_outputs(2088);
    layer3_outputs(1770) <= (layer2_outputs(2249)) and not (layer2_outputs(737));
    layer3_outputs(1771) <= not(layer2_outputs(2028)) or (layer2_outputs(2037));
    layer3_outputs(1772) <= layer2_outputs(644);
    layer3_outputs(1773) <= not((layer2_outputs(1831)) or (layer2_outputs(1044)));
    layer3_outputs(1774) <= (layer2_outputs(673)) and not (layer2_outputs(190));
    layer3_outputs(1775) <= not(layer2_outputs(1505)) or (layer2_outputs(2036));
    layer3_outputs(1776) <= (layer2_outputs(998)) and not (layer2_outputs(1485));
    layer3_outputs(1777) <= '1';
    layer3_outputs(1778) <= not(layer2_outputs(2258));
    layer3_outputs(1779) <= not(layer2_outputs(2302));
    layer3_outputs(1780) <= (layer2_outputs(2535)) and (layer2_outputs(2166));
    layer3_outputs(1781) <= not(layer2_outputs(2453));
    layer3_outputs(1782) <= layer2_outputs(165);
    layer3_outputs(1783) <= not(layer2_outputs(1878));
    layer3_outputs(1784) <= '0';
    layer3_outputs(1785) <= not(layer2_outputs(2195));
    layer3_outputs(1786) <= (layer2_outputs(53)) and not (layer2_outputs(292));
    layer3_outputs(1787) <= '0';
    layer3_outputs(1788) <= layer2_outputs(1137);
    layer3_outputs(1789) <= '1';
    layer3_outputs(1790) <= not(layer2_outputs(852));
    layer3_outputs(1791) <= not((layer2_outputs(2326)) or (layer2_outputs(1017)));
    layer3_outputs(1792) <= (layer2_outputs(2377)) and not (layer2_outputs(1645));
    layer3_outputs(1793) <= not(layer2_outputs(80)) or (layer2_outputs(2298));
    layer3_outputs(1794) <= (layer2_outputs(467)) and not (layer2_outputs(1936));
    layer3_outputs(1795) <= not(layer2_outputs(841));
    layer3_outputs(1796) <= not(layer2_outputs(702));
    layer3_outputs(1797) <= layer2_outputs(780);
    layer3_outputs(1798) <= not(layer2_outputs(983)) or (layer2_outputs(2451));
    layer3_outputs(1799) <= '0';
    layer3_outputs(1800) <= layer2_outputs(1806);
    layer3_outputs(1801) <= not(layer2_outputs(1827)) or (layer2_outputs(1590));
    layer3_outputs(1802) <= layer2_outputs(1794);
    layer3_outputs(1803) <= not(layer2_outputs(1990)) or (layer2_outputs(1233));
    layer3_outputs(1804) <= not(layer2_outputs(717));
    layer3_outputs(1805) <= layer2_outputs(1611);
    layer3_outputs(1806) <= layer2_outputs(1930);
    layer3_outputs(1807) <= '0';
    layer3_outputs(1808) <= not((layer2_outputs(2346)) or (layer2_outputs(1743)));
    layer3_outputs(1809) <= layer2_outputs(469);
    layer3_outputs(1810) <= not(layer2_outputs(1164)) or (layer2_outputs(1166));
    layer3_outputs(1811) <= '0';
    layer3_outputs(1812) <= not(layer2_outputs(2016));
    layer3_outputs(1813) <= '0';
    layer3_outputs(1814) <= not(layer2_outputs(1004));
    layer3_outputs(1815) <= not((layer2_outputs(160)) xor (layer2_outputs(694)));
    layer3_outputs(1816) <= not(layer2_outputs(1982));
    layer3_outputs(1817) <= not(layer2_outputs(1374));
    layer3_outputs(1818) <= not((layer2_outputs(1450)) or (layer2_outputs(95)));
    layer3_outputs(1819) <= not((layer2_outputs(645)) or (layer2_outputs(1107)));
    layer3_outputs(1820) <= not(layer2_outputs(1639));
    layer3_outputs(1821) <= (layer2_outputs(636)) and (layer2_outputs(681));
    layer3_outputs(1822) <= layer2_outputs(459);
    layer3_outputs(1823) <= not(layer2_outputs(1686)) or (layer2_outputs(1240));
    layer3_outputs(1824) <= '1';
    layer3_outputs(1825) <= layer2_outputs(121);
    layer3_outputs(1826) <= not((layer2_outputs(1654)) xor (layer2_outputs(571)));
    layer3_outputs(1827) <= '1';
    layer3_outputs(1828) <= layer2_outputs(719);
    layer3_outputs(1829) <= not(layer2_outputs(696)) or (layer2_outputs(17));
    layer3_outputs(1830) <= (layer2_outputs(960)) and not (layer2_outputs(1549));
    layer3_outputs(1831) <= layer2_outputs(2253);
    layer3_outputs(1832) <= not(layer2_outputs(1297)) or (layer2_outputs(994));
    layer3_outputs(1833) <= '0';
    layer3_outputs(1834) <= layer2_outputs(708);
    layer3_outputs(1835) <= not((layer2_outputs(1617)) and (layer2_outputs(1278)));
    layer3_outputs(1836) <= not((layer2_outputs(302)) or (layer2_outputs(1152)));
    layer3_outputs(1837) <= (layer2_outputs(130)) or (layer2_outputs(1109));
    layer3_outputs(1838) <= not(layer2_outputs(1654));
    layer3_outputs(1839) <= not(layer2_outputs(154));
    layer3_outputs(1840) <= not(layer2_outputs(1681));
    layer3_outputs(1841) <= layer2_outputs(85);
    layer3_outputs(1842) <= not(layer2_outputs(1319)) or (layer2_outputs(310));
    layer3_outputs(1843) <= layer2_outputs(595);
    layer3_outputs(1844) <= layer2_outputs(857);
    layer3_outputs(1845) <= layer2_outputs(1414);
    layer3_outputs(1846) <= (layer2_outputs(797)) and (layer2_outputs(2491));
    layer3_outputs(1847) <= layer2_outputs(147);
    layer3_outputs(1848) <= '0';
    layer3_outputs(1849) <= '1';
    layer3_outputs(1850) <= not(layer2_outputs(2455)) or (layer2_outputs(263));
    layer3_outputs(1851) <= '1';
    layer3_outputs(1852) <= (layer2_outputs(2118)) or (layer2_outputs(1920));
    layer3_outputs(1853) <= (layer2_outputs(56)) or (layer2_outputs(1173));
    layer3_outputs(1854) <= (layer2_outputs(2542)) xor (layer2_outputs(2214));
    layer3_outputs(1855) <= '1';
    layer3_outputs(1856) <= layer2_outputs(1626);
    layer3_outputs(1857) <= (layer2_outputs(2355)) and (layer2_outputs(16));
    layer3_outputs(1858) <= not(layer2_outputs(1824)) or (layer2_outputs(1982));
    layer3_outputs(1859) <= layer2_outputs(2181);
    layer3_outputs(1860) <= not((layer2_outputs(1954)) and (layer2_outputs(1977)));
    layer3_outputs(1861) <= (layer2_outputs(980)) and not (layer2_outputs(763));
    layer3_outputs(1862) <= not((layer2_outputs(2212)) xor (layer2_outputs(217)));
    layer3_outputs(1863) <= '0';
    layer3_outputs(1864) <= '0';
    layer3_outputs(1865) <= '1';
    layer3_outputs(1866) <= (layer2_outputs(2117)) and not (layer2_outputs(429));
    layer3_outputs(1867) <= not(layer2_outputs(45)) or (layer2_outputs(691));
    layer3_outputs(1868) <= not((layer2_outputs(2505)) and (layer2_outputs(2150)));
    layer3_outputs(1869) <= not((layer2_outputs(2241)) and (layer2_outputs(556)));
    layer3_outputs(1870) <= (layer2_outputs(978)) and not (layer2_outputs(1688));
    layer3_outputs(1871) <= not(layer2_outputs(1333)) or (layer2_outputs(2056));
    layer3_outputs(1872) <= layer2_outputs(2351);
    layer3_outputs(1873) <= not((layer2_outputs(1050)) and (layer2_outputs(135)));
    layer3_outputs(1874) <= (layer2_outputs(2520)) and not (layer2_outputs(1343));
    layer3_outputs(1875) <= '0';
    layer3_outputs(1876) <= '1';
    layer3_outputs(1877) <= '0';
    layer3_outputs(1878) <= (layer2_outputs(28)) and not (layer2_outputs(2426));
    layer3_outputs(1879) <= (layer2_outputs(1308)) and not (layer2_outputs(850));
    layer3_outputs(1880) <= (layer2_outputs(2309)) or (layer2_outputs(1913));
    layer3_outputs(1881) <= not(layer2_outputs(1300));
    layer3_outputs(1882) <= layer2_outputs(1408);
    layer3_outputs(1883) <= (layer2_outputs(698)) and not (layer2_outputs(1397));
    layer3_outputs(1884) <= (layer2_outputs(639)) and (layer2_outputs(1382));
    layer3_outputs(1885) <= '0';
    layer3_outputs(1886) <= '1';
    layer3_outputs(1887) <= (layer2_outputs(1824)) and not (layer2_outputs(1338));
    layer3_outputs(1888) <= not(layer2_outputs(1652)) or (layer2_outputs(1816));
    layer3_outputs(1889) <= (layer2_outputs(1106)) xor (layer2_outputs(1657));
    layer3_outputs(1890) <= '1';
    layer3_outputs(1891) <= layer2_outputs(382);
    layer3_outputs(1892) <= not(layer2_outputs(1729));
    layer3_outputs(1893) <= layer2_outputs(181);
    layer3_outputs(1894) <= not((layer2_outputs(1962)) or (layer2_outputs(1191)));
    layer3_outputs(1895) <= not(layer2_outputs(123));
    layer3_outputs(1896) <= not(layer2_outputs(1331));
    layer3_outputs(1897) <= (layer2_outputs(2438)) and not (layer2_outputs(1376));
    layer3_outputs(1898) <= not((layer2_outputs(539)) or (layer2_outputs(425)));
    layer3_outputs(1899) <= not(layer2_outputs(2420)) or (layer2_outputs(2200));
    layer3_outputs(1900) <= not(layer2_outputs(1420));
    layer3_outputs(1901) <= (layer2_outputs(1543)) and not (layer2_outputs(637));
    layer3_outputs(1902) <= not(layer2_outputs(1721));
    layer3_outputs(1903) <= (layer2_outputs(354)) and not (layer2_outputs(268));
    layer3_outputs(1904) <= (layer2_outputs(2411)) and (layer2_outputs(348));
    layer3_outputs(1905) <= not(layer2_outputs(718));
    layer3_outputs(1906) <= layer2_outputs(1946);
    layer3_outputs(1907) <= layer2_outputs(1232);
    layer3_outputs(1908) <= not((layer2_outputs(171)) and (layer2_outputs(1418)));
    layer3_outputs(1909) <= layer2_outputs(1802);
    layer3_outputs(1910) <= not(layer2_outputs(761)) or (layer2_outputs(874));
    layer3_outputs(1911) <= not(layer2_outputs(27));
    layer3_outputs(1912) <= not((layer2_outputs(2518)) xor (layer2_outputs(424)));
    layer3_outputs(1913) <= not(layer2_outputs(1020)) or (layer2_outputs(2303));
    layer3_outputs(1914) <= layer2_outputs(375);
    layer3_outputs(1915) <= layer2_outputs(570);
    layer3_outputs(1916) <= (layer2_outputs(1118)) or (layer2_outputs(1706));
    layer3_outputs(1917) <= (layer2_outputs(1867)) and not (layer2_outputs(1840));
    layer3_outputs(1918) <= layer2_outputs(2447);
    layer3_outputs(1919) <= not(layer2_outputs(402));
    layer3_outputs(1920) <= not(layer2_outputs(474)) or (layer2_outputs(1749));
    layer3_outputs(1921) <= (layer2_outputs(1724)) or (layer2_outputs(2402));
    layer3_outputs(1922) <= not(layer2_outputs(920)) or (layer2_outputs(1090));
    layer3_outputs(1923) <= not((layer2_outputs(2445)) or (layer2_outputs(1803)));
    layer3_outputs(1924) <= layer2_outputs(579);
    layer3_outputs(1925) <= (layer2_outputs(304)) and not (layer2_outputs(2210));
    layer3_outputs(1926) <= layer2_outputs(1969);
    layer3_outputs(1927) <= layer2_outputs(407);
    layer3_outputs(1928) <= layer2_outputs(428);
    layer3_outputs(1929) <= (layer2_outputs(2044)) xor (layer2_outputs(963));
    layer3_outputs(1930) <= layer2_outputs(1994);
    layer3_outputs(1931) <= not(layer2_outputs(738)) or (layer2_outputs(2483));
    layer3_outputs(1932) <= layer2_outputs(45);
    layer3_outputs(1933) <= not((layer2_outputs(2071)) and (layer2_outputs(466)));
    layer3_outputs(1934) <= not(layer2_outputs(1921));
    layer3_outputs(1935) <= '0';
    layer3_outputs(1936) <= (layer2_outputs(1672)) and not (layer2_outputs(1651));
    layer3_outputs(1937) <= '1';
    layer3_outputs(1938) <= not(layer2_outputs(684)) or (layer2_outputs(2414));
    layer3_outputs(1939) <= not(layer2_outputs(349));
    layer3_outputs(1940) <= (layer2_outputs(2328)) and not (layer2_outputs(1551));
    layer3_outputs(1941) <= not(layer2_outputs(811));
    layer3_outputs(1942) <= layer2_outputs(1553);
    layer3_outputs(1943) <= (layer2_outputs(953)) and not (layer2_outputs(616));
    layer3_outputs(1944) <= (layer2_outputs(2085)) and not (layer2_outputs(572));
    layer3_outputs(1945) <= not((layer2_outputs(2088)) or (layer2_outputs(677)));
    layer3_outputs(1946) <= (layer2_outputs(1208)) or (layer2_outputs(554));
    layer3_outputs(1947) <= not(layer2_outputs(4));
    layer3_outputs(1948) <= not(layer2_outputs(1238));
    layer3_outputs(1949) <= not(layer2_outputs(1498));
    layer3_outputs(1950) <= layer2_outputs(693);
    layer3_outputs(1951) <= (layer2_outputs(790)) and not (layer2_outputs(2024));
    layer3_outputs(1952) <= (layer2_outputs(2503)) and (layer2_outputs(211));
    layer3_outputs(1953) <= '1';
    layer3_outputs(1954) <= not(layer2_outputs(697));
    layer3_outputs(1955) <= layer2_outputs(809);
    layer3_outputs(1956) <= not((layer2_outputs(1353)) or (layer2_outputs(2369)));
    layer3_outputs(1957) <= layer2_outputs(1701);
    layer3_outputs(1958) <= not(layer2_outputs(962));
    layer3_outputs(1959) <= not(layer2_outputs(634));
    layer3_outputs(1960) <= (layer2_outputs(2542)) and not (layer2_outputs(1981));
    layer3_outputs(1961) <= not(layer2_outputs(323));
    layer3_outputs(1962) <= layer2_outputs(640);
    layer3_outputs(1963) <= not(layer2_outputs(2020));
    layer3_outputs(1964) <= layer2_outputs(1753);
    layer3_outputs(1965) <= (layer2_outputs(789)) and (layer2_outputs(1468));
    layer3_outputs(1966) <= not(layer2_outputs(2077)) or (layer2_outputs(2246));
    layer3_outputs(1967) <= layer2_outputs(2530);
    layer3_outputs(1968) <= not(layer2_outputs(1070));
    layer3_outputs(1969) <= (layer2_outputs(306)) and (layer2_outputs(1531));
    layer3_outputs(1970) <= layer2_outputs(778);
    layer3_outputs(1971) <= (layer2_outputs(1526)) and not (layer2_outputs(2310));
    layer3_outputs(1972) <= '1';
    layer3_outputs(1973) <= not(layer2_outputs(1268)) or (layer2_outputs(1267));
    layer3_outputs(1974) <= not(layer2_outputs(2288)) or (layer2_outputs(1287));
    layer3_outputs(1975) <= not((layer2_outputs(801)) xor (layer2_outputs(2206)));
    layer3_outputs(1976) <= layer2_outputs(2019);
    layer3_outputs(1977) <= (layer2_outputs(2065)) and not (layer2_outputs(1102));
    layer3_outputs(1978) <= layer2_outputs(2050);
    layer3_outputs(1979) <= (layer2_outputs(1054)) and (layer2_outputs(838));
    layer3_outputs(1980) <= layer2_outputs(336);
    layer3_outputs(1981) <= layer2_outputs(913);
    layer3_outputs(1982) <= (layer2_outputs(1007)) or (layer2_outputs(2009));
    layer3_outputs(1983) <= layer2_outputs(984);
    layer3_outputs(1984) <= (layer2_outputs(13)) or (layer2_outputs(2207));
    layer3_outputs(1985) <= not(layer2_outputs(1853));
    layer3_outputs(1986) <= '0';
    layer3_outputs(1987) <= layer2_outputs(1273);
    layer3_outputs(1988) <= layer2_outputs(1108);
    layer3_outputs(1989) <= (layer2_outputs(776)) and not (layer2_outputs(178));
    layer3_outputs(1990) <= not(layer2_outputs(2429));
    layer3_outputs(1991) <= not((layer2_outputs(1150)) and (layer2_outputs(271)));
    layer3_outputs(1992) <= '0';
    layer3_outputs(1993) <= not(layer2_outputs(1885));
    layer3_outputs(1994) <= '0';
    layer3_outputs(1995) <= not((layer2_outputs(1466)) and (layer2_outputs(1471)));
    layer3_outputs(1996) <= layer2_outputs(980);
    layer3_outputs(1997) <= not((layer2_outputs(1715)) and (layer2_outputs(808)));
    layer3_outputs(1998) <= '1';
    layer3_outputs(1999) <= (layer2_outputs(471)) or (layer2_outputs(2144));
    layer3_outputs(2000) <= layer2_outputs(621);
    layer3_outputs(2001) <= not((layer2_outputs(1957)) or (layer2_outputs(1513)));
    layer3_outputs(2002) <= not(layer2_outputs(546)) or (layer2_outputs(2439));
    layer3_outputs(2003) <= layer2_outputs(1207);
    layer3_outputs(2004) <= layer2_outputs(487);
    layer3_outputs(2005) <= (layer2_outputs(1781)) and (layer2_outputs(116));
    layer3_outputs(2006) <= (layer2_outputs(920)) or (layer2_outputs(641));
    layer3_outputs(2007) <= not(layer2_outputs(13)) or (layer2_outputs(88));
    layer3_outputs(2008) <= not((layer2_outputs(2158)) and (layer2_outputs(2512)));
    layer3_outputs(2009) <= not(layer2_outputs(380));
    layer3_outputs(2010) <= not(layer2_outputs(1332));
    layer3_outputs(2011) <= '0';
    layer3_outputs(2012) <= not((layer2_outputs(44)) or (layer2_outputs(76)));
    layer3_outputs(2013) <= layer2_outputs(1416);
    layer3_outputs(2014) <= not(layer2_outputs(1352));
    layer3_outputs(2015) <= not((layer2_outputs(301)) or (layer2_outputs(1473)));
    layer3_outputs(2016) <= (layer2_outputs(1438)) and not (layer2_outputs(126));
    layer3_outputs(2017) <= '0';
    layer3_outputs(2018) <= (layer2_outputs(1316)) and not (layer2_outputs(108));
    layer3_outputs(2019) <= (layer2_outputs(2257)) or (layer2_outputs(2550));
    layer3_outputs(2020) <= not((layer2_outputs(1281)) and (layer2_outputs(1580)));
    layer3_outputs(2021) <= not((layer2_outputs(585)) or (layer2_outputs(547)));
    layer3_outputs(2022) <= (layer2_outputs(191)) and (layer2_outputs(2273));
    layer3_outputs(2023) <= layer2_outputs(1448);
    layer3_outputs(2024) <= (layer2_outputs(1773)) and not (layer2_outputs(2550));
    layer3_outputs(2025) <= layer2_outputs(1079);
    layer3_outputs(2026) <= (layer2_outputs(757)) and not (layer2_outputs(862));
    layer3_outputs(2027) <= not(layer2_outputs(1238)) or (layer2_outputs(62));
    layer3_outputs(2028) <= not(layer2_outputs(1761));
    layer3_outputs(2029) <= not(layer2_outputs(142));
    layer3_outputs(2030) <= not((layer2_outputs(506)) or (layer2_outputs(1320)));
    layer3_outputs(2031) <= layer2_outputs(1902);
    layer3_outputs(2032) <= not(layer2_outputs(998));
    layer3_outputs(2033) <= layer2_outputs(519);
    layer3_outputs(2034) <= '1';
    layer3_outputs(2035) <= not(layer2_outputs(2440)) or (layer2_outputs(1210));
    layer3_outputs(2036) <= '0';
    layer3_outputs(2037) <= (layer2_outputs(1479)) and (layer2_outputs(198));
    layer3_outputs(2038) <= (layer2_outputs(573)) and not (layer2_outputs(1201));
    layer3_outputs(2039) <= layer2_outputs(2222);
    layer3_outputs(2040) <= layer2_outputs(2103);
    layer3_outputs(2041) <= not((layer2_outputs(829)) and (layer2_outputs(651)));
    layer3_outputs(2042) <= not(layer2_outputs(1897)) or (layer2_outputs(1820));
    layer3_outputs(2043) <= layer2_outputs(2090);
    layer3_outputs(2044) <= not(layer2_outputs(2101)) or (layer2_outputs(855));
    layer3_outputs(2045) <= (layer2_outputs(1660)) and not (layer2_outputs(2307));
    layer3_outputs(2046) <= (layer2_outputs(1074)) and not (layer2_outputs(533));
    layer3_outputs(2047) <= not(layer2_outputs(190));
    layer3_outputs(2048) <= (layer2_outputs(1716)) or (layer2_outputs(86));
    layer3_outputs(2049) <= not((layer2_outputs(1237)) xor (layer2_outputs(510)));
    layer3_outputs(2050) <= not((layer2_outputs(2387)) and (layer2_outputs(2547)));
    layer3_outputs(2051) <= not((layer2_outputs(1618)) or (layer2_outputs(811)));
    layer3_outputs(2052) <= not(layer2_outputs(2108)) or (layer2_outputs(245));
    layer3_outputs(2053) <= '0';
    layer3_outputs(2054) <= not(layer2_outputs(454)) or (layer2_outputs(308));
    layer3_outputs(2055) <= (layer2_outputs(2135)) and (layer2_outputs(1452));
    layer3_outputs(2056) <= not(layer2_outputs(416));
    layer3_outputs(2057) <= not(layer2_outputs(2433));
    layer3_outputs(2058) <= not((layer2_outputs(2320)) and (layer2_outputs(1063)));
    layer3_outputs(2059) <= '1';
    layer3_outputs(2060) <= layer2_outputs(1313);
    layer3_outputs(2061) <= not((layer2_outputs(853)) and (layer2_outputs(1015)));
    layer3_outputs(2062) <= (layer2_outputs(2491)) and not (layer2_outputs(78));
    layer3_outputs(2063) <= '0';
    layer3_outputs(2064) <= not(layer2_outputs(1180));
    layer3_outputs(2065) <= not((layer2_outputs(1966)) and (layer2_outputs(1375)));
    layer3_outputs(2066) <= not(layer2_outputs(1417));
    layer3_outputs(2067) <= not(layer2_outputs(484));
    layer3_outputs(2068) <= not(layer2_outputs(1892));
    layer3_outputs(2069) <= (layer2_outputs(656)) and not (layer2_outputs(1264));
    layer3_outputs(2070) <= '0';
    layer3_outputs(2071) <= not(layer2_outputs(685));
    layer3_outputs(2072) <= (layer2_outputs(1458)) and not (layer2_outputs(2530));
    layer3_outputs(2073) <= not(layer2_outputs(192));
    layer3_outputs(2074) <= layer2_outputs(1971);
    layer3_outputs(2075) <= '0';
    layer3_outputs(2076) <= (layer2_outputs(1350)) and (layer2_outputs(187));
    layer3_outputs(2077) <= '1';
    layer3_outputs(2078) <= not((layer2_outputs(2344)) or (layer2_outputs(669)));
    layer3_outputs(2079) <= (layer2_outputs(1276)) and not (layer2_outputs(894));
    layer3_outputs(2080) <= not(layer2_outputs(230));
    layer3_outputs(2081) <= layer2_outputs(1056);
    layer3_outputs(2082) <= (layer2_outputs(1748)) and not (layer2_outputs(1911));
    layer3_outputs(2083) <= (layer2_outputs(518)) or (layer2_outputs(2008));
    layer3_outputs(2084) <= not((layer2_outputs(1899)) or (layer2_outputs(58)));
    layer3_outputs(2085) <= (layer2_outputs(1081)) and not (layer2_outputs(1524));
    layer3_outputs(2086) <= not(layer2_outputs(1756)) or (layer2_outputs(2086));
    layer3_outputs(2087) <= layer2_outputs(49);
    layer3_outputs(2088) <= '1';
    layer3_outputs(2089) <= layer2_outputs(1159);
    layer3_outputs(2090) <= not((layer2_outputs(2115)) or (layer2_outputs(356)));
    layer3_outputs(2091) <= layer2_outputs(1273);
    layer3_outputs(2092) <= not((layer2_outputs(2105)) or (layer2_outputs(381)));
    layer3_outputs(2093) <= not((layer2_outputs(2252)) and (layer2_outputs(1695)));
    layer3_outputs(2094) <= '0';
    layer3_outputs(2095) <= not(layer2_outputs(1354)) or (layer2_outputs(2237));
    layer3_outputs(2096) <= (layer2_outputs(1360)) and not (layer2_outputs(856));
    layer3_outputs(2097) <= (layer2_outputs(2138)) xor (layer2_outputs(1595));
    layer3_outputs(2098) <= '1';
    layer3_outputs(2099) <= not((layer2_outputs(1986)) and (layer2_outputs(179)));
    layer3_outputs(2100) <= not(layer2_outputs(744));
    layer3_outputs(2101) <= layer2_outputs(492);
    layer3_outputs(2102) <= not(layer2_outputs(874));
    layer3_outputs(2103) <= not(layer2_outputs(1064));
    layer3_outputs(2104) <= (layer2_outputs(140)) and not (layer2_outputs(1077));
    layer3_outputs(2105) <= (layer2_outputs(2235)) and not (layer2_outputs(64));
    layer3_outputs(2106) <= (layer2_outputs(1679)) and not (layer2_outputs(1870));
    layer3_outputs(2107) <= (layer2_outputs(2470)) or (layer2_outputs(1789));
    layer3_outputs(2108) <= (layer2_outputs(2526)) or (layer2_outputs(1603));
    layer3_outputs(2109) <= (layer2_outputs(1715)) and (layer2_outputs(122));
    layer3_outputs(2110) <= (layer2_outputs(1682)) and (layer2_outputs(2549));
    layer3_outputs(2111) <= (layer2_outputs(2511)) and not (layer2_outputs(1572));
    layer3_outputs(2112) <= (layer2_outputs(2284)) and (layer2_outputs(455));
    layer3_outputs(2113) <= (layer2_outputs(678)) and (layer2_outputs(362));
    layer3_outputs(2114) <= (layer2_outputs(2441)) and (layer2_outputs(1476));
    layer3_outputs(2115) <= layer2_outputs(267);
    layer3_outputs(2116) <= (layer2_outputs(463)) and not (layer2_outputs(166));
    layer3_outputs(2117) <= (layer2_outputs(1873)) and not (layer2_outputs(1548));
    layer3_outputs(2118) <= '1';
    layer3_outputs(2119) <= (layer2_outputs(2094)) and (layer2_outputs(872));
    layer3_outputs(2120) <= '0';
    layer3_outputs(2121) <= layer2_outputs(1527);
    layer3_outputs(2122) <= layer2_outputs(2192);
    layer3_outputs(2123) <= '1';
    layer3_outputs(2124) <= layer2_outputs(1084);
    layer3_outputs(2125) <= (layer2_outputs(952)) and (layer2_outputs(1494));
    layer3_outputs(2126) <= (layer2_outputs(1209)) or (layer2_outputs(893));
    layer3_outputs(2127) <= '0';
    layer3_outputs(2128) <= (layer2_outputs(1398)) or (layer2_outputs(1661));
    layer3_outputs(2129) <= not((layer2_outputs(2398)) and (layer2_outputs(1348)));
    layer3_outputs(2130) <= not(layer2_outputs(206));
    layer3_outputs(2131) <= (layer2_outputs(512)) and not (layer2_outputs(331));
    layer3_outputs(2132) <= layer2_outputs(2031);
    layer3_outputs(2133) <= not((layer2_outputs(1215)) xor (layer2_outputs(2296)));
    layer3_outputs(2134) <= '0';
    layer3_outputs(2135) <= not(layer2_outputs(1635));
    layer3_outputs(2136) <= not((layer2_outputs(1580)) and (layer2_outputs(2148)));
    layer3_outputs(2137) <= (layer2_outputs(396)) and not (layer2_outputs(1248));
    layer3_outputs(2138) <= '1';
    layer3_outputs(2139) <= (layer2_outputs(1691)) and not (layer2_outputs(2495));
    layer3_outputs(2140) <= (layer2_outputs(851)) or (layer2_outputs(955));
    layer3_outputs(2141) <= not(layer2_outputs(2465));
    layer3_outputs(2142) <= (layer2_outputs(2485)) or (layer2_outputs(2174));
    layer3_outputs(2143) <= not(layer2_outputs(2036));
    layer3_outputs(2144) <= not(layer2_outputs(949)) or (layer2_outputs(1765));
    layer3_outputs(2145) <= (layer2_outputs(1141)) and not (layer2_outputs(30));
    layer3_outputs(2146) <= (layer2_outputs(993)) xor (layer2_outputs(1850));
    layer3_outputs(2147) <= '0';
    layer3_outputs(2148) <= (layer2_outputs(636)) and not (layer2_outputs(1370));
    layer3_outputs(2149) <= (layer2_outputs(1733)) and (layer2_outputs(1864));
    layer3_outputs(2150) <= not((layer2_outputs(1696)) and (layer2_outputs(1103)));
    layer3_outputs(2151) <= not(layer2_outputs(146)) or (layer2_outputs(721));
    layer3_outputs(2152) <= not((layer2_outputs(2548)) or (layer2_outputs(1835)));
    layer3_outputs(2153) <= layer2_outputs(1804);
    layer3_outputs(2154) <= (layer2_outputs(2111)) and (layer2_outputs(989));
    layer3_outputs(2155) <= layer2_outputs(1545);
    layer3_outputs(2156) <= not(layer2_outputs(699)) or (layer2_outputs(1391));
    layer3_outputs(2157) <= (layer2_outputs(1327)) or (layer2_outputs(1340));
    layer3_outputs(2158) <= (layer2_outputs(960)) and not (layer2_outputs(172));
    layer3_outputs(2159) <= layer2_outputs(1191);
    layer3_outputs(2160) <= '1';
    layer3_outputs(2161) <= (layer2_outputs(772)) and not (layer2_outputs(1392));
    layer3_outputs(2162) <= not(layer2_outputs(319)) or (layer2_outputs(2300));
    layer3_outputs(2163) <= not(layer2_outputs(415));
    layer3_outputs(2164) <= layer2_outputs(2473);
    layer3_outputs(2165) <= not(layer2_outputs(703)) or (layer2_outputs(2172));
    layer3_outputs(2166) <= not(layer2_outputs(2221));
    layer3_outputs(2167) <= '0';
    layer3_outputs(2168) <= '0';
    layer3_outputs(2169) <= '0';
    layer3_outputs(2170) <= not((layer2_outputs(1848)) xor (layer2_outputs(1362)));
    layer3_outputs(2171) <= (layer2_outputs(2509)) and not (layer2_outputs(2557));
    layer3_outputs(2172) <= not(layer2_outputs(2283)) or (layer2_outputs(1250));
    layer3_outputs(2173) <= layer2_outputs(2539);
    layer3_outputs(2174) <= not(layer2_outputs(1964));
    layer3_outputs(2175) <= (layer2_outputs(780)) or (layer2_outputs(2096));
    layer3_outputs(2176) <= not(layer2_outputs(1523)) or (layer2_outputs(496));
    layer3_outputs(2177) <= not(layer2_outputs(1941)) or (layer2_outputs(2126));
    layer3_outputs(2178) <= not(layer2_outputs(704)) or (layer2_outputs(1826));
    layer3_outputs(2179) <= (layer2_outputs(1895)) and (layer2_outputs(197));
    layer3_outputs(2180) <= (layer2_outputs(2374)) or (layer2_outputs(1722));
    layer3_outputs(2181) <= not(layer2_outputs(826));
    layer3_outputs(2182) <= layer2_outputs(591);
    layer3_outputs(2183) <= layer2_outputs(2082);
    layer3_outputs(2184) <= not(layer2_outputs(1692));
    layer3_outputs(2185) <= '0';
    layer3_outputs(2186) <= not(layer2_outputs(79)) or (layer2_outputs(279));
    layer3_outputs(2187) <= layer2_outputs(1012);
    layer3_outputs(2188) <= (layer2_outputs(840)) and not (layer2_outputs(711));
    layer3_outputs(2189) <= not((layer2_outputs(631)) or (layer2_outputs(1676)));
    layer3_outputs(2190) <= not((layer2_outputs(1991)) or (layer2_outputs(759)));
    layer3_outputs(2191) <= layer2_outputs(710);
    layer3_outputs(2192) <= '1';
    layer3_outputs(2193) <= '1';
    layer3_outputs(2194) <= (layer2_outputs(1937)) or (layer2_outputs(2033));
    layer3_outputs(2195) <= '1';
    layer3_outputs(2196) <= not(layer2_outputs(2400)) or (layer2_outputs(1678));
    layer3_outputs(2197) <= not(layer2_outputs(934));
    layer3_outputs(2198) <= not(layer2_outputs(1121));
    layer3_outputs(2199) <= layer2_outputs(1976);
    layer3_outputs(2200) <= '1';
    layer3_outputs(2201) <= not(layer2_outputs(837));
    layer3_outputs(2202) <= not(layer2_outputs(2430));
    layer3_outputs(2203) <= not(layer2_outputs(884));
    layer3_outputs(2204) <= (layer2_outputs(1333)) and (layer2_outputs(2364));
    layer3_outputs(2205) <= not(layer2_outputs(1309));
    layer3_outputs(2206) <= (layer2_outputs(824)) and (layer2_outputs(1141));
    layer3_outputs(2207) <= not(layer2_outputs(823));
    layer3_outputs(2208) <= not(layer2_outputs(1428)) or (layer2_outputs(2492));
    layer3_outputs(2209) <= not(layer2_outputs(2040));
    layer3_outputs(2210) <= (layer2_outputs(1702)) and not (layer2_outputs(2545));
    layer3_outputs(2211) <= not(layer2_outputs(2409)) or (layer2_outputs(369));
    layer3_outputs(2212) <= not((layer2_outputs(720)) xor (layer2_outputs(2032)));
    layer3_outputs(2213) <= layer2_outputs(1600);
    layer3_outputs(2214) <= not(layer2_outputs(2149));
    layer3_outputs(2215) <= not(layer2_outputs(1630)) or (layer2_outputs(1487));
    layer3_outputs(2216) <= '0';
    layer3_outputs(2217) <= not((layer2_outputs(729)) and (layer2_outputs(494)));
    layer3_outputs(2218) <= not(layer2_outputs(1145)) or (layer2_outputs(1390));
    layer3_outputs(2219) <= not(layer2_outputs(2405));
    layer3_outputs(2220) <= not(layer2_outputs(1698));
    layer3_outputs(2221) <= layer2_outputs(1403);
    layer3_outputs(2222) <= layer2_outputs(469);
    layer3_outputs(2223) <= (layer2_outputs(1786)) and (layer2_outputs(1226));
    layer3_outputs(2224) <= (layer2_outputs(2207)) and not (layer2_outputs(1364));
    layer3_outputs(2225) <= not(layer2_outputs(1828));
    layer3_outputs(2226) <= not(layer2_outputs(468));
    layer3_outputs(2227) <= layer2_outputs(1539);
    layer3_outputs(2228) <= not(layer2_outputs(814));
    layer3_outputs(2229) <= layer2_outputs(1362);
    layer3_outputs(2230) <= layer2_outputs(722);
    layer3_outputs(2231) <= layer2_outputs(120);
    layer3_outputs(2232) <= layer2_outputs(1724);
    layer3_outputs(2233) <= not(layer2_outputs(563)) or (layer2_outputs(1884));
    layer3_outputs(2234) <= (layer2_outputs(110)) or (layer2_outputs(286));
    layer3_outputs(2235) <= layer2_outputs(1236);
    layer3_outputs(2236) <= layer2_outputs(340);
    layer3_outputs(2237) <= (layer2_outputs(339)) and not (layer2_outputs(2130));
    layer3_outputs(2238) <= not(layer2_outputs(1520));
    layer3_outputs(2239) <= (layer2_outputs(1261)) and not (layer2_outputs(911));
    layer3_outputs(2240) <= not((layer2_outputs(1707)) and (layer2_outputs(1486)));
    layer3_outputs(2241) <= not(layer2_outputs(545)) or (layer2_outputs(686));
    layer3_outputs(2242) <= not(layer2_outputs(1705));
    layer3_outputs(2243) <= layer2_outputs(1035);
    layer3_outputs(2244) <= (layer2_outputs(1467)) and (layer2_outputs(968));
    layer3_outputs(2245) <= not(layer2_outputs(2448));
    layer3_outputs(2246) <= layer2_outputs(413);
    layer3_outputs(2247) <= layer2_outputs(1073);
    layer3_outputs(2248) <= layer2_outputs(1422);
    layer3_outputs(2249) <= layer2_outputs(113);
    layer3_outputs(2250) <= not(layer2_outputs(1877));
    layer3_outputs(2251) <= '1';
    layer3_outputs(2252) <= layer2_outputs(1436);
    layer3_outputs(2253) <= not(layer2_outputs(1833));
    layer3_outputs(2254) <= not(layer2_outputs(1174)) or (layer2_outputs(1542));
    layer3_outputs(2255) <= not((layer2_outputs(171)) xor (layer2_outputs(1847)));
    layer3_outputs(2256) <= layer2_outputs(183);
    layer3_outputs(2257) <= (layer2_outputs(900)) and not (layer2_outputs(1017));
    layer3_outputs(2258) <= '0';
    layer3_outputs(2259) <= (layer2_outputs(852)) and (layer2_outputs(2527));
    layer3_outputs(2260) <= not(layer2_outputs(1112));
    layer3_outputs(2261) <= not(layer2_outputs(101)) or (layer2_outputs(2559));
    layer3_outputs(2262) <= layer2_outputs(626);
    layer3_outputs(2263) <= not(layer2_outputs(557));
    layer3_outputs(2264) <= not(layer2_outputs(1517)) or (layer2_outputs(1794));
    layer3_outputs(2265) <= not(layer2_outputs(1051));
    layer3_outputs(2266) <= layer2_outputs(1589);
    layer3_outputs(2267) <= layer2_outputs(1541);
    layer3_outputs(2268) <= (layer2_outputs(464)) and not (layer2_outputs(1005));
    layer3_outputs(2269) <= layer2_outputs(2302);
    layer3_outputs(2270) <= '0';
    layer3_outputs(2271) <= (layer2_outputs(1351)) and (layer2_outputs(987));
    layer3_outputs(2272) <= (layer2_outputs(219)) or (layer2_outputs(2432));
    layer3_outputs(2273) <= not(layer2_outputs(1255)) or (layer2_outputs(235));
    layer3_outputs(2274) <= layer2_outputs(1820);
    layer3_outputs(2275) <= layer2_outputs(741);
    layer3_outputs(2276) <= (layer2_outputs(914)) and not (layer2_outputs(708));
    layer3_outputs(2277) <= not(layer2_outputs(2333));
    layer3_outputs(2278) <= '1';
    layer3_outputs(2279) <= (layer2_outputs(2286)) and not (layer2_outputs(3));
    layer3_outputs(2280) <= not(layer2_outputs(1836));
    layer3_outputs(2281) <= not((layer2_outputs(2113)) or (layer2_outputs(1745)));
    layer3_outputs(2282) <= layer2_outputs(2216);
    layer3_outputs(2283) <= (layer2_outputs(2167)) and (layer2_outputs(242));
    layer3_outputs(2284) <= (layer2_outputs(2032)) and not (layer2_outputs(1341));
    layer3_outputs(2285) <= (layer2_outputs(979)) and (layer2_outputs(1857));
    layer3_outputs(2286) <= layer2_outputs(1501);
    layer3_outputs(2287) <= not((layer2_outputs(1944)) and (layer2_outputs(48)));
    layer3_outputs(2288) <= (layer2_outputs(228)) and not (layer2_outputs(185));
    layer3_outputs(2289) <= (layer2_outputs(530)) and not (layer2_outputs(383));
    layer3_outputs(2290) <= (layer2_outputs(2376)) and not (layer2_outputs(971));
    layer3_outputs(2291) <= not((layer2_outputs(2204)) and (layer2_outputs(1985)));
    layer3_outputs(2292) <= not((layer2_outputs(2259)) and (layer2_outputs(1948)));
    layer3_outputs(2293) <= '1';
    layer3_outputs(2294) <= layer2_outputs(2046);
    layer3_outputs(2295) <= not(layer2_outputs(1701)) or (layer2_outputs(2029));
    layer3_outputs(2296) <= not(layer2_outputs(965)) or (layer2_outputs(1919));
    layer3_outputs(2297) <= not(layer2_outputs(1033)) or (layer2_outputs(2017));
    layer3_outputs(2298) <= (layer2_outputs(322)) and not (layer2_outputs(184));
    layer3_outputs(2299) <= not(layer2_outputs(418));
    layer3_outputs(2300) <= (layer2_outputs(1059)) or (layer2_outputs(914));
    layer3_outputs(2301) <= not(layer2_outputs(2005));
    layer3_outputs(2302) <= (layer2_outputs(295)) and (layer2_outputs(1653));
    layer3_outputs(2303) <= (layer2_outputs(758)) and not (layer2_outputs(2080));
    layer3_outputs(2304) <= (layer2_outputs(1369)) and not (layer2_outputs(497));
    layer3_outputs(2305) <= (layer2_outputs(937)) and not (layer2_outputs(1263));
    layer3_outputs(2306) <= (layer2_outputs(1906)) or (layer2_outputs(186));
    layer3_outputs(2307) <= not(layer2_outputs(2089)) or (layer2_outputs(2065));
    layer3_outputs(2308) <= layer2_outputs(374);
    layer3_outputs(2309) <= (layer2_outputs(2229)) and not (layer2_outputs(1686));
    layer3_outputs(2310) <= (layer2_outputs(1179)) xor (layer2_outputs(1011));
    layer3_outputs(2311) <= layer2_outputs(574);
    layer3_outputs(2312) <= (layer2_outputs(2510)) and not (layer2_outputs(1396));
    layer3_outputs(2313) <= layer2_outputs(2050);
    layer3_outputs(2314) <= (layer2_outputs(157)) and (layer2_outputs(1856));
    layer3_outputs(2315) <= not(layer2_outputs(2534));
    layer3_outputs(2316) <= layer2_outputs(813);
    layer3_outputs(2317) <= '0';
    layer3_outputs(2318) <= layer2_outputs(1579);
    layer3_outputs(2319) <= not(layer2_outputs(1304));
    layer3_outputs(2320) <= not(layer2_outputs(106)) or (layer2_outputs(1396));
    layer3_outputs(2321) <= not((layer2_outputs(368)) or (layer2_outputs(1833)));
    layer3_outputs(2322) <= '1';
    layer3_outputs(2323) <= layer2_outputs(2043);
    layer3_outputs(2324) <= not((layer2_outputs(35)) xor (layer2_outputs(1960)));
    layer3_outputs(2325) <= layer2_outputs(1536);
    layer3_outputs(2326) <= layer2_outputs(822);
    layer3_outputs(2327) <= (layer2_outputs(2052)) and not (layer2_outputs(244));
    layer3_outputs(2328) <= (layer2_outputs(1694)) or (layer2_outputs(706));
    layer3_outputs(2329) <= '1';
    layer3_outputs(2330) <= (layer2_outputs(213)) or (layer2_outputs(150));
    layer3_outputs(2331) <= (layer2_outputs(485)) and (layer2_outputs(34));
    layer3_outputs(2332) <= layer2_outputs(666);
    layer3_outputs(2333) <= '1';
    layer3_outputs(2334) <= not((layer2_outputs(1142)) or (layer2_outputs(279)));
    layer3_outputs(2335) <= not((layer2_outputs(229)) and (layer2_outputs(2446)));
    layer3_outputs(2336) <= layer2_outputs(1760);
    layer3_outputs(2337) <= not(layer2_outputs(1124));
    layer3_outputs(2338) <= layer2_outputs(2278);
    layer3_outputs(2339) <= not((layer2_outputs(1655)) and (layer2_outputs(617)));
    layer3_outputs(2340) <= not((layer2_outputs(591)) and (layer2_outputs(1288)));
    layer3_outputs(2341) <= not((layer2_outputs(821)) or (layer2_outputs(383)));
    layer3_outputs(2342) <= layer2_outputs(1665);
    layer3_outputs(2343) <= not((layer2_outputs(915)) and (layer2_outputs(1039)));
    layer3_outputs(2344) <= (layer2_outputs(613)) and (layer2_outputs(1761));
    layer3_outputs(2345) <= not(layer2_outputs(1034));
    layer3_outputs(2346) <= not(layer2_outputs(1047)) or (layer2_outputs(83));
    layer3_outputs(2347) <= not(layer2_outputs(226));
    layer3_outputs(2348) <= not(layer2_outputs(437)) or (layer2_outputs(2174));
    layer3_outputs(2349) <= layer2_outputs(221);
    layer3_outputs(2350) <= not((layer2_outputs(832)) xor (layer2_outputs(1974)));
    layer3_outputs(2351) <= not((layer2_outputs(1161)) xor (layer2_outputs(782)));
    layer3_outputs(2352) <= layer2_outputs(434);
    layer3_outputs(2353) <= '1';
    layer3_outputs(2354) <= layer2_outputs(959);
    layer3_outputs(2355) <= (layer2_outputs(733)) and (layer2_outputs(2448));
    layer3_outputs(2356) <= not(layer2_outputs(1098)) or (layer2_outputs(2327));
    layer3_outputs(2357) <= not(layer2_outputs(2010));
    layer3_outputs(2358) <= not((layer2_outputs(72)) xor (layer2_outputs(161)));
    layer3_outputs(2359) <= '0';
    layer3_outputs(2360) <= not(layer2_outputs(538)) or (layer2_outputs(535));
    layer3_outputs(2361) <= (layer2_outputs(333)) and not (layer2_outputs(1234));
    layer3_outputs(2362) <= '1';
    layer3_outputs(2363) <= not((layer2_outputs(2297)) or (layer2_outputs(2137)));
    layer3_outputs(2364) <= '0';
    layer3_outputs(2365) <= not(layer2_outputs(1295));
    layer3_outputs(2366) <= (layer2_outputs(2181)) and not (layer2_outputs(2055));
    layer3_outputs(2367) <= not(layer2_outputs(208));
    layer3_outputs(2368) <= not((layer2_outputs(1421)) and (layer2_outputs(1156)));
    layer3_outputs(2369) <= layer2_outputs(2319);
    layer3_outputs(2370) <= not(layer2_outputs(564)) or (layer2_outputs(2536));
    layer3_outputs(2371) <= (layer2_outputs(349)) and not (layer2_outputs(1966));
    layer3_outputs(2372) <= not(layer2_outputs(1107));
    layer3_outputs(2373) <= (layer2_outputs(2180)) and not (layer2_outputs(1123));
    layer3_outputs(2374) <= layer2_outputs(1409);
    layer3_outputs(2375) <= not(layer2_outputs(202));
    layer3_outputs(2376) <= layer2_outputs(644);
    layer3_outputs(2377) <= (layer2_outputs(2399)) and not (layer2_outputs(182));
    layer3_outputs(2378) <= (layer2_outputs(507)) and not (layer2_outputs(2055));
    layer3_outputs(2379) <= (layer2_outputs(2151)) or (layer2_outputs(1170));
    layer3_outputs(2380) <= not((layer2_outputs(1020)) and (layer2_outputs(826)));
    layer3_outputs(2381) <= not((layer2_outputs(2407)) and (layer2_outputs(2097)));
    layer3_outputs(2382) <= layer2_outputs(2234);
    layer3_outputs(2383) <= not((layer2_outputs(119)) or (layer2_outputs(1547)));
    layer3_outputs(2384) <= layer2_outputs(2311);
    layer3_outputs(2385) <= (layer2_outputs(1693)) and not (layer2_outputs(736));
    layer3_outputs(2386) <= layer2_outputs(898);
    layer3_outputs(2387) <= not(layer2_outputs(908)) or (layer2_outputs(1190));
    layer3_outputs(2388) <= layer2_outputs(2391);
    layer3_outputs(2389) <= layer2_outputs(713);
    layer3_outputs(2390) <= (layer2_outputs(1592)) and not (layer2_outputs(1522));
    layer3_outputs(2391) <= layer2_outputs(859);
    layer3_outputs(2392) <= not(layer2_outputs(2040));
    layer3_outputs(2393) <= (layer2_outputs(1018)) and not (layer2_outputs(91));
    layer3_outputs(2394) <= (layer2_outputs(2382)) or (layer2_outputs(1379));
    layer3_outputs(2395) <= not(layer2_outputs(69));
    layer3_outputs(2396) <= (layer2_outputs(2524)) or (layer2_outputs(412));
    layer3_outputs(2397) <= '0';
    layer3_outputs(2398) <= (layer2_outputs(1977)) and not (layer2_outputs(740));
    layer3_outputs(2399) <= not(layer2_outputs(337));
    layer3_outputs(2400) <= layer2_outputs(1792);
    layer3_outputs(2401) <= '0';
    layer3_outputs(2402) <= not(layer2_outputs(2480)) or (layer2_outputs(1813));
    layer3_outputs(2403) <= not(layer2_outputs(873));
    layer3_outputs(2404) <= layer2_outputs(1272);
    layer3_outputs(2405) <= '1';
    layer3_outputs(2406) <= (layer2_outputs(1038)) or (layer2_outputs(776));
    layer3_outputs(2407) <= layer2_outputs(1419);
    layer3_outputs(2408) <= not(layer2_outputs(1919));
    layer3_outputs(2409) <= (layer2_outputs(752)) and (layer2_outputs(1871));
    layer3_outputs(2410) <= not(layer2_outputs(1869)) or (layer2_outputs(75));
    layer3_outputs(2411) <= layer2_outputs(2372);
    layer3_outputs(2412) <= not(layer2_outputs(1013)) or (layer2_outputs(1138));
    layer3_outputs(2413) <= (layer2_outputs(1000)) and not (layer2_outputs(28));
    layer3_outputs(2414) <= (layer2_outputs(1658)) and not (layer2_outputs(2130));
    layer3_outputs(2415) <= (layer2_outputs(1916)) and not (layer2_outputs(880));
    layer3_outputs(2416) <= (layer2_outputs(1493)) or (layer2_outputs(2385));
    layer3_outputs(2417) <= (layer2_outputs(1758)) and (layer2_outputs(2247));
    layer3_outputs(2418) <= layer2_outputs(1075);
    layer3_outputs(2419) <= '1';
    layer3_outputs(2420) <= not(layer2_outputs(1519)) or (layer2_outputs(1606));
    layer3_outputs(2421) <= not(layer2_outputs(1672)) or (layer2_outputs(1247));
    layer3_outputs(2422) <= (layer2_outputs(215)) and not (layer2_outputs(1956));
    layer3_outputs(2423) <= layer2_outputs(568);
    layer3_outputs(2424) <= layer2_outputs(114);
    layer3_outputs(2425) <= '1';
    layer3_outputs(2426) <= not(layer2_outputs(609));
    layer3_outputs(2427) <= not((layer2_outputs(1467)) or (layer2_outputs(1501)));
    layer3_outputs(2428) <= layer2_outputs(2226);
    layer3_outputs(2429) <= (layer2_outputs(172)) and not (layer2_outputs(496));
    layer3_outputs(2430) <= (layer2_outputs(2338)) and not (layer2_outputs(1375));
    layer3_outputs(2431) <= (layer2_outputs(1968)) and (layer2_outputs(1928));
    layer3_outputs(2432) <= layer2_outputs(1013);
    layer3_outputs(2433) <= not(layer2_outputs(526));
    layer3_outputs(2434) <= (layer2_outputs(1002)) xor (layer2_outputs(1242));
    layer3_outputs(2435) <= '1';
    layer3_outputs(2436) <= not(layer2_outputs(997));
    layer3_outputs(2437) <= not(layer2_outputs(758));
    layer3_outputs(2438) <= not(layer2_outputs(2360)) or (layer2_outputs(2524));
    layer3_outputs(2439) <= layer2_outputs(2342);
    layer3_outputs(2440) <= not((layer2_outputs(87)) and (layer2_outputs(528)));
    layer3_outputs(2441) <= layer2_outputs(1062);
    layer3_outputs(2442) <= not(layer2_outputs(1465)) or (layer2_outputs(1157));
    layer3_outputs(2443) <= not(layer2_outputs(2220)) or (layer2_outputs(47));
    layer3_outputs(2444) <= (layer2_outputs(57)) and not (layer2_outputs(249));
    layer3_outputs(2445) <= not(layer2_outputs(1091));
    layer3_outputs(2446) <= not((layer2_outputs(1481)) or (layer2_outputs(143)));
    layer3_outputs(2447) <= not(layer2_outputs(1160));
    layer3_outputs(2448) <= layer2_outputs(88);
    layer3_outputs(2449) <= not(layer2_outputs(2092)) or (layer2_outputs(1800));
    layer3_outputs(2450) <= (layer2_outputs(1949)) and not (layer2_outputs(1584));
    layer3_outputs(2451) <= (layer2_outputs(1683)) or (layer2_outputs(2472));
    layer3_outputs(2452) <= layer2_outputs(1220);
    layer3_outputs(2453) <= '0';
    layer3_outputs(2454) <= layer2_outputs(1557);
    layer3_outputs(2455) <= not(layer2_outputs(1049));
    layer3_outputs(2456) <= (layer2_outputs(2501)) and (layer2_outputs(770));
    layer3_outputs(2457) <= not(layer2_outputs(2096));
    layer3_outputs(2458) <= not(layer2_outputs(338));
    layer3_outputs(2459) <= not((layer2_outputs(2066)) xor (layer2_outputs(1796)));
    layer3_outputs(2460) <= '1';
    layer3_outputs(2461) <= (layer2_outputs(1244)) xor (layer2_outputs(1762));
    layer3_outputs(2462) <= (layer2_outputs(1387)) and not (layer2_outputs(1518));
    layer3_outputs(2463) <= '1';
    layer3_outputs(2464) <= (layer2_outputs(1933)) or (layer2_outputs(1139));
    layer3_outputs(2465) <= (layer2_outputs(328)) and (layer2_outputs(1949));
    layer3_outputs(2466) <= (layer2_outputs(1808)) and not (layer2_outputs(1917));
    layer3_outputs(2467) <= (layer2_outputs(1742)) and not (layer2_outputs(2271));
    layer3_outputs(2468) <= (layer2_outputs(266)) and (layer2_outputs(1131));
    layer3_outputs(2469) <= (layer2_outputs(795)) or (layer2_outputs(10));
    layer3_outputs(2470) <= not(layer2_outputs(723));
    layer3_outputs(2471) <= not(layer2_outputs(1317));
    layer3_outputs(2472) <= '1';
    layer3_outputs(2473) <= not(layer2_outputs(1074));
    layer3_outputs(2474) <= layer2_outputs(2371);
    layer3_outputs(2475) <= layer2_outputs(1313);
    layer3_outputs(2476) <= layer2_outputs(756);
    layer3_outputs(2477) <= layer2_outputs(2014);
    layer3_outputs(2478) <= not(layer2_outputs(436)) or (layer2_outputs(1870));
    layer3_outputs(2479) <= '0';
    layer3_outputs(2480) <= not((layer2_outputs(2136)) or (layer2_outputs(1091)));
    layer3_outputs(2481) <= not(layer2_outputs(922));
    layer3_outputs(2482) <= layer2_outputs(367);
    layer3_outputs(2483) <= (layer2_outputs(240)) or (layer2_outputs(1643));
    layer3_outputs(2484) <= not(layer2_outputs(911)) or (layer2_outputs(56));
    layer3_outputs(2485) <= (layer2_outputs(1997)) and (layer2_outputs(1374));
    layer3_outputs(2486) <= (layer2_outputs(2367)) and (layer2_outputs(2103));
    layer3_outputs(2487) <= (layer2_outputs(738)) and not (layer2_outputs(373));
    layer3_outputs(2488) <= (layer2_outputs(2558)) and not (layer2_outputs(289));
    layer3_outputs(2489) <= (layer2_outputs(1669)) or (layer2_outputs(311));
    layer3_outputs(2490) <= not((layer2_outputs(1582)) or (layer2_outputs(36)));
    layer3_outputs(2491) <= (layer2_outputs(2449)) and not (layer2_outputs(611));
    layer3_outputs(2492) <= layer2_outputs(1777);
    layer3_outputs(2493) <= (layer2_outputs(1248)) or (layer2_outputs(2554));
    layer3_outputs(2494) <= layer2_outputs(188);
    layer3_outputs(2495) <= layer2_outputs(1690);
    layer3_outputs(2496) <= (layer2_outputs(425)) and not (layer2_outputs(243));
    layer3_outputs(2497) <= not(layer2_outputs(531));
    layer3_outputs(2498) <= (layer2_outputs(734)) and not (layer2_outputs(753));
    layer3_outputs(2499) <= (layer2_outputs(1212)) and not (layer2_outputs(1725));
    layer3_outputs(2500) <= (layer2_outputs(1314)) and not (layer2_outputs(2418));
    layer3_outputs(2501) <= not((layer2_outputs(179)) xor (layer2_outputs(2008)));
    layer3_outputs(2502) <= '1';
    layer3_outputs(2503) <= not(layer2_outputs(1451)) or (layer2_outputs(1358));
    layer3_outputs(2504) <= (layer2_outputs(613)) or (layer2_outputs(2348));
    layer3_outputs(2505) <= layer2_outputs(1055);
    layer3_outputs(2506) <= '0';
    layer3_outputs(2507) <= not((layer2_outputs(1279)) and (layer2_outputs(2136)));
    layer3_outputs(2508) <= '0';
    layer3_outputs(2509) <= not(layer2_outputs(785));
    layer3_outputs(2510) <= not(layer2_outputs(1604)) or (layer2_outputs(1515));
    layer3_outputs(2511) <= (layer2_outputs(1906)) and not (layer2_outputs(219));
    layer3_outputs(2512) <= (layer2_outputs(698)) and not (layer2_outputs(584));
    layer3_outputs(2513) <= not(layer2_outputs(1575)) or (layer2_outputs(745));
    layer3_outputs(2514) <= not(layer2_outputs(2020));
    layer3_outputs(2515) <= not((layer2_outputs(1844)) or (layer2_outputs(1183)));
    layer3_outputs(2516) <= (layer2_outputs(389)) and not (layer2_outputs(2460));
    layer3_outputs(2517) <= layer2_outputs(1195);
    layer3_outputs(2518) <= not(layer2_outputs(119)) or (layer2_outputs(867));
    layer3_outputs(2519) <= (layer2_outputs(1665)) xor (layer2_outputs(169));
    layer3_outputs(2520) <= '1';
    layer3_outputs(2521) <= '0';
    layer3_outputs(2522) <= not(layer2_outputs(1868)) or (layer2_outputs(50));
    layer3_outputs(2523) <= not(layer2_outputs(2203));
    layer3_outputs(2524) <= not(layer2_outputs(2294)) or (layer2_outputs(2345));
    layer3_outputs(2525) <= (layer2_outputs(1474)) and not (layer2_outputs(988));
    layer3_outputs(2526) <= not(layer2_outputs(1845));
    layer3_outputs(2527) <= layer2_outputs(2133);
    layer3_outputs(2528) <= not((layer2_outputs(2312)) and (layer2_outputs(1655)));
    layer3_outputs(2529) <= layer2_outputs(2079);
    layer3_outputs(2530) <= (layer2_outputs(2357)) and not (layer2_outputs(408));
    layer3_outputs(2531) <= not(layer2_outputs(2526)) or (layer2_outputs(2120));
    layer3_outputs(2532) <= '0';
    layer3_outputs(2533) <= not((layer2_outputs(133)) and (layer2_outputs(1)));
    layer3_outputs(2534) <= not(layer2_outputs(2078)) or (layer2_outputs(1197));
    layer3_outputs(2535) <= (layer2_outputs(238)) or (layer2_outputs(578));
    layer3_outputs(2536) <= (layer2_outputs(1403)) and not (layer2_outputs(534));
    layer3_outputs(2537) <= layer2_outputs(355);
    layer3_outputs(2538) <= (layer2_outputs(1585)) xor (layer2_outputs(441));
    layer3_outputs(2539) <= layer2_outputs(2289);
    layer3_outputs(2540) <= not(layer2_outputs(614));
    layer3_outputs(2541) <= not(layer2_outputs(92));
    layer3_outputs(2542) <= layer2_outputs(595);
    layer3_outputs(2543) <= (layer2_outputs(2322)) and (layer2_outputs(1612));
    layer3_outputs(2544) <= layer2_outputs(2378);
    layer3_outputs(2545) <= not(layer2_outputs(1492));
    layer3_outputs(2546) <= layer2_outputs(2315);
    layer3_outputs(2547) <= (layer2_outputs(547)) and not (layer2_outputs(280));
    layer3_outputs(2548) <= (layer2_outputs(801)) or (layer2_outputs(784));
    layer3_outputs(2549) <= layer2_outputs(1136);
    layer3_outputs(2550) <= layer2_outputs(511);
    layer3_outputs(2551) <= not((layer2_outputs(2354)) and (layer2_outputs(957)));
    layer3_outputs(2552) <= not(layer2_outputs(1151));
    layer3_outputs(2553) <= layer2_outputs(655);
    layer3_outputs(2554) <= layer2_outputs(746);
    layer3_outputs(2555) <= not((layer2_outputs(1752)) or (layer2_outputs(1232)));
    layer3_outputs(2556) <= not(layer2_outputs(1470));
    layer3_outputs(2557) <= not(layer2_outputs(0));
    layer3_outputs(2558) <= '1';
    layer3_outputs(2559) <= layer2_outputs(1712);
    layer4_outputs(0) <= not(layer3_outputs(266));
    layer4_outputs(1) <= not(layer3_outputs(1930)) or (layer3_outputs(2505));
    layer4_outputs(2) <= not(layer3_outputs(2525)) or (layer3_outputs(494));
    layer4_outputs(3) <= layer3_outputs(631);
    layer4_outputs(4) <= not(layer3_outputs(1299));
    layer4_outputs(5) <= (layer3_outputs(1985)) and not (layer3_outputs(1085));
    layer4_outputs(6) <= not((layer3_outputs(594)) xor (layer3_outputs(1164)));
    layer4_outputs(7) <= (layer3_outputs(1229)) and not (layer3_outputs(191));
    layer4_outputs(8) <= layer3_outputs(998);
    layer4_outputs(9) <= (layer3_outputs(1659)) and (layer3_outputs(1962));
    layer4_outputs(10) <= not((layer3_outputs(1853)) or (layer3_outputs(1855)));
    layer4_outputs(11) <= not(layer3_outputs(1933));
    layer4_outputs(12) <= layer3_outputs(735);
    layer4_outputs(13) <= (layer3_outputs(357)) or (layer3_outputs(2481));
    layer4_outputs(14) <= layer3_outputs(397);
    layer4_outputs(15) <= layer3_outputs(2493);
    layer4_outputs(16) <= '0';
    layer4_outputs(17) <= layer3_outputs(326);
    layer4_outputs(18) <= not(layer3_outputs(70));
    layer4_outputs(19) <= (layer3_outputs(150)) xor (layer3_outputs(1836));
    layer4_outputs(20) <= (layer3_outputs(2158)) or (layer3_outputs(61));
    layer4_outputs(21) <= not(layer3_outputs(2249));
    layer4_outputs(22) <= layer3_outputs(1595);
    layer4_outputs(23) <= layer3_outputs(2135);
    layer4_outputs(24) <= not(layer3_outputs(1011));
    layer4_outputs(25) <= not((layer3_outputs(1955)) and (layer3_outputs(327)));
    layer4_outputs(26) <= not((layer3_outputs(1114)) and (layer3_outputs(715)));
    layer4_outputs(27) <= not(layer3_outputs(1846)) or (layer3_outputs(1167));
    layer4_outputs(28) <= not(layer3_outputs(2238));
    layer4_outputs(29) <= not((layer3_outputs(2318)) and (layer3_outputs(2269)));
    layer4_outputs(30) <= '0';
    layer4_outputs(31) <= '1';
    layer4_outputs(32) <= (layer3_outputs(657)) xor (layer3_outputs(198));
    layer4_outputs(33) <= not(layer3_outputs(1788));
    layer4_outputs(34) <= not(layer3_outputs(2098));
    layer4_outputs(35) <= not(layer3_outputs(1747));
    layer4_outputs(36) <= '1';
    layer4_outputs(37) <= layer3_outputs(84);
    layer4_outputs(38) <= not(layer3_outputs(967));
    layer4_outputs(39) <= not((layer3_outputs(2504)) or (layer3_outputs(2241)));
    layer4_outputs(40) <= (layer3_outputs(1299)) and not (layer3_outputs(220));
    layer4_outputs(41) <= '1';
    layer4_outputs(42) <= not(layer3_outputs(1562));
    layer4_outputs(43) <= not(layer3_outputs(1298));
    layer4_outputs(44) <= not((layer3_outputs(2461)) xor (layer3_outputs(1789)));
    layer4_outputs(45) <= (layer3_outputs(1015)) or (layer3_outputs(445));
    layer4_outputs(46) <= not((layer3_outputs(636)) or (layer3_outputs(1804)));
    layer4_outputs(47) <= layer3_outputs(1345);
    layer4_outputs(48) <= '0';
    layer4_outputs(49) <= (layer3_outputs(1158)) xor (layer3_outputs(1127));
    layer4_outputs(50) <= layer3_outputs(1629);
    layer4_outputs(51) <= (layer3_outputs(659)) and (layer3_outputs(910));
    layer4_outputs(52) <= layer3_outputs(545);
    layer4_outputs(53) <= (layer3_outputs(1893)) xor (layer3_outputs(234));
    layer4_outputs(54) <= not(layer3_outputs(1753));
    layer4_outputs(55) <= (layer3_outputs(2174)) or (layer3_outputs(2129));
    layer4_outputs(56) <= (layer3_outputs(622)) and (layer3_outputs(2327));
    layer4_outputs(57) <= not((layer3_outputs(1694)) or (layer3_outputs(1870)));
    layer4_outputs(58) <= not(layer3_outputs(1737));
    layer4_outputs(59) <= '1';
    layer4_outputs(60) <= not(layer3_outputs(100));
    layer4_outputs(61) <= not((layer3_outputs(1290)) or (layer3_outputs(2130)));
    layer4_outputs(62) <= (layer3_outputs(2508)) and not (layer3_outputs(1808));
    layer4_outputs(63) <= layer3_outputs(1124);
    layer4_outputs(64) <= layer3_outputs(785);
    layer4_outputs(65) <= not(layer3_outputs(2282));
    layer4_outputs(66) <= layer3_outputs(1096);
    layer4_outputs(67) <= (layer3_outputs(1721)) or (layer3_outputs(518));
    layer4_outputs(68) <= not(layer3_outputs(969));
    layer4_outputs(69) <= '1';
    layer4_outputs(70) <= not(layer3_outputs(976));
    layer4_outputs(71) <= (layer3_outputs(78)) xor (layer3_outputs(12));
    layer4_outputs(72) <= (layer3_outputs(1752)) and not (layer3_outputs(1590));
    layer4_outputs(73) <= not((layer3_outputs(461)) and (layer3_outputs(737)));
    layer4_outputs(74) <= (layer3_outputs(1524)) xor (layer3_outputs(458));
    layer4_outputs(75) <= not(layer3_outputs(500));
    layer4_outputs(76) <= (layer3_outputs(1922)) xor (layer3_outputs(369));
    layer4_outputs(77) <= not(layer3_outputs(2367));
    layer4_outputs(78) <= (layer3_outputs(2140)) and (layer3_outputs(861));
    layer4_outputs(79) <= (layer3_outputs(585)) and not (layer3_outputs(1823));
    layer4_outputs(80) <= not(layer3_outputs(2542));
    layer4_outputs(81) <= layer3_outputs(1876);
    layer4_outputs(82) <= '1';
    layer4_outputs(83) <= layer3_outputs(1210);
    layer4_outputs(84) <= not(layer3_outputs(105));
    layer4_outputs(85) <= not((layer3_outputs(1794)) or (layer3_outputs(2395)));
    layer4_outputs(86) <= not((layer3_outputs(773)) and (layer3_outputs(1323)));
    layer4_outputs(87) <= layer3_outputs(2196);
    layer4_outputs(88) <= layer3_outputs(1680);
    layer4_outputs(89) <= not(layer3_outputs(2447)) or (layer3_outputs(1254));
    layer4_outputs(90) <= not(layer3_outputs(693));
    layer4_outputs(91) <= not(layer3_outputs(1924));
    layer4_outputs(92) <= not((layer3_outputs(1553)) or (layer3_outputs(978)));
    layer4_outputs(93) <= (layer3_outputs(857)) and not (layer3_outputs(1285));
    layer4_outputs(94) <= not(layer3_outputs(226)) or (layer3_outputs(2288));
    layer4_outputs(95) <= layer3_outputs(1786);
    layer4_outputs(96) <= (layer3_outputs(1688)) and not (layer3_outputs(1957));
    layer4_outputs(97) <= not(layer3_outputs(1097));
    layer4_outputs(98) <= '1';
    layer4_outputs(99) <= not(layer3_outputs(1195));
    layer4_outputs(100) <= not(layer3_outputs(1490));
    layer4_outputs(101) <= not(layer3_outputs(667));
    layer4_outputs(102) <= not(layer3_outputs(1026));
    layer4_outputs(103) <= (layer3_outputs(1943)) and (layer3_outputs(1337));
    layer4_outputs(104) <= not((layer3_outputs(1376)) and (layer3_outputs(1976)));
    layer4_outputs(105) <= layer3_outputs(941);
    layer4_outputs(106) <= layer3_outputs(2197);
    layer4_outputs(107) <= layer3_outputs(2457);
    layer4_outputs(108) <= not(layer3_outputs(1198));
    layer4_outputs(109) <= not(layer3_outputs(1832));
    layer4_outputs(110) <= layer3_outputs(1843);
    layer4_outputs(111) <= not(layer3_outputs(1707)) or (layer3_outputs(1129));
    layer4_outputs(112) <= (layer3_outputs(2202)) and not (layer3_outputs(1334));
    layer4_outputs(113) <= (layer3_outputs(401)) and (layer3_outputs(2201));
    layer4_outputs(114) <= not((layer3_outputs(2152)) and (layer3_outputs(1246)));
    layer4_outputs(115) <= (layer3_outputs(2347)) and not (layer3_outputs(447));
    layer4_outputs(116) <= not((layer3_outputs(1354)) or (layer3_outputs(770)));
    layer4_outputs(117) <= '1';
    layer4_outputs(118) <= layer3_outputs(2239);
    layer4_outputs(119) <= '1';
    layer4_outputs(120) <= not((layer3_outputs(421)) or (layer3_outputs(2200)));
    layer4_outputs(121) <= (layer3_outputs(763)) and not (layer3_outputs(438));
    layer4_outputs(122) <= layer3_outputs(468);
    layer4_outputs(123) <= not(layer3_outputs(1550));
    layer4_outputs(124) <= not(layer3_outputs(2468));
    layer4_outputs(125) <= not(layer3_outputs(1480));
    layer4_outputs(126) <= (layer3_outputs(634)) and not (layer3_outputs(1409));
    layer4_outputs(127) <= (layer3_outputs(154)) or (layer3_outputs(1424));
    layer4_outputs(128) <= '1';
    layer4_outputs(129) <= '0';
    layer4_outputs(130) <= (layer3_outputs(1776)) and not (layer3_outputs(1757));
    layer4_outputs(131) <= layer3_outputs(153);
    layer4_outputs(132) <= '0';
    layer4_outputs(133) <= not(layer3_outputs(1981));
    layer4_outputs(134) <= not(layer3_outputs(1284));
    layer4_outputs(135) <= layer3_outputs(97);
    layer4_outputs(136) <= not(layer3_outputs(2033));
    layer4_outputs(137) <= not(layer3_outputs(522));
    layer4_outputs(138) <= (layer3_outputs(1503)) and (layer3_outputs(2410));
    layer4_outputs(139) <= layer3_outputs(1135);
    layer4_outputs(140) <= not(layer3_outputs(2319));
    layer4_outputs(141) <= layer3_outputs(1170);
    layer4_outputs(142) <= layer3_outputs(184);
    layer4_outputs(143) <= (layer3_outputs(439)) and not (layer3_outputs(709));
    layer4_outputs(144) <= (layer3_outputs(915)) and not (layer3_outputs(367));
    layer4_outputs(145) <= not(layer3_outputs(209));
    layer4_outputs(146) <= not(layer3_outputs(1804));
    layer4_outputs(147) <= (layer3_outputs(2130)) and not (layer3_outputs(1879));
    layer4_outputs(148) <= not((layer3_outputs(656)) and (layer3_outputs(1129)));
    layer4_outputs(149) <= not((layer3_outputs(1275)) xor (layer3_outputs(874)));
    layer4_outputs(150) <= layer3_outputs(52);
    layer4_outputs(151) <= (layer3_outputs(670)) and (layer3_outputs(2061));
    layer4_outputs(152) <= not(layer3_outputs(943));
    layer4_outputs(153) <= '1';
    layer4_outputs(154) <= layer3_outputs(106);
    layer4_outputs(155) <= layer3_outputs(905);
    layer4_outputs(156) <= layer3_outputs(1041);
    layer4_outputs(157) <= (layer3_outputs(1112)) and not (layer3_outputs(2129));
    layer4_outputs(158) <= layer3_outputs(440);
    layer4_outputs(159) <= not(layer3_outputs(218));
    layer4_outputs(160) <= layer3_outputs(1997);
    layer4_outputs(161) <= layer3_outputs(1182);
    layer4_outputs(162) <= layer3_outputs(2421);
    layer4_outputs(163) <= not((layer3_outputs(275)) and (layer3_outputs(1821)));
    layer4_outputs(164) <= not(layer3_outputs(1594)) or (layer3_outputs(515));
    layer4_outputs(165) <= '0';
    layer4_outputs(166) <= not(layer3_outputs(2358));
    layer4_outputs(167) <= not(layer3_outputs(2428));
    layer4_outputs(168) <= not(layer3_outputs(478));
    layer4_outputs(169) <= layer3_outputs(1238);
    layer4_outputs(170) <= (layer3_outputs(1923)) and not (layer3_outputs(215));
    layer4_outputs(171) <= (layer3_outputs(982)) and not (layer3_outputs(851));
    layer4_outputs(172) <= '1';
    layer4_outputs(173) <= (layer3_outputs(2474)) and (layer3_outputs(750));
    layer4_outputs(174) <= layer3_outputs(719);
    layer4_outputs(175) <= (layer3_outputs(1451)) and (layer3_outputs(82));
    layer4_outputs(176) <= (layer3_outputs(2180)) and (layer3_outputs(2513));
    layer4_outputs(177) <= layer3_outputs(1819);
    layer4_outputs(178) <= (layer3_outputs(641)) and (layer3_outputs(519));
    layer4_outputs(179) <= not(layer3_outputs(1081)) or (layer3_outputs(1370));
    layer4_outputs(180) <= not(layer3_outputs(797));
    layer4_outputs(181) <= '0';
    layer4_outputs(182) <= layer3_outputs(2067);
    layer4_outputs(183) <= '0';
    layer4_outputs(184) <= (layer3_outputs(1858)) or (layer3_outputs(1282));
    layer4_outputs(185) <= not(layer3_outputs(1288)) or (layer3_outputs(2183));
    layer4_outputs(186) <= not(layer3_outputs(582));
    layer4_outputs(187) <= layer3_outputs(1463);
    layer4_outputs(188) <= layer3_outputs(1918);
    layer4_outputs(189) <= (layer3_outputs(1377)) or (layer3_outputs(41));
    layer4_outputs(190) <= not((layer3_outputs(2321)) and (layer3_outputs(1452)));
    layer4_outputs(191) <= not(layer3_outputs(246));
    layer4_outputs(192) <= not((layer3_outputs(75)) and (layer3_outputs(1733)));
    layer4_outputs(193) <= (layer3_outputs(943)) and not (layer3_outputs(625));
    layer4_outputs(194) <= (layer3_outputs(1853)) and (layer3_outputs(64));
    layer4_outputs(195) <= not((layer3_outputs(1075)) or (layer3_outputs(1655)));
    layer4_outputs(196) <= layer3_outputs(485);
    layer4_outputs(197) <= not(layer3_outputs(16)) or (layer3_outputs(8));
    layer4_outputs(198) <= not(layer3_outputs(1142)) or (layer3_outputs(1551));
    layer4_outputs(199) <= not(layer3_outputs(2158));
    layer4_outputs(200) <= (layer3_outputs(1632)) and not (layer3_outputs(944));
    layer4_outputs(201) <= layer3_outputs(1262);
    layer4_outputs(202) <= not(layer3_outputs(1413));
    layer4_outputs(203) <= '0';
    layer4_outputs(204) <= (layer3_outputs(1358)) and (layer3_outputs(1411));
    layer4_outputs(205) <= not(layer3_outputs(325));
    layer4_outputs(206) <= (layer3_outputs(232)) and (layer3_outputs(2417));
    layer4_outputs(207) <= layer3_outputs(2043);
    layer4_outputs(208) <= not(layer3_outputs(2218));
    layer4_outputs(209) <= not(layer3_outputs(166));
    layer4_outputs(210) <= layer3_outputs(2225);
    layer4_outputs(211) <= '0';
    layer4_outputs(212) <= '0';
    layer4_outputs(213) <= layer3_outputs(1585);
    layer4_outputs(214) <= (layer3_outputs(481)) and not (layer3_outputs(2284));
    layer4_outputs(215) <= (layer3_outputs(774)) or (layer3_outputs(1387));
    layer4_outputs(216) <= not(layer3_outputs(1592));
    layer4_outputs(217) <= layer3_outputs(545);
    layer4_outputs(218) <= not(layer3_outputs(2011)) or (layer3_outputs(1380));
    layer4_outputs(219) <= not(layer3_outputs(752));
    layer4_outputs(220) <= not(layer3_outputs(2354));
    layer4_outputs(221) <= layer3_outputs(2448);
    layer4_outputs(222) <= not(layer3_outputs(427));
    layer4_outputs(223) <= (layer3_outputs(2370)) or (layer3_outputs(2301));
    layer4_outputs(224) <= not(layer3_outputs(2105));
    layer4_outputs(225) <= not(layer3_outputs(1365)) or (layer3_outputs(1713));
    layer4_outputs(226) <= not(layer3_outputs(1964)) or (layer3_outputs(152));
    layer4_outputs(227) <= not(layer3_outputs(2494)) or (layer3_outputs(1312));
    layer4_outputs(228) <= not(layer3_outputs(1787));
    layer4_outputs(229) <= '0';
    layer4_outputs(230) <= not((layer3_outputs(2450)) or (layer3_outputs(14)));
    layer4_outputs(231) <= not(layer3_outputs(1306));
    layer4_outputs(232) <= layer3_outputs(1810);
    layer4_outputs(233) <= '0';
    layer4_outputs(234) <= (layer3_outputs(374)) or (layer3_outputs(1115));
    layer4_outputs(235) <= (layer3_outputs(243)) xor (layer3_outputs(280));
    layer4_outputs(236) <= not((layer3_outputs(1666)) or (layer3_outputs(1605)));
    layer4_outputs(237) <= (layer3_outputs(426)) and not (layer3_outputs(44));
    layer4_outputs(238) <= (layer3_outputs(2381)) or (layer3_outputs(5));
    layer4_outputs(239) <= (layer3_outputs(1317)) and not (layer3_outputs(1441));
    layer4_outputs(240) <= not(layer3_outputs(2534)) or (layer3_outputs(1633));
    layer4_outputs(241) <= not(layer3_outputs(2199));
    layer4_outputs(242) <= not(layer3_outputs(1123));
    layer4_outputs(243) <= (layer3_outputs(1728)) and (layer3_outputs(85));
    layer4_outputs(244) <= layer3_outputs(366);
    layer4_outputs(245) <= (layer3_outputs(666)) and not (layer3_outputs(92));
    layer4_outputs(246) <= '0';
    layer4_outputs(247) <= (layer3_outputs(2514)) and (layer3_outputs(119));
    layer4_outputs(248) <= not(layer3_outputs(1028));
    layer4_outputs(249) <= (layer3_outputs(2137)) xor (layer3_outputs(884));
    layer4_outputs(250) <= (layer3_outputs(1879)) or (layer3_outputs(779));
    layer4_outputs(251) <= (layer3_outputs(2363)) and not (layer3_outputs(550));
    layer4_outputs(252) <= not(layer3_outputs(430));
    layer4_outputs(253) <= not(layer3_outputs(1085));
    layer4_outputs(254) <= not(layer3_outputs(1378));
    layer4_outputs(255) <= (layer3_outputs(242)) and not (layer3_outputs(1868));
    layer4_outputs(256) <= layer3_outputs(721);
    layer4_outputs(257) <= not(layer3_outputs(1150)) or (layer3_outputs(995));
    layer4_outputs(258) <= layer3_outputs(2236);
    layer4_outputs(259) <= layer3_outputs(2277);
    layer4_outputs(260) <= not((layer3_outputs(2488)) and (layer3_outputs(473)));
    layer4_outputs(261) <= not(layer3_outputs(2065));
    layer4_outputs(262) <= not(layer3_outputs(1083)) or (layer3_outputs(274));
    layer4_outputs(263) <= layer3_outputs(1136);
    layer4_outputs(264) <= (layer3_outputs(2537)) or (layer3_outputs(213));
    layer4_outputs(265) <= not(layer3_outputs(1307)) or (layer3_outputs(1522));
    layer4_outputs(266) <= not(layer3_outputs(2492));
    layer4_outputs(267) <= not(layer3_outputs(1157));
    layer4_outputs(268) <= (layer3_outputs(329)) and not (layer3_outputs(2402));
    layer4_outputs(269) <= '1';
    layer4_outputs(270) <= '0';
    layer4_outputs(271) <= (layer3_outputs(1266)) and not (layer3_outputs(2117));
    layer4_outputs(272) <= layer3_outputs(262);
    layer4_outputs(273) <= not(layer3_outputs(1089));
    layer4_outputs(274) <= layer3_outputs(1764);
    layer4_outputs(275) <= not(layer3_outputs(586)) or (layer3_outputs(1375));
    layer4_outputs(276) <= layer3_outputs(2198);
    layer4_outputs(277) <= '0';
    layer4_outputs(278) <= not(layer3_outputs(2342));
    layer4_outputs(279) <= not(layer3_outputs(629));
    layer4_outputs(280) <= (layer3_outputs(1563)) xor (layer3_outputs(191));
    layer4_outputs(281) <= '0';
    layer4_outputs(282) <= layer3_outputs(960);
    layer4_outputs(283) <= not((layer3_outputs(1543)) and (layer3_outputs(1416)));
    layer4_outputs(284) <= '0';
    layer4_outputs(285) <= not((layer3_outputs(2049)) xor (layer3_outputs(2078)));
    layer4_outputs(286) <= layer3_outputs(84);
    layer4_outputs(287) <= (layer3_outputs(1217)) xor (layer3_outputs(2257));
    layer4_outputs(288) <= not((layer3_outputs(966)) and (layer3_outputs(1231)));
    layer4_outputs(289) <= not(layer3_outputs(194));
    layer4_outputs(290) <= layer3_outputs(2499);
    layer4_outputs(291) <= not(layer3_outputs(428));
    layer4_outputs(292) <= layer3_outputs(2436);
    layer4_outputs(293) <= not(layer3_outputs(63));
    layer4_outputs(294) <= layer3_outputs(798);
    layer4_outputs(295) <= not(layer3_outputs(533));
    layer4_outputs(296) <= '1';
    layer4_outputs(297) <= not((layer3_outputs(1688)) or (layer3_outputs(602)));
    layer4_outputs(298) <= not(layer3_outputs(2004));
    layer4_outputs(299) <= layer3_outputs(2066);
    layer4_outputs(300) <= layer3_outputs(1793);
    layer4_outputs(301) <= not(layer3_outputs(62));
    layer4_outputs(302) <= not(layer3_outputs(459)) or (layer3_outputs(538));
    layer4_outputs(303) <= layer3_outputs(1949);
    layer4_outputs(304) <= '1';
    layer4_outputs(305) <= not(layer3_outputs(677));
    layer4_outputs(306) <= not(layer3_outputs(2021)) or (layer3_outputs(542));
    layer4_outputs(307) <= (layer3_outputs(2449)) and not (layer3_outputs(480));
    layer4_outputs(308) <= layer3_outputs(499);
    layer4_outputs(309) <= layer3_outputs(958);
    layer4_outputs(310) <= not((layer3_outputs(2076)) and (layer3_outputs(1978)));
    layer4_outputs(311) <= not(layer3_outputs(2548)) or (layer3_outputs(555));
    layer4_outputs(312) <= (layer3_outputs(455)) and (layer3_outputs(2526));
    layer4_outputs(313) <= (layer3_outputs(266)) xor (layer3_outputs(948));
    layer4_outputs(314) <= (layer3_outputs(930)) or (layer3_outputs(2310));
    layer4_outputs(315) <= not((layer3_outputs(649)) or (layer3_outputs(1528)));
    layer4_outputs(316) <= '1';
    layer4_outputs(317) <= (layer3_outputs(1346)) xor (layer3_outputs(2460));
    layer4_outputs(318) <= layer3_outputs(1825);
    layer4_outputs(319) <= layer3_outputs(1034);
    layer4_outputs(320) <= not(layer3_outputs(2167)) or (layer3_outputs(219));
    layer4_outputs(321) <= (layer3_outputs(740)) and not (layer3_outputs(1024));
    layer4_outputs(322) <= layer3_outputs(946);
    layer4_outputs(323) <= not(layer3_outputs(1750));
    layer4_outputs(324) <= (layer3_outputs(2072)) and not (layer3_outputs(295));
    layer4_outputs(325) <= layer3_outputs(1499);
    layer4_outputs(326) <= layer3_outputs(1111);
    layer4_outputs(327) <= layer3_outputs(688);
    layer4_outputs(328) <= (layer3_outputs(2270)) and not (layer3_outputs(842));
    layer4_outputs(329) <= layer3_outputs(1780);
    layer4_outputs(330) <= layer3_outputs(2552);
    layer4_outputs(331) <= not((layer3_outputs(1291)) and (layer3_outputs(129)));
    layer4_outputs(332) <= layer3_outputs(1626);
    layer4_outputs(333) <= (layer3_outputs(1090)) and (layer3_outputs(1418));
    layer4_outputs(334) <= not((layer3_outputs(495)) and (layer3_outputs(580)));
    layer4_outputs(335) <= not(layer3_outputs(2459)) or (layer3_outputs(1491));
    layer4_outputs(336) <= (layer3_outputs(2351)) and not (layer3_outputs(1027));
    layer4_outputs(337) <= layer3_outputs(2319);
    layer4_outputs(338) <= (layer3_outputs(2317)) and (layer3_outputs(254));
    layer4_outputs(339) <= not((layer3_outputs(2345)) or (layer3_outputs(2161)));
    layer4_outputs(340) <= not((layer3_outputs(74)) and (layer3_outputs(1388)));
    layer4_outputs(341) <= not(layer3_outputs(2123)) or (layer3_outputs(1308));
    layer4_outputs(342) <= (layer3_outputs(365)) and not (layer3_outputs(2279));
    layer4_outputs(343) <= '1';
    layer4_outputs(344) <= not((layer3_outputs(1577)) and (layer3_outputs(510)));
    layer4_outputs(345) <= not((layer3_outputs(1547)) xor (layer3_outputs(37)));
    layer4_outputs(346) <= (layer3_outputs(1018)) or (layer3_outputs(170));
    layer4_outputs(347) <= not((layer3_outputs(614)) or (layer3_outputs(252)));
    layer4_outputs(348) <= '1';
    layer4_outputs(349) <= not((layer3_outputs(2245)) or (layer3_outputs(2288)));
    layer4_outputs(350) <= not(layer3_outputs(1748));
    layer4_outputs(351) <= not(layer3_outputs(1139));
    layer4_outputs(352) <= (layer3_outputs(1886)) or (layer3_outputs(1168));
    layer4_outputs(353) <= layer3_outputs(1466);
    layer4_outputs(354) <= not(layer3_outputs(1856));
    layer4_outputs(355) <= layer3_outputs(2207);
    layer4_outputs(356) <= not((layer3_outputs(892)) xor (layer3_outputs(463)));
    layer4_outputs(357) <= not((layer3_outputs(490)) and (layer3_outputs(1760)));
    layer4_outputs(358) <= layer3_outputs(334);
    layer4_outputs(359) <= not(layer3_outputs(217));
    layer4_outputs(360) <= (layer3_outputs(1427)) and not (layer3_outputs(413));
    layer4_outputs(361) <= (layer3_outputs(251)) and not (layer3_outputs(1051));
    layer4_outputs(362) <= not(layer3_outputs(1049));
    layer4_outputs(363) <= layer3_outputs(2321);
    layer4_outputs(364) <= not((layer3_outputs(1030)) or (layer3_outputs(432)));
    layer4_outputs(365) <= (layer3_outputs(1515)) and (layer3_outputs(261));
    layer4_outputs(366) <= not(layer3_outputs(263));
    layer4_outputs(367) <= (layer3_outputs(1639)) and not (layer3_outputs(835));
    layer4_outputs(368) <= not((layer3_outputs(710)) or (layer3_outputs(1938)));
    layer4_outputs(369) <= not(layer3_outputs(2445));
    layer4_outputs(370) <= layer3_outputs(850);
    layer4_outputs(371) <= (layer3_outputs(99)) or (layer3_outputs(573));
    layer4_outputs(372) <= not(layer3_outputs(341));
    layer4_outputs(373) <= not((layer3_outputs(975)) or (layer3_outputs(182)));
    layer4_outputs(374) <= layer3_outputs(1771);
    layer4_outputs(375) <= layer3_outputs(1319);
    layer4_outputs(376) <= layer3_outputs(2229);
    layer4_outputs(377) <= (layer3_outputs(214)) or (layer3_outputs(1264));
    layer4_outputs(378) <= layer3_outputs(1892);
    layer4_outputs(379) <= (layer3_outputs(2516)) xor (layer3_outputs(1705));
    layer4_outputs(380) <= '0';
    layer4_outputs(381) <= not(layer3_outputs(1664)) or (layer3_outputs(2164));
    layer4_outputs(382) <= (layer3_outputs(1196)) and not (layer3_outputs(1445));
    layer4_outputs(383) <= layer3_outputs(1223);
    layer4_outputs(384) <= '0';
    layer4_outputs(385) <= layer3_outputs(165);
    layer4_outputs(386) <= not(layer3_outputs(1528));
    layer4_outputs(387) <= not((layer3_outputs(268)) or (layer3_outputs(853)));
    layer4_outputs(388) <= '0';
    layer4_outputs(389) <= layer3_outputs(1531);
    layer4_outputs(390) <= '0';
    layer4_outputs(391) <= layer3_outputs(816);
    layer4_outputs(392) <= layer3_outputs(1648);
    layer4_outputs(393) <= (layer3_outputs(882)) and not (layer3_outputs(270));
    layer4_outputs(394) <= (layer3_outputs(2484)) and not (layer3_outputs(1598));
    layer4_outputs(395) <= not((layer3_outputs(2173)) and (layer3_outputs(2337)));
    layer4_outputs(396) <= not(layer3_outputs(868));
    layer4_outputs(397) <= not(layer3_outputs(2294));
    layer4_outputs(398) <= layer3_outputs(2539);
    layer4_outputs(399) <= '0';
    layer4_outputs(400) <= not(layer3_outputs(825));
    layer4_outputs(401) <= not(layer3_outputs(1455)) or (layer3_outputs(1134));
    layer4_outputs(402) <= (layer3_outputs(599)) and not (layer3_outputs(1296));
    layer4_outputs(403) <= layer3_outputs(804);
    layer4_outputs(404) <= layer3_outputs(465);
    layer4_outputs(405) <= not(layer3_outputs(2174));
    layer4_outputs(406) <= (layer3_outputs(496)) xor (layer3_outputs(2308));
    layer4_outputs(407) <= (layer3_outputs(1902)) and (layer3_outputs(640));
    layer4_outputs(408) <= not((layer3_outputs(624)) xor (layer3_outputs(1535)));
    layer4_outputs(409) <= layer3_outputs(144);
    layer4_outputs(410) <= (layer3_outputs(660)) and (layer3_outputs(1107));
    layer4_outputs(411) <= layer3_outputs(612);
    layer4_outputs(412) <= (layer3_outputs(418)) and not (layer3_outputs(1156));
    layer4_outputs(413) <= (layer3_outputs(1118)) and (layer3_outputs(33));
    layer4_outputs(414) <= '0';
    layer4_outputs(415) <= (layer3_outputs(1871)) and not (layer3_outputs(736));
    layer4_outputs(416) <= (layer3_outputs(1277)) or (layer3_outputs(1361));
    layer4_outputs(417) <= (layer3_outputs(48)) and not (layer3_outputs(531));
    layer4_outputs(418) <= (layer3_outputs(471)) xor (layer3_outputs(1942));
    layer4_outputs(419) <= (layer3_outputs(2228)) xor (layer3_outputs(560));
    layer4_outputs(420) <= (layer3_outputs(131)) and not (layer3_outputs(1442));
    layer4_outputs(421) <= not(layer3_outputs(1936)) or (layer3_outputs(292));
    layer4_outputs(422) <= not(layer3_outputs(1189));
    layer4_outputs(423) <= not(layer3_outputs(1333)) or (layer3_outputs(155));
    layer4_outputs(424) <= not((layer3_outputs(763)) or (layer3_outputs(315)));
    layer4_outputs(425) <= not((layer3_outputs(909)) and (layer3_outputs(235)));
    layer4_outputs(426) <= not(layer3_outputs(2323));
    layer4_outputs(427) <= not(layer3_outputs(1616));
    layer4_outputs(428) <= layer3_outputs(1579);
    layer4_outputs(429) <= (layer3_outputs(2242)) and not (layer3_outputs(1404));
    layer4_outputs(430) <= not(layer3_outputs(1124)) or (layer3_outputs(1660));
    layer4_outputs(431) <= layer3_outputs(1921);
    layer4_outputs(432) <= not(layer3_outputs(1918)) or (layer3_outputs(2311));
    layer4_outputs(433) <= layer3_outputs(469);
    layer4_outputs(434) <= (layer3_outputs(2252)) and (layer3_outputs(300));
    layer4_outputs(435) <= layer3_outputs(2366);
    layer4_outputs(436) <= not((layer3_outputs(2291)) or (layer3_outputs(785)));
    layer4_outputs(437) <= (layer3_outputs(1553)) and (layer3_outputs(985));
    layer4_outputs(438) <= '0';
    layer4_outputs(439) <= not(layer3_outputs(1792));
    layer4_outputs(440) <= not(layer3_outputs(1791));
    layer4_outputs(441) <= (layer3_outputs(1172)) and (layer3_outputs(972));
    layer4_outputs(442) <= (layer3_outputs(2396)) or (layer3_outputs(299));
    layer4_outputs(443) <= (layer3_outputs(704)) and not (layer3_outputs(1994));
    layer4_outputs(444) <= not(layer3_outputs(1014)) or (layer3_outputs(1829));
    layer4_outputs(445) <= layer3_outputs(368);
    layer4_outputs(446) <= not(layer3_outputs(364));
    layer4_outputs(447) <= not((layer3_outputs(1654)) and (layer3_outputs(1078)));
    layer4_outputs(448) <= not(layer3_outputs(25)) or (layer3_outputs(1923));
    layer4_outputs(449) <= layer3_outputs(2320);
    layer4_outputs(450) <= (layer3_outputs(1630)) and not (layer3_outputs(625));
    layer4_outputs(451) <= (layer3_outputs(1018)) or (layer3_outputs(1575));
    layer4_outputs(452) <= layer3_outputs(923);
    layer4_outputs(453) <= (layer3_outputs(1514)) and not (layer3_outputs(1039));
    layer4_outputs(454) <= layer3_outputs(2345);
    layer4_outputs(455) <= layer3_outputs(1382);
    layer4_outputs(456) <= not(layer3_outputs(1547));
    layer4_outputs(457) <= (layer3_outputs(2429)) or (layer3_outputs(807));
    layer4_outputs(458) <= (layer3_outputs(793)) or (layer3_outputs(2419));
    layer4_outputs(459) <= not((layer3_outputs(1909)) and (layer3_outputs(926)));
    layer4_outputs(460) <= not(layer3_outputs(912)) or (layer3_outputs(643));
    layer4_outputs(461) <= layer3_outputs(1116);
    layer4_outputs(462) <= not((layer3_outputs(1460)) or (layer3_outputs(361)));
    layer4_outputs(463) <= not(layer3_outputs(828));
    layer4_outputs(464) <= not(layer3_outputs(802)) or (layer3_outputs(344));
    layer4_outputs(465) <= not(layer3_outputs(2454));
    layer4_outputs(466) <= not(layer3_outputs(2173));
    layer4_outputs(467) <= (layer3_outputs(669)) and not (layer3_outputs(2324));
    layer4_outputs(468) <= layer3_outputs(712);
    layer4_outputs(469) <= (layer3_outputs(1748)) and not (layer3_outputs(929));
    layer4_outputs(470) <= (layer3_outputs(1981)) xor (layer3_outputs(1177));
    layer4_outputs(471) <= (layer3_outputs(1960)) and (layer3_outputs(1190));
    layer4_outputs(472) <= not(layer3_outputs(2133));
    layer4_outputs(473) <= not((layer3_outputs(2520)) and (layer3_outputs(734)));
    layer4_outputs(474) <= (layer3_outputs(39)) and (layer3_outputs(517));
    layer4_outputs(475) <= not(layer3_outputs(493)) or (layer3_outputs(215));
    layer4_outputs(476) <= not(layer3_outputs(1550)) or (layer3_outputs(1799));
    layer4_outputs(477) <= not((layer3_outputs(1680)) or (layer3_outputs(658)));
    layer4_outputs(478) <= (layer3_outputs(114)) or (layer3_outputs(481));
    layer4_outputs(479) <= '0';
    layer4_outputs(480) <= (layer3_outputs(1763)) and not (layer3_outputs(241));
    layer4_outputs(481) <= not(layer3_outputs(707));
    layer4_outputs(482) <= '0';
    layer4_outputs(483) <= not(layer3_outputs(541)) or (layer3_outputs(1827));
    layer4_outputs(484) <= not((layer3_outputs(1479)) and (layer3_outputs(356)));
    layer4_outputs(485) <= (layer3_outputs(1588)) and not (layer3_outputs(1240));
    layer4_outputs(486) <= not(layer3_outputs(316)) or (layer3_outputs(605));
    layer4_outputs(487) <= not(layer3_outputs(2122));
    layer4_outputs(488) <= (layer3_outputs(1769)) or (layer3_outputs(482));
    layer4_outputs(489) <= not(layer3_outputs(2367)) or (layer3_outputs(2285));
    layer4_outputs(490) <= (layer3_outputs(567)) and (layer3_outputs(754));
    layer4_outputs(491) <= not(layer3_outputs(2240));
    layer4_outputs(492) <= not((layer3_outputs(1500)) xor (layer3_outputs(908)));
    layer4_outputs(493) <= not((layer3_outputs(66)) and (layer3_outputs(2141)));
    layer4_outputs(494) <= layer3_outputs(1419);
    layer4_outputs(495) <= not(layer3_outputs(2144));
    layer4_outputs(496) <= (layer3_outputs(821)) and (layer3_outputs(1144));
    layer4_outputs(497) <= (layer3_outputs(1936)) and (layer3_outputs(156));
    layer4_outputs(498) <= (layer3_outputs(313)) or (layer3_outputs(1005));
    layer4_outputs(499) <= not((layer3_outputs(684)) or (layer3_outputs(604)));
    layer4_outputs(500) <= not(layer3_outputs(256));
    layer4_outputs(501) <= (layer3_outputs(1647)) and not (layer3_outputs(2398));
    layer4_outputs(502) <= (layer3_outputs(2404)) and (layer3_outputs(561));
    layer4_outputs(503) <= not(layer3_outputs(415)) or (layer3_outputs(511));
    layer4_outputs(504) <= layer3_outputs(2344);
    layer4_outputs(505) <= (layer3_outputs(1990)) and (layer3_outputs(168));
    layer4_outputs(506) <= not(layer3_outputs(117));
    layer4_outputs(507) <= not(layer3_outputs(2369));
    layer4_outputs(508) <= '0';
    layer4_outputs(509) <= (layer3_outputs(1541)) and not (layer3_outputs(741));
    layer4_outputs(510) <= not((layer3_outputs(424)) or (layer3_outputs(2107)));
    layer4_outputs(511) <= not(layer3_outputs(1));
    layer4_outputs(512) <= not(layer3_outputs(2057));
    layer4_outputs(513) <= layer3_outputs(924);
    layer4_outputs(514) <= layer3_outputs(248);
    layer4_outputs(515) <= (layer3_outputs(597)) or (layer3_outputs(364));
    layer4_outputs(516) <= '1';
    layer4_outputs(517) <= not(layer3_outputs(2060));
    layer4_outputs(518) <= not((layer3_outputs(2025)) or (layer3_outputs(1474)));
    layer4_outputs(519) <= (layer3_outputs(1249)) and not (layer3_outputs(1106));
    layer4_outputs(520) <= '0';
    layer4_outputs(521) <= (layer3_outputs(1755)) xor (layer3_outputs(391));
    layer4_outputs(522) <= layer3_outputs(2068);
    layer4_outputs(523) <= (layer3_outputs(64)) and (layer3_outputs(1349));
    layer4_outputs(524) <= layer3_outputs(1330);
    layer4_outputs(525) <= not(layer3_outputs(823));
    layer4_outputs(526) <= not(layer3_outputs(1191));
    layer4_outputs(527) <= layer3_outputs(2219);
    layer4_outputs(528) <= layer3_outputs(2275);
    layer4_outputs(529) <= layer3_outputs(2002);
    layer4_outputs(530) <= not((layer3_outputs(1774)) and (layer3_outputs(2430)));
    layer4_outputs(531) <= (layer3_outputs(230)) and not (layer3_outputs(1101));
    layer4_outputs(532) <= not(layer3_outputs(1503)) or (layer3_outputs(394));
    layer4_outputs(533) <= (layer3_outputs(305)) and not (layer3_outputs(1421));
    layer4_outputs(534) <= layer3_outputs(310);
    layer4_outputs(535) <= layer3_outputs(2342);
    layer4_outputs(536) <= not(layer3_outputs(136));
    layer4_outputs(537) <= not(layer3_outputs(1841));
    layer4_outputs(538) <= not(layer3_outputs(1295)) or (layer3_outputs(1534));
    layer4_outputs(539) <= not(layer3_outputs(229));
    layer4_outputs(540) <= (layer3_outputs(1386)) and not (layer3_outputs(2505));
    layer4_outputs(541) <= (layer3_outputs(1625)) and (layer3_outputs(1327));
    layer4_outputs(542) <= layer3_outputs(1057);
    layer4_outputs(543) <= not(layer3_outputs(2533));
    layer4_outputs(544) <= layer3_outputs(2553);
    layer4_outputs(545) <= not(layer3_outputs(1685)) or (layer3_outputs(2113));
    layer4_outputs(546) <= not(layer3_outputs(2441));
    layer4_outputs(547) <= (layer3_outputs(861)) and not (layer3_outputs(515));
    layer4_outputs(548) <= (layer3_outputs(1395)) and not (layer3_outputs(490));
    layer4_outputs(549) <= not(layer3_outputs(958));
    layer4_outputs(550) <= not(layer3_outputs(1489));
    layer4_outputs(551) <= not(layer3_outputs(949)) or (layer3_outputs(1708));
    layer4_outputs(552) <= (layer3_outputs(46)) or (layer3_outputs(1370));
    layer4_outputs(553) <= (layer3_outputs(1288)) or (layer3_outputs(977));
    layer4_outputs(554) <= layer3_outputs(824);
    layer4_outputs(555) <= layer3_outputs(2053);
    layer4_outputs(556) <= not(layer3_outputs(2425));
    layer4_outputs(557) <= (layer3_outputs(1433)) or (layer3_outputs(1096));
    layer4_outputs(558) <= not((layer3_outputs(1360)) or (layer3_outputs(2322)));
    layer4_outputs(559) <= (layer3_outputs(1719)) and not (layer3_outputs(1651));
    layer4_outputs(560) <= not(layer3_outputs(1381)) or (layer3_outputs(2205));
    layer4_outputs(561) <= (layer3_outputs(1056)) and not (layer3_outputs(1027));
    layer4_outputs(562) <= not(layer3_outputs(339)) or (layer3_outputs(566));
    layer4_outputs(563) <= '1';
    layer4_outputs(564) <= not(layer3_outputs(1394));
    layer4_outputs(565) <= '1';
    layer4_outputs(566) <= '0';
    layer4_outputs(567) <= layer3_outputs(695);
    layer4_outputs(568) <= not(layer3_outputs(821));
    layer4_outputs(569) <= not(layer3_outputs(675));
    layer4_outputs(570) <= (layer3_outputs(1711)) and not (layer3_outputs(1098));
    layer4_outputs(571) <= not((layer3_outputs(171)) or (layer3_outputs(439)));
    layer4_outputs(572) <= not(layer3_outputs(2035));
    layer4_outputs(573) <= '0';
    layer4_outputs(574) <= layer3_outputs(2539);
    layer4_outputs(575) <= layer3_outputs(2222);
    layer4_outputs(576) <= layer3_outputs(921);
    layer4_outputs(577) <= (layer3_outputs(399)) xor (layer3_outputs(1884));
    layer4_outputs(578) <= (layer3_outputs(2299)) and not (layer3_outputs(1941));
    layer4_outputs(579) <= not(layer3_outputs(918));
    layer4_outputs(580) <= not(layer3_outputs(1823));
    layer4_outputs(581) <= not((layer3_outputs(1928)) and (layer3_outputs(2498)));
    layer4_outputs(582) <= layer3_outputs(313);
    layer4_outputs(583) <= layer3_outputs(2121);
    layer4_outputs(584) <= layer3_outputs(744);
    layer4_outputs(585) <= (layer3_outputs(2125)) xor (layer3_outputs(1430));
    layer4_outputs(586) <= layer3_outputs(1658);
    layer4_outputs(587) <= not(layer3_outputs(653));
    layer4_outputs(588) <= (layer3_outputs(2449)) and (layer3_outputs(1812));
    layer4_outputs(589) <= '0';
    layer4_outputs(590) <= layer3_outputs(2267);
    layer4_outputs(591) <= layer3_outputs(1451);
    layer4_outputs(592) <= not(layer3_outputs(69)) or (layer3_outputs(379));
    layer4_outputs(593) <= '0';
    layer4_outputs(594) <= layer3_outputs(2455);
    layer4_outputs(595) <= (layer3_outputs(1197)) and (layer3_outputs(49));
    layer4_outputs(596) <= not(layer3_outputs(1995));
    layer4_outputs(597) <= (layer3_outputs(2309)) and (layer3_outputs(1132));
    layer4_outputs(598) <= not(layer3_outputs(177));
    layer4_outputs(599) <= not((layer3_outputs(483)) and (layer3_outputs(1796)));
    layer4_outputs(600) <= (layer3_outputs(205)) or (layer3_outputs(887));
    layer4_outputs(601) <= layer3_outputs(796);
    layer4_outputs(602) <= not((layer3_outputs(152)) or (layer3_outputs(101)));
    layer4_outputs(603) <= (layer3_outputs(118)) or (layer3_outputs(1716));
    layer4_outputs(604) <= layer3_outputs(876);
    layer4_outputs(605) <= '0';
    layer4_outputs(606) <= (layer3_outputs(340)) and (layer3_outputs(973));
    layer4_outputs(607) <= not((layer3_outputs(991)) and (layer3_outputs(491)));
    layer4_outputs(608) <= layer3_outputs(2401);
    layer4_outputs(609) <= not((layer3_outputs(1429)) or (layer3_outputs(462)));
    layer4_outputs(610) <= not((layer3_outputs(437)) xor (layer3_outputs(2155)));
    layer4_outputs(611) <= (layer3_outputs(2298)) and (layer3_outputs(240));
    layer4_outputs(612) <= not((layer3_outputs(272)) or (layer3_outputs(2116)));
    layer4_outputs(613) <= not((layer3_outputs(2109)) xor (layer3_outputs(1133)));
    layer4_outputs(614) <= not((layer3_outputs(787)) and (layer3_outputs(1418)));
    layer4_outputs(615) <= (layer3_outputs(2198)) xor (layer3_outputs(1348));
    layer4_outputs(616) <= layer3_outputs(127);
    layer4_outputs(617) <= '0';
    layer4_outputs(618) <= not(layer3_outputs(1700));
    layer4_outputs(619) <= not(layer3_outputs(903)) or (layer3_outputs(1535));
    layer4_outputs(620) <= not(layer3_outputs(1093));
    layer4_outputs(621) <= (layer3_outputs(922)) or (layer3_outputs(761));
    layer4_outputs(622) <= not(layer3_outputs(945));
    layer4_outputs(623) <= not((layer3_outputs(962)) and (layer3_outputs(42)));
    layer4_outputs(624) <= '1';
    layer4_outputs(625) <= not(layer3_outputs(840));
    layer4_outputs(626) <= not(layer3_outputs(693));
    layer4_outputs(627) <= not(layer3_outputs(210));
    layer4_outputs(628) <= not((layer3_outputs(417)) or (layer3_outputs(2521)));
    layer4_outputs(629) <= not((layer3_outputs(1331)) or (layer3_outputs(2348)));
    layer4_outputs(630) <= not(layer3_outputs(2491)) or (layer3_outputs(1044));
    layer4_outputs(631) <= '1';
    layer4_outputs(632) <= layer3_outputs(1583);
    layer4_outputs(633) <= not((layer3_outputs(1057)) and (layer3_outputs(804)));
    layer4_outputs(634) <= not(layer3_outputs(2156));
    layer4_outputs(635) <= (layer3_outputs(1709)) and not (layer3_outputs(403));
    layer4_outputs(636) <= (layer3_outputs(1283)) or (layer3_outputs(557));
    layer4_outputs(637) <= not(layer3_outputs(1350)) or (layer3_outputs(306));
    layer4_outputs(638) <= '0';
    layer4_outputs(639) <= not((layer3_outputs(2460)) xor (layer3_outputs(1422)));
    layer4_outputs(640) <= not(layer3_outputs(165));
    layer4_outputs(641) <= (layer3_outputs(1274)) and (layer3_outputs(1316));
    layer4_outputs(642) <= not(layer3_outputs(671)) or (layer3_outputs(357));
    layer4_outputs(643) <= (layer3_outputs(2029)) and not (layer3_outputs(2381));
    layer4_outputs(644) <= layer3_outputs(2211);
    layer4_outputs(645) <= not(layer3_outputs(1249));
    layer4_outputs(646) <= (layer3_outputs(1928)) and not (layer3_outputs(293));
    layer4_outputs(647) <= not(layer3_outputs(1065));
    layer4_outputs(648) <= not(layer3_outputs(1227));
    layer4_outputs(649) <= not(layer3_outputs(540));
    layer4_outputs(650) <= layer3_outputs(2529);
    layer4_outputs(651) <= (layer3_outputs(7)) and not (layer3_outputs(2384));
    layer4_outputs(652) <= not((layer3_outputs(1669)) xor (layer3_outputs(2528)));
    layer4_outputs(653) <= '1';
    layer4_outputs(654) <= layer3_outputs(175);
    layer4_outputs(655) <= layer3_outputs(1034);
    layer4_outputs(656) <= layer3_outputs(964);
    layer4_outputs(657) <= layer3_outputs(1826);
    layer4_outputs(658) <= not(layer3_outputs(2477)) or (layer3_outputs(944));
    layer4_outputs(659) <= not(layer3_outputs(2248)) or (layer3_outputs(1447));
    layer4_outputs(660) <= not(layer3_outputs(1383));
    layer4_outputs(661) <= not(layer3_outputs(168)) or (layer3_outputs(1652));
    layer4_outputs(662) <= not((layer3_outputs(635)) and (layer3_outputs(1578)));
    layer4_outputs(663) <= not((layer3_outputs(844)) or (layer3_outputs(1677)));
    layer4_outputs(664) <= (layer3_outputs(2254)) and not (layer3_outputs(484));
    layer4_outputs(665) <= (layer3_outputs(623)) or (layer3_outputs(2235));
    layer4_outputs(666) <= not(layer3_outputs(2312));
    layer4_outputs(667) <= '1';
    layer4_outputs(668) <= (layer3_outputs(1637)) or (layer3_outputs(396));
    layer4_outputs(669) <= layer3_outputs(118);
    layer4_outputs(670) <= layer3_outputs(1445);
    layer4_outputs(671) <= layer3_outputs(2518);
    layer4_outputs(672) <= not((layer3_outputs(1243)) or (layer3_outputs(1285)));
    layer4_outputs(673) <= not((layer3_outputs(1777)) or (layer3_outputs(2099)));
    layer4_outputs(674) <= (layer3_outputs(1638)) or (layer3_outputs(2255));
    layer4_outputs(675) <= not(layer3_outputs(669));
    layer4_outputs(676) <= '0';
    layer4_outputs(677) <= (layer3_outputs(872)) and (layer3_outputs(940));
    layer4_outputs(678) <= not(layer3_outputs(1577)) or (layer3_outputs(2148));
    layer4_outputs(679) <= (layer3_outputs(638)) or (layer3_outputs(2523));
    layer4_outputs(680) <= not(layer3_outputs(860));
    layer4_outputs(681) <= not(layer3_outputs(822));
    layer4_outputs(682) <= not(layer3_outputs(50)) or (layer3_outputs(22));
    layer4_outputs(683) <= '0';
    layer4_outputs(684) <= not(layer3_outputs(444));
    layer4_outputs(685) <= (layer3_outputs(2555)) or (layer3_outputs(700));
    layer4_outputs(686) <= (layer3_outputs(923)) and not (layer3_outputs(736));
    layer4_outputs(687) <= layer3_outputs(1297);
    layer4_outputs(688) <= not(layer3_outputs(456));
    layer4_outputs(689) <= not(layer3_outputs(1140)) or (layer3_outputs(2088));
    layer4_outputs(690) <= not(layer3_outputs(1305)) or (layer3_outputs(1848));
    layer4_outputs(691) <= (layer3_outputs(1038)) or (layer3_outputs(999));
    layer4_outputs(692) <= layer3_outputs(875);
    layer4_outputs(693) <= not((layer3_outputs(1542)) xor (layer3_outputs(1103)));
    layer4_outputs(694) <= (layer3_outputs(1920)) and not (layer3_outputs(1517));
    layer4_outputs(695) <= not(layer3_outputs(1859));
    layer4_outputs(696) <= layer3_outputs(771);
    layer4_outputs(697) <= not(layer3_outputs(6));
    layer4_outputs(698) <= not((layer3_outputs(1974)) or (layer3_outputs(297)));
    layer4_outputs(699) <= not(layer3_outputs(1724));
    layer4_outputs(700) <= not(layer3_outputs(2182));
    layer4_outputs(701) <= not(layer3_outputs(1580));
    layer4_outputs(702) <= not((layer3_outputs(125)) or (layer3_outputs(7)));
    layer4_outputs(703) <= not(layer3_outputs(2388));
    layer4_outputs(704) <= layer3_outputs(1328);
    layer4_outputs(705) <= (layer3_outputs(1876)) and not (layer3_outputs(2119));
    layer4_outputs(706) <= (layer3_outputs(323)) and not (layer3_outputs(346));
    layer4_outputs(707) <= (layer3_outputs(1393)) and (layer3_outputs(855));
    layer4_outputs(708) <= not(layer3_outputs(282));
    layer4_outputs(709) <= not(layer3_outputs(188)) or (layer3_outputs(1948));
    layer4_outputs(710) <= (layer3_outputs(1284)) xor (layer3_outputs(706));
    layer4_outputs(711) <= not(layer3_outputs(747));
    layer4_outputs(712) <= not(layer3_outputs(1996));
    layer4_outputs(713) <= layer3_outputs(1601);
    layer4_outputs(714) <= not(layer3_outputs(1128));
    layer4_outputs(715) <= not((layer3_outputs(453)) or (layer3_outputs(592)));
    layer4_outputs(716) <= '1';
    layer4_outputs(717) <= not(layer3_outputs(425));
    layer4_outputs(718) <= not((layer3_outputs(2071)) and (layer3_outputs(437)));
    layer4_outputs(719) <= (layer3_outputs(1614)) or (layer3_outputs(832));
    layer4_outputs(720) <= layer3_outputs(2069);
    layer4_outputs(721) <= not(layer3_outputs(1757));
    layer4_outputs(722) <= not(layer3_outputs(1201)) or (layer3_outputs(1493));
    layer4_outputs(723) <= not(layer3_outputs(1833));
    layer4_outputs(724) <= (layer3_outputs(531)) and (layer3_outputs(1886));
    layer4_outputs(725) <= not(layer3_outputs(281));
    layer4_outputs(726) <= not((layer3_outputs(2551)) xor (layer3_outputs(2262)));
    layer4_outputs(727) <= layer3_outputs(1795);
    layer4_outputs(728) <= not((layer3_outputs(2530)) and (layer3_outputs(897)));
    layer4_outputs(729) <= layer3_outputs(2039);
    layer4_outputs(730) <= not(layer3_outputs(1333)) or (layer3_outputs(2044));
    layer4_outputs(731) <= not(layer3_outputs(392));
    layer4_outputs(732) <= layer3_outputs(813);
    layer4_outputs(733) <= not(layer3_outputs(1677)) or (layer3_outputs(1831));
    layer4_outputs(734) <= layer3_outputs(1966);
    layer4_outputs(735) <= (layer3_outputs(846)) and not (layer3_outputs(372));
    layer4_outputs(736) <= not(layer3_outputs(206));
    layer4_outputs(737) <= not((layer3_outputs(1549)) and (layer3_outputs(1431)));
    layer4_outputs(738) <= layer3_outputs(1917);
    layer4_outputs(739) <= (layer3_outputs(589)) or (layer3_outputs(572));
    layer4_outputs(740) <= not(layer3_outputs(1692)) or (layer3_outputs(104));
    layer4_outputs(741) <= (layer3_outputs(2017)) xor (layer3_outputs(2264));
    layer4_outputs(742) <= not(layer3_outputs(2507)) or (layer3_outputs(959));
    layer4_outputs(743) <= not(layer3_outputs(1366)) or (layer3_outputs(642));
    layer4_outputs(744) <= not(layer3_outputs(404));
    layer4_outputs(745) <= (layer3_outputs(1174)) and not (layer3_outputs(2349));
    layer4_outputs(746) <= layer3_outputs(2213);
    layer4_outputs(747) <= (layer3_outputs(1657)) and not (layer3_outputs(796));
    layer4_outputs(748) <= not(layer3_outputs(2325)) or (layer3_outputs(2223));
    layer4_outputs(749) <= not((layer3_outputs(1406)) and (layer3_outputs(2355)));
    layer4_outputs(750) <= '1';
    layer4_outputs(751) <= not(layer3_outputs(1519));
    layer4_outputs(752) <= layer3_outputs(1444);
    layer4_outputs(753) <= layer3_outputs(1683);
    layer4_outputs(754) <= '1';
    layer4_outputs(755) <= not(layer3_outputs(2442)) or (layer3_outputs(1894));
    layer4_outputs(756) <= layer3_outputs(1861);
    layer4_outputs(757) <= not(layer3_outputs(1358)) or (layer3_outputs(620));
    layer4_outputs(758) <= layer3_outputs(2089);
    layer4_outputs(759) <= layer3_outputs(88);
    layer4_outputs(760) <= not((layer3_outputs(827)) or (layer3_outputs(1485)));
    layer4_outputs(761) <= not(layer3_outputs(2227));
    layer4_outputs(762) <= not((layer3_outputs(1896)) or (layer3_outputs(15)));
    layer4_outputs(763) <= layer3_outputs(1462);
    layer4_outputs(764) <= (layer3_outputs(1260)) xor (layer3_outputs(239));
    layer4_outputs(765) <= layer3_outputs(1934);
    layer4_outputs(766) <= layer3_outputs(1182);
    layer4_outputs(767) <= not(layer3_outputs(256));
    layer4_outputs(768) <= layer3_outputs(1485);
    layer4_outputs(769) <= layer3_outputs(1400);
    layer4_outputs(770) <= not((layer3_outputs(1364)) and (layer3_outputs(507)));
    layer4_outputs(771) <= not(layer3_outputs(1484));
    layer4_outputs(772) <= (layer3_outputs(1236)) or (layer3_outputs(888));
    layer4_outputs(773) <= (layer3_outputs(1278)) or (layer3_outputs(2153));
    layer4_outputs(774) <= (layer3_outputs(484)) and not (layer3_outputs(1638));
    layer4_outputs(775) <= not(layer3_outputs(839));
    layer4_outputs(776) <= not(layer3_outputs(1156)) or (layer3_outputs(869));
    layer4_outputs(777) <= (layer3_outputs(803)) and (layer3_outputs(2545));
    layer4_outputs(778) <= layer3_outputs(579);
    layer4_outputs(779) <= (layer3_outputs(1506)) and not (layer3_outputs(1740));
    layer4_outputs(780) <= not((layer3_outputs(1)) or (layer3_outputs(100)));
    layer4_outputs(781) <= not(layer3_outputs(2034));
    layer4_outputs(782) <= (layer3_outputs(2151)) and not (layer3_outputs(745));
    layer4_outputs(783) <= '0';
    layer4_outputs(784) <= (layer3_outputs(1192)) and (layer3_outputs(2442));
    layer4_outputs(785) <= not((layer3_outputs(679)) and (layer3_outputs(1891)));
    layer4_outputs(786) <= layer3_outputs(1170);
    layer4_outputs(787) <= not((layer3_outputs(98)) xor (layer3_outputs(517)));
    layer4_outputs(788) <= (layer3_outputs(166)) or (layer3_outputs(811));
    layer4_outputs(789) <= (layer3_outputs(1368)) and not (layer3_outputs(862));
    layer4_outputs(790) <= '1';
    layer4_outputs(791) <= not(layer3_outputs(2026));
    layer4_outputs(792) <= layer3_outputs(608);
    layer4_outputs(793) <= (layer3_outputs(1117)) and not (layer3_outputs(1016));
    layer4_outputs(794) <= '0';
    layer4_outputs(795) <= not(layer3_outputs(808)) or (layer3_outputs(181));
    layer4_outputs(796) <= (layer3_outputs(1835)) or (layer3_outputs(984));
    layer4_outputs(797) <= not(layer3_outputs(692));
    layer4_outputs(798) <= layer3_outputs(2466);
    layer4_outputs(799) <= (layer3_outputs(1044)) or (layer3_outputs(1351));
    layer4_outputs(800) <= not(layer3_outputs(34));
    layer4_outputs(801) <= not(layer3_outputs(2166)) or (layer3_outputs(2278));
    layer4_outputs(802) <= not((layer3_outputs(2358)) and (layer3_outputs(991)));
    layer4_outputs(803) <= not(layer3_outputs(311)) or (layer3_outputs(549));
    layer4_outputs(804) <= not((layer3_outputs(1775)) and (layer3_outputs(2239)));
    layer4_outputs(805) <= (layer3_outputs(67)) and not (layer3_outputs(470));
    layer4_outputs(806) <= (layer3_outputs(1579)) or (layer3_outputs(1177));
    layer4_outputs(807) <= not(layer3_outputs(1589));
    layer4_outputs(808) <= layer3_outputs(790);
    layer4_outputs(809) <= not(layer3_outputs(1389));
    layer4_outputs(810) <= (layer3_outputs(2329)) and not (layer3_outputs(1457));
    layer4_outputs(811) <= not(layer3_outputs(1676));
    layer4_outputs(812) <= (layer3_outputs(1656)) and (layer3_outputs(458));
    layer4_outputs(813) <= (layer3_outputs(781)) and not (layer3_outputs(2268));
    layer4_outputs(814) <= layer3_outputs(795);
    layer4_outputs(815) <= layer3_outputs(2275);
    layer4_outputs(816) <= (layer3_outputs(19)) and not (layer3_outputs(1155));
    layer4_outputs(817) <= layer3_outputs(1521);
    layer4_outputs(818) <= not(layer3_outputs(2246)) or (layer3_outputs(2396));
    layer4_outputs(819) <= not((layer3_outputs(980)) and (layer3_outputs(1080)));
    layer4_outputs(820) <= layer3_outputs(1697);
    layer4_outputs(821) <= not(layer3_outputs(998)) or (layer3_outputs(2187));
    layer4_outputs(822) <= (layer3_outputs(341)) and (layer3_outputs(2400));
    layer4_outputs(823) <= layer3_outputs(1063);
    layer4_outputs(824) <= (layer3_outputs(161)) and (layer3_outputs(347));
    layer4_outputs(825) <= not(layer3_outputs(301)) or (layer3_outputs(1984));
    layer4_outputs(826) <= not((layer3_outputs(234)) xor (layer3_outputs(788)));
    layer4_outputs(827) <= '0';
    layer4_outputs(828) <= not(layer3_outputs(1204));
    layer4_outputs(829) <= (layer3_outputs(596)) and (layer3_outputs(402));
    layer4_outputs(830) <= not(layer3_outputs(1440));
    layer4_outputs(831) <= layer3_outputs(2005);
    layer4_outputs(832) <= (layer3_outputs(876)) and not (layer3_outputs(1142));
    layer4_outputs(833) <= layer3_outputs(2326);
    layer4_outputs(834) <= '1';
    layer4_outputs(835) <= not((layer3_outputs(2206)) or (layer3_outputs(857)));
    layer4_outputs(836) <= (layer3_outputs(1915)) and not (layer3_outputs(1311));
    layer4_outputs(837) <= not(layer3_outputs(2404));
    layer4_outputs(838) <= layer3_outputs(2320);
    layer4_outputs(839) <= layer3_outputs(678);
    layer4_outputs(840) <= '1';
    layer4_outputs(841) <= not(layer3_outputs(920));
    layer4_outputs(842) <= not((layer3_outputs(1612)) or (layer3_outputs(229)));
    layer4_outputs(843) <= '0';
    layer4_outputs(844) <= not(layer3_outputs(454));
    layer4_outputs(845) <= not(layer3_outputs(2392));
    layer4_outputs(846) <= not(layer3_outputs(79)) or (layer3_outputs(1888));
    layer4_outputs(847) <= (layer3_outputs(2030)) and not (layer3_outputs(2542));
    layer4_outputs(848) <= layer3_outputs(660);
    layer4_outputs(849) <= not((layer3_outputs(489)) and (layer3_outputs(792)));
    layer4_outputs(850) <= layer3_outputs(762);
    layer4_outputs(851) <= not(layer3_outputs(1777));
    layer4_outputs(852) <= (layer3_outputs(611)) and not (layer3_outputs(2558));
    layer4_outputs(853) <= '1';
    layer4_outputs(854) <= not((layer3_outputs(2036)) and (layer3_outputs(537)));
    layer4_outputs(855) <= not((layer3_outputs(470)) and (layer3_outputs(1037)));
    layer4_outputs(856) <= layer3_outputs(1663);
    layer4_outputs(857) <= not(layer3_outputs(607));
    layer4_outputs(858) <= not(layer3_outputs(2096));
    layer4_outputs(859) <= not((layer3_outputs(2003)) and (layer3_outputs(2023)));
    layer4_outputs(860) <= (layer3_outputs(2443)) and not (layer3_outputs(855));
    layer4_outputs(861) <= not(layer3_outputs(1854));
    layer4_outputs(862) <= not(layer3_outputs(1022));
    layer4_outputs(863) <= (layer3_outputs(1267)) or (layer3_outputs(2513));
    layer4_outputs(864) <= (layer3_outputs(2378)) xor (layer3_outputs(541));
    layer4_outputs(865) <= layer3_outputs(1960);
    layer4_outputs(866) <= not(layer3_outputs(2124)) or (layer3_outputs(1513));
    layer4_outputs(867) <= not((layer3_outputs(815)) xor (layer3_outputs(2397)));
    layer4_outputs(868) <= not(layer3_outputs(1897));
    layer4_outputs(869) <= (layer3_outputs(2213)) and not (layer3_outputs(1786));
    layer4_outputs(870) <= not(layer3_outputs(1099)) or (layer3_outputs(554));
    layer4_outputs(871) <= (layer3_outputs(69)) and not (layer3_outputs(434));
    layer4_outputs(872) <= (layer3_outputs(117)) and not (layer3_outputs(135));
    layer4_outputs(873) <= '0';
    layer4_outputs(874) <= (layer3_outputs(1324)) and not (layer3_outputs(2178));
    layer4_outputs(875) <= '1';
    layer4_outputs(876) <= (layer3_outputs(1317)) and not (layer3_outputs(620));
    layer4_outputs(877) <= not(layer3_outputs(1347));
    layer4_outputs(878) <= layer3_outputs(592);
    layer4_outputs(879) <= layer3_outputs(43);
    layer4_outputs(880) <= (layer3_outputs(637)) xor (layer3_outputs(2525));
    layer4_outputs(881) <= not((layer3_outputs(1605)) or (layer3_outputs(2235)));
    layer4_outputs(882) <= layer3_outputs(2076);
    layer4_outputs(883) <= not(layer3_outputs(1775)) or (layer3_outputs(1105));
    layer4_outputs(884) <= '0';
    layer4_outputs(885) <= layer3_outputs(2047);
    layer4_outputs(886) <= not(layer3_outputs(1384));
    layer4_outputs(887) <= not(layer3_outputs(830));
    layer4_outputs(888) <= layer3_outputs(1476);
    layer4_outputs(889) <= not(layer3_outputs(1469)) or (layer3_outputs(1345));
    layer4_outputs(890) <= not((layer3_outputs(1063)) and (layer3_outputs(1464)));
    layer4_outputs(891) <= '0';
    layer4_outputs(892) <= not(layer3_outputs(697));
    layer4_outputs(893) <= (layer3_outputs(551)) and not (layer3_outputs(380));
    layer4_outputs(894) <= layer3_outputs(2506);
    layer4_outputs(895) <= not(layer3_outputs(2095));
    layer4_outputs(896) <= not(layer3_outputs(912)) or (layer3_outputs(353));
    layer4_outputs(897) <= '1';
    layer4_outputs(898) <= (layer3_outputs(443)) or (layer3_outputs(756));
    layer4_outputs(899) <= not((layer3_outputs(2010)) and (layer3_outputs(1292)));
    layer4_outputs(900) <= not(layer3_outputs(1084)) or (layer3_outputs(652));
    layer4_outputs(901) <= not(layer3_outputs(301)) or (layer3_outputs(1393));
    layer4_outputs(902) <= layer3_outputs(810);
    layer4_outputs(903) <= not((layer3_outputs(1815)) or (layer3_outputs(2382)));
    layer4_outputs(904) <= layer3_outputs(136);
    layer4_outputs(905) <= layer3_outputs(314);
    layer4_outputs(906) <= not((layer3_outputs(1592)) and (layer3_outputs(794)));
    layer4_outputs(907) <= (layer3_outputs(432)) or (layer3_outputs(1763));
    layer4_outputs(908) <= not(layer3_outputs(1881));
    layer4_outputs(909) <= not(layer3_outputs(1531)) or (layer3_outputs(1155));
    layer4_outputs(910) <= layer3_outputs(2490);
    layer4_outputs(911) <= not(layer3_outputs(627)) or (layer3_outputs(1119));
    layer4_outputs(912) <= layer3_outputs(2111);
    layer4_outputs(913) <= layer3_outputs(1233);
    layer4_outputs(914) <= (layer3_outputs(51)) and not (layer3_outputs(1294));
    layer4_outputs(915) <= layer3_outputs(1310);
    layer4_outputs(916) <= not(layer3_outputs(2031));
    layer4_outputs(917) <= not(layer3_outputs(2260));
    layer4_outputs(918) <= not(layer3_outputs(2016));
    layer4_outputs(919) <= layer3_outputs(2375);
    layer4_outputs(920) <= '1';
    layer4_outputs(921) <= '1';
    layer4_outputs(922) <= not((layer3_outputs(584)) or (layer3_outputs(2109)));
    layer4_outputs(923) <= layer3_outputs(294);
    layer4_outputs(924) <= not(layer3_outputs(1661));
    layer4_outputs(925) <= (layer3_outputs(748)) and not (layer3_outputs(312));
    layer4_outputs(926) <= '1';
    layer4_outputs(927) <= not(layer3_outputs(1691));
    layer4_outputs(928) <= not(layer3_outputs(1771));
    layer4_outputs(929) <= not(layer3_outputs(1515));
    layer4_outputs(930) <= not(layer3_outputs(1088));
    layer4_outputs(931) <= (layer3_outputs(1228)) or (layer3_outputs(1855));
    layer4_outputs(932) <= (layer3_outputs(2278)) and not (layer3_outputs(123));
    layer4_outputs(933) <= (layer3_outputs(860)) xor (layer3_outputs(1710));
    layer4_outputs(934) <= (layer3_outputs(638)) or (layer3_outputs(18));
    layer4_outputs(935) <= not((layer3_outputs(1813)) xor (layer3_outputs(2175)));
    layer4_outputs(936) <= (layer3_outputs(2206)) and not (layer3_outputs(1780));
    layer4_outputs(937) <= not(layer3_outputs(727));
    layer4_outputs(938) <= (layer3_outputs(1224)) and not (layer3_outputs(148));
    layer4_outputs(939) <= not(layer3_outputs(2314)) or (layer3_outputs(2346));
    layer4_outputs(940) <= not(layer3_outputs(2415));
    layer4_outputs(941) <= (layer3_outputs(2476)) or (layer3_outputs(701));
    layer4_outputs(942) <= '1';
    layer4_outputs(943) <= (layer3_outputs(1472)) and not (layer3_outputs(2549));
    layer4_outputs(944) <= not(layer3_outputs(2313));
    layer4_outputs(945) <= (layer3_outputs(947)) and (layer3_outputs(1365));
    layer4_outputs(946) <= '1';
    layer4_outputs(947) <= (layer3_outputs(1087)) or (layer3_outputs(1606));
    layer4_outputs(948) <= not((layer3_outputs(29)) and (layer3_outputs(281)));
    layer4_outputs(949) <= not(layer3_outputs(1770));
    layer4_outputs(950) <= not(layer3_outputs(1959));
    layer4_outputs(951) <= not((layer3_outputs(738)) xor (layer3_outputs(1095)));
    layer4_outputs(952) <= '1';
    layer4_outputs(953) <= layer3_outputs(473);
    layer4_outputs(954) <= not(layer3_outputs(1390)) or (layer3_outputs(844));
    layer4_outputs(955) <= not(layer3_outputs(2470));
    layer4_outputs(956) <= layer3_outputs(927);
    layer4_outputs(957) <= (layer3_outputs(1660)) and (layer3_outputs(2024));
    layer4_outputs(958) <= not(layer3_outputs(2)) or (layer3_outputs(1473));
    layer4_outputs(959) <= (layer3_outputs(1607)) or (layer3_outputs(901));
    layer4_outputs(960) <= (layer3_outputs(145)) or (layer3_outputs(886));
    layer4_outputs(961) <= not(layer3_outputs(1186)) or (layer3_outputs(852));
    layer4_outputs(962) <= (layer3_outputs(535)) or (layer3_outputs(292));
    layer4_outputs(963) <= (layer3_outputs(602)) and not (layer3_outputs(318));
    layer4_outputs(964) <= layer3_outputs(1584);
    layer4_outputs(965) <= layer3_outputs(694);
    layer4_outputs(966) <= not(layer3_outputs(1327)) or (layer3_outputs(385));
    layer4_outputs(967) <= layer3_outputs(1999);
    layer4_outputs(968) <= not(layer3_outputs(1836)) or (layer3_outputs(1435));
    layer4_outputs(969) <= not(layer3_outputs(1031)) or (layer3_outputs(1667));
    layer4_outputs(970) <= layer3_outputs(2399);
    layer4_outputs(971) <= not(layer3_outputs(1295));
    layer4_outputs(972) <= not((layer3_outputs(999)) or (layer3_outputs(544)));
    layer4_outputs(973) <= layer3_outputs(2353);
    layer4_outputs(974) <= layer3_outputs(869);
    layer4_outputs(975) <= not(layer3_outputs(2040));
    layer4_outputs(976) <= not(layer3_outputs(1901)) or (layer3_outputs(2405));
    layer4_outputs(977) <= layer3_outputs(467);
    layer4_outputs(978) <= not(layer3_outputs(267));
    layer4_outputs(979) <= layer3_outputs(2299);
    layer4_outputs(980) <= layer3_outputs(1769);
    layer4_outputs(981) <= (layer3_outputs(1806)) and not (layer3_outputs(971));
    layer4_outputs(982) <= (layer3_outputs(1893)) and (layer3_outputs(1900));
    layer4_outputs(983) <= not(layer3_outputs(1472));
    layer4_outputs(984) <= not(layer3_outputs(1497));
    layer4_outputs(985) <= layer3_outputs(2494);
    layer4_outputs(986) <= (layer3_outputs(1614)) or (layer3_outputs(394));
    layer4_outputs(987) <= layer3_outputs(2289);
    layer4_outputs(988) <= layer3_outputs(1662);
    layer4_outputs(989) <= (layer3_outputs(201)) and (layer3_outputs(263));
    layer4_outputs(990) <= (layer3_outputs(1280)) and not (layer3_outputs(695));
    layer4_outputs(991) <= (layer3_outputs(742)) or (layer3_outputs(849));
    layer4_outputs(992) <= (layer3_outputs(1712)) and not (layer3_outputs(1205));
    layer4_outputs(993) <= not((layer3_outputs(423)) and (layer3_outputs(1585)));
    layer4_outputs(994) <= (layer3_outputs(1220)) or (layer3_outputs(2264));
    layer4_outputs(995) <= layer3_outputs(1789);
    layer4_outputs(996) <= not(layer3_outputs(2469));
    layer4_outputs(997) <= layer3_outputs(762);
    layer4_outputs(998) <= not((layer3_outputs(1391)) and (layer3_outputs(376)));
    layer4_outputs(999) <= not(layer3_outputs(913));
    layer4_outputs(1000) <= not(layer3_outputs(222));
    layer4_outputs(1001) <= not(layer3_outputs(1275));
    layer4_outputs(1002) <= not(layer3_outputs(1022));
    layer4_outputs(1003) <= not(layer3_outputs(1097)) or (layer3_outputs(2056));
    layer4_outputs(1004) <= not(layer3_outputs(1021));
    layer4_outputs(1005) <= (layer3_outputs(383)) and not (layer3_outputs(1032));
    layer4_outputs(1006) <= (layer3_outputs(494)) and not (layer3_outputs(1809));
    layer4_outputs(1007) <= not((layer3_outputs(2176)) or (layer3_outputs(1818)));
    layer4_outputs(1008) <= not((layer3_outputs(1308)) or (layer3_outputs(1373)));
    layer4_outputs(1009) <= layer3_outputs(513);
    layer4_outputs(1010) <= not(layer3_outputs(1986)) or (layer3_outputs(291));
    layer4_outputs(1011) <= '0';
    layer4_outputs(1012) <= (layer3_outputs(2148)) or (layer3_outputs(2166));
    layer4_outputs(1013) <= (layer3_outputs(1343)) and (layer3_outputs(2390));
    layer4_outputs(1014) <= (layer3_outputs(1145)) or (layer3_outputs(57));
    layer4_outputs(1015) <= layer3_outputs(1439);
    layer4_outputs(1016) <= (layer3_outputs(269)) and not (layer3_outputs(2393));
    layer4_outputs(1017) <= not(layer3_outputs(486));
    layer4_outputs(1018) <= '0';
    layer4_outputs(1019) <= not(layer3_outputs(854));
    layer4_outputs(1020) <= '0';
    layer4_outputs(1021) <= not(layer3_outputs(920)) or (layer3_outputs(1537));
    layer4_outputs(1022) <= not(layer3_outputs(565));
    layer4_outputs(1023) <= (layer3_outputs(653)) or (layer3_outputs(167));
    layer4_outputs(1024) <= (layer3_outputs(2104)) and (layer3_outputs(1846));
    layer4_outputs(1025) <= layer3_outputs(2330);
    layer4_outputs(1026) <= layer3_outputs(2554);
    layer4_outputs(1027) <= layer3_outputs(2361);
    layer4_outputs(1028) <= (layer3_outputs(2401)) and not (layer3_outputs(193));
    layer4_outputs(1029) <= not(layer3_outputs(2458));
    layer4_outputs(1030) <= layer3_outputs(1800);
    layer4_outputs(1031) <= '1';
    layer4_outputs(1032) <= (layer3_outputs(711)) and not (layer3_outputs(1067));
    layer4_outputs(1033) <= '1';
    layer4_outputs(1034) <= not(layer3_outputs(219));
    layer4_outputs(1035) <= not(layer3_outputs(2142));
    layer4_outputs(1036) <= layer3_outputs(1747);
    layer4_outputs(1037) <= not(layer3_outputs(1621));
    layer4_outputs(1038) <= not(layer3_outputs(1252)) or (layer3_outputs(1318));
    layer4_outputs(1039) <= (layer3_outputs(2407)) and (layer3_outputs(1937));
    layer4_outputs(1040) <= not(layer3_outputs(271));
    layer4_outputs(1041) <= not(layer3_outputs(1977)) or (layer3_outputs(1824));
    layer4_outputs(1042) <= (layer3_outputs(806)) and not (layer3_outputs(2159));
    layer4_outputs(1043) <= layer3_outputs(700);
    layer4_outputs(1044) <= '1';
    layer4_outputs(1045) <= not(layer3_outputs(731));
    layer4_outputs(1046) <= layer3_outputs(706);
    layer4_outputs(1047) <= layer3_outputs(755);
    layer4_outputs(1048) <= (layer3_outputs(776)) or (layer3_outputs(1121));
    layer4_outputs(1049) <= not(layer3_outputs(2300)) or (layer3_outputs(1159));
    layer4_outputs(1050) <= (layer3_outputs(271)) or (layer3_outputs(1171));
    layer4_outputs(1051) <= not(layer3_outputs(163)) or (layer3_outputs(1367));
    layer4_outputs(1052) <= layer3_outputs(2509);
    layer4_outputs(1053) <= layer3_outputs(1734);
    layer4_outputs(1054) <= layer3_outputs(1173);
    layer4_outputs(1055) <= layer3_outputs(1564);
    layer4_outputs(1056) <= (layer3_outputs(2103)) or (layer3_outputs(814));
    layer4_outputs(1057) <= (layer3_outputs(2463)) and not (layer3_outputs(956));
    layer4_outputs(1058) <= layer3_outputs(2041);
    layer4_outputs(1059) <= not(layer3_outputs(953));
    layer4_outputs(1060) <= not(layer3_outputs(1621));
    layer4_outputs(1061) <= not(layer3_outputs(1586));
    layer4_outputs(1062) <= not(layer3_outputs(1453));
    layer4_outputs(1063) <= not(layer3_outputs(29)) or (layer3_outputs(2027));
    layer4_outputs(1064) <= (layer3_outputs(1714)) or (layer3_outputs(2469));
    layer4_outputs(1065) <= '0';
    layer4_outputs(1066) <= (layer3_outputs(2303)) and not (layer3_outputs(216));
    layer4_outputs(1067) <= not(layer3_outputs(1735));
    layer4_outputs(1068) <= layer3_outputs(1889);
    layer4_outputs(1069) <= layer3_outputs(2000);
    layer4_outputs(1070) <= (layer3_outputs(836)) and not (layer3_outputs(397));
    layer4_outputs(1071) <= '0';
    layer4_outputs(1072) <= not(layer3_outputs(1221));
    layer4_outputs(1073) <= not(layer3_outputs(1648)) or (layer3_outputs(1185));
    layer4_outputs(1074) <= layer3_outputs(1193);
    layer4_outputs(1075) <= (layer3_outputs(634)) and not (layer3_outputs(1423));
    layer4_outputs(1076) <= layer3_outputs(1845);
    layer4_outputs(1077) <= (layer3_outputs(1989)) and not (layer3_outputs(2498));
    layer4_outputs(1078) <= not(layer3_outputs(2448));
    layer4_outputs(1079) <= not(layer3_outputs(245));
    layer4_outputs(1080) <= not((layer3_outputs(1474)) and (layer3_outputs(2052)));
    layer4_outputs(1081) <= layer3_outputs(1339);
    layer4_outputs(1082) <= '0';
    layer4_outputs(1083) <= '0';
    layer4_outputs(1084) <= layer3_outputs(1505);
    layer4_outputs(1085) <= layer3_outputs(1758);
    layer4_outputs(1086) <= not(layer3_outputs(395));
    layer4_outputs(1087) <= not(layer3_outputs(1484));
    layer4_outputs(1088) <= not((layer3_outputs(1047)) xor (layer3_outputs(1927)));
    layer4_outputs(1089) <= '1';
    layer4_outputs(1090) <= '0';
    layer4_outputs(1091) <= not(layer3_outputs(503));
    layer4_outputs(1092) <= (layer3_outputs(546)) and not (layer3_outputs(27));
    layer4_outputs(1093) <= not((layer3_outputs(963)) and (layer3_outputs(738)));
    layer4_outputs(1094) <= '1';
    layer4_outputs(1095) <= (layer3_outputs(2046)) or (layer3_outputs(199));
    layer4_outputs(1096) <= not((layer3_outputs(1597)) and (layer3_outputs(1477)));
    layer4_outputs(1097) <= not(layer3_outputs(1754));
    layer4_outputs(1098) <= layer3_outputs(570);
    layer4_outputs(1099) <= not(layer3_outputs(1988));
    layer4_outputs(1100) <= layer3_outputs(315);
    layer4_outputs(1101) <= (layer3_outputs(2489)) and (layer3_outputs(1762));
    layer4_outputs(1102) <= '1';
    layer4_outputs(1103) <= (layer3_outputs(925)) and not (layer3_outputs(2136));
    layer4_outputs(1104) <= (layer3_outputs(409)) or (layer3_outputs(607));
    layer4_outputs(1105) <= not(layer3_outputs(2557));
    layer4_outputs(1106) <= (layer3_outputs(2222)) and not (layer3_outputs(1153));
    layer4_outputs(1107) <= not(layer3_outputs(403));
    layer4_outputs(1108) <= not((layer3_outputs(1562)) or (layer3_outputs(822)));
    layer4_outputs(1109) <= not(layer3_outputs(2018));
    layer4_outputs(1110) <= not(layer3_outputs(658));
    layer4_outputs(1111) <= not(layer3_outputs(1999));
    layer4_outputs(1112) <= '0';
    layer4_outputs(1113) <= (layer3_outputs(1867)) or (layer3_outputs(838));
    layer4_outputs(1114) <= not(layer3_outputs(588)) or (layer3_outputs(1827));
    layer4_outputs(1115) <= not(layer3_outputs(317)) or (layer3_outputs(365));
    layer4_outputs(1116) <= layer3_outputs(1749);
    layer4_outputs(1117) <= (layer3_outputs(1708)) and (layer3_outputs(632));
    layer4_outputs(1118) <= (layer3_outputs(867)) or (layer3_outputs(1281));
    layer4_outputs(1119) <= not((layer3_outputs(2383)) or (layer3_outputs(1302)));
    layer4_outputs(1120) <= (layer3_outputs(60)) or (layer3_outputs(195));
    layer4_outputs(1121) <= layer3_outputs(2177);
    layer4_outputs(1122) <= layer3_outputs(1293);
    layer4_outputs(1123) <= not((layer3_outputs(2180)) or (layer3_outputs(199)));
    layer4_outputs(1124) <= not(layer3_outputs(1331));
    layer4_outputs(1125) <= '0';
    layer4_outputs(1126) <= not(layer3_outputs(456));
    layer4_outputs(1127) <= not(layer3_outputs(1954));
    layer4_outputs(1128) <= '0';
    layer4_outputs(1129) <= layer3_outputs(1287);
    layer4_outputs(1130) <= (layer3_outputs(1784)) and (layer3_outputs(1031));
    layer4_outputs(1131) <= (layer3_outputs(941)) and not (layer3_outputs(2066));
    layer4_outputs(1132) <= layer3_outputs(491);
    layer4_outputs(1133) <= '1';
    layer4_outputs(1134) <= '0';
    layer4_outputs(1135) <= not(layer3_outputs(337));
    layer4_outputs(1136) <= not(layer3_outputs(1094));
    layer4_outputs(1137) <= not((layer3_outputs(6)) or (layer3_outputs(670)));
    layer4_outputs(1138) <= '1';
    layer4_outputs(1139) <= (layer3_outputs(698)) xor (layer3_outputs(1475));
    layer4_outputs(1140) <= (layer3_outputs(1774)) xor (layer3_outputs(465));
    layer4_outputs(1141) <= not(layer3_outputs(1055)) or (layer3_outputs(1866));
    layer4_outputs(1142) <= (layer3_outputs(95)) and (layer3_outputs(312));
    layer4_outputs(1143) <= not(layer3_outputs(2371)) or (layer3_outputs(498));
    layer4_outputs(1144) <= not(layer3_outputs(1407)) or (layer3_outputs(1967));
    layer4_outputs(1145) <= '0';
    layer4_outputs(1146) <= not(layer3_outputs(1665));
    layer4_outputs(1147) <= (layer3_outputs(512)) and not (layer3_outputs(694));
    layer4_outputs(1148) <= layer3_outputs(2054);
    layer4_outputs(1149) <= (layer3_outputs(858)) xor (layer3_outputs(1513));
    layer4_outputs(1150) <= '0';
    layer4_outputs(1151) <= '0';
    layer4_outputs(1152) <= layer3_outputs(440);
    layer4_outputs(1153) <= not((layer3_outputs(1412)) and (layer3_outputs(1362)));
    layer4_outputs(1154) <= not(layer3_outputs(2227));
    layer4_outputs(1155) <= not(layer3_outputs(1220));
    layer4_outputs(1156) <= (layer3_outputs(254)) and (layer3_outputs(2327));
    layer4_outputs(1157) <= (layer3_outputs(1850)) and not (layer3_outputs(2330));
    layer4_outputs(1158) <= layer3_outputs(883);
    layer4_outputs(1159) <= layer3_outputs(2373);
    layer4_outputs(1160) <= not(layer3_outputs(795));
    layer4_outputs(1161) <= '0';
    layer4_outputs(1162) <= (layer3_outputs(1896)) and not (layer3_outputs(419));
    layer4_outputs(1163) <= not((layer3_outputs(163)) and (layer3_outputs(2256)));
    layer4_outputs(1164) <= not(layer3_outputs(730)) or (layer3_outputs(2154));
    layer4_outputs(1165) <= '0';
    layer4_outputs(1166) <= layer3_outputs(2464);
    layer4_outputs(1167) <= not(layer3_outputs(1671));
    layer4_outputs(1168) <= layer3_outputs(11);
    layer4_outputs(1169) <= not(layer3_outputs(1417));
    layer4_outputs(1170) <= not((layer3_outputs(633)) and (layer3_outputs(139)));
    layer4_outputs(1171) <= (layer3_outputs(775)) and (layer3_outputs(1857));
    layer4_outputs(1172) <= not(layer3_outputs(1138));
    layer4_outputs(1173) <= not(layer3_outputs(2164));
    layer4_outputs(1174) <= (layer3_outputs(1256)) or (layer3_outputs(2020));
    layer4_outputs(1175) <= layer3_outputs(2048);
    layer4_outputs(1176) <= not(layer3_outputs(1883));
    layer4_outputs(1177) <= layer3_outputs(2236);
    layer4_outputs(1178) <= (layer3_outputs(613)) and (layer3_outputs(319));
    layer4_outputs(1179) <= layer3_outputs(1309);
    layer4_outputs(1180) <= layer3_outputs(399);
    layer4_outputs(1181) <= not(layer3_outputs(590));
    layer4_outputs(1182) <= not((layer3_outputs(1848)) and (layer3_outputs(865)));
    layer4_outputs(1183) <= layer3_outputs(1970);
    layer4_outputs(1184) <= not((layer3_outputs(1989)) or (layer3_outputs(556)));
    layer4_outputs(1185) <= layer3_outputs(485);
    layer4_outputs(1186) <= (layer3_outputs(2386)) and not (layer3_outputs(2552));
    layer4_outputs(1187) <= not(layer3_outputs(2304)) or (layer3_outputs(1973));
    layer4_outputs(1188) <= not((layer3_outputs(564)) xor (layer3_outputs(381)));
    layer4_outputs(1189) <= not((layer3_outputs(535)) and (layer3_outputs(1902)));
    layer4_outputs(1190) <= (layer3_outputs(1230)) or (layer3_outputs(1414));
    layer4_outputs(1191) <= not(layer3_outputs(1241));
    layer4_outputs(1192) <= layer3_outputs(2295);
    layer4_outputs(1193) <= layer3_outputs(1891);
    layer4_outputs(1194) <= not(layer3_outputs(2437));
    layer4_outputs(1195) <= layer3_outputs(1340);
    layer4_outputs(1196) <= layer3_outputs(436);
    layer4_outputs(1197) <= (layer3_outputs(2115)) xor (layer3_outputs(926));
    layer4_outputs(1198) <= layer3_outputs(11);
    layer4_outputs(1199) <= '1';
    layer4_outputs(1200) <= not(layer3_outputs(316)) or (layer3_outputs(333));
    layer4_outputs(1201) <= not(layer3_outputs(189)) or (layer3_outputs(416));
    layer4_outputs(1202) <= (layer3_outputs(214)) or (layer3_outputs(1991));
    layer4_outputs(1203) <= not(layer3_outputs(2516)) or (layer3_outputs(1043));
    layer4_outputs(1204) <= layer3_outputs(2246);
    layer4_outputs(1205) <= layer3_outputs(1597);
    layer4_outputs(1206) <= layer3_outputs(1086);
    layer4_outputs(1207) <= '1';
    layer4_outputs(1208) <= layer3_outputs(2382);
    layer4_outputs(1209) <= layer3_outputs(739);
    layer4_outputs(1210) <= not((layer3_outputs(324)) and (layer3_outputs(1172)));
    layer4_outputs(1211) <= not(layer3_outputs(2479));
    layer4_outputs(1212) <= not(layer3_outputs(388));
    layer4_outputs(1213) <= not(layer3_outputs(889)) or (layer3_outputs(1436));
    layer4_outputs(1214) <= (layer3_outputs(1619)) and not (layer3_outputs(570));
    layer4_outputs(1215) <= not(layer3_outputs(334));
    layer4_outputs(1216) <= not((layer3_outputs(764)) xor (layer3_outputs(1146)));
    layer4_outputs(1217) <= not((layer3_outputs(1286)) or (layer3_outputs(713)));
    layer4_outputs(1218) <= not((layer3_outputs(2033)) and (layer3_outputs(1122)));
    layer4_outputs(1219) <= (layer3_outputs(1573)) and (layer3_outputs(2335));
    layer4_outputs(1220) <= not(layer3_outputs(1082));
    layer4_outputs(1221) <= layer3_outputs(1461);
    layer4_outputs(1222) <= '1';
    layer4_outputs(1223) <= layer3_outputs(1812);
    layer4_outputs(1224) <= (layer3_outputs(1434)) and not (layer3_outputs(87));
    layer4_outputs(1225) <= not(layer3_outputs(2245)) or (layer3_outputs(1279));
    layer4_outputs(1226) <= (layer3_outputs(749)) and not (layer3_outputs(1974));
    layer4_outputs(1227) <= not((layer3_outputs(2406)) or (layer3_outputs(1446)));
    layer4_outputs(1228) <= layer3_outputs(482);
    layer4_outputs(1229) <= (layer3_outputs(2420)) or (layer3_outputs(1201));
    layer4_outputs(1230) <= '1';
    layer4_outputs(1231) <= layer3_outputs(133);
    layer4_outputs(1232) <= not(layer3_outputs(1772));
    layer4_outputs(1233) <= '0';
    layer4_outputs(1234) <= (layer3_outputs(771)) and not (layer3_outputs(1131));
    layer4_outputs(1235) <= (layer3_outputs(1036)) or (layer3_outputs(951));
    layer4_outputs(1236) <= not((layer3_outputs(1641)) and (layer3_outputs(2466)));
    layer4_outputs(1237) <= (layer3_outputs(1558)) or (layer3_outputs(1988));
    layer4_outputs(1238) <= '0';
    layer4_outputs(1239) <= layer3_outputs(2014);
    layer4_outputs(1240) <= (layer3_outputs(1723)) and (layer3_outputs(890));
    layer4_outputs(1241) <= not(layer3_outputs(2152)) or (layer3_outputs(981));
    layer4_outputs(1242) <= not(layer3_outputs(2424));
    layer4_outputs(1243) <= not((layer3_outputs(1617)) or (layer3_outputs(328)));
    layer4_outputs(1244) <= not(layer3_outputs(1352)) or (layer3_outputs(945));
    layer4_outputs(1245) <= (layer3_outputs(1552)) xor (layer3_outputs(2432));
    layer4_outputs(1246) <= layer3_outputs(1008);
    layer4_outputs(1247) <= not(layer3_outputs(914));
    layer4_outputs(1248) <= layer3_outputs(2009);
    layer4_outputs(1249) <= '1';
    layer4_outputs(1250) <= not(layer3_outputs(1658));
    layer4_outputs(1251) <= (layer3_outputs(818)) and not (layer3_outputs(1525));
    layer4_outputs(1252) <= layer3_outputs(1019);
    layer4_outputs(1253) <= layer3_outputs(1023);
    layer4_outputs(1254) <= not((layer3_outputs(1190)) or (layer3_outputs(891)));
    layer4_outputs(1255) <= '1';
    layer4_outputs(1256) <= layer3_outputs(2153);
    layer4_outputs(1257) <= layer3_outputs(1136);
    layer4_outputs(1258) <= not(layer3_outputs(2380)) or (layer3_outputs(563));
    layer4_outputs(1259) <= not(layer3_outputs(443));
    layer4_outputs(1260) <= (layer3_outputs(2318)) or (layer3_outputs(164));
    layer4_outputs(1261) <= not(layer3_outputs(2438));
    layer4_outputs(1262) <= layer3_outputs(2473);
    layer4_outputs(1263) <= (layer3_outputs(35)) xor (layer3_outputs(530));
    layer4_outputs(1264) <= not(layer3_outputs(1646));
    layer4_outputs(1265) <= (layer3_outputs(1968)) and not (layer3_outputs(204));
    layer4_outputs(1266) <= not((layer3_outputs(410)) and (layer3_outputs(714)));
    layer4_outputs(1267) <= not(layer3_outputs(1247));
    layer4_outputs(1268) <= '1';
    layer4_outputs(1269) <= not(layer3_outputs(780)) or (layer3_outputs(1637));
    layer4_outputs(1270) <= not(layer3_outputs(1634));
    layer4_outputs(1271) <= (layer3_outputs(22)) and (layer3_outputs(2412));
    layer4_outputs(1272) <= not(layer3_outputs(2131));
    layer4_outputs(1273) <= not(layer3_outputs(207));
    layer4_outputs(1274) <= (layer3_outputs(218)) and not (layer3_outputs(1992));
    layer4_outputs(1275) <= not((layer3_outputs(1341)) or (layer3_outputs(597)));
    layer4_outputs(1276) <= '1';
    layer4_outputs(1277) <= not((layer3_outputs(2553)) and (layer3_outputs(1273)));
    layer4_outputs(1278) <= not(layer3_outputs(319)) or (layer3_outputs(47));
    layer4_outputs(1279) <= not(layer3_outputs(1970));
    layer4_outputs(1280) <= not(layer3_outputs(650)) or (layer3_outputs(1860));
    layer4_outputs(1281) <= '1';
    layer4_outputs(1282) <= not(layer3_outputs(1080)) or (layer3_outputs(123));
    layer4_outputs(1283) <= layer3_outputs(2418);
    layer4_outputs(1284) <= (layer3_outputs(1978)) and (layer3_outputs(387));
    layer4_outputs(1285) <= layer3_outputs(190);
    layer4_outputs(1286) <= not(layer3_outputs(1095));
    layer4_outputs(1287) <= not((layer3_outputs(1252)) or (layer3_outputs(2207)));
    layer4_outputs(1288) <= (layer3_outputs(2214)) or (layer3_outputs(55));
    layer4_outputs(1289) <= layer3_outputs(2465);
    layer4_outputs(1290) <= (layer3_outputs(2193)) and not (layer3_outputs(1489));
    layer4_outputs(1291) <= (layer3_outputs(278)) and (layer3_outputs(891));
    layer4_outputs(1292) <= not(layer3_outputs(70));
    layer4_outputs(1293) <= layer3_outputs(361);
    layer4_outputs(1294) <= layer3_outputs(1224);
    layer4_outputs(1295) <= not((layer3_outputs(309)) and (layer3_outputs(277)));
    layer4_outputs(1296) <= '1';
    layer4_outputs(1297) <= not(layer3_outputs(265)) or (layer3_outputs(83));
    layer4_outputs(1298) <= not((layer3_outputs(1955)) or (layer3_outputs(143)));
    layer4_outputs(1299) <= (layer3_outputs(2412)) or (layer3_outputs(863));
    layer4_outputs(1300) <= not(layer3_outputs(727));
    layer4_outputs(1301) <= not((layer3_outputs(1668)) or (layer3_outputs(784)));
    layer4_outputs(1302) <= layer3_outputs(1314);
    layer4_outputs(1303) <= '1';
    layer4_outputs(1304) <= layer3_outputs(934);
    layer4_outputs(1305) <= layer3_outputs(2291);
    layer4_outputs(1306) <= not(layer3_outputs(2183)) or (layer3_outputs(2488));
    layer4_outputs(1307) <= not(layer3_outputs(734));
    layer4_outputs(1308) <= (layer3_outputs(1752)) and not (layer3_outputs(654));
    layer4_outputs(1309) <= layer3_outputs(834);
    layer4_outputs(1310) <= not(layer3_outputs(1339));
    layer4_outputs(1311) <= not((layer3_outputs(726)) or (layer3_outputs(1035)));
    layer4_outputs(1312) <= not(layer3_outputs(2203));
    layer4_outputs(1313) <= layer3_outputs(575);
    layer4_outputs(1314) <= (layer3_outputs(1014)) or (layer3_outputs(1650));
    layer4_outputs(1315) <= (layer3_outputs(1123)) and (layer3_outputs(509));
    layer4_outputs(1316) <= not((layer3_outputs(1005)) or (layer3_outputs(50)));
    layer4_outputs(1317) <= layer3_outputs(523);
    layer4_outputs(1318) <= not(layer3_outputs(294)) or (layer3_outputs(974));
    layer4_outputs(1319) <= layer3_outputs(1998);
    layer4_outputs(1320) <= not(layer3_outputs(961));
    layer4_outputs(1321) <= (layer3_outputs(1534)) and not (layer3_outputs(791));
    layer4_outputs(1322) <= layer3_outputs(444);
    layer4_outputs(1323) <= (layer3_outputs(890)) and not (layer3_outputs(737));
    layer4_outputs(1324) <= (layer3_outputs(1163)) and not (layer3_outputs(702));
    layer4_outputs(1325) <= not(layer3_outputs(2204));
    layer4_outputs(1326) <= (layer3_outputs(76)) or (layer3_outputs(1511));
    layer4_outputs(1327) <= not(layer3_outputs(1788));
    layer4_outputs(1328) <= layer3_outputs(2194);
    layer4_outputs(1329) <= not(layer3_outputs(82));
    layer4_outputs(1330) <= (layer3_outputs(1467)) or (layer3_outputs(59));
    layer4_outputs(1331) <= layer3_outputs(2301);
    layer4_outputs(1332) <= '0';
    layer4_outputs(1333) <= (layer3_outputs(532)) or (layer3_outputs(283));
    layer4_outputs(1334) <= (layer3_outputs(1912)) xor (layer3_outputs(1906));
    layer4_outputs(1335) <= (layer3_outputs(2362)) or (layer3_outputs(2069));
    layer4_outputs(1336) <= layer3_outputs(2107);
    layer4_outputs(1337) <= not(layer3_outputs(1042)) or (layer3_outputs(2034));
    layer4_outputs(1338) <= not((layer3_outputs(210)) or (layer3_outputs(615)));
    layer4_outputs(1339) <= '0';
    layer4_outputs(1340) <= (layer3_outputs(1002)) and (layer3_outputs(883));
    layer4_outputs(1341) <= layer3_outputs(718);
    layer4_outputs(1342) <= (layer3_outputs(2495)) and (layer3_outputs(2549));
    layer4_outputs(1343) <= not(layer3_outputs(2237));
    layer4_outputs(1344) <= layer3_outputs(2001);
    layer4_outputs(1345) <= layer3_outputs(2012);
    layer4_outputs(1346) <= not(layer3_outputs(665));
    layer4_outputs(1347) <= not(layer3_outputs(151));
    layer4_outputs(1348) <= not(layer3_outputs(677));
    layer4_outputs(1349) <= not(layer3_outputs(1403)) or (layer3_outputs(1256));
    layer4_outputs(1350) <= not(layer3_outputs(1754)) or (layer3_outputs(1452));
    layer4_outputs(1351) <= not(layer3_outputs(179)) or (layer3_outputs(391));
    layer4_outputs(1352) <= not(layer3_outputs(2339)) or (layer3_outputs(1328));
    layer4_outputs(1353) <= not((layer3_outputs(983)) and (layer3_outputs(2303)));
    layer4_outputs(1354) <= not(layer3_outputs(3));
    layer4_outputs(1355) <= not(layer3_outputs(2430));
    layer4_outputs(1356) <= '1';
    layer4_outputs(1357) <= layer3_outputs(2452);
    layer4_outputs(1358) <= not(layer3_outputs(293));
    layer4_outputs(1359) <= (layer3_outputs(847)) and not (layer3_outputs(611));
    layer4_outputs(1360) <= not(layer3_outputs(1915));
    layer4_outputs(1361) <= (layer3_outputs(1458)) xor (layer3_outputs(871));
    layer4_outputs(1362) <= layer3_outputs(2154);
    layer4_outputs(1363) <= not(layer3_outputs(579));
    layer4_outputs(1364) <= not((layer3_outputs(733)) or (layer3_outputs(350)));
    layer4_outputs(1365) <= (layer3_outputs(1572)) xor (layer3_outputs(2544));
    layer4_outputs(1366) <= layer3_outputs(1947);
    layer4_outputs(1367) <= (layer3_outputs(1815)) or (layer3_outputs(1058));
    layer4_outputs(1368) <= layer3_outputs(81);
    layer4_outputs(1369) <= (layer3_outputs(872)) or (layer3_outputs(1003));
    layer4_outputs(1370) <= not(layer3_outputs(179));
    layer4_outputs(1371) <= not(layer3_outputs(990)) or (layer3_outputs(595));
    layer4_outputs(1372) <= '0';
    layer4_outputs(1373) <= (layer3_outputs(596)) or (layer3_outputs(1768));
    layer4_outputs(1374) <= not(layer3_outputs(1524));
    layer4_outputs(1375) <= (layer3_outputs(1062)) and (layer3_outputs(161));
    layer4_outputs(1376) <= not(layer3_outputs(521)) or (layer3_outputs(453));
    layer4_outputs(1377) <= not(layer3_outputs(1971));
    layer4_outputs(1378) <= layer3_outputs(2163);
    layer4_outputs(1379) <= not(layer3_outputs(129)) or (layer3_outputs(320));
    layer4_outputs(1380) <= not(layer3_outputs(1171));
    layer4_outputs(1381) <= layer3_outputs(2170);
    layer4_outputs(1382) <= layer3_outputs(1116);
    layer4_outputs(1383) <= layer3_outputs(1237);
    layer4_outputs(1384) <= not((layer3_outputs(526)) or (layer3_outputs(2063)));
    layer4_outputs(1385) <= '1';
    layer4_outputs(1386) <= not(layer3_outputs(323));
    layer4_outputs(1387) <= not((layer3_outputs(1833)) and (layer3_outputs(2281)));
    layer4_outputs(1388) <= layer3_outputs(2340);
    layer4_outputs(1389) <= layer3_outputs(1271);
    layer4_outputs(1390) <= layer3_outputs(2200);
    layer4_outputs(1391) <= '1';
    layer4_outputs(1392) <= not(layer3_outputs(343));
    layer4_outputs(1393) <= (layer3_outputs(2383)) or (layer3_outputs(2485));
    layer4_outputs(1394) <= (layer3_outputs(182)) or (layer3_outputs(115));
    layer4_outputs(1395) <= not(layer3_outputs(450)) or (layer3_outputs(1732));
    layer4_outputs(1396) <= (layer3_outputs(2287)) or (layer3_outputs(2464));
    layer4_outputs(1397) <= not(layer3_outputs(1001));
    layer4_outputs(1398) <= not(layer3_outputs(1108)) or (layer3_outputs(1221));
    layer4_outputs(1399) <= (layer3_outputs(2445)) and not (layer3_outputs(1767));
    layer4_outputs(1400) <= not((layer3_outputs(662)) and (layer3_outputs(2437)));
    layer4_outputs(1401) <= '0';
    layer4_outputs(1402) <= not(layer3_outputs(1878));
    layer4_outputs(1403) <= not(layer3_outputs(336));
    layer4_outputs(1404) <= layer3_outputs(1536);
    layer4_outputs(1405) <= not((layer3_outputs(516)) or (layer3_outputs(1307)));
    layer4_outputs(1406) <= (layer3_outputs(1779)) and not (layer3_outputs(449));
    layer4_outputs(1407) <= not(layer3_outputs(812));
    layer4_outputs(1408) <= (layer3_outputs(1431)) or (layer3_outputs(302));
    layer4_outputs(1409) <= (layer3_outputs(2247)) and (layer3_outputs(1510));
    layer4_outputs(1410) <= not(layer3_outputs(916));
    layer4_outputs(1411) <= not(layer3_outputs(1913));
    layer4_outputs(1412) <= not((layer3_outputs(2144)) or (layer3_outputs(65)));
    layer4_outputs(1413) <= not((layer3_outputs(977)) and (layer3_outputs(2297)));
    layer4_outputs(1414) <= layer3_outputs(2453);
    layer4_outputs(1415) <= layer3_outputs(1636);
    layer4_outputs(1416) <= not(layer3_outputs(128));
    layer4_outputs(1417) <= not(layer3_outputs(578)) or (layer3_outputs(2073));
    layer4_outputs(1418) <= (layer3_outputs(2388)) or (layer3_outputs(2355));
    layer4_outputs(1419) <= (layer3_outputs(2157)) and not (layer3_outputs(591));
    layer4_outputs(1420) <= (layer3_outputs(1153)) or (layer3_outputs(2370));
    layer4_outputs(1421) <= (layer3_outputs(1847)) and not (layer3_outputs(1496));
    layer4_outputs(1422) <= not(layer3_outputs(536));
    layer4_outputs(1423) <= (layer3_outputs(103)) xor (layer3_outputs(1392));
    layer4_outputs(1424) <= layer3_outputs(212);
    layer4_outputs(1425) <= layer3_outputs(1919);
    layer4_outputs(1426) <= (layer3_outputs(2307)) or (layer3_outputs(1352));
    layer4_outputs(1427) <= not(layer3_outputs(769));
    layer4_outputs(1428) <= layer3_outputs(120);
    layer4_outputs(1429) <= (layer3_outputs(8)) and not (layer3_outputs(974));
    layer4_outputs(1430) <= not(layer3_outputs(729));
    layer4_outputs(1431) <= layer3_outputs(2092);
    layer4_outputs(1432) <= layer3_outputs(1672);
    layer4_outputs(1433) <= layer3_outputs(1332);
    layer4_outputs(1434) <= not(layer3_outputs(2122));
    layer4_outputs(1435) <= (layer3_outputs(377)) or (layer3_outputs(852));
    layer4_outputs(1436) <= (layer3_outputs(115)) and not (layer3_outputs(88));
    layer4_outputs(1437) <= not((layer3_outputs(1128)) or (layer3_outputs(1842)));
    layer4_outputs(1438) <= not(layer3_outputs(1516));
    layer4_outputs(1439) <= not(layer3_outputs(2077)) or (layer3_outputs(1187));
    layer4_outputs(1440) <= (layer3_outputs(2191)) and not (layer3_outputs(2006));
    layer4_outputs(1441) <= not((layer3_outputs(2357)) or (layer3_outputs(1600)));
    layer4_outputs(1442) <= not((layer3_outputs(2328)) and (layer3_outputs(1972)));
    layer4_outputs(1443) <= not(layer3_outputs(2243));
    layer4_outputs(1444) <= (layer3_outputs(1315)) and (layer3_outputs(2165));
    layer4_outputs(1445) <= not(layer3_outputs(1193));
    layer4_outputs(1446) <= layer3_outputs(671);
    layer4_outputs(1447) <= (layer3_outputs(648)) and not (layer3_outputs(2273));
    layer4_outputs(1448) <= not(layer3_outputs(2295));
    layer4_outputs(1449) <= layer3_outputs(1508);
    layer4_outputs(1450) <= layer3_outputs(1538);
    layer4_outputs(1451) <= not(layer3_outputs(512));
    layer4_outputs(1452) <= layer3_outputs(2111);
    layer4_outputs(1453) <= not(layer3_outputs(894));
    layer4_outputs(1454) <= layer3_outputs(2075);
    layer4_outputs(1455) <= layer3_outputs(1265);
    layer4_outputs(1456) <= not(layer3_outputs(1872));
    layer4_outputs(1457) <= (layer3_outputs(655)) or (layer3_outputs(503));
    layer4_outputs(1458) <= not(layer3_outputs(268));
    layer4_outputs(1459) <= layer3_outputs(354);
    layer4_outputs(1460) <= not(layer3_outputs(1581));
    layer4_outputs(1461) <= not(layer3_outputs(176));
    layer4_outputs(1462) <= (layer3_outputs(1916)) or (layer3_outputs(1259));
    layer4_outputs(1463) <= layer3_outputs(1052);
    layer4_outputs(1464) <= not((layer3_outputs(468)) or (layer3_outputs(2543)));
    layer4_outputs(1465) <= not(layer3_outputs(1961));
    layer4_outputs(1466) <= not((layer3_outputs(2131)) and (layer3_outputs(144)));
    layer4_outputs(1467) <= not(layer3_outputs(1743)) or (layer3_outputs(1590));
    layer4_outputs(1468) <= layer3_outputs(1052);
    layer4_outputs(1469) <= layer3_outputs(390);
    layer4_outputs(1470) <= '1';
    layer4_outputs(1471) <= layer3_outputs(1071);
    layer4_outputs(1472) <= layer3_outputs(2369);
    layer4_outputs(1473) <= not(layer3_outputs(697));
    layer4_outputs(1474) <= not(layer3_outputs(1546));
    layer4_outputs(1475) <= (layer3_outputs(1903)) xor (layer3_outputs(1834));
    layer4_outputs(1476) <= not(layer3_outputs(1157));
    layer4_outputs(1477) <= not(layer3_outputs(488));
    layer4_outputs(1478) <= (layer3_outputs(173)) xor (layer3_outputs(2493));
    layer4_outputs(1479) <= not(layer3_outputs(2403));
    layer4_outputs(1480) <= layer3_outputs(1703);
    layer4_outputs(1481) <= not((layer3_outputs(259)) xor (layer3_outputs(2499)));
    layer4_outputs(1482) <= not((layer3_outputs(1668)) and (layer3_outputs(2090)));
    layer4_outputs(1483) <= (layer3_outputs(1766)) xor (layer3_outputs(1023));
    layer4_outputs(1484) <= (layer3_outputs(538)) and not (layer3_outputs(732));
    layer4_outputs(1485) <= (layer3_outputs(2060)) and not (layer3_outputs(2006));
    layer4_outputs(1486) <= not(layer3_outputs(1225));
    layer4_outputs(1487) <= not((layer3_outputs(1258)) and (layer3_outputs(1913)));
    layer4_outputs(1488) <= (layer3_outputs(2133)) xor (layer3_outputs(1194));
    layer4_outputs(1489) <= layer3_outputs(1438);
    layer4_outputs(1490) <= (layer3_outputs(2521)) and not (layer3_outputs(832));
    layer4_outputs(1491) <= not(layer3_outputs(2323));
    layer4_outputs(1492) <= layer3_outputs(1622);
    layer4_outputs(1493) <= layer3_outputs(175);
    layer4_outputs(1494) <= '0';
    layer4_outputs(1495) <= not(layer3_outputs(509));
    layer4_outputs(1496) <= layer3_outputs(1897);
    layer4_outputs(1497) <= '0';
    layer4_outputs(1498) <= not(layer3_outputs(733));
    layer4_outputs(1499) <= (layer3_outputs(2231)) xor (layer3_outputs(2279));
    layer4_outputs(1500) <= '1';
    layer4_outputs(1501) <= layer3_outputs(728);
    layer4_outputs(1502) <= not(layer3_outputs(603));
    layer4_outputs(1503) <= (layer3_outputs(1215)) and not (layer3_outputs(2248));
    layer4_outputs(1504) <= not(layer3_outputs(1919));
    layer4_outputs(1505) <= layer3_outputs(2333);
    layer4_outputs(1506) <= not(layer3_outputs(1141)) or (layer3_outputs(1461));
    layer4_outputs(1507) <= '1';
    layer4_outputs(1508) <= not((layer3_outputs(2378)) xor (layer3_outputs(348)));
    layer4_outputs(1509) <= not(layer3_outputs(1874));
    layer4_outputs(1510) <= not(layer3_outputs(180));
    layer4_outputs(1511) <= not((layer3_outputs(363)) or (layer3_outputs(2147)));
    layer4_outputs(1512) <= not((layer3_outputs(2284)) or (layer3_outputs(1716)));
    layer4_outputs(1513) <= not(layer3_outputs(911));
    layer4_outputs(1514) <= not(layer3_outputs(417));
    layer4_outputs(1515) <= (layer3_outputs(1232)) or (layer3_outputs(720));
    layer4_outputs(1516) <= layer3_outputs(1272);
    layer4_outputs(1517) <= (layer3_outputs(1061)) and (layer3_outputs(1268));
    layer4_outputs(1518) <= not(layer3_outputs(2261)) or (layer3_outputs(2375));
    layer4_outputs(1519) <= (layer3_outputs(810)) xor (layer3_outputs(1604));
    layer4_outputs(1520) <= not((layer3_outputs(1593)) and (layer3_outputs(2160)));
    layer4_outputs(1521) <= layer3_outputs(1805);
    layer4_outputs(1522) <= '1';
    layer4_outputs(1523) <= layer3_outputs(1519);
    layer4_outputs(1524) <= not(layer3_outputs(249)) or (layer3_outputs(2083));
    layer4_outputs(1525) <= layer3_outputs(2182);
    layer4_outputs(1526) <= '1';
    layer4_outputs(1527) <= not((layer3_outputs(1795)) xor (layer3_outputs(2205)));
    layer4_outputs(1528) <= (layer3_outputs(2436)) xor (layer3_outputs(604));
    layer4_outputs(1529) <= not((layer3_outputs(338)) and (layer3_outputs(1343)));
    layer4_outputs(1530) <= not((layer3_outputs(934)) or (layer3_outputs(2186)));
    layer4_outputs(1531) <= not((layer3_outputs(2193)) or (layer3_outputs(2233)));
    layer4_outputs(1532) <= (layer3_outputs(2244)) and (layer3_outputs(1048));
    layer4_outputs(1533) <= not(layer3_outputs(2064));
    layer4_outputs(1534) <= layer3_outputs(687);
    layer4_outputs(1535) <= layer3_outputs(1140);
    layer4_outputs(1536) <= (layer3_outputs(1397)) and not (layer3_outputs(1119));
    layer4_outputs(1537) <= (layer3_outputs(2094)) and not (layer3_outputs(2451));
    layer4_outputs(1538) <= (layer3_outputs(109)) and (layer3_outputs(676));
    layer4_outputs(1539) <= layer3_outputs(237);
    layer4_outputs(1540) <= layer3_outputs(1426);
    layer4_outputs(1541) <= (layer3_outputs(217)) and not (layer3_outputs(1854));
    layer4_outputs(1542) <= '1';
    layer4_outputs(1543) <= not(layer3_outputs(1447));
    layer4_outputs(1544) <= not(layer3_outputs(1591)) or (layer3_outputs(1806));
    layer4_outputs(1545) <= (layer3_outputs(684)) and not (layer3_outputs(936));
    layer4_outputs(1546) <= not(layer3_outputs(1214)) or (layer3_outputs(932));
    layer4_outputs(1547) <= '1';
    layer4_outputs(1548) <= not((layer3_outputs(408)) or (layer3_outputs(2392)));
    layer4_outputs(1549) <= not(layer3_outputs(803)) or (layer3_outputs(990));
    layer4_outputs(1550) <= (layer3_outputs(130)) and not (layer3_outputs(1130));
    layer4_outputs(1551) <= not((layer3_outputs(308)) and (layer3_outputs(587)));
    layer4_outputs(1552) <= not(layer3_outputs(1399)) or (layer3_outputs(225));
    layer4_outputs(1553) <= not(layer3_outputs(1606)) or (layer3_outputs(1178));
    layer4_outputs(1554) <= (layer3_outputs(1518)) and (layer3_outputs(460));
    layer4_outputs(1555) <= layer3_outputs(1059);
    layer4_outputs(1556) <= layer3_outputs(2276);
    layer4_outputs(1557) <= not(layer3_outputs(1228));
    layer4_outputs(1558) <= layer3_outputs(2250);
    layer4_outputs(1559) <= (layer3_outputs(298)) and not (layer3_outputs(1699));
    layer4_outputs(1560) <= layer3_outputs(2234);
    layer4_outputs(1561) <= '0';
    layer4_outputs(1562) <= not(layer3_outputs(2185));
    layer4_outputs(1563) <= not(layer3_outputs(2065)) or (layer3_outputs(1570));
    layer4_outputs(1564) <= not(layer3_outputs(1134)) or (layer3_outputs(1301));
    layer4_outputs(1565) <= not(layer3_outputs(599));
    layer4_outputs(1566) <= not((layer3_outputs(416)) xor (layer3_outputs(1640)));
    layer4_outputs(1567) <= not(layer3_outputs(1718));
    layer4_outputs(1568) <= (layer3_outputs(2274)) and not (layer3_outputs(550));
    layer4_outputs(1569) <= (layer3_outputs(562)) and not (layer3_outputs(1234));
    layer4_outputs(1570) <= not(layer3_outputs(1969));
    layer4_outputs(1571) <= '1';
    layer4_outputs(1572) <= not(layer3_outputs(2045));
    layer4_outputs(1573) <= not((layer3_outputs(2309)) or (layer3_outputs(2316)));
    layer4_outputs(1574) <= not(layer3_outputs(9));
    layer4_outputs(1575) <= not(layer3_outputs(76)) or (layer3_outputs(1965));
    layer4_outputs(1576) <= (layer3_outputs(405)) and (layer3_outputs(2433));
    layer4_outputs(1577) <= not(layer3_outputs(2001)) or (layer3_outputs(283));
    layer4_outputs(1578) <= '0';
    layer4_outputs(1579) <= not((layer3_outputs(777)) and (layer3_outputs(2191)));
    layer4_outputs(1580) <= (layer3_outputs(793)) and (layer3_outputs(2468));
    layer4_outputs(1581) <= not((layer3_outputs(2550)) xor (layer3_outputs(1189)));
    layer4_outputs(1582) <= (layer3_outputs(135)) and not (layer3_outputs(1003));
    layer4_outputs(1583) <= (layer3_outputs(424)) and (layer3_outputs(1106));
    layer4_outputs(1584) <= layer3_outputs(2497);
    layer4_outputs(1585) <= not((layer3_outputs(1207)) and (layer3_outputs(513)));
    layer4_outputs(1586) <= not((layer3_outputs(89)) or (layer3_outputs(1009)));
    layer4_outputs(1587) <= layer3_outputs(1811);
    layer4_outputs(1588) <= not(layer3_outputs(1282));
    layer4_outputs(1589) <= not(layer3_outputs(502));
    layer4_outputs(1590) <= (layer3_outputs(899)) and not (layer3_outputs(2307));
    layer4_outputs(1591) <= (layer3_outputs(2302)) and not (layer3_outputs(1910));
    layer4_outputs(1592) <= '0';
    layer4_outputs(1593) <= layer3_outputs(1956);
    layer4_outputs(1594) <= '1';
    layer4_outputs(1595) <= (layer3_outputs(1074)) or (layer3_outputs(2171));
    layer4_outputs(1596) <= layer3_outputs(1873);
    layer4_outputs(1597) <= not(layer3_outputs(1290));
    layer4_outputs(1598) <= layer3_outputs(213);
    layer4_outputs(1599) <= (layer3_outputs(2038)) and not (layer3_outputs(1718));
    layer4_outputs(1600) <= (layer3_outputs(139)) and not (layer3_outputs(2423));
    layer4_outputs(1601) <= layer3_outputs(2486);
    layer4_outputs(1602) <= layer3_outputs(824);
    layer4_outputs(1603) <= (layer3_outputs(295)) and not (layer3_outputs(92));
    layer4_outputs(1604) <= layer3_outputs(1086);
    layer4_outputs(1605) <= layer3_outputs(864);
    layer4_outputs(1606) <= layer3_outputs(1828);
    layer4_outputs(1607) <= not((layer3_outputs(2400)) xor (layer3_outputs(1587)));
    layer4_outputs(1608) <= '0';
    layer4_outputs(1609) <= layer3_outputs(284);
    layer4_outputs(1610) <= layer3_outputs(732);
    layer4_outputs(1611) <= not(layer3_outputs(774));
    layer4_outputs(1612) <= not(layer3_outputs(2252));
    layer4_outputs(1613) <= '1';
    layer4_outputs(1614) <= not(layer3_outputs(1021));
    layer4_outputs(1615) <= (layer3_outputs(1388)) and (layer3_outputs(159));
    layer4_outputs(1616) <= not(layer3_outputs(2512));
    layer4_outputs(1617) <= layer3_outputs(992);
    layer4_outputs(1618) <= (layer3_outputs(1567)) and (layer3_outputs(2292));
    layer4_outputs(1619) <= layer3_outputs(1111);
    layer4_outputs(1620) <= (layer3_outputs(574)) or (layer3_outputs(1572));
    layer4_outputs(1621) <= layer3_outputs(1131);
    layer4_outputs(1622) <= layer3_outputs(1847);
    layer4_outputs(1623) <= not(layer3_outputs(1759));
    layer4_outputs(1624) <= layer3_outputs(1514);
    layer4_outputs(1625) <= not(layer3_outputs(1030)) or (layer3_outputs(1935));
    layer4_outputs(1626) <= layer3_outputs(1235);
    layer4_outputs(1627) <= not(layer3_outputs(2331));
    layer4_outputs(1628) <= '1';
    layer4_outputs(1629) <= '1';
    layer4_outputs(1630) <= layer3_outputs(1548);
    layer4_outputs(1631) <= not(layer3_outputs(1432));
    layer4_outputs(1632) <= '1';
    layer4_outputs(1633) <= (layer3_outputs(1782)) and not (layer3_outputs(755));
    layer4_outputs(1634) <= layer3_outputs(79);
    layer4_outputs(1635) <= layer3_outputs(492);
    layer4_outputs(1636) <= not(layer3_outputs(552)) or (layer3_outputs(1073));
    layer4_outputs(1637) <= (layer3_outputs(1778)) and not (layer3_outputs(1880));
    layer4_outputs(1638) <= not((layer3_outputs(194)) or (layer3_outputs(1409)));
    layer4_outputs(1639) <= not(layer3_outputs(2165));
    layer4_outputs(1640) <= not(layer3_outputs(2538));
    layer4_outputs(1641) <= not(layer3_outputs(1045)) or (layer3_outputs(1818));
    layer4_outputs(1642) <= not(layer3_outputs(309));
    layer4_outputs(1643) <= not((layer3_outputs(1781)) and (layer3_outputs(2216)));
    layer4_outputs(1644) <= layer3_outputs(2547);
    layer4_outputs(1645) <= layer3_outputs(98);
    layer4_outputs(1646) <= not(layer3_outputs(474));
    layer4_outputs(1647) <= (layer3_outputs(2090)) and (layer3_outputs(54));
    layer4_outputs(1648) <= layer3_outputs(2456);
    layer4_outputs(1649) <= not(layer3_outputs(1961));
    layer4_outputs(1650) <= (layer3_outputs(1965)) xor (layer3_outputs(1363));
    layer4_outputs(1651) <= (layer3_outputs(1581)) and not (layer3_outputs(345));
    layer4_outputs(1652) <= not(layer3_outputs(735));
    layer4_outputs(1653) <= (layer3_outputs(1937)) or (layer3_outputs(2551));
    layer4_outputs(1654) <= '1';
    layer4_outputs(1655) <= layer3_outputs(748);
    layer4_outputs(1656) <= '0';
    layer4_outputs(1657) <= not(layer3_outputs(1674));
    layer4_outputs(1658) <= '0';
    layer4_outputs(1659) <= layer3_outputs(2347);
    layer4_outputs(1660) <= not(layer3_outputs(546));
    layer4_outputs(1661) <= layer3_outputs(1236);
    layer4_outputs(1662) <= not(layer3_outputs(1176));
    layer4_outputs(1663) <= not(layer3_outputs(1864)) or (layer3_outputs(228));
    layer4_outputs(1664) <= not(layer3_outputs(1179)) or (layer3_outputs(630));
    layer4_outputs(1665) <= layer3_outputs(2007);
    layer4_outputs(1666) <= (layer3_outputs(1405)) and (layer3_outputs(1533));
    layer4_outputs(1667) <= layer3_outputs(178);
    layer4_outputs(1668) <= layer3_outputs(109);
    layer4_outputs(1669) <= layer3_outputs(134);
    layer4_outputs(1670) <= (layer3_outputs(237)) and not (layer3_outputs(1199));
    layer4_outputs(1671) <= not(layer3_outputs(815)) or (layer3_outputs(1687));
    layer4_outputs(1672) <= not((layer3_outputs(53)) xor (layer3_outputs(211)));
    layer4_outputs(1673) <= layer3_outputs(1376);
    layer4_outputs(1674) <= not(layer3_outputs(705));
    layer4_outputs(1675) <= (layer3_outputs(2126)) or (layer3_outputs(1334));
    layer4_outputs(1676) <= layer3_outputs(576);
    layer4_outputs(1677) <= (layer3_outputs(2462)) and not (layer3_outputs(1425));
    layer4_outputs(1678) <= '1';
    layer4_outputs(1679) <= not(layer3_outputs(1033));
    layer4_outputs(1680) <= (layer3_outputs(1442)) and not (layer3_outputs(2016));
    layer4_outputs(1681) <= (layer3_outputs(56)) and not (layer3_outputs(2112));
    layer4_outputs(1682) <= (layer3_outputs(895)) and not (layer3_outputs(386));
    layer4_outputs(1683) <= not(layer3_outputs(2403)) or (layer3_outputs(1502));
    layer4_outputs(1684) <= layer3_outputs(277);
    layer4_outputs(1685) <= (layer3_outputs(619)) and (layer3_outputs(157));
    layer4_outputs(1686) <= not(layer3_outputs(155));
    layer4_outputs(1687) <= not(layer3_outputs(2056));
    layer4_outputs(1688) <= not(layer3_outputs(709)) or (layer3_outputs(1985));
    layer4_outputs(1689) <= (layer3_outputs(1047)) and not (layer3_outputs(751));
    layer4_outputs(1690) <= (layer3_outputs(145)) and not (layer3_outputs(1364));
    layer4_outputs(1691) <= not(layer3_outputs(1053)) or (layer3_outputs(2277));
    layer4_outputs(1692) <= not(layer3_outputs(2159)) or (layer3_outputs(1329));
    layer4_outputs(1693) <= not((layer3_outputs(547)) xor (layer3_outputs(288)));
    layer4_outputs(1694) <= not(layer3_outputs(1440)) or (layer3_outputs(722));
    layer4_outputs(1695) <= not(layer3_outputs(1143));
    layer4_outputs(1696) <= not(layer3_outputs(406)) or (layer3_outputs(1659));
    layer4_outputs(1697) <= not(layer3_outputs(132));
    layer4_outputs(1698) <= layer3_outputs(901);
    layer4_outputs(1699) <= not(layer3_outputs(2523));
    layer4_outputs(1700) <= layer3_outputs(2255);
    layer4_outputs(1701) <= not((layer3_outputs(1151)) and (layer3_outputs(2091)));
    layer4_outputs(1702) <= not(layer3_outputs(1398));
    layer4_outputs(1703) <= layer3_outputs(2028);
    layer4_outputs(1704) <= not(layer3_outputs(2189));
    layer4_outputs(1705) <= not(layer3_outputs(2003));
    layer4_outputs(1706) <= not(layer3_outputs(1852));
    layer4_outputs(1707) <= not((layer3_outputs(1401)) or (layer3_outputs(1741)));
    layer4_outputs(1708) <= layer3_outputs(947);
    layer4_outputs(1709) <= (layer3_outputs(269)) and (layer3_outputs(2502));
    layer4_outputs(1710) <= not(layer3_outputs(337)) or (layer3_outputs(1049));
    layer4_outputs(1711) <= (layer3_outputs(1770)) and not (layer3_outputs(2135));
    layer4_outputs(1712) <= not((layer3_outputs(1693)) xor (layer3_outputs(806)));
    layer4_outputs(1713) <= (layer3_outputs(2097)) and (layer3_outputs(559));
    layer4_outputs(1714) <= not(layer3_outputs(970)) or (layer3_outputs(2184));
    layer4_outputs(1715) <= (layer3_outputs(2377)) and (layer3_outputs(1448));
    layer4_outputs(1716) <= '1';
    layer4_outputs(1717) <= (layer3_outputs(745)) xor (layer3_outputs(409));
    layer4_outputs(1718) <= layer3_outputs(717);
    layer4_outputs(1719) <= not((layer3_outputs(454)) and (layer3_outputs(2343)));
    layer4_outputs(1720) <= layer3_outputs(1082);
    layer4_outputs(1721) <= not((layer3_outputs(1880)) or (layer3_outputs(986)));
    layer4_outputs(1722) <= '0';
    layer4_outputs(1723) <= not(layer3_outputs(223));
    layer4_outputs(1724) <= layer3_outputs(1261);
    layer4_outputs(1725) <= (layer3_outputs(553)) and (layer3_outputs(68));
    layer4_outputs(1726) <= not((layer3_outputs(1396)) and (layer3_outputs(1250)));
    layer4_outputs(1727) <= layer3_outputs(679);
    layer4_outputs(1728) <= (layer3_outputs(881)) and not (layer3_outputs(1008));
    layer4_outputs(1729) <= (layer3_outputs(725)) or (layer3_outputs(2389));
    layer4_outputs(1730) <= not(layer3_outputs(332));
    layer4_outputs(1731) <= layer3_outputs(1971);
    layer4_outputs(1732) <= layer3_outputs(2084);
    layer4_outputs(1733) <= (layer3_outputs(898)) and not (layer3_outputs(112));
    layer4_outputs(1734) <= layer3_outputs(370);
    layer4_outputs(1735) <= (layer3_outputs(584)) and not (layer3_outputs(2455));
    layer4_outputs(1736) <= layer3_outputs(1809);
    layer4_outputs(1737) <= not(layer3_outputs(2365));
    layer4_outputs(1738) <= not((layer3_outputs(2203)) and (layer3_outputs(1822)));
    layer4_outputs(1739) <= not(layer3_outputs(534)) or (layer3_outputs(1216));
    layer4_outputs(1740) <= not(layer3_outputs(2452));
    layer4_outputs(1741) <= (layer3_outputs(1536)) or (layer3_outputs(1137));
    layer4_outputs(1742) <= not(layer3_outputs(540));
    layer4_outputs(1743) <= '1';
    layer4_outputs(1744) <= not(layer3_outputs(1785));
    layer4_outputs(1745) <= not(layer3_outputs(1610)) or (layer3_outputs(1078));
    layer4_outputs(1746) <= not(layer3_outputs(2457));
    layer4_outputs(1747) <= (layer3_outputs(1208)) and not (layer3_outputs(749));
    layer4_outputs(1748) <= '1';
    layer4_outputs(1749) <= not(layer3_outputs(1244)) or (layer3_outputs(1225));
    layer4_outputs(1750) <= not(layer3_outputs(2519));
    layer4_outputs(1751) <= not(layer3_outputs(682)) or (layer3_outputs(725));
    layer4_outputs(1752) <= layer3_outputs(2313);
    layer4_outputs(1753) <= (layer3_outputs(933)) xor (layer3_outputs(2495));
    layer4_outputs(1754) <= '1';
    layer4_outputs(1755) <= (layer3_outputs(1762)) and not (layer3_outputs(2104));
    layer4_outputs(1756) <= not(layer3_outputs(340));
    layer4_outputs(1757) <= (layer3_outputs(1165)) and not (layer3_outputs(724));
    layer4_outputs(1758) <= layer3_outputs(2483);
    layer4_outputs(1759) <= layer3_outputs(1532);
    layer4_outputs(1760) <= layer3_outputs(2350);
    layer4_outputs(1761) <= not(layer3_outputs(643));
    layer4_outputs(1762) <= not((layer3_outputs(270)) or (layer3_outputs(2038)));
    layer4_outputs(1763) <= not((layer3_outputs(504)) and (layer3_outputs(446)));
    layer4_outputs(1764) <= not(layer3_outputs(1567));
    layer4_outputs(1765) <= not((layer3_outputs(2172)) and (layer3_outputs(680)));
    layer4_outputs(1766) <= layer3_outputs(2456);
    layer4_outputs(1767) <= not((layer3_outputs(1488)) and (layer3_outputs(2212)));
    layer4_outputs(1768) <= not((layer3_outputs(2353)) xor (layer3_outputs(661)));
    layer4_outputs(1769) <= (layer3_outputs(565)) or (layer3_outputs(1799));
    layer4_outputs(1770) <= not((layer3_outputs(829)) and (layer3_outputs(290)));
    layer4_outputs(1771) <= '1';
    layer4_outputs(1772) <= not(layer3_outputs(1493)) or (layer3_outputs(2517));
    layer4_outputs(1773) <= layer3_outputs(972);
    layer4_outputs(1774) <= '1';
    layer4_outputs(1775) <= '1';
    layer4_outputs(1776) <= not((layer3_outputs(1025)) xor (layer3_outputs(1325)));
    layer4_outputs(1777) <= not(layer3_outputs(2428));
    layer4_outputs(1778) <= not(layer3_outputs(1728));
    layer4_outputs(1779) <= layer3_outputs(528);
    layer4_outputs(1780) <= not(layer3_outputs(2350));
    layer4_outputs(1781) <= (layer3_outputs(501)) and not (layer3_outputs(2441));
    layer4_outputs(1782) <= layer3_outputs(2434);
    layer4_outputs(1783) <= not(layer3_outputs(36));
    layer4_outputs(1784) <= (layer3_outputs(289)) and not (layer3_outputs(90));
    layer4_outputs(1785) <= not(layer3_outputs(1646)) or (layer3_outputs(480));
    layer4_outputs(1786) <= not(layer3_outputs(1542));
    layer4_outputs(1787) <= layer3_outputs(335);
    layer4_outputs(1788) <= '0';
    layer4_outputs(1789) <= '1';
    layer4_outputs(1790) <= not((layer3_outputs(255)) or (layer3_outputs(742)));
    layer4_outputs(1791) <= layer3_outputs(703);
    layer4_outputs(1792) <= layer3_outputs(138);
    layer4_outputs(1793) <= layer3_outputs(1929);
    layer4_outputs(1794) <= layer3_outputs(1185);
    layer4_outputs(1795) <= (layer3_outputs(2373)) and not (layer3_outputs(1664));
    layer4_outputs(1796) <= (layer3_outputs(1251)) or (layer3_outputs(1744));
    layer4_outputs(1797) <= (layer3_outputs(1588)) and not (layer3_outputs(768));
    layer4_outputs(1798) <= '1';
    layer4_outputs(1799) <= layer3_outputs(108);
    layer4_outputs(1800) <= not(layer3_outputs(296));
    layer4_outputs(1801) <= layer3_outputs(1066);
    layer4_outputs(1802) <= not(layer3_outputs(672));
    layer4_outputs(1803) <= (layer3_outputs(1731)) and not (layer3_outputs(1801));
    layer4_outputs(1804) <= (layer3_outputs(488)) and not (layer3_outputs(1545));
    layer4_outputs(1805) <= not(layer3_outputs(1894));
    layer4_outputs(1806) <= not(layer3_outputs(1501));
    layer4_outputs(1807) <= not(layer3_outputs(1644)) or (layer3_outputs(2115));
    layer4_outputs(1808) <= not(layer3_outputs(1013));
    layer4_outputs(1809) <= not(layer3_outputs(2073));
    layer4_outputs(1810) <= not(layer3_outputs(716));
    layer4_outputs(1811) <= not(layer3_outputs(2530));
    layer4_outputs(1812) <= not((layer3_outputs(379)) xor (layer3_outputs(1168)));
    layer4_outputs(1813) <= (layer3_outputs(0)) and not (layer3_outputs(2251));
    layer4_outputs(1814) <= not(layer3_outputs(1500)) or (layer3_outputs(1873));
    layer4_outputs(1815) <= not(layer3_outputs(975));
    layer4_outputs(1816) <= not((layer3_outputs(845)) and (layer3_outputs(1410)));
    layer4_outputs(1817) <= layer3_outputs(350);
    layer4_outputs(1818) <= not(layer3_outputs(1077)) or (layer3_outputs(464));
    layer4_outputs(1819) <= layer3_outputs(299);
    layer4_outputs(1820) <= '1';
    layer4_outputs(1821) <= (layer3_outputs(1371)) or (layer3_outputs(988));
    layer4_outputs(1822) <= not(layer3_outputs(67));
    layer4_outputs(1823) <= not(layer3_outputs(2427));
    layer4_outputs(1824) <= not((layer3_outputs(519)) and (layer3_outputs(521)));
    layer4_outputs(1825) <= not(layer3_outputs(1681)) or (layer3_outputs(247));
    layer4_outputs(1826) <= (layer3_outputs(1132)) or (layer3_outputs(1530));
    layer4_outputs(1827) <= layer3_outputs(1532);
    layer4_outputs(1828) <= '1';
    layer4_outputs(1829) <= not((layer3_outputs(249)) xor (layer3_outputs(2147)));
    layer4_outputs(1830) <= not((layer3_outputs(557)) and (layer3_outputs(421)));
    layer4_outputs(1831) <= layer3_outputs(2274);
    layer4_outputs(1832) <= layer3_outputs(593);
    layer4_outputs(1833) <= not(layer3_outputs(906));
    layer4_outputs(1834) <= not(layer3_outputs(1561)) or (layer3_outputs(707));
    layer4_outputs(1835) <= layer3_outputs(1595);
    layer4_outputs(1836) <= not(layer3_outputs(668)) or (layer3_outputs(842));
    layer4_outputs(1837) <= '0';
    layer4_outputs(1838) <= layer3_outputs(1865);
    layer4_outputs(1839) <= (layer3_outputs(1160)) and (layer3_outputs(1326));
    layer4_outputs(1840) <= layer3_outputs(854);
    layer4_outputs(1841) <= (layer3_outputs(1860)) xor (layer3_outputs(284));
    layer4_outputs(1842) <= layer3_outputs(906);
    layer4_outputs(1843) <= not(layer3_outputs(1389));
    layer4_outputs(1844) <= not((layer3_outputs(2280)) or (layer3_outputs(1158)));
    layer4_outputs(1845) <= not((layer3_outputs(358)) and (layer3_outputs(1026)));
    layer4_outputs(1846) <= (layer3_outputs(2543)) and (layer3_outputs(1359));
    layer4_outputs(1847) <= not(layer3_outputs(2338));
    layer4_outputs(1848) <= not(layer3_outputs(1094)) or (layer3_outputs(937));
    layer4_outputs(1849) <= layer3_outputs(298);
    layer4_outputs(1850) <= (layer3_outputs(2426)) and not (layer3_outputs(335));
    layer4_outputs(1851) <= (layer3_outputs(1412)) xor (layer3_outputs(551));
    layer4_outputs(1852) <= layer3_outputs(621);
    layer4_outputs(1853) <= (layer3_outputs(1126)) and not (layer3_outputs(126));
    layer4_outputs(1854) <= not((layer3_outputs(1958)) xor (layer3_outputs(1966)));
    layer4_outputs(1855) <= not(layer3_outputs(1291));
    layer4_outputs(1856) <= not(layer3_outputs(1734));
    layer4_outputs(1857) <= not(layer3_outputs(2414)) or (layer3_outputs(231));
    layer4_outputs(1858) <= (layer3_outputs(2170)) or (layer3_outputs(988));
    layer4_outputs(1859) <= not((layer3_outputs(1191)) or (layer3_outputs(2032)));
    layer4_outputs(1860) <= not(layer3_outputs(278));
    layer4_outputs(1861) <= (layer3_outputs(373)) or (layer3_outputs(1169));
    layer4_outputs(1862) <= '1';
    layer4_outputs(1863) <= not(layer3_outputs(590)) or (layer3_outputs(419));
    layer4_outputs(1864) <= not(layer3_outputs(2474));
    layer4_outputs(1865) <= layer3_outputs(1209);
    layer4_outputs(1866) <= (layer3_outputs(1184)) xor (layer3_outputs(1443));
    layer4_outputs(1867) <= not(layer3_outputs(2352));
    layer4_outputs(1868) <= not(layer3_outputs(1615));
    layer4_outputs(1869) <= (layer3_outputs(1673)) and not (layer3_outputs(2253));
    layer4_outputs(1870) <= (layer3_outputs(2086)) and not (layer3_outputs(1192));
    layer4_outputs(1871) <= not(layer3_outputs(1420));
    layer4_outputs(1872) <= not((layer3_outputs(1832)) or (layer3_outputs(1076)));
    layer4_outputs(1873) <= layer3_outputs(224);
    layer4_outputs(1874) <= not(layer3_outputs(1297)) or (layer3_outputs(2101));
    layer4_outputs(1875) <= layer3_outputs(2124);
    layer4_outputs(1876) <= layer3_outputs(2356);
    layer4_outputs(1877) <= (layer3_outputs(2286)) or (layer3_outputs(2338));
    layer4_outputs(1878) <= not(layer3_outputs(1541));
    layer4_outputs(1879) <= not(layer3_outputs(2360)) or (layer3_outputs(908));
    layer4_outputs(1880) <= layer3_outputs(233);
    layer4_outputs(1881) <= not(layer3_outputs(2022));
    layer4_outputs(1882) <= layer3_outputs(1467);
    layer4_outputs(1883) <= layer3_outputs(382);
    layer4_outputs(1884) <= not(layer3_outputs(775));
    layer4_outputs(1885) <= not(layer3_outputs(401));
    layer4_outputs(1886) <= (layer3_outputs(176)) xor (layer3_outputs(2422));
    layer4_outputs(1887) <= not(layer3_outputs(982));
    layer4_outputs(1888) <= not(layer3_outputs(688));
    layer4_outputs(1889) <= not(layer3_outputs(1102)) or (layer3_outputs(2389));
    layer4_outputs(1890) <= not((layer3_outputs(2184)) or (layer3_outputs(603)));
    layer4_outputs(1891) <= not((layer3_outputs(699)) or (layer3_outputs(28)));
    layer4_outputs(1892) <= not(layer3_outputs(849)) or (layer3_outputs(995));
    layer4_outputs(1893) <= (layer3_outputs(1353)) and not (layer3_outputs(1742));
    layer4_outputs(1894) <= (layer3_outputs(2527)) and (layer3_outputs(2106));
    layer4_outputs(1895) <= not(layer3_outputs(2167)) or (layer3_outputs(4));
    layer4_outputs(1896) <= not((layer3_outputs(349)) and (layer3_outputs(44)));
    layer4_outputs(1897) <= not(layer3_outputs(837));
    layer4_outputs(1898) <= (layer3_outputs(200)) and not (layer3_outputs(2141));
    layer4_outputs(1899) <= (layer3_outputs(2005)) xor (layer3_outputs(1814));
    layer4_outputs(1900) <= not(layer3_outputs(10));
    layer4_outputs(1901) <= (layer3_outputs(1226)) or (layer3_outputs(1710));
    layer4_outputs(1902) <= not(layer3_outputs(128));
    layer4_outputs(1903) <= not(layer3_outputs(623));
    layer4_outputs(1904) <= not((layer3_outputs(132)) xor (layer3_outputs(196)));
    layer4_outputs(1905) <= (layer3_outputs(356)) and not (layer3_outputs(2089));
    layer4_outputs(1906) <= not(layer3_outputs(1962));
    layer4_outputs(1907) <= not(layer3_outputs(1476));
    layer4_outputs(1908) <= not(layer3_outputs(2425));
    layer4_outputs(1909) <= layer3_outputs(96);
    layer4_outputs(1910) <= layer3_outputs(1135);
    layer4_outputs(1911) <= layer3_outputs(813);
    layer4_outputs(1912) <= layer3_outputs(1667);
    layer4_outputs(1913) <= layer3_outputs(2559);
    layer4_outputs(1914) <= not((layer3_outputs(307)) or (layer3_outputs(2541)));
    layer4_outputs(1915) <= not((layer3_outputs(2341)) xor (layer3_outputs(1781)));
    layer4_outputs(1916) <= layer3_outputs(1038);
    layer4_outputs(1917) <= layer3_outputs(372);
    layer4_outputs(1918) <= not(layer3_outputs(2117)) or (layer3_outputs(1843));
    layer4_outputs(1919) <= (layer3_outputs(400)) and (layer3_outputs(248));
    layer4_outputs(1920) <= (layer3_outputs(149)) and (layer3_outputs(892));
    layer4_outputs(1921) <= layer3_outputs(72);
    layer4_outputs(1922) <= not(layer3_outputs(1717));
    layer4_outputs(1923) <= not((layer3_outputs(992)) and (layer3_outputs(1425)));
    layer4_outputs(1924) <= '1';
    layer4_outputs(1925) <= layer3_outputs(1293);
    layer4_outputs(1926) <= layer3_outputs(1706);
    layer4_outputs(1927) <= (layer3_outputs(2380)) and not (layer3_outputs(2266));
    layer4_outputs(1928) <= not(layer3_outputs(794));
    layer4_outputs(1929) <= '0';
    layer4_outputs(1930) <= not(layer3_outputs(149));
    layer4_outputs(1931) <= (layer3_outputs(635)) or (layer3_outputs(646));
    layer4_outputs(1932) <= layer3_outputs(717);
    layer4_outputs(1933) <= layer3_outputs(1045);
    layer4_outputs(1934) <= (layer3_outputs(2098)) and (layer3_outputs(850));
    layer4_outputs(1935) <= not((layer3_outputs(696)) or (layer3_outputs(1953)));
    layer4_outputs(1936) <= (layer3_outputs(1261)) and (layer3_outputs(231));
    layer4_outputs(1937) <= layer3_outputs(1457);
    layer4_outputs(1938) <= not(layer3_outputs(2229));
    layer4_outputs(1939) <= not(layer3_outputs(1952));
    layer4_outputs(1940) <= '0';
    layer4_outputs(1941) <= not((layer3_outputs(1355)) and (layer3_outputs(672)));
    layer4_outputs(1942) <= not(layer3_outputs(1276)) or (layer3_outputs(2517));
    layer4_outputs(1943) <= not((layer3_outputs(1529)) or (layer3_outputs(1160)));
    layer4_outputs(1944) <= not(layer3_outputs(1655));
    layer4_outputs(1945) <= '1';
    layer4_outputs(1946) <= (layer3_outputs(378)) and not (layer3_outputs(1817));
    layer4_outputs(1947) <= layer3_outputs(1380);
    layer4_outputs(1948) <= (layer3_outputs(1456)) and not (layer3_outputs(230));
    layer4_outputs(1949) <= not((layer3_outputs(966)) and (layer3_outputs(525)));
    layer4_outputs(1950) <= not(layer3_outputs(716));
    layer4_outputs(1951) <= (layer3_outputs(1360)) or (layer3_outputs(239));
    layer4_outputs(1952) <= (layer3_outputs(2)) and (layer3_outputs(1245));
    layer4_outputs(1953) <= (layer3_outputs(2325)) and not (layer3_outputs(915));
    layer4_outputs(1954) <= '1';
    layer4_outputs(1955) <= layer3_outputs(1093);
    layer4_outputs(1956) <= layer3_outputs(1907);
    layer4_outputs(1957) <= (layer3_outputs(1481)) xor (layer3_outputs(2328));
    layer4_outputs(1958) <= (layer3_outputs(2329)) or (layer3_outputs(2348));
    layer4_outputs(1959) <= not((layer3_outputs(1465)) and (layer3_outputs(548)));
    layer4_outputs(1960) <= '1';
    layer4_outputs(1961) <= (layer3_outputs(2128)) and (layer3_outputs(398));
    layer4_outputs(1962) <= not(layer3_outputs(2374));
    layer4_outputs(1963) <= layer3_outputs(2079);
    layer4_outputs(1964) <= not(layer3_outputs(2503));
    layer4_outputs(1965) <= not(layer3_outputs(1792)) or (layer3_outputs(877));
    layer4_outputs(1966) <= not((layer3_outputs(1248)) and (layer3_outputs(1888)));
    layer4_outputs(1967) <= (layer3_outputs(1826)) and not (layer3_outputs(668));
    layer4_outputs(1968) <= layer3_outputs(2454);
    layer4_outputs(1969) <= not(layer3_outputs(575));
    layer4_outputs(1970) <= not((layer3_outputs(21)) xor (layer3_outputs(265)));
    layer4_outputs(1971) <= layer3_outputs(402);
    layer4_outputs(1972) <= '0';
    layer4_outputs(1973) <= '0';
    layer4_outputs(1974) <= not((layer3_outputs(1939)) and (layer3_outputs(1206)));
    layer4_outputs(1975) <= '1';
    layer4_outputs(1976) <= '0';
    layer4_outputs(1977) <= layer3_outputs(1069);
    layer4_outputs(1978) <= not((layer3_outputs(93)) or (layer3_outputs(1751)));
    layer4_outputs(1979) <= not(layer3_outputs(2547)) or (layer3_outputs(3));
    layer4_outputs(1980) <= layer3_outputs(27);
    layer4_outputs(1981) <= not(layer3_outputs(675)) or (layer3_outputs(1766));
    layer4_outputs(1982) <= not(layer3_outputs(1778));
    layer4_outputs(1983) <= '0';
    layer4_outputs(1984) <= layer3_outputs(1269);
    layer4_outputs(1985) <= (layer3_outputs(2459)) and not (layer3_outputs(113));
    layer4_outputs(1986) <= '1';
    layer4_outputs(1987) <= not(layer3_outputs(154)) or (layer3_outputs(111));
    layer4_outputs(1988) <= not(layer3_outputs(143)) or (layer3_outputs(224));
    layer4_outputs(1989) <= (layer3_outputs(2029)) and (layer3_outputs(1108));
    layer4_outputs(1990) <= '1';
    layer4_outputs(1991) <= not(layer3_outputs(1125)) or (layer3_outputs(329));
    layer4_outputs(1992) <= '1';
    layer4_outputs(1993) <= (layer3_outputs(1250)) and not (layer3_outputs(628));
    layer4_outputs(1994) <= (layer3_outputs(1347)) and not (layer3_outputs(1269));
    layer4_outputs(1995) <= not(layer3_outputs(1730));
    layer4_outputs(1996) <= layer3_outputs(1706);
    layer4_outputs(1997) <= '0';
    layer4_outputs(1998) <= (layer3_outputs(961)) or (layer3_outputs(1222));
    layer4_outputs(1999) <= not(layer3_outputs(647));
    layer4_outputs(2000) <= (layer3_outputs(1631)) xor (layer3_outputs(1016));
    layer4_outputs(2001) <= layer3_outputs(1395);
    layer4_outputs(2002) <= (layer3_outputs(37)) or (layer3_outputs(201));
    layer4_outputs(2003) <= not(layer3_outputs(2411));
    layer4_outputs(2004) <= not(layer3_outputs(1029)) or (layer3_outputs(1144));
    layer4_outputs(2005) <= layer3_outputs(2432);
    layer4_outputs(2006) <= '0';
    layer4_outputs(2007) <= '0';
    layer4_outputs(2008) <= (layer3_outputs(1329)) and not (layer3_outputs(2535));
    layer4_outputs(2009) <= layer3_outputs(162);
    layer4_outputs(2010) <= layer3_outputs(581);
    layer4_outputs(2011) <= not(layer3_outputs(423)) or (layer3_outputs(1598));
    layer4_outputs(2012) <= '1';
    layer4_outputs(2013) <= (layer3_outputs(1932)) and not (layer3_outputs(1623));
    layer4_outputs(2014) <= not((layer3_outputs(2224)) and (layer3_outputs(2359)));
    layer4_outputs(2015) <= (layer3_outputs(841)) and not (layer3_outputs(2214));
    layer4_outputs(2016) <= layer3_outputs(1591);
    layer4_outputs(2017) <= layer3_outputs(1679);
    layer4_outputs(2018) <= not((layer3_outputs(200)) or (layer3_outputs(1276)));
    layer4_outputs(2019) <= (layer3_outputs(1320)) and not (layer3_outputs(2271));
    layer4_outputs(2020) <= (layer3_outputs(1837)) and (layer3_outputs(2012));
    layer4_outputs(2021) <= layer3_outputs(1696);
    layer4_outputs(2022) <= '0';
    layer4_outputs(2023) <= '1';
    layer4_outputs(2024) <= not((layer3_outputs(2156)) or (layer3_outputs(206)));
    layer4_outputs(2025) <= (layer3_outputs(2011)) and (layer3_outputs(997));
    layer4_outputs(2026) <= '0';
    layer4_outputs(2027) <= not((layer3_outputs(1154)) and (layer3_outputs(761)));
    layer4_outputs(2028) <= not(layer3_outputs(1363)) or (layer3_outputs(2137));
    layer4_outputs(2029) <= not((layer3_outputs(1947)) or (layer3_outputs(600)));
    layer4_outputs(2030) <= not(layer3_outputs(2336)) or (layer3_outputs(1361));
    layer4_outputs(2031) <= layer3_outputs(1765);
    layer4_outputs(2032) <= not(layer3_outputs(1558));
    layer4_outputs(2033) <= layer3_outputs(508);
    layer4_outputs(2034) <= (layer3_outputs(1120)) and not (layer3_outputs(2337));
    layer4_outputs(2035) <= not(layer3_outputs(1726)) or (layer3_outputs(1039));
    layer4_outputs(2036) <= not(layer3_outputs(1369));
    layer4_outputs(2037) <= not((layer3_outputs(1645)) and (layer3_outputs(2075)));
    layer4_outputs(2038) <= layer3_outputs(2043);
    layer4_outputs(2039) <= (layer3_outputs(1865)) xor (layer3_outputs(893));
    layer4_outputs(2040) <= not(layer3_outputs(114)) or (layer3_outputs(246));
    layer4_outputs(2041) <= layer3_outputs(2296);
    layer4_outputs(2042) <= (layer3_outputs(24)) and not (layer3_outputs(1993));
    layer4_outputs(2043) <= not(layer3_outputs(183));
    layer4_outputs(2044) <= layer3_outputs(1750);
    layer4_outputs(2045) <= layer3_outputs(847);
    layer4_outputs(2046) <= (layer3_outputs(1011)) and (layer3_outputs(1072));
    layer4_outputs(2047) <= not(layer3_outputs(2444)) or (layer3_outputs(279));
    layer4_outputs(2048) <= (layer3_outputs(497)) and not (layer3_outputs(1202));
    layer4_outputs(2049) <= not(layer3_outputs(2192)) or (layer3_outputs(151));
    layer4_outputs(2050) <= layer3_outputs(89);
    layer4_outputs(2051) <= not((layer3_outputs(355)) and (layer3_outputs(430)));
    layer4_outputs(2052) <= layer3_outputs(661);
    layer4_outputs(2053) <= not(layer3_outputs(2544));
    layer4_outputs(2054) <= (layer3_outputs(2008)) and not (layer3_outputs(650));
    layer4_outputs(2055) <= not(layer3_outputs(2085));
    layer4_outputs(2056) <= layer3_outputs(472);
    layer4_outputs(2057) <= not(layer3_outputs(1280)) or (layer3_outputs(1704));
    layer4_outputs(2058) <= '0';
    layer4_outputs(2059) <= '1';
    layer4_outputs(2060) <= not(layer3_outputs(802)) or (layer3_outputs(1007));
    layer4_outputs(2061) <= not(layer3_outputs(1507));
    layer4_outputs(2062) <= layer3_outputs(2335);
    layer4_outputs(2063) <= not(layer3_outputs(1723));
    layer4_outputs(2064) <= not(layer3_outputs(1578));
    layer4_outputs(2065) <= (layer3_outputs(651)) and not (layer3_outputs(127));
    layer4_outputs(2066) <= (layer3_outputs(1337)) and not (layer3_outputs(1138));
    layer4_outputs(2067) <= not(layer3_outputs(1509));
    layer4_outputs(2068) <= not(layer3_outputs(2211)) or (layer3_outputs(1878));
    layer4_outputs(2069) <= '1';
    layer4_outputs(2070) <= (layer3_outputs(885)) and not (layer3_outputs(800));
    layer4_outputs(2071) <= '0';
    layer4_outputs(2072) <= '0';
    layer4_outputs(2073) <= (layer3_outputs(38)) and not (layer3_outputs(57));
    layer4_outputs(2074) <= '0';
    layer4_outputs(2075) <= (layer3_outputs(1141)) and not (layer3_outputs(1219));
    layer4_outputs(2076) <= (layer3_outputs(1682)) and not (layer3_outputs(404));
    layer4_outputs(2077) <= layer3_outputs(1725);
    layer4_outputs(2078) <= '0';
    layer4_outputs(2079) <= not(layer3_outputs(2431)) or (layer3_outputs(1556));
    layer4_outputs(2080) <= layer3_outputs(2241);
    layer4_outputs(2081) <= not((layer3_outputs(496)) or (layer3_outputs(2263)));
    layer4_outputs(2082) <= not(layer3_outputs(1931)) or (layer3_outputs(1410));
    layer4_outputs(2083) <= not(layer3_outputs(1421)) or (layer3_outputs(664));
    layer4_outputs(2084) <= (layer3_outputs(940)) and not (layer3_outputs(358));
    layer4_outputs(2085) <= (layer3_outputs(1315)) and (layer3_outputs(2508));
    layer4_outputs(2086) <= layer3_outputs(1040);
    layer4_outputs(2087) <= not((layer3_outputs(1229)) and (layer3_outputs(728)));
    layer4_outputs(2088) <= not(layer3_outputs(1839)) or (layer3_outputs(1316));
    layer4_outputs(2089) <= not((layer3_outputs(1324)) xor (layer3_outputs(1449)));
    layer4_outputs(2090) <= (layer3_outputs(1219)) and not (layer3_outputs(1609));
    layer4_outputs(2091) <= (layer3_outputs(2491)) and not (layer3_outputs(577));
    layer4_outputs(2092) <= not((layer3_outputs(2087)) and (layer3_outputs(220)));
    layer4_outputs(2093) <= '1';
    layer4_outputs(2094) <= (layer3_outputs(840)) and not (layer3_outputs(1724));
    layer4_outputs(2095) <= layer3_outputs(1147);
    layer4_outputs(2096) <= layer3_outputs(1654);
    layer4_outputs(2097) <= not(layer3_outputs(1675));
    layer4_outputs(2098) <= not((layer3_outputs(177)) and (layer3_outputs(1977)));
    layer4_outputs(2099) <= '1';
    layer4_outputs(2100) <= layer3_outputs(1372);
    layer4_outputs(2101) <= layer3_outputs(1504);
    layer4_outputs(2102) <= (layer3_outputs(96)) or (layer3_outputs(1497));
    layer4_outputs(2103) <= layer3_outputs(1850);
    layer4_outputs(2104) <= layer3_outputs(2486);
    layer4_outputs(2105) <= not((layer3_outputs(17)) and (layer3_outputs(1114)));
    layer4_outputs(2106) <= layer3_outputs(2031);
    layer4_outputs(2107) <= layer3_outputs(2522);
    layer4_outputs(2108) <= not((layer3_outputs(1494)) and (layer3_outputs(1684)));
    layer4_outputs(2109) <= layer3_outputs(1401);
    layer4_outputs(2110) <= not(layer3_outputs(172));
    layer4_outputs(2111) <= layer3_outputs(1941);
    layer4_outputs(2112) <= not(layer3_outputs(846)) or (layer3_outputs(1468));
    layer4_outputs(2113) <= '1';
    layer4_outputs(2114) <= (layer3_outputs(2514)) and not (layer3_outputs(769));
    layer4_outputs(2115) <= layer3_outputs(2216);
    layer4_outputs(2116) <= layer3_outputs(1907);
    layer4_outputs(2117) <= (layer3_outputs(1552)) and not (layer3_outputs(1204));
    layer4_outputs(2118) <= not(layer3_outputs(225));
    layer4_outputs(2119) <= layer3_outputs(1258);
    layer4_outputs(2120) <= not(layer3_outputs(1845));
    layer4_outputs(2121) <= not(layer3_outputs(2142));
    layer4_outputs(2122) <= (layer3_outputs(787)) or (layer3_outputs(1230));
    layer4_outputs(2123) <= layer3_outputs(2471);
    layer4_outputs(2124) <= (layer3_outputs(1844)) and (layer3_outputs(1555));
    layer4_outputs(2125) <= (layer3_outputs(1715)) and not (layer3_outputs(2268));
    layer4_outputs(2126) <= layer3_outputs(1510);
    layer4_outputs(2127) <= not(layer3_outputs(1456));
    layer4_outputs(2128) <= layer3_outputs(1589);
    layer4_outputs(2129) <= layer3_outputs(1992);
    layer4_outputs(2130) <= not(layer3_outputs(2231));
    layer4_outputs(2131) <= not((layer3_outputs(105)) xor (layer3_outputs(193)));
    layer4_outputs(2132) <= layer3_outputs(692);
    layer4_outputs(2133) <= layer3_outputs(1573);
    layer4_outputs(2134) <= layer3_outputs(1872);
    layer4_outputs(2135) <= (layer3_outputs(2002)) and not (layer3_outputs(43));
    layer4_outputs(2136) <= not(layer3_outputs(142));
    layer4_outputs(2137) <= (layer3_outputs(2204)) and not (layer3_outputs(678));
    layer4_outputs(2138) <= (layer3_outputs(235)) and (layer3_outputs(1820));
    layer4_outputs(2139) <= layer3_outputs(1313);
    layer4_outputs(2140) <= layer3_outputs(1620);
    layer4_outputs(2141) <= not(layer3_outputs(1294));
    layer4_outputs(2142) <= (layer3_outputs(1254)) and (layer3_outputs(4));
    layer4_outputs(2143) <= not(layer3_outputs(759)) or (layer3_outputs(99));
    layer4_outputs(2144) <= not(layer3_outputs(703)) or (layer3_outputs(1481));
    layer4_outputs(2145) <= '0';
    layer4_outputs(2146) <= '1';
    layer4_outputs(2147) <= not((layer3_outputs(878)) or (layer3_outputs(2101)));
    layer4_outputs(2148) <= layer3_outputs(624);
    layer4_outputs(2149) <= not(layer3_outputs(345)) or (layer3_outputs(2497));
    layer4_outputs(2150) <= layer3_outputs(1689);
    layer4_outputs(2151) <= not(layer3_outputs(1051)) or (layer3_outputs(1188));
    layer4_outputs(2152) <= not((layer3_outputs(1468)) and (layer3_outputs(1050)));
    layer4_outputs(2153) <= '1';
    layer4_outputs(2154) <= not(layer3_outputs(1679));
    layer4_outputs(2155) <= not(layer3_outputs(2217)) or (layer3_outputs(902));
    layer4_outputs(2156) <= not(layer3_outputs(1914)) or (layer3_outputs(2049));
    layer4_outputs(2157) <= (layer3_outputs(466)) and not (layer3_outputs(1772));
    layer4_outputs(2158) <= not((layer3_outputs(2376)) or (layer3_outputs(983)));
    layer4_outputs(2159) <= '0';
    layer4_outputs(2160) <= not(layer3_outputs(2541)) or (layer3_outputs(61));
    layer4_outputs(2161) <= '1';
    layer4_outputs(2162) <= not(layer3_outputs(46)) or (layer3_outputs(1369));
    layer4_outputs(2163) <= not(layer3_outputs(1356));
    layer4_outputs(2164) <= (layer3_outputs(2509)) and (layer3_outputs(1428));
    layer4_outputs(2165) <= (layer3_outputs(1396)) and (layer3_outputs(183));
    layer4_outputs(2166) <= layer3_outputs(1540);
    layer4_outputs(2167) <= not(layer3_outputs(449)) or (layer3_outputs(24));
    layer4_outputs(2168) <= layer3_outputs(1064);
    layer4_outputs(2169) <= not((layer3_outputs(320)) and (layer3_outputs(1163)));
    layer4_outputs(2170) <= not(layer3_outputs(2112)) or (layer3_outputs(1738));
    layer4_outputs(2171) <= '0';
    layer4_outputs(2172) <= '1';
    layer4_outputs(2173) <= not(layer3_outputs(2143));
    layer4_outputs(2174) <= '0';
    layer4_outputs(2175) <= layer3_outputs(612);
    layer4_outputs(2176) <= '1';
    layer4_outputs(2177) <= (layer3_outputs(121)) and (layer3_outputs(708));
    layer4_outputs(2178) <= layer3_outputs(1029);
    layer4_outputs(2179) <= not(layer3_outputs(1642)) or (layer3_outputs(2100));
    layer4_outputs(2180) <= not(layer3_outputs(1362)) or (layer3_outputs(1482));
    layer4_outputs(2181) <= layer3_outputs(366);
    layer4_outputs(2182) <= (layer3_outputs(789)) xor (layer3_outputs(1736));
    layer4_outputs(2183) <= not(layer3_outputs(407)) or (layer3_outputs(884));
    layer4_outputs(2184) <= layer3_outputs(359);
    layer4_outputs(2185) <= layer3_outputs(133);
    layer4_outputs(2186) <= '1';
    layer4_outputs(2187) <= (layer3_outputs(814)) and not (layer3_outputs(770));
    layer4_outputs(2188) <= '0';
    layer4_outputs(2189) <= layer3_outputs(1104);
    layer4_outputs(2190) <= (layer3_outputs(610)) and (layer3_outputs(1222));
    layer4_outputs(2191) <= (layer3_outputs(1217)) xor (layer3_outputs(53));
    layer4_outputs(2192) <= '1';
    layer4_outputs(2193) <= (layer3_outputs(462)) and (layer3_outputs(1945));
    layer4_outputs(2194) <= layer3_outputs(389);
    layer4_outputs(2195) <= not((layer3_outputs(1350)) or (layer3_outputs(776)));
    layer4_outputs(2196) <= (layer3_outputs(2212)) and not (layer3_outputs(2132));
    layer4_outputs(2197) <= not((layer3_outputs(2407)) or (layer3_outputs(186)));
    layer4_outputs(2198) <= not(layer3_outputs(1247));
    layer4_outputs(2199) <= (layer3_outputs(1839)) or (layer3_outputs(304));
    layer4_outputs(2200) <= not((layer3_outputs(30)) or (layer3_outputs(1320)));
    layer4_outputs(2201) <= (layer3_outputs(817)) or (layer3_outputs(924));
    layer4_outputs(2202) <= (layer3_outputs(2110)) xor (layer3_outputs(1554));
    layer4_outputs(2203) <= (layer3_outputs(2439)) and (layer3_outputs(102));
    layer4_outputs(2204) <= layer3_outputs(1357);
    layer4_outputs(2205) <= not(layer3_outputs(888));
    layer4_outputs(2206) <= (layer3_outputs(1079)) and not (layer3_outputs(1948));
    layer4_outputs(2207) <= layer3_outputs(2155);
    layer4_outputs(2208) <= '1';
    layer4_outputs(2209) <= layer3_outputs(819);
    layer4_outputs(2210) <= not(layer3_outputs(756));
    layer4_outputs(2211) <= not(layer3_outputs(222));
    layer4_outputs(2212) <= (layer3_outputs(2372)) and not (layer3_outputs(1197));
    layer4_outputs(2213) <= layer3_outputs(2371);
    layer4_outputs(2214) <= layer3_outputs(1107);
    layer4_outputs(2215) <= not(layer3_outputs(2149));
    layer4_outputs(2216) <= (layer3_outputs(1495)) and not (layer3_outputs(1568));
    layer4_outputs(2217) <= not((layer3_outputs(1819)) and (layer3_outputs(1004)));
    layer4_outputs(2218) <= not((layer3_outputs(23)) or (layer3_outputs(696)));
    layer4_outputs(2219) <= (layer3_outputs(87)) and (layer3_outputs(54));
    layer4_outputs(2220) <= not((layer3_outputs(1882)) or (layer3_outputs(1824)));
    layer4_outputs(2221) <= layer3_outputs(2045);
    layer4_outputs(2222) <= layer3_outputs(157);
    layer4_outputs(2223) <= layer3_outputs(2019);
    layer4_outputs(2224) <= (layer3_outputs(1831)) and not (layer3_outputs(1828));
    layer4_outputs(2225) <= (layer3_outputs(1212)) or (layer3_outputs(375));
    layer4_outputs(2226) <= not((layer3_outputs(1385)) and (layer3_outputs(1944)));
    layer4_outputs(2227) <= not(layer3_outputs(97));
    layer4_outputs(2228) <= '1';
    layer4_outputs(2229) <= not((layer3_outputs(238)) xor (layer3_outputs(2438)));
    layer4_outputs(2230) <= not((layer3_outputs(862)) and (layer3_outputs(834)));
    layer4_outputs(2231) <= not(layer3_outputs(1311)) or (layer3_outputs(83));
    layer4_outputs(2232) <= not(layer3_outputs(112));
    layer4_outputs(2233) <= not(layer3_outputs(1972));
    layer4_outputs(2234) <= layer3_outputs(1911);
    layer4_outputs(2235) <= (layer3_outputs(789)) and (layer3_outputs(1242));
    layer4_outputs(2236) <= not(layer3_outputs(957));
    layer4_outputs(2237) <= not(layer3_outputs(1099));
    layer4_outputs(2238) <= layer3_outputs(457);
    layer4_outputs(2239) <= not((layer3_outputs(2168)) xor (layer3_outputs(2219)));
    layer4_outputs(2240) <= not((layer3_outputs(65)) xor (layer3_outputs(1437)));
    layer4_outputs(2241) <= not((layer3_outputs(1335)) and (layer3_outputs(2470)));
    layer4_outputs(2242) <= not(layer3_outputs(987)) or (layer3_outputs(524));
    layer4_outputs(2243) <= not((layer3_outputs(493)) xor (layer3_outputs(2500)));
    layer4_outputs(2244) <= (layer3_outputs(1544)) xor (layer3_outputs(1346));
    layer4_outputs(2245) <= not(layer3_outputs(2556)) or (layer3_outputs(2000));
    layer4_outputs(2246) <= not(layer3_outputs(2431));
    layer4_outputs(2247) <= not(layer3_outputs(598)) or (layer3_outputs(1384));
    layer4_outputs(2248) <= (layer3_outputs(1300)) and not (layer3_outputs(1943));
    layer4_outputs(2249) <= (layer3_outputs(1674)) and (layer3_outputs(296));
    layer4_outputs(2250) <= layer3_outputs(1797);
    layer4_outputs(2251) <= not((layer3_outputs(164)) or (layer3_outputs(122)));
    layer4_outputs(2252) <= layer3_outputs(2518);
    layer4_outputs(2253) <= not((layer3_outputs(1110)) xor (layer3_outputs(1423)));
    layer4_outputs(2254) <= not(layer3_outputs(2471));
    layer4_outputs(2255) <= (layer3_outputs(103)) and not (layer3_outputs(120));
    layer4_outputs(2256) <= not(layer3_outputs(506));
    layer4_outputs(2257) <= layer3_outputs(1904);
    layer4_outputs(2258) <= (layer3_outputs(645)) xor (layer3_outputs(1166));
    layer4_outputs(2259) <= '0';
    layer4_outputs(2260) <= not(layer3_outputs(874));
    layer4_outputs(2261) <= layer3_outputs(370);
    layer4_outputs(2262) <= not(layer3_outputs(1074));
    layer4_outputs(2263) <= layer3_outputs(1649);
    layer4_outputs(2264) <= (layer3_outputs(31)) and (layer3_outputs(1180));
    layer4_outputs(2265) <= not(layer3_outputs(1628)) or (layer3_outputs(2296));
    layer4_outputs(2266) <= not(layer3_outputs(613));
    layer4_outputs(2267) <= not(layer3_outputs(2035));
    layer4_outputs(2268) <= layer3_outputs(2146);
    layer4_outputs(2269) <= layer3_outputs(1686);
    layer4_outputs(2270) <= not(layer3_outputs(808)) or (layer3_outputs(536));
    layer4_outputs(2271) <= not(layer3_outputs(1545));
    layer4_outputs(2272) <= layer3_outputs(568);
    layer4_outputs(2273) <= (layer3_outputs(2181)) and not (layer3_outputs(450));
    layer4_outputs(2274) <= not(layer3_outputs(1386));
    layer4_outputs(2275) <= not(layer3_outputs(917));
    layer4_outputs(2276) <= not(layer3_outputs(534)) or (layer3_outputs(192));
    layer4_outputs(2277) <= layer3_outputs(1749);
    layer4_outputs(2278) <= '1';
    layer4_outputs(2279) <= '0';
    layer4_outputs(2280) <= layer3_outputs(752);
    layer4_outputs(2281) <= not(layer3_outputs(2506)) or (layer3_outputs(1257));
    layer4_outputs(2282) <= layer3_outputs(1829);
    layer4_outputs(2283) <= layer3_outputs(1214);
    layer4_outputs(2284) <= not(layer3_outputs(2102));
    layer4_outputs(2285) <= not(layer3_outputs(1768)) or (layer3_outputs(1283));
    layer4_outputs(2286) <= not((layer3_outputs(2139)) and (layer3_outputs(2080)));
    layer4_outputs(2287) <= '1';
    layer4_outputs(2288) <= '1';
    layer4_outputs(2289) <= not(layer3_outputs(704));
    layer4_outputs(2290) <= not(layer3_outputs(2377)) or (layer3_outputs(2435));
    layer4_outputs(2291) <= (layer3_outputs(2558)) or (layer3_outputs(16));
    layer4_outputs(2292) <= layer3_outputs(1126);
    layer4_outputs(2293) <= layer3_outputs(1301);
    layer4_outputs(2294) <= not(layer3_outputs(2228));
    layer4_outputs(2295) <= (layer3_outputs(1898)) and not (layer3_outputs(1231));
    layer4_outputs(2296) <= not(layer3_outputs(352)) or (layer3_outputs(442));
    layer4_outputs(2297) <= not((layer3_outputs(925)) and (layer3_outputs(993)));
    layer4_outputs(2298) <= layer3_outputs(1332);
    layer4_outputs(2299) <= '1';
    layer4_outputs(2300) <= not(layer3_outputs(264));
    layer4_outputs(2301) <= not(layer3_outputs(1004));
    layer4_outputs(2302) <= (layer3_outputs(1520)) or (layer3_outputs(1238));
    layer4_outputs(2303) <= not(layer3_outputs(1599));
    layer4_outputs(2304) <= not((layer3_outputs(1991)) or (layer3_outputs(1835)));
    layer4_outputs(2305) <= (layer3_outputs(553)) or (layer3_outputs(1455));
    layer4_outputs(2306) <= (layer3_outputs(1584)) and not (layer3_outputs(1783));
    layer4_outputs(2307) <= not((layer3_outputs(900)) and (layer3_outputs(2087)));
    layer4_outputs(2308) <= layer3_outputs(325);
    layer4_outputs(2309) <= (layer3_outputs(721)) or (layer3_outputs(106));
    layer4_outputs(2310) <= (layer3_outputs(2461)) and not (layer3_outputs(1559));
    layer4_outputs(2311) <= (layer3_outputs(1758)) or (layer3_outputs(589));
    layer4_outputs(2312) <= layer3_outputs(1856);
    layer4_outputs(2313) <= not((layer3_outputs(1736)) and (layer3_outputs(1794)));
    layer4_outputs(2314) <= layer3_outputs(618);
    layer4_outputs(2315) <= not(layer3_outputs(1487)) or (layer3_outputs(963));
    layer4_outputs(2316) <= (layer3_outputs(1090)) and not (layer3_outputs(2480));
    layer4_outputs(2317) <= not((layer3_outputs(919)) and (layer3_outputs(1569)));
    layer4_outputs(2318) <= not((layer3_outputs(1302)) and (layer3_outputs(674)));
    layer4_outputs(2319) <= (layer3_outputs(1841)) and not (layer3_outputs(529));
    layer4_outputs(2320) <= (layer3_outputs(250)) and (layer3_outputs(1260));
    layer4_outputs(2321) <= (layer3_outputs(2064)) and not (layer3_outputs(1373));
    layer4_outputs(2322) <= not(layer3_outputs(2357)) or (layer3_outputs(322));
    layer4_outputs(2323) <= not(layer3_outputs(1602));
    layer4_outputs(2324) <= (layer3_outputs(146)) or (layer3_outputs(2238));
    layer4_outputs(2325) <= not(layer3_outputs(1700));
    layer4_outputs(2326) <= (layer3_outputs(2224)) and (layer3_outputs(1402));
    layer4_outputs(2327) <= not(layer3_outputs(0));
    layer4_outputs(2328) <= (layer3_outputs(412)) and not (layer3_outputs(606));
    layer4_outputs(2329) <= '1';
    layer4_outputs(2330) <= (layer3_outputs(477)) and not (layer3_outputs(502));
    layer4_outputs(2331) <= (layer3_outputs(56)) or (layer3_outputs(1330));
    layer4_outputs(2332) <= (layer3_outputs(25)) and not (layer3_outputs(2467));
    layer4_outputs(2333) <= not(layer3_outputs(2305));
    layer4_outputs(2334) <= not(layer3_outputs(2532)) or (layer3_outputs(367));
    layer4_outputs(2335) <= not(layer3_outputs(2258)) or (layer3_outputs(1070));
    layer4_outputs(2336) <= not(layer3_outputs(10));
    layer4_outputs(2337) <= not(layer3_outputs(686));
    layer4_outputs(2338) <= not((layer3_outputs(1020)) or (layer3_outputs(276)));
    layer4_outputs(2339) <= not(layer3_outputs(2258)) or (layer3_outputs(718));
    layer4_outputs(2340) <= (layer3_outputs(435)) and not (layer3_outputs(2234));
    layer4_outputs(2341) <= (layer3_outputs(317)) and not (layer3_outputs(1939));
    layer4_outputs(2342) <= not(layer3_outputs(1356));
    layer4_outputs(2343) <= (layer3_outputs(45)) and not (layer3_outputs(595));
    layer4_outputs(2344) <= not(layer3_outputs(1807)) or (layer3_outputs(1213));
    layer4_outputs(2345) <= not(layer3_outputs(1068)) or (layer3_outputs(172));
    layer4_outputs(2346) <= not((layer3_outputs(300)) or (layer3_outputs(930)));
    layer4_outputs(2347) <= not(layer3_outputs(1884)) or (layer3_outputs(1024));
    layer4_outputs(2348) <= not(layer3_outputs(1720));
    layer4_outputs(2349) <= not(layer3_outputs(1499));
    layer4_outputs(2350) <= not(layer3_outputs(80)) or (layer3_outputs(1810));
    layer4_outputs(2351) <= (layer3_outputs(1458)) and not (layer3_outputs(158));
    layer4_outputs(2352) <= (layer3_outputs(400)) and (layer3_outputs(352));
    layer4_outputs(2353) <= not(layer3_outputs(1341));
    layer4_outputs(2354) <= not(layer3_outputs(407)) or (layer3_outputs(2501));
    layer4_outputs(2355) <= not((layer3_outputs(1448)) and (layer3_outputs(1475)));
    layer4_outputs(2356) <= layer3_outputs(2209);
    layer4_outputs(2357) <= not(layer3_outputs(997)) or (layer3_outputs(1507));
    layer4_outputs(2358) <= not(layer3_outputs(631));
    layer4_outputs(2359) <= layer3_outputs(1314);
    layer4_outputs(2360) <= not(layer3_outputs(1340));
    layer4_outputs(2361) <= (layer3_outputs(2121)) or (layer3_outputs(1580));
    layer4_outputs(2362) <= not((layer3_outputs(1382)) xor (layer3_outputs(2273)));
    layer4_outputs(2363) <= not(layer3_outputs(1184));
    layer4_outputs(2364) <= not(layer3_outputs(2559));
    layer4_outputs(2365) <= layer3_outputs(1237);
    layer4_outputs(2366) <= not(layer3_outputs(1707));
    layer4_outputs(2367) <= (layer3_outputs(1162)) and (layer3_outputs(898));
    layer4_outputs(2368) <= not(layer3_outputs(2125));
    layer4_outputs(2369) <= not(layer3_outputs(431));
    layer4_outputs(2370) <= not((layer3_outputs(377)) xor (layer3_outputs(1864)));
    layer4_outputs(2371) <= not(layer3_outputs(1234));
    layer4_outputs(2372) <= not(layer3_outputs(2548));
    layer4_outputs(2373) <= (layer3_outputs(156)) and not (layer3_outputs(393));
    layer4_outputs(2374) <= not(layer3_outputs(363));
    layer4_outputs(2375) <= not((layer3_outputs(2028)) and (layer3_outputs(559)));
    layer4_outputs(2376) <= (layer3_outputs(1207)) and not (layer3_outputs(630));
    layer4_outputs(2377) <= layer3_outputs(2391);
    layer4_outputs(2378) <= not(layer3_outputs(2477)) or (layer3_outputs(1704));
    layer4_outputs(2379) <= not(layer3_outputs(1625));
    layer4_outputs(2380) <= '0';
    layer4_outputs(2381) <= (layer3_outputs(1908)) or (layer3_outputs(1640));
    layer4_outputs(2382) <= not(layer3_outputs(1091)) or (layer3_outputs(1040));
    layer4_outputs(2383) <= '1';
    layer4_outputs(2384) <= not(layer3_outputs(71)) or (layer3_outputs(2082));
    layer4_outputs(2385) <= (layer3_outputs(1209)) and (layer3_outputs(1486));
    layer4_outputs(2386) <= not(layer3_outputs(1069));
    layer4_outputs(2387) <= layer3_outputs(1722);
    layer4_outputs(2388) <= '1';
    layer4_outputs(2389) <= not(layer3_outputs(1415));
    layer4_outputs(2390) <= '0';
    layer4_outputs(2391) <= layer3_outputs(729);
    layer4_outputs(2392) <= (layer3_outputs(1859)) or (layer3_outputs(1842));
    layer4_outputs(2393) <= (layer3_outputs(1643)) and not (layer3_outputs(2079));
    layer4_outputs(2394) <= not(layer3_outputs(2221));
    layer4_outputs(2395) <= not(layer3_outputs(2042)) or (layer3_outputs(1427));
    layer4_outputs(2396) <= '0';
    layer4_outputs(2397) <= (layer3_outputs(1950)) and not (layer3_outputs(336));
    layer4_outputs(2398) <= not((layer3_outputs(1407)) and (layer3_outputs(2366)));
    layer4_outputs(2399) <= not(layer3_outputs(681));
    layer4_outputs(2400) <= '1';
    layer4_outputs(2401) <= (layer3_outputs(1406)) or (layer3_outputs(2439));
    layer4_outputs(2402) <= not(layer3_outputs(757));
    layer4_outputs(2403) <= layer3_outputs(1441);
    layer4_outputs(2404) <= not(layer3_outputs(2385));
    layer4_outputs(2405) <= not(layer3_outputs(359));
    layer4_outputs(2406) <= '0';
    layer4_outputs(2407) <= not(layer3_outputs(1450));
    layer4_outputs(2408) <= not((layer3_outputs(809)) xor (layer3_outputs(642)));
    layer4_outputs(2409) <= not((layer3_outputs(1259)) or (layer3_outputs(628)));
    layer4_outputs(2410) <= (layer3_outputs(1357)) and not (layer3_outputs(1565));
    layer4_outputs(2411) <= not(layer3_outputs(1958));
    layer4_outputs(2412) <= (layer3_outputs(1422)) and not (layer3_outputs(1342));
    layer4_outputs(2413) <= not((layer3_outputs(1729)) xor (layer3_outputs(116)));
    layer4_outputs(2414) <= not((layer3_outputs(2406)) and (layer3_outputs(261)));
    layer4_outputs(2415) <= '1';
    layer4_outputs(2416) <= (layer3_outputs(663)) and not (layer3_outputs(410));
    layer4_outputs(2417) <= layer3_outputs(2189);
    layer4_outputs(2418) <= layer3_outputs(322);
    layer4_outputs(2419) <= not(layer3_outputs(2402)) or (layer3_outputs(2557));
    layer4_outputs(2420) <= not(layer3_outputs(2294));
    layer4_outputs(2421) <= (layer3_outputs(1387)) xor (layer3_outputs(853));
    layer4_outputs(2422) <= layer3_outputs(122);
    layer4_outputs(2423) <= not((layer3_outputs(2482)) and (layer3_outputs(1738)));
    layer4_outputs(2424) <= not((layer3_outputs(2181)) or (layer3_outputs(1914)));
    layer4_outputs(2425) <= (layer3_outputs(837)) and (layer3_outputs(245));
    layer4_outputs(2426) <= layer3_outputs(2103);
    layer4_outputs(2427) <= '1';
    layer4_outputs(2428) <= not(layer3_outputs(1527));
    layer4_outputs(2429) <= (layer3_outputs(580)) and not (layer3_outputs(1411));
    layer4_outputs(2430) <= not((layer3_outputs(2419)) or (layer3_outputs(2510)));
    layer4_outputs(2431) <= (layer3_outputs(667)) and not (layer3_outputs(251));
    layer4_outputs(2432) <= (layer3_outputs(264)) and not (layer3_outputs(1089));
    layer4_outputs(2433) <= not((layer3_outputs(1946)) or (layer3_outputs(2450)));
    layer4_outputs(2434) <= (layer3_outputs(591)) xor (layer3_outputs(478));
    layer4_outputs(2435) <= not(layer3_outputs(1613));
    layer4_outputs(2436) <= not((layer3_outputs(1993)) or (layer3_outputs(441)));
    layer4_outputs(2437) <= not(layer3_outputs(952));
    layer4_outputs(2438) <= not(layer3_outputs(2209));
    layer4_outputs(2439) <= (layer3_outputs(2145)) and not (layer3_outputs(866));
    layer4_outputs(2440) <= layer3_outputs(659);
    layer4_outputs(2441) <= (layer3_outputs(2440)) or (layer3_outputs(474));
    layer4_outputs(2442) <= not(layer3_outputs(287)) or (layer3_outputs(2422));
    layer4_outputs(2443) <= layer3_outputs(2546);
    layer4_outputs(2444) <= (layer3_outputs(1482)) and (layer3_outputs(508));
    layer4_outputs(2445) <= (layer3_outputs(2368)) or (layer3_outputs(2306));
    layer4_outputs(2446) <= (layer3_outputs(2093)) or (layer3_outputs(20));
    layer4_outputs(2447) <= layer3_outputs(2485);
    layer4_outputs(2448) <= (layer3_outputs(751)) xor (layer3_outputs(1587));
    layer4_outputs(2449) <= (layer3_outputs(2510)) and (layer3_outputs(627));
    layer4_outputs(2450) <= not(layer3_outputs(1496)) or (layer3_outputs(2062));
    layer4_outputs(2451) <= layer3_outputs(1883);
    layer4_outputs(2452) <= not(layer3_outputs(1713));
    layer4_outputs(2453) <= not(layer3_outputs(2276));
    layer4_outputs(2454) <= (layer3_outputs(80)) and not (layer3_outputs(2186));
    layer4_outputs(2455) <= (layer3_outputs(554)) and not (layer3_outputs(368));
    layer4_outputs(2456) <= (layer3_outputs(864)) and not (layer3_outputs(26));
    layer4_outputs(2457) <= '0';
    layer4_outputs(2458) <= not(layer3_outputs(487));
    layer4_outputs(2459) <= '0';
    layer4_outputs(2460) <= '1';
    layer4_outputs(2461) <= layer3_outputs(124);
    layer4_outputs(2462) <= layer3_outputs(1530);
    layer4_outputs(2463) <= '0';
    layer4_outputs(2464) <= not(layer3_outputs(1109)) or (layer3_outputs(212));
    layer4_outputs(2465) <= not(layer3_outputs(1226));
    layer4_outputs(2466) <= (layer3_outputs(782)) and not (layer3_outputs(77));
    layer4_outputs(2467) <= '0';
    layer4_outputs(2468) <= layer3_outputs(349);
    layer4_outputs(2469) <= not(layer3_outputs(119));
    layer4_outputs(2470) <= (layer3_outputs(326)) and (layer3_outputs(2257));
    layer4_outputs(2471) <= layer3_outputs(434);
    layer4_outputs(2472) <= (layer3_outputs(1200)) and (layer3_outputs(2531));
    layer4_outputs(2473) <= (layer3_outputs(1874)) and not (layer3_outputs(2435));
    layer4_outputs(2474) <= not(layer3_outputs(461));
    layer4_outputs(2475) <= not(layer3_outputs(1215)) or (layer3_outputs(2023));
    layer4_outputs(2476) <= '1';
    layer4_outputs(2477) <= layer3_outputs(2119);
    layer4_outputs(2478) <= (layer3_outputs(1840)) or (layer3_outputs(20));
    layer4_outputs(2479) <= (layer3_outputs(2482)) and not (layer3_outputs(5));
    layer4_outputs(2480) <= (layer3_outputs(2185)) and (layer3_outputs(2243));
    layer4_outputs(2481) <= layer3_outputs(433);
    layer4_outputs(2482) <= (layer3_outputs(1235)) and (layer3_outputs(2364));
    layer4_outputs(2483) <= layer3_outputs(569);
    layer4_outputs(2484) <= not(layer3_outputs(2512)) or (layer3_outputs(1012));
    layer4_outputs(2485) <= layer3_outputs(406);
    layer4_outputs(2486) <= not(layer3_outputs(495)) or (layer3_outputs(131));
    layer4_outputs(2487) <= not(layer3_outputs(1344));
    layer4_outputs(2488) <= layer3_outputs(1081);
    layer4_outputs(2489) <= not(layer3_outputs(1875));
    layer4_outputs(2490) <= layer3_outputs(1372);
    layer4_outputs(2491) <= not(layer3_outputs(1719)) or (layer3_outputs(1571));
    layer4_outputs(2492) <= (layer3_outputs(1982)) or (layer3_outputs(2414));
    layer4_outputs(2493) <= not(layer3_outputs(1984));
    layer4_outputs(2494) <= not(layer3_outputs(823));
    layer4_outputs(2495) <= layer3_outputs(1987);
    layer4_outputs(2496) <= (layer3_outputs(1239)) and not (layer3_outputs(1575));
    layer4_outputs(2497) <= layer3_outputs(395);
    layer4_outputs(2498) <= not(layer3_outputs(544));
    layer4_outputs(2499) <= '0';
    layer4_outputs(2500) <= (layer3_outputs(817)) and (layer3_outputs(2201));
    layer4_outputs(2501) <= '0';
    layer4_outputs(2502) <= (layer3_outputs(760)) or (layer3_outputs(104));
    layer4_outputs(2503) <= layer3_outputs(346);
    layer4_outputs(2504) <= not(layer3_outputs(1702)) or (layer3_outputs(2223));
    layer4_outputs(2505) <= (layer3_outputs(523)) xor (layer3_outputs(948));
    layer4_outputs(2506) <= (layer3_outputs(205)) and not (layer3_outputs(568));
    layer4_outputs(2507) <= not(layer3_outputs(826)) or (layer3_outputs(2266));
    layer4_outputs(2508) <= not(layer3_outputs(451)) or (layer3_outputs(723));
    layer4_outputs(2509) <= '0';
    layer4_outputs(2510) <= not(layer3_outputs(1814));
    layer4_outputs(2511) <= not(layer3_outputs(2527));
    layer4_outputs(2512) <= (layer3_outputs(2088)) and not (layer3_outputs(101));
    layer4_outputs(2513) <= not(layer3_outputs(1019));
    layer4_outputs(2514) <= layer3_outputs(2300);
    layer4_outputs(2515) <= '1';
    layer4_outputs(2516) <= (layer3_outputs(1935)) xor (layer3_outputs(1398));
    layer4_outputs(2517) <= '0';
    layer4_outputs(2518) <= layer3_outputs(2376);
    layer4_outputs(2519) <= not(layer3_outputs(2315));
    layer4_outputs(2520) <= '0';
    layer4_outputs(2521) <= '1';
    layer4_outputs(2522) <= '1';
    layer4_outputs(2523) <= not(layer3_outputs(1183));
    layer4_outputs(2524) <= not(layer3_outputs(1310));
    layer4_outputs(2525) <= layer3_outputs(825);
    layer4_outputs(2526) <= layer3_outputs(712);
    layer4_outputs(2527) <= not(layer3_outputs(1521));
    layer4_outputs(2528) <= layer3_outputs(2462);
    layer4_outputs(2529) <= layer3_outputs(2057);
    layer4_outputs(2530) <= not(layer3_outputs(2110)) or (layer3_outputs(2416));
    layer4_outputs(2531) <= '1';
    layer4_outputs(2532) <= not(layer3_outputs(1926));
    layer4_outputs(2533) <= not((layer3_outputs(873)) and (layer3_outputs(548)));
    layer4_outputs(2534) <= layer3_outputs(2018);
    layer4_outputs(2535) <= not((layer3_outputs(715)) xor (layer3_outputs(1980)));
    layer4_outputs(2536) <= layer3_outputs(1164);
    layer4_outputs(2537) <= (layer3_outputs(1967)) and (layer3_outputs(185));
    layer4_outputs(2538) <= layer3_outputs(1378);
    layer4_outputs(2539) <= not(layer3_outputs(1698)) or (layer3_outputs(2226));
    layer4_outputs(2540) <= not(layer3_outputs(2237)) or (layer3_outputs(2394));
    layer4_outputs(2541) <= layer3_outputs(1571);
    layer4_outputs(2542) <= not(layer3_outputs(1516));
    layer4_outputs(2543) <= (layer3_outputs(1159)) and (layer3_outputs(2283));
    layer4_outputs(2544) <= '0';
    layer4_outputs(2545) <= not((layer3_outputs(1615)) and (layer3_outputs(911)));
    layer4_outputs(2546) <= not((layer3_outputs(1176)) or (layer3_outputs(2190)));
    layer4_outputs(2547) <= (layer3_outputs(1905)) xor (layer3_outputs(1557));
    layer4_outputs(2548) <= not(layer3_outputs(1424)) or (layer3_outputs(1459));
    layer4_outputs(2549) <= '1';
    layer4_outputs(2550) <= not((layer3_outputs(2467)) and (layer3_outputs(2105)));
    layer4_outputs(2551) <= '1';
    layer4_outputs(2552) <= layer3_outputs(504);
    layer4_outputs(2553) <= not(layer3_outputs(1210)) or (layer3_outputs(274));
    layer4_outputs(2554) <= layer3_outputs(2160);
    layer4_outputs(2555) <= not(layer3_outputs(954)) or (layer3_outputs(1246));
    layer4_outputs(2556) <= (layer3_outputs(1689)) and not (layer3_outputs(2429));
    layer4_outputs(2557) <= not((layer3_outputs(687)) and (layer3_outputs(38)));
    layer4_outputs(2558) <= not(layer3_outputs(150));
    layer4_outputs(2559) <= not(layer3_outputs(2490));
    layer5_outputs(0) <= '0';
    layer5_outputs(1) <= (layer4_outputs(1688)) and not (layer4_outputs(917));
    layer5_outputs(2) <= not(layer4_outputs(2180));
    layer5_outputs(3) <= not(layer4_outputs(551));
    layer5_outputs(4) <= not(layer4_outputs(1263)) or (layer4_outputs(965));
    layer5_outputs(5) <= layer4_outputs(1635);
    layer5_outputs(6) <= not((layer4_outputs(740)) or (layer4_outputs(1034)));
    layer5_outputs(7) <= not(layer4_outputs(2426));
    layer5_outputs(8) <= not(layer4_outputs(451));
    layer5_outputs(9) <= layer4_outputs(1278);
    layer5_outputs(10) <= '0';
    layer5_outputs(11) <= not(layer4_outputs(667)) or (layer4_outputs(889));
    layer5_outputs(12) <= layer4_outputs(688);
    layer5_outputs(13) <= (layer4_outputs(1150)) and not (layer4_outputs(1041));
    layer5_outputs(14) <= (layer4_outputs(581)) and not (layer4_outputs(1541));
    layer5_outputs(15) <= not(layer4_outputs(384)) or (layer4_outputs(1135));
    layer5_outputs(16) <= not(layer4_outputs(1169)) or (layer4_outputs(6));
    layer5_outputs(17) <= (layer4_outputs(1191)) and not (layer4_outputs(790));
    layer5_outputs(18) <= layer4_outputs(370);
    layer5_outputs(19) <= layer4_outputs(105);
    layer5_outputs(20) <= (layer4_outputs(2327)) xor (layer4_outputs(1579));
    layer5_outputs(21) <= not((layer4_outputs(1583)) or (layer4_outputs(549)));
    layer5_outputs(22) <= not(layer4_outputs(1574));
    layer5_outputs(23) <= (layer4_outputs(2392)) and not (layer4_outputs(343));
    layer5_outputs(24) <= layer4_outputs(926);
    layer5_outputs(25) <= not(layer4_outputs(507));
    layer5_outputs(26) <= (layer4_outputs(2301)) or (layer4_outputs(2373));
    layer5_outputs(27) <= not((layer4_outputs(1758)) xor (layer4_outputs(1021)));
    layer5_outputs(28) <= layer4_outputs(2333);
    layer5_outputs(29) <= not((layer4_outputs(1927)) or (layer4_outputs(255)));
    layer5_outputs(30) <= layer4_outputs(2371);
    layer5_outputs(31) <= (layer4_outputs(1797)) and (layer4_outputs(1517));
    layer5_outputs(32) <= not(layer4_outputs(113));
    layer5_outputs(33) <= layer4_outputs(406);
    layer5_outputs(34) <= layer4_outputs(1206);
    layer5_outputs(35) <= (layer4_outputs(2551)) and not (layer4_outputs(68));
    layer5_outputs(36) <= not(layer4_outputs(1404));
    layer5_outputs(37) <= layer4_outputs(678);
    layer5_outputs(38) <= layer4_outputs(1197);
    layer5_outputs(39) <= '1';
    layer5_outputs(40) <= layer4_outputs(2236);
    layer5_outputs(41) <= layer4_outputs(1877);
    layer5_outputs(42) <= not(layer4_outputs(2371));
    layer5_outputs(43) <= not(layer4_outputs(46)) or (layer4_outputs(138));
    layer5_outputs(44) <= not(layer4_outputs(2215));
    layer5_outputs(45) <= layer4_outputs(1213);
    layer5_outputs(46) <= not(layer4_outputs(1500));
    layer5_outputs(47) <= not(layer4_outputs(2409)) or (layer4_outputs(2502));
    layer5_outputs(48) <= layer4_outputs(1869);
    layer5_outputs(49) <= not(layer4_outputs(376));
    layer5_outputs(50) <= not(layer4_outputs(1371)) or (layer4_outputs(2527));
    layer5_outputs(51) <= layer4_outputs(116);
    layer5_outputs(52) <= not(layer4_outputs(65));
    layer5_outputs(53) <= not(layer4_outputs(2057));
    layer5_outputs(54) <= '0';
    layer5_outputs(55) <= not(layer4_outputs(648));
    layer5_outputs(56) <= layer4_outputs(1928);
    layer5_outputs(57) <= (layer4_outputs(776)) and not (layer4_outputs(1533));
    layer5_outputs(58) <= (layer4_outputs(225)) and not (layer4_outputs(1927));
    layer5_outputs(59) <= not(layer4_outputs(51));
    layer5_outputs(60) <= layer4_outputs(19);
    layer5_outputs(61) <= layer4_outputs(151);
    layer5_outputs(62) <= not(layer4_outputs(2234));
    layer5_outputs(63) <= not(layer4_outputs(1704));
    layer5_outputs(64) <= not(layer4_outputs(738));
    layer5_outputs(65) <= not(layer4_outputs(1480)) or (layer4_outputs(1231));
    layer5_outputs(66) <= (layer4_outputs(2370)) and (layer4_outputs(2093));
    layer5_outputs(67) <= not(layer4_outputs(1518));
    layer5_outputs(68) <= layer4_outputs(485);
    layer5_outputs(69) <= layer4_outputs(900);
    layer5_outputs(70) <= not((layer4_outputs(1458)) or (layer4_outputs(2357)));
    layer5_outputs(71) <= layer4_outputs(1671);
    layer5_outputs(72) <= (layer4_outputs(2004)) and not (layer4_outputs(2188));
    layer5_outputs(73) <= not(layer4_outputs(2189));
    layer5_outputs(74) <= not((layer4_outputs(1449)) xor (layer4_outputs(1135)));
    layer5_outputs(75) <= not((layer4_outputs(1609)) or (layer4_outputs(1755)));
    layer5_outputs(76) <= layer4_outputs(97);
    layer5_outputs(77) <= not(layer4_outputs(1436));
    layer5_outputs(78) <= not(layer4_outputs(1115));
    layer5_outputs(79) <= '1';
    layer5_outputs(80) <= (layer4_outputs(1713)) xor (layer4_outputs(979));
    layer5_outputs(81) <= layer4_outputs(836);
    layer5_outputs(82) <= not((layer4_outputs(1586)) xor (layer4_outputs(2342)));
    layer5_outputs(83) <= not(layer4_outputs(1498));
    layer5_outputs(84) <= not(layer4_outputs(1565));
    layer5_outputs(85) <= not(layer4_outputs(2292));
    layer5_outputs(86) <= layer4_outputs(2017);
    layer5_outputs(87) <= not((layer4_outputs(2228)) xor (layer4_outputs(1740)));
    layer5_outputs(88) <= not(layer4_outputs(649));
    layer5_outputs(89) <= not(layer4_outputs(212));
    layer5_outputs(90) <= layer4_outputs(282);
    layer5_outputs(91) <= not(layer4_outputs(1856));
    layer5_outputs(92) <= layer4_outputs(1284);
    layer5_outputs(93) <= layer4_outputs(150);
    layer5_outputs(94) <= not(layer4_outputs(424));
    layer5_outputs(95) <= not(layer4_outputs(1985)) or (layer4_outputs(2069));
    layer5_outputs(96) <= not(layer4_outputs(1462));
    layer5_outputs(97) <= layer4_outputs(1664);
    layer5_outputs(98) <= layer4_outputs(246);
    layer5_outputs(99) <= '1';
    layer5_outputs(100) <= not((layer4_outputs(1428)) or (layer4_outputs(488)));
    layer5_outputs(101) <= (layer4_outputs(118)) or (layer4_outputs(494));
    layer5_outputs(102) <= layer4_outputs(2075);
    layer5_outputs(103) <= layer4_outputs(2138);
    layer5_outputs(104) <= not(layer4_outputs(1375)) or (layer4_outputs(2012));
    layer5_outputs(105) <= not(layer4_outputs(1333));
    layer5_outputs(106) <= not((layer4_outputs(1025)) xor (layer4_outputs(2048)));
    layer5_outputs(107) <= not(layer4_outputs(80));
    layer5_outputs(108) <= (layer4_outputs(1784)) xor (layer4_outputs(11));
    layer5_outputs(109) <= layer4_outputs(575);
    layer5_outputs(110) <= not((layer4_outputs(1692)) or (layer4_outputs(1083)));
    layer5_outputs(111) <= (layer4_outputs(1276)) xor (layer4_outputs(735));
    layer5_outputs(112) <= not(layer4_outputs(1974)) or (layer4_outputs(398));
    layer5_outputs(113) <= not((layer4_outputs(2167)) and (layer4_outputs(1851)));
    layer5_outputs(114) <= (layer4_outputs(385)) xor (layer4_outputs(2150));
    layer5_outputs(115) <= (layer4_outputs(1136)) xor (layer4_outputs(2134));
    layer5_outputs(116) <= not(layer4_outputs(112));
    layer5_outputs(117) <= not(layer4_outputs(1996));
    layer5_outputs(118) <= not((layer4_outputs(1373)) xor (layer4_outputs(1247)));
    layer5_outputs(119) <= (layer4_outputs(1746)) or (layer4_outputs(1469));
    layer5_outputs(120) <= not(layer4_outputs(1359));
    layer5_outputs(121) <= not(layer4_outputs(97)) or (layer4_outputs(2002));
    layer5_outputs(122) <= (layer4_outputs(1185)) and (layer4_outputs(1958));
    layer5_outputs(123) <= not((layer4_outputs(814)) or (layer4_outputs(1183)));
    layer5_outputs(124) <= layer4_outputs(204);
    layer5_outputs(125) <= not(layer4_outputs(2165));
    layer5_outputs(126) <= (layer4_outputs(506)) and (layer4_outputs(545));
    layer5_outputs(127) <= '1';
    layer5_outputs(128) <= not((layer4_outputs(1971)) or (layer4_outputs(1503)));
    layer5_outputs(129) <= (layer4_outputs(818)) xor (layer4_outputs(256));
    layer5_outputs(130) <= (layer4_outputs(781)) and not (layer4_outputs(2460));
    layer5_outputs(131) <= (layer4_outputs(1223)) and (layer4_outputs(1217));
    layer5_outputs(132) <= not(layer4_outputs(778));
    layer5_outputs(133) <= (layer4_outputs(2124)) and (layer4_outputs(1291));
    layer5_outputs(134) <= layer4_outputs(1804);
    layer5_outputs(135) <= not(layer4_outputs(2123));
    layer5_outputs(136) <= not(layer4_outputs(2440));
    layer5_outputs(137) <= not((layer4_outputs(887)) xor (layer4_outputs(1474)));
    layer5_outputs(138) <= not(layer4_outputs(887));
    layer5_outputs(139) <= layer4_outputs(714);
    layer5_outputs(140) <= not(layer4_outputs(863));
    layer5_outputs(141) <= (layer4_outputs(347)) xor (layer4_outputs(1117));
    layer5_outputs(142) <= not((layer4_outputs(598)) and (layer4_outputs(199)));
    layer5_outputs(143) <= layer4_outputs(2511);
    layer5_outputs(144) <= not(layer4_outputs(23));
    layer5_outputs(145) <= layer4_outputs(1987);
    layer5_outputs(146) <= (layer4_outputs(729)) or (layer4_outputs(2541));
    layer5_outputs(147) <= layer4_outputs(1838);
    layer5_outputs(148) <= layer4_outputs(938);
    layer5_outputs(149) <= not(layer4_outputs(1478));
    layer5_outputs(150) <= layer4_outputs(1122);
    layer5_outputs(151) <= layer4_outputs(280);
    layer5_outputs(152) <= not((layer4_outputs(58)) or (layer4_outputs(1793)));
    layer5_outputs(153) <= (layer4_outputs(588)) and (layer4_outputs(1783));
    layer5_outputs(154) <= not(layer4_outputs(2133));
    layer5_outputs(155) <= not((layer4_outputs(1633)) and (layer4_outputs(1918)));
    layer5_outputs(156) <= not((layer4_outputs(693)) or (layer4_outputs(407)));
    layer5_outputs(157) <= not(layer4_outputs(1624));
    layer5_outputs(158) <= not(layer4_outputs(2497)) or (layer4_outputs(404));
    layer5_outputs(159) <= not(layer4_outputs(982));
    layer5_outputs(160) <= layer4_outputs(2032);
    layer5_outputs(161) <= not(layer4_outputs(1189)) or (layer4_outputs(1428));
    layer5_outputs(162) <= not(layer4_outputs(2401));
    layer5_outputs(163) <= not(layer4_outputs(2432));
    layer5_outputs(164) <= not(layer4_outputs(584)) or (layer4_outputs(2549));
    layer5_outputs(165) <= layer4_outputs(1723);
    layer5_outputs(166) <= not((layer4_outputs(696)) xor (layer4_outputs(1330)));
    layer5_outputs(167) <= not(layer4_outputs(1646));
    layer5_outputs(168) <= not(layer4_outputs(328));
    layer5_outputs(169) <= not((layer4_outputs(2014)) and (layer4_outputs(710)));
    layer5_outputs(170) <= '1';
    layer5_outputs(171) <= not(layer4_outputs(197)) or (layer4_outputs(879));
    layer5_outputs(172) <= layer4_outputs(1079);
    layer5_outputs(173) <= layer4_outputs(935);
    layer5_outputs(174) <= layer4_outputs(2149);
    layer5_outputs(175) <= (layer4_outputs(236)) and not (layer4_outputs(1099));
    layer5_outputs(176) <= not(layer4_outputs(1841));
    layer5_outputs(177) <= (layer4_outputs(477)) and (layer4_outputs(2243));
    layer5_outputs(178) <= (layer4_outputs(1525)) or (layer4_outputs(66));
    layer5_outputs(179) <= layer4_outputs(1741);
    layer5_outputs(180) <= layer4_outputs(928);
    layer5_outputs(181) <= not(layer4_outputs(583));
    layer5_outputs(182) <= (layer4_outputs(94)) and (layer4_outputs(1484));
    layer5_outputs(183) <= layer4_outputs(1309);
    layer5_outputs(184) <= layer4_outputs(1421);
    layer5_outputs(185) <= not(layer4_outputs(2308));
    layer5_outputs(186) <= '0';
    layer5_outputs(187) <= '0';
    layer5_outputs(188) <= (layer4_outputs(2166)) and not (layer4_outputs(638));
    layer5_outputs(189) <= (layer4_outputs(2038)) and (layer4_outputs(1691));
    layer5_outputs(190) <= layer4_outputs(168);
    layer5_outputs(191) <= not((layer4_outputs(1864)) or (layer4_outputs(349)));
    layer5_outputs(192) <= layer4_outputs(974);
    layer5_outputs(193) <= not(layer4_outputs(1753));
    layer5_outputs(194) <= layer4_outputs(938);
    layer5_outputs(195) <= layer4_outputs(424);
    layer5_outputs(196) <= not(layer4_outputs(2378));
    layer5_outputs(197) <= not((layer4_outputs(1286)) and (layer4_outputs(504)));
    layer5_outputs(198) <= layer4_outputs(1380);
    layer5_outputs(199) <= not(layer4_outputs(1951));
    layer5_outputs(200) <= not(layer4_outputs(1084)) or (layer4_outputs(247));
    layer5_outputs(201) <= (layer4_outputs(1252)) and not (layer4_outputs(2452));
    layer5_outputs(202) <= (layer4_outputs(1726)) and (layer4_outputs(2266));
    layer5_outputs(203) <= not((layer4_outputs(2240)) xor (layer4_outputs(883)));
    layer5_outputs(204) <= layer4_outputs(209);
    layer5_outputs(205) <= not(layer4_outputs(2019));
    layer5_outputs(206) <= not((layer4_outputs(2539)) or (layer4_outputs(2287)));
    layer5_outputs(207) <= not((layer4_outputs(2066)) xor (layer4_outputs(1962)));
    layer5_outputs(208) <= not(layer4_outputs(314)) or (layer4_outputs(1479));
    layer5_outputs(209) <= (layer4_outputs(710)) or (layer4_outputs(1686));
    layer5_outputs(210) <= (layer4_outputs(213)) and not (layer4_outputs(1960));
    layer5_outputs(211) <= (layer4_outputs(2297)) and not (layer4_outputs(0));
    layer5_outputs(212) <= not(layer4_outputs(593)) or (layer4_outputs(102));
    layer5_outputs(213) <= not(layer4_outputs(22));
    layer5_outputs(214) <= layer4_outputs(1836);
    layer5_outputs(215) <= layer4_outputs(966);
    layer5_outputs(216) <= not(layer4_outputs(1762));
    layer5_outputs(217) <= '1';
    layer5_outputs(218) <= not(layer4_outputs(1824)) or (layer4_outputs(1459));
    layer5_outputs(219) <= '0';
    layer5_outputs(220) <= layer4_outputs(904);
    layer5_outputs(221) <= not((layer4_outputs(1514)) and (layer4_outputs(773)));
    layer5_outputs(222) <= not(layer4_outputs(1212));
    layer5_outputs(223) <= not(layer4_outputs(701));
    layer5_outputs(224) <= (layer4_outputs(2054)) or (layer4_outputs(1889));
    layer5_outputs(225) <= (layer4_outputs(1847)) and not (layer4_outputs(1173));
    layer5_outputs(226) <= not((layer4_outputs(2109)) xor (layer4_outputs(1325)));
    layer5_outputs(227) <= not(layer4_outputs(339));
    layer5_outputs(228) <= not((layer4_outputs(2091)) and (layer4_outputs(2188)));
    layer5_outputs(229) <= (layer4_outputs(1226)) xor (layer4_outputs(2184));
    layer5_outputs(230) <= layer4_outputs(666);
    layer5_outputs(231) <= not(layer4_outputs(2207));
    layer5_outputs(232) <= not(layer4_outputs(1186)) or (layer4_outputs(319));
    layer5_outputs(233) <= layer4_outputs(1750);
    layer5_outputs(234) <= (layer4_outputs(464)) and not (layer4_outputs(2178));
    layer5_outputs(235) <= layer4_outputs(2006);
    layer5_outputs(236) <= (layer4_outputs(826)) xor (layer4_outputs(91));
    layer5_outputs(237) <= (layer4_outputs(1645)) and (layer4_outputs(2037));
    layer5_outputs(238) <= (layer4_outputs(169)) xor (layer4_outputs(628));
    layer5_outputs(239) <= not(layer4_outputs(1734));
    layer5_outputs(240) <= not((layer4_outputs(2473)) xor (layer4_outputs(2232)));
    layer5_outputs(241) <= not(layer4_outputs(1465)) or (layer4_outputs(1623));
    layer5_outputs(242) <= not(layer4_outputs(648));
    layer5_outputs(243) <= not(layer4_outputs(1164));
    layer5_outputs(244) <= layer4_outputs(304);
    layer5_outputs(245) <= not(layer4_outputs(841));
    layer5_outputs(246) <= layer4_outputs(984);
    layer5_outputs(247) <= not((layer4_outputs(1952)) xor (layer4_outputs(419)));
    layer5_outputs(248) <= '1';
    layer5_outputs(249) <= layer4_outputs(1628);
    layer5_outputs(250) <= (layer4_outputs(98)) and not (layer4_outputs(519));
    layer5_outputs(251) <= layer4_outputs(250);
    layer5_outputs(252) <= not(layer4_outputs(1601));
    layer5_outputs(253) <= layer4_outputs(2483);
    layer5_outputs(254) <= layer4_outputs(1244);
    layer5_outputs(255) <= not((layer4_outputs(1343)) or (layer4_outputs(1382)));
    layer5_outputs(256) <= '0';
    layer5_outputs(257) <= not(layer4_outputs(2399));
    layer5_outputs(258) <= not(layer4_outputs(811)) or (layer4_outputs(631));
    layer5_outputs(259) <= not(layer4_outputs(2507));
    layer5_outputs(260) <= not((layer4_outputs(1656)) and (layer4_outputs(1467)));
    layer5_outputs(261) <= layer4_outputs(1578);
    layer5_outputs(262) <= layer4_outputs(2256);
    layer5_outputs(263) <= '1';
    layer5_outputs(264) <= not(layer4_outputs(508)) or (layer4_outputs(890));
    layer5_outputs(265) <= (layer4_outputs(745)) and not (layer4_outputs(1771));
    layer5_outputs(266) <= layer4_outputs(1053);
    layer5_outputs(267) <= (layer4_outputs(844)) or (layer4_outputs(2277));
    layer5_outputs(268) <= not(layer4_outputs(1786));
    layer5_outputs(269) <= layer4_outputs(1417);
    layer5_outputs(270) <= (layer4_outputs(1086)) and not (layer4_outputs(2177));
    layer5_outputs(271) <= (layer4_outputs(1707)) or (layer4_outputs(263));
    layer5_outputs(272) <= not(layer4_outputs(1614)) or (layer4_outputs(1964));
    layer5_outputs(273) <= not(layer4_outputs(318)) or (layer4_outputs(2235));
    layer5_outputs(274) <= layer4_outputs(2284);
    layer5_outputs(275) <= not((layer4_outputs(1393)) or (layer4_outputs(2019)));
    layer5_outputs(276) <= layer4_outputs(1074);
    layer5_outputs(277) <= not((layer4_outputs(530)) and (layer4_outputs(2543)));
    layer5_outputs(278) <= (layer4_outputs(1364)) and not (layer4_outputs(484));
    layer5_outputs(279) <= not((layer4_outputs(1225)) xor (layer4_outputs(926)));
    layer5_outputs(280) <= not(layer4_outputs(2223));
    layer5_outputs(281) <= not(layer4_outputs(1978)) or (layer4_outputs(1233));
    layer5_outputs(282) <= layer4_outputs(1258);
    layer5_outputs(283) <= layer4_outputs(1322);
    layer5_outputs(284) <= (layer4_outputs(550)) and not (layer4_outputs(365));
    layer5_outputs(285) <= (layer4_outputs(753)) and not (layer4_outputs(1363));
    layer5_outputs(286) <= not(layer4_outputs(1050)) or (layer4_outputs(1953));
    layer5_outputs(287) <= not(layer4_outputs(1761)) or (layer4_outputs(1420));
    layer5_outputs(288) <= (layer4_outputs(2495)) xor (layer4_outputs(1118));
    layer5_outputs(289) <= not((layer4_outputs(2398)) or (layer4_outputs(1810)));
    layer5_outputs(290) <= not((layer4_outputs(2498)) and (layer4_outputs(1063)));
    layer5_outputs(291) <= not(layer4_outputs(1979));
    layer5_outputs(292) <= (layer4_outputs(1659)) and not (layer4_outputs(2544));
    layer5_outputs(293) <= not(layer4_outputs(1298));
    layer5_outputs(294) <= layer4_outputs(633);
    layer5_outputs(295) <= (layer4_outputs(106)) and (layer4_outputs(766));
    layer5_outputs(296) <= layer4_outputs(895);
    layer5_outputs(297) <= not((layer4_outputs(1708)) and (layer4_outputs(15)));
    layer5_outputs(298) <= layer4_outputs(1871);
    layer5_outputs(299) <= (layer4_outputs(903)) xor (layer4_outputs(1510));
    layer5_outputs(300) <= not(layer4_outputs(412));
    layer5_outputs(301) <= not((layer4_outputs(2151)) and (layer4_outputs(2153)));
    layer5_outputs(302) <= not(layer4_outputs(127));
    layer5_outputs(303) <= (layer4_outputs(2)) and not (layer4_outputs(1738));
    layer5_outputs(304) <= layer4_outputs(2083);
    layer5_outputs(305) <= not(layer4_outputs(298)) or (layer4_outputs(646));
    layer5_outputs(306) <= layer4_outputs(1646);
    layer5_outputs(307) <= (layer4_outputs(1408)) or (layer4_outputs(2115));
    layer5_outputs(308) <= not((layer4_outputs(2013)) xor (layer4_outputs(366)));
    layer5_outputs(309) <= not((layer4_outputs(1015)) xor (layer4_outputs(691)));
    layer5_outputs(310) <= (layer4_outputs(2506)) and not (layer4_outputs(1741));
    layer5_outputs(311) <= layer4_outputs(1698);
    layer5_outputs(312) <= '1';
    layer5_outputs(313) <= not((layer4_outputs(262)) and (layer4_outputs(616)));
    layer5_outputs(314) <= layer4_outputs(639);
    layer5_outputs(315) <= not(layer4_outputs(2558));
    layer5_outputs(316) <= not(layer4_outputs(1727));
    layer5_outputs(317) <= not(layer4_outputs(2133)) or (layer4_outputs(1193));
    layer5_outputs(318) <= layer4_outputs(1640);
    layer5_outputs(319) <= (layer4_outputs(2463)) and not (layer4_outputs(1620));
    layer5_outputs(320) <= not((layer4_outputs(57)) or (layer4_outputs(1849)));
    layer5_outputs(321) <= (layer4_outputs(228)) xor (layer4_outputs(2002));
    layer5_outputs(322) <= (layer4_outputs(1720)) and not (layer4_outputs(1966));
    layer5_outputs(323) <= not((layer4_outputs(531)) xor (layer4_outputs(2031)));
    layer5_outputs(324) <= not(layer4_outputs(1002));
    layer5_outputs(325) <= (layer4_outputs(1140)) xor (layer4_outputs(2015));
    layer5_outputs(326) <= layer4_outputs(1996);
    layer5_outputs(327) <= layer4_outputs(658);
    layer5_outputs(328) <= not(layer4_outputs(1852)) or (layer4_outputs(1262));
    layer5_outputs(329) <= not(layer4_outputs(1833));
    layer5_outputs(330) <= (layer4_outputs(1785)) and not (layer4_outputs(1003));
    layer5_outputs(331) <= (layer4_outputs(1983)) xor (layer4_outputs(796));
    layer5_outputs(332) <= (layer4_outputs(1024)) and not (layer4_outputs(808));
    layer5_outputs(333) <= not(layer4_outputs(2154));
    layer5_outputs(334) <= not(layer4_outputs(1184));
    layer5_outputs(335) <= not(layer4_outputs(784));
    layer5_outputs(336) <= not(layer4_outputs(1192));
    layer5_outputs(337) <= not(layer4_outputs(908));
    layer5_outputs(338) <= (layer4_outputs(2373)) and (layer4_outputs(580));
    layer5_outputs(339) <= not(layer4_outputs(2283));
    layer5_outputs(340) <= not(layer4_outputs(2303));
    layer5_outputs(341) <= layer4_outputs(1670);
    layer5_outputs(342) <= not(layer4_outputs(1809)) or (layer4_outputs(558));
    layer5_outputs(343) <= layer4_outputs(1188);
    layer5_outputs(344) <= (layer4_outputs(2415)) or (layer4_outputs(605));
    layer5_outputs(345) <= not(layer4_outputs(1721)) or (layer4_outputs(1611));
    layer5_outputs(346) <= '0';
    layer5_outputs(347) <= not(layer4_outputs(1407));
    layer5_outputs(348) <= (layer4_outputs(1412)) or (layer4_outputs(1691));
    layer5_outputs(349) <= '0';
    layer5_outputs(350) <= not(layer4_outputs(1220)) or (layer4_outputs(1626));
    layer5_outputs(351) <= '0';
    layer5_outputs(352) <= not(layer4_outputs(840));
    layer5_outputs(353) <= (layer4_outputs(2443)) and not (layer4_outputs(1757));
    layer5_outputs(354) <= (layer4_outputs(1029)) and not (layer4_outputs(2179));
    layer5_outputs(355) <= layer4_outputs(1218);
    layer5_outputs(356) <= layer4_outputs(2076);
    layer5_outputs(357) <= layer4_outputs(672);
    layer5_outputs(358) <= not(layer4_outputs(2386));
    layer5_outputs(359) <= not((layer4_outputs(2517)) xor (layer4_outputs(1687)));
    layer5_outputs(360) <= layer4_outputs(1442);
    layer5_outputs(361) <= not(layer4_outputs(504));
    layer5_outputs(362) <= layer4_outputs(1912);
    layer5_outputs(363) <= not(layer4_outputs(394));
    layer5_outputs(364) <= '0';
    layer5_outputs(365) <= (layer4_outputs(1112)) and not (layer4_outputs(1467));
    layer5_outputs(366) <= layer4_outputs(2168);
    layer5_outputs(367) <= not(layer4_outputs(48));
    layer5_outputs(368) <= not((layer4_outputs(577)) and (layer4_outputs(1032)));
    layer5_outputs(369) <= layer4_outputs(1282);
    layer5_outputs(370) <= (layer4_outputs(236)) xor (layer4_outputs(2099));
    layer5_outputs(371) <= layer4_outputs(252);
    layer5_outputs(372) <= layer4_outputs(319);
    layer5_outputs(373) <= not(layer4_outputs(1145));
    layer5_outputs(374) <= '1';
    layer5_outputs(375) <= layer4_outputs(2127);
    layer5_outputs(376) <= not((layer4_outputs(324)) and (layer4_outputs(2095)));
    layer5_outputs(377) <= layer4_outputs(499);
    layer5_outputs(378) <= (layer4_outputs(2341)) and not (layer4_outputs(882));
    layer5_outputs(379) <= not(layer4_outputs(3));
    layer5_outputs(380) <= (layer4_outputs(1710)) xor (layer4_outputs(2367));
    layer5_outputs(381) <= (layer4_outputs(136)) and not (layer4_outputs(2493));
    layer5_outputs(382) <= (layer4_outputs(1440)) and not (layer4_outputs(2152));
    layer5_outputs(383) <= not((layer4_outputs(670)) xor (layer4_outputs(852)));
    layer5_outputs(384) <= not((layer4_outputs(930)) xor (layer4_outputs(458)));
    layer5_outputs(385) <= layer4_outputs(1302);
    layer5_outputs(386) <= layer4_outputs(369);
    layer5_outputs(387) <= (layer4_outputs(729)) or (layer4_outputs(1600));
    layer5_outputs(388) <= not(layer4_outputs(456)) or (layer4_outputs(2540));
    layer5_outputs(389) <= not(layer4_outputs(2029));
    layer5_outputs(390) <= (layer4_outputs(645)) and not (layer4_outputs(611));
    layer5_outputs(391) <= (layer4_outputs(1006)) and (layer4_outputs(792));
    layer5_outputs(392) <= not(layer4_outputs(1234));
    layer5_outputs(393) <= (layer4_outputs(483)) and (layer4_outputs(12));
    layer5_outputs(394) <= not(layer4_outputs(1998));
    layer5_outputs(395) <= not((layer4_outputs(75)) and (layer4_outputs(2144)));
    layer5_outputs(396) <= (layer4_outputs(91)) and not (layer4_outputs(2146));
    layer5_outputs(397) <= not(layer4_outputs(432)) or (layer4_outputs(302));
    layer5_outputs(398) <= layer4_outputs(168);
    layer5_outputs(399) <= not(layer4_outputs(786));
    layer5_outputs(400) <= not((layer4_outputs(193)) xor (layer4_outputs(662)));
    layer5_outputs(401) <= not(layer4_outputs(937));
    layer5_outputs(402) <= not(layer4_outputs(2116));
    layer5_outputs(403) <= not(layer4_outputs(1516));
    layer5_outputs(404) <= layer4_outputs(2020);
    layer5_outputs(405) <= (layer4_outputs(1386)) and not (layer4_outputs(2257));
    layer5_outputs(406) <= not((layer4_outputs(1668)) and (layer4_outputs(1026)));
    layer5_outputs(407) <= layer4_outputs(1524);
    layer5_outputs(408) <= layer4_outputs(2385);
    layer5_outputs(409) <= not(layer4_outputs(351));
    layer5_outputs(410) <= (layer4_outputs(1)) and not (layer4_outputs(1293));
    layer5_outputs(411) <= layer4_outputs(325);
    layer5_outputs(412) <= layer4_outputs(572);
    layer5_outputs(413) <= not((layer4_outputs(578)) and (layer4_outputs(2170)));
    layer5_outputs(414) <= (layer4_outputs(2363)) or (layer4_outputs(1051));
    layer5_outputs(415) <= not((layer4_outputs(1010)) xor (layer4_outputs(382)));
    layer5_outputs(416) <= not((layer4_outputs(665)) xor (layer4_outputs(1902)));
    layer5_outputs(417) <= layer4_outputs(998);
    layer5_outputs(418) <= layer4_outputs(1490);
    layer5_outputs(419) <= layer4_outputs(755);
    layer5_outputs(420) <= not(layer4_outputs(1630));
    layer5_outputs(421) <= layer4_outputs(521);
    layer5_outputs(422) <= (layer4_outputs(1883)) and not (layer4_outputs(2092));
    layer5_outputs(423) <= (layer4_outputs(378)) and not (layer4_outputs(1149));
    layer5_outputs(424) <= layer4_outputs(2244);
    layer5_outputs(425) <= not(layer4_outputs(145));
    layer5_outputs(426) <= not(layer4_outputs(1676));
    layer5_outputs(427) <= layer4_outputs(1589);
    layer5_outputs(428) <= '1';
    layer5_outputs(429) <= (layer4_outputs(737)) and not (layer4_outputs(1794));
    layer5_outputs(430) <= (layer4_outputs(743)) or (layer4_outputs(2024));
    layer5_outputs(431) <= not(layer4_outputs(1926));
    layer5_outputs(432) <= not((layer4_outputs(60)) or (layer4_outputs(2408)));
    layer5_outputs(433) <= layer4_outputs(2376);
    layer5_outputs(434) <= (layer4_outputs(1172)) xor (layer4_outputs(942));
    layer5_outputs(435) <= '0';
    layer5_outputs(436) <= (layer4_outputs(2103)) xor (layer4_outputs(131));
    layer5_outputs(437) <= not(layer4_outputs(204));
    layer5_outputs(438) <= (layer4_outputs(410)) and not (layer4_outputs(182));
    layer5_outputs(439) <= (layer4_outputs(1209)) xor (layer4_outputs(1503));
    layer5_outputs(440) <= (layer4_outputs(2007)) and not (layer4_outputs(1712));
    layer5_outputs(441) <= layer4_outputs(2298);
    layer5_outputs(442) <= layer4_outputs(647);
    layer5_outputs(443) <= not(layer4_outputs(1546));
    layer5_outputs(444) <= not((layer4_outputs(697)) or (layer4_outputs(1324)));
    layer5_outputs(445) <= (layer4_outputs(1203)) xor (layer4_outputs(706));
    layer5_outputs(446) <= not(layer4_outputs(624));
    layer5_outputs(447) <= not((layer4_outputs(395)) xor (layer4_outputs(746)));
    layer5_outputs(448) <= (layer4_outputs(345)) or (layer4_outputs(646));
    layer5_outputs(449) <= not((layer4_outputs(1413)) and (layer4_outputs(0)));
    layer5_outputs(450) <= not(layer4_outputs(1045)) or (layer4_outputs(351));
    layer5_outputs(451) <= '1';
    layer5_outputs(452) <= not(layer4_outputs(1867));
    layer5_outputs(453) <= '0';
    layer5_outputs(454) <= not((layer4_outputs(1731)) xor (layer4_outputs(361)));
    layer5_outputs(455) <= layer4_outputs(2089);
    layer5_outputs(456) <= not(layer4_outputs(2005));
    layer5_outputs(457) <= not((layer4_outputs(943)) and (layer4_outputs(1148)));
    layer5_outputs(458) <= layer4_outputs(2462);
    layer5_outputs(459) <= layer4_outputs(1742);
    layer5_outputs(460) <= (layer4_outputs(2294)) or (layer4_outputs(1199));
    layer5_outputs(461) <= layer4_outputs(1125);
    layer5_outputs(462) <= not(layer4_outputs(526));
    layer5_outputs(463) <= '1';
    layer5_outputs(464) <= (layer4_outputs(1639)) and not (layer4_outputs(1446));
    layer5_outputs(465) <= (layer4_outputs(907)) xor (layer4_outputs(411));
    layer5_outputs(466) <= not((layer4_outputs(1181)) and (layer4_outputs(1310)));
    layer5_outputs(467) <= not(layer4_outputs(426));
    layer5_outputs(468) <= not(layer4_outputs(925));
    layer5_outputs(469) <= layer4_outputs(615);
    layer5_outputs(470) <= (layer4_outputs(2286)) and not (layer4_outputs(1165));
    layer5_outputs(471) <= not((layer4_outputs(1230)) or (layer4_outputs(1222)));
    layer5_outputs(472) <= layer4_outputs(1424);
    layer5_outputs(473) <= layer4_outputs(197);
    layer5_outputs(474) <= layer4_outputs(857);
    layer5_outputs(475) <= not(layer4_outputs(741));
    layer5_outputs(476) <= layer4_outputs(2132);
    layer5_outputs(477) <= (layer4_outputs(1526)) and not (layer4_outputs(809));
    layer5_outputs(478) <= (layer4_outputs(148)) and not (layer4_outputs(1925));
    layer5_outputs(479) <= (layer4_outputs(2524)) and (layer4_outputs(2246));
    layer5_outputs(480) <= (layer4_outputs(2534)) and (layer4_outputs(466));
    layer5_outputs(481) <= not(layer4_outputs(2219));
    layer5_outputs(482) <= not(layer4_outputs(1724));
    layer5_outputs(483) <= (layer4_outputs(761)) and not (layer4_outputs(2403));
    layer5_outputs(484) <= (layer4_outputs(238)) and not (layer4_outputs(876));
    layer5_outputs(485) <= not((layer4_outputs(54)) xor (layer4_outputs(2243)));
    layer5_outputs(486) <= not(layer4_outputs(754)) or (layer4_outputs(1178));
    layer5_outputs(487) <= '0';
    layer5_outputs(488) <= '1';
    layer5_outputs(489) <= '1';
    layer5_outputs(490) <= not(layer4_outputs(1537));
    layer5_outputs(491) <= layer4_outputs(1893);
    layer5_outputs(492) <= '1';
    layer5_outputs(493) <= not(layer4_outputs(1676));
    layer5_outputs(494) <= not(layer4_outputs(2394));
    layer5_outputs(495) <= layer4_outputs(520);
    layer5_outputs(496) <= layer4_outputs(744);
    layer5_outputs(497) <= layer4_outputs(1345);
    layer5_outputs(498) <= layer4_outputs(792);
    layer5_outputs(499) <= layer4_outputs(1744);
    layer5_outputs(500) <= '0';
    layer5_outputs(501) <= (layer4_outputs(1567)) and not (layer4_outputs(416));
    layer5_outputs(502) <= layer4_outputs(167);
    layer5_outputs(503) <= not((layer4_outputs(1399)) or (layer4_outputs(136)));
    layer5_outputs(504) <= layer4_outputs(702);
    layer5_outputs(505) <= '1';
    layer5_outputs(506) <= layer4_outputs(1406);
    layer5_outputs(507) <= (layer4_outputs(2471)) and (layer4_outputs(1812));
    layer5_outputs(508) <= not((layer4_outputs(285)) or (layer4_outputs(1688)));
    layer5_outputs(509) <= not(layer4_outputs(2485)) or (layer4_outputs(2021));
    layer5_outputs(510) <= not(layer4_outputs(834)) or (layer4_outputs(2316));
    layer5_outputs(511) <= (layer4_outputs(440)) or (layer4_outputs(1133));
    layer5_outputs(512) <= layer4_outputs(2553);
    layer5_outputs(513) <= not(layer4_outputs(1684)) or (layer4_outputs(1486));
    layer5_outputs(514) <= not(layer4_outputs(766));
    layer5_outputs(515) <= not(layer4_outputs(2041));
    layer5_outputs(516) <= layer4_outputs(705);
    layer5_outputs(517) <= not(layer4_outputs(549)) or (layer4_outputs(1204));
    layer5_outputs(518) <= not(layer4_outputs(1209));
    layer5_outputs(519) <= not(layer4_outputs(88)) or (layer4_outputs(13));
    layer5_outputs(520) <= not(layer4_outputs(159));
    layer5_outputs(521) <= not(layer4_outputs(1732));
    layer5_outputs(522) <= layer4_outputs(849);
    layer5_outputs(523) <= not(layer4_outputs(318));
    layer5_outputs(524) <= not(layer4_outputs(2001)) or (layer4_outputs(1594));
    layer5_outputs(525) <= (layer4_outputs(1511)) xor (layer4_outputs(367));
    layer5_outputs(526) <= layer4_outputs(503);
    layer5_outputs(527) <= not((layer4_outputs(985)) or (layer4_outputs(366)));
    layer5_outputs(528) <= not(layer4_outputs(249));
    layer5_outputs(529) <= '1';
    layer5_outputs(530) <= not(layer4_outputs(1186));
    layer5_outputs(531) <= (layer4_outputs(2380)) or (layer4_outputs(1541));
    layer5_outputs(532) <= not(layer4_outputs(524));
    layer5_outputs(533) <= layer4_outputs(528);
    layer5_outputs(534) <= (layer4_outputs(345)) and not (layer4_outputs(2355));
    layer5_outputs(535) <= (layer4_outputs(475)) or (layer4_outputs(727));
    layer5_outputs(536) <= (layer4_outputs(2512)) and not (layer4_outputs(2156));
    layer5_outputs(537) <= (layer4_outputs(2552)) and not (layer4_outputs(2357));
    layer5_outputs(538) <= layer4_outputs(579);
    layer5_outputs(539) <= layer4_outputs(2284);
    layer5_outputs(540) <= layer4_outputs(1625);
    layer5_outputs(541) <= not(layer4_outputs(1217));
    layer5_outputs(542) <= '0';
    layer5_outputs(543) <= not(layer4_outputs(1806)) or (layer4_outputs(2447));
    layer5_outputs(544) <= not((layer4_outputs(2070)) or (layer4_outputs(612)));
    layer5_outputs(545) <= not((layer4_outputs(1821)) or (layer4_outputs(1666)));
    layer5_outputs(546) <= not(layer4_outputs(1078));
    layer5_outputs(547) <= not(layer4_outputs(2280));
    layer5_outputs(548) <= not(layer4_outputs(1453)) or (layer4_outputs(2307));
    layer5_outputs(549) <= not(layer4_outputs(331));
    layer5_outputs(550) <= not(layer4_outputs(2271));
    layer5_outputs(551) <= not((layer4_outputs(429)) and (layer4_outputs(683)));
    layer5_outputs(552) <= layer4_outputs(1492);
    layer5_outputs(553) <= (layer4_outputs(1038)) or (layer4_outputs(1531));
    layer5_outputs(554) <= (layer4_outputs(184)) and (layer4_outputs(1727));
    layer5_outputs(555) <= not((layer4_outputs(417)) xor (layer4_outputs(89)));
    layer5_outputs(556) <= (layer4_outputs(1509)) xor (layer4_outputs(1040));
    layer5_outputs(557) <= (layer4_outputs(1670)) and (layer4_outputs(1288));
    layer5_outputs(558) <= layer4_outputs(2548);
    layer5_outputs(559) <= '0';
    layer5_outputs(560) <= not(layer4_outputs(1574)) or (layer4_outputs(2328));
    layer5_outputs(561) <= layer4_outputs(1166);
    layer5_outputs(562) <= (layer4_outputs(1965)) and (layer4_outputs(1842));
    layer5_outputs(563) <= not(layer4_outputs(749)) or (layer4_outputs(325));
    layer5_outputs(564) <= not(layer4_outputs(1860)) or (layer4_outputs(203));
    layer5_outputs(565) <= layer4_outputs(1212);
    layer5_outputs(566) <= (layer4_outputs(1398)) and (layer4_outputs(259));
    layer5_outputs(567) <= layer4_outputs(2209);
    layer5_outputs(568) <= (layer4_outputs(859)) xor (layer4_outputs(860));
    layer5_outputs(569) <= not(layer4_outputs(83)) or (layer4_outputs(393));
    layer5_outputs(570) <= (layer4_outputs(1657)) xor (layer4_outputs(2343));
    layer5_outputs(571) <= layer4_outputs(558);
    layer5_outputs(572) <= (layer4_outputs(286)) xor (layer4_outputs(1450));
    layer5_outputs(573) <= not((layer4_outputs(2454)) or (layer4_outputs(186)));
    layer5_outputs(574) <= not((layer4_outputs(1390)) xor (layer4_outputs(894)));
    layer5_outputs(575) <= '1';
    layer5_outputs(576) <= not(layer4_outputs(724)) or (layer4_outputs(1021));
    layer5_outputs(577) <= (layer4_outputs(682)) xor (layer4_outputs(2214));
    layer5_outputs(578) <= not(layer4_outputs(616));
    layer5_outputs(579) <= not((layer4_outputs(703)) xor (layer4_outputs(2352)));
    layer5_outputs(580) <= not(layer4_outputs(2238));
    layer5_outputs(581) <= not(layer4_outputs(1476)) or (layer4_outputs(686));
    layer5_outputs(582) <= not(layer4_outputs(1411));
    layer5_outputs(583) <= (layer4_outputs(869)) and (layer4_outputs(1968));
    layer5_outputs(584) <= not(layer4_outputs(2277)) or (layer4_outputs(2535));
    layer5_outputs(585) <= (layer4_outputs(853)) and not (layer4_outputs(2175));
    layer5_outputs(586) <= not(layer4_outputs(2456));
    layer5_outputs(587) <= (layer4_outputs(948)) and not (layer4_outputs(1073));
    layer5_outputs(588) <= not(layer4_outputs(1941)) or (layer4_outputs(2524));
    layer5_outputs(589) <= not(layer4_outputs(1466));
    layer5_outputs(590) <= not(layer4_outputs(1463)) or (layer4_outputs(431));
    layer5_outputs(591) <= not(layer4_outputs(2420));
    layer5_outputs(592) <= layer4_outputs(2142);
    layer5_outputs(593) <= (layer4_outputs(1572)) and (layer4_outputs(2359));
    layer5_outputs(594) <= layer4_outputs(1350);
    layer5_outputs(595) <= layer4_outputs(1095);
    layer5_outputs(596) <= not(layer4_outputs(791));
    layer5_outputs(597) <= (layer4_outputs(57)) and not (layer4_outputs(1158));
    layer5_outputs(598) <= not(layer4_outputs(761)) or (layer4_outputs(2289));
    layer5_outputs(599) <= (layer4_outputs(531)) and not (layer4_outputs(870));
    layer5_outputs(600) <= '1';
    layer5_outputs(601) <= '1';
    layer5_outputs(602) <= not(layer4_outputs(898));
    layer5_outputs(603) <= not(layer4_outputs(953));
    layer5_outputs(604) <= layer4_outputs(2185);
    layer5_outputs(605) <= (layer4_outputs(119)) and not (layer4_outputs(1069));
    layer5_outputs(606) <= (layer4_outputs(1667)) and not (layer4_outputs(587));
    layer5_outputs(607) <= layer4_outputs(1280);
    layer5_outputs(608) <= not((layer4_outputs(569)) or (layer4_outputs(1736)));
    layer5_outputs(609) <= layer4_outputs(1702);
    layer5_outputs(610) <= layer4_outputs(1037);
    layer5_outputs(611) <= (layer4_outputs(1812)) and not (layer4_outputs(599));
    layer5_outputs(612) <= layer4_outputs(2155);
    layer5_outputs(613) <= (layer4_outputs(2218)) and not (layer4_outputs(1227));
    layer5_outputs(614) <= layer4_outputs(1273);
    layer5_outputs(615) <= not(layer4_outputs(1677));
    layer5_outputs(616) <= '1';
    layer5_outputs(617) <= layer4_outputs(2455);
    layer5_outputs(618) <= not(layer4_outputs(1284));
    layer5_outputs(619) <= not(layer4_outputs(237)) or (layer4_outputs(2258));
    layer5_outputs(620) <= layer4_outputs(41);
    layer5_outputs(621) <= layer4_outputs(1469);
    layer5_outputs(622) <= (layer4_outputs(437)) and not (layer4_outputs(2491));
    layer5_outputs(623) <= '1';
    layer5_outputs(624) <= not(layer4_outputs(133)) or (layer4_outputs(1405));
    layer5_outputs(625) <= (layer4_outputs(722)) or (layer4_outputs(1269));
    layer5_outputs(626) <= layer4_outputs(1220);
    layer5_outputs(627) <= not(layer4_outputs(1599));
    layer5_outputs(628) <= not(layer4_outputs(1489));
    layer5_outputs(629) <= layer4_outputs(219);
    layer5_outputs(630) <= not(layer4_outputs(975)) or (layer4_outputs(321));
    layer5_outputs(631) <= (layer4_outputs(2241)) or (layer4_outputs(2131));
    layer5_outputs(632) <= not((layer4_outputs(1086)) and (layer4_outputs(1047)));
    layer5_outputs(633) <= (layer4_outputs(1888)) or (layer4_outputs(1697));
    layer5_outputs(634) <= not((layer4_outputs(42)) and (layer4_outputs(906)));
    layer5_outputs(635) <= layer4_outputs(1539);
    layer5_outputs(636) <= not((layer4_outputs(461)) xor (layer4_outputs(2397)));
    layer5_outputs(637) <= not(layer4_outputs(1886));
    layer5_outputs(638) <= not(layer4_outputs(1436)) or (layer4_outputs(377));
    layer5_outputs(639) <= (layer4_outputs(1791)) or (layer4_outputs(390));
    layer5_outputs(640) <= (layer4_outputs(2242)) and not (layer4_outputs(570));
    layer5_outputs(641) <= layer4_outputs(2450);
    layer5_outputs(642) <= not((layer4_outputs(821)) and (layer4_outputs(1847)));
    layer5_outputs(643) <= layer4_outputs(162);
    layer5_outputs(644) <= (layer4_outputs(2466)) or (layer4_outputs(543));
    layer5_outputs(645) <= '0';
    layer5_outputs(646) <= not((layer4_outputs(1225)) and (layer4_outputs(1649)));
    layer5_outputs(647) <= not(layer4_outputs(1764));
    layer5_outputs(648) <= layer4_outputs(2283);
    layer5_outputs(649) <= (layer4_outputs(2530)) and not (layer4_outputs(2474));
    layer5_outputs(650) <= not(layer4_outputs(375));
    layer5_outputs(651) <= (layer4_outputs(69)) and not (layer4_outputs(650));
    layer5_outputs(652) <= layer4_outputs(1512);
    layer5_outputs(653) <= (layer4_outputs(352)) or (layer4_outputs(886));
    layer5_outputs(654) <= (layer4_outputs(1585)) and (layer4_outputs(1513));
    layer5_outputs(655) <= not(layer4_outputs(2237)) or (layer4_outputs(1714));
    layer5_outputs(656) <= '1';
    layer5_outputs(657) <= layer4_outputs(955);
    layer5_outputs(658) <= (layer4_outputs(1750)) and not (layer4_outputs(959));
    layer5_outputs(659) <= not((layer4_outputs(746)) and (layer4_outputs(1392)));
    layer5_outputs(660) <= not((layer4_outputs(338)) and (layer4_outputs(1700)));
    layer5_outputs(661) <= (layer4_outputs(265)) and (layer4_outputs(713));
    layer5_outputs(662) <= (layer4_outputs(2259)) and not (layer4_outputs(1692));
    layer5_outputs(663) <= layer4_outputs(292);
    layer5_outputs(664) <= (layer4_outputs(628)) or (layer4_outputs(2480));
    layer5_outputs(665) <= layer4_outputs(1897);
    layer5_outputs(666) <= (layer4_outputs(663)) and not (layer4_outputs(881));
    layer5_outputs(667) <= not((layer4_outputs(2384)) and (layer4_outputs(496)));
    layer5_outputs(668) <= (layer4_outputs(15)) xor (layer4_outputs(690));
    layer5_outputs(669) <= (layer4_outputs(2098)) and not (layer4_outputs(951));
    layer5_outputs(670) <= layer4_outputs(267);
    layer5_outputs(671) <= (layer4_outputs(1829)) and not (layer4_outputs(2323));
    layer5_outputs(672) <= (layer4_outputs(178)) or (layer4_outputs(2140));
    layer5_outputs(673) <= (layer4_outputs(889)) or (layer4_outputs(631));
    layer5_outputs(674) <= not((layer4_outputs(1331)) and (layer4_outputs(59)));
    layer5_outputs(675) <= (layer4_outputs(1627)) and not (layer4_outputs(637));
    layer5_outputs(676) <= (layer4_outputs(2113)) xor (layer4_outputs(860));
    layer5_outputs(677) <= not(layer4_outputs(2106));
    layer5_outputs(678) <= not((layer4_outputs(2502)) or (layer4_outputs(1944)));
    layer5_outputs(679) <= not((layer4_outputs(355)) or (layer4_outputs(1110)));
    layer5_outputs(680) <= (layer4_outputs(161)) and (layer4_outputs(297));
    layer5_outputs(681) <= (layer4_outputs(1656)) xor (layer4_outputs(1336));
    layer5_outputs(682) <= layer4_outputs(2262);
    layer5_outputs(683) <= layer4_outputs(1139);
    layer5_outputs(684) <= '1';
    layer5_outputs(685) <= (layer4_outputs(336)) and not (layer4_outputs(1410));
    layer5_outputs(686) <= (layer4_outputs(2457)) xor (layer4_outputs(678));
    layer5_outputs(687) <= not(layer4_outputs(2186)) or (layer4_outputs(363));
    layer5_outputs(688) <= not(layer4_outputs(2205));
    layer5_outputs(689) <= not(layer4_outputs(1532));
    layer5_outputs(690) <= not(layer4_outputs(2212)) or (layer4_outputs(2406));
    layer5_outputs(691) <= (layer4_outputs(442)) xor (layer4_outputs(1819));
    layer5_outputs(692) <= (layer4_outputs(634)) xor (layer4_outputs(1075));
    layer5_outputs(693) <= (layer4_outputs(1651)) xor (layer4_outputs(485));
    layer5_outputs(694) <= (layer4_outputs(2101)) and (layer4_outputs(1815));
    layer5_outputs(695) <= (layer4_outputs(2285)) and not (layer4_outputs(1419));
    layer5_outputs(696) <= not(layer4_outputs(896));
    layer5_outputs(697) <= (layer4_outputs(1877)) or (layer4_outputs(225));
    layer5_outputs(698) <= layer4_outputs(1083);
    layer5_outputs(699) <= not(layer4_outputs(493));
    layer5_outputs(700) <= not(layer4_outputs(1384)) or (layer4_outputs(1904));
    layer5_outputs(701) <= not((layer4_outputs(885)) xor (layer4_outputs(1344)));
    layer5_outputs(702) <= layer4_outputs(2130);
    layer5_outputs(703) <= not((layer4_outputs(50)) or (layer4_outputs(2287)));
    layer5_outputs(704) <= not(layer4_outputs(1880));
    layer5_outputs(705) <= not(layer4_outputs(1775));
    layer5_outputs(706) <= not(layer4_outputs(1433));
    layer5_outputs(707) <= not((layer4_outputs(1815)) xor (layer4_outputs(1082)));
    layer5_outputs(708) <= '1';
    layer5_outputs(709) <= layer4_outputs(1543);
    layer5_outputs(710) <= layer4_outputs(458);
    layer5_outputs(711) <= not((layer4_outputs(916)) and (layer4_outputs(951)));
    layer5_outputs(712) <= (layer4_outputs(492)) or (layer4_outputs(1903));
    layer5_outputs(713) <= not(layer4_outputs(1312));
    layer5_outputs(714) <= layer4_outputs(2107);
    layer5_outputs(715) <= not(layer4_outputs(349)) or (layer4_outputs(357));
    layer5_outputs(716) <= layer4_outputs(915);
    layer5_outputs(717) <= (layer4_outputs(2021)) xor (layer4_outputs(1684));
    layer5_outputs(718) <= layer4_outputs(1366);
    layer5_outputs(719) <= (layer4_outputs(1016)) and (layer4_outputs(663));
    layer5_outputs(720) <= not((layer4_outputs(1358)) or (layer4_outputs(2383)));
    layer5_outputs(721) <= not(layer4_outputs(2200)) or (layer4_outputs(2476));
    layer5_outputs(722) <= (layer4_outputs(2162)) and not (layer4_outputs(2252));
    layer5_outputs(723) <= not(layer4_outputs(2365));
    layer5_outputs(724) <= (layer4_outputs(219)) and (layer4_outputs(2065));
    layer5_outputs(725) <= not(layer4_outputs(308)) or (layer4_outputs(1461));
    layer5_outputs(726) <= (layer4_outputs(1277)) and not (layer4_outputs(2132));
    layer5_outputs(727) <= (layer4_outputs(651)) and not (layer4_outputs(1925));
    layer5_outputs(728) <= (layer4_outputs(963)) or (layer4_outputs(2310));
    layer5_outputs(729) <= layer4_outputs(1385);
    layer5_outputs(730) <= (layer4_outputs(578)) and not (layer4_outputs(422));
    layer5_outputs(731) <= layer4_outputs(1470);
    layer5_outputs(732) <= not(layer4_outputs(1899));
    layer5_outputs(733) <= not((layer4_outputs(2400)) and (layer4_outputs(1181)));
    layer5_outputs(734) <= (layer4_outputs(1455)) or (layer4_outputs(194));
    layer5_outputs(735) <= not(layer4_outputs(208)) or (layer4_outputs(1939));
    layer5_outputs(736) <= not(layer4_outputs(1329));
    layer5_outputs(737) <= (layer4_outputs(1886)) and not (layer4_outputs(806));
    layer5_outputs(738) <= not(layer4_outputs(350));
    layer5_outputs(739) <= (layer4_outputs(323)) and not (layer4_outputs(1326));
    layer5_outputs(740) <= not(layer4_outputs(2545));
    layer5_outputs(741) <= not(layer4_outputs(1770));
    layer5_outputs(742) <= not(layer4_outputs(1527));
    layer5_outputs(743) <= (layer4_outputs(1232)) and (layer4_outputs(2551));
    layer5_outputs(744) <= not(layer4_outputs(2056)) or (layer4_outputs(1924));
    layer5_outputs(745) <= not(layer4_outputs(108)) or (layer4_outputs(1252));
    layer5_outputs(746) <= layer4_outputs(842);
    layer5_outputs(747) <= layer4_outputs(2314);
    layer5_outputs(748) <= not(layer4_outputs(2087));
    layer5_outputs(749) <= not(layer4_outputs(2040));
    layer5_outputs(750) <= layer4_outputs(2136);
    layer5_outputs(751) <= (layer4_outputs(1179)) and (layer4_outputs(662));
    layer5_outputs(752) <= (layer4_outputs(994)) and not (layer4_outputs(654));
    layer5_outputs(753) <= (layer4_outputs(1091)) and not (layer4_outputs(1264));
    layer5_outputs(754) <= layer4_outputs(669);
    layer5_outputs(755) <= layer4_outputs(2290);
    layer5_outputs(756) <= not(layer4_outputs(1057));
    layer5_outputs(757) <= not(layer4_outputs(886)) or (layer4_outputs(1610));
    layer5_outputs(758) <= layer4_outputs(182);
    layer5_outputs(759) <= layer4_outputs(1718);
    layer5_outputs(760) <= (layer4_outputs(671)) and not (layer4_outputs(271));
    layer5_outputs(761) <= not(layer4_outputs(991));
    layer5_outputs(762) <= not((layer4_outputs(2135)) or (layer4_outputs(1215)));
    layer5_outputs(763) <= '1';
    layer5_outputs(764) <= not(layer4_outputs(1618));
    layer5_outputs(765) <= (layer4_outputs(1365)) xor (layer4_outputs(141));
    layer5_outputs(766) <= (layer4_outputs(2547)) xor (layer4_outputs(2053));
    layer5_outputs(767) <= not((layer4_outputs(536)) and (layer4_outputs(1879)));
    layer5_outputs(768) <= not(layer4_outputs(833));
    layer5_outputs(769) <= not(layer4_outputs(1930));
    layer5_outputs(770) <= layer4_outputs(2226);
    layer5_outputs(771) <= layer4_outputs(2289);
    layer5_outputs(772) <= not(layer4_outputs(1052));
    layer5_outputs(773) <= not(layer4_outputs(931)) or (layer4_outputs(552));
    layer5_outputs(774) <= (layer4_outputs(1312)) and not (layer4_outputs(571));
    layer5_outputs(775) <= not(layer4_outputs(1589)) or (layer4_outputs(391));
    layer5_outputs(776) <= not(layer4_outputs(595)) or (layer4_outputs(2090));
    layer5_outputs(777) <= layer4_outputs(2333);
    layer5_outputs(778) <= layer4_outputs(337);
    layer5_outputs(779) <= layer4_outputs(1664);
    layer5_outputs(780) <= layer4_outputs(27);
    layer5_outputs(781) <= not(layer4_outputs(1361)) or (layer4_outputs(1838));
    layer5_outputs(782) <= not(layer4_outputs(574));
    layer5_outputs(783) <= not(layer4_outputs(103));
    layer5_outputs(784) <= (layer4_outputs(1116)) xor (layer4_outputs(843));
    layer5_outputs(785) <= layer4_outputs(2203);
    layer5_outputs(786) <= layer4_outputs(1025);
    layer5_outputs(787) <= layer4_outputs(149);
    layer5_outputs(788) <= layer4_outputs(1934);
    layer5_outputs(789) <= layer4_outputs(867);
    layer5_outputs(790) <= (layer4_outputs(1894)) and not (layer4_outputs(816));
    layer5_outputs(791) <= (layer4_outputs(2195)) and not (layer4_outputs(1313));
    layer5_outputs(792) <= not((layer4_outputs(812)) xor (layer4_outputs(947)));
    layer5_outputs(793) <= not(layer4_outputs(2253));
    layer5_outputs(794) <= not(layer4_outputs(567));
    layer5_outputs(795) <= layer4_outputs(1746);
    layer5_outputs(796) <= layer4_outputs(582);
    layer5_outputs(797) <= (layer4_outputs(891)) xor (layer4_outputs(2536));
    layer5_outputs(798) <= not(layer4_outputs(240)) or (layer4_outputs(2027));
    layer5_outputs(799) <= not((layer4_outputs(191)) xor (layer4_outputs(1983)));
    layer5_outputs(800) <= layer4_outputs(986);
    layer5_outputs(801) <= not((layer4_outputs(580)) xor (layer4_outputs(1468)));
    layer5_outputs(802) <= not((layer4_outputs(1187)) xor (layer4_outputs(1856)));
    layer5_outputs(803) <= not((layer4_outputs(591)) and (layer4_outputs(2296)));
    layer5_outputs(804) <= layer4_outputs(1544);
    layer5_outputs(805) <= (layer4_outputs(1416)) and not (layer4_outputs(22));
    layer5_outputs(806) <= (layer4_outputs(2334)) xor (layer4_outputs(2484));
    layer5_outputs(807) <= (layer4_outputs(460)) and not (layer4_outputs(1969));
    layer5_outputs(808) <= '0';
    layer5_outputs(809) <= layer4_outputs(777);
    layer5_outputs(810) <= not(layer4_outputs(2389));
    layer5_outputs(811) <= layer4_outputs(514);
    layer5_outputs(812) <= layer4_outputs(557);
    layer5_outputs(813) <= not(layer4_outputs(1433));
    layer5_outputs(814) <= layer4_outputs(444);
    layer5_outputs(815) <= layer4_outputs(1126);
    layer5_outputs(816) <= layer4_outputs(2430);
    layer5_outputs(817) <= not(layer4_outputs(949));
    layer5_outputs(818) <= not(layer4_outputs(759));
    layer5_outputs(819) <= (layer4_outputs(793)) or (layer4_outputs(1799));
    layer5_outputs(820) <= not((layer4_outputs(2051)) or (layer4_outputs(1207)));
    layer5_outputs(821) <= layer4_outputs(2137);
    layer5_outputs(822) <= layer4_outputs(90);
    layer5_outputs(823) <= not(layer4_outputs(2101));
    layer5_outputs(824) <= not((layer4_outputs(602)) and (layer4_outputs(1972)));
    layer5_outputs(825) <= not(layer4_outputs(1133));
    layer5_outputs(826) <= not(layer4_outputs(538));
    layer5_outputs(827) <= layer4_outputs(1454);
    layer5_outputs(828) <= not((layer4_outputs(2252)) or (layer4_outputs(784)));
    layer5_outputs(829) <= layer4_outputs(2071);
    layer5_outputs(830) <= (layer4_outputs(983)) and not (layer4_outputs(1358));
    layer5_outputs(831) <= not((layer4_outputs(857)) xor (layer4_outputs(1914)));
    layer5_outputs(832) <= not((layer4_outputs(81)) xor (layer4_outputs(1350)));
    layer5_outputs(833) <= not(layer4_outputs(2417));
    layer5_outputs(834) <= (layer4_outputs(2016)) and not (layer4_outputs(310));
    layer5_outputs(835) <= not((layer4_outputs(379)) and (layer4_outputs(508)));
    layer5_outputs(836) <= (layer4_outputs(2537)) xor (layer4_outputs(45));
    layer5_outputs(837) <= not(layer4_outputs(1529));
    layer5_outputs(838) <= not((layer4_outputs(712)) or (layer4_outputs(1612)));
    layer5_outputs(839) <= not(layer4_outputs(1992));
    layer5_outputs(840) <= layer4_outputs(1776);
    layer5_outputs(841) <= (layer4_outputs(1359)) xor (layer4_outputs(1992));
    layer5_outputs(842) <= not(layer4_outputs(559));
    layer5_outputs(843) <= (layer4_outputs(1321)) xor (layer4_outputs(1577));
    layer5_outputs(844) <= not((layer4_outputs(449)) or (layer4_outputs(439)));
    layer5_outputs(845) <= not((layer4_outputs(1807)) or (layer4_outputs(193)));
    layer5_outputs(846) <= '0';
    layer5_outputs(847) <= (layer4_outputs(1337)) or (layer4_outputs(896));
    layer5_outputs(848) <= not(layer4_outputs(1394));
    layer5_outputs(849) <= (layer4_outputs(1141)) and not (layer4_outputs(1781));
    layer5_outputs(850) <= layer4_outputs(1845);
    layer5_outputs(851) <= not((layer4_outputs(1022)) and (layer4_outputs(279)));
    layer5_outputs(852) <= not((layer4_outputs(1720)) and (layer4_outputs(1733)));
    layer5_outputs(853) <= layer4_outputs(1276);
    layer5_outputs(854) <= (layer4_outputs(2048)) xor (layer4_outputs(1548));
    layer5_outputs(855) <= (layer4_outputs(2322)) and (layer4_outputs(2360));
    layer5_outputs(856) <= not(layer4_outputs(2194));
    layer5_outputs(857) <= (layer4_outputs(927)) and not (layer4_outputs(1174));
    layer5_outputs(858) <= not(layer4_outputs(445));
    layer5_outputs(859) <= not((layer4_outputs(2469)) or (layer4_outputs(329)));
    layer5_outputs(860) <= (layer4_outputs(327)) and not (layer4_outputs(656));
    layer5_outputs(861) <= not((layer4_outputs(1922)) or (layer4_outputs(685)));
    layer5_outputs(862) <= layer4_outputs(308);
    layer5_outputs(863) <= (layer4_outputs(2204)) and not (layer4_outputs(2245));
    layer5_outputs(864) <= (layer4_outputs(1591)) xor (layer4_outputs(1710));
    layer5_outputs(865) <= (layer4_outputs(2117)) and not (layer4_outputs(2520));
    layer5_outputs(866) <= (layer4_outputs(2389)) and (layer4_outputs(1587));
    layer5_outputs(867) <= layer4_outputs(755);
    layer5_outputs(868) <= (layer4_outputs(1781)) and not (layer4_outputs(1224));
    layer5_outputs(869) <= not((layer4_outputs(301)) xor (layer4_outputs(1446)));
    layer5_outputs(870) <= layer4_outputs(2369);
    layer5_outputs(871) <= not(layer4_outputs(326));
    layer5_outputs(872) <= not((layer4_outputs(449)) or (layer4_outputs(145)));
    layer5_outputs(873) <= not((layer4_outputs(125)) xor (layer4_outputs(446)));
    layer5_outputs(874) <= (layer4_outputs(830)) and not (layer4_outputs(275));
    layer5_outputs(875) <= not(layer4_outputs(1495)) or (layer4_outputs(1800));
    layer5_outputs(876) <= layer4_outputs(1521);
    layer5_outputs(877) <= (layer4_outputs(625)) and (layer4_outputs(276));
    layer5_outputs(878) <= (layer4_outputs(1928)) and not (layer4_outputs(664));
    layer5_outputs(879) <= (layer4_outputs(1177)) and not (layer4_outputs(190));
    layer5_outputs(880) <= not((layer4_outputs(1506)) xor (layer4_outputs(1993)));
    layer5_outputs(881) <= layer4_outputs(1377);
    layer5_outputs(882) <= not(layer4_outputs(1624)) or (layer4_outputs(636));
    layer5_outputs(883) <= not(layer4_outputs(77)) or (layer4_outputs(250));
    layer5_outputs(884) <= not((layer4_outputs(301)) or (layer4_outputs(29)));
    layer5_outputs(885) <= not(layer4_outputs(1703));
    layer5_outputs(886) <= not(layer4_outputs(393));
    layer5_outputs(887) <= (layer4_outputs(129)) and not (layer4_outputs(499));
    layer5_outputs(888) <= not(layer4_outputs(1491));
    layer5_outputs(889) <= not(layer4_outputs(1591)) or (layer4_outputs(316));
    layer5_outputs(890) <= '1';
    layer5_outputs(891) <= layer4_outputs(166);
    layer5_outputs(892) <= layer4_outputs(198);
    layer5_outputs(893) <= '0';
    layer5_outputs(894) <= not(layer4_outputs(2282));
    layer5_outputs(895) <= (layer4_outputs(1913)) and not (layer4_outputs(2506));
    layer5_outputs(896) <= layer4_outputs(2431);
    layer5_outputs(897) <= not(layer4_outputs(2049));
    layer5_outputs(898) <= (layer4_outputs(609)) and (layer4_outputs(159));
    layer5_outputs(899) <= (layer4_outputs(172)) and not (layer4_outputs(1933));
    layer5_outputs(900) <= not(layer4_outputs(1521));
    layer5_outputs(901) <= (layer4_outputs(481)) and (layer4_outputs(2520));
    layer5_outputs(902) <= layer4_outputs(1300);
    layer5_outputs(903) <= (layer4_outputs(394)) and (layer4_outputs(1372));
    layer5_outputs(904) <= (layer4_outputs(1906)) and (layer4_outputs(187));
    layer5_outputs(905) <= not((layer4_outputs(2255)) and (layer4_outputs(2263)));
    layer5_outputs(906) <= not(layer4_outputs(465));
    layer5_outputs(907) <= (layer4_outputs(1309)) and (layer4_outputs(877));
    layer5_outputs(908) <= (layer4_outputs(1074)) and (layer4_outputs(1738));
    layer5_outputs(909) <= '0';
    layer5_outputs(910) <= layer4_outputs(971);
    layer5_outputs(911) <= (layer4_outputs(146)) or (layer4_outputs(1606));
    layer5_outputs(912) <= not(layer4_outputs(1909));
    layer5_outputs(913) <= layer4_outputs(700);
    layer5_outputs(914) <= (layer4_outputs(180)) and (layer4_outputs(2475));
    layer5_outputs(915) <= not(layer4_outputs(1485)) or (layer4_outputs(1865));
    layer5_outputs(916) <= layer4_outputs(2121);
    layer5_outputs(917) <= not(layer4_outputs(862));
    layer5_outputs(918) <= layer4_outputs(1243);
    layer5_outputs(919) <= not(layer4_outputs(1337));
    layer5_outputs(920) <= not(layer4_outputs(16));
    layer5_outputs(921) <= not(layer4_outputs(1600));
    layer5_outputs(922) <= not(layer4_outputs(1806));
    layer5_outputs(923) <= not(layer4_outputs(2476));
    layer5_outputs(924) <= not(layer4_outputs(1536)) or (layer4_outputs(830));
    layer5_outputs(925) <= (layer4_outputs(132)) xor (layer4_outputs(521));
    layer5_outputs(926) <= (layer4_outputs(1895)) or (layer4_outputs(317));
    layer5_outputs(927) <= not(layer4_outputs(721));
    layer5_outputs(928) <= not((layer4_outputs(2324)) xor (layer4_outputs(294)));
    layer5_outputs(929) <= (layer4_outputs(1043)) or (layer4_outputs(12));
    layer5_outputs(930) <= (layer4_outputs(824)) or (layer4_outputs(392));
    layer5_outputs(931) <= (layer4_outputs(2078)) xor (layer4_outputs(235));
    layer5_outputs(932) <= '0';
    layer5_outputs(933) <= not(layer4_outputs(2508));
    layer5_outputs(934) <= not((layer4_outputs(166)) and (layer4_outputs(523)));
    layer5_outputs(935) <= not(layer4_outputs(622));
    layer5_outputs(936) <= (layer4_outputs(1052)) and not (layer4_outputs(1049));
    layer5_outputs(937) <= layer4_outputs(739);
    layer5_outputs(938) <= not(layer4_outputs(2255));
    layer5_outputs(939) <= not((layer4_outputs(1229)) and (layer4_outputs(1805)));
    layer5_outputs(940) <= not((layer4_outputs(18)) and (layer4_outputs(819)));
    layer5_outputs(941) <= not(layer4_outputs(1974)) or (layer4_outputs(1648));
    layer5_outputs(942) <= not(layer4_outputs(527));
    layer5_outputs(943) <= not(layer4_outputs(988)) or (layer4_outputs(1164));
    layer5_outputs(944) <= not(layer4_outputs(1672));
    layer5_outputs(945) <= layer4_outputs(1257);
    layer5_outputs(946) <= (layer4_outputs(2372)) xor (layer4_outputs(120));
    layer5_outputs(947) <= (layer4_outputs(465)) and (layer4_outputs(903));
    layer5_outputs(948) <= layer4_outputs(1321);
    layer5_outputs(949) <= not(layer4_outputs(2202));
    layer5_outputs(950) <= layer4_outputs(1761);
    layer5_outputs(951) <= not(layer4_outputs(2016)) or (layer4_outputs(1245));
    layer5_outputs(952) <= not(layer4_outputs(1319)) or (layer4_outputs(1317));
    layer5_outputs(953) <= not(layer4_outputs(2213));
    layer5_outputs(954) <= (layer4_outputs(258)) and (layer4_outputs(2481));
    layer5_outputs(955) <= not(layer4_outputs(1569));
    layer5_outputs(956) <= (layer4_outputs(189)) and (layer4_outputs(641));
    layer5_outputs(957) <= '1';
    layer5_outputs(958) <= not(layer4_outputs(364));
    layer5_outputs(959) <= layer4_outputs(771);
    layer5_outputs(960) <= layer4_outputs(513);
    layer5_outputs(961) <= not(layer4_outputs(418));
    layer5_outputs(962) <= (layer4_outputs(2091)) xor (layer4_outputs(186));
    layer5_outputs(963) <= (layer4_outputs(1346)) and not (layer4_outputs(2415));
    layer5_outputs(964) <= layer4_outputs(654);
    layer5_outputs(965) <= '0';
    layer5_outputs(966) <= not(layer4_outputs(1518));
    layer5_outputs(967) <= not(layer4_outputs(1618));
    layer5_outputs(968) <= layer4_outputs(2542);
    layer5_outputs(969) <= layer4_outputs(123);
    layer5_outputs(970) <= not(layer4_outputs(408)) or (layer4_outputs(2445));
    layer5_outputs(971) <= layer4_outputs(1056);
    layer5_outputs(972) <= (layer4_outputs(2017)) or (layer4_outputs(1859));
    layer5_outputs(973) <= not(layer4_outputs(1663)) or (layer4_outputs(233));
    layer5_outputs(974) <= layer4_outputs(2457);
    layer5_outputs(975) <= not((layer4_outputs(1427)) and (layer4_outputs(1354)));
    layer5_outputs(976) <= not(layer4_outputs(613));
    layer5_outputs(977) <= '0';
    layer5_outputs(978) <= layer4_outputs(1652);
    layer5_outputs(979) <= not((layer4_outputs(1699)) or (layer4_outputs(526)));
    layer5_outputs(980) <= not(layer4_outputs(497)) or (layer4_outputs(899));
    layer5_outputs(981) <= '0';
    layer5_outputs(982) <= not(layer4_outputs(1605)) or (layer4_outputs(1328));
    layer5_outputs(983) <= layer4_outputs(2362);
    layer5_outputs(984) <= not(layer4_outputs(1523));
    layer5_outputs(985) <= (layer4_outputs(115)) and not (layer4_outputs(655));
    layer5_outputs(986) <= not(layer4_outputs(1905));
    layer5_outputs(987) <= (layer4_outputs(1647)) and not (layer4_outputs(1816));
    layer5_outputs(988) <= (layer4_outputs(871)) and not (layer4_outputs(121));
    layer5_outputs(989) <= layer4_outputs(119);
    layer5_outputs(990) <= layer4_outputs(2266);
    layer5_outputs(991) <= (layer4_outputs(2112)) and not (layer4_outputs(676));
    layer5_outputs(992) <= not(layer4_outputs(1822)) or (layer4_outputs(468));
    layer5_outputs(993) <= (layer4_outputs(1248)) and not (layer4_outputs(691));
    layer5_outputs(994) <= not(layer4_outputs(179)) or (layer4_outputs(619));
    layer5_outputs(995) <= '1';
    layer5_outputs(996) <= layer4_outputs(978);
    layer5_outputs(997) <= layer4_outputs(2555);
    layer5_outputs(998) <= '0';
    layer5_outputs(999) <= not(layer4_outputs(1218)) or (layer4_outputs(626));
    layer5_outputs(1000) <= (layer4_outputs(1641)) and not (layer4_outputs(922));
    layer5_outputs(1001) <= layer4_outputs(1808);
    layer5_outputs(1002) <= '1';
    layer5_outputs(1003) <= not(layer4_outputs(2345));
    layer5_outputs(1004) <= layer4_outputs(1409);
    layer5_outputs(1005) <= (layer4_outputs(1481)) and (layer4_outputs(1608));
    layer5_outputs(1006) <= '1';
    layer5_outputs(1007) <= not(layer4_outputs(2072)) or (layer4_outputs(214));
    layer5_outputs(1008) <= layer4_outputs(1798);
    layer5_outputs(1009) <= not((layer4_outputs(2241)) and (layer4_outputs(195)));
    layer5_outputs(1010) <= not(layer4_outputs(673));
    layer5_outputs(1011) <= not((layer4_outputs(954)) and (layer4_outputs(2063)));
    layer5_outputs(1012) <= not(layer4_outputs(1797));
    layer5_outputs(1013) <= not(layer4_outputs(2251));
    layer5_outputs(1014) <= not(layer4_outputs(1172));
    layer5_outputs(1015) <= not((layer4_outputs(757)) and (layer4_outputs(2076)));
    layer5_outputs(1016) <= layer4_outputs(834);
    layer5_outputs(1017) <= not(layer4_outputs(1155)) or (layer4_outputs(2429));
    layer5_outputs(1018) <= not((layer4_outputs(1416)) or (layer4_outputs(1302)));
    layer5_outputs(1019) <= not((layer4_outputs(1582)) or (layer4_outputs(434)));
    layer5_outputs(1020) <= '0';
    layer5_outputs(1021) <= layer4_outputs(1557);
    layer5_outputs(1022) <= (layer4_outputs(355)) or (layer4_outputs(2516));
    layer5_outputs(1023) <= (layer4_outputs(2199)) or (layer4_outputs(2549));
    layer5_outputs(1024) <= not(layer4_outputs(1875));
    layer5_outputs(1025) <= not(layer4_outputs(2307));
    layer5_outputs(1026) <= not(layer4_outputs(2244));
    layer5_outputs(1027) <= not((layer4_outputs(2095)) xor (layer4_outputs(854)));
    layer5_outputs(1028) <= not(layer4_outputs(1441));
    layer5_outputs(1029) <= not((layer4_outputs(2295)) or (layer4_outputs(2197)));
    layer5_outputs(1030) <= (layer4_outputs(2555)) and not (layer4_outputs(943));
    layer5_outputs(1031) <= not(layer4_outputs(67));
    layer5_outputs(1032) <= not(layer4_outputs(715)) or (layer4_outputs(344));
    layer5_outputs(1033) <= (layer4_outputs(2270)) and (layer4_outputs(2052));
    layer5_outputs(1034) <= not(layer4_outputs(760)) or (layer4_outputs(1553));
    layer5_outputs(1035) <= not(layer4_outputs(573)) or (layer4_outputs(1010));
    layer5_outputs(1036) <= (layer4_outputs(679)) and (layer4_outputs(1362));
    layer5_outputs(1037) <= layer4_outputs(1875);
    layer5_outputs(1038) <= (layer4_outputs(2088)) and (layer4_outputs(1176));
    layer5_outputs(1039) <= not(layer4_outputs(1261));
    layer5_outputs(1040) <= not((layer4_outputs(1679)) xor (layer4_outputs(368)));
    layer5_outputs(1041) <= layer4_outputs(260);
    layer5_outputs(1042) <= (layer4_outputs(2125)) and not (layer4_outputs(1861));
    layer5_outputs(1043) <= layer4_outputs(1885);
    layer5_outputs(1044) <= (layer4_outputs(1108)) or (layer4_outputs(1170));
    layer5_outputs(1045) <= not(layer4_outputs(1515));
    layer5_outputs(1046) <= layer4_outputs(514);
    layer5_outputs(1047) <= not(layer4_outputs(838));
    layer5_outputs(1048) <= layer4_outputs(220);
    layer5_outputs(1049) <= not((layer4_outputs(1818)) xor (layer4_outputs(677)));
    layer5_outputs(1050) <= not(layer4_outputs(1262));
    layer5_outputs(1051) <= not(layer4_outputs(1162));
    layer5_outputs(1052) <= not((layer4_outputs(14)) xor (layer4_outputs(969)));
    layer5_outputs(1053) <= (layer4_outputs(1743)) and (layer4_outputs(490));
    layer5_outputs(1054) <= (layer4_outputs(998)) xor (layer4_outputs(900));
    layer5_outputs(1055) <= '1';
    layer5_outputs(1056) <= layer4_outputs(1501);
    layer5_outputs(1057) <= not(layer4_outputs(1050)) or (layer4_outputs(417));
    layer5_outputs(1058) <= layer4_outputs(2337);
    layer5_outputs(1059) <= (layer4_outputs(7)) and not (layer4_outputs(1620));
    layer5_outputs(1060) <= not(layer4_outputs(2354)) or (layer4_outputs(1426));
    layer5_outputs(1061) <= layer4_outputs(789);
    layer5_outputs(1062) <= layer4_outputs(451);
    layer5_outputs(1063) <= '0';
    layer5_outputs(1064) <= (layer4_outputs(2240)) and (layer4_outputs(443));
    layer5_outputs(1065) <= not((layer4_outputs(1378)) xor (layer4_outputs(71)));
    layer5_outputs(1066) <= not(layer4_outputs(708));
    layer5_outputs(1067) <= not(layer4_outputs(2157)) or (layer4_outputs(137));
    layer5_outputs(1068) <= not(layer4_outputs(802));
    layer5_outputs(1069) <= not(layer4_outputs(2198));
    layer5_outputs(1070) <= layer4_outputs(1404);
    layer5_outputs(1071) <= '0';
    layer5_outputs(1072) <= layer4_outputs(1051);
    layer5_outputs(1073) <= not(layer4_outputs(1780)) or (layer4_outputs(164));
    layer5_outputs(1074) <= not((layer4_outputs(1039)) xor (layer4_outputs(1277)));
    layer5_outputs(1075) <= not((layer4_outputs(2325)) and (layer4_outputs(154)));
    layer5_outputs(1076) <= (layer4_outputs(24)) and not (layer4_outputs(609));
    layer5_outputs(1077) <= layer4_outputs(2442);
    layer5_outputs(1078) <= not(layer4_outputs(1182));
    layer5_outputs(1079) <= (layer4_outputs(2183)) and not (layer4_outputs(139));
    layer5_outputs(1080) <= not((layer4_outputs(2170)) or (layer4_outputs(433)));
    layer5_outputs(1081) <= (layer4_outputs(2514)) or (layer4_outputs(2501));
    layer5_outputs(1082) <= layer4_outputs(139);
    layer5_outputs(1083) <= layer4_outputs(2126);
    layer5_outputs(1084) <= (layer4_outputs(5)) xor (layer4_outputs(2225));
    layer5_outputs(1085) <= not(layer4_outputs(1896));
    layer5_outputs(1086) <= not(layer4_outputs(2425));
    layer5_outputs(1087) <= '0';
    layer5_outputs(1088) <= (layer4_outputs(24)) and not (layer4_outputs(1795));
    layer5_outputs(1089) <= layer4_outputs(239);
    layer5_outputs(1090) <= not((layer4_outputs(495)) or (layer4_outputs(3)));
    layer5_outputs(1091) <= not(layer4_outputs(445));
    layer5_outputs(1092) <= '0';
    layer5_outputs(1093) <= not((layer4_outputs(880)) or (layer4_outputs(2030)));
    layer5_outputs(1094) <= not(layer4_outputs(864));
    layer5_outputs(1095) <= not(layer4_outputs(1434));
    layer5_outputs(1096) <= not(layer4_outputs(1347));
    layer5_outputs(1097) <= layer4_outputs(1712);
    layer5_outputs(1098) <= layer4_outputs(1425);
    layer5_outputs(1099) <= (layer4_outputs(1384)) and not (layer4_outputs(1747));
    layer5_outputs(1100) <= not(layer4_outputs(1090)) or (layer4_outputs(49));
    layer5_outputs(1101) <= not(layer4_outputs(140));
    layer5_outputs(1102) <= layer4_outputs(1841);
    layer5_outputs(1103) <= (layer4_outputs(1176)) and not (layer4_outputs(2008));
    layer5_outputs(1104) <= (layer4_outputs(2302)) xor (layer4_outputs(604));
    layer5_outputs(1105) <= not(layer4_outputs(2558));
    layer5_outputs(1106) <= not(layer4_outputs(2174));
    layer5_outputs(1107) <= not((layer4_outputs(1029)) or (layer4_outputs(423)));
    layer5_outputs(1108) <= not(layer4_outputs(2428)) or (layer4_outputs(1214));
    layer5_outputs(1109) <= not((layer4_outputs(1195)) or (layer4_outputs(559)));
    layer5_outputs(1110) <= (layer4_outputs(1580)) xor (layer4_outputs(469));
    layer5_outputs(1111) <= layer4_outputs(1884);
    layer5_outputs(1112) <= layer4_outputs(427);
    layer5_outputs(1113) <= not(layer4_outputs(1173));
    layer5_outputs(1114) <= layer4_outputs(2317);
    layer5_outputs(1115) <= (layer4_outputs(2309)) and not (layer4_outputs(2393));
    layer5_outputs(1116) <= (layer4_outputs(1982)) or (layer4_outputs(1981));
    layer5_outputs(1117) <= layer4_outputs(777);
    layer5_outputs(1118) <= not((layer4_outputs(1472)) xor (layer4_outputs(2047)));
    layer5_outputs(1119) <= layer4_outputs(2462);
    layer5_outputs(1120) <= layer4_outputs(888);
    layer5_outputs(1121) <= (layer4_outputs(2514)) and not (layer4_outputs(692));
    layer5_outputs(1122) <= not((layer4_outputs(2062)) xor (layer4_outputs(62)));
    layer5_outputs(1123) <= not((layer4_outputs(730)) xor (layer4_outputs(793)));
    layer5_outputs(1124) <= (layer4_outputs(306)) and not (layer4_outputs(2500));
    layer5_outputs(1125) <= layer4_outputs(1100);
    layer5_outputs(1126) <= (layer4_outputs(1009)) and not (layer4_outputs(995));
    layer5_outputs(1127) <= layer4_outputs(2419);
    layer5_outputs(1128) <= layer4_outputs(1430);
    layer5_outputs(1129) <= not(layer4_outputs(141));
    layer5_outputs(1130) <= not(layer4_outputs(1848));
    layer5_outputs(1131) <= not((layer4_outputs(1833)) or (layer4_outputs(56)));
    layer5_outputs(1132) <= (layer4_outputs(866)) and (layer4_outputs(788));
    layer5_outputs(1133) <= layer4_outputs(1103);
    layer5_outputs(1134) <= not((layer4_outputs(1852)) and (layer4_outputs(1402)));
    layer5_outputs(1135) <= (layer4_outputs(85)) xor (layer4_outputs(251));
    layer5_outputs(1136) <= (layer4_outputs(2263)) xor (layer4_outputs(2275));
    layer5_outputs(1137) <= (layer4_outputs(2238)) and not (layer4_outputs(1198));
    layer5_outputs(1138) <= layer4_outputs(977);
    layer5_outputs(1139) <= (layer4_outputs(546)) and (layer4_outputs(1732));
    layer5_outputs(1140) <= layer4_outputs(783);
    layer5_outputs(1141) <= not(layer4_outputs(155));
    layer5_outputs(1142) <= not(layer4_outputs(562)) or (layer4_outputs(117));
    layer5_outputs(1143) <= not(layer4_outputs(76));
    layer5_outputs(1144) <= not((layer4_outputs(1060)) or (layer4_outputs(2374)));
    layer5_outputs(1145) <= (layer4_outputs(2483)) and not (layer4_outputs(623));
    layer5_outputs(1146) <= not(layer4_outputs(2366));
    layer5_outputs(1147) <= (layer4_outputs(1557)) and not (layer4_outputs(1923));
    layer5_outputs(1148) <= layer4_outputs(47);
    layer5_outputs(1149) <= layer4_outputs(1131);
    layer5_outputs(1150) <= (layer4_outputs(2425)) or (layer4_outputs(1219));
    layer5_outputs(1151) <= not((layer4_outputs(602)) and (layer4_outputs(79)));
    layer5_outputs(1152) <= '0';
    layer5_outputs(1153) <= layer4_outputs(273);
    layer5_outputs(1154) <= layer4_outputs(282);
    layer5_outputs(1155) <= not((layer4_outputs(2254)) or (layer4_outputs(769)));
    layer5_outputs(1156) <= not((layer4_outputs(1122)) xor (layer4_outputs(2327)));
    layer5_outputs(1157) <= (layer4_outputs(2407)) or (layer4_outputs(87));
    layer5_outputs(1158) <= not(layer4_outputs(2308));
    layer5_outputs(1159) <= layer4_outputs(1000);
    layer5_outputs(1160) <= layer4_outputs(2055);
    layer5_outputs(1161) <= not(layer4_outputs(1473));
    layer5_outputs(1162) <= not(layer4_outputs(234));
    layer5_outputs(1163) <= layer4_outputs(135);
    layer5_outputs(1164) <= not(layer4_outputs(1889));
    layer5_outputs(1165) <= layer4_outputs(2490);
    layer5_outputs(1166) <= not(layer4_outputs(1711));
    layer5_outputs(1167) <= not(layer4_outputs(170));
    layer5_outputs(1168) <= (layer4_outputs(2305)) and (layer4_outputs(72));
    layer5_outputs(1169) <= not(layer4_outputs(115));
    layer5_outputs(1170) <= layer4_outputs(515);
    layer5_outputs(1171) <= not(layer4_outputs(64));
    layer5_outputs(1172) <= not(layer4_outputs(2314)) or (layer4_outputs(1672));
    layer5_outputs(1173) <= layer4_outputs(1650);
    layer5_outputs(1174) <= '1';
    layer5_outputs(1175) <= layer4_outputs(1768);
    layer5_outputs(1176) <= not((layer4_outputs(1824)) or (layer4_outputs(2247)));
    layer5_outputs(1177) <= not(layer4_outputs(374)) or (layer4_outputs(1331));
    layer5_outputs(1178) <= (layer4_outputs(1245)) and not (layer4_outputs(2108));
    layer5_outputs(1179) <= not(layer4_outputs(2440));
    layer5_outputs(1180) <= not((layer4_outputs(2120)) xor (layer4_outputs(1696)));
    layer5_outputs(1181) <= not((layer4_outputs(1108)) or (layer4_outputs(1240)));
    layer5_outputs(1182) <= (layer4_outputs(873)) xor (layer4_outputs(2180));
    layer5_outputs(1183) <= layer4_outputs(1607);
    layer5_outputs(1184) <= not((layer4_outputs(607)) xor (layer4_outputs(440)));
    layer5_outputs(1185) <= (layer4_outputs(585)) and not (layer4_outputs(1315));
    layer5_outputs(1186) <= not(layer4_outputs(1783));
    layer5_outputs(1187) <= not((layer4_outputs(2212)) xor (layer4_outputs(405)));
    layer5_outputs(1188) <= layer4_outputs(26);
    layer5_outputs(1189) <= not(layer4_outputs(1980));
    layer5_outputs(1190) <= not(layer4_outputs(1427));
    layer5_outputs(1191) <= layer4_outputs(681);
    layer5_outputs(1192) <= layer4_outputs(528);
    layer5_outputs(1193) <= (layer4_outputs(853)) xor (layer4_outputs(427));
    layer5_outputs(1194) <= not((layer4_outputs(1634)) and (layer4_outputs(192)));
    layer5_outputs(1195) <= not(layer4_outputs(2394));
    layer5_outputs(1196) <= not((layer4_outputs(972)) xor (layer4_outputs(2139)));
    layer5_outputs(1197) <= layer4_outputs(2526);
    layer5_outputs(1198) <= layer4_outputs(436);
    layer5_outputs(1199) <= not(layer4_outputs(2453));
    layer5_outputs(1200) <= not(layer4_outputs(944));
    layer5_outputs(1201) <= layer4_outputs(1460);
    layer5_outputs(1202) <= (layer4_outputs(1403)) and not (layer4_outputs(1177));
    layer5_outputs(1203) <= layer4_outputs(1905);
    layer5_outputs(1204) <= not(layer4_outputs(623));
    layer5_outputs(1205) <= layer4_outputs(1787);
    layer5_outputs(1206) <= (layer4_outputs(1658)) and not (layer4_outputs(1241));
    layer5_outputs(1207) <= (layer4_outputs(953)) and not (layer4_outputs(1956));
    layer5_outputs(1208) <= layer4_outputs(2088);
    layer5_outputs(1209) <= not(layer4_outputs(844));
    layer5_outputs(1210) <= (layer4_outputs(1749)) and not (layer4_outputs(954));
    layer5_outputs(1211) <= not(layer4_outputs(709));
    layer5_outputs(1212) <= not((layer4_outputs(1821)) and (layer4_outputs(1950)));
    layer5_outputs(1213) <= not(layer4_outputs(1223));
    layer5_outputs(1214) <= layer4_outputs(1998);
    layer5_outputs(1215) <= (layer4_outputs(1264)) or (layer4_outputs(2410));
    layer5_outputs(1216) <= not((layer4_outputs(657)) xor (layer4_outputs(1830)));
    layer5_outputs(1217) <= layer4_outputs(816);
    layer5_outputs(1218) <= layer4_outputs(2529);
    layer5_outputs(1219) <= layer4_outputs(2122);
    layer5_outputs(1220) <= not(layer4_outputs(510));
    layer5_outputs(1221) <= not(layer4_outputs(1601));
    layer5_outputs(1222) <= not(layer4_outputs(429)) or (layer4_outputs(764));
    layer5_outputs(1223) <= layer4_outputs(386);
    layer5_outputs(1224) <= (layer4_outputs(1826)) xor (layer4_outputs(2326));
    layer5_outputs(1225) <= (layer4_outputs(137)) and not (layer4_outputs(397));
    layer5_outputs(1226) <= layer4_outputs(1619);
    layer5_outputs(1227) <= not((layer4_outputs(2260)) and (layer4_outputs(820)));
    layer5_outputs(1228) <= layer4_outputs(757);
    layer5_outputs(1229) <= (layer4_outputs(2217)) xor (layer4_outputs(1242));
    layer5_outputs(1230) <= '0';
    layer5_outputs(1231) <= not(layer4_outputs(1665)) or (layer4_outputs(865));
    layer5_outputs(1232) <= not(layer4_outputs(64));
    layer5_outputs(1233) <= (layer4_outputs(295)) and not (layer4_outputs(730));
    layer5_outputs(1234) <= not(layer4_outputs(1760));
    layer5_outputs(1235) <= '0';
    layer5_outputs(1236) <= (layer4_outputs(1473)) and not (layer4_outputs(1429));
    layer5_outputs(1237) <= not(layer4_outputs(2519));
    layer5_outputs(1238) <= layer4_outputs(1102);
    layer5_outputs(1239) <= not(layer4_outputs(55)) or (layer4_outputs(1784));
    layer5_outputs(1240) <= not(layer4_outputs(731));
    layer5_outputs(1241) <= (layer4_outputs(551)) and not (layer4_outputs(547));
    layer5_outputs(1242) <= layer4_outputs(249);
    layer5_outputs(1243) <= layer4_outputs(2391);
    layer5_outputs(1244) <= not(layer4_outputs(2487));
    layer5_outputs(1245) <= layer4_outputs(1876);
    layer5_outputs(1246) <= (layer4_outputs(2538)) and not (layer4_outputs(2005));
    layer5_outputs(1247) <= not(layer4_outputs(1562));
    layer5_outputs(1248) <= not(layer4_outputs(79));
    layer5_outputs(1249) <= (layer4_outputs(125)) and not (layer4_outputs(1316));
    layer5_outputs(1250) <= not(layer4_outputs(1858));
    layer5_outputs(1251) <= layer4_outputs(1777);
    layer5_outputs(1252) <= not(layer4_outputs(542));
    layer5_outputs(1253) <= layer4_outputs(112);
    layer5_outputs(1254) <= (layer4_outputs(1693)) or (layer4_outputs(2158));
    layer5_outputs(1255) <= not(layer4_outputs(1406));
    layer5_outputs(1256) <= (layer4_outputs(1272)) or (layer4_outputs(1776));
    layer5_outputs(1257) <= (layer4_outputs(2148)) and not (layer4_outputs(1870));
    layer5_outputs(1258) <= layer4_outputs(583);
    layer5_outputs(1259) <= not((layer4_outputs(310)) or (layer4_outputs(1538)));
    layer5_outputs(1260) <= not((layer4_outputs(2121)) or (layer4_outputs(1892)));
    layer5_outputs(1261) <= layer4_outputs(1938);
    layer5_outputs(1262) <= (layer4_outputs(605)) or (layer4_outputs(2424));
    layer5_outputs(1263) <= not(layer4_outputs(340));
    layer5_outputs(1264) <= (layer4_outputs(2168)) and not (layer4_outputs(553));
    layer5_outputs(1265) <= not(layer4_outputs(1752));
    layer5_outputs(1266) <= (layer4_outputs(1867)) and not (layer4_outputs(399));
    layer5_outputs(1267) <= not(layer4_outputs(1997)) or (layer4_outputs(130));
    layer5_outputs(1268) <= not((layer4_outputs(1040)) xor (layer4_outputs(2201)));
    layer5_outputs(1269) <= not(layer4_outputs(1367)) or (layer4_outputs(1307));
    layer5_outputs(1270) <= not(layer4_outputs(1493));
    layer5_outputs(1271) <= layer4_outputs(1273);
    layer5_outputs(1272) <= (layer4_outputs(29)) and (layer4_outputs(303));
    layer5_outputs(1273) <= layer4_outputs(190);
    layer5_outputs(1274) <= not(layer4_outputs(1017));
    layer5_outputs(1275) <= '0';
    layer5_outputs(1276) <= not((layer4_outputs(222)) and (layer4_outputs(1878)));
    layer5_outputs(1277) <= layer4_outputs(606);
    layer5_outputs(1278) <= '1';
    layer5_outputs(1279) <= not((layer4_outputs(1411)) and (layer4_outputs(1121)));
    layer5_outputs(1280) <= not((layer4_outputs(1782)) and (layer4_outputs(1046)));
    layer5_outputs(1281) <= not(layer4_outputs(412));
    layer5_outputs(1282) <= not((layer4_outputs(1238)) and (layer4_outputs(1973)));
    layer5_outputs(1283) <= not(layer4_outputs(1964));
    layer5_outputs(1284) <= '1';
    layer5_outputs(1285) <= layer4_outputs(1216);
    layer5_outputs(1286) <= (layer4_outputs(2193)) and (layer4_outputs(1313));
    layer5_outputs(1287) <= not(layer4_outputs(2103));
    layer5_outputs(1288) <= not(layer4_outputs(786));
    layer5_outputs(1289) <= not(layer4_outputs(14));
    layer5_outputs(1290) <= not(layer4_outputs(2416)) or (layer4_outputs(750));
    layer5_outputs(1291) <= not(layer4_outputs(2399));
    layer5_outputs(1292) <= not((layer4_outputs(357)) xor (layer4_outputs(1849)));
    layer5_outputs(1293) <= (layer4_outputs(826)) and not (layer4_outputs(2349));
    layer5_outputs(1294) <= not((layer4_outputs(934)) xor (layer4_outputs(929)));
    layer5_outputs(1295) <= not(layer4_outputs(788));
    layer5_outputs(1296) <= not(layer4_outputs(1693));
    layer5_outputs(1297) <= not((layer4_outputs(986)) xor (layer4_outputs(1341)));
    layer5_outputs(1298) <= layer4_outputs(2391);
    layer5_outputs(1299) <= not((layer4_outputs(1769)) xor (layer4_outputs(772)));
    layer5_outputs(1300) <= layer4_outputs(2247);
    layer5_outputs(1301) <= not(layer4_outputs(291));
    layer5_outputs(1302) <= layer4_outputs(1440);
    layer5_outputs(1303) <= not((layer4_outputs(711)) or (layer4_outputs(1575)));
    layer5_outputs(1304) <= layer4_outputs(295);
    layer5_outputs(1305) <= not((layer4_outputs(1752)) and (layer4_outputs(1775)));
    layer5_outputs(1306) <= layer4_outputs(2477);
    layer5_outputs(1307) <= layer4_outputs(421);
    layer5_outputs(1308) <= (layer4_outputs(2361)) and (layer4_outputs(376));
    layer5_outputs(1309) <= layer4_outputs(1661);
    layer5_outputs(1310) <= layer4_outputs(2111);
    layer5_outputs(1311) <= not((layer4_outputs(1091)) or (layer4_outputs(2043)));
    layer5_outputs(1312) <= not(layer4_outputs(1475));
    layer5_outputs(1313) <= not(layer4_outputs(575));
    layer5_outputs(1314) <= (layer4_outputs(1986)) and (layer4_outputs(2262));
    layer5_outputs(1315) <= not(layer4_outputs(832)) or (layer4_outputs(73));
    layer5_outputs(1316) <= not((layer4_outputs(428)) xor (layer4_outputs(317)));
    layer5_outputs(1317) <= layer4_outputs(2201);
    layer5_outputs(1318) <= not(layer4_outputs(2098)) or (layer4_outputs(2253));
    layer5_outputs(1319) <= layer4_outputs(2339);
    layer5_outputs(1320) <= not((layer4_outputs(2141)) and (layer4_outputs(1437)));
    layer5_outputs(1321) <= '0';
    layer5_outputs(1322) <= not(layer4_outputs(1850)) or (layer4_outputs(1716));
    layer5_outputs(1323) <= not((layer4_outputs(1884)) and (layer4_outputs(2043)));
    layer5_outputs(1324) <= not(layer4_outputs(1092));
    layer5_outputs(1325) <= (layer4_outputs(232)) and not (layer4_outputs(2092));
    layer5_outputs(1326) <= (layer4_outputs(1389)) or (layer4_outputs(1772));
    layer5_outputs(1327) <= not(layer4_outputs(1449)) or (layer4_outputs(1159));
    layer5_outputs(1328) <= not(layer4_outputs(1301));
    layer5_outputs(1329) <= not((layer4_outputs(529)) xor (layer4_outputs(718)));
    layer5_outputs(1330) <= layer4_outputs(2468);
    layer5_outputs(1331) <= not(layer4_outputs(171));
    layer5_outputs(1332) <= not(layer4_outputs(2042)) or (layer4_outputs(1399));
    layer5_outputs(1333) <= (layer4_outputs(1946)) or (layer4_outputs(1093));
    layer5_outputs(1334) <= not(layer4_outputs(1921)) or (layer4_outputs(1419));
    layer5_outputs(1335) <= (layer4_outputs(173)) and not (layer4_outputs(597));
    layer5_outputs(1336) <= '0';
    layer5_outputs(1337) <= not(layer4_outputs(1356)) or (layer4_outputs(904));
    layer5_outputs(1338) <= layer4_outputs(787);
    layer5_outputs(1339) <= not(layer4_outputs(2225)) or (layer4_outputs(518));
    layer5_outputs(1340) <= '1';
    layer5_outputs(1341) <= not(layer4_outputs(330)) or (layer4_outputs(1755));
    layer5_outputs(1342) <= layer4_outputs(1986);
    layer5_outputs(1343) <= (layer4_outputs(878)) and (layer4_outputs(894));
    layer5_outputs(1344) <= not(layer4_outputs(1043));
    layer5_outputs(1345) <= not(layer4_outputs(2063)) or (layer4_outputs(1961));
    layer5_outputs(1346) <= not(layer4_outputs(1085));
    layer5_outputs(1347) <= not((layer4_outputs(2381)) and (layer4_outputs(657)));
    layer5_outputs(1348) <= not(layer4_outputs(419));
    layer5_outputs(1349) <= not(layer4_outputs(910));
    layer5_outputs(1350) <= layer4_outputs(1632);
    layer5_outputs(1351) <= not(layer4_outputs(2245));
    layer5_outputs(1352) <= '0';
    layer5_outputs(1353) <= (layer4_outputs(801)) or (layer4_outputs(2051));
    layer5_outputs(1354) <= (layer4_outputs(1238)) xor (layer4_outputs(1584));
    layer5_outputs(1355) <= layer4_outputs(2230);
    layer5_outputs(1356) <= not((layer4_outputs(833)) xor (layer4_outputs(2190)));
    layer5_outputs(1357) <= layer4_outputs(346);
    layer5_outputs(1358) <= layer4_outputs(1851);
    layer5_outputs(1359) <= layer4_outputs(614);
    layer5_outputs(1360) <= not((layer4_outputs(470)) xor (layer4_outputs(814)));
    layer5_outputs(1361) <= not((layer4_outputs(1641)) and (layer4_outputs(154)));
    layer5_outputs(1362) <= '1';
    layer5_outputs(1363) <= not(layer4_outputs(1626)) or (layer4_outputs(2153));
    layer5_outputs(1364) <= not(layer4_outputs(2331));
    layer5_outputs(1365) <= not(layer4_outputs(681)) or (layer4_outputs(768));
    layer5_outputs(1366) <= not((layer4_outputs(1023)) and (layer4_outputs(1942)));
    layer5_outputs(1367) <= not(layer4_outputs(1817));
    layer5_outputs(1368) <= not(layer4_outputs(2513));
    layer5_outputs(1369) <= not(layer4_outputs(2321));
    layer5_outputs(1370) <= '0';
    layer5_outputs(1371) <= layer4_outputs(2173);
    layer5_outputs(1372) <= (layer4_outputs(1610)) or (layer4_outputs(2449));
    layer5_outputs(1373) <= layer4_outputs(568);
    layer5_outputs(1374) <= (layer4_outputs(414)) xor (layer4_outputs(2256));
    layer5_outputs(1375) <= layer4_outputs(1623);
    layer5_outputs(1376) <= layer4_outputs(471);
    layer5_outputs(1377) <= layer4_outputs(1980);
    layer5_outputs(1378) <= layer4_outputs(1289);
    layer5_outputs(1379) <= not(layer4_outputs(1285)) or (layer4_outputs(1516));
    layer5_outputs(1380) <= (layer4_outputs(1759)) and not (layer4_outputs(138));
    layer5_outputs(1381) <= not((layer4_outputs(1538)) and (layer4_outputs(2390)));
    layer5_outputs(1382) <= (layer4_outputs(1228)) and not (layer4_outputs(1549));
    layer5_outputs(1383) <= not(layer4_outputs(1463)) or (layer4_outputs(124));
    layer5_outputs(1384) <= not(layer4_outputs(891));
    layer5_outputs(1385) <= layer4_outputs(242);
    layer5_outputs(1386) <= (layer4_outputs(1174)) xor (layer4_outputs(290));
    layer5_outputs(1387) <= not(layer4_outputs(1811));
    layer5_outputs(1388) <= (layer4_outputs(1035)) or (layer4_outputs(2351));
    layer5_outputs(1389) <= '0';
    layer5_outputs(1390) <= (layer4_outputs(1097)) or (layer4_outputs(1106));
    layer5_outputs(1391) <= layer4_outputs(736);
    layer5_outputs(1392) <= not(layer4_outputs(2518));
    layer5_outputs(1393) <= not((layer4_outputs(353)) and (layer4_outputs(1910)));
    layer5_outputs(1394) <= not((layer4_outputs(71)) or (layer4_outputs(2290)));
    layer5_outputs(1395) <= not(layer4_outputs(1311));
    layer5_outputs(1396) <= layer4_outputs(560);
    layer5_outputs(1397) <= (layer4_outputs(2183)) and (layer4_outputs(2358));
    layer5_outputs(1398) <= (layer4_outputs(373)) and not (layer4_outputs(846));
    layer5_outputs(1399) <= layer4_outputs(2325);
    layer5_outputs(1400) <= not(layer4_outputs(2525));
    layer5_outputs(1401) <= (layer4_outputs(548)) and (layer4_outputs(639));
    layer5_outputs(1402) <= (layer4_outputs(270)) and not (layer4_outputs(520));
    layer5_outputs(1403) <= layer4_outputs(1256);
    layer5_outputs(1404) <= not((layer4_outputs(2340)) or (layer4_outputs(1338)));
    layer5_outputs(1405) <= layer4_outputs(2319);
    layer5_outputs(1406) <= not((layer4_outputs(1968)) and (layer4_outputs(2293)));
    layer5_outputs(1407) <= layer4_outputs(1766);
    layer5_outputs(1408) <= not(layer4_outputs(1662));
    layer5_outputs(1409) <= not((layer4_outputs(408)) or (layer4_outputs(192)));
    layer5_outputs(1410) <= not(layer4_outputs(160));
    layer5_outputs(1411) <= layer4_outputs(1899);
    layer5_outputs(1412) <= (layer4_outputs(170)) and (layer4_outputs(2512));
    layer5_outputs(1413) <= layer4_outputs(2035);
    layer5_outputs(1414) <= not(layer4_outputs(497));
    layer5_outputs(1415) <= not(layer4_outputs(142)) or (layer4_outputs(1701));
    layer5_outputs(1416) <= not(layer4_outputs(1147)) or (layer4_outputs(500));
    layer5_outputs(1417) <= not(layer4_outputs(1380));
    layer5_outputs(1418) <= not(layer4_outputs(999));
    layer5_outputs(1419) <= layer4_outputs(1865);
    layer5_outputs(1420) <= (layer4_outputs(39)) and not (layer4_outputs(1642));
    layer5_outputs(1421) <= layer4_outputs(1489);
    layer5_outputs(1422) <= not((layer4_outputs(63)) or (layer4_outputs(764)));
    layer5_outputs(1423) <= not(layer4_outputs(1745)) or (layer4_outputs(2395));
    layer5_outputs(1424) <= layer4_outputs(1840);
    layer5_outputs(1425) <= not(layer4_outputs(61));
    layer5_outputs(1426) <= (layer4_outputs(2340)) and (layer4_outputs(93));
    layer5_outputs(1427) <= layer4_outputs(2081);
    layer5_outputs(1428) <= '1';
    layer5_outputs(1429) <= layer4_outputs(1378);
    layer5_outputs(1430) <= layer4_outputs(2426);
    layer5_outputs(1431) <= (layer4_outputs(244)) and not (layer4_outputs(2164));
    layer5_outputs(1432) <= not(layer4_outputs(89));
    layer5_outputs(1433) <= layer4_outputs(822);
    layer5_outputs(1434) <= layer4_outputs(867);
    layer5_outputs(1435) <= layer4_outputs(254);
    layer5_outputs(1436) <= layer4_outputs(2453);
    layer5_outputs(1437) <= not(layer4_outputs(568));
    layer5_outputs(1438) <= not(layer4_outputs(1275));
    layer5_outputs(1439) <= (layer4_outputs(1405)) and (layer4_outputs(2423));
    layer5_outputs(1440) <= (layer4_outputs(2531)) xor (layer4_outputs(2398));
    layer5_outputs(1441) <= (layer4_outputs(453)) and not (layer4_outputs(2249));
    layer5_outputs(1442) <= not((layer4_outputs(1526)) and (layer4_outputs(1519)));
    layer5_outputs(1443) <= layer4_outputs(720);
    layer5_outputs(1444) <= not((layer4_outputs(52)) and (layer4_outputs(2145)));
    layer5_outputs(1445) <= layer4_outputs(2559);
    layer5_outputs(1446) <= not((layer4_outputs(1155)) or (layer4_outputs(1033)));
    layer5_outputs(1447) <= not(layer4_outputs(487));
    layer5_outputs(1448) <= not(layer4_outputs(527));
    layer5_outputs(1449) <= (layer4_outputs(200)) and not (layer4_outputs(1914));
    layer5_outputs(1450) <= layer4_outputs(131);
    layer5_outputs(1451) <= layer4_outputs(1458);
    layer5_outputs(1452) <= not((layer4_outputs(2458)) or (layer4_outputs(19)));
    layer5_outputs(1453) <= not(layer4_outputs(448));
    layer5_outputs(1454) <= not(layer4_outputs(2110));
    layer5_outputs(1455) <= '0';
    layer5_outputs(1456) <= not((layer4_outputs(798)) xor (layer4_outputs(2298)));
    layer5_outputs(1457) <= (layer4_outputs(958)) or (layer4_outputs(1990));
    layer5_outputs(1458) <= not((layer4_outputs(2337)) or (layer4_outputs(2130)));
    layer5_outputs(1459) <= not(layer4_outputs(80));
    layer5_outputs(1460) <= (layer4_outputs(1758)) and (layer4_outputs(1198));
    layer5_outputs(1461) <= not((layer4_outputs(1565)) and (layer4_outputs(2336)));
    layer5_outputs(1462) <= not(layer4_outputs(1072));
    layer5_outputs(1463) <= not(layer4_outputs(202)) or (layer4_outputs(362));
    layer5_outputs(1464) <= (layer4_outputs(1049)) and not (layer4_outputs(415));
    layer5_outputs(1465) <= layer4_outputs(1711);
    layer5_outputs(1466) <= not(layer4_outputs(2044));
    layer5_outputs(1467) <= not(layer4_outputs(807));
    layer5_outputs(1468) <= not(layer4_outputs(1753)) or (layer4_outputs(1304));
    layer5_outputs(1469) <= not(layer4_outputs(967));
    layer5_outputs(1470) <= not((layer4_outputs(1695)) xor (layer4_outputs(1137)));
    layer5_outputs(1471) <= not(layer4_outputs(1687));
    layer5_outputs(1472) <= not(layer4_outputs(813));
    layer5_outputs(1473) <= layer4_outputs(1659);
    layer5_outputs(1474) <= (layer4_outputs(329)) and (layer4_outputs(1119));
    layer5_outputs(1475) <= not((layer4_outputs(1146)) xor (layer4_outputs(83)));
    layer5_outputs(1476) <= not(layer4_outputs(2450));
    layer5_outputs(1477) <= layer4_outputs(2402);
    layer5_outputs(1478) <= layer4_outputs(561);
    layer5_outputs(1479) <= layer4_outputs(771);
    layer5_outputs(1480) <= not((layer4_outputs(1197)) or (layer4_outputs(2)));
    layer5_outputs(1481) <= (layer4_outputs(1945)) and (layer4_outputs(1132));
    layer5_outputs(1482) <= layer4_outputs(705);
    layer5_outputs(1483) <= not(layer4_outputs(1058));
    layer5_outputs(1484) <= layer4_outputs(668);
    layer5_outputs(1485) <= not((layer4_outputs(762)) xor (layer4_outputs(770)));
    layer5_outputs(1486) <= not(layer4_outputs(2347)) or (layer4_outputs(2272));
    layer5_outputs(1487) <= layer4_outputs(775);
    layer5_outputs(1488) <= not((layer4_outputs(1290)) or (layer4_outputs(1887)));
    layer5_outputs(1489) <= not(layer4_outputs(2125)) or (layer4_outputs(395));
    layer5_outputs(1490) <= not(layer4_outputs(2190)) or (layer4_outputs(2172));
    layer5_outputs(1491) <= (layer4_outputs(836)) and not (layer4_outputs(741));
    layer5_outputs(1492) <= layer4_outputs(246);
    layer5_outputs(1493) <= '0';
    layer5_outputs(1494) <= not((layer4_outputs(342)) xor (layer4_outputs(1567)));
    layer5_outputs(1495) <= not(layer4_outputs(1251));
    layer5_outputs(1496) <= '0';
    layer5_outputs(1497) <= not(layer4_outputs(491)) or (layer4_outputs(1098));
    layer5_outputs(1498) <= (layer4_outputs(553)) and (layer4_outputs(2382));
    layer5_outputs(1499) <= '0';
    layer5_outputs(1500) <= not(layer4_outputs(2556));
    layer5_outputs(1501) <= layer4_outputs(328);
    layer5_outputs(1502) <= layer4_outputs(1564);
    layer5_outputs(1503) <= layer4_outputs(1482);
    layer5_outputs(1504) <= (layer4_outputs(1553)) and not (layer4_outputs(259));
    layer5_outputs(1505) <= (layer4_outputs(742)) and (layer4_outputs(316));
    layer5_outputs(1506) <= not(layer4_outputs(350));
    layer5_outputs(1507) <= not(layer4_outputs(1981));
    layer5_outputs(1508) <= not(layer4_outputs(162));
    layer5_outputs(1509) <= layer4_outputs(751);
    layer5_outputs(1510) <= not((layer4_outputs(309)) xor (layer4_outputs(2026)));
    layer5_outputs(1511) <= (layer4_outputs(2249)) and not (layer4_outputs(501));
    layer5_outputs(1512) <= not((layer4_outputs(2261)) or (layer4_outputs(854)));
    layer5_outputs(1513) <= not(layer4_outputs(1706));
    layer5_outputs(1514) <= not(layer4_outputs(1308)) or (layer4_outputs(2313));
    layer5_outputs(1515) <= (layer4_outputs(1450)) xor (layer4_outputs(215));
    layer5_outputs(1516) <= not(layer4_outputs(2437));
    layer5_outputs(1517) <= (layer4_outputs(36)) and (layer4_outputs(507));
    layer5_outputs(1518) <= (layer4_outputs(2239)) xor (layer4_outputs(1390));
    layer5_outputs(1519) <= not(layer4_outputs(1042)) or (layer4_outputs(100));
    layer5_outputs(1520) <= not(layer4_outputs(594));
    layer5_outputs(1521) <= (layer4_outputs(1603)) xor (layer4_outputs(2516));
    layer5_outputs(1522) <= not((layer4_outputs(1178)) and (layer4_outputs(298)));
    layer5_outputs(1523) <= not(layer4_outputs(1552)) or (layer4_outputs(44));
    layer5_outputs(1524) <= not(layer4_outputs(274));
    layer5_outputs(1525) <= (layer4_outputs(1668)) or (layer4_outputs(1160));
    layer5_outputs(1526) <= layer4_outputs(2100);
    layer5_outputs(1527) <= layer4_outputs(2488);
    layer5_outputs(1528) <= not(layer4_outputs(532));
    layer5_outputs(1529) <= (layer4_outputs(1179)) and (layer4_outputs(665));
    layer5_outputs(1530) <= (layer4_outputs(2222)) xor (layer4_outputs(1965));
    layer5_outputs(1531) <= not((layer4_outputs(798)) and (layer4_outputs(371)));
    layer5_outputs(1532) <= layer4_outputs(105);
    layer5_outputs(1533) <= not(layer4_outputs(2060));
    layer5_outputs(1534) <= (layer4_outputs(825)) and not (layer4_outputs(289));
    layer5_outputs(1535) <= (layer4_outputs(1151)) and (layer4_outputs(183));
    layer5_outputs(1536) <= layer4_outputs(538);
    layer5_outputs(1537) <= not(layer4_outputs(1532)) or (layer4_outputs(973));
    layer5_outputs(1538) <= not((layer4_outputs(377)) and (layer4_outputs(785)));
    layer5_outputs(1539) <= '1';
    layer5_outputs(1540) <= layer4_outputs(906);
    layer5_outputs(1541) <= not(layer4_outputs(723));
    layer5_outputs(1542) <= (layer4_outputs(120)) and not (layer4_outputs(1101));
    layer5_outputs(1543) <= layer4_outputs(1871);
    layer5_outputs(1544) <= not(layer4_outputs(277)) or (layer4_outputs(1242));
    layer5_outputs(1545) <= not(layer4_outputs(1731));
    layer5_outputs(1546) <= not((layer4_outputs(410)) xor (layer4_outputs(1677)));
    layer5_outputs(1547) <= not(layer4_outputs(1324));
    layer5_outputs(1548) <= (layer4_outputs(400)) or (layer4_outputs(1077));
    layer5_outputs(1549) <= not((layer4_outputs(9)) or (layer4_outputs(1615)));
    layer5_outputs(1550) <= (layer4_outputs(2037)) and not (layer4_outputs(2499));
    layer5_outputs(1551) <= not(layer4_outputs(1315));
    layer5_outputs(1552) <= not((layer4_outputs(919)) and (layer4_outputs(306)));
    layer5_outputs(1553) <= not(layer4_outputs(339));
    layer5_outputs(1554) <= not(layer4_outputs(821));
    layer5_outputs(1555) <= (layer4_outputs(1673)) or (layer4_outputs(1977));
    layer5_outputs(1556) <= layer4_outputs(1257);
    layer5_outputs(1557) <= not(layer4_outputs(1604));
    layer5_outputs(1558) <= (layer4_outputs(1447)) and not (layer4_outputs(401));
    layer5_outputs(1559) <= not((layer4_outputs(2485)) xor (layer4_outputs(1587)));
    layer5_outputs(1560) <= '1';
    layer5_outputs(1561) <= layer4_outputs(899);
    layer5_outputs(1562) <= (layer4_outputs(1438)) or (layer4_outputs(2310));
    layer5_outputs(1563) <= not(layer4_outputs(1131));
    layer5_outputs(1564) <= not(layer4_outputs(234));
    layer5_outputs(1565) <= layer4_outputs(671);
    layer5_outputs(1566) <= (layer4_outputs(799)) xor (layer4_outputs(188));
    layer5_outputs(1567) <= not(layer4_outputs(1336));
    layer5_outputs(1568) <= layer4_outputs(135);
    layer5_outputs(1569) <= '1';
    layer5_outputs(1570) <= not(layer4_outputs(1560)) or (layer4_outputs(940));
    layer5_outputs(1571) <= (layer4_outputs(1648)) and not (layer4_outputs(493));
    layer5_outputs(1572) <= not((layer4_outputs(1310)) xor (layer4_outputs(831)));
    layer5_outputs(1573) <= not(layer4_outputs(121));
    layer5_outputs(1574) <= (layer4_outputs(147)) xor (layer4_outputs(1901));
    layer5_outputs(1575) <= not(layer4_outputs(767));
    layer5_outputs(1576) <= (layer4_outputs(2332)) xor (layer4_outputs(1757));
    layer5_outputs(1577) <= not(layer4_outputs(2147));
    layer5_outputs(1578) <= (layer4_outputs(2083)) xor (layer4_outputs(1477));
    layer5_outputs(1579) <= not((layer4_outputs(778)) or (layer4_outputs(617)));
    layer5_outputs(1580) <= layer4_outputs(1206);
    layer5_outputs(1581) <= (layer4_outputs(1496)) and not (layer4_outputs(813));
    layer5_outputs(1582) <= layer4_outputs(1832);
    layer5_outputs(1583) <= layer4_outputs(1267);
    layer5_outputs(1584) <= (layer4_outputs(1305)) and not (layer4_outputs(147));
    layer5_outputs(1585) <= not((layer4_outputs(309)) and (layer4_outputs(2361)));
    layer5_outputs(1586) <= layer4_outputs(674);
    layer5_outputs(1587) <= not(layer4_outputs(626));
    layer5_outputs(1588) <= (layer4_outputs(1334)) and (layer4_outputs(991));
    layer5_outputs(1589) <= not(layer4_outputs(2496));
    layer5_outputs(1590) <= not(layer4_outputs(1881));
    layer5_outputs(1591) <= not(layer4_outputs(1434));
    layer5_outputs(1592) <= not(layer4_outputs(2246));
    layer5_outputs(1593) <= (layer4_outputs(1874)) and not (layer4_outputs(2315));
    layer5_outputs(1594) <= (layer4_outputs(839)) or (layer4_outputs(1152));
    layer5_outputs(1595) <= not((layer4_outputs(1170)) or (layer4_outputs(505)));
    layer5_outputs(1596) <= layer4_outputs(2077);
    layer5_outputs(1597) <= (layer4_outputs(620)) and (layer4_outputs(2372));
    layer5_outputs(1598) <= layer4_outputs(643);
    layer5_outputs(1599) <= not((layer4_outputs(1196)) or (layer4_outputs(1671)));
    layer5_outputs(1600) <= not((layer4_outputs(4)) and (layer4_outputs(1682)));
    layer5_outputs(1601) <= layer4_outputs(544);
    layer5_outputs(1602) <= layer4_outputs(11);
    layer5_outputs(1603) <= layer4_outputs(1333);
    layer5_outputs(1604) <= (layer4_outputs(1151)) and not (layer4_outputs(2231));
    layer5_outputs(1605) <= '0';
    layer5_outputs(1606) <= layer4_outputs(61);
    layer5_outputs(1607) <= layer4_outputs(1811);
    layer5_outputs(1608) <= layer4_outputs(111);
    layer5_outputs(1609) <= not((layer4_outputs(494)) or (layer4_outputs(430)));
    layer5_outputs(1610) <= (layer4_outputs(320)) and not (layer4_outputs(1878));
    layer5_outputs(1611) <= (layer4_outputs(1418)) and (layer4_outputs(1283));
    layer5_outputs(1612) <= '1';
    layer5_outputs(1613) <= not((layer4_outputs(479)) and (layer4_outputs(1644)));
    layer5_outputs(1614) <= '0';
    layer5_outputs(1615) <= not((layer4_outputs(1813)) or (layer4_outputs(1304)));
    layer5_outputs(1616) <= layer4_outputs(1205);
    layer5_outputs(1617) <= layer4_outputs(2064);
    layer5_outputs(1618) <= layer4_outputs(1937);
    layer5_outputs(1619) <= not((layer4_outputs(98)) or (layer4_outputs(2475)));
    layer5_outputs(1620) <= layer4_outputs(2316);
    layer5_outputs(1621) <= not(layer4_outputs(912)) or (layer4_outputs(1004));
    layer5_outputs(1622) <= (layer4_outputs(227)) and not (layer4_outputs(1790));
    layer5_outputs(1623) <= layer4_outputs(409);
    layer5_outputs(1624) <= layer4_outputs(1293);
    layer5_outputs(1625) <= not(layer4_outputs(1190)) or (layer4_outputs(389));
    layer5_outputs(1626) <= not(layer4_outputs(1588));
    layer5_outputs(1627) <= not(layer4_outputs(1363)) or (layer4_outputs(140));
    layer5_outputs(1628) <= not(layer4_outputs(208));
    layer5_outputs(1629) <= not(layer4_outputs(2437));
    layer5_outputs(1630) <= not((layer4_outputs(1917)) or (layer4_outputs(2177)));
    layer5_outputs(1631) <= not(layer4_outputs(2525));
    layer5_outputs(1632) <= not((layer4_outputs(1233)) and (layer4_outputs(920)));
    layer5_outputs(1633) <= (layer4_outputs(1001)) and (layer4_outputs(694));
    layer5_outputs(1634) <= not((layer4_outputs(1920)) or (layer4_outputs(1528)));
    layer5_outputs(1635) <= layer4_outputs(2039);
    layer5_outputs(1636) <= not(layer4_outputs(845));
    layer5_outputs(1637) <= layer4_outputs(2377);
    layer5_outputs(1638) <= not(layer4_outputs(66));
    layer5_outputs(1639) <= not(layer4_outputs(2356)) or (layer4_outputs(1756));
    layer5_outputs(1640) <= layer4_outputs(593);
    layer5_outputs(1641) <= not((layer4_outputs(930)) xor (layer4_outputs(144)));
    layer5_outputs(1642) <= not(layer4_outputs(1704)) or (layer4_outputs(241));
    layer5_outputs(1643) <= not((layer4_outputs(567)) or (layer4_outputs(2496)));
    layer5_outputs(1644) <= not(layer4_outputs(2293));
    layer5_outputs(1645) <= not(layer4_outputs(1874));
    layer5_outputs(1646) <= layer4_outputs(1802);
    layer5_outputs(1647) <= layer4_outputs(2089);
    layer5_outputs(1648) <= not((layer4_outputs(1027)) xor (layer4_outputs(890)));
    layer5_outputs(1649) <= not((layer4_outputs(840)) and (layer4_outputs(1294)));
    layer5_outputs(1650) <= (layer4_outputs(2517)) xor (layer4_outputs(876));
    layer5_outputs(1651) <= (layer4_outputs(964)) and not (layer4_outputs(1580));
    layer5_outputs(1652) <= layer4_outputs(461);
    layer5_outputs(1653) <= layer4_outputs(402);
    layer5_outputs(1654) <= '1';
    layer5_outputs(1655) <= not(layer4_outputs(815));
    layer5_outputs(1656) <= layer4_outputs(1047);
    layer5_outputs(1657) <= layer4_outputs(1169);
    layer5_outputs(1658) <= layer4_outputs(517);
    layer5_outputs(1659) <= '1';
    layer5_outputs(1660) <= layer4_outputs(2189);
    layer5_outputs(1661) <= (layer4_outputs(505)) and (layer4_outputs(2433));
    layer5_outputs(1662) <= (layer4_outputs(1542)) xor (layer4_outputs(1660));
    layer5_outputs(1663) <= layer4_outputs(1868);
    layer5_outputs(1664) <= layer4_outputs(2271);
    layer5_outputs(1665) <= (layer4_outputs(238)) and not (layer4_outputs(1369));
    layer5_outputs(1666) <= layer4_outputs(1383);
    layer5_outputs(1667) <= layer4_outputs(158);
    layer5_outputs(1668) <= layer4_outputs(817);
    layer5_outputs(1669) <= (layer4_outputs(1628)) xor (layer4_outputs(1002));
    layer5_outputs(1670) <= (layer4_outputs(165)) and (layer4_outputs(1669));
    layer5_outputs(1671) <= not(layer4_outputs(2487));
    layer5_outputs(1672) <= (layer4_outputs(2196)) and not (layer4_outputs(1639));
    layer5_outputs(1673) <= not((layer4_outputs(1597)) or (layer4_outputs(941)));
    layer5_outputs(1674) <= layer4_outputs(2355);
    layer5_outputs(1675) <= not((layer4_outputs(9)) or (layer4_outputs(1008)));
    layer5_outputs(1676) <= layer4_outputs(482);
    layer5_outputs(1677) <= not((layer4_outputs(2059)) xor (layer4_outputs(489)));
    layer5_outputs(1678) <= not(layer4_outputs(1167));
    layer5_outputs(1679) <= layer4_outputs(2120);
    layer5_outputs(1680) <= not((layer4_outputs(161)) xor (layer4_outputs(1087)));
    layer5_outputs(1681) <= (layer4_outputs(1554)) and (layer4_outputs(367));
    layer5_outputs(1682) <= layer4_outputs(2218);
    layer5_outputs(1683) <= not(layer4_outputs(1819));
    layer5_outputs(1684) <= (layer4_outputs(1930)) and not (layer4_outputs(686));
    layer5_outputs(1685) <= not(layer4_outputs(1185));
    layer5_outputs(1686) <= not((layer4_outputs(620)) and (layer4_outputs(689)));
    layer5_outputs(1687) <= layer4_outputs(2128);
    layer5_outputs(1688) <= layer4_outputs(2009);
    layer5_outputs(1689) <= not((layer4_outputs(502)) or (layer4_outputs(2428)));
    layer5_outputs(1690) <= not(layer4_outputs(1562));
    layer5_outputs(1691) <= (layer4_outputs(1272)) or (layer4_outputs(2023));
    layer5_outputs(1692) <= (layer4_outputs(2086)) or (layer4_outputs(1144));
    layer5_outputs(1693) <= not(layer4_outputs(726));
    layer5_outputs(1694) <= not(layer4_outputs(1346)) or (layer4_outputs(2451));
    layer5_outputs(1695) <= (layer4_outputs(2040)) and not (layer4_outputs(229));
    layer5_outputs(1696) <= (layer4_outputs(1127)) and (layer4_outputs(827));
    layer5_outputs(1697) <= not(layer4_outputs(1779)) or (layer4_outputs(1673));
    layer5_outputs(1698) <= (layer4_outputs(2464)) xor (layer4_outputs(1522));
    layer5_outputs(1699) <= not((layer4_outputs(670)) xor (layer4_outputs(1332)));
    layer5_outputs(1700) <= layer4_outputs(1827);
    layer5_outputs(1701) <= not((layer4_outputs(1124)) or (layer4_outputs(2538)));
    layer5_outputs(1702) <= not(layer4_outputs(453));
    layer5_outputs(1703) <= not((layer4_outputs(126)) or (layer4_outputs(1559)));
    layer5_outputs(1704) <= (layer4_outputs(965)) and not (layer4_outputs(254));
    layer5_outputs(1705) <= not(layer4_outputs(1748)) or (layer4_outputs(1564));
    layer5_outputs(1706) <= layer4_outputs(2057);
    layer5_outputs(1707) <= layer4_outputs(1485);
    layer5_outputs(1708) <= '1';
    layer5_outputs(1709) <= not(layer4_outputs(1527));
    layer5_outputs(1710) <= not(layer4_outputs(297));
    layer5_outputs(1711) <= not((layer4_outputs(2441)) xor (layer4_outputs(1724)));
    layer5_outputs(1712) <= layer4_outputs(1413);
    layer5_outputs(1713) <= layer4_outputs(872);
    layer5_outputs(1714) <= not((layer4_outputs(437)) xor (layer4_outputs(914)));
    layer5_outputs(1715) <= not(layer4_outputs(1003));
    layer5_outputs(1716) <= not(layer4_outputs(1306));
    layer5_outputs(1717) <= (layer4_outputs(1357)) and (layer4_outputs(1767));
    layer5_outputs(1718) <= not((layer4_outputs(2155)) and (layer4_outputs(1366)));
    layer5_outputs(1719) <= layer4_outputs(478);
    layer5_outputs(1720) <= (layer4_outputs(2087)) and not (layer4_outputs(1690));
    layer5_outputs(1721) <= layer4_outputs(44);
    layer5_outputs(1722) <= not((layer4_outputs(1274)) and (layer4_outputs(2489)));
    layer5_outputs(1723) <= (layer4_outputs(1540)) and not (layer4_outputs(1547));
    layer5_outputs(1724) <= not(layer4_outputs(148));
    layer5_outputs(1725) <= not(layer4_outputs(290));
    layer5_outputs(1726) <= not(layer4_outputs(2458));
    layer5_outputs(1727) <= (layer4_outputs(606)) and not (layer4_outputs(2467));
    layer5_outputs(1728) <= '0';
    layer5_outputs(1729) <= (layer4_outputs(2550)) and not (layer4_outputs(95));
    layer5_outputs(1730) <= (layer4_outputs(1524)) or (layer4_outputs(1199));
    layer5_outputs(1731) <= not(layer4_outputs(1932));
    layer5_outputs(1732) <= not(layer4_outputs(1637));
    layer5_outputs(1733) <= not((layer4_outputs(2344)) xor (layer4_outputs(226)));
    layer5_outputs(1734) <= not(layer4_outputs(724));
    layer5_outputs(1735) <= (layer4_outputs(1129)) xor (layer4_outputs(1012));
    layer5_outputs(1736) <= not(layer4_outputs(1519)) or (layer4_outputs(849));
    layer5_outputs(1737) <= not(layer4_outputs(396)) or (layer4_outputs(1410));
    layer5_outputs(1738) <= not((layer4_outputs(1137)) or (layer4_outputs(1472)));
    layer5_outputs(1739) <= not(layer4_outputs(1362));
    layer5_outputs(1740) <= not(layer4_outputs(1804));
    layer5_outputs(1741) <= (layer4_outputs(333)) xor (layer4_outputs(199));
    layer5_outputs(1742) <= layer4_outputs(582);
    layer5_outputs(1743) <= not(layer4_outputs(477));
    layer5_outputs(1744) <= not(layer4_outputs(512));
    layer5_outputs(1745) <= not((layer4_outputs(67)) xor (layer4_outputs(1193)));
    layer5_outputs(1746) <= layer4_outputs(1814);
    layer5_outputs(1747) <= not((layer4_outputs(2126)) xor (layer4_outputs(1595)));
    layer5_outputs(1748) <= (layer4_outputs(981)) and not (layer4_outputs(1999));
    layer5_outputs(1749) <= not(layer4_outputs(2116));
    layer5_outputs(1750) <= layer4_outputs(127);
    layer5_outputs(1751) <= layer4_outputs(271);
    layer5_outputs(1752) <= (layer4_outputs(1498)) xor (layer4_outputs(1573));
    layer5_outputs(1753) <= not(layer4_outputs(1062));
    layer5_outputs(1754) <= not((layer4_outputs(823)) and (layer4_outputs(997)));
    layer5_outputs(1755) <= layer4_outputs(2392);
    layer5_outputs(1756) <= not((layer4_outputs(1550)) and (layer4_outputs(1013)));
    layer5_outputs(1757) <= not(layer4_outputs(2559));
    layer5_outputs(1758) <= not((layer4_outputs(2018)) xor (layer4_outputs(156)));
    layer5_outputs(1759) <= not(layer4_outputs(1694));
    layer5_outputs(1760) <= layer4_outputs(180);
    layer5_outputs(1761) <= '0';
    layer5_outputs(1762) <= '0';
    layer5_outputs(1763) <= not((layer4_outputs(779)) or (layer4_outputs(149)));
    layer5_outputs(1764) <= not(layer4_outputs(1028));
    layer5_outputs(1765) <= not(layer4_outputs(2479));
    layer5_outputs(1766) <= (layer4_outputs(1987)) and not (layer4_outputs(2469));
    layer5_outputs(1767) <= not(layer4_outputs(2036)) or (layer4_outputs(1915));
    layer5_outputs(1768) <= not((layer4_outputs(1795)) and (layer4_outputs(1963)));
    layer5_outputs(1769) <= (layer4_outputs(962)) and not (layer4_outputs(2295));
    layer5_outputs(1770) <= not(layer4_outputs(369));
    layer5_outputs(1771) <= not(layer4_outputs(108));
    layer5_outputs(1772) <= not((layer4_outputs(2028)) xor (layer4_outputs(564)));
    layer5_outputs(1773) <= '0';
    layer5_outputs(1774) <= not(layer4_outputs(519));
    layer5_outputs(1775) <= (layer4_outputs(2179)) or (layer4_outputs(2214));
    layer5_outputs(1776) <= not(layer4_outputs(1081));
    layer5_outputs(1777) <= not(layer4_outputs(248));
    layer5_outputs(1778) <= layer4_outputs(1689);
    layer5_outputs(1779) <= layer4_outputs(2300);
    layer5_outputs(1780) <= not((layer4_outputs(1743)) and (layer4_outputs(898)));
    layer5_outputs(1781) <= (layer4_outputs(837)) or (layer4_outputs(1432));
    layer5_outputs(1782) <= layer4_outputs(1214);
    layer5_outputs(1783) <= layer4_outputs(2494);
    layer5_outputs(1784) <= '0';
    layer5_outputs(1785) <= not(layer4_outputs(2105));
    layer5_outputs(1786) <= '1';
    layer5_outputs(1787) <= (layer4_outputs(1107)) xor (layer4_outputs(702));
    layer5_outputs(1788) <= not(layer4_outputs(2503));
    layer5_outputs(1789) <= layer4_outputs(2364);
    layer5_outputs(1790) <= not(layer4_outputs(1103)) or (layer4_outputs(1166));
    layer5_outputs(1791) <= not(layer4_outputs(1984)) or (layer4_outputs(107));
    layer5_outputs(1792) <= not((layer4_outputs(2452)) or (layer4_outputs(2104)));
    layer5_outputs(1793) <= (layer4_outputs(852)) and (layer4_outputs(435));
    layer5_outputs(1794) <= layer4_outputs(187);
    layer5_outputs(1795) <= (layer4_outputs(1062)) and not (layer4_outputs(441));
    layer5_outputs(1796) <= layer4_outputs(1988);
    layer5_outputs(1797) <= (layer4_outputs(101)) and (layer4_outputs(905));
    layer5_outputs(1798) <= (layer4_outputs(2447)) xor (layer4_outputs(2119));
    layer5_outputs(1799) <= (layer4_outputs(1154)) xor (layer4_outputs(1948));
    layer5_outputs(1800) <= not((layer4_outputs(2362)) or (layer4_outputs(1268)));
    layer5_outputs(1801) <= layer4_outputs(2221);
    layer5_outputs(1802) <= not(layer4_outputs(1606));
    layer5_outputs(1803) <= not(layer4_outputs(1106));
    layer5_outputs(1804) <= not((layer4_outputs(638)) xor (layer4_outputs(428)));
    layer5_outputs(1805) <= not(layer4_outputs(1585));
    layer5_outputs(1806) <= not((layer4_outputs(2159)) xor (layer4_outputs(1742)));
    layer5_outputs(1807) <= layer4_outputs(2527);
    layer5_outputs(1808) <= (layer4_outputs(1046)) and (layer4_outputs(1771));
    layer5_outputs(1809) <= layer4_outputs(2122);
    layer5_outputs(1810) <= not(layer4_outputs(645));
    layer5_outputs(1811) <= (layer4_outputs(1969)) or (layer4_outputs(2198));
    layer5_outputs(1812) <= not(layer4_outputs(47));
    layer5_outputs(1813) <= layer4_outputs(908);
    layer5_outputs(1814) <= (layer4_outputs(929)) or (layer4_outputs(163));
    layer5_outputs(1815) <= not(layer4_outputs(356)) or (layer4_outputs(2171));
    layer5_outputs(1816) <= not(layer4_outputs(1019));
    layer5_outputs(1817) <= (layer4_outputs(1213)) and not (layer4_outputs(1507));
    layer5_outputs(1818) <= not(layer4_outputs(1602));
    layer5_outputs(1819) <= not(layer4_outputs(1256));
    layer5_outputs(1820) <= not((layer4_outputs(1778)) and (layer4_outputs(379)));
    layer5_outputs(1821) <= layer4_outputs(99);
    layer5_outputs(1822) <= layer4_outputs(2254);
    layer5_outputs(1823) <= (layer4_outputs(2204)) and not (layer4_outputs(1368));
    layer5_outputs(1824) <= not(layer4_outputs(547));
    layer5_outputs(1825) <= layer4_outputs(2354);
    layer5_outputs(1826) <= layer4_outputs(697);
    layer5_outputs(1827) <= '0';
    layer5_outputs(1828) <= not((layer4_outputs(2003)) and (layer4_outputs(2237)));
    layer5_outputs(1829) <= (layer4_outputs(37)) and not (layer4_outputs(690));
    layer5_outputs(1830) <= not((layer4_outputs(660)) and (layer4_outputs(1937)));
    layer5_outputs(1831) <= (layer4_outputs(1502)) and not (layer4_outputs(1402));
    layer5_outputs(1832) <= layer4_outputs(1933);
    layer5_outputs(1833) <= not((layer4_outputs(539)) xor (layer4_outputs(104)));
    layer5_outputs(1834) <= '1';
    layer5_outputs(1835) <= (layer4_outputs(892)) and not (layer4_outputs(633));
    layer5_outputs(1836) <= not(layer4_outputs(332));
    layer5_outputs(1837) <= not(layer4_outputs(1994));
    layer5_outputs(1838) <= not(layer4_outputs(570));
    layer5_outputs(1839) <= layer4_outputs(2384);
    layer5_outputs(1840) <= not(layer4_outputs(2359));
    layer5_outputs(1841) <= (layer4_outputs(2319)) xor (layer4_outputs(218));
    layer5_outputs(1842) <= (layer4_outputs(1308)) or (layer4_outputs(476));
    layer5_outputs(1843) <= (layer4_outputs(2191)) and (layer4_outputs(2032));
    layer5_outputs(1844) <= not((layer4_outputs(1954)) xor (layer4_outputs(758)));
    layer5_outputs(1845) <= not(layer4_outputs(1118)) or (layer4_outputs(919));
    layer5_outputs(1846) <= (layer4_outputs(2523)) and not (layer4_outputs(699));
    layer5_outputs(1847) <= (layer4_outputs(2264)) and not (layer4_outputs(273));
    layer5_outputs(1848) <= not((layer4_outputs(2491)) and (layer4_outputs(1573)));
    layer5_outputs(1849) <= not(layer4_outputs(1706));
    layer5_outputs(1850) <= not(layer4_outputs(2353));
    layer5_outputs(1851) <= not(layer4_outputs(1520));
    layer5_outputs(1852) <= (layer4_outputs(971)) and not (layer4_outputs(512));
    layer5_outputs(1853) <= (layer4_outputs(1258)) and not (layer4_outputs(381));
    layer5_outputs(1854) <= layer4_outputs(231);
    layer5_outputs(1855) <= (layer4_outputs(2482)) and not (layer4_outputs(1111));
    layer5_outputs(1856) <= not(layer4_outputs(1158));
    layer5_outputs(1857) <= not(layer4_outputs(1699));
    layer5_outputs(1858) <= not((layer4_outputs(600)) and (layer4_outputs(2131)));
    layer5_outputs(1859) <= (layer4_outputs(709)) or (layer4_outputs(1979));
    layer5_outputs(1860) <= not((layer4_outputs(102)) or (layer4_outputs(909)));
    layer5_outputs(1861) <= not(layer4_outputs(1533)) or (layer4_outputs(2369));
    layer5_outputs(1862) <= not(layer4_outputs(2041));
    layer5_outputs(1863) <= (layer4_outputs(363)) and (layer4_outputs(874));
    layer5_outputs(1864) <= (layer4_outputs(1477)) and (layer4_outputs(467));
    layer5_outputs(1865) <= not((layer4_outputs(2313)) xor (layer4_outputs(156)));
    layer5_outputs(1866) <= not(layer4_outputs(447));
    layer5_outputs(1867) <= not(layer4_outputs(1650));
    layer5_outputs(1868) <= (layer4_outputs(1142)) or (layer4_outputs(1338));
    layer5_outputs(1869) <= '0';
    layer5_outputs(1870) <= (layer4_outputs(2424)) or (layer4_outputs(590));
    layer5_outputs(1871) <= (layer4_outputs(1818)) or (layer4_outputs(1154));
    layer5_outputs(1872) <= (layer4_outputs(2377)) and (layer4_outputs(2154));
    layer5_outputs(1873) <= '0';
    layer5_outputs(1874) <= not(layer4_outputs(1247));
    layer5_outputs(1875) <= '0';
    layer5_outputs(1876) <= layer4_outputs(717);
    layer5_outputs(1877) <= not((layer4_outputs(627)) and (layer4_outputs(1709)));
    layer5_outputs(1878) <= (layer4_outputs(2515)) xor (layer4_outputs(1360));
    layer5_outputs(1879) <= not(layer4_outputs(464)) or (layer4_outputs(1393));
    layer5_outputs(1880) <= not(layer4_outputs(563));
    layer5_outputs(1881) <= layer4_outputs(1560);
    layer5_outputs(1882) <= not(layer4_outputs(1556));
    layer5_outputs(1883) <= layer4_outputs(2345);
    layer5_outputs(1884) <= layer4_outputs(1215);
    layer5_outputs(1885) <= layer4_outputs(2158);
    layer5_outputs(1886) <= not(layer4_outputs(2541)) or (layer4_outputs(838));
    layer5_outputs(1887) <= not((layer4_outputs(659)) xor (layer4_outputs(1343)));
    layer5_outputs(1888) <= not(layer4_outputs(2260));
    layer5_outputs(1889) <= not((layer4_outputs(936)) and (layer4_outputs(1250)));
    layer5_outputs(1890) <= (layer4_outputs(1509)) or (layer4_outputs(743));
    layer5_outputs(1891) <= not(layer4_outputs(40)) or (layer4_outputs(1976));
    layer5_outputs(1892) <= not(layer4_outputs(185));
    layer5_outputs(1893) <= not(layer4_outputs(1991));
    layer5_outputs(1894) <= layer4_outputs(550);
    layer5_outputs(1895) <= not(layer4_outputs(1846));
    layer5_outputs(1896) <= layer4_outputs(1802);
    layer5_outputs(1897) <= (layer4_outputs(268)) and not (layer4_outputs(806));
    layer5_outputs(1898) <= not(layer4_outputs(1105));
    layer5_outputs(1899) <= (layer4_outputs(1940)) and (layer4_outputs(621));
    layer5_outputs(1900) <= not(layer4_outputs(205));
    layer5_outputs(1901) <= not((layer4_outputs(2223)) or (layer4_outputs(1126)));
    layer5_outputs(1902) <= layer4_outputs(632);
    layer5_outputs(1903) <= not(layer4_outputs(396)) or (layer4_outputs(731));
    layer5_outputs(1904) <= (layer4_outputs(1018)) xor (layer4_outputs(572));
    layer5_outputs(1905) <= not((layer4_outputs(1698)) and (layer4_outputs(1690)));
    layer5_outputs(1906) <= layer4_outputs(253);
    layer5_outputs(1907) <= (layer4_outputs(248)) or (layer4_outputs(1907));
    layer5_outputs(1908) <= not(layer4_outputs(1168));
    layer5_outputs(1909) <= layer4_outputs(201);
    layer5_outputs(1910) <= (layer4_outputs(43)) and (layer4_outputs(2320));
    layer5_outputs(1911) <= not(layer4_outputs(2321));
    layer5_outputs(1912) <= not(layer4_outputs(1342));
    layer5_outputs(1913) <= '1';
    layer5_outputs(1914) <= layer4_outputs(1018);
    layer5_outputs(1915) <= (layer4_outputs(655)) and not (layer4_outputs(1550));
    layer5_outputs(1916) <= not((layer4_outputs(2178)) or (layer4_outputs(2038)));
    layer5_outputs(1917) <= not(layer4_outputs(1799));
    layer5_outputs(1918) <= layer4_outputs(1977);
    layer5_outputs(1919) <= not((layer4_outputs(674)) or (layer4_outputs(780)));
    layer5_outputs(1920) <= not(layer4_outputs(202));
    layer5_outputs(1921) <= layer4_outputs(543);
    layer5_outputs(1922) <= not(layer4_outputs(751));
    layer5_outputs(1923) <= (layer4_outputs(535)) and not (layer4_outputs(1876));
    layer5_outputs(1924) <= not(layer4_outputs(1912));
    layer5_outputs(1925) <= not((layer4_outputs(517)) or (layer4_outputs(990)));
    layer5_outputs(1926) <= layer4_outputs(454);
    layer5_outputs(1927) <= layer4_outputs(1011);
    layer5_outputs(1928) <= layer4_outputs(2503);
    layer5_outputs(1929) <= not((layer4_outputs(392)) and (layer4_outputs(924)));
    layer5_outputs(1930) <= (layer4_outputs(1266)) and (layer4_outputs(8));
    layer5_outputs(1931) <= layer4_outputs(1661);
    layer5_outputs(1932) <= '0';
    layer5_outputs(1933) <= not(layer4_outputs(637));
    layer5_outputs(1934) <= not(layer4_outputs(2375)) or (layer4_outputs(1007));
    layer5_outputs(1935) <= not((layer4_outputs(980)) xor (layer4_outputs(1588)));
    layer5_outputs(1936) <= not(layer4_outputs(364)) or (layer4_outputs(1613));
    layer5_outputs(1937) <= not(layer4_outputs(2067));
    layer5_outputs(1938) <= not((layer4_outputs(414)) or (layer4_outputs(1854)));
    layer5_outputs(1939) <= not(layer4_outputs(801));
    layer5_outputs(1940) <= (layer4_outputs(1008)) xor (layer4_outputs(2468));
    layer5_outputs(1941) <= layer4_outputs(18);
    layer5_outputs(1942) <= layer4_outputs(1906);
    layer5_outputs(1943) <= '1';
    layer5_outputs(1944) <= not((layer4_outputs(439)) xor (layer4_outputs(768)));
    layer5_outputs(1945) <= layer4_outputs(2317);
    layer5_outputs(1946) <= not((layer4_outputs(2472)) or (layer4_outputs(554)));
    layer5_outputs(1947) <= not((layer4_outputs(2118)) and (layer4_outputs(765)));
    layer5_outputs(1948) <= layer4_outputs(1066);
    layer5_outputs(1949) <= not(layer4_outputs(347));
    layer5_outputs(1950) <= not(layer4_outputs(1801));
    layer5_outputs(1951) <= (layer4_outputs(191)) and (layer4_outputs(1001));
    layer5_outputs(1952) <= not((layer4_outputs(2385)) and (layer4_outputs(1592)));
    layer5_outputs(1953) <= layer4_outputs(1488);
    layer5_outputs(1954) <= not((layer4_outputs(747)) or (layer4_outputs(2107)));
    layer5_outputs(1955) <= layer4_outputs(1465);
    layer5_outputs(1956) <= layer4_outputs(1708);
    layer5_outputs(1957) <= not(layer4_outputs(1621));
    layer5_outputs(1958) <= (layer4_outputs(330)) and not (layer4_outputs(584));
    layer5_outputs(1959) <= not(layer4_outputs(2510));
    layer5_outputs(1960) <= layer4_outputs(262);
    layer5_outputs(1961) <= layer4_outputs(2210);
    layer5_outputs(1962) <= (layer4_outputs(2414)) and not (layer4_outputs(1078));
    layer5_outputs(1963) <= not(layer4_outputs(2471));
    layer5_outputs(1964) <= layer4_outputs(1279);
    layer5_outputs(1965) <= not((layer4_outputs(1935)) or (layer4_outputs(1297)));
    layer5_outputs(1966) <= not(layer4_outputs(744));
    layer5_outputs(1967) <= (layer4_outputs(2206)) or (layer4_outputs(1396));
    layer5_outputs(1968) <= layer4_outputs(2123);
    layer5_outputs(1969) <= (layer4_outputs(625)) and not (layer4_outputs(1636));
    layer5_outputs(1970) <= (layer4_outputs(128)) and (layer4_outputs(2140));
    layer5_outputs(1971) <= (layer4_outputs(2135)) and not (layer4_outputs(1682));
    layer5_outputs(1972) <= '1';
    layer5_outputs(1973) <= not(layer4_outputs(1161));
    layer5_outputs(1974) <= layer4_outputs(554);
    layer5_outputs(1975) <= not(layer4_outputs(1015));
    layer5_outputs(1976) <= not(layer4_outputs(478)) or (layer4_outputs(990));
    layer5_outputs(1977) <= not(layer4_outputs(2288));
    layer5_outputs(1978) <= layer4_outputs(274);
    layer5_outputs(1979) <= not(layer4_outputs(2306));
    layer5_outputs(1980) <= not(layer4_outputs(2149));
    layer5_outputs(1981) <= not((layer4_outputs(1864)) xor (layer4_outputs(2186)));
    layer5_outputs(1982) <= not(layer4_outputs(1031));
    layer5_outputs(1983) <= '1';
    layer5_outputs(1984) <= not(layer4_outputs(1360));
    layer5_outputs(1985) <= not(layer4_outputs(487)) or (layer4_outputs(791));
    layer5_outputs(1986) <= (layer4_outputs(457)) xor (layer4_outputs(2113));
    layer5_outputs(1987) <= not((layer4_outputs(375)) and (layer4_outputs(912)));
    layer5_outputs(1988) <= (layer4_outputs(763)) xor (layer4_outputs(2250));
    layer5_outputs(1989) <= (layer4_outputs(1243)) and (layer4_outputs(2315));
    layer5_outputs(1990) <= not(layer4_outputs(1152)) or (layer4_outputs(1136));
    layer5_outputs(1991) <= not((layer4_outputs(627)) or (layer4_outputs(88)));
    layer5_outputs(1992) <= not((layer4_outputs(2136)) xor (layer4_outputs(1619)));
    layer5_outputs(1993) <= not(layer4_outputs(1967));
    layer5_outputs(1994) <= layer4_outputs(1079);
    layer5_outputs(1995) <= not((layer4_outputs(2224)) or (layer4_outputs(488)));
    layer5_outputs(1996) <= (layer4_outputs(111)) and not (layer4_outputs(966));
    layer5_outputs(1997) <= (layer4_outputs(1662)) and not (layer4_outputs(374));
    layer5_outputs(1998) <= (layer4_outputs(2061)) and not (layer4_outputs(1857));
    layer5_outputs(1999) <= not(layer4_outputs(360));
    layer5_outputs(2000) <= (layer4_outputs(586)) or (layer4_outputs(2119));
    layer5_outputs(2001) <= not(layer4_outputs(1351));
    layer5_outputs(2002) <= not(layer4_outputs(1978)) or (layer4_outputs(1470));
    layer5_outputs(2003) <= layer4_outputs(452);
    layer5_outputs(2004) <= not((layer4_outputs(1796)) xor (layer4_outputs(2028)));
    layer5_outputs(2005) <= not(layer4_outputs(1345));
    layer5_outputs(2006) <= not(layer4_outputs(1910)) or (layer4_outputs(2433));
    layer5_outputs(2007) <= layer4_outputs(650);
    layer5_outputs(2008) <= (layer4_outputs(848)) or (layer4_outputs(1239));
    layer5_outputs(2009) <= not(layer4_outputs(372));
    layer5_outputs(2010) <= '0';
    layer5_outputs(2011) <= not((layer4_outputs(1224)) or (layer4_outputs(1219)));
    layer5_outputs(2012) <= (layer4_outputs(278)) or (layer4_outputs(2329));
    layer5_outputs(2013) <= not(layer4_outputs(909));
    layer5_outputs(2014) <= (layer4_outputs(1617)) and (layer4_outputs(1454));
    layer5_outputs(2015) <= not(layer4_outputs(982));
    layer5_outputs(2016) <= layer4_outputs(2356);
    layer5_outputs(2017) <= layer4_outputs(2050);
    layer5_outputs(2018) <= not(layer4_outputs(90));
    layer5_outputs(2019) <= (layer4_outputs(1765)) or (layer4_outputs(472));
    layer5_outputs(2020) <= not(layer4_outputs(2500));
    layer5_outputs(2021) <= (layer4_outputs(1576)) and not (layer4_outputs(265));
    layer5_outputs(2022) <= (layer4_outputs(1922)) or (layer4_outputs(1407));
    layer5_outputs(2023) <= not(layer4_outputs(892));
    layer5_outputs(2024) <= (layer4_outputs(913)) or (layer4_outputs(2045));
    layer5_outputs(2025) <= not(layer4_outputs(157)) or (layer4_outputs(1080));
    layer5_outputs(2026) <= not(layer4_outputs(1194));
    layer5_outputs(2027) <= layer4_outputs(2300);
    layer5_outputs(2028) <= not(layer4_outputs(1006));
    layer5_outputs(2029) <= not(layer4_outputs(1490)) or (layer4_outputs(1160));
    layer5_outputs(2030) <= (layer4_outputs(1163)) and not (layer4_outputs(2434));
    layer5_outputs(2031) <= (layer4_outputs(2115)) and not (layer4_outputs(1063));
    layer5_outputs(2032) <= (layer4_outputs(972)) and not (layer4_outputs(1791));
    layer5_outputs(2033) <= not(layer4_outputs(1216));
    layer5_outputs(2034) <= (layer4_outputs(1296)) or (layer4_outputs(769));
    layer5_outputs(2035) <= layer4_outputs(1432);
    layer5_outputs(2036) <= not(layer4_outputs(745));
    layer5_outputs(2037) <= not((layer4_outputs(2532)) and (layer4_outputs(1785)));
    layer5_outputs(2038) <= not((layer4_outputs(444)) and (layer4_outputs(1210)));
    layer5_outputs(2039) <= not(layer4_outputs(2110)) or (layer4_outputs(1097));
    layer5_outputs(2040) <= not(layer4_outputs(1777));
    layer5_outputs(2041) <= not((layer4_outputs(177)) xor (layer4_outputs(1941)));
    layer5_outputs(2042) <= (layer4_outputs(1326)) and (layer4_outputs(70));
    layer5_outputs(2043) <= layer4_outputs(1848);
    layer5_outputs(2044) <= (layer4_outputs(920)) xor (layer4_outputs(804));
    layer5_outputs(2045) <= not(layer4_outputs(261));
    layer5_outputs(2046) <= (layer4_outputs(1080)) and not (layer4_outputs(2257));
    layer5_outputs(2047) <= not(layer4_outputs(1483));
    layer5_outputs(2048) <= layer4_outputs(1014);
    layer5_outputs(2049) <= layer4_outputs(2152);
    layer5_outputs(2050) <= (layer4_outputs(1632)) or (layer4_outputs(152));
    layer5_outputs(2051) <= not(layer4_outputs(2268));
    layer5_outputs(2052) <= layer4_outputs(1715);
    layer5_outputs(2053) <= layer4_outputs(196);
    layer5_outputs(2054) <= not((layer4_outputs(2221)) or (layer4_outputs(763)));
    layer5_outputs(2055) <= (layer4_outputs(157)) and not (layer4_outputs(1316));
    layer5_outputs(2056) <= (layer4_outputs(292)) xor (layer4_outputs(973));
    layer5_outputs(2057) <= '1';
    layer5_outputs(2058) <= (layer4_outputs(1680)) and (layer4_outputs(1613));
    layer5_outputs(2059) <= (layer4_outputs(884)) and (layer4_outputs(754));
    layer5_outputs(2060) <= (layer4_outputs(1542)) and (layer4_outputs(1762));
    layer5_outputs(2061) <= not((layer4_outputs(1423)) or (layer4_outputs(1654)));
    layer5_outputs(2062) <= '1';
    layer5_outputs(2063) <= (layer4_outputs(928)) and (layer4_outputs(1967));
    layer5_outputs(2064) <= not(layer4_outputs(313));
    layer5_outputs(2065) <= (layer4_outputs(2085)) and not (layer4_outputs(1836));
    layer5_outputs(2066) <= not(layer4_outputs(2505)) or (layer4_outputs(134));
    layer5_outputs(2067) <= not((layer4_outputs(579)) and (layer4_outputs(2145)));
    layer5_outputs(2068) <= not(layer4_outputs(2330)) or (layer4_outputs(2072));
    layer5_outputs(2069) <= layer4_outputs(1817);
    layer5_outputs(2070) <= layer4_outputs(1475);
    layer5_outputs(2071) <= not(layer4_outputs(1887));
    layer5_outputs(2072) <= not(layer4_outputs(1794));
    layer5_outputs(2073) <= not((layer4_outputs(1187)) xor (layer4_outputs(320)));
    layer5_outputs(2074) <= layer4_outputs(576);
    layer5_outputs(2075) <= not(layer4_outputs(1962)) or (layer4_outputs(1005));
    layer5_outputs(2076) <= (layer4_outputs(1894)) and not (layer4_outputs(207));
    layer5_outputs(2077) <= (layer4_outputs(21)) or (layer4_outputs(1660));
    layer5_outputs(2078) <= (layer4_outputs(1652)) and (layer4_outputs(2096));
    layer5_outputs(2079) <= not(layer4_outputs(482));
    layer5_outputs(2080) <= layer4_outputs(2233);
    layer5_outputs(2081) <= not((layer4_outputs(1444)) and (layer4_outputs(1921)));
    layer5_outputs(2082) <= '0';
    layer5_outputs(2083) <= (layer4_outputs(2518)) and not (layer4_outputs(1054));
    layer5_outputs(2084) <= not(layer4_outputs(968));
    layer5_outputs(2085) <= layer4_outputs(2291);
    layer5_outputs(2086) <= not((layer4_outputs(353)) or (layer4_outputs(489)));
    layer5_outputs(2087) <= layer4_outputs(927);
    layer5_outputs(2088) <= layer4_outputs(940);
    layer5_outputs(2089) <= not((layer4_outputs(1093)) and (layer4_outputs(113)));
    layer5_outputs(2090) <= not(layer4_outputs(1355)) or (layer4_outputs(1048));
    layer5_outputs(2091) <= not(layer4_outputs(1551));
    layer5_outputs(2092) <= not((layer4_outputs(2465)) xor (layer4_outputs(1593)));
    layer5_outputs(2093) <= layer4_outputs(1859);
    layer5_outputs(2094) <= layer4_outputs(1971);
    layer5_outputs(2095) <= not(layer4_outputs(2537)) or (layer4_outputs(1249));
    layer5_outputs(2096) <= (layer4_outputs(502)) and (layer4_outputs(1267));
    layer5_outputs(2097) <= layer4_outputs(2259);
    layer5_outputs(2098) <= (layer4_outputs(2134)) xor (layer4_outputs(359));
    layer5_outputs(2099) <= layer4_outputs(923);
    layer5_outputs(2100) <= not(layer4_outputs(27));
    layer5_outputs(2101) <= layer4_outputs(415);
    layer5_outputs(2102) <= layer4_outputs(530);
    layer5_outputs(2103) <= not(layer4_outputs(244));
    layer5_outputs(2104) <= (layer4_outputs(921)) or (layer4_outputs(809));
    layer5_outputs(2105) <= not(layer4_outputs(2405));
    layer5_outputs(2106) <= layer4_outputs(1840);
    layer5_outputs(2107) <= not(layer4_outputs(1244));
    layer5_outputs(2108) <= (layer4_outputs(803)) xor (layer4_outputs(872));
    layer5_outputs(2109) <= not((layer4_outputs(312)) xor (layer4_outputs(178)));
    layer5_outputs(2110) <= (layer4_outputs(1435)) xor (layer4_outputs(321));
    layer5_outputs(2111) <= (layer4_outputs(533)) xor (layer4_outputs(380));
    layer5_outputs(2112) <= (layer4_outputs(1647)) and not (layer4_outputs(1858));
    layer5_outputs(2113) <= not(layer4_outputs(815));
    layer5_outputs(2114) <= (layer4_outputs(996)) and (layer4_outputs(1820));
    layer5_outputs(2115) <= layer4_outputs(506);
    layer5_outputs(2116) <= (layer4_outputs(2219)) xor (layer4_outputs(109));
    layer5_outputs(2117) <= not((layer4_outputs(450)) xor (layer4_outputs(1726)));
    layer5_outputs(2118) <= not((layer4_outputs(1823)) or (layer4_outputs(695)));
    layer5_outputs(2119) <= not(layer4_outputs(1975));
    layer5_outputs(2120) <= layer4_outputs(936);
    layer5_outputs(2121) <= not((layer4_outputs(341)) or (layer4_outputs(1959)));
    layer5_outputs(2122) <= (layer4_outputs(1000)) and (layer4_outputs(486));
    layer5_outputs(2123) <= (layer4_outputs(1088)) xor (layer4_outputs(1825));
    layer5_outputs(2124) <= not(layer4_outputs(2044));
    layer5_outputs(2125) <= layer4_outputs(1320);
    layer5_outputs(2126) <= not((layer4_outputs(775)) xor (layer4_outputs(2380)));
    layer5_outputs(2127) <= not(layer4_outputs(1744)) or (layer4_outputs(2421));
    layer5_outputs(2128) <= (layer4_outputs(610)) and (layer4_outputs(1456));
    layer5_outputs(2129) <= '1';
    layer5_outputs(2130) <= '0';
    layer5_outputs(2131) <= layer4_outputs(2081);
    layer5_outputs(2132) <= not(layer4_outputs(284));
    layer5_outputs(2133) <= not(layer4_outputs(1342));
    layer5_outputs(2134) <= not(layer4_outputs(2144));
    layer5_outputs(2135) <= (layer4_outputs(933)) xor (layer4_outputs(1559));
    layer5_outputs(2136) <= not(layer4_outputs(2174)) or (layer4_outputs(123));
    layer5_outputs(2137) <= layer4_outputs(1468);
    layer5_outputs(2138) <= layer4_outputs(1235);
    layer5_outputs(2139) <= not((layer4_outputs(1201)) or (layer4_outputs(1087)));
    layer5_outputs(2140) <= (layer4_outputs(501)) or (layer4_outputs(2554));
    layer5_outputs(2141) <= not(layer4_outputs(2543));
    layer5_outputs(2142) <= (layer4_outputs(116)) xor (layer4_outputs(799));
    layer5_outputs(2143) <= not(layer4_outputs(918));
    layer5_outputs(2144) <= not(layer4_outputs(946)) or (layer4_outputs(2523));
    layer5_outputs(2145) <= layer4_outputs(39);
    layer5_outputs(2146) <= not((layer4_outputs(1347)) or (layer4_outputs(245)));
    layer5_outputs(2147) <= not(layer4_outputs(1957));
    layer5_outputs(2148) <= not(layer4_outputs(1466)) or (layer4_outputs(1096));
    layer5_outputs(2149) <= (layer4_outputs(326)) and not (layer4_outputs(1970));
    layer5_outputs(2150) <= not(layer4_outputs(1779)) or (layer4_outputs(1250));
    layer5_outputs(2151) <= (layer4_outputs(1722)) xor (layer4_outputs(828));
    layer5_outputs(2152) <= (layer4_outputs(1678)) xor (layer4_outputs(2383));
    layer5_outputs(2153) <= '1';
    layer5_outputs(2154) <= (layer4_outputs(737)) xor (layer4_outputs(264));
    layer5_outputs(2155) <= not(layer4_outputs(205));
    layer5_outputs(2156) <= layer4_outputs(2444);
    layer5_outputs(2157) <= '0';
    layer5_outputs(2158) <= not(layer4_outputs(76));
    layer5_outputs(2159) <= layer4_outputs(1348);
    layer5_outputs(2160) <= not(layer4_outputs(425));
    layer5_outputs(2161) <= not((layer4_outputs(423)) and (layer4_outputs(1956)));
    layer5_outputs(2162) <= not(layer4_outputs(1188)) or (layer4_outputs(343));
    layer5_outputs(2163) <= not((layer4_outputs(787)) xor (layer4_outputs(1953)));
    layer5_outputs(2164) <= layer4_outputs(2456);
    layer5_outputs(2165) <= layer4_outputs(45);
    layer5_outputs(2166) <= layer4_outputs(1952);
    layer5_outputs(2167) <= '0';
    layer5_outputs(2168) <= layer4_outputs(525);
    layer5_outputs(2169) <= layer4_outputs(2164);
    layer5_outputs(2170) <= (layer4_outputs(322)) and (layer4_outputs(1737));
    layer5_outputs(2171) <= (layer4_outputs(1099)) xor (layer4_outputs(2381));
    layer5_outputs(2172) <= (layer4_outputs(1512)) or (layer4_outputs(1576));
    layer5_outputs(2173) <= layer4_outputs(2546);
    layer5_outputs(2174) <= not(layer4_outputs(1479));
    layer5_outputs(2175) <= (layer4_outputs(661)) xor (layer4_outputs(721));
    layer5_outputs(2176) <= not((layer4_outputs(287)) or (layer4_outputs(1955)));
    layer5_outputs(2177) <= '1';
    layer5_outputs(2178) <= not(layer4_outputs(1544));
    layer5_outputs(2179) <= not((layer4_outputs(1679)) xor (layer4_outputs(1371)));
    layer5_outputs(2180) <= not(layer4_outputs(32));
    layer5_outputs(2181) <= (layer4_outputs(2009)) or (layer4_outputs(2142));
    layer5_outputs(2182) <= layer4_outputs(1530);
    layer5_outputs(2183) <= (layer4_outputs(256)) or (layer4_outputs(968));
    layer5_outputs(2184) <= not(layer4_outputs(21));
    layer5_outputs(2185) <= layer4_outputs(2349);
    layer5_outputs(2186) <= not(layer4_outputs(660)) or (layer4_outputs(1595));
    layer5_outputs(2187) <= layer4_outputs(2230);
    layer5_outputs(2188) <= (layer4_outputs(1681)) and not (layer4_outputs(1085));
    layer5_outputs(2189) <= not((layer4_outputs(1127)) xor (layer4_outputs(1140)));
    layer5_outputs(2190) <= layer4_outputs(1863);
    layer5_outputs(2191) <= not(layer4_outputs(1780));
    layer5_outputs(2192) <= layer4_outputs(2403);
    layer5_outputs(2193) <= (layer4_outputs(1130)) and not (layer4_outputs(1207));
    layer5_outputs(2194) <= not(layer4_outputs(2084)) or (layer4_outputs(1094));
    layer5_outputs(2195) <= layer4_outputs(1770);
    layer5_outputs(2196) <= not(layer4_outputs(2080));
    layer5_outputs(2197) <= layer4_outputs(878);
    layer5_outputs(2198) <= not(layer4_outputs(2000)) or (layer4_outputs(2093));
    layer5_outputs(2199) <= layer4_outputs(1230);
    layer5_outputs(2200) <= not((layer4_outputs(2274)) or (layer4_outputs(114)));
    layer5_outputs(2201) <= (layer4_outputs(2501)) and not (layer4_outputs(1975));
    layer5_outputs(2202) <= not(layer4_outputs(1853)) or (layer4_outputs(682));
    layer5_outputs(2203) <= not(layer4_outputs(32));
    layer5_outputs(2204) <= '1';
    layer5_outputs(2205) <= '1';
    layer5_outputs(2206) <= (layer4_outputs(874)) and not (layer4_outputs(1280));
    layer5_outputs(2207) <= not(layer4_outputs(2460));
    layer5_outputs(2208) <= not(layer4_outputs(612));
    layer5_outputs(2209) <= not(layer4_outputs(1592)) or (layer4_outputs(931));
    layer5_outputs(2210) <= not(layer4_outputs(1703));
    layer5_outputs(2211) <= '0';
    layer5_outputs(2212) <= not(layer4_outputs(2226)) or (layer4_outputs(253));
    layer5_outputs(2213) <= not((layer4_outputs(114)) xor (layer4_outputs(49)));
    layer5_outputs(2214) <= not((layer4_outputs(2033)) or (layer4_outputs(1514)));
    layer5_outputs(2215) <= (layer4_outputs(817)) and not (layer4_outputs(243));
    layer5_outputs(2216) <= (layer4_outputs(1839)) or (layer4_outputs(2464));
    layer5_outputs(2217) <= (layer4_outputs(1149)) and not (layer4_outputs(533));
    layer5_outputs(2218) <= not(layer4_outputs(2162));
    layer5_outputs(2219) <= not((layer4_outputs(2031)) and (layer4_outputs(959)));
    layer5_outputs(2220) <= not(layer4_outputs(1311));
    layer5_outputs(2221) <= layer4_outputs(1495);
    layer5_outputs(2222) <= layer4_outputs(1471);
    layer5_outputs(2223) <= layer4_outputs(403);
    layer5_outputs(2224) <= not((layer4_outputs(38)) and (layer4_outputs(2353)));
    layer5_outputs(2225) <= not((layer4_outputs(2111)) xor (layer4_outputs(534)));
    layer5_outputs(2226) <= (layer4_outputs(1329)) xor (layer4_outputs(621));
    layer5_outputs(2227) <= layer4_outputs(365);
    layer5_outputs(2228) <= layer4_outputs(688);
    layer5_outputs(2229) <= (layer4_outputs(1125)) and not (layer4_outputs(1237));
    layer5_outputs(2230) <= not((layer4_outputs(436)) or (layer4_outputs(1730)));
    layer5_outputs(2231) <= not(layer4_outputs(841));
    layer5_outputs(2232) <= layer4_outputs(979);
    layer5_outputs(2233) <= not(layer4_outputs(2479)) or (layer4_outputs(2413));
    layer5_outputs(2234) <= not(layer4_outputs(1598));
    layer5_outputs(2235) <= not(layer4_outputs(359)) or (layer4_outputs(1234));
    layer5_outputs(2236) <= (layer4_outputs(720)) or (layer4_outputs(53));
    layer5_outputs(2237) <= layer4_outputs(1121);
    layer5_outputs(2238) <= not(layer4_outputs(1236));
    layer5_outputs(2239) <= (layer4_outputs(269)) xor (layer4_outputs(544));
    layer5_outputs(2240) <= not(layer4_outputs(1534)) or (layer4_outputs(1004));
    layer5_outputs(2241) <= layer4_outputs(2073);
    layer5_outputs(2242) <= (layer4_outputs(1054)) or (layer4_outputs(1548));
    layer5_outputs(2243) <= layer4_outputs(2233);
    layer5_outputs(2244) <= not((layer4_outputs(1957)) xor (layer4_outputs(676)));
    layer5_outputs(2245) <= not((layer4_outputs(1528)) xor (layer4_outputs(1382)));
    layer5_outputs(2246) <= not((layer4_outputs(2014)) and (layer4_outputs(1104)));
    layer5_outputs(2247) <= not(layer4_outputs(2082)) or (layer4_outputs(473));
    layer5_outputs(2248) <= not(layer4_outputs(537));
    layer5_outputs(2249) <= (layer4_outputs(210)) and (layer4_outputs(230));
    layer5_outputs(2250) <= (layer4_outputs(592)) and (layer4_outputs(2265));
    layer5_outputs(2251) <= '0';
    layer5_outputs(2252) <= not(layer4_outputs(1950));
    layer5_outputs(2253) <= (layer4_outputs(918)) or (layer4_outputs(1702));
    layer5_outputs(2254) <= (layer4_outputs(2350)) or (layer4_outputs(565));
    layer5_outputs(2255) <= not(layer4_outputs(1612));
    layer5_outputs(2256) <= (layer4_outputs(2519)) and (layer4_outputs(1254));
    layer5_outputs(2257) <= not(layer4_outputs(571)) or (layer4_outputs(1558));
    layer5_outputs(2258) <= (layer4_outputs(421)) and (layer4_outputs(1045));
    layer5_outputs(2259) <= (layer4_outputs(911)) and not (layer4_outputs(332));
    layer5_outputs(2260) <= not(layer4_outputs(1369));
    layer5_outputs(2261) <= not(layer4_outputs(492));
    layer5_outputs(2262) <= (layer4_outputs(589)) xor (layer4_outputs(1381));
    layer5_outputs(2263) <= not(layer4_outputs(910)) or (layer4_outputs(546));
    layer5_outputs(2264) <= not((layer4_outputs(1201)) xor (layer4_outputs(1394)));
    layer5_outputs(2265) <= not(layer4_outputs(1529));
    layer5_outputs(2266) <= not(layer4_outputs(1988));
    layer5_outputs(2267) <= layer4_outputs(496);
    layer5_outputs(2268) <= not(layer4_outputs(733)) or (layer4_outputs(2231));
    layer5_outputs(2269) <= not(layer4_outputs(736));
    layer5_outputs(2270) <= not(layer4_outputs(1653));
    layer5_outputs(2271) <= layer4_outputs(1556);
    layer5_outputs(2272) <= not(layer4_outputs(344));
    layer5_outputs(2273) <= not(layer4_outputs(110));
    layer5_outputs(2274) <= not(layer4_outputs(2242));
    layer5_outputs(2275) <= not(layer4_outputs(2272));
    layer5_outputs(2276) <= not((layer4_outputs(522)) or (layer4_outputs(122)));
    layer5_outputs(2277) <= (layer4_outputs(211)) and (layer4_outputs(573));
    layer5_outputs(2278) <= layer4_outputs(2278);
    layer5_outputs(2279) <= layer4_outputs(1850);
    layer5_outputs(2280) <= (layer4_outputs(1940)) xor (layer4_outputs(1084));
    layer5_outputs(2281) <= layer4_outputs(2494);
    layer5_outputs(2282) <= layer4_outputs(732);
    layer5_outputs(2283) <= not((layer4_outputs(300)) or (layer4_outputs(2166)));
    layer5_outputs(2284) <= not(layer4_outputs(2001));
    layer5_outputs(2285) <= not(layer4_outputs(245)) or (layer4_outputs(1268));
    layer5_outputs(2286) <= not((layer4_outputs(513)) and (layer4_outputs(1486)));
    layer5_outputs(2287) <= not(layer4_outputs(217));
    layer5_outputs(2288) <= not((layer4_outputs(1484)) or (layer4_outputs(4)));
    layer5_outputs(2289) <= not((layer4_outputs(2435)) xor (layer4_outputs(169)));
    layer5_outputs(2290) <= not((layer4_outputs(1058)) or (layer4_outputs(725)));
    layer5_outputs(2291) <= (layer4_outputs(1327)) and not (layer4_outputs(2055));
    layer5_outputs(2292) <= (layer4_outputs(1997)) and not (layer4_outputs(1023));
    layer5_outputs(2293) <= not((layer4_outputs(2470)) and (layer4_outputs(1658)));
    layer5_outputs(2294) <= (layer4_outputs(742)) and not (layer4_outputs(307));
    layer5_outputs(2295) <= (layer4_outputs(2015)) and not (layer4_outputs(442));
    layer5_outputs(2296) <= (layer4_outputs(756)) and not (layer4_outputs(223));
    layer5_outputs(2297) <= (layer4_outputs(454)) and (layer4_outputs(2489));
    layer5_outputs(2298) <= not(layer4_outputs(1291));
    layer5_outputs(2299) <= not((layer4_outputs(845)) xor (layer4_outputs(1261)));
    layer5_outputs(2300) <= (layer4_outputs(1397)) and (layer4_outputs(1723));
    layer5_outputs(2301) <= layer4_outputs(640);
    layer5_outputs(2302) <= not(layer4_outputs(2182)) or (layer4_outputs(2331));
    layer5_outputs(2303) <= not((layer4_outputs(1918)) or (layer4_outputs(70)));
    layer5_outputs(2304) <= layer4_outputs(1246);
    layer5_outputs(2305) <= not(layer4_outputs(1782)) or (layer4_outputs(1055));
    layer5_outputs(2306) <= layer4_outputs(1295);
    layer5_outputs(2307) <= not(layer4_outputs(448));
    layer5_outputs(2308) <= layer4_outputs(1026);
    layer5_outputs(2309) <= (layer4_outputs(2429)) and not (layer4_outputs(1701));
    layer5_outputs(2310) <= '0';
    layer5_outputs(2311) <= not((layer4_outputs(2217)) xor (layer4_outputs(2084)));
    layer5_outputs(2312) <= not(layer4_outputs(1483));
    layer5_outputs(2313) <= not((layer4_outputs(107)) xor (layer4_outputs(16)));
    layer5_outputs(2314) <= (layer4_outputs(46)) and (layer4_outputs(917));
    layer5_outputs(2315) <= '1';
    layer5_outputs(2316) <= (layer4_outputs(1401)) and not (layer4_outputs(1064));
    layer5_outputs(2317) <= not(layer4_outputs(797));
    layer5_outputs(2318) <= (layer4_outputs(468)) and not (layer4_outputs(2504));
    layer5_outputs(2319) <= not(layer4_outputs(2058));
    layer5_outputs(2320) <= layer4_outputs(1096);
    layer5_outputs(2321) <= not((layer4_outputs(1697)) or (layer4_outputs(75)));
    layer5_outputs(2322) <= not(layer4_outputs(1722));
    layer5_outputs(2323) <= (layer4_outputs(1633)) and not (layer4_outputs(610));
    layer5_outputs(2324) <= layer4_outputs(1035);
    layer5_outputs(2325) <= layer4_outputs(939);
    layer5_outputs(2326) <= not((layer4_outputs(42)) and (layer4_outputs(1295)));
    layer5_outputs(2327) <= not(layer4_outputs(782)) or (layer4_outputs(2276));
    layer5_outputs(2328) <= not(layer4_outputs(532));
    layer5_outputs(2329) <= (layer4_outputs(1787)) or (layer4_outputs(1116));
    layer5_outputs(2330) <= not((layer4_outputs(1970)) xor (layer4_outputs(2309)));
    layer5_outputs(2331) <= not(layer4_outputs(2096));
    layer5_outputs(2332) <= not(layer4_outputs(1248)) or (layer4_outputs(534));
    layer5_outputs(2333) <= not(layer4_outputs(1424));
    layer5_outputs(2334) <= not(layer4_outputs(1081));
    layer5_outputs(2335) <= '0';
    layer5_outputs(2336) <= (layer4_outputs(1339)) and (layer4_outputs(1226));
    layer5_outputs(2337) <= layer4_outputs(397);
    layer5_outputs(2338) <= not(layer4_outputs(1076));
    layer5_outputs(2339) <= not(layer4_outputs(481));
    layer5_outputs(2340) <= not(layer4_outputs(658));
    layer5_outputs(2341) <= not(layer4_outputs(1189));
    layer5_outputs(2342) <= (layer4_outputs(1442)) or (layer4_outputs(1289));
    layer5_outputs(2343) <= not(layer4_outputs(56));
    layer5_outputs(2344) <= not((layer4_outputs(1425)) or (layer4_outputs(1117)));
    layer5_outputs(2345) <= '0';
    layer5_outputs(2346) <= layer4_outputs(2234);
    layer5_outputs(2347) <= (layer4_outputs(1095)) xor (layer4_outputs(2370));
    layer5_outputs(2348) <= layer4_outputs(1370);
    layer5_outputs(2349) <= not((layer4_outputs(2097)) and (layer4_outputs(2545)));
    layer5_outputs(2350) <= layer4_outputs(1279);
    layer5_outputs(2351) <= (layer4_outputs(2052)) or (layer4_outputs(2528));
    layer5_outputs(2352) <= layer4_outputs(221);
    layer5_outputs(2353) <= layer4_outputs(133);
    layer5_outputs(2354) <= not((layer4_outputs(950)) or (layer4_outputs(1949)));
    layer5_outputs(2355) <= not(layer4_outputs(823));
    layer5_outputs(2356) <= (layer4_outputs(1275)) and not (layer4_outputs(952));
    layer5_outputs(2357) <= (layer4_outputs(807)) and not (layer4_outputs(2236));
    layer5_outputs(2358) <= not(layer4_outputs(1913));
    layer5_outputs(2359) <= (layer4_outputs(565)) xor (layer4_outputs(1013));
    layer5_outputs(2360) <= not(layer4_outputs(1734));
    layer5_outputs(2361) <= not(layer4_outputs(870)) or (layer4_outputs(2365));
    layer5_outputs(2362) <= (layer4_outputs(2302)) and not (layer4_outputs(835));
    layer5_outputs(2363) <= not(layer4_outputs(1616));
    layer5_outputs(2364) <= not(layer4_outputs(2215)) or (layer4_outputs(2058));
    layer5_outputs(2365) <= not((layer4_outputs(603)) or (layer4_outputs(280)));
    layer5_outputs(2366) <= not(layer4_outputs(1183)) or (layer4_outputs(495));
    layer5_outputs(2367) <= not(layer4_outputs(1259));
    layer5_outputs(2368) <= layer4_outputs(1946);
    layer5_outputs(2369) <= not(layer4_outputs(1028));
    layer5_outputs(2370) <= (layer4_outputs(420)) or (layer4_outputs(1842));
    layer5_outputs(2371) <= not(layer4_outputs(2165));
    layer5_outputs(2372) <= not(layer4_outputs(635));
    layer5_outputs(2373) <= layer4_outputs(708);
    layer5_outputs(2374) <= (layer4_outputs(252)) and (layer4_outputs(1499));
    layer5_outputs(2375) <= not(layer4_outputs(278)) or (layer4_outputs(407));
    layer5_outputs(2376) <= layer4_outputs(1555);
    layer5_outputs(2377) <= not(layer4_outputs(994));
    layer5_outputs(2378) <= not(layer4_outputs(1129)) or (layer4_outputs(305));
    layer5_outputs(2379) <= (layer4_outputs(2077)) and not (layer4_outputs(556));
    layer5_outputs(2380) <= not((layer4_outputs(1839)) and (layer4_outputs(1200)));
    layer5_outputs(2381) <= not(layer4_outputs(2417));
    layer5_outputs(2382) <= layer4_outputs(6);
    layer5_outputs(2383) <= not(layer4_outputs(1866)) or (layer4_outputs(1351));
    layer5_outputs(2384) <= layer4_outputs(1772);
    layer5_outputs(2385) <= not(layer4_outputs(2477)) or (layer4_outputs(2070));
    layer5_outputs(2386) <= layer4_outputs(1105);
    layer5_outputs(2387) <= (layer4_outputs(279)) or (layer4_outputs(961));
    layer5_outputs(2388) <= (layer4_outputs(1123)) xor (layer4_outputs(944));
    layer5_outputs(2389) <= not((layer4_outputs(370)) or (layer4_outputs(1982)));
    layer5_outputs(2390) <= (layer4_outputs(879)) or (layer4_outputs(2455));
    layer5_outputs(2391) <= not(layer4_outputs(2280));
    layer5_outputs(2392) <= layer4_outputs(334);
    layer5_outputs(2393) <= (layer4_outputs(1631)) and not (layer4_outputs(1683));
    layer5_outputs(2394) <= '0';
    layer5_outputs(2395) <= (layer4_outputs(2161)) or (layer4_outputs(868));
    layer5_outputs(2396) <= not(layer4_outputs(945)) or (layer4_outputs(569));
    layer5_outputs(2397) <= (layer4_outputs(1299)) and not (layer4_outputs(1523));
    layer5_outputs(2398) <= not(layer4_outputs(869)) or (layer4_outputs(1766));
    layer5_outputs(2399) <= not(layer4_outputs(1844));
    layer5_outputs(2400) <= '0';
    layer5_outputs(2401) <= not(layer4_outputs(656));
    layer5_outputs(2402) <= not(layer4_outputs(438)) or (layer4_outputs(175));
    layer5_outputs(2403) <= layer4_outputs(2336);
    layer5_outputs(2404) <= not(layer4_outputs(1422));
    layer5_outputs(2405) <= not(layer4_outputs(2082));
    layer5_outputs(2406) <= not((layer4_outputs(498)) and (layer4_outputs(1190)));
    layer5_outputs(2407) <= not((layer4_outputs(480)) and (layer4_outputs(1019)));
    layer5_outputs(2408) <= layer4_outputs(1604);
    layer5_outputs(2409) <= layer4_outputs(1939);
    layer5_outputs(2410) <= not((layer4_outputs(1893)) or (layer4_outputs(590)));
    layer5_outputs(2411) <= layer4_outputs(1398);
    layer5_outputs(2412) <= not(layer4_outputs(1032)) or (layer4_outputs(1057));
    layer5_outputs(2413) <= not(layer4_outputs(400)) or (layer4_outputs(1778));
    layer5_outputs(2414) <= layer4_outputs(409);
    layer5_outputs(2415) <= not(layer4_outputs(2159));
    layer5_outputs(2416) <= not((layer4_outputs(1318)) and (layer4_outputs(1502)));
    layer5_outputs(2417) <= not(layer4_outputs(848));
    layer5_outputs(2418) <= (layer4_outputs(358)) and not (layer4_outputs(2499));
    layer5_outputs(2419) <= not(layer4_outputs(77));
    layer5_outputs(2420) <= layer4_outputs(257);
    layer5_outputs(2421) <= layer4_outputs(452);
    layer5_outputs(2422) <= (layer4_outputs(644)) and (layer4_outputs(785));
    layer5_outputs(2423) <= not((layer4_outputs(805)) and (layer4_outputs(855)));
    layer5_outputs(2424) <= not(layer4_outputs(293));
    layer5_outputs(2425) <= layer4_outputs(599);
    layer5_outputs(2426) <= (layer4_outputs(608)) and (layer4_outputs(1414));
    layer5_outputs(2427) <= (layer4_outputs(594)) and not (layer4_outputs(1680));
    layer5_outputs(2428) <= not(layer4_outputs(1555));
    layer5_outputs(2429) <= (layer4_outputs(810)) and not (layer4_outputs(1566));
    layer5_outputs(2430) <= '1';
    layer5_outputs(2431) <= layer4_outputs(2335);
    layer5_outputs(2432) <= not((layer4_outputs(1208)) xor (layer4_outputs(476)));
    layer5_outputs(2433) <= layer4_outputs(529);
    layer5_outputs(2434) <= not(layer4_outputs(211)) or (layer4_outputs(2413));
    layer5_outputs(2435) <= not(layer4_outputs(1845));
    layer5_outputs(2436) <= (layer4_outputs(2432)) xor (layer4_outputs(811));
    layer5_outputs(2437) <= layer4_outputs(1482);
    layer5_outputs(2438) <= not(layer4_outputs(165)) or (layer4_outputs(2526));
    layer5_outputs(2439) <= not(layer4_outputs(1571));
    layer5_outputs(2440) <= not(layer4_outputs(466));
    layer5_outputs(2441) <= not(layer4_outputs(629));
    layer5_outputs(2442) <= (layer4_outputs(1719)) and not (layer4_outputs(185));
    layer5_outputs(2443) <= not((layer4_outputs(1675)) or (layer4_outputs(2445)));
    layer5_outputs(2444) <= not((layer4_outputs(164)) and (layer4_outputs(1464)));
    layer5_outputs(2445) <= not(layer4_outputs(2265)) or (layer4_outputs(2550));
    layer5_outputs(2446) <= not((layer4_outputs(1882)) and (layer4_outputs(2106)));
    layer5_outputs(2447) <= (layer4_outputs(1305)) and not (layer4_outputs(2542));
    layer5_outputs(2448) <= (layer4_outputs(239)) and (layer4_outputs(649));
    layer5_outputs(2449) <= not((layer4_outputs(251)) xor (layer4_outputs(2395)));
    layer5_outputs(2450) <= layer4_outputs(523);
    layer5_outputs(2451) <= (layer4_outputs(198)) and not (layer4_outputs(596));
    layer5_outputs(2452) <= (layer4_outputs(1195)) and not (layer4_outputs(935));
    layer5_outputs(2453) <= not(layer4_outputs(2129));
    layer5_outputs(2454) <= not(layer4_outputs(1448));
    layer5_outputs(2455) <= not(layer4_outputs(1685)) or (layer4_outputs(194));
    layer5_outputs(2456) <= (layer4_outputs(209)) xor (layer4_outputs(1504));
    layer5_outputs(2457) <= (layer4_outputs(780)) and (layer4_outputs(1898));
    layer5_outputs(2458) <= not((layer4_outputs(2169)) xor (layer4_outputs(1332)));
    layer5_outputs(2459) <= layer4_outputs(789);
    layer5_outputs(2460) <= layer4_outputs(51);
    layer5_outputs(2461) <= not((layer4_outputs(893)) xor (layer4_outputs(1549)));
    layer5_outputs(2462) <= not(layer4_outputs(1735));
    layer5_outputs(2463) <= layer4_outputs(373);
    layer5_outputs(2464) <= not((layer4_outputs(591)) xor (layer4_outputs(1554)));
    layer5_outputs(2465) <= layer4_outputs(536);
    layer5_outputs(2466) <= (layer4_outputs(1030)) xor (layer4_outputs(264));
    layer5_outputs(2467) <= (layer4_outputs(1756)) and not (layer4_outputs(1109));
    layer5_outputs(2468) <= not((layer4_outputs(263)) or (layer4_outputs(1039)));
    layer5_outputs(2469) <= not(layer4_outputs(818));
    layer5_outputs(2470) <= (layer4_outputs(1132)) and not (layer4_outputs(607));
    layer5_outputs(2471) <= (layer4_outputs(2338)) and not (layer4_outputs(1760));
    layer5_outputs(2472) <= not(layer4_outputs(2351));
    layer5_outputs(2473) <= not(layer4_outputs(1092)) or (layer4_outputs(2368));
    layer5_outputs(2474) <= layer4_outputs(882);
    layer5_outputs(2475) <= (layer4_outputs(1237)) and (layer4_outputs(914));
    layer5_outputs(2476) <= (layer4_outputs(303)) and (layer4_outputs(723));
    layer5_outputs(2477) <= (layer4_outputs(382)) and (layer4_outputs(2530));
    layer5_outputs(2478) <= not(layer4_outputs(1739));
    layer5_outputs(2479) <= (layer4_outputs(1251)) or (layer4_outputs(1966));
    layer5_outputs(2480) <= '0';
    layer5_outputs(2481) <= (layer4_outputs(850)) xor (layer4_outputs(1270));
    layer5_outputs(2482) <= (layer4_outputs(216)) and not (layer4_outputs(2311));
    layer5_outputs(2483) <= layer4_outputs(2463);
    layer5_outputs(2484) <= (layer4_outputs(1803)) xor (layer4_outputs(1443));
    layer5_outputs(2485) <= not((layer4_outputs(1111)) and (layer4_outputs(635)));
    layer5_outputs(2486) <= not(layer4_outputs(2033)) or (layer4_outputs(1908));
    layer5_outputs(2487) <= (layer4_outputs(1290)) and not (layer4_outputs(1834));
    layer5_outputs(2488) <= not(layer4_outputs(459));
    layer5_outputs(2489) <= not(layer4_outputs(2510));
    layer5_outputs(2490) <= layer4_outputs(957);
    layer5_outputs(2491) <= layer4_outputs(1932);
    layer5_outputs(2492) <= layer4_outputs(272);
    layer5_outputs(2493) <= not((layer4_outputs(96)) and (layer4_outputs(223)));
    layer5_outputs(2494) <= layer4_outputs(1014);
    layer5_outputs(2495) <= (layer4_outputs(484)) xor (layer4_outputs(696));
    layer5_outputs(2496) <= not((layer4_outputs(2306)) and (layer4_outputs(2251)));
    layer5_outputs(2497) <= not(layer4_outputs(243));
    layer5_outputs(2498) <= not((layer4_outputs(511)) or (layer4_outputs(810)));
    layer5_outputs(2499) <= not(layer4_outputs(2274)) or (layer4_outputs(1053));
    layer5_outputs(2500) <= '1';
    layer5_outputs(2501) <= not(layer4_outputs(747));
    layer5_outputs(2502) <= (layer4_outputs(2157)) and not (layer4_outputs(2446));
    layer5_outputs(2503) <= layer4_outputs(1590);
    layer5_outputs(2504) <= not(layer4_outputs(1729));
    layer5_outputs(2505) <= (layer4_outputs(2160)) or (layer4_outputs(717));
    layer5_outputs(2506) <= (layer4_outputs(2192)) and not (layer4_outputs(2546));
    layer5_outputs(2507) <= layer4_outputs(1292);
    layer5_outputs(2508) <= (layer4_outputs(237)) or (layer4_outputs(459));
    layer5_outputs(2509) <= layer4_outputs(383);
    layer5_outputs(2510) <= (layer4_outputs(1602)) and not (layer4_outputs(1421));
    layer5_outputs(2511) <= layer4_outputs(509);
    layer5_outputs(2512) <= layer4_outputs(884);
    layer5_outputs(2513) <= (layer4_outputs(981)) and (layer4_outputs(331));
    layer5_outputs(2514) <= not(layer4_outputs(378));
    layer5_outputs(2515) <= (layer4_outputs(1629)) and not (layer4_outputs(1621));
    layer5_outputs(2516) <= not(layer4_outputs(405));
    layer5_outputs(2517) <= not(layer4_outputs(1180));
    layer5_outputs(2518) <= (layer4_outputs(420)) xor (layer4_outputs(28));
    layer5_outputs(2519) <= (layer4_outputs(2018)) and not (layer4_outputs(1947));
    layer5_outputs(2520) <= not(layer4_outputs(1638)) or (layer4_outputs(901));
    layer5_outputs(2521) <= '1';
    layer5_outputs(2522) <= layer4_outputs(1314);
    layer5_outputs(2523) <= not((layer4_outputs(1636)) and (layer4_outputs(1814)));
    layer5_outputs(2524) <= layer4_outputs(2035);
    layer5_outputs(2525) <= (layer4_outputs(2332)) and (layer4_outputs(1943));
    layer5_outputs(2526) <= not(layer4_outputs(1089));
    layer5_outputs(2527) <= layer4_outputs(470);
    layer5_outputs(2528) <= not(layer4_outputs(2422));
    layer5_outputs(2529) <= '0';
    layer5_outputs(2530) <= not(layer4_outputs(861));
    layer5_outputs(2531) <= not(layer4_outputs(1481));
    layer5_outputs(2532) <= layer4_outputs(134);
    layer5_outputs(2533) <= not(layer4_outputs(1517)) or (layer4_outputs(1354));
    layer5_outputs(2534) <= not((layer4_outputs(179)) and (layer4_outputs(2036)));
    layer5_outputs(2535) <= not(layer4_outputs(2250));
    layer5_outputs(2536) <= '1';
    layer5_outputs(2537) <= '0';
    layer5_outputs(2538) <= (layer4_outputs(469)) and (layer4_outputs(380));
    layer5_outputs(2539) <= (layer4_outputs(664)) and not (layer4_outputs(472));
    layer5_outputs(2540) <= not(layer4_outputs(524));
    layer5_outputs(2541) <= (layer4_outputs(1898)) xor (layer4_outputs(1364));
    layer5_outputs(2542) <= layer4_outputs(2338);
    layer5_outputs(2543) <= layer4_outputs(222);
    layer5_outputs(2544) <= (layer4_outputs(1353)) and not (layer4_outputs(855));
    layer5_outputs(2545) <= layer4_outputs(642);
    layer5_outputs(2546) <= (layer4_outputs(2529)) or (layer4_outputs(1773));
    layer5_outputs(2547) <= not(layer4_outputs(1769));
    layer5_outputs(2548) <= not((layer4_outputs(1713)) and (layer4_outputs(592)));
    layer5_outputs(2549) <= (layer4_outputs(902)) and not (layer4_outputs(78));
    layer5_outputs(2550) <= not(layer4_outputs(2304));
    layer5_outputs(2551) <= not(layer4_outputs(283));
    layer5_outputs(2552) <= (layer4_outputs(1561)) and not (layer4_outputs(1462));
    layer5_outputs(2553) <= not((layer4_outputs(1476)) and (layer4_outputs(1543)));
    layer5_outputs(2554) <= (layer4_outputs(2482)) or (layer4_outputs(1786));
    layer5_outputs(2555) <= not(layer4_outputs(2191));
    layer5_outputs(2556) <= (layer4_outputs(992)) or (layer4_outputs(634));
    layer5_outputs(2557) <= layer4_outputs(2404);
    layer5_outputs(2558) <= layer4_outputs(474);
    layer5_outputs(2559) <= not(layer4_outputs(1286));
    layer6_outputs(0) <= not(layer5_outputs(1079));
    layer6_outputs(1) <= layer5_outputs(367);
    layer6_outputs(2) <= not(layer5_outputs(706));
    layer6_outputs(3) <= not((layer5_outputs(2068)) or (layer5_outputs(1490)));
    layer6_outputs(4) <= not((layer5_outputs(1278)) or (layer5_outputs(313)));
    layer6_outputs(5) <= not((layer5_outputs(724)) xor (layer5_outputs(2407)));
    layer6_outputs(6) <= layer5_outputs(139);
    layer6_outputs(7) <= not((layer5_outputs(1324)) xor (layer5_outputs(81)));
    layer6_outputs(8) <= not((layer5_outputs(745)) and (layer5_outputs(493)));
    layer6_outputs(9) <= not(layer5_outputs(1966));
    layer6_outputs(10) <= layer5_outputs(568);
    layer6_outputs(11) <= not((layer5_outputs(652)) and (layer5_outputs(1154)));
    layer6_outputs(12) <= layer5_outputs(581);
    layer6_outputs(13) <= not((layer5_outputs(1936)) xor (layer5_outputs(1324)));
    layer6_outputs(14) <= (layer5_outputs(217)) xor (layer5_outputs(343));
    layer6_outputs(15) <= not((layer5_outputs(233)) xor (layer5_outputs(442)));
    layer6_outputs(16) <= not(layer5_outputs(2313));
    layer6_outputs(17) <= not(layer5_outputs(1942));
    layer6_outputs(18) <= not((layer5_outputs(1789)) or (layer5_outputs(536)));
    layer6_outputs(19) <= not(layer5_outputs(306));
    layer6_outputs(20) <= (layer5_outputs(2541)) or (layer5_outputs(2280));
    layer6_outputs(21) <= layer5_outputs(1868);
    layer6_outputs(22) <= (layer5_outputs(1757)) and (layer5_outputs(30));
    layer6_outputs(23) <= not(layer5_outputs(1341));
    layer6_outputs(24) <= layer5_outputs(1437);
    layer6_outputs(25) <= layer5_outputs(868);
    layer6_outputs(26) <= not(layer5_outputs(2287));
    layer6_outputs(27) <= not(layer5_outputs(569));
    layer6_outputs(28) <= layer5_outputs(1317);
    layer6_outputs(29) <= layer5_outputs(394);
    layer6_outputs(30) <= (layer5_outputs(981)) xor (layer5_outputs(1925));
    layer6_outputs(31) <= (layer5_outputs(1693)) and (layer5_outputs(2147));
    layer6_outputs(32) <= '0';
    layer6_outputs(33) <= not(layer5_outputs(220));
    layer6_outputs(34) <= not(layer5_outputs(1209));
    layer6_outputs(35) <= not(layer5_outputs(1584));
    layer6_outputs(36) <= layer5_outputs(1261);
    layer6_outputs(37) <= not(layer5_outputs(112));
    layer6_outputs(38) <= not(layer5_outputs(9));
    layer6_outputs(39) <= layer5_outputs(2325);
    layer6_outputs(40) <= layer5_outputs(316);
    layer6_outputs(41) <= (layer5_outputs(635)) and not (layer5_outputs(348));
    layer6_outputs(42) <= (layer5_outputs(1436)) or (layer5_outputs(856));
    layer6_outputs(43) <= (layer5_outputs(1098)) xor (layer5_outputs(1737));
    layer6_outputs(44) <= (layer5_outputs(667)) and not (layer5_outputs(762));
    layer6_outputs(45) <= layer5_outputs(2433);
    layer6_outputs(46) <= not(layer5_outputs(1291)) or (layer5_outputs(1593));
    layer6_outputs(47) <= not(layer5_outputs(626));
    layer6_outputs(48) <= not(layer5_outputs(2482));
    layer6_outputs(49) <= layer5_outputs(1348);
    layer6_outputs(50) <= (layer5_outputs(1714)) xor (layer5_outputs(926));
    layer6_outputs(51) <= layer5_outputs(914);
    layer6_outputs(52) <= not(layer5_outputs(1156));
    layer6_outputs(53) <= layer5_outputs(474);
    layer6_outputs(54) <= not(layer5_outputs(42));
    layer6_outputs(55) <= layer5_outputs(636);
    layer6_outputs(56) <= (layer5_outputs(615)) or (layer5_outputs(423));
    layer6_outputs(57) <= layer5_outputs(2048);
    layer6_outputs(58) <= not(layer5_outputs(1731));
    layer6_outputs(59) <= layer5_outputs(1945);
    layer6_outputs(60) <= not((layer5_outputs(2260)) xor (layer5_outputs(1100)));
    layer6_outputs(61) <= (layer5_outputs(1361)) and not (layer5_outputs(814));
    layer6_outputs(62) <= (layer5_outputs(1353)) and (layer5_outputs(428));
    layer6_outputs(63) <= not((layer5_outputs(690)) xor (layer5_outputs(1606)));
    layer6_outputs(64) <= (layer5_outputs(1577)) and not (layer5_outputs(1318));
    layer6_outputs(65) <= not(layer5_outputs(383)) or (layer5_outputs(29));
    layer6_outputs(66) <= (layer5_outputs(2269)) and not (layer5_outputs(1401));
    layer6_outputs(67) <= (layer5_outputs(1387)) and not (layer5_outputs(2298));
    layer6_outputs(68) <= not(layer5_outputs(906));
    layer6_outputs(69) <= not(layer5_outputs(1007));
    layer6_outputs(70) <= not(layer5_outputs(2239));
    layer6_outputs(71) <= (layer5_outputs(1792)) and (layer5_outputs(1395));
    layer6_outputs(72) <= layer5_outputs(468);
    layer6_outputs(73) <= layer5_outputs(647);
    layer6_outputs(74) <= not(layer5_outputs(140));
    layer6_outputs(75) <= not((layer5_outputs(1991)) and (layer5_outputs(1947)));
    layer6_outputs(76) <= layer5_outputs(341);
    layer6_outputs(77) <= layer5_outputs(1928);
    layer6_outputs(78) <= not(layer5_outputs(425)) or (layer5_outputs(307));
    layer6_outputs(79) <= not((layer5_outputs(1068)) and (layer5_outputs(2458)));
    layer6_outputs(80) <= (layer5_outputs(240)) or (layer5_outputs(268));
    layer6_outputs(81) <= not(layer5_outputs(1653));
    layer6_outputs(82) <= layer5_outputs(1333);
    layer6_outputs(83) <= not((layer5_outputs(2421)) or (layer5_outputs(956)));
    layer6_outputs(84) <= not(layer5_outputs(909)) or (layer5_outputs(2054));
    layer6_outputs(85) <= layer5_outputs(189);
    layer6_outputs(86) <= not(layer5_outputs(22));
    layer6_outputs(87) <= not(layer5_outputs(1235));
    layer6_outputs(88) <= (layer5_outputs(1529)) xor (layer5_outputs(255));
    layer6_outputs(89) <= layer5_outputs(672);
    layer6_outputs(90) <= layer5_outputs(2178);
    layer6_outputs(91) <= not((layer5_outputs(5)) xor (layer5_outputs(807)));
    layer6_outputs(92) <= (layer5_outputs(2219)) or (layer5_outputs(527));
    layer6_outputs(93) <= not((layer5_outputs(1559)) or (layer5_outputs(424)));
    layer6_outputs(94) <= not((layer5_outputs(1968)) xor (layer5_outputs(1865)));
    layer6_outputs(95) <= not((layer5_outputs(202)) and (layer5_outputs(1950)));
    layer6_outputs(96) <= not(layer5_outputs(1163));
    layer6_outputs(97) <= not(layer5_outputs(1749));
    layer6_outputs(98) <= (layer5_outputs(1544)) or (layer5_outputs(2411));
    layer6_outputs(99) <= not(layer5_outputs(2068)) or (layer5_outputs(234));
    layer6_outputs(100) <= (layer5_outputs(2454)) or (layer5_outputs(2128));
    layer6_outputs(101) <= (layer5_outputs(731)) and not (layer5_outputs(35));
    layer6_outputs(102) <= (layer5_outputs(1448)) and not (layer5_outputs(413));
    layer6_outputs(103) <= not(layer5_outputs(358));
    layer6_outputs(104) <= layer5_outputs(1646);
    layer6_outputs(105) <= layer5_outputs(209);
    layer6_outputs(106) <= '1';
    layer6_outputs(107) <= not((layer5_outputs(1927)) xor (layer5_outputs(169)));
    layer6_outputs(108) <= not((layer5_outputs(1878)) or (layer5_outputs(2334)));
    layer6_outputs(109) <= '1';
    layer6_outputs(110) <= (layer5_outputs(1666)) and not (layer5_outputs(2229));
    layer6_outputs(111) <= not((layer5_outputs(1957)) and (layer5_outputs(1935)));
    layer6_outputs(112) <= not((layer5_outputs(2011)) or (layer5_outputs(1701)));
    layer6_outputs(113) <= layer5_outputs(1959);
    layer6_outputs(114) <= (layer5_outputs(200)) and not (layer5_outputs(1679));
    layer6_outputs(115) <= not((layer5_outputs(1752)) or (layer5_outputs(1046)));
    layer6_outputs(116) <= not(layer5_outputs(976));
    layer6_outputs(117) <= not((layer5_outputs(1673)) or (layer5_outputs(899)));
    layer6_outputs(118) <= not(layer5_outputs(1434));
    layer6_outputs(119) <= layer5_outputs(2333);
    layer6_outputs(120) <= not(layer5_outputs(159));
    layer6_outputs(121) <= layer5_outputs(2276);
    layer6_outputs(122) <= layer5_outputs(421);
    layer6_outputs(123) <= not((layer5_outputs(2154)) or (layer5_outputs(2216)));
    layer6_outputs(124) <= not((layer5_outputs(730)) or (layer5_outputs(2149)));
    layer6_outputs(125) <= layer5_outputs(1900);
    layer6_outputs(126) <= (layer5_outputs(973)) xor (layer5_outputs(1262));
    layer6_outputs(127) <= layer5_outputs(85);
    layer6_outputs(128) <= not(layer5_outputs(1088));
    layer6_outputs(129) <= (layer5_outputs(1334)) and not (layer5_outputs(2394));
    layer6_outputs(130) <= not(layer5_outputs(2151));
    layer6_outputs(131) <= not((layer5_outputs(2015)) or (layer5_outputs(9)));
    layer6_outputs(132) <= layer5_outputs(1662);
    layer6_outputs(133) <= not((layer5_outputs(2311)) or (layer5_outputs(2372)));
    layer6_outputs(134) <= not(layer5_outputs(1476));
    layer6_outputs(135) <= not(layer5_outputs(364));
    layer6_outputs(136) <= not(layer5_outputs(2376));
    layer6_outputs(137) <= layer5_outputs(937);
    layer6_outputs(138) <= layer5_outputs(2468);
    layer6_outputs(139) <= not(layer5_outputs(930)) or (layer5_outputs(951));
    layer6_outputs(140) <= not((layer5_outputs(198)) and (layer5_outputs(680)));
    layer6_outputs(141) <= not(layer5_outputs(824)) or (layer5_outputs(484));
    layer6_outputs(142) <= '0';
    layer6_outputs(143) <= not((layer5_outputs(1796)) xor (layer5_outputs(1953)));
    layer6_outputs(144) <= not(layer5_outputs(1637));
    layer6_outputs(145) <= layer5_outputs(1600);
    layer6_outputs(146) <= not(layer5_outputs(1379));
    layer6_outputs(147) <= layer5_outputs(827);
    layer6_outputs(148) <= not(layer5_outputs(1946));
    layer6_outputs(149) <= (layer5_outputs(2160)) xor (layer5_outputs(2165));
    layer6_outputs(150) <= '1';
    layer6_outputs(151) <= layer5_outputs(654);
    layer6_outputs(152) <= layer5_outputs(1395);
    layer6_outputs(153) <= not(layer5_outputs(1501));
    layer6_outputs(154) <= (layer5_outputs(715)) xor (layer5_outputs(1380));
    layer6_outputs(155) <= not(layer5_outputs(1810)) or (layer5_outputs(498));
    layer6_outputs(156) <= not((layer5_outputs(259)) and (layer5_outputs(1336)));
    layer6_outputs(157) <= (layer5_outputs(2008)) and (layer5_outputs(1379));
    layer6_outputs(158) <= layer5_outputs(1977);
    layer6_outputs(159) <= (layer5_outputs(1739)) xor (layer5_outputs(2397));
    layer6_outputs(160) <= not(layer5_outputs(1399));
    layer6_outputs(161) <= (layer5_outputs(1447)) xor (layer5_outputs(2136));
    layer6_outputs(162) <= layer5_outputs(357);
    layer6_outputs(163) <= not(layer5_outputs(894));
    layer6_outputs(164) <= layer5_outputs(1958);
    layer6_outputs(165) <= not((layer5_outputs(988)) or (layer5_outputs(1954)));
    layer6_outputs(166) <= not((layer5_outputs(1196)) and (layer5_outputs(296)));
    layer6_outputs(167) <= not(layer5_outputs(1370)) or (layer5_outputs(45));
    layer6_outputs(168) <= not(layer5_outputs(2379));
    layer6_outputs(169) <= not(layer5_outputs(1463));
    layer6_outputs(170) <= not(layer5_outputs(1742)) or (layer5_outputs(152));
    layer6_outputs(171) <= layer5_outputs(891);
    layer6_outputs(172) <= layer5_outputs(2486);
    layer6_outputs(173) <= layer5_outputs(1968);
    layer6_outputs(174) <= not(layer5_outputs(33)) or (layer5_outputs(471));
    layer6_outputs(175) <= not(layer5_outputs(27));
    layer6_outputs(176) <= not(layer5_outputs(852));
    layer6_outputs(177) <= layer5_outputs(1017);
    layer6_outputs(178) <= not(layer5_outputs(500)) or (layer5_outputs(2225));
    layer6_outputs(179) <= not(layer5_outputs(1848)) or (layer5_outputs(1630));
    layer6_outputs(180) <= not(layer5_outputs(1333));
    layer6_outputs(181) <= not((layer5_outputs(115)) and (layer5_outputs(1841)));
    layer6_outputs(182) <= layer5_outputs(1467);
    layer6_outputs(183) <= layer5_outputs(1518);
    layer6_outputs(184) <= layer5_outputs(278);
    layer6_outputs(185) <= '1';
    layer6_outputs(186) <= not(layer5_outputs(1369));
    layer6_outputs(187) <= not(layer5_outputs(1309));
    layer6_outputs(188) <= layer5_outputs(25);
    layer6_outputs(189) <= not(layer5_outputs(2328));
    layer6_outputs(190) <= (layer5_outputs(1085)) and not (layer5_outputs(644));
    layer6_outputs(191) <= not(layer5_outputs(1661));
    layer6_outputs(192) <= (layer5_outputs(315)) and (layer5_outputs(2488));
    layer6_outputs(193) <= (layer5_outputs(2099)) and not (layer5_outputs(1617));
    layer6_outputs(194) <= layer5_outputs(686);
    layer6_outputs(195) <= (layer5_outputs(2100)) and not (layer5_outputs(2341));
    layer6_outputs(196) <= not(layer5_outputs(1095));
    layer6_outputs(197) <= (layer5_outputs(1199)) xor (layer5_outputs(2505));
    layer6_outputs(198) <= not(layer5_outputs(2152)) or (layer5_outputs(2401));
    layer6_outputs(199) <= not(layer5_outputs(676));
    layer6_outputs(200) <= (layer5_outputs(1283)) or (layer5_outputs(726));
    layer6_outputs(201) <= not(layer5_outputs(1740));
    layer6_outputs(202) <= layer5_outputs(2018);
    layer6_outputs(203) <= layer5_outputs(1800);
    layer6_outputs(204) <= layer5_outputs(2537);
    layer6_outputs(205) <= not(layer5_outputs(553)) or (layer5_outputs(2174));
    layer6_outputs(206) <= not((layer5_outputs(479)) or (layer5_outputs(870)));
    layer6_outputs(207) <= not(layer5_outputs(520));
    layer6_outputs(208) <= (layer5_outputs(652)) and (layer5_outputs(2464));
    layer6_outputs(209) <= not((layer5_outputs(2348)) xor (layer5_outputs(2347)));
    layer6_outputs(210) <= not(layer5_outputs(1354)) or (layer5_outputs(2455));
    layer6_outputs(211) <= layer5_outputs(1795);
    layer6_outputs(212) <= not(layer5_outputs(812));
    layer6_outputs(213) <= not(layer5_outputs(927));
    layer6_outputs(214) <= not((layer5_outputs(335)) and (layer5_outputs(2405)));
    layer6_outputs(215) <= (layer5_outputs(2167)) and not (layer5_outputs(800));
    layer6_outputs(216) <= not((layer5_outputs(1819)) xor (layer5_outputs(365)));
    layer6_outputs(217) <= layer5_outputs(2548);
    layer6_outputs(218) <= not(layer5_outputs(1280));
    layer6_outputs(219) <= not((layer5_outputs(1059)) or (layer5_outputs(330)));
    layer6_outputs(220) <= not(layer5_outputs(2032));
    layer6_outputs(221) <= not(layer5_outputs(804));
    layer6_outputs(222) <= not(layer5_outputs(330));
    layer6_outputs(223) <= layer5_outputs(1946);
    layer6_outputs(224) <= (layer5_outputs(2277)) xor (layer5_outputs(314));
    layer6_outputs(225) <= not(layer5_outputs(863));
    layer6_outputs(226) <= layer5_outputs(1543);
    layer6_outputs(227) <= layer5_outputs(462);
    layer6_outputs(228) <= layer5_outputs(674);
    layer6_outputs(229) <= (layer5_outputs(2461)) and not (layer5_outputs(1678));
    layer6_outputs(230) <= not(layer5_outputs(1815));
    layer6_outputs(231) <= not(layer5_outputs(1643));
    layer6_outputs(232) <= (layer5_outputs(1256)) xor (layer5_outputs(503));
    layer6_outputs(233) <= not(layer5_outputs(2439)) or (layer5_outputs(975));
    layer6_outputs(234) <= (layer5_outputs(2022)) and not (layer5_outputs(1276));
    layer6_outputs(235) <= not(layer5_outputs(1076));
    layer6_outputs(236) <= not((layer5_outputs(1722)) and (layer5_outputs(1336)));
    layer6_outputs(237) <= not(layer5_outputs(1411));
    layer6_outputs(238) <= (layer5_outputs(532)) and (layer5_outputs(1813));
    layer6_outputs(239) <= layer5_outputs(324);
    layer6_outputs(240) <= not((layer5_outputs(130)) xor (layer5_outputs(403)));
    layer6_outputs(241) <= not((layer5_outputs(2492)) xor (layer5_outputs(2017)));
    layer6_outputs(242) <= layer5_outputs(2406);
    layer6_outputs(243) <= layer5_outputs(2255);
    layer6_outputs(244) <= not(layer5_outputs(1307)) or (layer5_outputs(2389));
    layer6_outputs(245) <= not(layer5_outputs(1328));
    layer6_outputs(246) <= not(layer5_outputs(641));
    layer6_outputs(247) <= not(layer5_outputs(1383));
    layer6_outputs(248) <= layer5_outputs(203);
    layer6_outputs(249) <= not(layer5_outputs(1866));
    layer6_outputs(250) <= not(layer5_outputs(743));
    layer6_outputs(251) <= layer5_outputs(287);
    layer6_outputs(252) <= not(layer5_outputs(1104)) or (layer5_outputs(1073));
    layer6_outputs(253) <= (layer5_outputs(38)) or (layer5_outputs(1057));
    layer6_outputs(254) <= (layer5_outputs(1686)) and (layer5_outputs(1313));
    layer6_outputs(255) <= not(layer5_outputs(1061));
    layer6_outputs(256) <= layer5_outputs(625);
    layer6_outputs(257) <= not(layer5_outputs(709)) or (layer5_outputs(63));
    layer6_outputs(258) <= (layer5_outputs(954)) xor (layer5_outputs(221));
    layer6_outputs(259) <= layer5_outputs(2150);
    layer6_outputs(260) <= not(layer5_outputs(1963));
    layer6_outputs(261) <= not(layer5_outputs(2396)) or (layer5_outputs(433));
    layer6_outputs(262) <= layer5_outputs(262);
    layer6_outputs(263) <= (layer5_outputs(874)) xor (layer5_outputs(1164));
    layer6_outputs(264) <= layer5_outputs(2516);
    layer6_outputs(265) <= not(layer5_outputs(2130)) or (layer5_outputs(85));
    layer6_outputs(266) <= (layer5_outputs(2304)) xor (layer5_outputs(2061));
    layer6_outputs(267) <= layer5_outputs(1203);
    layer6_outputs(268) <= layer5_outputs(942);
    layer6_outputs(269) <= layer5_outputs(390);
    layer6_outputs(270) <= not(layer5_outputs(510)) or (layer5_outputs(2162));
    layer6_outputs(271) <= not((layer5_outputs(623)) xor (layer5_outputs(1314)));
    layer6_outputs(272) <= not((layer5_outputs(40)) and (layer5_outputs(714)));
    layer6_outputs(273) <= layer5_outputs(1826);
    layer6_outputs(274) <= layer5_outputs(1364);
    layer6_outputs(275) <= layer5_outputs(2006);
    layer6_outputs(276) <= layer5_outputs(1368);
    layer6_outputs(277) <= not(layer5_outputs(295));
    layer6_outputs(278) <= (layer5_outputs(1611)) and (layer5_outputs(348));
    layer6_outputs(279) <= (layer5_outputs(1694)) xor (layer5_outputs(1233));
    layer6_outputs(280) <= not((layer5_outputs(760)) or (layer5_outputs(1186)));
    layer6_outputs(281) <= layer5_outputs(2228);
    layer6_outputs(282) <= (layer5_outputs(1035)) and not (layer5_outputs(1517));
    layer6_outputs(283) <= not(layer5_outputs(1883));
    layer6_outputs(284) <= not(layer5_outputs(736));
    layer6_outputs(285) <= not((layer5_outputs(1028)) xor (layer5_outputs(395)));
    layer6_outputs(286) <= layer5_outputs(2210);
    layer6_outputs(287) <= layer5_outputs(1149);
    layer6_outputs(288) <= not(layer5_outputs(2413));
    layer6_outputs(289) <= (layer5_outputs(1916)) or (layer5_outputs(966));
    layer6_outputs(290) <= layer5_outputs(1009);
    layer6_outputs(291) <= not(layer5_outputs(1660));
    layer6_outputs(292) <= not(layer5_outputs(962));
    layer6_outputs(293) <= not(layer5_outputs(468));
    layer6_outputs(294) <= not((layer5_outputs(825)) xor (layer5_outputs(1562)));
    layer6_outputs(295) <= layer5_outputs(936);
    layer6_outputs(296) <= not((layer5_outputs(1525)) and (layer5_outputs(2257)));
    layer6_outputs(297) <= layer5_outputs(1554);
    layer6_outputs(298) <= layer5_outputs(1103);
    layer6_outputs(299) <= not((layer5_outputs(1432)) or (layer5_outputs(2448)));
    layer6_outputs(300) <= not(layer5_outputs(2089));
    layer6_outputs(301) <= not((layer5_outputs(1414)) or (layer5_outputs(518)));
    layer6_outputs(302) <= layer5_outputs(1725);
    layer6_outputs(303) <= not(layer5_outputs(1281));
    layer6_outputs(304) <= not(layer5_outputs(296)) or (layer5_outputs(786));
    layer6_outputs(305) <= layer5_outputs(1909);
    layer6_outputs(306) <= layer5_outputs(986);
    layer6_outputs(307) <= not(layer5_outputs(402)) or (layer5_outputs(190));
    layer6_outputs(308) <= layer5_outputs(1522);
    layer6_outputs(309) <= (layer5_outputs(2461)) xor (layer5_outputs(341));
    layer6_outputs(310) <= not(layer5_outputs(1903));
    layer6_outputs(311) <= layer5_outputs(1555);
    layer6_outputs(312) <= not((layer5_outputs(822)) xor (layer5_outputs(1696)));
    layer6_outputs(313) <= layer5_outputs(2063);
    layer6_outputs(314) <= (layer5_outputs(274)) and not (layer5_outputs(2048));
    layer6_outputs(315) <= (layer5_outputs(1377)) xor (layer5_outputs(2140));
    layer6_outputs(316) <= not(layer5_outputs(1015)) or (layer5_outputs(907));
    layer6_outputs(317) <= not(layer5_outputs(116));
    layer6_outputs(318) <= not(layer5_outputs(2488)) or (layer5_outputs(1133));
    layer6_outputs(319) <= (layer5_outputs(1654)) and (layer5_outputs(292));
    layer6_outputs(320) <= layer5_outputs(1309);
    layer6_outputs(321) <= '0';
    layer6_outputs(322) <= not(layer5_outputs(276));
    layer6_outputs(323) <= not((layer5_outputs(1510)) and (layer5_outputs(2343)));
    layer6_outputs(324) <= not(layer5_outputs(1523));
    layer6_outputs(325) <= not((layer5_outputs(470)) xor (layer5_outputs(2183)));
    layer6_outputs(326) <= not(layer5_outputs(108)) or (layer5_outputs(364));
    layer6_outputs(327) <= layer5_outputs(165);
    layer6_outputs(328) <= layer5_outputs(2024);
    layer6_outputs(329) <= layer5_outputs(1222);
    layer6_outputs(330) <= layer5_outputs(2100);
    layer6_outputs(331) <= not((layer5_outputs(1948)) and (layer5_outputs(2405)));
    layer6_outputs(332) <= not(layer5_outputs(215));
    layer6_outputs(333) <= layer5_outputs(1846);
    layer6_outputs(334) <= layer5_outputs(707);
    layer6_outputs(335) <= layer5_outputs(107);
    layer6_outputs(336) <= layer5_outputs(49);
    layer6_outputs(337) <= (layer5_outputs(357)) or (layer5_outputs(1121));
    layer6_outputs(338) <= (layer5_outputs(2115)) and not (layer5_outputs(1855));
    layer6_outputs(339) <= layer5_outputs(1265);
    layer6_outputs(340) <= layer5_outputs(1443);
    layer6_outputs(341) <= not((layer5_outputs(1790)) xor (layer5_outputs(1650)));
    layer6_outputs(342) <= (layer5_outputs(2080)) and (layer5_outputs(1873));
    layer6_outputs(343) <= (layer5_outputs(1710)) and not (layer5_outputs(333));
    layer6_outputs(344) <= (layer5_outputs(1638)) and not (layer5_outputs(737));
    layer6_outputs(345) <= not(layer5_outputs(1955));
    layer6_outputs(346) <= not((layer5_outputs(2244)) xor (layer5_outputs(31)));
    layer6_outputs(347) <= not(layer5_outputs(621));
    layer6_outputs(348) <= not(layer5_outputs(1360));
    layer6_outputs(349) <= layer5_outputs(177);
    layer6_outputs(350) <= layer5_outputs(19);
    layer6_outputs(351) <= (layer5_outputs(1921)) and not (layer5_outputs(1586));
    layer6_outputs(352) <= (layer5_outputs(1725)) or (layer5_outputs(1298));
    layer6_outputs(353) <= not((layer5_outputs(1847)) xor (layer5_outputs(1041)));
    layer6_outputs(354) <= not(layer5_outputs(351)) or (layer5_outputs(566));
    layer6_outputs(355) <= (layer5_outputs(2530)) and not (layer5_outputs(172));
    layer6_outputs(356) <= not((layer5_outputs(933)) and (layer5_outputs(2367)));
    layer6_outputs(357) <= layer5_outputs(875);
    layer6_outputs(358) <= layer5_outputs(1086);
    layer6_outputs(359) <= not(layer5_outputs(1468)) or (layer5_outputs(888));
    layer6_outputs(360) <= layer5_outputs(2045);
    layer6_outputs(361) <= (layer5_outputs(1269)) and not (layer5_outputs(2440));
    layer6_outputs(362) <= not(layer5_outputs(1667));
    layer6_outputs(363) <= layer5_outputs(1619);
    layer6_outputs(364) <= not((layer5_outputs(1190)) or (layer5_outputs(1784)));
    layer6_outputs(365) <= layer5_outputs(323);
    layer6_outputs(366) <= layer5_outputs(1072);
    layer6_outputs(367) <= (layer5_outputs(1264)) or (layer5_outputs(1636));
    layer6_outputs(368) <= layer5_outputs(2147);
    layer6_outputs(369) <= not(layer5_outputs(2393));
    layer6_outputs(370) <= not(layer5_outputs(315));
    layer6_outputs(371) <= not(layer5_outputs(1203));
    layer6_outputs(372) <= not(layer5_outputs(1471)) or (layer5_outputs(1213));
    layer6_outputs(373) <= layer5_outputs(2312);
    layer6_outputs(374) <= layer5_outputs(900);
    layer6_outputs(375) <= layer5_outputs(234);
    layer6_outputs(376) <= (layer5_outputs(2515)) xor (layer5_outputs(452));
    layer6_outputs(377) <= layer5_outputs(2145);
    layer6_outputs(378) <= not(layer5_outputs(431)) or (layer5_outputs(2113));
    layer6_outputs(379) <= not(layer5_outputs(1181));
    layer6_outputs(380) <= (layer5_outputs(1964)) and not (layer5_outputs(461));
    layer6_outputs(381) <= layer5_outputs(940);
    layer6_outputs(382) <= not((layer5_outputs(1393)) and (layer5_outputs(1268)));
    layer6_outputs(383) <= (layer5_outputs(486)) and (layer5_outputs(1285));
    layer6_outputs(384) <= not(layer5_outputs(1665));
    layer6_outputs(385) <= not((layer5_outputs(1453)) and (layer5_outputs(885)));
    layer6_outputs(386) <= not(layer5_outputs(52));
    layer6_outputs(387) <= not(layer5_outputs(2399)) or (layer5_outputs(1721));
    layer6_outputs(388) <= (layer5_outputs(1350)) and not (layer5_outputs(220));
    layer6_outputs(389) <= not((layer5_outputs(1045)) or (layer5_outputs(1783)));
    layer6_outputs(390) <= (layer5_outputs(1469)) and (layer5_outputs(570));
    layer6_outputs(391) <= not(layer5_outputs(1514)) or (layer5_outputs(1400));
    layer6_outputs(392) <= layer5_outputs(19);
    layer6_outputs(393) <= (layer5_outputs(68)) xor (layer5_outputs(305));
    layer6_outputs(394) <= not(layer5_outputs(1431));
    layer6_outputs(395) <= layer5_outputs(1270);
    layer6_outputs(396) <= (layer5_outputs(735)) and not (layer5_outputs(2293));
    layer6_outputs(397) <= not(layer5_outputs(1864)) or (layer5_outputs(1983));
    layer6_outputs(398) <= '1';
    layer6_outputs(399) <= not(layer5_outputs(328));
    layer6_outputs(400) <= not((layer5_outputs(2056)) xor (layer5_outputs(1805)));
    layer6_outputs(401) <= layer5_outputs(1920);
    layer6_outputs(402) <= (layer5_outputs(65)) xor (layer5_outputs(213));
    layer6_outputs(403) <= not(layer5_outputs(1410)) or (layer5_outputs(2235));
    layer6_outputs(404) <= layer5_outputs(2115);
    layer6_outputs(405) <= layer5_outputs(788);
    layer6_outputs(406) <= not(layer5_outputs(64));
    layer6_outputs(407) <= layer5_outputs(293);
    layer6_outputs(408) <= (layer5_outputs(2009)) xor (layer5_outputs(258));
    layer6_outputs(409) <= not(layer5_outputs(1265)) or (layer5_outputs(1037));
    layer6_outputs(410) <= (layer5_outputs(1193)) and (layer5_outputs(1078));
    layer6_outputs(411) <= not(layer5_outputs(311));
    layer6_outputs(412) <= layer5_outputs(752);
    layer6_outputs(413) <= layer5_outputs(2500);
    layer6_outputs(414) <= layer5_outputs(255);
    layer6_outputs(415) <= layer5_outputs(484);
    layer6_outputs(416) <= layer5_outputs(2232);
    layer6_outputs(417) <= not((layer5_outputs(1202)) and (layer5_outputs(2424)));
    layer6_outputs(418) <= (layer5_outputs(2158)) or (layer5_outputs(733));
    layer6_outputs(419) <= (layer5_outputs(312)) and not (layer5_outputs(153));
    layer6_outputs(420) <= layer5_outputs(163);
    layer6_outputs(421) <= layer5_outputs(1380);
    layer6_outputs(422) <= (layer5_outputs(297)) or (layer5_outputs(2146));
    layer6_outputs(423) <= layer5_outputs(2556);
    layer6_outputs(424) <= not(layer5_outputs(41));
    layer6_outputs(425) <= layer5_outputs(1592);
    layer6_outputs(426) <= not(layer5_outputs(964));
    layer6_outputs(427) <= not(layer5_outputs(681));
    layer6_outputs(428) <= (layer5_outputs(1901)) xor (layer5_outputs(263));
    layer6_outputs(429) <= layer5_outputs(2508);
    layer6_outputs(430) <= (layer5_outputs(2448)) or (layer5_outputs(1327));
    layer6_outputs(431) <= layer5_outputs(2035);
    layer6_outputs(432) <= (layer5_outputs(2314)) or (layer5_outputs(1797));
    layer6_outputs(433) <= not(layer5_outputs(1892));
    layer6_outputs(434) <= layer5_outputs(2350);
    layer6_outputs(435) <= not(layer5_outputs(1274)) or (layer5_outputs(1857));
    layer6_outputs(436) <= not(layer5_outputs(131));
    layer6_outputs(437) <= not((layer5_outputs(1243)) xor (layer5_outputs(2052)));
    layer6_outputs(438) <= not(layer5_outputs(1322));
    layer6_outputs(439) <= layer5_outputs(784);
    layer6_outputs(440) <= not((layer5_outputs(1887)) and (layer5_outputs(1473)));
    layer6_outputs(441) <= layer5_outputs(2064);
    layer6_outputs(442) <= layer5_outputs(946);
    layer6_outputs(443) <= layer5_outputs(1403);
    layer6_outputs(444) <= layer5_outputs(1482);
    layer6_outputs(445) <= not(layer5_outputs(2028));
    layer6_outputs(446) <= (layer5_outputs(355)) or (layer5_outputs(648));
    layer6_outputs(447) <= layer5_outputs(1061);
    layer6_outputs(448) <= not((layer5_outputs(33)) or (layer5_outputs(859)));
    layer6_outputs(449) <= layer5_outputs(1806);
    layer6_outputs(450) <= (layer5_outputs(40)) and (layer5_outputs(2114));
    layer6_outputs(451) <= not((layer5_outputs(1569)) xor (layer5_outputs(1862)));
    layer6_outputs(452) <= not(layer5_outputs(1760));
    layer6_outputs(453) <= not(layer5_outputs(546));
    layer6_outputs(454) <= layer5_outputs(2351);
    layer6_outputs(455) <= '1';
    layer6_outputs(456) <= not((layer5_outputs(1587)) or (layer5_outputs(2094)));
    layer6_outputs(457) <= not((layer5_outputs(599)) xor (layer5_outputs(918)));
    layer6_outputs(458) <= layer5_outputs(15);
    layer6_outputs(459) <= (layer5_outputs(737)) xor (layer5_outputs(1049));
    layer6_outputs(460) <= layer5_outputs(602);
    layer6_outputs(461) <= not(layer5_outputs(576));
    layer6_outputs(462) <= not(layer5_outputs(1074)) or (layer5_outputs(257));
    layer6_outputs(463) <= not(layer5_outputs(2065));
    layer6_outputs(464) <= layer5_outputs(749);
    layer6_outputs(465) <= not(layer5_outputs(313)) or (layer5_outputs(197));
    layer6_outputs(466) <= layer5_outputs(1840);
    layer6_outputs(467) <= layer5_outputs(2148);
    layer6_outputs(468) <= layer5_outputs(614);
    layer6_outputs(469) <= not((layer5_outputs(279)) xor (layer5_outputs(2445)));
    layer6_outputs(470) <= not((layer5_outputs(1437)) xor (layer5_outputs(2315)));
    layer6_outputs(471) <= not((layer5_outputs(1751)) or (layer5_outputs(1779)));
    layer6_outputs(472) <= layer5_outputs(1563);
    layer6_outputs(473) <= layer5_outputs(2019);
    layer6_outputs(474) <= not(layer5_outputs(2189)) or (layer5_outputs(88));
    layer6_outputs(475) <= layer5_outputs(1398);
    layer6_outputs(476) <= (layer5_outputs(1694)) and not (layer5_outputs(285));
    layer6_outputs(477) <= (layer5_outputs(266)) and (layer5_outputs(1364));
    layer6_outputs(478) <= (layer5_outputs(1572)) and not (layer5_outputs(237));
    layer6_outputs(479) <= not(layer5_outputs(139));
    layer6_outputs(480) <= (layer5_outputs(2182)) and not (layer5_outputs(1465));
    layer6_outputs(481) <= layer5_outputs(2532);
    layer6_outputs(482) <= not(layer5_outputs(1914));
    layer6_outputs(483) <= not((layer5_outputs(370)) xor (layer5_outputs(1487)));
    layer6_outputs(484) <= not(layer5_outputs(211));
    layer6_outputs(485) <= not(layer5_outputs(76)) or (layer5_outputs(965));
    layer6_outputs(486) <= layer5_outputs(2234);
    layer6_outputs(487) <= (layer5_outputs(629)) xor (layer5_outputs(2368));
    layer6_outputs(488) <= not((layer5_outputs(2044)) xor (layer5_outputs(2206)));
    layer6_outputs(489) <= layer5_outputs(199);
    layer6_outputs(490) <= not((layer5_outputs(1632)) xor (layer5_outputs(1538)));
    layer6_outputs(491) <= (layer5_outputs(2549)) or (layer5_outputs(191));
    layer6_outputs(492) <= (layer5_outputs(1729)) and (layer5_outputs(883));
    layer6_outputs(493) <= not(layer5_outputs(1687));
    layer6_outputs(494) <= not(layer5_outputs(1627)) or (layer5_outputs(1581));
    layer6_outputs(495) <= not(layer5_outputs(243)) or (layer5_outputs(2132));
    layer6_outputs(496) <= not(layer5_outputs(1732)) or (layer5_outputs(424));
    layer6_outputs(497) <= not(layer5_outputs(2360));
    layer6_outputs(498) <= not(layer5_outputs(1669));
    layer6_outputs(499) <= not(layer5_outputs(984));
    layer6_outputs(500) <= not((layer5_outputs(28)) xor (layer5_outputs(490)));
    layer6_outputs(501) <= (layer5_outputs(2170)) xor (layer5_outputs(722));
    layer6_outputs(502) <= layer5_outputs(2231);
    layer6_outputs(503) <= not(layer5_outputs(134));
    layer6_outputs(504) <= layer5_outputs(1297);
    layer6_outputs(505) <= layer5_outputs(1724);
    layer6_outputs(506) <= not(layer5_outputs(685));
    layer6_outputs(507) <= (layer5_outputs(1240)) and not (layer5_outputs(1841));
    layer6_outputs(508) <= layer5_outputs(1554);
    layer6_outputs(509) <= layer5_outputs(1077);
    layer6_outputs(510) <= layer5_outputs(597);
    layer6_outputs(511) <= not(layer5_outputs(766)) or (layer5_outputs(117));
    layer6_outputs(512) <= not(layer5_outputs(277));
    layer6_outputs(513) <= not((layer5_outputs(403)) or (layer5_outputs(228)));
    layer6_outputs(514) <= not(layer5_outputs(2332));
    layer6_outputs(515) <= (layer5_outputs(1215)) xor (layer5_outputs(1455));
    layer6_outputs(516) <= not(layer5_outputs(275));
    layer6_outputs(517) <= not((layer5_outputs(1726)) and (layer5_outputs(1807)));
    layer6_outputs(518) <= (layer5_outputs(1050)) xor (layer5_outputs(372));
    layer6_outputs(519) <= not((layer5_outputs(433)) or (layer5_outputs(1847)));
    layer6_outputs(520) <= (layer5_outputs(1021)) xor (layer5_outputs(272));
    layer6_outputs(521) <= not(layer5_outputs(1459));
    layer6_outputs(522) <= not(layer5_outputs(133));
    layer6_outputs(523) <= not(layer5_outputs(1019));
    layer6_outputs(524) <= not(layer5_outputs(129));
    layer6_outputs(525) <= not(layer5_outputs(454));
    layer6_outputs(526) <= not(layer5_outputs(1412)) or (layer5_outputs(2408));
    layer6_outputs(527) <= not((layer5_outputs(290)) or (layer5_outputs(2305)));
    layer6_outputs(528) <= not(layer5_outputs(360));
    layer6_outputs(529) <= (layer5_outputs(1018)) and not (layer5_outputs(2087));
    layer6_outputs(530) <= (layer5_outputs(1808)) and not (layer5_outputs(1303));
    layer6_outputs(531) <= not(layer5_outputs(257)) or (layer5_outputs(1793));
    layer6_outputs(532) <= not(layer5_outputs(977));
    layer6_outputs(533) <= (layer5_outputs(1031)) and not (layer5_outputs(2369));
    layer6_outputs(534) <= (layer5_outputs(1488)) or (layer5_outputs(129));
    layer6_outputs(535) <= (layer5_outputs(204)) and not (layer5_outputs(794));
    layer6_outputs(536) <= (layer5_outputs(1106)) xor (layer5_outputs(1195));
    layer6_outputs(537) <= layer5_outputs(948);
    layer6_outputs(538) <= (layer5_outputs(455)) and not (layer5_outputs(1919));
    layer6_outputs(539) <= (layer5_outputs(1124)) and (layer5_outputs(705));
    layer6_outputs(540) <= not((layer5_outputs(2196)) xor (layer5_outputs(182)));
    layer6_outputs(541) <= not((layer5_outputs(1721)) xor (layer5_outputs(1233)));
    layer6_outputs(542) <= (layer5_outputs(822)) xor (layer5_outputs(354));
    layer6_outputs(543) <= '1';
    layer6_outputs(544) <= not(layer5_outputs(1896)) or (layer5_outputs(2344));
    layer6_outputs(545) <= not((layer5_outputs(344)) or (layer5_outputs(481)));
    layer6_outputs(546) <= (layer5_outputs(182)) or (layer5_outputs(2235));
    layer6_outputs(547) <= not(layer5_outputs(1076));
    layer6_outputs(548) <= not(layer5_outputs(663));
    layer6_outputs(549) <= not(layer5_outputs(241)) or (layer5_outputs(2297));
    layer6_outputs(550) <= not(layer5_outputs(1385));
    layer6_outputs(551) <= not(layer5_outputs(265));
    layer6_outputs(552) <= not((layer5_outputs(1251)) or (layer5_outputs(1695)));
    layer6_outputs(553) <= not(layer5_outputs(2107));
    layer6_outputs(554) <= layer5_outputs(333);
    layer6_outputs(555) <= layer5_outputs(2101);
    layer6_outputs(556) <= not(layer5_outputs(1005)) or (layer5_outputs(2415));
    layer6_outputs(557) <= (layer5_outputs(51)) and (layer5_outputs(1761));
    layer6_outputs(558) <= (layer5_outputs(289)) and not (layer5_outputs(1775));
    layer6_outputs(559) <= layer5_outputs(1766);
    layer6_outputs(560) <= not(layer5_outputs(1939)) or (layer5_outputs(458));
    layer6_outputs(561) <= not(layer5_outputs(1792));
    layer6_outputs(562) <= layer5_outputs(524);
    layer6_outputs(563) <= not(layer5_outputs(2320));
    layer6_outputs(564) <= not(layer5_outputs(894));
    layer6_outputs(565) <= (layer5_outputs(2191)) and (layer5_outputs(503));
    layer6_outputs(566) <= layer5_outputs(2133);
    layer6_outputs(567) <= not(layer5_outputs(2049)) or (layer5_outputs(1937));
    layer6_outputs(568) <= (layer5_outputs(824)) and not (layer5_outputs(875));
    layer6_outputs(569) <= '0';
    layer6_outputs(570) <= not(layer5_outputs(1071)) or (layer5_outputs(496));
    layer6_outputs(571) <= not((layer5_outputs(1929)) and (layer5_outputs(2490)));
    layer6_outputs(572) <= not(layer5_outputs(252));
    layer6_outputs(573) <= not(layer5_outputs(515));
    layer6_outputs(574) <= not(layer5_outputs(1303)) or (layer5_outputs(709));
    layer6_outputs(575) <= '0';
    layer6_outputs(576) <= layer5_outputs(2484);
    layer6_outputs(577) <= layer5_outputs(1244);
    layer6_outputs(578) <= not(layer5_outputs(142));
    layer6_outputs(579) <= not(layer5_outputs(741));
    layer6_outputs(580) <= (layer5_outputs(29)) and (layer5_outputs(1820));
    layer6_outputs(581) <= layer5_outputs(2351);
    layer6_outputs(582) <= not(layer5_outputs(785));
    layer6_outputs(583) <= not(layer5_outputs(99)) or (layer5_outputs(712));
    layer6_outputs(584) <= not(layer5_outputs(2104));
    layer6_outputs(585) <= not(layer5_outputs(201));
    layer6_outputs(586) <= not(layer5_outputs(2553));
    layer6_outputs(587) <= not((layer5_outputs(1347)) or (layer5_outputs(1533)));
    layer6_outputs(588) <= not(layer5_outputs(2355));
    layer6_outputs(589) <= (layer5_outputs(1537)) and not (layer5_outputs(681));
    layer6_outputs(590) <= not(layer5_outputs(610)) or (layer5_outputs(2433));
    layer6_outputs(591) <= not(layer5_outputs(939));
    layer6_outputs(592) <= not(layer5_outputs(508));
    layer6_outputs(593) <= (layer5_outputs(2513)) and (layer5_outputs(768));
    layer6_outputs(594) <= layer5_outputs(2353);
    layer6_outputs(595) <= layer5_outputs(608);
    layer6_outputs(596) <= not(layer5_outputs(651));
    layer6_outputs(597) <= not(layer5_outputs(1768)) or (layer5_outputs(1154));
    layer6_outputs(598) <= layer5_outputs(2168);
    layer6_outputs(599) <= layer5_outputs(1978);
    layer6_outputs(600) <= layer5_outputs(196);
    layer6_outputs(601) <= not(layer5_outputs(620));
    layer6_outputs(602) <= layer5_outputs(432);
    layer6_outputs(603) <= not(layer5_outputs(644));
    layer6_outputs(604) <= (layer5_outputs(2373)) or (layer5_outputs(550));
    layer6_outputs(605) <= not(layer5_outputs(2498));
    layer6_outputs(606) <= layer5_outputs(125);
    layer6_outputs(607) <= layer5_outputs(922);
    layer6_outputs(608) <= not(layer5_outputs(588));
    layer6_outputs(609) <= not(layer5_outputs(485));
    layer6_outputs(610) <= (layer5_outputs(1442)) xor (layer5_outputs(2303));
    layer6_outputs(611) <= (layer5_outputs(877)) and not (layer5_outputs(204));
    layer6_outputs(612) <= not(layer5_outputs(1897));
    layer6_outputs(613) <= not((layer5_outputs(1982)) xor (layer5_outputs(50)));
    layer6_outputs(614) <= not(layer5_outputs(904));
    layer6_outputs(615) <= not(layer5_outputs(2525)) or (layer5_outputs(693));
    layer6_outputs(616) <= not(layer5_outputs(393));
    layer6_outputs(617) <= layer5_outputs(471);
    layer6_outputs(618) <= layer5_outputs(1836);
    layer6_outputs(619) <= not(layer5_outputs(863)) or (layer5_outputs(1664));
    layer6_outputs(620) <= not(layer5_outputs(1375));
    layer6_outputs(621) <= layer5_outputs(1585);
    layer6_outputs(622) <= (layer5_outputs(645)) xor (layer5_outputs(1339));
    layer6_outputs(623) <= not(layer5_outputs(2338));
    layer6_outputs(624) <= layer5_outputs(476);
    layer6_outputs(625) <= layer5_outputs(102);
    layer6_outputs(626) <= not(layer5_outputs(972));
    layer6_outputs(627) <= layer5_outputs(1994);
    layer6_outputs(628) <= not(layer5_outputs(1139));
    layer6_outputs(629) <= not(layer5_outputs(1297));
    layer6_outputs(630) <= not(layer5_outputs(2181));
    layer6_outputs(631) <= not(layer5_outputs(1041)) or (layer5_outputs(207));
    layer6_outputs(632) <= not((layer5_outputs(478)) xor (layer5_outputs(2289)));
    layer6_outputs(633) <= layer5_outputs(2336);
    layer6_outputs(634) <= not(layer5_outputs(317));
    layer6_outputs(635) <= layer5_outputs(437);
    layer6_outputs(636) <= layer5_outputs(2045);
    layer6_outputs(637) <= (layer5_outputs(543)) and (layer5_outputs(714));
    layer6_outputs(638) <= not(layer5_outputs(2007));
    layer6_outputs(639) <= not(layer5_outputs(1682));
    layer6_outputs(640) <= layer5_outputs(861);
    layer6_outputs(641) <= not(layer5_outputs(1489)) or (layer5_outputs(1970));
    layer6_outputs(642) <= not(layer5_outputs(66));
    layer6_outputs(643) <= not(layer5_outputs(1030));
    layer6_outputs(644) <= not((layer5_outputs(167)) xor (layer5_outputs(2381)));
    layer6_outputs(645) <= (layer5_outputs(655)) and not (layer5_outputs(2281));
    layer6_outputs(646) <= layer5_outputs(2320);
    layer6_outputs(647) <= not(layer5_outputs(1647));
    layer6_outputs(648) <= (layer5_outputs(1556)) xor (layer5_outputs(622));
    layer6_outputs(649) <= layer5_outputs(2317);
    layer6_outputs(650) <= not(layer5_outputs(1286)) or (layer5_outputs(373));
    layer6_outputs(651) <= layer5_outputs(2158);
    layer6_outputs(652) <= (layer5_outputs(1279)) and (layer5_outputs(1288));
    layer6_outputs(653) <= layer5_outputs(841);
    layer6_outputs(654) <= layer5_outputs(1854);
    layer6_outputs(655) <= layer5_outputs(592);
    layer6_outputs(656) <= (layer5_outputs(1735)) and (layer5_outputs(1108));
    layer6_outputs(657) <= (layer5_outputs(2087)) or (layer5_outputs(69));
    layer6_outputs(658) <= layer5_outputs(2078);
    layer6_outputs(659) <= (layer5_outputs(1561)) and not (layer5_outputs(1845));
    layer6_outputs(660) <= not(layer5_outputs(1837)) or (layer5_outputs(799));
    layer6_outputs(661) <= not(layer5_outputs(1427)) or (layer5_outputs(557));
    layer6_outputs(662) <= (layer5_outputs(1880)) xor (layer5_outputs(1175));
    layer6_outputs(663) <= layer5_outputs(1318);
    layer6_outputs(664) <= not(layer5_outputs(1857));
    layer6_outputs(665) <= layer5_outputs(955);
    layer6_outputs(666) <= not(layer5_outputs(385));
    layer6_outputs(667) <= (layer5_outputs(527)) xor (layer5_outputs(2233));
    layer6_outputs(668) <= layer5_outputs(1931);
    layer6_outputs(669) <= not(layer5_outputs(2232));
    layer6_outputs(670) <= layer5_outputs(45);
    layer6_outputs(671) <= not((layer5_outputs(2457)) xor (layer5_outputs(282)));
    layer6_outputs(672) <= (layer5_outputs(2419)) and (layer5_outputs(2559));
    layer6_outputs(673) <= (layer5_outputs(2498)) and not (layer5_outputs(1973));
    layer6_outputs(674) <= '0';
    layer6_outputs(675) <= layer5_outputs(1645);
    layer6_outputs(676) <= not(layer5_outputs(1325));
    layer6_outputs(677) <= not((layer5_outputs(1279)) xor (layer5_outputs(73)));
    layer6_outputs(678) <= not((layer5_outputs(637)) and (layer5_outputs(743)));
    layer6_outputs(679) <= not(layer5_outputs(2102));
    layer6_outputs(680) <= not(layer5_outputs(2092));
    layer6_outputs(681) <= not((layer5_outputs(959)) or (layer5_outputs(2396)));
    layer6_outputs(682) <= layer5_outputs(1115);
    layer6_outputs(683) <= (layer5_outputs(1373)) or (layer5_outputs(2339));
    layer6_outputs(684) <= layer5_outputs(1995);
    layer6_outputs(685) <= (layer5_outputs(1590)) xor (layer5_outputs(1216));
    layer6_outputs(686) <= (layer5_outputs(1052)) and (layer5_outputs(2468));
    layer6_outputs(687) <= not((layer5_outputs(828)) and (layer5_outputs(2447)));
    layer6_outputs(688) <= not(layer5_outputs(1902)) or (layer5_outputs(642));
    layer6_outputs(689) <= not(layer5_outputs(402));
    layer6_outputs(690) <= not(layer5_outputs(1898));
    layer6_outputs(691) <= not(layer5_outputs(181));
    layer6_outputs(692) <= not(layer5_outputs(2539));
    layer6_outputs(693) <= (layer5_outputs(2381)) or (layer5_outputs(1166));
    layer6_outputs(694) <= not(layer5_outputs(2170)) or (layer5_outputs(810));
    layer6_outputs(695) <= (layer5_outputs(1494)) xor (layer5_outputs(588));
    layer6_outputs(696) <= (layer5_outputs(1350)) and (layer5_outputs(2538));
    layer6_outputs(697) <= (layer5_outputs(287)) or (layer5_outputs(2423));
    layer6_outputs(698) <= layer5_outputs(2554);
    layer6_outputs(699) <= layer5_outputs(766);
    layer6_outputs(700) <= '0';
    layer6_outputs(701) <= (layer5_outputs(1428)) or (layer5_outputs(998));
    layer6_outputs(702) <= (layer5_outputs(140)) xor (layer5_outputs(781));
    layer6_outputs(703) <= not((layer5_outputs(1252)) xor (layer5_outputs(2447)));
    layer6_outputs(704) <= not(layer5_outputs(2185));
    layer6_outputs(705) <= not(layer5_outputs(501));
    layer6_outputs(706) <= not(layer5_outputs(2253));
    layer6_outputs(707) <= layer5_outputs(393);
    layer6_outputs(708) <= not((layer5_outputs(1993)) and (layer5_outputs(2210)));
    layer6_outputs(709) <= not((layer5_outputs(2076)) xor (layer5_outputs(1136)));
    layer6_outputs(710) <= not((layer5_outputs(2416)) and (layer5_outputs(601)));
    layer6_outputs(711) <= (layer5_outputs(1659)) and (layer5_outputs(48));
    layer6_outputs(712) <= layer5_outputs(2117);
    layer6_outputs(713) <= layer5_outputs(1503);
    layer6_outputs(714) <= layer5_outputs(1722);
    layer6_outputs(715) <= not(layer5_outputs(718));
    layer6_outputs(716) <= not(layer5_outputs(2319)) or (layer5_outputs(260));
    layer6_outputs(717) <= not((layer5_outputs(1239)) xor (layer5_outputs(157)));
    layer6_outputs(718) <= not((layer5_outputs(862)) xor (layer5_outputs(1025)));
    layer6_outputs(719) <= not(layer5_outputs(2201)) or (layer5_outputs(1172));
    layer6_outputs(720) <= not((layer5_outputs(1347)) or (layer5_outputs(2227)));
    layer6_outputs(721) <= (layer5_outputs(715)) xor (layer5_outputs(1407));
    layer6_outputs(722) <= layer5_outputs(2009);
    layer6_outputs(723) <= not(layer5_outputs(1216));
    layer6_outputs(724) <= not(layer5_outputs(323));
    layer6_outputs(725) <= not((layer5_outputs(1248)) or (layer5_outputs(2110)));
    layer6_outputs(726) <= not(layer5_outputs(1386));
    layer6_outputs(727) <= layer5_outputs(301);
    layer6_outputs(728) <= layer5_outputs(2172);
    layer6_outputs(729) <= layer5_outputs(2033);
    layer6_outputs(730) <= (layer5_outputs(2467)) and not (layer5_outputs(1716));
    layer6_outputs(731) <= layer5_outputs(1992);
    layer6_outputs(732) <= not((layer5_outputs(249)) or (layer5_outputs(559)));
    layer6_outputs(733) <= not(layer5_outputs(200));
    layer6_outputs(734) <= (layer5_outputs(1877)) and not (layer5_outputs(1704));
    layer6_outputs(735) <= not(layer5_outputs(2547)) or (layer5_outputs(2067));
    layer6_outputs(736) <= layer5_outputs(310);
    layer6_outputs(737) <= '1';
    layer6_outputs(738) <= (layer5_outputs(67)) or (layer5_outputs(149));
    layer6_outputs(739) <= not(layer5_outputs(2534)) or (layer5_outputs(318));
    layer6_outputs(740) <= (layer5_outputs(2550)) xor (layer5_outputs(1980));
    layer6_outputs(741) <= not(layer5_outputs(1374));
    layer6_outputs(742) <= (layer5_outputs(2300)) or (layer5_outputs(2500));
    layer6_outputs(743) <= not((layer5_outputs(552)) xor (layer5_outputs(630)));
    layer6_outputs(744) <= layer5_outputs(2099);
    layer6_outputs(745) <= layer5_outputs(565);
    layer6_outputs(746) <= not((layer5_outputs(1275)) xor (layer5_outputs(789)));
    layer6_outputs(747) <= layer5_outputs(1217);
    layer6_outputs(748) <= layer5_outputs(2221);
    layer6_outputs(749) <= layer5_outputs(60);
    layer6_outputs(750) <= not(layer5_outputs(2066));
    layer6_outputs(751) <= not(layer5_outputs(1770));
    layer6_outputs(752) <= (layer5_outputs(1356)) and not (layer5_outputs(1218));
    layer6_outputs(753) <= not(layer5_outputs(2178));
    layer6_outputs(754) <= layer5_outputs(684);
    layer6_outputs(755) <= not(layer5_outputs(2149));
    layer6_outputs(756) <= not(layer5_outputs(1192));
    layer6_outputs(757) <= (layer5_outputs(1062)) and not (layer5_outputs(759));
    layer6_outputs(758) <= not((layer5_outputs(291)) or (layer5_outputs(225)));
    layer6_outputs(759) <= layer5_outputs(794);
    layer6_outputs(760) <= not(layer5_outputs(1407));
    layer6_outputs(761) <= (layer5_outputs(1941)) xor (layer5_outputs(1833));
    layer6_outputs(762) <= not(layer5_outputs(1820));
    layer6_outputs(763) <= (layer5_outputs(1528)) and not (layer5_outputs(2020));
    layer6_outputs(764) <= not(layer5_outputs(1928));
    layer6_outputs(765) <= (layer5_outputs(340)) or (layer5_outputs(2133));
    layer6_outputs(766) <= layer5_outputs(609);
    layer6_outputs(767) <= not(layer5_outputs(1801)) or (layer5_outputs(1164));
    layer6_outputs(768) <= not((layer5_outputs(453)) xor (layer5_outputs(2236)));
    layer6_outputs(769) <= layer5_outputs(641);
    layer6_outputs(770) <= layer5_outputs(1959);
    layer6_outputs(771) <= (layer5_outputs(358)) and not (layer5_outputs(2462));
    layer6_outputs(772) <= layer5_outputs(332);
    layer6_outputs(773) <= layer5_outputs(127);
    layer6_outputs(774) <= not((layer5_outputs(2311)) or (layer5_outputs(1346)));
    layer6_outputs(775) <= not(layer5_outputs(2040)) or (layer5_outputs(1504));
    layer6_outputs(776) <= not(layer5_outputs(2039));
    layer6_outputs(777) <= not((layer5_outputs(1399)) or (layer5_outputs(1146)));
    layer6_outputs(778) <= not(layer5_outputs(924));
    layer6_outputs(779) <= layer5_outputs(107);
    layer6_outputs(780) <= layer5_outputs(569);
    layer6_outputs(781) <= layer5_outputs(1602);
    layer6_outputs(782) <= (layer5_outputs(620)) and not (layer5_outputs(1158));
    layer6_outputs(783) <= not(layer5_outputs(483));
    layer6_outputs(784) <= layer5_outputs(1984);
    layer6_outputs(785) <= layer5_outputs(2008);
    layer6_outputs(786) <= layer5_outputs(899);
    layer6_outputs(787) <= not(layer5_outputs(37));
    layer6_outputs(788) <= not(layer5_outputs(135));
    layer6_outputs(789) <= layer5_outputs(2398);
    layer6_outputs(790) <= not(layer5_outputs(489));
    layer6_outputs(791) <= layer5_outputs(1561);
    layer6_outputs(792) <= not(layer5_outputs(1144)) or (layer5_outputs(2437));
    layer6_outputs(793) <= not(layer5_outputs(2203));
    layer6_outputs(794) <= not(layer5_outputs(1551));
    layer6_outputs(795) <= '1';
    layer6_outputs(796) <= not((layer5_outputs(1934)) and (layer5_outputs(167)));
    layer6_outputs(797) <= not(layer5_outputs(2175));
    layer6_outputs(798) <= not(layer5_outputs(801));
    layer6_outputs(799) <= layer5_outputs(1418);
    layer6_outputs(800) <= not(layer5_outputs(836));
    layer6_outputs(801) <= layer5_outputs(2108);
    layer6_outputs(802) <= not(layer5_outputs(2329));
    layer6_outputs(803) <= not(layer5_outputs(1289));
    layer6_outputs(804) <= layer5_outputs(2475);
    layer6_outputs(805) <= layer5_outputs(1676);
    layer6_outputs(806) <= layer5_outputs(2337);
    layer6_outputs(807) <= not((layer5_outputs(1458)) xor (layer5_outputs(684)));
    layer6_outputs(808) <= (layer5_outputs(1320)) and (layer5_outputs(1888));
    layer6_outputs(809) <= layer5_outputs(1812);
    layer6_outputs(810) <= layer5_outputs(1569);
    layer6_outputs(811) <= layer5_outputs(530);
    layer6_outputs(812) <= not((layer5_outputs(319)) and (layer5_outputs(1644)));
    layer6_outputs(813) <= (layer5_outputs(1524)) or (layer5_outputs(322));
    layer6_outputs(814) <= layer5_outputs(435);
    layer6_outputs(815) <= not(layer5_outputs(2458));
    layer6_outputs(816) <= '0';
    layer6_outputs(817) <= not((layer5_outputs(223)) and (layer5_outputs(1565)));
    layer6_outputs(818) <= not(layer5_outputs(1563));
    layer6_outputs(819) <= layer5_outputs(441);
    layer6_outputs(820) <= not(layer5_outputs(2275));
    layer6_outputs(821) <= (layer5_outputs(1680)) and not (layer5_outputs(1052));
    layer6_outputs(822) <= not(layer5_outputs(1527)) or (layer5_outputs(760));
    layer6_outputs(823) <= not(layer5_outputs(1199)) or (layer5_outputs(1748));
    layer6_outputs(824) <= (layer5_outputs(1966)) or (layer5_outputs(2240));
    layer6_outputs(825) <= not(layer5_outputs(1084));
    layer6_outputs(826) <= not(layer5_outputs(756));
    layer6_outputs(827) <= layer5_outputs(2078);
    layer6_outputs(828) <= not((layer5_outputs(1642)) or (layer5_outputs(834)));
    layer6_outputs(829) <= layer5_outputs(531);
    layer6_outputs(830) <= not(layer5_outputs(67));
    layer6_outputs(831) <= not(layer5_outputs(886));
    layer6_outputs(832) <= layer5_outputs(626);
    layer6_outputs(833) <= '1';
    layer6_outputs(834) <= (layer5_outputs(1924)) and not (layer5_outputs(740));
    layer6_outputs(835) <= not(layer5_outputs(2388));
    layer6_outputs(836) <= not(layer5_outputs(1116));
    layer6_outputs(837) <= layer5_outputs(823);
    layer6_outputs(838) <= not(layer5_outputs(2176));
    layer6_outputs(839) <= (layer5_outputs(636)) or (layer5_outputs(1082));
    layer6_outputs(840) <= not((layer5_outputs(1232)) or (layer5_outputs(1455)));
    layer6_outputs(841) <= layer5_outputs(2013);
    layer6_outputs(842) <= not(layer5_outputs(134)) or (layer5_outputs(778));
    layer6_outputs(843) <= '1';
    layer6_outputs(844) <= not(layer5_outputs(2364)) or (layer5_outputs(2427));
    layer6_outputs(845) <= not(layer5_outputs(244)) or (layer5_outputs(656));
    layer6_outputs(846) <= not(layer5_outputs(1855));
    layer6_outputs(847) <= not((layer5_outputs(1102)) or (layer5_outputs(1709)));
    layer6_outputs(848) <= not(layer5_outputs(1505));
    layer6_outputs(849) <= not(layer5_outputs(1595)) or (layer5_outputs(2123));
    layer6_outputs(850) <= not(layer5_outputs(2040));
    layer6_outputs(851) <= (layer5_outputs(1111)) and not (layer5_outputs(1807));
    layer6_outputs(852) <= not((layer5_outputs(1341)) or (layer5_outputs(675)));
    layer6_outputs(853) <= (layer5_outputs(806)) xor (layer5_outputs(1231));
    layer6_outputs(854) <= not((layer5_outputs(1180)) and (layer5_outputs(2268)));
    layer6_outputs(855) <= not(layer5_outputs(911));
    layer6_outputs(856) <= not((layer5_outputs(730)) xor (layer5_outputs(2274)));
    layer6_outputs(857) <= layer5_outputs(1226);
    layer6_outputs(858) <= layer5_outputs(2371);
    layer6_outputs(859) <= not(layer5_outputs(396));
    layer6_outputs(860) <= not(layer5_outputs(34));
    layer6_outputs(861) <= layer5_outputs(1965);
    layer6_outputs(862) <= not(layer5_outputs(1127));
    layer6_outputs(863) <= (layer5_outputs(2382)) and (layer5_outputs(1207));
    layer6_outputs(864) <= layer5_outputs(970);
    layer6_outputs(865) <= not((layer5_outputs(1475)) and (layer5_outputs(1176)));
    layer6_outputs(866) <= layer5_outputs(1884);
    layer6_outputs(867) <= not(layer5_outputs(2088));
    layer6_outputs(868) <= (layer5_outputs(1015)) and (layer5_outputs(797));
    layer6_outputs(869) <= not(layer5_outputs(2240)) or (layer5_outputs(1006));
    layer6_outputs(870) <= (layer5_outputs(881)) and not (layer5_outputs(2469));
    layer6_outputs(871) <= not((layer5_outputs(165)) and (layer5_outputs(1948)));
    layer6_outputs(872) <= layer5_outputs(1433);
    layer6_outputs(873) <= layer5_outputs(1178);
    layer6_outputs(874) <= layer5_outputs(2460);
    layer6_outputs(875) <= not(layer5_outputs(2090)) or (layer5_outputs(2330));
    layer6_outputs(876) <= (layer5_outputs(720)) and not (layer5_outputs(1359));
    layer6_outputs(877) <= not(layer5_outputs(133));
    layer6_outputs(878) <= not((layer5_outputs(411)) or (layer5_outputs(1897)));
    layer6_outputs(879) <= layer5_outputs(2326);
    layer6_outputs(880) <= not(layer5_outputs(688));
    layer6_outputs(881) <= not(layer5_outputs(2344));
    layer6_outputs(882) <= not(layer5_outputs(473)) or (layer5_outputs(2110));
    layer6_outputs(883) <= layer5_outputs(1707);
    layer6_outputs(884) <= not(layer5_outputs(418));
    layer6_outputs(885) <= layer5_outputs(431);
    layer6_outputs(886) <= not(layer5_outputs(2222));
    layer6_outputs(887) <= layer5_outputs(1771);
    layer6_outputs(888) <= not(layer5_outputs(2443));
    layer6_outputs(889) <= layer5_outputs(2027);
    layer6_outputs(890) <= layer5_outputs(1507);
    layer6_outputs(891) <= not(layer5_outputs(858));
    layer6_outputs(892) <= (layer5_outputs(374)) xor (layer5_outputs(1330));
    layer6_outputs(893) <= not((layer5_outputs(929)) or (layer5_outputs(277)));
    layer6_outputs(894) <= not(layer5_outputs(469));
    layer6_outputs(895) <= not(layer5_outputs(2337));
    layer6_outputs(896) <= layer5_outputs(189);
    layer6_outputs(897) <= not(layer5_outputs(2426));
    layer6_outputs(898) <= not(layer5_outputs(1556));
    layer6_outputs(899) <= layer5_outputs(991);
    layer6_outputs(900) <= not(layer5_outputs(2295)) or (layer5_outputs(586));
    layer6_outputs(901) <= (layer5_outputs(1259)) or (layer5_outputs(1468));
    layer6_outputs(902) <= not((layer5_outputs(239)) or (layer5_outputs(2109)));
    layer6_outputs(903) <= layer5_outputs(833);
    layer6_outputs(904) <= layer5_outputs(1574);
    layer6_outputs(905) <= (layer5_outputs(1274)) xor (layer5_outputs(396));
    layer6_outputs(906) <= not((layer5_outputs(1867)) or (layer5_outputs(2361)));
    layer6_outputs(907) <= layer5_outputs(488);
    layer6_outputs(908) <= (layer5_outputs(2426)) xor (layer5_outputs(1398));
    layer6_outputs(909) <= (layer5_outputs(1549)) xor (layer5_outputs(397));
    layer6_outputs(910) <= (layer5_outputs(1837)) and (layer5_outputs(1918));
    layer6_outputs(911) <= not(layer5_outputs(1301));
    layer6_outputs(912) <= not((layer5_outputs(2128)) xor (layer5_outputs(1719)));
    layer6_outputs(913) <= layer5_outputs(1161);
    layer6_outputs(914) <= (layer5_outputs(512)) xor (layer5_outputs(2315));
    layer6_outputs(915) <= not((layer5_outputs(256)) xor (layer5_outputs(1036)));
    layer6_outputs(916) <= not(layer5_outputs(1660));
    layer6_outputs(917) <= layer5_outputs(1236);
    layer6_outputs(918) <= not(layer5_outputs(2135));
    layer6_outputs(919) <= (layer5_outputs(1743)) and not (layer5_outputs(1397));
    layer6_outputs(920) <= not((layer5_outputs(1267)) or (layer5_outputs(2304)));
    layer6_outputs(921) <= not(layer5_outputs(1130)) or (layer5_outputs(1915));
    layer6_outputs(922) <= not(layer5_outputs(603)) or (layer5_outputs(347));
    layer6_outputs(923) <= not(layer5_outputs(2419));
    layer6_outputs(924) <= not(layer5_outputs(1272)) or (layer5_outputs(2233));
    layer6_outputs(925) <= not((layer5_outputs(54)) and (layer5_outputs(1879)));
    layer6_outputs(926) <= (layer5_outputs(1116)) or (layer5_outputs(1198));
    layer6_outputs(927) <= (layer5_outputs(463)) xor (layer5_outputs(1388));
    layer6_outputs(928) <= not((layer5_outputs(1454)) xor (layer5_outputs(866)));
    layer6_outputs(929) <= (layer5_outputs(673)) or (layer5_outputs(1538));
    layer6_outputs(930) <= not(layer5_outputs(2263));
    layer6_outputs(931) <= not(layer5_outputs(1904)) or (layer5_outputs(1583));
    layer6_outputs(932) <= layer5_outputs(404);
    layer6_outputs(933) <= layer5_outputs(2248);
    layer6_outputs(934) <= not(layer5_outputs(2220)) or (layer5_outputs(2164));
    layer6_outputs(935) <= not(layer5_outputs(850));
    layer6_outputs(936) <= not((layer5_outputs(1353)) and (layer5_outputs(2168)));
    layer6_outputs(937) <= (layer5_outputs(1463)) or (layer5_outputs(2029));
    layer6_outputs(938) <= not(layer5_outputs(2074));
    layer6_outputs(939) <= (layer5_outputs(2230)) and not (layer5_outputs(779));
    layer6_outputs(940) <= not(layer5_outputs(1981));
    layer6_outputs(941) <= not((layer5_outputs(1122)) or (layer5_outputs(858)));
    layer6_outputs(942) <= not(layer5_outputs(708));
    layer6_outputs(943) <= not((layer5_outputs(997)) xor (layer5_outputs(1331)));
    layer6_outputs(944) <= not((layer5_outputs(902)) and (layer5_outputs(1672)));
    layer6_outputs(945) <= (layer5_outputs(2095)) xor (layer5_outputs(59));
    layer6_outputs(946) <= not(layer5_outputs(1366));
    layer6_outputs(947) <= layer5_outputs(993);
    layer6_outputs(948) <= layer5_outputs(2317);
    layer6_outputs(949) <= (layer5_outputs(1787)) xor (layer5_outputs(352));
    layer6_outputs(950) <= (layer5_outputs(1367)) xor (layer5_outputs(1478));
    layer6_outputs(951) <= not(layer5_outputs(1753));
    layer6_outputs(952) <= layer5_outputs(337);
    layer6_outputs(953) <= not(layer5_outputs(697));
    layer6_outputs(954) <= (layer5_outputs(1356)) and (layer5_outputs(389));
    layer6_outputs(955) <= layer5_outputs(1014);
    layer6_outputs(956) <= not(layer5_outputs(1371));
    layer6_outputs(957) <= layer5_outputs(350);
    layer6_outputs(958) <= not(layer5_outputs(2428));
    layer6_outputs(959) <= layer5_outputs(2021);
    layer6_outputs(960) <= '0';
    layer6_outputs(961) <= not((layer5_outputs(2215)) or (layer5_outputs(1186)));
    layer6_outputs(962) <= not(layer5_outputs(2474));
    layer6_outputs(963) <= (layer5_outputs(650)) and (layer5_outputs(1234));
    layer6_outputs(964) <= not((layer5_outputs(1372)) xor (layer5_outputs(1814)));
    layer6_outputs(965) <= not((layer5_outputs(1521)) and (layer5_outputs(994)));
    layer6_outputs(966) <= not(layer5_outputs(1069));
    layer6_outputs(967) <= '0';
    layer6_outputs(968) <= (layer5_outputs(2271)) and not (layer5_outputs(128));
    layer6_outputs(969) <= layer5_outputs(1304);
    layer6_outputs(970) <= not(layer5_outputs(1552));
    layer6_outputs(971) <= (layer5_outputs(1844)) and not (layer5_outputs(1882));
    layer6_outputs(972) <= layer5_outputs(216);
    layer6_outputs(973) <= layer5_outputs(2531);
    layer6_outputs(974) <= layer5_outputs(2456);
    layer6_outputs(975) <= not(layer5_outputs(213));
    layer6_outputs(976) <= (layer5_outputs(1295)) xor (layer5_outputs(2278));
    layer6_outputs(977) <= layer5_outputs(301);
    layer6_outputs(978) <= (layer5_outputs(855)) and not (layer5_outputs(879));
    layer6_outputs(979) <= layer5_outputs(624);
    layer6_outputs(980) <= (layer5_outputs(1285)) or (layer5_outputs(1389));
    layer6_outputs(981) <= layer5_outputs(190);
    layer6_outputs(982) <= not(layer5_outputs(787));
    layer6_outputs(983) <= layer5_outputs(1492);
    layer6_outputs(984) <= not((layer5_outputs(703)) xor (layer5_outputs(171)));
    layer6_outputs(985) <= (layer5_outputs(246)) xor (layer5_outputs(1035));
    layer6_outputs(986) <= not(layer5_outputs(1695));
    layer6_outputs(987) <= (layer5_outputs(1420)) and not (layer5_outputs(2288));
    layer6_outputs(988) <= layer5_outputs(1392);
    layer6_outputs(989) <= not(layer5_outputs(2524));
    layer6_outputs(990) <= layer5_outputs(533);
    layer6_outputs(991) <= layer5_outputs(639);
    layer6_outputs(992) <= not(layer5_outputs(1570));
    layer6_outputs(993) <= (layer5_outputs(1895)) and not (layer5_outputs(1655));
    layer6_outputs(994) <= not(layer5_outputs(1519));
    layer6_outputs(995) <= not((layer5_outputs(1055)) xor (layer5_outputs(1390)));
    layer6_outputs(996) <= not((layer5_outputs(1597)) and (layer5_outputs(2143)));
    layer6_outputs(997) <= not((layer5_outputs(2392)) or (layer5_outputs(23)));
    layer6_outputs(998) <= not(layer5_outputs(1153));
    layer6_outputs(999) <= layer5_outputs(640);
    layer6_outputs(1000) <= layer5_outputs(1422);
    layer6_outputs(1001) <= not(layer5_outputs(989)) or (layer5_outputs(758));
    layer6_outputs(1002) <= not(layer5_outputs(723));
    layer6_outputs(1003) <= not(layer5_outputs(1328));
    layer6_outputs(1004) <= (layer5_outputs(2122)) xor (layer5_outputs(903));
    layer6_outputs(1005) <= not((layer5_outputs(1680)) and (layer5_outputs(1462)));
    layer6_outputs(1006) <= not((layer5_outputs(787)) and (layer5_outputs(662)));
    layer6_outputs(1007) <= not(layer5_outputs(1949));
    layer6_outputs(1008) <= not(layer5_outputs(1922));
    layer6_outputs(1009) <= not((layer5_outputs(963)) xor (layer5_outputs(361)));
    layer6_outputs(1010) <= (layer5_outputs(2002)) xor (layer5_outputs(245));
    layer6_outputs(1011) <= (layer5_outputs(898)) and not (layer5_outputs(208));
    layer6_outputs(1012) <= not(layer5_outputs(613));
    layer6_outputs(1013) <= layer5_outputs(1430);
    layer6_outputs(1014) <= not(layer5_outputs(700)) or (layer5_outputs(1651));
    layer6_outputs(1015) <= (layer5_outputs(2036)) xor (layer5_outputs(1373));
    layer6_outputs(1016) <= layer5_outputs(1911);
    layer6_outputs(1017) <= (layer5_outputs(173)) and (layer5_outputs(1305));
    layer6_outputs(1018) <= not((layer5_outputs(1590)) or (layer5_outputs(416)));
    layer6_outputs(1019) <= layer5_outputs(551);
    layer6_outputs(1020) <= not((layer5_outputs(520)) and (layer5_outputs(801)));
    layer6_outputs(1021) <= not((layer5_outputs(1541)) or (layer5_outputs(1688)));
    layer6_outputs(1022) <= layer5_outputs(2408);
    layer6_outputs(1023) <= (layer5_outputs(1532)) or (layer5_outputs(1943));
    layer6_outputs(1024) <= not(layer5_outputs(1191));
    layer6_outputs(1025) <= layer5_outputs(303);
    layer6_outputs(1026) <= (layer5_outputs(1079)) xor (layer5_outputs(2383));
    layer6_outputs(1027) <= not(layer5_outputs(849));
    layer6_outputs(1028) <= layer5_outputs(1571);
    layer6_outputs(1029) <= layer5_outputs(1862);
    layer6_outputs(1030) <= layer5_outputs(21);
    layer6_outputs(1031) <= (layer5_outputs(2512)) xor (layer5_outputs(907));
    layer6_outputs(1032) <= not(layer5_outputs(1097));
    layer6_outputs(1033) <= layer5_outputs(1507);
    layer6_outputs(1034) <= layer5_outputs(757);
    layer6_outputs(1035) <= '0';
    layer6_outputs(1036) <= layer5_outputs(2221);
    layer6_outputs(1037) <= (layer5_outputs(350)) xor (layer5_outputs(1160));
    layer6_outputs(1038) <= layer5_outputs(132);
    layer6_outputs(1039) <= layer5_outputs(2220);
    layer6_outputs(1040) <= (layer5_outputs(2494)) and not (layer5_outputs(286));
    layer6_outputs(1041) <= not((layer5_outputs(1224)) xor (layer5_outputs(1802)));
    layer6_outputs(1042) <= not(layer5_outputs(502));
    layer6_outputs(1043) <= not(layer5_outputs(1047));
    layer6_outputs(1044) <= layer5_outputs(1132);
    layer6_outputs(1045) <= layer5_outputs(2187);
    layer6_outputs(1046) <= layer5_outputs(1639);
    layer6_outputs(1047) <= not(layer5_outputs(1951));
    layer6_outputs(1048) <= layer5_outputs(2105);
    layer6_outputs(1049) <= not((layer5_outputs(2080)) xor (layer5_outputs(1999)));
    layer6_outputs(1050) <= not(layer5_outputs(269));
    layer6_outputs(1051) <= not(layer5_outputs(1355));
    layer6_outputs(1052) <= not(layer5_outputs(1976));
    layer6_outputs(1053) <= layer5_outputs(2411);
    layer6_outputs(1054) <= layer5_outputs(1405);
    layer6_outputs(1055) <= not((layer5_outputs(414)) xor (layer5_outputs(1893)));
    layer6_outputs(1056) <= (layer5_outputs(66)) and (layer5_outputs(1457));
    layer6_outputs(1057) <= layer5_outputs(843);
    layer6_outputs(1058) <= layer5_outputs(1675);
    layer6_outputs(1059) <= not(layer5_outputs(1498));
    layer6_outputs(1060) <= layer5_outputs(562);
    layer6_outputs(1061) <= layer5_outputs(1572);
    layer6_outputs(1062) <= not(layer5_outputs(1346));
    layer6_outputs(1063) <= not(layer5_outputs(1549));
    layer6_outputs(1064) <= not((layer5_outputs(1224)) and (layer5_outputs(121)));
    layer6_outputs(1065) <= layer5_outputs(247);
    layer6_outputs(1066) <= layer5_outputs(62);
    layer6_outputs(1067) <= not(layer5_outputs(1157)) or (layer5_outputs(2124));
    layer6_outputs(1068) <= layer5_outputs(1734);
    layer6_outputs(1069) <= (layer5_outputs(2300)) and not (layer5_outputs(1409));
    layer6_outputs(1070) <= layer5_outputs(160);
    layer6_outputs(1071) <= not((layer5_outputs(1367)) xor (layer5_outputs(2341)));
    layer6_outputs(1072) <= layer5_outputs(2390);
    layer6_outputs(1073) <= not(layer5_outputs(153)) or (layer5_outputs(1910));
    layer6_outputs(1074) <= not(layer5_outputs(1860));
    layer6_outputs(1075) <= (layer5_outputs(1039)) or (layer5_outputs(1814));
    layer6_outputs(1076) <= layer5_outputs(122);
    layer6_outputs(1077) <= not(layer5_outputs(1143));
    layer6_outputs(1078) <= layer5_outputs(647);
    layer6_outputs(1079) <= (layer5_outputs(598)) or (layer5_outputs(970));
    layer6_outputs(1080) <= (layer5_outputs(224)) or (layer5_outputs(237));
    layer6_outputs(1081) <= layer5_outputs(1738);
    layer6_outputs(1082) <= layer5_outputs(1991);
    layer6_outputs(1083) <= (layer5_outputs(2077)) and not (layer5_outputs(1727));
    layer6_outputs(1084) <= (layer5_outputs(441)) and (layer5_outputs(2501));
    layer6_outputs(1085) <= not(layer5_outputs(515));
    layer6_outputs(1086) <= layer5_outputs(498);
    layer6_outputs(1087) <= layer5_outputs(2218);
    layer6_outputs(1088) <= not(layer5_outputs(1205));
    layer6_outputs(1089) <= not(layer5_outputs(1253)) or (layer5_outputs(1096));
    layer6_outputs(1090) <= layer5_outputs(2441);
    layer6_outputs(1091) <= not(layer5_outputs(889)) or (layer5_outputs(2350));
    layer6_outputs(1092) <= (layer5_outputs(6)) and not (layer5_outputs(1548));
    layer6_outputs(1093) <= not(layer5_outputs(1241));
    layer6_outputs(1094) <= layer5_outputs(1459);
    layer6_outputs(1095) <= (layer5_outputs(573)) xor (layer5_outputs(306));
    layer6_outputs(1096) <= layer5_outputs(548);
    layer6_outputs(1097) <= not(layer5_outputs(109));
    layer6_outputs(1098) <= (layer5_outputs(661)) xor (layer5_outputs(826));
    layer6_outputs(1099) <= (layer5_outputs(2394)) and not (layer5_outputs(2205));
    layer6_outputs(1100) <= layer5_outputs(2031);
    layer6_outputs(1101) <= not(layer5_outputs(741));
    layer6_outputs(1102) <= not((layer5_outputs(2552)) or (layer5_outputs(335)));
    layer6_outputs(1103) <= not(layer5_outputs(2525));
    layer6_outputs(1104) <= not(layer5_outputs(2338));
    layer6_outputs(1105) <= (layer5_outputs(1605)) or (layer5_outputs(1396));
    layer6_outputs(1106) <= not(layer5_outputs(1480));
    layer6_outputs(1107) <= (layer5_outputs(1416)) and not (layer5_outputs(1371));
    layer6_outputs(1108) <= layer5_outputs(1300);
    layer6_outputs(1109) <= layer5_outputs(84);
    layer6_outputs(1110) <= not(layer5_outputs(971));
    layer6_outputs(1111) <= not(layer5_outputs(823));
    layer6_outputs(1112) <= layer5_outputs(1895);
    layer6_outputs(1113) <= (layer5_outputs(698)) and not (layer5_outputs(1034));
    layer6_outputs(1114) <= not(layer5_outputs(734));
    layer6_outputs(1115) <= layer5_outputs(1516);
    layer6_outputs(1116) <= layer5_outputs(978);
    layer6_outputs(1117) <= not(layer5_outputs(425));
    layer6_outputs(1118) <= layer5_outputs(1818);
    layer6_outputs(1119) <= not(layer5_outputs(2185));
    layer6_outputs(1120) <= not((layer5_outputs(44)) or (layer5_outputs(1942)));
    layer6_outputs(1121) <= (layer5_outputs(884)) and not (layer5_outputs(887));
    layer6_outputs(1122) <= not(layer5_outputs(1638));
    layer6_outputs(1123) <= not(layer5_outputs(1369)) or (layer5_outputs(162));
    layer6_outputs(1124) <= layer5_outputs(1903);
    layer6_outputs(1125) <= (layer5_outputs(2155)) and not (layer5_outputs(1957));
    layer6_outputs(1126) <= (layer5_outputs(2542)) and not (layer5_outputs(1641));
    layer6_outputs(1127) <= not(layer5_outputs(1335)) or (layer5_outputs(1256));
    layer6_outputs(1128) <= layer5_outputs(2184);
    layer6_outputs(1129) <= not(layer5_outputs(941));
    layer6_outputs(1130) <= (layer5_outputs(2449)) or (layer5_outputs(1558));
    layer6_outputs(1131) <= not(layer5_outputs(465));
    layer6_outputs(1132) <= not(layer5_outputs(1388));
    layer6_outputs(1133) <= layer5_outputs(1477);
    layer6_outputs(1134) <= not(layer5_outputs(2106));
    layer6_outputs(1135) <= not(layer5_outputs(854));
    layer6_outputs(1136) <= layer5_outputs(695);
    layer6_outputs(1137) <= not(layer5_outputs(1358));
    layer6_outputs(1138) <= '0';
    layer6_outputs(1139) <= (layer5_outputs(491)) xor (layer5_outputs(2340));
    layer6_outputs(1140) <= not(layer5_outputs(847));
    layer6_outputs(1141) <= not((layer5_outputs(2268)) and (layer5_outputs(919)));
    layer6_outputs(1142) <= not(layer5_outputs(2374));
    layer6_outputs(1143) <= layer5_outputs(1142);
    layer6_outputs(1144) <= layer5_outputs(2404);
    layer6_outputs(1145) <= not((layer5_outputs(1711)) xor (layer5_outputs(779)));
    layer6_outputs(1146) <= '1';
    layer6_outputs(1147) <= layer5_outputs(353);
    layer6_outputs(1148) <= layer5_outputs(2324);
    layer6_outputs(1149) <= (layer5_outputs(1115)) and not (layer5_outputs(1705));
    layer6_outputs(1150) <= not(layer5_outputs(37));
    layer6_outputs(1151) <= layer5_outputs(1351);
    layer6_outputs(1152) <= not(layer5_outputs(120));
    layer6_outputs(1153) <= not(layer5_outputs(1874));
    layer6_outputs(1154) <= not((layer5_outputs(1266)) xor (layer5_outputs(410)));
    layer6_outputs(1155) <= layer5_outputs(2339);
    layer6_outputs(1156) <= layer5_outputs(151);
    layer6_outputs(1157) <= not(layer5_outputs(839));
    layer6_outputs(1158) <= not((layer5_outputs(1244)) or (layer5_outputs(2485)));
    layer6_outputs(1159) <= not(layer5_outputs(2345));
    layer6_outputs(1160) <= layer5_outputs(1989);
    layer6_outputs(1161) <= not(layer5_outputs(1093)) or (layer5_outputs(850));
    layer6_outputs(1162) <= not((layer5_outputs(377)) or (layer5_outputs(2340)));
    layer6_outputs(1163) <= (layer5_outputs(2409)) and (layer5_outputs(1183));
    layer6_outputs(1164) <= not(layer5_outputs(799));
    layer6_outputs(1165) <= not(layer5_outputs(197));
    layer6_outputs(1166) <= not((layer5_outputs(1378)) xor (layer5_outputs(604)));
    layer6_outputs(1167) <= not(layer5_outputs(1668));
    layer6_outputs(1168) <= not(layer5_outputs(452));
    layer6_outputs(1169) <= layer5_outputs(1145);
    layer6_outputs(1170) <= not((layer5_outputs(1534)) and (layer5_outputs(1289)));
    layer6_outputs(1171) <= not((layer5_outputs(1684)) xor (layer5_outputs(1496)));
    layer6_outputs(1172) <= not((layer5_outputs(1070)) or (layer5_outputs(2229)));
    layer6_outputs(1173) <= (layer5_outputs(765)) or (layer5_outputs(137));
    layer6_outputs(1174) <= layer5_outputs(2358);
    layer6_outputs(1175) <= (layer5_outputs(214)) xor (layer5_outputs(1746));
    layer6_outputs(1176) <= not(layer5_outputs(2188));
    layer6_outputs(1177) <= (layer5_outputs(1789)) and (layer5_outputs(1363));
    layer6_outputs(1178) <= not(layer5_outputs(1424)) or (layer5_outputs(1620));
    layer6_outputs(1179) <= not(layer5_outputs(1762)) or (layer5_outputs(170));
    layer6_outputs(1180) <= layer5_outputs(2418);
    layer6_outputs(1181) <= (layer5_outputs(1989)) xor (layer5_outputs(2002));
    layer6_outputs(1182) <= not(layer5_outputs(747));
    layer6_outputs(1183) <= layer5_outputs(2367);
    layer6_outputs(1184) <= not((layer5_outputs(2137)) xor (layer5_outputs(2545)));
    layer6_outputs(1185) <= (layer5_outputs(1571)) xor (layer5_outputs(186));
    layer6_outputs(1186) <= not(layer5_outputs(1082)) or (layer5_outputs(1391));
    layer6_outputs(1187) <= (layer5_outputs(697)) and not (layer5_outputs(2362));
    layer6_outputs(1188) <= not(layer5_outputs(2502));
    layer6_outputs(1189) <= '1';
    layer6_outputs(1190) <= not(layer5_outputs(2527)) or (layer5_outputs(2278));
    layer6_outputs(1191) <= not((layer5_outputs(2504)) or (layer5_outputs(1385)));
    layer6_outputs(1192) <= not(layer5_outputs(754)) or (layer5_outputs(60));
    layer6_outputs(1193) <= not(layer5_outputs(1631));
    layer6_outputs(1194) <= layer5_outputs(702);
    layer6_outputs(1195) <= layer5_outputs(1272);
    layer6_outputs(1196) <= (layer5_outputs(2507)) or (layer5_outputs(1631));
    layer6_outputs(1197) <= layer5_outputs(2323);
    layer6_outputs(1198) <= layer5_outputs(1712);
    layer6_outputs(1199) <= not(layer5_outputs(2208));
    layer6_outputs(1200) <= not(layer5_outputs(530));
    layer6_outputs(1201) <= '0';
    layer6_outputs(1202) <= not(layer5_outputs(56));
    layer6_outputs(1203) <= layer5_outputs(531);
    layer6_outputs(1204) <= (layer5_outputs(1476)) or (layer5_outputs(2113));
    layer6_outputs(1205) <= not(layer5_outputs(16)) or (layer5_outputs(1718));
    layer6_outputs(1206) <= (layer5_outputs(2547)) xor (layer5_outputs(579));
    layer6_outputs(1207) <= (layer5_outputs(2380)) and (layer5_outputs(116));
    layer6_outputs(1208) <= not(layer5_outputs(69)) or (layer5_outputs(2144));
    layer6_outputs(1209) <= not((layer5_outputs(830)) xor (layer5_outputs(771)));
    layer6_outputs(1210) <= not((layer5_outputs(126)) or (layer5_outputs(2267)));
    layer6_outputs(1211) <= layer5_outputs(3);
    layer6_outputs(1212) <= layer5_outputs(2250);
    layer6_outputs(1213) <= layer5_outputs(2037);
    layer6_outputs(1214) <= (layer5_outputs(2374)) and not (layer5_outputs(1045));
    layer6_outputs(1215) <= not(layer5_outputs(1685));
    layer6_outputs(1216) <= (layer5_outputs(124)) and not (layer5_outputs(534));
    layer6_outputs(1217) <= not(layer5_outputs(1998)) or (layer5_outputs(851));
    layer6_outputs(1218) <= not(layer5_outputs(1027));
    layer6_outputs(1219) <= layer5_outputs(1460);
    layer6_outputs(1220) <= not(layer5_outputs(506));
    layer6_outputs(1221) <= '1';
    layer6_outputs(1222) <= not(layer5_outputs(250));
    layer6_outputs(1223) <= (layer5_outputs(1774)) and (layer5_outputs(1913));
    layer6_outputs(1224) <= not((layer5_outputs(1044)) and (layer5_outputs(63)));
    layer6_outputs(1225) <= layer5_outputs(774);
    layer6_outputs(1226) <= layer5_outputs(2375);
    layer6_outputs(1227) <= (layer5_outputs(2207)) xor (layer5_outputs(137));
    layer6_outputs(1228) <= (layer5_outputs(2420)) and not (layer5_outputs(812));
    layer6_outputs(1229) <= not((layer5_outputs(2470)) xor (layer5_outputs(2051)));
    layer6_outputs(1230) <= not(layer5_outputs(725)) or (layer5_outputs(1596));
    layer6_outputs(1231) <= layer5_outputs(2094);
    layer6_outputs(1232) <= layer5_outputs(53);
    layer6_outputs(1233) <= not((layer5_outputs(706)) or (layer5_outputs(749)));
    layer6_outputs(1234) <= layer5_outputs(2271);
    layer6_outputs(1235) <= not(layer5_outputs(383));
    layer6_outputs(1236) <= not(layer5_outputs(2124));
    layer6_outputs(1237) <= layer5_outputs(593);
    layer6_outputs(1238) <= layer5_outputs(563);
    layer6_outputs(1239) <= not(layer5_outputs(1671));
    layer6_outputs(1240) <= not((layer5_outputs(1384)) and (layer5_outputs(1956)));
    layer6_outputs(1241) <= not((layer5_outputs(2446)) xor (layer5_outputs(187)));
    layer6_outputs(1242) <= not(layer5_outputs(93));
    layer6_outputs(1243) <= not(layer5_outputs(1713));
    layer6_outputs(1244) <= layer5_outputs(1858);
    layer6_outputs(1245) <= (layer5_outputs(1001)) and not (layer5_outputs(430));
    layer6_outputs(1246) <= layer5_outputs(1992);
    layer6_outputs(1247) <= (layer5_outputs(2042)) xor (layer5_outputs(2264));
    layer6_outputs(1248) <= (layer5_outputs(2082)) xor (layer5_outputs(472));
    layer6_outputs(1249) <= not(layer5_outputs(2090));
    layer6_outputs(1250) <= layer5_outputs(1311);
    layer6_outputs(1251) <= not(layer5_outputs(109));
    layer6_outputs(1252) <= (layer5_outputs(1625)) xor (layer5_outputs(1532));
    layer6_outputs(1253) <= layer5_outputs(1038);
    layer6_outputs(1254) <= (layer5_outputs(331)) and (layer5_outputs(161));
    layer6_outputs(1255) <= not(layer5_outputs(1430));
    layer6_outputs(1256) <= not(layer5_outputs(2279)) or (layer5_outputs(1885));
    layer6_outputs(1257) <= (layer5_outputs(391)) or (layer5_outputs(1131));
    layer6_outputs(1258) <= not((layer5_outputs(278)) or (layer5_outputs(124)));
    layer6_outputs(1259) <= not(layer5_outputs(711));
    layer6_outputs(1260) <= not((layer5_outputs(866)) xor (layer5_outputs(2020)));
    layer6_outputs(1261) <= (layer5_outputs(2056)) and not (layer5_outputs(844));
    layer6_outputs(1262) <= not((layer5_outputs(1326)) and (layer5_outputs(694)));
    layer6_outputs(1263) <= layer5_outputs(2098);
    layer6_outputs(1264) <= (layer5_outputs(319)) xor (layer5_outputs(1524));
    layer6_outputs(1265) <= not(layer5_outputs(696)) or (layer5_outputs(2515));
    layer6_outputs(1266) <= not(layer5_outputs(2174));
    layer6_outputs(1267) <= (layer5_outputs(678)) and not (layer5_outputs(1513));
    layer6_outputs(1268) <= not(layer5_outputs(1458)) or (layer5_outputs(1545));
    layer6_outputs(1269) <= layer5_outputs(669);
    layer6_outputs(1270) <= layer5_outputs(1004);
    layer6_outputs(1271) <= not((layer5_outputs(1550)) or (layer5_outputs(725)));
    layer6_outputs(1272) <= (layer5_outputs(2201)) and not (layer5_outputs(529));
    layer6_outputs(1273) <= not((layer5_outputs(2364)) and (layer5_outputs(74)));
    layer6_outputs(1274) <= not(layer5_outputs(871));
    layer6_outputs(1275) <= (layer5_outputs(1170)) and (layer5_outputs(2543));
    layer6_outputs(1276) <= not(layer5_outputs(1169));
    layer6_outputs(1277) <= layer5_outputs(669);
    layer6_outputs(1278) <= not(layer5_outputs(475));
    layer6_outputs(1279) <= not((layer5_outputs(1100)) xor (layer5_outputs(262)));
    layer6_outputs(1280) <= not(layer5_outputs(1083));
    layer6_outputs(1281) <= (layer5_outputs(2214)) and (layer5_outputs(1316));
    layer6_outputs(1282) <= not(layer5_outputs(475));
    layer6_outputs(1283) <= layer5_outputs(2156);
    layer6_outputs(1284) <= layer5_outputs(1453);
    layer6_outputs(1285) <= layer5_outputs(1118);
    layer6_outputs(1286) <= not((layer5_outputs(2299)) and (layer5_outputs(1445)));
    layer6_outputs(1287) <= (layer5_outputs(2272)) and not (layer5_outputs(931));
    layer6_outputs(1288) <= layer5_outputs(558);
    layer6_outputs(1289) <= not(layer5_outputs(2047));
    layer6_outputs(1290) <= (layer5_outputs(294)) xor (layer5_outputs(1512));
    layer6_outputs(1291) <= layer5_outputs(878);
    layer6_outputs(1292) <= layer5_outputs(596);
    layer6_outputs(1293) <= not(layer5_outputs(72));
    layer6_outputs(1294) <= not((layer5_outputs(2403)) xor (layer5_outputs(983)));
    layer6_outputs(1295) <= not((layer5_outputs(1767)) and (layer5_outputs(1842)));
    layer6_outputs(1296) <= layer5_outputs(662);
    layer6_outputs(1297) <= (layer5_outputs(428)) xor (layer5_outputs(1818));
    layer6_outputs(1298) <= layer5_outputs(1575);
    layer6_outputs(1299) <= not(layer5_outputs(380));
    layer6_outputs(1300) <= not(layer5_outputs(603));
    layer6_outputs(1301) <= not(layer5_outputs(2246));
    layer6_outputs(1302) <= not(layer5_outputs(1745));
    layer6_outputs(1303) <= (layer5_outputs(1954)) and (layer5_outputs(1148));
    layer6_outputs(1304) <= layer5_outputs(1657);
    layer6_outputs(1305) <= not((layer5_outputs(1581)) or (layer5_outputs(1979)));
    layer6_outputs(1306) <= (layer5_outputs(1997)) xor (layer5_outputs(58));
    layer6_outputs(1307) <= not(layer5_outputs(2445));
    layer6_outputs(1308) <= not(layer5_outputs(1423));
    layer6_outputs(1309) <= (layer5_outputs(17)) xor (layer5_outputs(2363));
    layer6_outputs(1310) <= '1';
    layer6_outputs(1311) <= layer5_outputs(2386);
    layer6_outputs(1312) <= (layer5_outputs(290)) xor (layer5_outputs(973));
    layer6_outputs(1313) <= not(layer5_outputs(1918));
    layer6_outputs(1314) <= layer5_outputs(2266);
    layer6_outputs(1315) <= not((layer5_outputs(2536)) xor (layer5_outputs(467)));
    layer6_outputs(1316) <= (layer5_outputs(1614)) or (layer5_outputs(2163));
    layer6_outputs(1317) <= not(layer5_outputs(1984));
    layer6_outputs(1318) <= (layer5_outputs(1505)) and (layer5_outputs(549));
    layer6_outputs(1319) <= (layer5_outputs(901)) xor (layer5_outputs(1578));
    layer6_outputs(1320) <= (layer5_outputs(764)) and (layer5_outputs(1881));
    layer6_outputs(1321) <= not(layer5_outputs(1295));
    layer6_outputs(1322) <= not(layer5_outputs(1578));
    layer6_outputs(1323) <= not((layer5_outputs(227)) and (layer5_outputs(2481)));
    layer6_outputs(1324) <= not((layer5_outputs(1962)) xor (layer5_outputs(1690)));
    layer6_outputs(1325) <= not(layer5_outputs(1331));
    layer6_outputs(1326) <= layer5_outputs(1011);
    layer6_outputs(1327) <= not(layer5_outputs(436)) or (layer5_outputs(284));
    layer6_outputs(1328) <= layer5_outputs(1283);
    layer6_outputs(1329) <= (layer5_outputs(1794)) and not (layer5_outputs(97));
    layer6_outputs(1330) <= layer5_outputs(1197);
    layer6_outputs(1331) <= layer5_outputs(2369);
    layer6_outputs(1332) <= not(layer5_outputs(398));
    layer6_outputs(1333) <= not(layer5_outputs(2186)) or (layer5_outputs(1406));
    layer6_outputs(1334) <= (layer5_outputs(881)) and not (layer5_outputs(1623));
    layer6_outputs(1335) <= not((layer5_outputs(1240)) xor (layer5_outputs(2325)));
    layer6_outputs(1336) <= not(layer5_outputs(1649)) or (layer5_outputs(1777));
    layer6_outputs(1337) <= not((layer5_outputs(2554)) or (layer5_outputs(103)));
    layer6_outputs(1338) <= (layer5_outputs(2227)) and (layer5_outputs(876));
    layer6_outputs(1339) <= layer5_outputs(411);
    layer6_outputs(1340) <= (layer5_outputs(2366)) and not (layer5_outputs(75));
    layer6_outputs(1341) <= not(layer5_outputs(2476));
    layer6_outputs(1342) <= not(layer5_outputs(915));
    layer6_outputs(1343) <= not((layer5_outputs(1726)) xor (layer5_outputs(1604)));
    layer6_outputs(1344) <= not(layer5_outputs(539));
    layer6_outputs(1345) <= not((layer5_outputs(540)) and (layer5_outputs(559)));
    layer6_outputs(1346) <= not(layer5_outputs(1929)) or (layer5_outputs(2370));
    layer6_outputs(1347) <= layer5_outputs(1821);
    layer6_outputs(1348) <= not(layer5_outputs(447));
    layer6_outputs(1349) <= not(layer5_outputs(1525));
    layer6_outputs(1350) <= not((layer5_outputs(1778)) and (layer5_outputs(1270)));
    layer6_outputs(1351) <= layer5_outputs(385);
    layer6_outputs(1352) <= not(layer5_outputs(2212));
    layer6_outputs(1353) <= not(layer5_outputs(1119));
    layer6_outputs(1354) <= (layer5_outputs(796)) and (layer5_outputs(144));
    layer6_outputs(1355) <= layer5_outputs(2025);
    layer6_outputs(1356) <= not(layer5_outputs(1446));
    layer6_outputs(1357) <= (layer5_outputs(1690)) xor (layer5_outputs(2026));
    layer6_outputs(1358) <= not(layer5_outputs(1514));
    layer6_outputs(1359) <= not((layer5_outputs(1781)) and (layer5_outputs(984)));
    layer6_outputs(1360) <= not(layer5_outputs(456));
    layer6_outputs(1361) <= layer5_outputs(583);
    layer6_outputs(1362) <= not(layer5_outputs(466));
    layer6_outputs(1363) <= not(layer5_outputs(57));
    layer6_outputs(1364) <= layer5_outputs(554);
    layer6_outputs(1365) <= layer5_outputs(2284);
    layer6_outputs(1366) <= not(layer5_outputs(674)) or (layer5_outputs(936));
    layer6_outputs(1367) <= not((layer5_outputs(640)) or (layer5_outputs(1647)));
    layer6_outputs(1368) <= layer5_outputs(38);
    layer6_outputs(1369) <= layer5_outputs(2275);
    layer6_outputs(1370) <= not(layer5_outputs(1947));
    layer6_outputs(1371) <= not((layer5_outputs(2119)) xor (layer5_outputs(1537)));
    layer6_outputs(1372) <= not(layer5_outputs(2342));
    layer6_outputs(1373) <= not(layer5_outputs(2509));
    layer6_outputs(1374) <= not(layer5_outputs(230));
    layer6_outputs(1375) <= layer5_outputs(2159);
    layer6_outputs(1376) <= not(layer5_outputs(1299)) or (layer5_outputs(210));
    layer6_outputs(1377) <= layer5_outputs(1925);
    layer6_outputs(1378) <= layer5_outputs(1826);
    layer6_outputs(1379) <= (layer5_outputs(2523)) and not (layer5_outputs(339));
    layer6_outputs(1380) <= not(layer5_outputs(1287)) or (layer5_outputs(2309));
    layer6_outputs(1381) <= layer5_outputs(150);
    layer6_outputs(1382) <= (layer5_outputs(554)) and (layer5_outputs(1171));
    layer6_outputs(1383) <= (layer5_outputs(2127)) and not (layer5_outputs(1175));
    layer6_outputs(1384) <= (layer5_outputs(89)) xor (layer5_outputs(1113));
    layer6_outputs(1385) <= (layer5_outputs(103)) and not (layer5_outputs(1273));
    layer6_outputs(1386) <= not((layer5_outputs(1296)) or (layer5_outputs(782)));
    layer6_outputs(1387) <= layer5_outputs(1376);
    layer6_outputs(1388) <= not(layer5_outputs(130));
    layer6_outputs(1389) <= layer5_outputs(2004);
    layer6_outputs(1390) <= layer5_outputs(202);
    layer6_outputs(1391) <= not(layer5_outputs(557));
    layer6_outputs(1392) <= layer5_outputs(1308);
    layer6_outputs(1393) <= (layer5_outputs(214)) xor (layer5_outputs(1910));
    layer6_outputs(1394) <= layer5_outputs(941);
    layer6_outputs(1395) <= (layer5_outputs(1273)) and not (layer5_outputs(2248));
    layer6_outputs(1396) <= (layer5_outputs(1692)) xor (layer5_outputs(614));
    layer6_outputs(1397) <= not(layer5_outputs(1506));
    layer6_outputs(1398) <= layer5_outputs(516);
    layer6_outputs(1399) <= '0';
    layer6_outputs(1400) <= layer5_outputs(2262);
    layer6_outputs(1401) <= not(layer5_outputs(1081));
    layer6_outputs(1402) <= (layer5_outputs(2063)) and not (layer5_outputs(2194));
    layer6_outputs(1403) <= layer5_outputs(111);
    layer6_outputs(1404) <= layer5_outputs(1217);
    layer6_outputs(1405) <= not(layer5_outputs(905));
    layer6_outputs(1406) <= not(layer5_outputs(2243)) or (layer5_outputs(71));
    layer6_outputs(1407) <= not(layer5_outputs(373));
    layer6_outputs(1408) <= (layer5_outputs(221)) and not (layer5_outputs(1200));
    layer6_outputs(1409) <= (layer5_outputs(1652)) and (layer5_outputs(327));
    layer6_outputs(1410) <= not((layer5_outputs(1823)) xor (layer5_outputs(1748)));
    layer6_outputs(1411) <= (layer5_outputs(494)) and not (layer5_outputs(1671));
    layer6_outputs(1412) <= not(layer5_outputs(2429));
    layer6_outputs(1413) <= not(layer5_outputs(2225));
    layer6_outputs(1414) <= not(layer5_outputs(2298));
    layer6_outputs(1415) <= not(layer5_outputs(1714));
    layer6_outputs(1416) <= not(layer5_outputs(1835));
    layer6_outputs(1417) <= (layer5_outputs(839)) xor (layer5_outputs(695));
    layer6_outputs(1418) <= layer5_outputs(978);
    layer6_outputs(1419) <= not(layer5_outputs(1709));
    layer6_outputs(1420) <= (layer5_outputs(1550)) or (layer5_outputs(1594));
    layer6_outputs(1421) <= not((layer5_outputs(2075)) xor (layer5_outputs(1493)));
    layer6_outputs(1422) <= layer5_outputs(1728);
    layer6_outputs(1423) <= (layer5_outputs(1607)) xor (layer5_outputs(2400));
    layer6_outputs(1424) <= not((layer5_outputs(969)) xor (layer5_outputs(1969)));
    layer6_outputs(1425) <= (layer5_outputs(2512)) xor (layer5_outputs(1311));
    layer6_outputs(1426) <= (layer5_outputs(2412)) or (layer5_outputs(1886));
    layer6_outputs(1427) <= (layer5_outputs(1848)) xor (layer5_outputs(1130));
    layer6_outputs(1428) <= layer5_outputs(1609);
    layer6_outputs(1429) <= (layer5_outputs(1247)) or (layer5_outputs(2378));
    layer6_outputs(1430) <= layer5_outputs(1187);
    layer6_outputs(1431) <= (layer5_outputs(1904)) and (layer5_outputs(1985));
    layer6_outputs(1432) <= layer5_outputs(1004);
    layer6_outputs(1433) <= layer5_outputs(867);
    layer6_outputs(1434) <= not(layer5_outputs(2499));
    layer6_outputs(1435) <= (layer5_outputs(453)) xor (layer5_outputs(1070));
    layer6_outputs(1436) <= layer5_outputs(2155);
    layer6_outputs(1437) <= layer5_outputs(1390);
    layer6_outputs(1438) <= not((layer5_outputs(21)) or (layer5_outputs(772)));
    layer6_outputs(1439) <= not(layer5_outputs(1194));
    layer6_outputs(1440) <= not(layer5_outputs(1906));
    layer6_outputs(1441) <= '1';
    layer6_outputs(1442) <= not(layer5_outputs(1499)) or (layer5_outputs(171));
    layer6_outputs(1443) <= not(layer5_outputs(300));
    layer6_outputs(1444) <= layer5_outputs(1460);
    layer6_outputs(1445) <= not((layer5_outputs(2462)) and (layer5_outputs(2530)));
    layer6_outputs(1446) <= layer5_outputs(1827);
    layer6_outputs(1447) <= (layer5_outputs(950)) and (layer5_outputs(2451));
    layer6_outputs(1448) <= layer5_outputs(911);
    layer6_outputs(1449) <= (layer5_outputs(1754)) and not (layer5_outputs(1956));
    layer6_outputs(1450) <= not((layer5_outputs(1090)) xor (layer5_outputs(586)));
    layer6_outputs(1451) <= not(layer5_outputs(1091));
    layer6_outputs(1452) <= not(layer5_outputs(924));
    layer6_outputs(1453) <= layer5_outputs(594);
    layer6_outputs(1454) <= not(layer5_outputs(1716));
    layer6_outputs(1455) <= not(layer5_outputs(2224)) or (layer5_outputs(1471));
    layer6_outputs(1456) <= (layer5_outputs(1670)) xor (layer5_outputs(106));
    layer6_outputs(1457) <= not(layer5_outputs(1245));
    layer6_outputs(1458) <= layer5_outputs(2062);
    layer6_outputs(1459) <= not(layer5_outputs(859));
    layer6_outputs(1460) <= layer5_outputs(632);
    layer6_outputs(1461) <= not((layer5_outputs(942)) or (layer5_outputs(792)));
    layer6_outputs(1462) <= not((layer5_outputs(192)) xor (layer5_outputs(141)));
    layer6_outputs(1463) <= not((layer5_outputs(2378)) or (layer5_outputs(1446)));
    layer6_outputs(1464) <= (layer5_outputs(2506)) xor (layer5_outputs(1158));
    layer6_outputs(1465) <= '1';
    layer6_outputs(1466) <= layer5_outputs(251);
    layer6_outputs(1467) <= not((layer5_outputs(1397)) xor (layer5_outputs(1495)));
    layer6_outputs(1468) <= not(layer5_outputs(558));
    layer6_outputs(1469) <= (layer5_outputs(1899)) and (layer5_outputs(2387));
    layer6_outputs(1470) <= (layer5_outputs(1728)) or (layer5_outputs(665));
    layer6_outputs(1471) <= (layer5_outputs(1944)) xor (layer5_outputs(2327));
    layer6_outputs(1472) <= not(layer5_outputs(1885)) or (layer5_outputs(903));
    layer6_outputs(1473) <= (layer5_outputs(36)) and (layer5_outputs(1497));
    layer6_outputs(1474) <= not((layer5_outputs(223)) or (layer5_outputs(369)));
    layer6_outputs(1475) <= not(layer5_outputs(2475)) or (layer5_outputs(673));
    layer6_outputs(1476) <= not(layer5_outputs(606));
    layer6_outputs(1477) <= not((layer5_outputs(670)) or (layer5_outputs(1699)));
    layer6_outputs(1478) <= layer5_outputs(739);
    layer6_outputs(1479) <= not(layer5_outputs(2522));
    layer6_outputs(1480) <= not(layer5_outputs(897));
    layer6_outputs(1481) <= not(layer5_outputs(1519));
    layer6_outputs(1482) <= layer5_outputs(76);
    layer6_outputs(1483) <= layer5_outputs(1452);
    layer6_outputs(1484) <= (layer5_outputs(740)) or (layer5_outputs(2444));
    layer6_outputs(1485) <= not(layer5_outputs(1843));
    layer6_outputs(1486) <= not(layer5_outputs(605)) or (layer5_outputs(718));
    layer6_outputs(1487) <= layer5_outputs(951);
    layer6_outputs(1488) <= not(layer5_outputs(1557));
    layer6_outputs(1489) <= not(layer5_outputs(2382)) or (layer5_outputs(838));
    layer6_outputs(1490) <= (layer5_outputs(1189)) and not (layer5_outputs(909));
    layer6_outputs(1491) <= layer5_outputs(648);
    layer6_outputs(1492) <= layer5_outputs(1737);
    layer6_outputs(1493) <= (layer5_outputs(675)) and not (layer5_outputs(499));
    layer6_outputs(1494) <= layer5_outputs(1679);
    layer6_outputs(1495) <= not(layer5_outputs(77));
    layer6_outputs(1496) <= not((layer5_outputs(2058)) and (layer5_outputs(2259)));
    layer6_outputs(1497) <= not(layer5_outputs(738)) or (layer5_outputs(2285));
    layer6_outputs(1498) <= not(layer5_outputs(1738)) or (layer5_outputs(979));
    layer6_outputs(1499) <= (layer5_outputs(1609)) and (layer5_outputs(2285));
    layer6_outputs(1500) <= (layer5_outputs(998)) and not (layer5_outputs(1221));
    layer6_outputs(1501) <= not(layer5_outputs(1882));
    layer6_outputs(1502) <= not((layer5_outputs(77)) and (layer5_outputs(1930)));
    layer6_outputs(1503) <= not(layer5_outputs(1799));
    layer6_outputs(1504) <= layer5_outputs(242);
    layer6_outputs(1505) <= not(layer5_outputs(776));
    layer6_outputs(1506) <= layer5_outputs(1648);
    layer6_outputs(1507) <= (layer5_outputs(664)) xor (layer5_outputs(696));
    layer6_outputs(1508) <= (layer5_outputs(923)) xor (layer5_outputs(1072));
    layer6_outputs(1509) <= not(layer5_outputs(83)) or (layer5_outputs(1703));
    layer6_outputs(1510) <= not(layer5_outputs(86));
    layer6_outputs(1511) <= not(layer5_outputs(443));
    layer6_outputs(1512) <= not(layer5_outputs(2377)) or (layer5_outputs(580));
    layer6_outputs(1513) <= (layer5_outputs(211)) xor (layer5_outputs(1856));
    layer6_outputs(1514) <= layer5_outputs(1260);
    layer6_outputs(1515) <= layer5_outputs(128);
    layer6_outputs(1516) <= layer5_outputs(1828);
    layer6_outputs(1517) <= not((layer5_outputs(1212)) xor (layer5_outputs(499)));
    layer6_outputs(1518) <= not(layer5_outputs(1795));
    layer6_outputs(1519) <= layer5_outputs(2503);
    layer6_outputs(1520) <= layer5_outputs(1119);
    layer6_outputs(1521) <= layer5_outputs(329);
    layer6_outputs(1522) <= not(layer5_outputs(2442));
    layer6_outputs(1523) <= not(layer5_outputs(355));
    layer6_outputs(1524) <= not(layer5_outputs(1803)) or (layer5_outputs(578));
    layer6_outputs(1525) <= (layer5_outputs(2553)) and not (layer5_outputs(842));
    layer6_outputs(1526) <= '1';
    layer6_outputs(1527) <= not(layer5_outputs(394));
    layer6_outputs(1528) <= layer5_outputs(761);
    layer6_outputs(1529) <= not(layer5_outputs(1473));
    layer6_outputs(1530) <= not(layer5_outputs(2397));
    layer6_outputs(1531) <= (layer5_outputs(2452)) or (layer5_outputs(815));
    layer6_outputs(1532) <= not(layer5_outputs(817));
    layer6_outputs(1533) <= not(layer5_outputs(2069));
    layer6_outputs(1534) <= not((layer5_outputs(1529)) or (layer5_outputs(1908)));
    layer6_outputs(1535) <= (layer5_outputs(1639)) and not (layer5_outputs(996));
    layer6_outputs(1536) <= (layer5_outputs(41)) xor (layer5_outputs(1698));
    layer6_outputs(1537) <= (layer5_outputs(809)) xor (layer5_outputs(2557));
    layer6_outputs(1538) <= layer5_outputs(1711);
    layer6_outputs(1539) <= (layer5_outputs(1568)) xor (layer5_outputs(2081));
    layer6_outputs(1540) <= layer5_outputs(2279);
    layer6_outputs(1541) <= (layer5_outputs(2105)) and (layer5_outputs(271));
    layer6_outputs(1542) <= layer5_outputs(1249);
    layer6_outputs(1543) <= not(layer5_outputs(872));
    layer6_outputs(1544) <= not(layer5_outputs(1172));
    layer6_outputs(1545) <= not(layer5_outputs(819));
    layer6_outputs(1546) <= (layer5_outputs(46)) xor (layer5_outputs(2016));
    layer6_outputs(1547) <= not(layer5_outputs(1287));
    layer6_outputs(1548) <= layer5_outputs(222);
    layer6_outputs(1549) <= '0';
    layer6_outputs(1550) <= not((layer5_outputs(493)) xor (layer5_outputs(1178)));
    layer6_outputs(1551) <= not(layer5_outputs(1767)) or (layer5_outputs(2204));
    layer6_outputs(1552) <= not((layer5_outputs(2064)) and (layer5_outputs(1081)));
    layer6_outputs(1553) <= layer5_outputs(704);
    layer6_outputs(1554) <= layer5_outputs(113);
    layer6_outputs(1555) <= not((layer5_outputs(2463)) xor (layer5_outputs(369)));
    layer6_outputs(1556) <= layer5_outputs(893);
    layer6_outputs(1557) <= layer5_outputs(2030);
    layer6_outputs(1558) <= not(layer5_outputs(2365)) or (layer5_outputs(47));
    layer6_outputs(1559) <= (layer5_outputs(2332)) and (layer5_outputs(1327));
    layer6_outputs(1560) <= (layer5_outputs(1898)) and (layer5_outputs(627));
    layer6_outputs(1561) <= layer5_outputs(687);
    layer6_outputs(1562) <= layer5_outputs(1056);
    layer6_outputs(1563) <= layer5_outputs(1209);
    layer6_outputs(1564) <= (layer5_outputs(473)) xor (layer5_outputs(2517));
    layer6_outputs(1565) <= (layer5_outputs(1734)) and not (layer5_outputs(1188));
    layer6_outputs(1566) <= not(layer5_outputs(2192));
    layer6_outputs(1567) <= (layer5_outputs(857)) xor (layer5_outputs(151));
    layer6_outputs(1568) <= not(layer5_outputs(1355));
    layer6_outputs(1569) <= (layer5_outputs(53)) xor (layer5_outputs(1661));
    layer6_outputs(1570) <= not((layer5_outputs(2200)) xor (layer5_outputs(1613)));
    layer6_outputs(1571) <= (layer5_outputs(94)) xor (layer5_outputs(860));
    layer6_outputs(1572) <= not((layer5_outputs(1863)) and (layer5_outputs(811)));
    layer6_outputs(1573) <= not(layer5_outputs(2187));
    layer6_outputs(1574) <= (layer5_outputs(2508)) and not (layer5_outputs(1724));
    layer6_outputs(1575) <= not((layer5_outputs(1937)) xor (layer5_outputs(2431)));
    layer6_outputs(1576) <= layer5_outputs(1189);
    layer6_outputs(1577) <= (layer5_outputs(368)) xor (layer5_outputs(2044));
    layer6_outputs(1578) <= not(layer5_outputs(3));
    layer6_outputs(1579) <= not(layer5_outputs(1448)) or (layer5_outputs(1401));
    layer6_outputs(1580) <= layer5_outputs(1488);
    layer6_outputs(1581) <= not((layer5_outputs(6)) xor (layer5_outputs(1223)));
    layer6_outputs(1582) <= (layer5_outputs(884)) and (layer5_outputs(2086));
    layer6_outputs(1583) <= (layer5_outputs(1306)) or (layer5_outputs(1491));
    layer6_outputs(1584) <= not(layer5_outputs(1774));
    layer6_outputs(1585) <= layer5_outputs(882);
    layer6_outputs(1586) <= (layer5_outputs(853)) xor (layer5_outputs(1762));
    layer6_outputs(1587) <= (layer5_outputs(479)) and not (layer5_outputs(702));
    layer6_outputs(1588) <= layer5_outputs(1975);
    layer6_outputs(1589) <= not(layer5_outputs(1212));
    layer6_outputs(1590) <= not(layer5_outputs(44));
    layer6_outputs(1591) <= (layer5_outputs(2306)) or (layer5_outputs(995));
    layer6_outputs(1592) <= layer5_outputs(217);
    layer6_outputs(1593) <= (layer5_outputs(1365)) xor (layer5_outputs(813));
    layer6_outputs(1594) <= (layer5_outputs(2485)) xor (layer5_outputs(905));
    layer6_outputs(1595) <= not(layer5_outputs(390));
    layer6_outputs(1596) <= not(layer5_outputs(659));
    layer6_outputs(1597) <= not(layer5_outputs(1610));
    layer6_outputs(1598) <= not(layer5_outputs(943));
    layer6_outputs(1599) <= (layer5_outputs(427)) and not (layer5_outputs(1037));
    layer6_outputs(1600) <= layer5_outputs(661);
    layer6_outputs(1601) <= layer5_outputs(1414);
    layer6_outputs(1602) <= not((layer5_outputs(1222)) xor (layer5_outputs(2406)));
    layer6_outputs(1603) <= layer5_outputs(1894);
    layer6_outputs(1604) <= layer5_outputs(260);
    layer6_outputs(1605) <= not(layer5_outputs(716));
    layer6_outputs(1606) <= not(layer5_outputs(58));
    layer6_outputs(1607) <= not((layer5_outputs(365)) and (layer5_outputs(932)));
    layer6_outputs(1608) <= (layer5_outputs(2474)) and (layer5_outputs(2083));
    layer6_outputs(1609) <= not(layer5_outputs(2432));
    layer6_outputs(1610) <= layer5_outputs(1891);
    layer6_outputs(1611) <= (layer5_outputs(786)) or (layer5_outputs(419));
    layer6_outputs(1612) <= not((layer5_outputs(843)) xor (layer5_outputs(328)));
    layer6_outputs(1613) <= not(layer5_outputs(831));
    layer6_outputs(1614) <= layer5_outputs(138);
    layer6_outputs(1615) <= not(layer5_outputs(2423)) or (layer5_outputs(2388));
    layer6_outputs(1616) <= not(layer5_outputs(2559));
    layer6_outputs(1617) <= not(layer5_outputs(1191));
    layer6_outputs(1618) <= layer5_outputs(412);
    layer6_outputs(1619) <= not((layer5_outputs(1745)) and (layer5_outputs(2255)));
    layer6_outputs(1620) <= not((layer5_outputs(757)) and (layer5_outputs(366)));
    layer6_outputs(1621) <= not((layer5_outputs(2212)) and (layer5_outputs(541)));
    layer6_outputs(1622) <= (layer5_outputs(119)) xor (layer5_outputs(8));
    layer6_outputs(1623) <= not(layer5_outputs(159));
    layer6_outputs(1624) <= (layer5_outputs(460)) and (layer5_outputs(1686));
    layer6_outputs(1625) <= layer5_outputs(1836);
    layer6_outputs(1626) <= not(layer5_outputs(1955));
    layer6_outputs(1627) <= (layer5_outputs(2016)) and not (layer5_outputs(253));
    layer6_outputs(1628) <= layer5_outputs(710);
    layer6_outputs(1629) <= '1';
    layer6_outputs(1630) <= layer5_outputs(1881);
    layer6_outputs(1631) <= '1';
    layer6_outputs(1632) <= layer5_outputs(1658);
    layer6_outputs(1633) <= layer5_outputs(1418);
    layer6_outputs(1634) <= not(layer5_outputs(1701));
    layer6_outputs(1635) <= (layer5_outputs(945)) and (layer5_outputs(1608));
    layer6_outputs(1636) <= not(layer5_outputs(1205)) or (layer5_outputs(298));
    layer6_outputs(1637) <= layer5_outputs(1334);
    layer6_outputs(1638) <= not((layer5_outputs(1184)) or (layer5_outputs(1167)));
    layer6_outputs(1639) <= not(layer5_outputs(584));
    layer6_outputs(1640) <= not((layer5_outputs(1103)) or (layer5_outputs(1906)));
    layer6_outputs(1641) <= (layer5_outputs(742)) and (layer5_outputs(1442));
    layer6_outputs(1642) <= not((layer5_outputs(112)) and (layer5_outputs(659)));
    layer6_outputs(1643) <= not(layer5_outputs(1595));
    layer6_outputs(1644) <= layer5_outputs(242);
    layer6_outputs(1645) <= not(layer5_outputs(845));
    layer6_outputs(1646) <= not(layer5_outputs(1840));
    layer6_outputs(1647) <= not(layer5_outputs(971)) or (layer5_outputs(2296));
    layer6_outputs(1648) <= layer5_outputs(834);
    layer6_outputs(1649) <= not(layer5_outputs(710));
    layer6_outputs(1650) <= layer5_outputs(2098);
    layer6_outputs(1651) <= not((layer5_outputs(1489)) xor (layer5_outputs(840)));
    layer6_outputs(1652) <= (layer5_outputs(1477)) or (layer5_outputs(646));
    layer6_outputs(1653) <= (layer5_outputs(1329)) and (layer5_outputs(2096));
    layer6_outputs(1654) <= (layer5_outputs(745)) and (layer5_outputs(224));
    layer6_outputs(1655) <= not(layer5_outputs(2188)) or (layer5_outputs(934));
    layer6_outputs(1656) <= layer5_outputs(727);
    layer6_outputs(1657) <= layer5_outputs(1502);
    layer6_outputs(1658) <= not(layer5_outputs(158));
    layer6_outputs(1659) <= layer5_outputs(634);
    layer6_outputs(1660) <= not(layer5_outputs(1257));
    layer6_outputs(1661) <= (layer5_outputs(1500)) or (layer5_outputs(1128));
    layer6_outputs(1662) <= layer5_outputs(95);
    layer6_outputs(1663) <= (layer5_outputs(1666)) and (layer5_outputs(1490));
    layer6_outputs(1664) <= (layer5_outputs(406)) xor (layer5_outputs(1916));
    layer6_outputs(1665) <= not(layer5_outputs(1466));
    layer6_outputs(1666) <= not(layer5_outputs(2534));
    layer6_outputs(1667) <= (layer5_outputs(865)) or (layer5_outputs(910));
    layer6_outputs(1668) <= (layer5_outputs(553)) and not (layer5_outputs(1594));
    layer6_outputs(1669) <= not(layer5_outputs(1749));
    layer6_outputs(1670) <= layer5_outputs(92);
    layer6_outputs(1671) <= (layer5_outputs(216)) and not (layer5_outputs(1564));
    layer6_outputs(1672) <= (layer5_outputs(476)) or (layer5_outputs(61));
    layer6_outputs(1673) <= (layer5_outputs(1484)) and (layer5_outputs(148));
    layer6_outputs(1674) <= not(layer5_outputs(885));
    layer6_outputs(1675) <= not(layer5_outputs(609));
    layer6_outputs(1676) <= (layer5_outputs(2195)) and not (layer5_outputs(2256));
    layer6_outputs(1677) <= not(layer5_outputs(555));
    layer6_outputs(1678) <= not(layer5_outputs(1806));
    layer6_outputs(1679) <= (layer5_outputs(206)) xor (layer5_outputs(1951));
    layer6_outputs(1680) <= (layer5_outputs(994)) and not (layer5_outputs(1717));
    layer6_outputs(1681) <= not((layer5_outputs(1067)) xor (layer5_outputs(999)));
    layer6_outputs(1682) <= not(layer5_outputs(1280)) or (layer5_outputs(1425));
    layer6_outputs(1683) <= (layer5_outputs(1753)) and not (layer5_outputs(1911));
    layer6_outputs(1684) <= not(layer5_outputs(1325)) or (layer5_outputs(218));
    layer6_outputs(1685) <= layer5_outputs(1971);
    layer6_outputs(1686) <= layer5_outputs(1713);
    layer6_outputs(1687) <= layer5_outputs(25);
    layer6_outputs(1688) <= not(layer5_outputs(800));
    layer6_outputs(1689) <= layer5_outputs(1056);
    layer6_outputs(1690) <= not((layer5_outputs(2193)) and (layer5_outputs(2477)));
    layer6_outputs(1691) <= layer5_outputs(629);
    layer6_outputs(1692) <= (layer5_outputs(416)) xor (layer5_outputs(100));
    layer6_outputs(1693) <= not((layer5_outputs(1759)) or (layer5_outputs(317)));
    layer6_outputs(1694) <= layer5_outputs(426);
    layer6_outputs(1695) <= (layer5_outputs(1622)) or (layer5_outputs(84));
    layer6_outputs(1696) <= (layer5_outputs(2482)) or (layer5_outputs(802));
    layer6_outputs(1697) <= (layer5_outputs(1900)) and not (layer5_outputs(946));
    layer6_outputs(1698) <= not(layer5_outputs(649));
    layer6_outputs(1699) <= layer5_outputs(1750);
    layer6_outputs(1700) <= '1';
    layer6_outputs(1701) <= layer5_outputs(1349);
    layer6_outputs(1702) <= not(layer5_outputs(1370)) or (layer5_outputs(2505));
    layer6_outputs(1703) <= not(layer5_outputs(1752));
    layer6_outputs(1704) <= not((layer5_outputs(2308)) xor (layer5_outputs(1990)));
    layer6_outputs(1705) <= not(layer5_outputs(528));
    layer6_outputs(1706) <= not((layer5_outputs(935)) and (layer5_outputs(363)));
    layer6_outputs(1707) <= layer5_outputs(1567);
    layer6_outputs(1708) <= layer5_outputs(1242);
    layer6_outputs(1709) <= (layer5_outputs(302)) xor (layer5_outputs(2502));
    layer6_outputs(1710) <= (layer5_outputs(2432)) and not (layer5_outputs(82));
    layer6_outputs(1711) <= layer5_outputs(910);
    layer6_outputs(1712) <= not(layer5_outputs(1348));
    layer6_outputs(1713) <= '0';
    layer6_outputs(1714) <= layer5_outputs(1587);
    layer6_outputs(1715) <= layer5_outputs(1583);
    layer6_outputs(1716) <= layer5_outputs(2266);
    layer6_outputs(1717) <= (layer5_outputs(2283)) and (layer5_outputs(1456));
    layer6_outputs(1718) <= (layer5_outputs(1829)) and (layer5_outputs(2085));
    layer6_outputs(1719) <= not(layer5_outputs(2377)) or (layer5_outputs(621));
    layer6_outputs(1720) <= layer5_outputs(628);
    layer6_outputs(1721) <= layer5_outputs(2545);
    layer6_outputs(1722) <= not(layer5_outputs(91));
    layer6_outputs(1723) <= (layer5_outputs(1861)) and (layer5_outputs(1315));
    layer6_outputs(1724) <= not(layer5_outputs(806));
    layer6_outputs(1725) <= layer5_outputs(1715);
    layer6_outputs(1726) <= (layer5_outputs(465)) and not (layer5_outputs(1431));
    layer6_outputs(1727) <= layer5_outputs(1354);
    layer6_outputs(1728) <= not(layer5_outputs(904));
    layer6_outputs(1729) <= not(layer5_outputs(871));
    layer6_outputs(1730) <= layer5_outputs(1019);
    layer6_outputs(1731) <= not(layer5_outputs(596));
    layer6_outputs(1732) <= not(layer5_outputs(1424));
    layer6_outputs(1733) <= not(layer5_outputs(1237)) or (layer5_outputs(399));
    layer6_outputs(1734) <= not(layer5_outputs(356));
    layer6_outputs(1735) <= not(layer5_outputs(906));
    layer6_outputs(1736) <= not((layer5_outputs(2125)) or (layer5_outputs(595)));
    layer6_outputs(1737) <= (layer5_outputs(780)) and not (layer5_outputs(1227));
    layer6_outputs(1738) <= (layer5_outputs(1565)) or (layer5_outputs(547));
    layer6_outputs(1739) <= not((layer5_outputs(2546)) and (layer5_outputs(1648)));
    layer6_outputs(1740) <= not((layer5_outputs(203)) and (layer5_outputs(2028)));
    layer6_outputs(1741) <= not((layer5_outputs(2241)) or (layer5_outputs(114)));
    layer6_outputs(1742) <= not(layer5_outputs(2410));
    layer6_outputs(1743) <= not((layer5_outputs(1517)) xor (layer5_outputs(1953)));
    layer6_outputs(1744) <= not((layer5_outputs(1675)) and (layer5_outputs(1611)));
    layer6_outputs(1745) <= not((layer5_outputs(960)) xor (layer5_outputs(1268)));
    layer6_outputs(1746) <= not(layer5_outputs(784));
    layer6_outputs(1747) <= (layer5_outputs(46)) or (layer5_outputs(606));
    layer6_outputs(1748) <= not((layer5_outputs(1235)) xor (layer5_outputs(1156)));
    layer6_outputs(1749) <= layer5_outputs(7);
    layer6_outputs(1750) <= layer5_outputs(1044);
    layer6_outputs(1751) <= layer5_outputs(2118);
    layer6_outputs(1752) <= layer5_outputs(1150);
    layer6_outputs(1753) <= not((layer5_outputs(960)) xor (layer5_outputs(525)));
    layer6_outputs(1754) <= (layer5_outputs(1522)) and not (layer5_outputs(665));
    layer6_outputs(1755) <= not(layer5_outputs(1655));
    layer6_outputs(1756) <= layer5_outputs(964);
    layer6_outputs(1757) <= layer5_outputs(972);
    layer6_outputs(1758) <= (layer5_outputs(2049)) and not (layer5_outputs(2003));
    layer6_outputs(1759) <= (layer5_outputs(155)) xor (layer5_outputs(187));
    layer6_outputs(1760) <= not((layer5_outputs(123)) and (layer5_outputs(71)));
    layer6_outputs(1761) <= (layer5_outputs(2353)) or (layer5_outputs(1823));
    layer6_outputs(1762) <= layer5_outputs(990);
    layer6_outputs(1763) <= not(layer5_outputs(682));
    layer6_outputs(1764) <= (layer5_outputs(1384)) xor (layer5_outputs(2529));
    layer6_outputs(1765) <= not((layer5_outputs(2101)) or (layer5_outputs(1159)));
    layer6_outputs(1766) <= (layer5_outputs(284)) and not (layer5_outputs(1785));
    layer6_outputs(1767) <= (layer5_outputs(2287)) or (layer5_outputs(2544));
    layer6_outputs(1768) <= (layer5_outputs(2329)) and (layer5_outputs(1548));
    layer6_outputs(1769) <= (layer5_outputs(486)) and not (layer5_outputs(1148));
    layer6_outputs(1770) <= layer5_outputs(1850);
    layer6_outputs(1771) <= not((layer5_outputs(1712)) xor (layer5_outputs(2129)));
    layer6_outputs(1772) <= not((layer5_outputs(292)) and (layer5_outputs(1856)));
    layer6_outputs(1773) <= (layer5_outputs(1877)) and (layer5_outputs(12));
    layer6_outputs(1774) <= not(layer5_outputs(1107));
    layer6_outputs(1775) <= not((layer5_outputs(1269)) and (layer5_outputs(1765)));
    layer6_outputs(1776) <= (layer5_outputs(2038)) and not (layer5_outputs(2473));
    layer6_outputs(1777) <= (layer5_outputs(2181)) and not (layer5_outputs(985));
    layer6_outputs(1778) <= layer5_outputs(1994);
    layer6_outputs(1779) <= layer5_outputs(241);
    layer6_outputs(1780) <= not(layer5_outputs(2390));
    layer6_outputs(1781) <= (layer5_outputs(2533)) and not (layer5_outputs(18));
    layer6_outputs(1782) <= (layer5_outputs(1766)) and (layer5_outputs(272));
    layer6_outputs(1783) <= not((layer5_outputs(293)) or (layer5_outputs(585)));
    layer6_outputs(1784) <= not((layer5_outputs(1470)) xor (layer5_outputs(2289)));
    layer6_outputs(1785) <= not(layer5_outputs(253));
    layer6_outputs(1786) <= not(layer5_outputs(2195)) or (layer5_outputs(2125));
    layer6_outputs(1787) <= layer5_outputs(183);
    layer6_outputs(1788) <= layer5_outputs(2422);
    layer6_outputs(1789) <= (layer5_outputs(782)) and not (layer5_outputs(592));
    layer6_outputs(1790) <= layer5_outputs(917);
    layer6_outputs(1791) <= layer5_outputs(119);
    layer6_outputs(1792) <= not(layer5_outputs(1000));
    layer6_outputs(1793) <= not(layer5_outputs(2141));
    layer6_outputs(1794) <= (layer5_outputs(916)) or (layer5_outputs(1177));
    layer6_outputs(1795) <= (layer5_outputs(795)) or (layer5_outputs(2253));
    layer6_outputs(1796) <= (layer5_outputs(2472)) and not (layer5_outputs(1865));
    layer6_outputs(1797) <= not(layer5_outputs(371));
    layer6_outputs(1798) <= not(layer5_outputs(2523)) or (layer5_outputs(36));
    layer6_outputs(1799) <= layer5_outputs(1421);
    layer6_outputs(1800) <= not(layer5_outputs(1067)) or (layer5_outputs(2018));
    layer6_outputs(1801) <= (layer5_outputs(2450)) or (layer5_outputs(1834));
    layer6_outputs(1802) <= not(layer5_outputs(308));
    layer6_outputs(1803) <= not(layer5_outputs(1776));
    layer6_outputs(1804) <= not((layer5_outputs(2478)) xor (layer5_outputs(726)));
    layer6_outputs(1805) <= layer5_outputs(343);
    layer6_outputs(1806) <= not(layer5_outputs(2022)) or (layer5_outputs(1717));
    layer6_outputs(1807) <= (layer5_outputs(501)) and not (layer5_outputs(1426));
    layer6_outputs(1808) <= not((layer5_outputs(1267)) and (layer5_outputs(1057)));
    layer6_outputs(1809) <= layer5_outputs(1449);
    layer6_outputs(1810) <= not((layer5_outputs(102)) xor (layer5_outputs(541)));
    layer6_outputs(1811) <= not(layer5_outputs(686));
    layer6_outputs(1812) <= layer5_outputs(667);
    layer6_outputs(1813) <= layer5_outputs(2435);
    layer6_outputs(1814) <= not((layer5_outputs(1450)) xor (layer5_outputs(2215)));
    layer6_outputs(1815) <= not(layer5_outputs(870));
    layer6_outputs(1816) <= not((layer5_outputs(1292)) xor (layer5_outputs(2349)));
    layer6_outputs(1817) <= layer5_outputs(1039);
    layer6_outputs(1818) <= layer5_outputs(205);
    layer6_outputs(1819) <= not(layer5_outputs(514));
    layer6_outputs(1820) <= layer5_outputs(1998);
    layer6_outputs(1821) <= not((layer5_outputs(1649)) or (layer5_outputs(2379)));
    layer6_outputs(1822) <= not((layer5_outputs(2510)) or (layer5_outputs(2299)));
    layer6_outputs(1823) <= not(layer5_outputs(1727));
    layer6_outputs(1824) <= not(layer5_outputs(690)) or (layer5_outputs(1001));
    layer6_outputs(1825) <= layer5_outputs(2106);
    layer6_outputs(1826) <= (layer5_outputs(126)) or (layer5_outputs(1769));
    layer6_outputs(1827) <= not(layer5_outputs(1313));
    layer6_outputs(1828) <= layer5_outputs(2417);
    layer6_outputs(1829) <= not(layer5_outputs(1162));
    layer6_outputs(1830) <= layer5_outputs(1520);
    layer6_outputs(1831) <= not(layer5_outputs(732));
    layer6_outputs(1832) <= not(layer5_outputs(1096));
    layer6_outputs(1833) <= layer5_outputs(1335);
    layer6_outputs(1834) <= not(layer5_outputs(2202)) or (layer5_outputs(2159));
    layer6_outputs(1835) <= not(layer5_outputs(1747));
    layer6_outputs(1836) <= layer5_outputs(2336);
    layer6_outputs(1837) <= (layer5_outputs(1938)) and not (layer5_outputs(1526));
    layer6_outputs(1838) <= layer5_outputs(362);
    layer6_outputs(1839) <= layer5_outputs(2241);
    layer6_outputs(1840) <= layer5_outputs(2343);
    layer6_outputs(1841) <= layer5_outputs(359);
    layer6_outputs(1842) <= layer5_outputs(2252);
    layer6_outputs(1843) <= not(layer5_outputs(1557));
    layer6_outputs(1844) <= not((layer5_outputs(886)) or (layer5_outputs(2492)));
    layer6_outputs(1845) <= (layer5_outputs(754)) and not (layer5_outputs(2436));
    layer6_outputs(1846) <= not(layer5_outputs(1159)) or (layer5_outputs(157));
    layer6_outputs(1847) <= (layer5_outputs(1110)) and not (layer5_outputs(775));
    layer6_outputs(1848) <= (layer5_outputs(2031)) and (layer5_outputs(1419));
    layer6_outputs(1849) <= layer5_outputs(2089);
    layer6_outputs(1850) <= not(layer5_outputs(2541));
    layer6_outputs(1851) <= layer5_outputs(2436);
    layer6_outputs(1852) <= (layer5_outputs(1131)) or (layer5_outputs(2260));
    layer6_outputs(1853) <= not((layer5_outputs(325)) and (layer5_outputs(1588)));
    layer6_outputs(1854) <= layer5_outputs(544);
    layer6_outputs(1855) <= layer5_outputs(1963);
    layer6_outputs(1856) <= (layer5_outputs(1393)) and not (layer5_outputs(2497));
    layer6_outputs(1857) <= not(layer5_outputs(2276));
    layer6_outputs(1858) <= (layer5_outputs(1102)) and not (layer5_outputs(322));
    layer6_outputs(1859) <= not(layer5_outputs(628)) or (layer5_outputs(450));
    layer6_outputs(1860) <= not(layer5_outputs(2273));
    layer6_outputs(1861) <= not(layer5_outputs(1315)) or (layer5_outputs(2213));
    layer6_outputs(1862) <= not(layer5_outputs(1949)) or (layer5_outputs(793));
    layer6_outputs(1863) <= not(layer5_outputs(280));
    layer6_outputs(1864) <= not(layer5_outputs(1729)) or (layer5_outputs(2451));
    layer6_outputs(1865) <= layer5_outputs(1281);
    layer6_outputs(1866) <= layer5_outputs(579);
    layer6_outputs(1867) <= not((layer5_outputs(1114)) xor (layer5_outputs(477)));
    layer6_outputs(1868) <= not(layer5_outputs(1387)) or (layer5_outputs(2310));
    layer6_outputs(1869) <= layer5_outputs(1121);
    layer6_outputs(1870) <= not((layer5_outputs(1382)) xor (layer5_outputs(2366)));
    layer6_outputs(1871) <= not(layer5_outputs(576));
    layer6_outputs(1872) <= layer5_outputs(90);
    layer6_outputs(1873) <= not(layer5_outputs(1165));
    layer6_outputs(1874) <= not(layer5_outputs(352)) or (layer5_outputs(600));
    layer6_outputs(1875) <= not(layer5_outputs(1843));
    layer6_outputs(1876) <= not(layer5_outputs(827));
    layer6_outputs(1877) <= layer5_outputs(483);
    layer6_outputs(1878) <= layer5_outputs(1662);
    layer6_outputs(1879) <= not(layer5_outputs(371));
    layer6_outputs(1880) <= not((layer5_outputs(1263)) or (layer5_outputs(925)));
    layer6_outputs(1881) <= not(layer5_outputs(2558)) or (layer5_outputs(1930));
    layer6_outputs(1882) <= (layer5_outputs(1271)) and (layer5_outputs(1972));
    layer6_outputs(1883) <= (layer5_outputs(2075)) and (layer5_outputs(1509));
    layer6_outputs(1884) <= not((layer5_outputs(2294)) and (layer5_outputs(148)));
    layer6_outputs(1885) <= not(layer5_outputs(386));
    layer6_outputs(1886) <= not((layer5_outputs(24)) or (layer5_outputs(1135)));
    layer6_outputs(1887) <= (layer5_outputs(487)) xor (layer5_outputs(1720));
    layer6_outputs(1888) <= not((layer5_outputs(1742)) and (layer5_outputs(1105)));
    layer6_outputs(1889) <= not(layer5_outputs(1150));
    layer6_outputs(1890) <= (layer5_outputs(288)) and not (layer5_outputs(2384));
    layer6_outputs(1891) <= not(layer5_outputs(1988));
    layer6_outputs(1892) <= not(layer5_outputs(855));
    layer6_outputs(1893) <= not(layer5_outputs(2302));
    layer6_outputs(1894) <= not((layer5_outputs(457)) and (layer5_outputs(914)));
    layer6_outputs(1895) <= not(layer5_outputs(2409));
    layer6_outputs(1896) <= not(layer5_outputs(2091));
    layer6_outputs(1897) <= not((layer5_outputs(1718)) xor (layer5_outputs(2501)));
    layer6_outputs(1898) <= layer5_outputs(442);
    layer6_outputs(1899) <= layer5_outputs(1779);
    layer6_outputs(1900) <= layer5_outputs(2352);
    layer6_outputs(1901) <= not(layer5_outputs(818)) or (layer5_outputs(790));
    layer6_outputs(1902) <= not(layer5_outputs(731));
    layer6_outputs(1903) <= not((layer5_outputs(1323)) and (layer5_outputs(456)));
    layer6_outputs(1904) <= layer5_outputs(196);
    layer6_outputs(1905) <= layer5_outputs(2258);
    layer6_outputs(1906) <= (layer5_outputs(847)) xor (layer5_outputs(959));
    layer6_outputs(1907) <= layer5_outputs(1682);
    layer6_outputs(1908) <= layer5_outputs(2349);
    layer6_outputs(1909) <= not(layer5_outputs(81));
    layer6_outputs(1910) <= not(layer5_outputs(1723)) or (layer5_outputs(1801));
    layer6_outputs(1911) <= layer5_outputs(634);
    layer6_outputs(1912) <= (layer5_outputs(372)) and not (layer5_outputs(2357));
    layer6_outputs(1913) <= layer5_outputs(300);
    layer6_outputs(1914) <= (layer5_outputs(1708)) and not (layer5_outputs(467));
    layer6_outputs(1915) <= (layer5_outputs(803)) xor (layer5_outputs(1575));
    layer6_outputs(1916) <= layer5_outputs(150);
    layer6_outputs(1917) <= layer5_outputs(2531);
    layer6_outputs(1918) <= (layer5_outputs(464)) and not (layer5_outputs(1705));
    layer6_outputs(1919) <= '1';
    layer6_outputs(1920) <= (layer5_outputs(1101)) and not (layer5_outputs(1893));
    layer6_outputs(1921) <= (layer5_outputs(2355)) and not (layer5_outputs(1504));
    layer6_outputs(1922) <= not((layer5_outputs(1677)) and (layer5_outputs(637)));
    layer6_outputs(1923) <= not(layer5_outputs(1670)) or (layer5_outputs(2286));
    layer6_outputs(1924) <= layer5_outputs(420);
    layer6_outputs(1925) <= not((layer5_outputs(1210)) xor (layer5_outputs(1241)));
    layer6_outputs(1926) <= not(layer5_outputs(896));
    layer6_outputs(1927) <= not(layer5_outputs(2282));
    layer6_outputs(1928) <= not((layer5_outputs(504)) and (layer5_outputs(1447)));
    layer6_outputs(1929) <= not(layer5_outputs(307));
    layer6_outputs(1930) <= not(layer5_outputs(2209));
    layer6_outputs(1931) <= not(layer5_outputs(1607));
    layer6_outputs(1932) <= (layer5_outputs(1616)) or (layer5_outputs(1168));
    layer6_outputs(1933) <= (layer5_outputs(2380)) and (layer5_outputs(11));
    layer6_outputs(1934) <= not(layer5_outputs(156));
    layer6_outputs(1935) <= not(layer5_outputs(2391));
    layer6_outputs(1936) <= not((layer5_outputs(359)) and (layer5_outputs(957)));
    layer6_outputs(1937) <= (layer5_outputs(188)) and not (layer5_outputs(1402));
    layer6_outputs(1938) <= layer5_outputs(549);
    layer6_outputs(1939) <= not(layer5_outputs(788));
    layer6_outputs(1940) <= not(layer5_outputs(417));
    layer6_outputs(1941) <= not((layer5_outputs(790)) xor (layer5_outputs(1439)));
    layer6_outputs(1942) <= (layer5_outputs(449)) xor (layer5_outputs(1635));
    layer6_outputs(1943) <= not((layer5_outputs(933)) and (layer5_outputs(1710)));
    layer6_outputs(1944) <= not(layer5_outputs(2273));
    layer6_outputs(1945) <= (layer5_outputs(2552)) xor (layer5_outputs(1669));
    layer6_outputs(1946) <= '1';
    layer6_outputs(1947) <= not(layer5_outputs(2166)) or (layer5_outputs(771));
    layer6_outputs(1948) <= not(layer5_outputs(2511)) or (layer5_outputs(303));
    layer6_outputs(1949) <= not(layer5_outputs(633));
    layer6_outputs(1950) <= (layer5_outputs(2146)) and not (layer5_outputs(1433));
    layer6_outputs(1951) <= not((layer5_outputs(1086)) xor (layer5_outputs(2327)));
    layer6_outputs(1952) <= not(layer5_outputs(807));
    layer6_outputs(1953) <= not(layer5_outputs(944)) or (layer5_outputs(2459));
    layer6_outputs(1954) <= (layer5_outputs(1456)) and not (layer5_outputs(1332));
    layer6_outputs(1955) <= layer5_outputs(897);
    layer6_outputs(1956) <= not(layer5_outputs(517));
    layer6_outputs(1957) <= layer5_outputs(1009);
    layer6_outputs(1958) <= (layer5_outputs(1876)) xor (layer5_outputs(1940));
    layer6_outputs(1959) <= (layer5_outputs(563)) xor (layer5_outputs(312));
    layer6_outputs(1960) <= '0';
    layer6_outputs(1961) <= not((layer5_outputs(1266)) or (layer5_outputs(1804)));
    layer6_outputs(1962) <= not(layer5_outputs(1372)) or (layer5_outputs(1643));
    layer6_outputs(1963) <= layer5_outputs(1546);
    layer6_outputs(1964) <= '1';
    layer6_outputs(1965) <= not(layer5_outputs(1077));
    layer6_outputs(1966) <= not(layer5_outputs(459));
    layer6_outputs(1967) <= (layer5_outputs(1299)) xor (layer5_outputs(289));
    layer6_outputs(1968) <= '1';
    layer6_outputs(1969) <= not((layer5_outputs(368)) and (layer5_outputs(1706)));
    layer6_outputs(1970) <= '1';
    layer6_outputs(1971) <= not(layer5_outputs(1101));
    layer6_outputs(1972) <= not(layer5_outputs(2307));
    layer6_outputs(1973) <= layer5_outputs(1261);
    layer6_outputs(1974) <= not(layer5_outputs(2499));
    layer6_outputs(1975) <= layer5_outputs(836);
    layer6_outputs(1976) <= not((layer5_outputs(2491)) xor (layer5_outputs(1402)));
    layer6_outputs(1977) <= not(layer5_outputs(701));
    layer6_outputs(1978) <= not(layer5_outputs(1008));
    layer6_outputs(1979) <= layer5_outputs(1731);
    layer6_outputs(1980) <= not((layer5_outputs(1120)) or (layer5_outputs(1046)));
    layer6_outputs(1981) <= not((layer5_outputs(2484)) or (layer5_outputs(2430)));
    layer6_outputs(1982) <= (layer5_outputs(1874)) xor (layer5_outputs(1612));
    layer6_outputs(1983) <= layer5_outputs(1282);
    layer6_outputs(1984) <= not(layer5_outputs(207));
    layer6_outputs(1985) <= (layer5_outputs(1599)) xor (layer5_outputs(2083));
    layer6_outputs(1986) <= not((layer5_outputs(1012)) xor (layer5_outputs(1852)));
    layer6_outputs(1987) <= not((layer5_outputs(291)) or (layer5_outputs(1180)));
    layer6_outputs(1988) <= not((layer5_outputs(506)) xor (layer5_outputs(1485)));
    layer6_outputs(1989) <= layer5_outputs(1685);
    layer6_outputs(1990) <= not(layer5_outputs(1787));
    layer6_outputs(1991) <= layer5_outputs(0);
    layer6_outputs(1992) <= not(layer5_outputs(1940)) or (layer5_outputs(321));
    layer6_outputs(1993) <= not((layer5_outputs(1396)) and (layer5_outputs(2489)));
    layer6_outputs(1994) <= not((layer5_outputs(382)) or (layer5_outputs(2511)));
    layer6_outputs(1995) <= layer5_outputs(399);
    layer6_outputs(1996) <= not((layer5_outputs(362)) or (layer5_outputs(567)));
    layer6_outputs(1997) <= not((layer5_outputs(720)) and (layer5_outputs(1871)));
    layer6_outputs(1998) <= (layer5_outputs(2291)) and not (layer5_outputs(232));
    layer6_outputs(1999) <= not(layer5_outputs(231));
    layer6_outputs(2000) <= layer5_outputs(1000);
    layer6_outputs(2001) <= not((layer5_outputs(887)) or (layer5_outputs(1262)));
    layer6_outputs(2002) <= (layer5_outputs(860)) xor (layer5_outputs(145));
    layer6_outputs(2003) <= not((layer5_outputs(1627)) or (layer5_outputs(185)));
    layer6_outputs(2004) <= not(layer5_outputs(1054)) or (layer5_outputs(1091));
    layer6_outputs(2005) <= not((layer5_outputs(382)) or (layer5_outputs(682)));
    layer6_outputs(2006) <= not(layer5_outputs(1496)) or (layer5_outputs(2055));
    layer6_outputs(2007) <= not(layer5_outputs(1486)) or (layer5_outputs(693));
    layer6_outputs(2008) <= (layer5_outputs(2131)) and not (layer5_outputs(888));
    layer6_outputs(2009) <= layer5_outputs(1810);
    layer6_outputs(2010) <= layer5_outputs(2135);
    layer6_outputs(2011) <= not(layer5_outputs(1099));
    layer6_outputs(2012) <= not((layer5_outputs(1879)) xor (layer5_outputs(1849)));
    layer6_outputs(2013) <= not((layer5_outputs(1120)) xor (layer5_outputs(509)));
    layer6_outputs(2014) <= not(layer5_outputs(318));
    layer6_outputs(2015) <= (layer5_outputs(208)) xor (layer5_outputs(1741));
    layer6_outputs(2016) <= '1';
    layer6_outputs(2017) <= not(layer5_outputs(2460)) or (layer5_outputs(206));
    layer6_outputs(2018) <= layer5_outputs(900);
    layer6_outputs(2019) <= (layer5_outputs(1736)) and (layer5_outputs(1981));
    layer6_outputs(2020) <= not(layer5_outputs(977));
    layer6_outputs(2021) <= not(layer5_outputs(1924));
    layer6_outputs(2022) <= layer5_outputs(1510);
    layer6_outputs(2023) <= not(layer5_outputs(1345));
    layer6_outputs(2024) <= not(layer5_outputs(966));
    layer6_outputs(2025) <= (layer5_outputs(2428)) xor (layer5_outputs(23));
    layer6_outputs(2026) <= not(layer5_outputs(1574));
    layer6_outputs(2027) <= layer5_outputs(1854);
    layer6_outputs(2028) <= '0';
    layer6_outputs(2029) <= layer5_outputs(2465);
    layer6_outputs(2030) <= layer5_outputs(1588);
    layer6_outputs(2031) <= layer5_outputs(1513);
    layer6_outputs(2032) <= not(layer5_outputs(2161));
    layer6_outputs(2033) <= not(layer5_outputs(1772)) or (layer5_outputs(1875));
    layer6_outputs(2034) <= (layer5_outputs(1080)) and not (layer5_outputs(2205));
    layer6_outputs(2035) <= not(layer5_outputs(813));
    layer6_outputs(2036) <= not(layer5_outputs(1308));
    layer6_outputs(2037) <= '0';
    layer6_outputs(2038) <= not(layer5_outputs(1162));
    layer6_outputs(2039) <= not(layer5_outputs(922));
    layer6_outputs(2040) <= not(layer5_outputs(758));
    layer6_outputs(2041) <= layer5_outputs(587);
    layer6_outputs(2042) <= not(layer5_outputs(1029)) or (layer5_outputs(155));
    layer6_outputs(2043) <= layer5_outputs(2218);
    layer6_outputs(2044) <= layer5_outputs(2231);
    layer6_outputs(2045) <= (layer5_outputs(513)) and (layer5_outputs(513));
    layer6_outputs(2046) <= not((layer5_outputs(2424)) and (layer5_outputs(2006)));
    layer6_outputs(2047) <= not(layer5_outputs(1702));
    layer6_outputs(2048) <= not(layer5_outputs(792)) or (layer5_outputs(2041));
    layer6_outputs(2049) <= not((layer5_outputs(491)) xor (layer5_outputs(618)));
    layer6_outputs(2050) <= (layer5_outputs(1064)) and not (layer5_outputs(1824));
    layer6_outputs(2051) <= not(layer5_outputs(270));
    layer6_outputs(2052) <= (layer5_outputs(1664)) and (layer5_outputs(2263));
    layer6_outputs(2053) <= (layer5_outputs(92)) and not (layer5_outputs(2086));
    layer6_outputs(2054) <= layer5_outputs(176);
    layer6_outputs(2055) <= (layer5_outputs(1730)) xor (layer5_outputs(49));
    layer6_outputs(2056) <= not(layer5_outputs(968));
    layer6_outputs(2057) <= not(layer5_outputs(1551)) or (layer5_outputs(1917));
    layer6_outputs(2058) <= not(layer5_outputs(916));
    layer6_outputs(2059) <= layer5_outputs(2540);
    layer6_outputs(2060) <= (layer5_outputs(947)) and not (layer5_outputs(789));
    layer6_outputs(2061) <= not(layer5_outputs(269));
    layer6_outputs(2062) <= not(layer5_outputs(689));
    layer6_outputs(2063) <= not((layer5_outputs(429)) or (layer5_outputs(1651)));
    layer6_outputs(2064) <= (layer5_outputs(1889)) xor (layer5_outputs(976));
    layer6_outputs(2065) <= not(layer5_outputs(1252)) or (layer5_outputs(773));
    layer6_outputs(2066) <= not(layer5_outputs(2091)) or (layer5_outputs(753));
    layer6_outputs(2067) <= not((layer5_outputs(1884)) and (layer5_outputs(865)));
    layer6_outputs(2068) <= (layer5_outputs(1641)) and not (layer5_outputs(1012));
    layer6_outputs(2069) <= not(layer5_outputs(222));
    layer6_outputs(2070) <= not((layer5_outputs(2471)) xor (layer5_outputs(2328)));
    layer6_outputs(2071) <= not(layer5_outputs(945));
    layer6_outputs(2072) <= (layer5_outputs(917)) and (layer5_outputs(415));
    layer6_outputs(2073) <= layer5_outputs(1773);
    layer6_outputs(2074) <= not(layer5_outputs(953));
    layer6_outputs(2075) <= not(layer5_outputs(2027));
    layer6_outputs(2076) <= (layer5_outputs(492)) or (layer5_outputs(1830));
    layer6_outputs(2077) <= not((layer5_outputs(1210)) xor (layer5_outputs(864)));
    layer6_outputs(2078) <= not((layer5_outputs(538)) or (layer5_outputs(954)));
    layer6_outputs(2079) <= not((layer5_outputs(1089)) or (layer5_outputs(1582)));
    layer6_outputs(2080) <= not(layer5_outputs(1613));
    layer6_outputs(2081) <= '1';
    layer6_outputs(2082) <= not(layer5_outputs(534));
    layer6_outputs(2083) <= not(layer5_outputs(1838)) or (layer5_outputs(2011));
    layer6_outputs(2084) <= not(layer5_outputs(683));
    layer6_outputs(2085) <= not(layer5_outputs(1075));
    layer6_outputs(2086) <= not(layer5_outputs(521)) or (layer5_outputs(1978));
    layer6_outputs(2087) <= not((layer5_outputs(1630)) and (layer5_outputs(12)));
    layer6_outputs(2088) <= not(layer5_outputs(1228)) or (layer5_outputs(2302));
    layer6_outputs(2089) <= (layer5_outputs(1866)) xor (layer5_outputs(2001));
    layer6_outputs(2090) <= (layer5_outputs(2361)) xor (layer5_outputs(1579));
    layer6_outputs(2091) <= not(layer5_outputs(1464));
    layer6_outputs(2092) <= layer5_outputs(929);
    layer6_outputs(2093) <= layer5_outputs(2142);
    layer6_outputs(2094) <= not(layer5_outputs(273));
    layer6_outputs(2095) <= layer5_outputs(1633);
    layer6_outputs(2096) <= not((layer5_outputs(370)) xor (layer5_outputs(1225)));
    layer6_outputs(2097) <= (layer5_outputs(443)) and not (layer5_outputs(16));
    layer6_outputs(2098) <= not((layer5_outputs(117)) xor (layer5_outputs(2061)));
    layer6_outputs(2099) <= layer5_outputs(297);
    layer6_outputs(2100) <= layer5_outputs(2376);
    layer6_outputs(2101) <= not(layer5_outputs(316));
    layer6_outputs(2102) <= not(layer5_outputs(1275));
    layer6_outputs(2103) <= not(layer5_outputs(1258));
    layer6_outputs(2104) <= not(layer5_outputs(769));
    layer6_outputs(2105) <= not(layer5_outputs(546));
    layer6_outputs(2106) <= not((layer5_outputs(1470)) xor (layer5_outputs(141)));
    layer6_outputs(2107) <= not(layer5_outputs(2539));
    layer6_outputs(2108) <= layer5_outputs(1192);
    layer6_outputs(2109) <= not((layer5_outputs(380)) xor (layer5_outputs(24)));
    layer6_outputs(2110) <= not(layer5_outputs(2245));
    layer6_outputs(2111) <= not(layer5_outputs(1780));
    layer6_outputs(2112) <= not((layer5_outputs(561)) xor (layer5_outputs(1094)));
    layer6_outputs(2113) <= not((layer5_outputs(2333)) xor (layer5_outputs(2296)));
    layer6_outputs(2114) <= (layer5_outputs(1851)) xor (layer5_outputs(564));
    layer6_outputs(2115) <= not(layer5_outputs(566));
    layer6_outputs(2116) <= layer5_outputs(1144);
    layer6_outputs(2117) <= not((layer5_outputs(451)) or (layer5_outputs(2079)));
    layer6_outputs(2118) <= not((layer5_outputs(703)) or (layer5_outputs(1425)));
    layer6_outputs(2119) <= layer5_outputs(797);
    layer6_outputs(2120) <= not((layer5_outputs(989)) or (layer5_outputs(2543)));
    layer6_outputs(2121) <= layer5_outputs(2322);
    layer6_outputs(2122) <= layer5_outputs(1326);
    layer6_outputs(2123) <= not((layer5_outputs(2251)) xor (layer5_outputs(161)));
    layer6_outputs(2124) <= layer5_outputs(497);
    layer6_outputs(2125) <= not((layer5_outputs(1905)) and (layer5_outputs(193)));
    layer6_outputs(2126) <= layer5_outputs(2265);
    layer6_outputs(2127) <= not((layer5_outputs(1511)) xor (layer5_outputs(985)));
    layer6_outputs(2128) <= layer5_outputs(2272);
    layer6_outputs(2129) <= not((layer5_outputs(1122)) xor (layer5_outputs(590)));
    layer6_outputs(2130) <= layer5_outputs(1603);
    layer6_outputs(2131) <= not((layer5_outputs(610)) xor (layer5_outputs(584)));
    layer6_outputs(2132) <= layer5_outputs(1135);
    layer6_outputs(2133) <= not(layer5_outputs(1615));
    layer6_outputs(2134) <= (layer5_outputs(1831)) and (layer5_outputs(2179));
    layer6_outputs(2135) <= layer5_outputs(259);
    layer6_outputs(2136) <= not((layer5_outputs(597)) and (layer5_outputs(1996)));
    layer6_outputs(2137) <= layer5_outputs(1688);
    layer6_outputs(2138) <= layer5_outputs(1145);
    layer6_outputs(2139) <= not((layer5_outputs(2117)) or (layer5_outputs(552)));
    layer6_outputs(2140) <= layer5_outputs(1084);
    layer6_outputs(2141) <= not(layer5_outputs(1472));
    layer6_outputs(2142) <= not(layer5_outputs(721));
    layer6_outputs(2143) <= layer5_outputs(691);
    layer6_outputs(2144) <= layer5_outputs(2331);
    layer6_outputs(2145) <= not((layer5_outputs(1597)) xor (layer5_outputs(2177)));
    layer6_outputs(2146) <= layer5_outputs(2331);
    layer6_outputs(2147) <= not(layer5_outputs(1656)) or (layer5_outputs(808));
    layer6_outputs(2148) <= not(layer5_outputs(1508));
    layer6_outputs(2149) <= not((layer5_outputs(1939)) xor (layer5_outputs(1141)));
    layer6_outputs(2150) <= (layer5_outputs(2537)) xor (layer5_outputs(1445));
    layer6_outputs(2151) <= (layer5_outputs(176)) and not (layer5_outputs(581));
    layer6_outputs(2152) <= (layer5_outputs(1010)) xor (layer5_outputs(1271));
    layer6_outputs(2153) <= (layer5_outputs(1125)) or (layer5_outputs(1975));
    layer6_outputs(2154) <= not((layer5_outputs(1621)) xor (layer5_outputs(1824)));
    layer6_outputs(2155) <= not(layer5_outputs(2389)) or (layer5_outputs(131));
    layer6_outputs(2156) <= layer5_outputs(2335);
    layer6_outputs(2157) <= layer5_outputs(1207);
    layer6_outputs(2158) <= layer5_outputs(1558);
    layer6_outputs(2159) <= (layer5_outputs(422)) and (layer5_outputs(2071));
    layer6_outputs(2160) <= (layer5_outputs(2342)) and (layer5_outputs(1090));
    layer6_outputs(2161) <= (layer5_outputs(2509)) or (layer5_outputs(1620));
    layer6_outputs(2162) <= layer5_outputs(34);
    layer6_outputs(2163) <= layer5_outputs(1905);
    layer6_outputs(2164) <= (layer5_outputs(2175)) xor (layer5_outputs(191));
    layer6_outputs(2165) <= not(layer5_outputs(229));
    layer6_outputs(2166) <= not((layer5_outputs(88)) xor (layer5_outputs(180)));
    layer6_outputs(2167) <= (layer5_outputs(226)) or (layer5_outputs(1357));
    layer6_outputs(2168) <= not((layer5_outputs(43)) and (layer5_outputs(817)));
    layer6_outputs(2169) <= (layer5_outputs(2425)) and (layer5_outputs(1307));
    layer6_outputs(2170) <= layer5_outputs(1585);
    layer6_outputs(2171) <= (layer5_outputs(239)) xor (layer5_outputs(2208));
    layer6_outputs(2172) <= (layer5_outputs(624)) xor (layer5_outputs(2230));
    layer6_outputs(2173) <= not((layer5_outputs(405)) and (layer5_outputs(677)));
    layer6_outputs(2174) <= not((layer5_outputs(2395)) or (layer5_outputs(1055)));
    layer6_outputs(2175) <= layer5_outputs(1229);
    layer6_outputs(2176) <= layer5_outputs(751);
    layer6_outputs(2177) <= layer5_outputs(2066);
    layer6_outputs(2178) <= not(layer5_outputs(1707));
    layer6_outputs(2179) <= not(layer5_outputs(747));
    layer6_outputs(2180) <= (layer5_outputs(755)) and (layer5_outputs(1886));
    layer6_outputs(2181) <= (layer5_outputs(2417)) and not (layer5_outputs(1254));
    layer6_outputs(2182) <= layer5_outputs(154);
    layer6_outputs(2183) <= not(layer5_outputs(1361));
    layer6_outputs(2184) <= not(layer5_outputs(2167));
    layer6_outputs(2185) <= not(layer5_outputs(928));
    layer6_outputs(2186) <= not(layer5_outputs(1883));
    layer6_outputs(2187) <= (layer5_outputs(1650)) and not (layer5_outputs(1601));
    layer6_outputs(2188) <= layer5_outputs(361);
    layer6_outputs(2189) <= layer5_outputs(761);
    layer6_outputs(2190) <= not(layer5_outputs(295));
    layer6_outputs(2191) <= not(layer5_outputs(921)) or (layer5_outputs(1306));
    layer6_outputs(2192) <= (layer5_outputs(1586)) and (layer5_outputs(1229));
    layer6_outputs(2193) <= not((layer5_outputs(389)) and (layer5_outputs(407)));
    layer6_outputs(2194) <= (layer5_outputs(13)) xor (layer5_outputs(2223));
    layer6_outputs(2195) <= (layer5_outputs(2249)) or (layer5_outputs(1933));
    layer6_outputs(2196) <= not(layer5_outputs(2051));
    layer6_outputs(2197) <= layer5_outputs(1816);
    layer6_outputs(2198) <= layer5_outputs(448);
    layer6_outputs(2199) <= layer5_outputs(2425);
    layer6_outputs(2200) <= layer5_outputs(891);
    layer6_outputs(2201) <= (layer5_outputs(1979)) or (layer5_outputs(613));
    layer6_outputs(2202) <= not((layer5_outputs(2456)) and (layer5_outputs(928)));
    layer6_outputs(2203) <= (layer5_outputs(2384)) and (layer5_outputs(2150));
    layer6_outputs(2204) <= layer5_outputs(1290);
    layer6_outputs(2205) <= not((layer5_outputs(1936)) xor (layer5_outputs(1783)));
    layer6_outputs(2206) <= not((layer5_outputs(611)) or (layer5_outputs(1441)));
    layer6_outputs(2207) <= not(layer5_outputs(2053));
    layer6_outputs(2208) <= (layer5_outputs(1104)) or (layer5_outputs(679));
    layer6_outputs(2209) <= not(layer5_outputs(2503));
    layer6_outputs(2210) <= not((layer5_outputs(1251)) or (layer5_outputs(780)));
    layer6_outputs(2211) <= layer5_outputs(1221);
    layer6_outputs(2212) <= '0';
    layer6_outputs(2213) <= layer5_outputs(90);
    layer6_outputs(2214) <= layer5_outputs(841);
    layer6_outputs(2215) <= not(layer5_outputs(135));
    layer6_outputs(2216) <= not((layer5_outputs(1922)) xor (layer5_outputs(1793)));
    layer6_outputs(2217) <= layer5_outputs(111);
    layer6_outputs(2218) <= layer5_outputs(2282);
    layer6_outputs(2219) <= (layer5_outputs(2490)) xor (layer5_outputs(54));
    layer6_outputs(2220) <= not(layer5_outputs(1589)) or (layer5_outputs(2535));
    layer6_outputs(2221) <= layer5_outputs(1413);
    layer6_outputs(2222) <= not(layer5_outputs(279));
    layer6_outputs(2223) <= layer5_outputs(2527);
    layer6_outputs(2224) <= layer5_outputs(1169);
    layer6_outputs(2225) <= (layer5_outputs(556)) xor (layer5_outputs(1123));
    layer6_outputs(2226) <= layer5_outputs(633);
    layer6_outputs(2227) <= layer5_outputs(1858);
    layer6_outputs(2228) <= layer5_outputs(254);
    layer6_outputs(2229) <= not((layer5_outputs(2259)) xor (layer5_outputs(1697)));
    layer6_outputs(2230) <= not(layer5_outputs(1259));
    layer6_outputs(2231) <= not(layer5_outputs(405));
    layer6_outputs(2232) <= not(layer5_outputs(91));
    layer6_outputs(2233) <= not(layer5_outputs(612));
    layer6_outputs(2234) <= not((layer5_outputs(31)) xor (layer5_outputs(2410)));
    layer6_outputs(2235) <= layer5_outputs(1800);
    layer6_outputs(2236) <= (layer5_outputs(1835)) or (layer5_outputs(997));
    layer6_outputs(2237) <= not(layer5_outputs(523));
    layer6_outputs(2238) <= layer5_outputs(1464);
    layer6_outputs(2239) <= (layer5_outputs(474)) xor (layer5_outputs(22));
    layer6_outputs(2240) <= layer5_outputs(2473);
    layer6_outputs(2241) <= not(layer5_outputs(940));
    layer6_outputs(2242) <= (layer5_outputs(1187)) and not (layer5_outputs(838));
    layer6_outputs(2243) <= layer5_outputs(1204);
    layer6_outputs(2244) <= not(layer5_outputs(982)) or (layer5_outputs(1735));
    layer6_outputs(2245) <= not((layer5_outputs(2465)) and (layer5_outputs(1811)));
    layer6_outputs(2246) <= not(layer5_outputs(1541));
    layer6_outputs(2247) <= layer5_outputs(2107);
    layer6_outputs(2248) <= layer5_outputs(2324);
    layer6_outputs(2249) <= not((layer5_outputs(2510)) xor (layer5_outputs(1786)));
    layer6_outputs(2250) <= not((layer5_outputs(802)) xor (layer5_outputs(1206)));
    layer6_outputs(2251) <= not((layer5_outputs(469)) xor (layer5_outputs(511)));
    layer6_outputs(2252) <= layer5_outputs(327);
    layer6_outputs(2253) <= (layer5_outputs(1859)) xor (layer5_outputs(538));
    layer6_outputs(2254) <= layer5_outputs(1065);
    layer6_outputs(2255) <= '1';
    layer6_outputs(2256) <= not(layer5_outputs(852));
    layer6_outputs(2257) <= not((layer5_outputs(2151)) xor (layer5_outputs(104)));
    layer6_outputs(2258) <= (layer5_outputs(1658)) xor (layer5_outputs(535));
    layer6_outputs(2259) <= layer5_outputs(651);
    layer6_outputs(2260) <= not((layer5_outputs(570)) and (layer5_outputs(1194)));
    layer6_outputs(2261) <= not(layer5_outputs(1255));
    layer6_outputs(2262) <= not(layer5_outputs(1435));
    layer6_outputs(2263) <= not(layer5_outputs(1435));
    layer6_outputs(2264) <= not(layer5_outputs(185));
    layer6_outputs(2265) <= (layer5_outputs(1568)) and not (layer5_outputs(1693));
    layer6_outputs(2266) <= (layer5_outputs(1098)) and not (layer5_outputs(1704));
    layer6_outputs(2267) <= not((layer5_outputs(2464)) xor (layer5_outputs(2119)));
    layer6_outputs(2268) <= not(layer5_outputs(1921));
    layer6_outputs(2269) <= not((layer5_outputs(2459)) and (layer5_outputs(1022)));
    layer6_outputs(2270) <= '1';
    layer6_outputs(2271) <= not(layer5_outputs(699)) or (layer5_outputs(1389));
    layer6_outputs(2272) <= not(layer5_outputs(440)) or (layer5_outputs(1523));
    layer6_outputs(2273) <= not(layer5_outputs(1844));
    layer6_outputs(2274) <= layer5_outputs(381);
    layer6_outputs(2275) <= not(layer5_outputs(1439));
    layer6_outputs(2276) <= not(layer5_outputs(969));
    layer6_outputs(2277) <= layer5_outputs(1849);
    layer6_outputs(2278) <= layer5_outputs(20);
    layer6_outputs(2279) <= layer5_outputs(118);
    layer6_outputs(2280) <= layer5_outputs(1360);
    layer6_outputs(2281) <= not(layer5_outputs(2190));
    layer6_outputs(2282) <= not((layer5_outputs(1912)) and (layer5_outputs(2060)));
    layer6_outputs(2283) <= not(layer5_outputs(2030));
    layer6_outputs(2284) <= not(layer5_outputs(913)) or (layer5_outputs(267));
    layer6_outputs(2285) <= layer5_outputs(582);
    layer6_outputs(2286) <= not(layer5_outputs(1788));
    layer6_outputs(2287) <= layer5_outputs(660);
    layer6_outputs(2288) <= not((layer5_outputs(2244)) or (layer5_outputs(1466)));
    layer6_outputs(2289) <= not(layer5_outputs(2171));
    layer6_outputs(2290) <= layer5_outputs(86);
    layer6_outputs(2291) <= layer5_outputs(472);
    layer6_outputs(2292) <= not(layer5_outputs(643));
    layer6_outputs(2293) <= not(layer5_outputs(2413));
    layer6_outputs(2294) <= not(layer5_outputs(1454));
    layer6_outputs(2295) <= not(layer5_outputs(935));
    layer6_outputs(2296) <= not(layer5_outputs(2141));
    layer6_outputs(2297) <= not((layer5_outputs(51)) xor (layer5_outputs(2207)));
    layer6_outputs(2298) <= layer5_outputs(2047);
    layer6_outputs(2299) <= not((layer5_outputs(1450)) and (layer5_outputs(1432)));
    layer6_outputs(2300) <= not(layer5_outputs(1934));
    layer6_outputs(2301) <= not(layer5_outputs(108)) or (layer5_outputs(1377));
    layer6_outputs(2302) <= layer5_outputs(247);
    layer6_outputs(2303) <= not(layer5_outputs(1715)) or (layer5_outputs(477));
    layer6_outputs(2304) <= not(layer5_outputs(2391));
    layer6_outputs(2305) <= layer5_outputs(302);
    layer6_outputs(2306) <= layer5_outputs(1118);
    layer6_outputs(2307) <= not((layer5_outputs(767)) and (layer5_outputs(701)));
    layer6_outputs(2308) <= layer5_outputs(728);
    layer6_outputs(2309) <= not(layer5_outputs(459));
    layer6_outputs(2310) <= not(layer5_outputs(342));
    layer6_outputs(2311) <= not(layer5_outputs(1580));
    layer6_outputs(2312) <= not(layer5_outputs(1969));
    layer6_outputs(2313) <= layer5_outputs(1610);
    layer6_outputs(2314) <= not(layer5_outputs(1970));
    layer6_outputs(2315) <= layer5_outputs(1596);
    layer6_outputs(2316) <= (layer5_outputs(1915)) xor (layer5_outputs(351));
    layer6_outputs(2317) <= (layer5_outputs(876)) or (layer5_outputs(1228));
    layer6_outputs(2318) <= not(layer5_outputs(533));
    layer6_outputs(2319) <= '0';
    layer6_outputs(2320) <= not(layer5_outputs(1023)) or (layer5_outputs(1246));
    layer6_outputs(2321) <= layer5_outputs(2163);
    layer6_outputs(2322) <= not(layer5_outputs(1699));
    layer6_outputs(2323) <= (layer5_outputs(470)) or (layer5_outputs(374));
    layer6_outputs(2324) <= not((layer5_outputs(685)) and (layer5_outputs(1838)));
    layer6_outputs(2325) <= layer5_outputs(174);
    layer6_outputs(2326) <= not((layer5_outputs(1938)) and (layer5_outputs(2046)));
    layer6_outputs(2327) <= not(layer5_outputs(2467));
    layer6_outputs(2328) <= not(layer5_outputs(1842));
    layer6_outputs(2329) <= layer5_outputs(2069);
    layer6_outputs(2330) <= layer5_outputs(1657);
    layer6_outputs(2331) <= not((layer5_outputs(1048)) xor (layer5_outputs(798)));
    layer6_outputs(2332) <= not((layer5_outputs(746)) xor (layer5_outputs(2421)));
    layer6_outputs(2333) <= layer5_outputs(413);
    layer6_outputs(2334) <= not(layer5_outputs(650));
    layer6_outputs(2335) <= not(layer5_outputs(1171)) or (layer5_outputs(2176));
    layer6_outputs(2336) <= layer5_outputs(1403);
    layer6_outputs(2337) <= not((layer5_outputs(2549)) or (layer5_outputs(218)));
    layer6_outputs(2338) <= layer5_outputs(1646);
    layer6_outputs(2339) <= not(layer5_outputs(198));
    layer6_outputs(2340) <= not(layer5_outputs(723));
    layer6_outputs(2341) <= layer5_outputs(2313);
    layer6_outputs(2342) <= not(layer5_outputs(1250));
    layer6_outputs(2343) <= layer5_outputs(2013);
    layer6_outputs(2344) <= not((layer5_outputs(2352)) xor (layer5_outputs(258)));
    layer6_outputs(2345) <= not(layer5_outputs(384));
    layer6_outputs(2346) <= not(layer5_outputs(1474));
    layer6_outputs(2347) <= not(layer5_outputs(2079));
    layer6_outputs(2348) <= layer5_outputs(229);
    layer6_outputs(2349) <= layer5_outputs(2144);
    layer6_outputs(2350) <= not((layer5_outputs(175)) xor (layer5_outputs(2479)));
    layer6_outputs(2351) <= layer5_outputs(1022);
    layer6_outputs(2352) <= (layer5_outputs(2345)) xor (layer5_outputs(805));
    layer6_outputs(2353) <= layer5_outputs(1066);
    layer6_outputs(2354) <= (layer5_outputs(2219)) and not (layer5_outputs(1797));
    layer6_outputs(2355) <= not((layer5_outputs(1092)) xor (layer5_outputs(518)));
    layer6_outputs(2356) <= (layer5_outputs(339)) and not (layer5_outputs(854));
    layer6_outputs(2357) <= (layer5_outputs(808)) and not (layer5_outputs(937));
    layer6_outputs(2358) <= not(layer5_outputs(1802));
    layer6_outputs(2359) <= (layer5_outputs(2489)) and (layer5_outputs(1461));
    layer6_outputs(2360) <= layer5_outputs(1257);
    layer6_outputs(2361) <= layer5_outputs(1791);
    layer6_outputs(2362) <= (layer5_outputs(2226)) or (layer5_outputs(844));
    layer6_outputs(2363) <= not((layer5_outputs(1421)) and (layer5_outputs(811)));
    layer6_outputs(2364) <= layer5_outputs(1394);
    layer6_outputs(2365) <= not(layer5_outputs(1467));
    layer6_outputs(2366) <= layer5_outputs(573);
    layer6_outputs(2367) <= layer5_outputs(510);
    layer6_outputs(2368) <= not(layer5_outputs(1813));
    layer6_outputs(2369) <= layer5_outputs(1423);
    layer6_outputs(2370) <= (layer5_outputs(1967)) and not (layer5_outputs(653));
    layer6_outputs(2371) <= not((layer5_outputs(1974)) or (layer5_outputs(1054)));
    layer6_outputs(2372) <= not(layer5_outputs(1555)) or (layer5_outputs(535));
    layer6_outputs(2373) <= not(layer5_outputs(692));
    layer6_outputs(2374) <= layer5_outputs(1771);
    layer6_outputs(2375) <= (layer5_outputs(1545)) or (layer5_outputs(582));
    layer6_outputs(2376) <= (layer5_outputs(50)) and not (layer5_outputs(1520));
    layer6_outputs(2377) <= not(layer5_outputs(1760));
    layer6_outputs(2378) <= layer5_outputs(2414);
    layer6_outputs(2379) <= not(layer5_outputs(419));
    layer6_outputs(2380) <= (layer5_outputs(645)) xor (layer5_outputs(337));
    layer6_outputs(2381) <= not(layer5_outputs(883));
    layer6_outputs(2382) <= not(layer5_outputs(254));
    layer6_outputs(2383) <= layer5_outputs(2385);
    layer6_outputs(2384) <= (layer5_outputs(2161)) and (layer5_outputs(1896));
    layer6_outputs(2385) <= layer5_outputs(379);
    layer6_outputs(2386) <= not(layer5_outputs(1479));
    layer6_outputs(2387) <= not((layer5_outputs(1412)) and (layer5_outputs(2142)));
    layer6_outputs(2388) <= not(layer5_outputs(543));
    layer6_outputs(2389) <= not((layer5_outputs(65)) xor (layer5_outputs(1330)));
    layer6_outputs(2390) <= (layer5_outputs(1996)) or (layer5_outputs(2538));
    layer6_outputs(2391) <= not(layer5_outputs(75));
    layer6_outputs(2392) <= not(layer5_outputs(1042));
    layer6_outputs(2393) <= not(layer5_outputs(2524)) or (layer5_outputs(1850));
    layer6_outputs(2394) <= (layer5_outputs(172)) or (layer5_outputs(1926));
    layer6_outputs(2395) <= '1';
    layer6_outputs(2396) <= layer5_outputs(1500);
    layer6_outputs(2397) <= (layer5_outputs(329)) and not (layer5_outputs(2179));
    layer6_outputs(2398) <= not((layer5_outputs(2023)) and (layer5_outputs(1547)));
    layer6_outputs(2399) <= not((layer5_outputs(1962)) and (layer5_outputs(1785)));
    layer6_outputs(2400) <= not(layer5_outputs(1097));
    layer6_outputs(2401) <= (layer5_outputs(2400)) or (layer5_outputs(1584));
    layer6_outputs(2402) <= not(layer5_outputs(178));
    layer6_outputs(2403) <= layer5_outputs(32);
    layer6_outputs(2404) <= (layer5_outputs(1577)) and not (layer5_outputs(354));
    layer6_outputs(2405) <= not(layer5_outputs(1277));
    layer6_outputs(2406) <= not((layer5_outputs(2533)) xor (layer5_outputs(225)));
    layer6_outputs(2407) <= '0';
    layer6_outputs(2408) <= not(layer5_outputs(1914));
    layer6_outputs(2409) <= (layer5_outputs(338)) xor (layer5_outputs(481));
    layer6_outputs(2410) <= not((layer5_outputs(2015)) xor (layer5_outputs(1195)));
    layer6_outputs(2411) <= not(layer5_outputs(1185)) or (layer5_outputs(1378));
    layer6_outputs(2412) <= (layer5_outputs(1264)) and not (layer5_outputs(631));
    layer6_outputs(2413) <= not(layer5_outputs(2270));
    layer6_outputs(2414) <= (layer5_outputs(285)) and not (layer5_outputs(2082));
    layer6_outputs(2415) <= not(layer5_outputs(687));
    layer6_outputs(2416) <= (layer5_outputs(463)) xor (layer5_outputs(1069));
    layer6_outputs(2417) <= layer5_outputs(1310);
    layer6_outputs(2418) <= not(layer5_outputs(1011));
    layer6_outputs(2419) <= not(layer5_outputs(87)) or (layer5_outputs(1917));
    layer6_outputs(2420) <= not(layer5_outputs(1291));
    layer6_outputs(2421) <= not(layer5_outputs(193));
    layer6_outputs(2422) <= layer5_outputs(1845);
    layer6_outputs(2423) <= not((layer5_outputs(2214)) and (layer5_outputs(1434)));
    layer6_outputs(2424) <= (layer5_outputs(2362)) and not (layer5_outputs(274));
    layer6_outputs(2425) <= not(layer5_outputs(169));
    layer6_outputs(2426) <= not(layer5_outputs(1427));
    layer6_outputs(2427) <= not(layer5_outputs(857));
    layer6_outputs(2428) <= layer5_outputs(1197);
    layer6_outputs(2429) <= layer5_outputs(1107);
    layer6_outputs(2430) <= layer5_outputs(1508);
    layer6_outputs(2431) <= not(layer5_outputs(1288));
    layer6_outputs(2432) <= not(layer5_outputs(1033));
    layer6_outputs(2433) <= layer5_outputs(2007);
    layer6_outputs(2434) <= not((layer5_outputs(2291)) xor (layer5_outputs(993)));
    layer6_outputs(2435) <= not((layer5_outputs(1053)) xor (layer5_outputs(577)));
    layer6_outputs(2436) <= layer5_outputs(281);
    layer6_outputs(2437) <= not(layer5_outputs(1344));
    layer6_outputs(2438) <= not(layer5_outputs(462));
    layer6_outputs(2439) <= (layer5_outputs(1645)) and (layer5_outputs(446));
    layer6_outputs(2440) <= (layer5_outputs(2070)) and not (layer5_outputs(1497));
    layer6_outputs(2441) <= not((layer5_outputs(1128)) or (layer5_outputs(2192)));
    layer6_outputs(2442) <= layer5_outputs(1051);
    layer6_outputs(2443) <= '0';
    layer6_outputs(2444) <= '0';
    layer6_outputs(2445) <= not(layer5_outputs(97));
    layer6_outputs(2446) <= (layer5_outputs(366)) xor (layer5_outputs(832));
    layer6_outputs(2447) <= not(layer5_outputs(1706));
    layer6_outputs(2448) <= not((layer5_outputs(2112)) xor (layer5_outputs(2321)));
    layer6_outputs(2449) <= not(layer5_outputs(677));
    layer6_outputs(2450) <= (layer5_outputs(2139)) xor (layer5_outputs(1987));
    layer6_outputs(2451) <= not(layer5_outputs(1534));
    layer6_outputs(2452) <= not(layer5_outputs(539));
    layer6_outputs(2453) <= (layer5_outputs(923)) xor (layer5_outputs(1213));
    layer6_outputs(2454) <= not(layer5_outputs(1506));
    layer6_outputs(2455) <= not(layer5_outputs(1678)) or (layer5_outputs(2203));
    layer6_outputs(2456) <= (layer5_outputs(1374)) and not (layer5_outputs(1198));
    layer6_outputs(2457) <= (layer5_outputs(305)) xor (layer5_outputs(1092));
    layer6_outputs(2458) <= not(layer5_outputs(2004));
    layer6_outputs(2459) <= not(layer5_outputs(1509));
    layer6_outputs(2460) <= layer5_outputs(2267);
    layer6_outputs(2461) <= not(layer5_outputs(101));
    layer6_outputs(2462) <= layer5_outputs(52);
    layer6_outputs(2463) <= (layer5_outputs(991)) xor (layer5_outputs(2270));
    layer6_outputs(2464) <= not(layer5_outputs(548));
    layer6_outputs(2465) <= layer5_outputs(336);
    layer6_outputs(2466) <= (layer5_outputs(447)) and not (layer5_outputs(810));
    layer6_outputs(2467) <= not(layer5_outputs(990)) or (layer5_outputs(1133));
    layer6_outputs(2468) <= layer5_outputs(7);
    layer6_outputs(2469) <= not(layer5_outputs(1417));
    layer6_outputs(2470) <= not(layer5_outputs(1400)) or (layer5_outputs(2491));
    layer6_outputs(2471) <= not(layer5_outputs(2556)) or (layer5_outputs(1740));
    layer6_outputs(2472) <= not(layer5_outputs(2526));
    layer6_outputs(2473) <= not(layer5_outputs(1860)) or (layer5_outputs(1698));
    layer6_outputs(2474) <= layer5_outputs(1683);
    layer6_outputs(2475) <= layer5_outputs(83);
    layer6_outputs(2476) <= layer5_outputs(160);
    layer6_outputs(2477) <= (layer5_outputs(96)) and not (layer5_outputs(47));
    layer6_outputs(2478) <= layer5_outputs(1700);
    layer6_outputs(2479) <= not(layer5_outputs(1536));
    layer6_outputs(2480) <= layer5_outputs(896);
    layer6_outputs(2481) <= not((layer5_outputs(183)) xor (layer5_outputs(132)));
    layer6_outputs(2482) <= layer5_outputs(2148);
    layer6_outputs(2483) <= layer5_outputs(867);
    layer6_outputs(2484) <= not(layer5_outputs(210)) or (layer5_outputs(1750));
    layer6_outputs(2485) <= not(layer5_outputs(422));
    layer6_outputs(2486) <= not(layer5_outputs(1908));
    layer6_outputs(2487) <= layer5_outputs(2358);
    layer6_outputs(2488) <= not(layer5_outputs(1782)) or (layer5_outputs(2254));
    layer6_outputs(2489) <= layer5_outputs(1634);
    layer6_outputs(2490) <= not(layer5_outputs(2060));
    layer6_outputs(2491) <= not((layer5_outputs(1784)) and (layer5_outputs(1676)));
    layer6_outputs(2492) <= '0';
    layer6_outputs(2493) <= not(layer5_outputs(938));
    layer6_outputs(2494) <= layer5_outputs(1809);
    layer6_outputs(2495) <= not(layer5_outputs(2165));
    layer6_outputs(2496) <= layer5_outputs(965);
    layer6_outputs(2497) <= (layer5_outputs(1304)) and not (layer5_outputs(1245));
    layer6_outputs(2498) <= (layer5_outputs(1163)) or (layer5_outputs(2347));
    layer6_outputs(2499) <= (layer5_outputs(256)) and (layer5_outputs(1869));
    layer6_outputs(2500) <= not(layer5_outputs(2528));
    layer6_outputs(2501) <= not(layer5_outputs(692));
    layer6_outputs(2502) <= layer5_outputs(1980);
    layer6_outputs(2503) <= (layer5_outputs(1822)) and not (layer5_outputs(878));
    layer6_outputs(2504) <= not(layer5_outputs(2504));
    layer6_outputs(2505) <= not(layer5_outputs(1494));
    layer6_outputs(2506) <= (layer5_outputs(2416)) and not (layer5_outputs(1051));
    layer6_outputs(2507) <= layer5_outputs(1111);
    layer6_outputs(2508) <= not(layer5_outputs(454));
    layer6_outputs(2509) <= layer5_outputs(2481);
    layer6_outputs(2510) <= not(layer5_outputs(2216)) or (layer5_outputs(2171));
    layer6_outputs(2511) <= not((layer5_outputs(1756)) and (layer5_outputs(2532)));
    layer6_outputs(2512) <= (layer5_outputs(1382)) xor (layer5_outputs(1683));
    layer6_outputs(2513) <= not(layer5_outputs(1700));
    layer6_outputs(2514) <= layer5_outputs(439);
    layer6_outputs(2515) <= '0';
    layer6_outputs(2516) <= not(layer5_outputs(1653)) or (layer5_outputs(48));
    layer6_outputs(2517) <= not((layer5_outputs(1391)) and (layer5_outputs(387)));
    layer6_outputs(2518) <= (layer5_outputs(391)) and (layer5_outputs(378));
    layer6_outputs(2519) <= (layer5_outputs(1479)) and not (layer5_outputs(1238));
    layer6_outputs(2520) <= not((layer5_outputs(632)) and (layer5_outputs(1527)));
    layer6_outputs(2521) <= not((layer5_outputs(2043)) and (layer5_outputs(2072)));
    layer6_outputs(2522) <= not((layer5_outputs(1208)) and (layer5_outputs(2262)));
    layer6_outputs(2523) <= not(layer5_outputs(2126));
    layer6_outputs(2524) <= not(layer5_outputs(1043)) or (layer5_outputs(2162));
    layer6_outputs(2525) <= not(layer5_outputs(1831));
    layer6_outputs(2526) <= not(layer5_outputs(502));
    layer6_outputs(2527) <= '0';
    layer6_outputs(2528) <= not((layer5_outputs(526)) xor (layer5_outputs(2555)));
    layer6_outputs(2529) <= (layer5_outputs(2)) and not (layer5_outputs(1160));
    layer6_outputs(2530) <= (layer5_outputs(489)) xor (layer5_outputs(73));
    layer6_outputs(2531) <= layer5_outputs(2516);
    layer6_outputs(2532) <= not(layer5_outputs(967)) or (layer5_outputs(245));
    layer6_outputs(2533) <= not(layer5_outputs(1146)) or (layer5_outputs(931));
    layer6_outputs(2534) <= layer5_outputs(1338);
    layer6_outputs(2535) <= layer5_outputs(1352);
    layer6_outputs(2536) <= (layer5_outputs(1733)) xor (layer5_outputs(261));
    layer6_outputs(2537) <= not(layer5_outputs(1149));
    layer6_outputs(2538) <= (layer5_outputs(1756)) and not (layer5_outputs(2466));
    layer6_outputs(2539) <= not((layer5_outputs(1888)) and (layer5_outputs(575)));
    layer6_outputs(2540) <= layer5_outputs(2242);
    layer6_outputs(2541) <= layer5_outputs(1933);
    layer6_outputs(2542) <= not(layer5_outputs(1340)) or (layer5_outputs(1227));
    layer6_outputs(2543) <= layer5_outputs(1744);
    layer6_outputs(2544) <= not(layer5_outputs(168));
    layer6_outputs(2545) <= (layer5_outputs(346)) and not (layer5_outputs(2224));
    layer6_outputs(2546) <= not((layer5_outputs(1964)) xor (layer5_outputs(2012)));
    layer6_outputs(2547) <= (layer5_outputs(1859)) xor (layer5_outputs(1246));
    layer6_outputs(2548) <= not((layer5_outputs(1629)) xor (layer5_outputs(856)));
    layer6_outputs(2549) <= not(layer5_outputs(1935));
    layer6_outputs(2550) <= not(layer5_outputs(1173));
    layer6_outputs(2551) <= layer5_outputs(138);
    layer6_outputs(2552) <= not(layer5_outputs(271));
    layer6_outputs(2553) <= (layer5_outputs(2307)) and (layer5_outputs(426));
    layer6_outputs(2554) <= not((layer5_outputs(1592)) and (layer5_outputs(2493)));
    layer6_outputs(2555) <= not(layer5_outputs(1005)) or (layer5_outputs(642));
    layer6_outputs(2556) <= not(layer5_outputs(1739));
    layer6_outputs(2557) <= not((layer5_outputs(1576)) xor (layer5_outputs(926)));
    layer6_outputs(2558) <= (layer5_outputs(438)) or (layer5_outputs(430));
    layer6_outputs(2559) <= not(layer5_outputs(2029)) or (layer5_outputs(1553));
    outputs(0) <= (layer6_outputs(749)) xor (layer6_outputs(1991));
    outputs(1) <= layer6_outputs(1492);
    outputs(2) <= not(layer6_outputs(1913));
    outputs(3) <= layer6_outputs(2304);
    outputs(4) <= not(layer6_outputs(1648));
    outputs(5) <= not(layer6_outputs(186));
    outputs(6) <= layer6_outputs(962);
    outputs(7) <= layer6_outputs(841);
    outputs(8) <= layer6_outputs(1034);
    outputs(9) <= layer6_outputs(523);
    outputs(10) <= layer6_outputs(1561);
    outputs(11) <= (layer6_outputs(1660)) xor (layer6_outputs(939));
    outputs(12) <= layer6_outputs(763);
    outputs(13) <= not((layer6_outputs(1993)) or (layer6_outputs(1939)));
    outputs(14) <= layer6_outputs(1457);
    outputs(15) <= layer6_outputs(2356);
    outputs(16) <= not(layer6_outputs(518));
    outputs(17) <= layer6_outputs(2208);
    outputs(18) <= layer6_outputs(2232);
    outputs(19) <= layer6_outputs(1237);
    outputs(20) <= not((layer6_outputs(367)) xor (layer6_outputs(376)));
    outputs(21) <= not(layer6_outputs(1432));
    outputs(22) <= layer6_outputs(1625);
    outputs(23) <= layer6_outputs(1065);
    outputs(24) <= not((layer6_outputs(283)) and (layer6_outputs(1410)));
    outputs(25) <= not(layer6_outputs(1573));
    outputs(26) <= not(layer6_outputs(838));
    outputs(27) <= not(layer6_outputs(621));
    outputs(28) <= layer6_outputs(847);
    outputs(29) <= not(layer6_outputs(984));
    outputs(30) <= layer6_outputs(654);
    outputs(31) <= layer6_outputs(1150);
    outputs(32) <= not(layer6_outputs(733));
    outputs(33) <= not(layer6_outputs(1409));
    outputs(34) <= not(layer6_outputs(2540));
    outputs(35) <= not((layer6_outputs(776)) xor (layer6_outputs(2072)));
    outputs(36) <= not(layer6_outputs(1616));
    outputs(37) <= layer6_outputs(1699);
    outputs(38) <= layer6_outputs(1492);
    outputs(39) <= (layer6_outputs(1036)) and not (layer6_outputs(2442));
    outputs(40) <= not(layer6_outputs(100));
    outputs(41) <= not(layer6_outputs(235));
    outputs(42) <= layer6_outputs(2377);
    outputs(43) <= layer6_outputs(2462);
    outputs(44) <= not(layer6_outputs(1731));
    outputs(45) <= not(layer6_outputs(2393));
    outputs(46) <= layer6_outputs(662);
    outputs(47) <= not(layer6_outputs(1210));
    outputs(48) <= not(layer6_outputs(2292));
    outputs(49) <= layer6_outputs(758);
    outputs(50) <= not((layer6_outputs(1908)) xor (layer6_outputs(1750)));
    outputs(51) <= (layer6_outputs(265)) and (layer6_outputs(1825));
    outputs(52) <= not(layer6_outputs(2317));
    outputs(53) <= (layer6_outputs(526)) xor (layer6_outputs(1031));
    outputs(54) <= layer6_outputs(2063);
    outputs(55) <= not(layer6_outputs(255));
    outputs(56) <= (layer6_outputs(1597)) and not (layer6_outputs(2300));
    outputs(57) <= not(layer6_outputs(335));
    outputs(58) <= not((layer6_outputs(1361)) or (layer6_outputs(2176)));
    outputs(59) <= not(layer6_outputs(65));
    outputs(60) <= not(layer6_outputs(774));
    outputs(61) <= layer6_outputs(660);
    outputs(62) <= not(layer6_outputs(605));
    outputs(63) <= layer6_outputs(1661);
    outputs(64) <= (layer6_outputs(828)) xor (layer6_outputs(136));
    outputs(65) <= not((layer6_outputs(1286)) and (layer6_outputs(1993)));
    outputs(66) <= layer6_outputs(41);
    outputs(67) <= layer6_outputs(452);
    outputs(68) <= layer6_outputs(284);
    outputs(69) <= not((layer6_outputs(1526)) xor (layer6_outputs(1005)));
    outputs(70) <= layer6_outputs(1852);
    outputs(71) <= not(layer6_outputs(974));
    outputs(72) <= (layer6_outputs(1953)) and (layer6_outputs(312));
    outputs(73) <= layer6_outputs(1466);
    outputs(74) <= layer6_outputs(1207);
    outputs(75) <= not(layer6_outputs(1165));
    outputs(76) <= (layer6_outputs(1489)) and (layer6_outputs(1936));
    outputs(77) <= layer6_outputs(1372);
    outputs(78) <= not(layer6_outputs(995));
    outputs(79) <= not(layer6_outputs(240));
    outputs(80) <= not(layer6_outputs(2337));
    outputs(81) <= layer6_outputs(823);
    outputs(82) <= layer6_outputs(523);
    outputs(83) <= not((layer6_outputs(65)) xor (layer6_outputs(902)));
    outputs(84) <= layer6_outputs(2187);
    outputs(85) <= not(layer6_outputs(549));
    outputs(86) <= layer6_outputs(1311);
    outputs(87) <= not(layer6_outputs(2163));
    outputs(88) <= not(layer6_outputs(1048));
    outputs(89) <= layer6_outputs(192);
    outputs(90) <= not(layer6_outputs(2446)) or (layer6_outputs(2301));
    outputs(91) <= not(layer6_outputs(2223));
    outputs(92) <= not(layer6_outputs(2362));
    outputs(93) <= not(layer6_outputs(498));
    outputs(94) <= layer6_outputs(868);
    outputs(95) <= (layer6_outputs(2235)) xor (layer6_outputs(1503));
    outputs(96) <= not(layer6_outputs(881));
    outputs(97) <= not(layer6_outputs(1373)) or (layer6_outputs(1095));
    outputs(98) <= not((layer6_outputs(2057)) or (layer6_outputs(1378)));
    outputs(99) <= (layer6_outputs(1903)) and not (layer6_outputs(1683));
    outputs(100) <= layer6_outputs(1180);
    outputs(101) <= layer6_outputs(1139);
    outputs(102) <= not(layer6_outputs(253));
    outputs(103) <= layer6_outputs(1534);
    outputs(104) <= layer6_outputs(1054);
    outputs(105) <= layer6_outputs(417);
    outputs(106) <= not(layer6_outputs(2456));
    outputs(107) <= (layer6_outputs(1591)) and not (layer6_outputs(881));
    outputs(108) <= not(layer6_outputs(1224));
    outputs(109) <= not((layer6_outputs(1761)) or (layer6_outputs(2174)));
    outputs(110) <= (layer6_outputs(1986)) or (layer6_outputs(1208));
    outputs(111) <= not(layer6_outputs(378));
    outputs(112) <= layer6_outputs(2543);
    outputs(113) <= layer6_outputs(1401);
    outputs(114) <= layer6_outputs(1931);
    outputs(115) <= layer6_outputs(1965);
    outputs(116) <= not(layer6_outputs(1234));
    outputs(117) <= not(layer6_outputs(371));
    outputs(118) <= not(layer6_outputs(1787));
    outputs(119) <= not(layer6_outputs(415));
    outputs(120) <= layer6_outputs(1292);
    outputs(121) <= (layer6_outputs(639)) and (layer6_outputs(197));
    outputs(122) <= not(layer6_outputs(2051));
    outputs(123) <= layer6_outputs(1695);
    outputs(124) <= not(layer6_outputs(638));
    outputs(125) <= layer6_outputs(1811);
    outputs(126) <= layer6_outputs(690);
    outputs(127) <= not(layer6_outputs(2039));
    outputs(128) <= not(layer6_outputs(2332));
    outputs(129) <= not(layer6_outputs(886));
    outputs(130) <= (layer6_outputs(642)) and not (layer6_outputs(25));
    outputs(131) <= not(layer6_outputs(1723));
    outputs(132) <= not((layer6_outputs(1220)) xor (layer6_outputs(659)));
    outputs(133) <= (layer6_outputs(1965)) xor (layer6_outputs(1713));
    outputs(134) <= not(layer6_outputs(273));
    outputs(135) <= layer6_outputs(1479);
    outputs(136) <= not(layer6_outputs(316));
    outputs(137) <= not(layer6_outputs(731));
    outputs(138) <= (layer6_outputs(1495)) or (layer6_outputs(1087));
    outputs(139) <= layer6_outputs(2041);
    outputs(140) <= not(layer6_outputs(283));
    outputs(141) <= (layer6_outputs(1057)) xor (layer6_outputs(859));
    outputs(142) <= layer6_outputs(1354);
    outputs(143) <= layer6_outputs(1796);
    outputs(144) <= not((layer6_outputs(1332)) or (layer6_outputs(1459)));
    outputs(145) <= layer6_outputs(2135);
    outputs(146) <= layer6_outputs(933);
    outputs(147) <= layer6_outputs(1104);
    outputs(148) <= not(layer6_outputs(2524)) or (layer6_outputs(1769));
    outputs(149) <= not(layer6_outputs(293));
    outputs(150) <= layer6_outputs(1433);
    outputs(151) <= layer6_outputs(160);
    outputs(152) <= layer6_outputs(587);
    outputs(153) <= layer6_outputs(993);
    outputs(154) <= layer6_outputs(1882);
    outputs(155) <= not(layer6_outputs(1440)) or (layer6_outputs(1549));
    outputs(156) <= layer6_outputs(658);
    outputs(157) <= not(layer6_outputs(2234));
    outputs(158) <= not((layer6_outputs(1691)) or (layer6_outputs(1595)));
    outputs(159) <= not(layer6_outputs(1911));
    outputs(160) <= not((layer6_outputs(1343)) xor (layer6_outputs(1970)));
    outputs(161) <= not(layer6_outputs(194));
    outputs(162) <= not(layer6_outputs(2445));
    outputs(163) <= (layer6_outputs(409)) and (layer6_outputs(68));
    outputs(164) <= layer6_outputs(519);
    outputs(165) <= (layer6_outputs(246)) or (layer6_outputs(973));
    outputs(166) <= not(layer6_outputs(1584));
    outputs(167) <= layer6_outputs(383);
    outputs(168) <= layer6_outputs(1012);
    outputs(169) <= not((layer6_outputs(178)) xor (layer6_outputs(1637)));
    outputs(170) <= not(layer6_outputs(817));
    outputs(171) <= not((layer6_outputs(1140)) xor (layer6_outputs(1963)));
    outputs(172) <= not(layer6_outputs(2485));
    outputs(173) <= not((layer6_outputs(903)) or (layer6_outputs(971)));
    outputs(174) <= layer6_outputs(1209);
    outputs(175) <= (layer6_outputs(2545)) or (layer6_outputs(2414));
    outputs(176) <= not(layer6_outputs(1730));
    outputs(177) <= not((layer6_outputs(2452)) or (layer6_outputs(2388)));
    outputs(178) <= not(layer6_outputs(2157));
    outputs(179) <= not(layer6_outputs(549));
    outputs(180) <= not(layer6_outputs(1849)) or (layer6_outputs(1737));
    outputs(181) <= not(layer6_outputs(2403));
    outputs(182) <= not(layer6_outputs(1268));
    outputs(183) <= (layer6_outputs(715)) and (layer6_outputs(514));
    outputs(184) <= (layer6_outputs(2158)) or (layer6_outputs(2349));
    outputs(185) <= not(layer6_outputs(44));
    outputs(186) <= not(layer6_outputs(2101));
    outputs(187) <= layer6_outputs(224);
    outputs(188) <= not((layer6_outputs(1628)) xor (layer6_outputs(2053)));
    outputs(189) <= not(layer6_outputs(1644));
    outputs(190) <= not((layer6_outputs(1531)) xor (layer6_outputs(1547)));
    outputs(191) <= not(layer6_outputs(1780));
    outputs(192) <= (layer6_outputs(515)) xor (layer6_outputs(2538));
    outputs(193) <= not(layer6_outputs(693));
    outputs(194) <= not(layer6_outputs(2333));
    outputs(195) <= not(layer6_outputs(1364));
    outputs(196) <= not((layer6_outputs(1269)) or (layer6_outputs(1320)));
    outputs(197) <= layer6_outputs(1187);
    outputs(198) <= not((layer6_outputs(442)) xor (layer6_outputs(1995)));
    outputs(199) <= (layer6_outputs(1343)) and not (layer6_outputs(1621));
    outputs(200) <= not(layer6_outputs(2360));
    outputs(201) <= not(layer6_outputs(1058));
    outputs(202) <= (layer6_outputs(2283)) and not (layer6_outputs(2475));
    outputs(203) <= layer6_outputs(2277);
    outputs(204) <= (layer6_outputs(2486)) and not (layer6_outputs(1230));
    outputs(205) <= layer6_outputs(1260);
    outputs(206) <= not(layer6_outputs(1172));
    outputs(207) <= (layer6_outputs(2383)) and not (layer6_outputs(240));
    outputs(208) <= (layer6_outputs(1280)) and not (layer6_outputs(1094));
    outputs(209) <= not(layer6_outputs(2421));
    outputs(210) <= not((layer6_outputs(2082)) xor (layer6_outputs(1645)));
    outputs(211) <= not(layer6_outputs(2009));
    outputs(212) <= not(layer6_outputs(2457));
    outputs(213) <= not((layer6_outputs(2394)) xor (layer6_outputs(204)));
    outputs(214) <= not(layer6_outputs(1287));
    outputs(215) <= not(layer6_outputs(1460));
    outputs(216) <= layer6_outputs(196);
    outputs(217) <= (layer6_outputs(153)) xor (layer6_outputs(1102));
    outputs(218) <= layer6_outputs(2291);
    outputs(219) <= not(layer6_outputs(54));
    outputs(220) <= not(layer6_outputs(1906));
    outputs(221) <= not((layer6_outputs(557)) or (layer6_outputs(1137)));
    outputs(222) <= not((layer6_outputs(258)) and (layer6_outputs(1558)));
    outputs(223) <= not(layer6_outputs(1589));
    outputs(224) <= not(layer6_outputs(1812));
    outputs(225) <= not(layer6_outputs(1024));
    outputs(226) <= layer6_outputs(1678);
    outputs(227) <= not(layer6_outputs(1774)) or (layer6_outputs(303));
    outputs(228) <= layer6_outputs(1590);
    outputs(229) <= not(layer6_outputs(2021));
    outputs(230) <= not(layer6_outputs(502));
    outputs(231) <= not(layer6_outputs(2231));
    outputs(232) <= not(layer6_outputs(698));
    outputs(233) <= layer6_outputs(422);
    outputs(234) <= not((layer6_outputs(1164)) and (layer6_outputs(222)));
    outputs(235) <= layer6_outputs(2115);
    outputs(236) <= not(layer6_outputs(863));
    outputs(237) <= not(layer6_outputs(1951));
    outputs(238) <= (layer6_outputs(1133)) and not (layer6_outputs(580));
    outputs(239) <= not(layer6_outputs(880));
    outputs(240) <= layer6_outputs(445);
    outputs(241) <= not(layer6_outputs(2022));
    outputs(242) <= (layer6_outputs(2368)) and not (layer6_outputs(1038));
    outputs(243) <= layer6_outputs(305);
    outputs(244) <= (layer6_outputs(1657)) xor (layer6_outputs(2155));
    outputs(245) <= not(layer6_outputs(261));
    outputs(246) <= (layer6_outputs(2221)) and not (layer6_outputs(77));
    outputs(247) <= not(layer6_outputs(1255));
    outputs(248) <= (layer6_outputs(230)) and not (layer6_outputs(2146));
    outputs(249) <= not(layer6_outputs(1302));
    outputs(250) <= layer6_outputs(2367);
    outputs(251) <= not(layer6_outputs(2198));
    outputs(252) <= (layer6_outputs(2327)) xor (layer6_outputs(2559));
    outputs(253) <= (layer6_outputs(708)) and not (layer6_outputs(1334));
    outputs(254) <= not((layer6_outputs(701)) xor (layer6_outputs(234)));
    outputs(255) <= layer6_outputs(689);
    outputs(256) <= not(layer6_outputs(1109));
    outputs(257) <= not(layer6_outputs(2298)) or (layer6_outputs(1439));
    outputs(258) <= not((layer6_outputs(1496)) xor (layer6_outputs(47)));
    outputs(259) <= (layer6_outputs(169)) and (layer6_outputs(359));
    outputs(260) <= layer6_outputs(2245);
    outputs(261) <= layer6_outputs(427);
    outputs(262) <= not(layer6_outputs(344));
    outputs(263) <= not(layer6_outputs(181));
    outputs(264) <= not(layer6_outputs(2230));
    outputs(265) <= layer6_outputs(93);
    outputs(266) <= not(layer6_outputs(1795));
    outputs(267) <= not(layer6_outputs(2213));
    outputs(268) <= layer6_outputs(1939);
    outputs(269) <= (layer6_outputs(88)) and not (layer6_outputs(1999));
    outputs(270) <= not((layer6_outputs(2120)) xor (layer6_outputs(2283)));
    outputs(271) <= not(layer6_outputs(1034));
    outputs(272) <= layer6_outputs(287);
    outputs(273) <= not(layer6_outputs(749));
    outputs(274) <= not(layer6_outputs(821));
    outputs(275) <= (layer6_outputs(1102)) and not (layer6_outputs(32));
    outputs(276) <= layer6_outputs(461);
    outputs(277) <= layer6_outputs(1528);
    outputs(278) <= not(layer6_outputs(1243));
    outputs(279) <= not(layer6_outputs(522));
    outputs(280) <= not(layer6_outputs(2367));
    outputs(281) <= (layer6_outputs(963)) and not (layer6_outputs(1737));
    outputs(282) <= not(layer6_outputs(1105));
    outputs(283) <= not(layer6_outputs(1468));
    outputs(284) <= (layer6_outputs(1498)) and not (layer6_outputs(757));
    outputs(285) <= layer6_outputs(1980);
    outputs(286) <= layer6_outputs(686);
    outputs(287) <= (layer6_outputs(954)) and (layer6_outputs(1329));
    outputs(288) <= not(layer6_outputs(422));
    outputs(289) <= not(layer6_outputs(206));
    outputs(290) <= (layer6_outputs(328)) and (layer6_outputs(1726));
    outputs(291) <= not((layer6_outputs(2434)) or (layer6_outputs(2058)));
    outputs(292) <= layer6_outputs(2171);
    outputs(293) <= layer6_outputs(1088);
    outputs(294) <= not(layer6_outputs(1899));
    outputs(295) <= (layer6_outputs(1879)) xor (layer6_outputs(2559));
    outputs(296) <= layer6_outputs(37);
    outputs(297) <= layer6_outputs(149);
    outputs(298) <= not((layer6_outputs(1679)) xor (layer6_outputs(2056)));
    outputs(299) <= (layer6_outputs(2033)) and not (layer6_outputs(40));
    outputs(300) <= not(layer6_outputs(1144));
    outputs(301) <= (layer6_outputs(411)) and not (layer6_outputs(339));
    outputs(302) <= layer6_outputs(2242);
    outputs(303) <= not(layer6_outputs(531));
    outputs(304) <= layer6_outputs(989);
    outputs(305) <= layer6_outputs(2145);
    outputs(306) <= not((layer6_outputs(2527)) or (layer6_outputs(1306)));
    outputs(307) <= layer6_outputs(176);
    outputs(308) <= layer6_outputs(1379);
    outputs(309) <= not((layer6_outputs(236)) xor (layer6_outputs(2320)));
    outputs(310) <= (layer6_outputs(713)) xor (layer6_outputs(877));
    outputs(311) <= not(layer6_outputs(1509));
    outputs(312) <= (layer6_outputs(1931)) and (layer6_outputs(631));
    outputs(313) <= not(layer6_outputs(1013));
    outputs(314) <= layer6_outputs(2095);
    outputs(315) <= layer6_outputs(2100);
    outputs(316) <= not((layer6_outputs(497)) xor (layer6_outputs(2236)));
    outputs(317) <= (layer6_outputs(182)) and not (layer6_outputs(760));
    outputs(318) <= (layer6_outputs(2364)) xor (layer6_outputs(1692));
    outputs(319) <= not((layer6_outputs(1047)) or (layer6_outputs(757)));
    outputs(320) <= not((layer6_outputs(1271)) xor (layer6_outputs(340)));
    outputs(321) <= not(layer6_outputs(1103));
    outputs(322) <= (layer6_outputs(891)) and not (layer6_outputs(117));
    outputs(323) <= not((layer6_outputs(248)) or (layer6_outputs(1718)));
    outputs(324) <= not(layer6_outputs(2004));
    outputs(325) <= layer6_outputs(77);
    outputs(326) <= layer6_outputs(334);
    outputs(327) <= (layer6_outputs(382)) and not (layer6_outputs(1782));
    outputs(328) <= (layer6_outputs(836)) and not (layer6_outputs(596));
    outputs(329) <= layer6_outputs(2396);
    outputs(330) <= not(layer6_outputs(1242));
    outputs(331) <= (layer6_outputs(561)) and (layer6_outputs(384));
    outputs(332) <= (layer6_outputs(173)) and (layer6_outputs(1572));
    outputs(333) <= layer6_outputs(2071);
    outputs(334) <= not((layer6_outputs(2364)) xor (layer6_outputs(2450)));
    outputs(335) <= not(layer6_outputs(765));
    outputs(336) <= (layer6_outputs(449)) and (layer6_outputs(2157));
    outputs(337) <= not(layer6_outputs(553));
    outputs(338) <= not((layer6_outputs(990)) xor (layer6_outputs(1207)));
    outputs(339) <= not((layer6_outputs(1990)) and (layer6_outputs(781)));
    outputs(340) <= not(layer6_outputs(747));
    outputs(341) <= not(layer6_outputs(1242));
    outputs(342) <= layer6_outputs(1194);
    outputs(343) <= not(layer6_outputs(2547));
    outputs(344) <= (layer6_outputs(509)) and not (layer6_outputs(1131));
    outputs(345) <= not((layer6_outputs(1882)) or (layer6_outputs(2019)));
    outputs(346) <= not(layer6_outputs(1532));
    outputs(347) <= (layer6_outputs(1266)) xor (layer6_outputs(2040));
    outputs(348) <= not((layer6_outputs(1788)) xor (layer6_outputs(1399)));
    outputs(349) <= (layer6_outputs(349)) and (layer6_outputs(302));
    outputs(350) <= layer6_outputs(456);
    outputs(351) <= not(layer6_outputs(1989));
    outputs(352) <= not(layer6_outputs(1650));
    outputs(353) <= not((layer6_outputs(1992)) xor (layer6_outputs(1213)));
    outputs(354) <= not((layer6_outputs(2455)) and (layer6_outputs(1129)));
    outputs(355) <= (layer6_outputs(393)) and not (layer6_outputs(1481));
    outputs(356) <= not(layer6_outputs(2434));
    outputs(357) <= layer6_outputs(2381);
    outputs(358) <= (layer6_outputs(418)) xor (layer6_outputs(52));
    outputs(359) <= layer6_outputs(2262);
    outputs(360) <= not(layer6_outputs(1078));
    outputs(361) <= not(layer6_outputs(1080));
    outputs(362) <= layer6_outputs(2222);
    outputs(363) <= not(layer6_outputs(1685));
    outputs(364) <= layer6_outputs(2553);
    outputs(365) <= not((layer6_outputs(2551)) or (layer6_outputs(1352)));
    outputs(366) <= (layer6_outputs(2215)) and not (layer6_outputs(2047));
    outputs(367) <= not((layer6_outputs(1337)) or (layer6_outputs(738)));
    outputs(368) <= (layer6_outputs(2247)) and not (layer6_outputs(850));
    outputs(369) <= not((layer6_outputs(1837)) xor (layer6_outputs(2107)));
    outputs(370) <= not(layer6_outputs(1359));
    outputs(371) <= layer6_outputs(1158);
    outputs(372) <= not(layer6_outputs(320));
    outputs(373) <= (layer6_outputs(1983)) xor (layer6_outputs(298));
    outputs(374) <= layer6_outputs(1381);
    outputs(375) <= layer6_outputs(2296);
    outputs(376) <= not(layer6_outputs(559));
    outputs(377) <= not(layer6_outputs(1979));
    outputs(378) <= layer6_outputs(885);
    outputs(379) <= not(layer6_outputs(1466));
    outputs(380) <= (layer6_outputs(86)) and not (layer6_outputs(2008));
    outputs(381) <= (layer6_outputs(2261)) xor (layer6_outputs(242));
    outputs(382) <= not(layer6_outputs(1103));
    outputs(383) <= layer6_outputs(2053);
    outputs(384) <= not(layer6_outputs(739));
    outputs(385) <= layer6_outputs(1267);
    outputs(386) <= (layer6_outputs(94)) and (layer6_outputs(2136));
    outputs(387) <= not(layer6_outputs(1948));
    outputs(388) <= (layer6_outputs(1943)) xor (layer6_outputs(1388));
    outputs(389) <= not((layer6_outputs(2061)) xor (layer6_outputs(2325)));
    outputs(390) <= layer6_outputs(138);
    outputs(391) <= layer6_outputs(1933);
    outputs(392) <= layer6_outputs(840);
    outputs(393) <= (layer6_outputs(2556)) xor (layer6_outputs(699));
    outputs(394) <= not(layer6_outputs(1319));
    outputs(395) <= layer6_outputs(1839);
    outputs(396) <= not(layer6_outputs(341));
    outputs(397) <= layer6_outputs(275);
    outputs(398) <= not(layer6_outputs(2383));
    outputs(399) <= (layer6_outputs(564)) or (layer6_outputs(863));
    outputs(400) <= layer6_outputs(1958);
    outputs(401) <= not(layer6_outputs(926));
    outputs(402) <= not(layer6_outputs(517));
    outputs(403) <= (layer6_outputs(1136)) and not (layer6_outputs(1985));
    outputs(404) <= (layer6_outputs(2286)) and (layer6_outputs(235));
    outputs(405) <= layer6_outputs(64);
    outputs(406) <= layer6_outputs(804);
    outputs(407) <= layer6_outputs(2216);
    outputs(408) <= (layer6_outputs(1330)) xor (layer6_outputs(1662));
    outputs(409) <= not((layer6_outputs(232)) xor (layer6_outputs(508)));
    outputs(410) <= layer6_outputs(681);
    outputs(411) <= not(layer6_outputs(1656));
    outputs(412) <= (layer6_outputs(2293)) and (layer6_outputs(1705));
    outputs(413) <= (layer6_outputs(332)) and not (layer6_outputs(114));
    outputs(414) <= layer6_outputs(1309);
    outputs(415) <= layer6_outputs(1028);
    outputs(416) <= (layer6_outputs(185)) and not (layer6_outputs(1750));
    outputs(417) <= not(layer6_outputs(600));
    outputs(418) <= (layer6_outputs(676)) xor (layer6_outputs(1962));
    outputs(419) <= not(layer6_outputs(796));
    outputs(420) <= (layer6_outputs(1517)) and not (layer6_outputs(1613));
    outputs(421) <= layer6_outputs(37);
    outputs(422) <= (layer6_outputs(1483)) and not (layer6_outputs(968));
    outputs(423) <= layer6_outputs(1274);
    outputs(424) <= not(layer6_outputs(765));
    outputs(425) <= (layer6_outputs(1148)) and (layer6_outputs(2151));
    outputs(426) <= not(layer6_outputs(33));
    outputs(427) <= not(layer6_outputs(2197));
    outputs(428) <= not(layer6_outputs(541));
    outputs(429) <= not(layer6_outputs(1684));
    outputs(430) <= not((layer6_outputs(41)) or (layer6_outputs(2525)));
    outputs(431) <= not((layer6_outputs(2479)) or (layer6_outputs(2314)));
    outputs(432) <= not(layer6_outputs(101));
    outputs(433) <= not(layer6_outputs(1830));
    outputs(434) <= not((layer6_outputs(1098)) xor (layer6_outputs(2212)));
    outputs(435) <= not((layer6_outputs(1313)) xor (layer6_outputs(864)));
    outputs(436) <= (layer6_outputs(1322)) and not (layer6_outputs(1800));
    outputs(437) <= (layer6_outputs(1670)) and (layer6_outputs(827));
    outputs(438) <= layer6_outputs(1241);
    outputs(439) <= not((layer6_outputs(902)) or (layer6_outputs(385)));
    outputs(440) <= (layer6_outputs(2212)) xor (layer6_outputs(1603));
    outputs(441) <= layer6_outputs(2179);
    outputs(442) <= not(layer6_outputs(652));
    outputs(443) <= not(layer6_outputs(693));
    outputs(444) <= not((layer6_outputs(795)) xor (layer6_outputs(2225)));
    outputs(445) <= layer6_outputs(2216);
    outputs(446) <= layer6_outputs(1810);
    outputs(447) <= (layer6_outputs(50)) xor (layer6_outputs(2120));
    outputs(448) <= layer6_outputs(1381);
    outputs(449) <= layer6_outputs(1463);
    outputs(450) <= layer6_outputs(2295);
    outputs(451) <= not(layer6_outputs(506));
    outputs(452) <= (layer6_outputs(1930)) xor (layer6_outputs(761));
    outputs(453) <= (layer6_outputs(2086)) and (layer6_outputs(2355));
    outputs(454) <= (layer6_outputs(264)) and (layer6_outputs(1152));
    outputs(455) <= layer6_outputs(1732);
    outputs(456) <= not(layer6_outputs(1643));
    outputs(457) <= (layer6_outputs(2384)) xor (layer6_outputs(2274));
    outputs(458) <= not(layer6_outputs(525));
    outputs(459) <= layer6_outputs(1777);
    outputs(460) <= (layer6_outputs(627)) and not (layer6_outputs(1273));
    outputs(461) <= (layer6_outputs(1704)) and not (layer6_outputs(18));
    outputs(462) <= (layer6_outputs(2463)) xor (layer6_outputs(1141));
    outputs(463) <= layer6_outputs(561);
    outputs(464) <= not((layer6_outputs(2389)) xor (layer6_outputs(1410)));
    outputs(465) <= layer6_outputs(953);
    outputs(466) <= not((layer6_outputs(2450)) or (layer6_outputs(758)));
    outputs(467) <= (layer6_outputs(403)) xor (layer6_outputs(413));
    outputs(468) <= (layer6_outputs(1438)) and not (layer6_outputs(688));
    outputs(469) <= layer6_outputs(1284);
    outputs(470) <= (layer6_outputs(2340)) xor (layer6_outputs(1588));
    outputs(471) <= layer6_outputs(1940);
    outputs(472) <= (layer6_outputs(31)) and (layer6_outputs(547));
    outputs(473) <= (layer6_outputs(612)) and not (layer6_outputs(2324));
    outputs(474) <= layer6_outputs(1548);
    outputs(475) <= not((layer6_outputs(492)) and (layer6_outputs(1607)));
    outputs(476) <= layer6_outputs(1618);
    outputs(477) <= not(layer6_outputs(2346));
    outputs(478) <= layer6_outputs(67);
    outputs(479) <= not((layer6_outputs(805)) or (layer6_outputs(544)));
    outputs(480) <= layer6_outputs(971);
    outputs(481) <= not(layer6_outputs(472));
    outputs(482) <= (layer6_outputs(2052)) and not (layer6_outputs(131));
    outputs(483) <= not(layer6_outputs(1522));
    outputs(484) <= not((layer6_outputs(2420)) xor (layer6_outputs(2464)));
    outputs(485) <= not((layer6_outputs(1847)) xor (layer6_outputs(315)));
    outputs(486) <= not(layer6_outputs(2172));
    outputs(487) <= layer6_outputs(296);
    outputs(488) <= (layer6_outputs(123)) or (layer6_outputs(995));
    outputs(489) <= not((layer6_outputs(886)) xor (layer6_outputs(458)));
    outputs(490) <= (layer6_outputs(2008)) xor (layer6_outputs(1840));
    outputs(491) <= layer6_outputs(2104);
    outputs(492) <= not(layer6_outputs(2476));
    outputs(493) <= (layer6_outputs(2256)) xor (layer6_outputs(1500));
    outputs(494) <= not(layer6_outputs(228));
    outputs(495) <= layer6_outputs(1766);
    outputs(496) <= not(layer6_outputs(889));
    outputs(497) <= (layer6_outputs(1042)) and not (layer6_outputs(1937));
    outputs(498) <= (layer6_outputs(1523)) and not (layer6_outputs(2106));
    outputs(499) <= layer6_outputs(1250);
    outputs(500) <= layer6_outputs(1303);
    outputs(501) <= layer6_outputs(1424);
    outputs(502) <= (layer6_outputs(2106)) xor (layer6_outputs(2558));
    outputs(503) <= layer6_outputs(1185);
    outputs(504) <= not(layer6_outputs(57));
    outputs(505) <= (layer6_outputs(890)) and not (layer6_outputs(1530));
    outputs(506) <= layer6_outputs(1335);
    outputs(507) <= not((layer6_outputs(824)) xor (layer6_outputs(988)));
    outputs(508) <= not((layer6_outputs(346)) or (layer6_outputs(190)));
    outputs(509) <= layer6_outputs(920);
    outputs(510) <= layer6_outputs(1975);
    outputs(511) <= not(layer6_outputs(1472));
    outputs(512) <= (layer6_outputs(917)) xor (layer6_outputs(269));
    outputs(513) <= not((layer6_outputs(1043)) xor (layer6_outputs(1472)));
    outputs(514) <= not((layer6_outputs(2075)) or (layer6_outputs(876)));
    outputs(515) <= layer6_outputs(17);
    outputs(516) <= (layer6_outputs(708)) and (layer6_outputs(66));
    outputs(517) <= not((layer6_outputs(2276)) xor (layer6_outputs(543)));
    outputs(518) <= layer6_outputs(17);
    outputs(519) <= not(layer6_outputs(46)) or (layer6_outputs(533));
    outputs(520) <= (layer6_outputs(2324)) and not (layer6_outputs(1060));
    outputs(521) <= not(layer6_outputs(72));
    outputs(522) <= layer6_outputs(623);
    outputs(523) <= layer6_outputs(151);
    outputs(524) <= not(layer6_outputs(1181));
    outputs(525) <= not(layer6_outputs(620));
    outputs(526) <= layer6_outputs(1725);
    outputs(527) <= layer6_outputs(602);
    outputs(528) <= not(layer6_outputs(15));
    outputs(529) <= (layer6_outputs(822)) and not (layer6_outputs(1921));
    outputs(530) <= not(layer6_outputs(1709));
    outputs(531) <= layer6_outputs(1781);
    outputs(532) <= not(layer6_outputs(2512));
    outputs(533) <= not(layer6_outputs(323));
    outputs(534) <= layer6_outputs(1282);
    outputs(535) <= not(layer6_outputs(1122));
    outputs(536) <= not(layer6_outputs(1487));
    outputs(537) <= layer6_outputs(81);
    outputs(538) <= (layer6_outputs(289)) xor (layer6_outputs(1217));
    outputs(539) <= layer6_outputs(488);
    outputs(540) <= not((layer6_outputs(1176)) xor (layer6_outputs(631)));
    outputs(541) <= not(layer6_outputs(287));
    outputs(542) <= not((layer6_outputs(291)) and (layer6_outputs(1785)));
    outputs(543) <= not(layer6_outputs(241));
    outputs(544) <= not(layer6_outputs(1857));
    outputs(545) <= layer6_outputs(1845);
    outputs(546) <= (layer6_outputs(1676)) and not (layer6_outputs(1304));
    outputs(547) <= not(layer6_outputs(502)) or (layer6_outputs(342));
    outputs(548) <= not(layer6_outputs(1218));
    outputs(549) <= layer6_outputs(2035);
    outputs(550) <= not(layer6_outputs(1119));
    outputs(551) <= (layer6_outputs(1758)) xor (layer6_outputs(2299));
    outputs(552) <= not(layer6_outputs(2059));
    outputs(553) <= not(layer6_outputs(2069));
    outputs(554) <= (layer6_outputs(2191)) and not (layer6_outputs(411));
    outputs(555) <= (layer6_outputs(1423)) and not (layer6_outputs(1167));
    outputs(556) <= not((layer6_outputs(1082)) xor (layer6_outputs(845)));
    outputs(557) <= layer6_outputs(317);
    outputs(558) <= not(layer6_outputs(684));
    outputs(559) <= (layer6_outputs(496)) xor (layer6_outputs(1871));
    outputs(560) <= (layer6_outputs(155)) xor (layer6_outputs(1815));
    outputs(561) <= not(layer6_outputs(274));
    outputs(562) <= not(layer6_outputs(1800));
    outputs(563) <= (layer6_outputs(649)) xor (layer6_outputs(1813));
    outputs(564) <= not((layer6_outputs(2438)) or (layer6_outputs(1030)));
    outputs(565) <= layer6_outputs(1755);
    outputs(566) <= not(layer6_outputs(913));
    outputs(567) <= not(layer6_outputs(1165));
    outputs(568) <= layer6_outputs(189);
    outputs(569) <= (layer6_outputs(2418)) and not (layer6_outputs(958));
    outputs(570) <= layer6_outputs(121);
    outputs(571) <= layer6_outputs(2416);
    outputs(572) <= layer6_outputs(1728);
    outputs(573) <= not(layer6_outputs(2210));
    outputs(574) <= not(layer6_outputs(375)) or (layer6_outputs(2113));
    outputs(575) <= layer6_outputs(1548);
    outputs(576) <= not(layer6_outputs(1088));
    outputs(577) <= not(layer6_outputs(1677));
    outputs(578) <= layer6_outputs(889);
    outputs(579) <= not(layer6_outputs(1163));
    outputs(580) <= (layer6_outputs(1416)) and not (layer6_outputs(978));
    outputs(581) <= not((layer6_outputs(2382)) xor (layer6_outputs(2122)));
    outputs(582) <= layer6_outputs(1193);
    outputs(583) <= not(layer6_outputs(2411));
    outputs(584) <= not((layer6_outputs(455)) xor (layer6_outputs(1747)));
    outputs(585) <= not((layer6_outputs(537)) xor (layer6_outputs(2255)));
    outputs(586) <= not(layer6_outputs(1877));
    outputs(587) <= layer6_outputs(956);
    outputs(588) <= layer6_outputs(348);
    outputs(589) <= layer6_outputs(2505);
    outputs(590) <= layer6_outputs(602);
    outputs(591) <= (layer6_outputs(781)) and (layer6_outputs(48));
    outputs(592) <= layer6_outputs(1040);
    outputs(593) <= not(layer6_outputs(2330));
    outputs(594) <= layer6_outputs(1029);
    outputs(595) <= layer6_outputs(950);
    outputs(596) <= layer6_outputs(647);
    outputs(597) <= not(layer6_outputs(75));
    outputs(598) <= not(layer6_outputs(512));
    outputs(599) <= not(layer6_outputs(2522));
    outputs(600) <= layer6_outputs(2321);
    outputs(601) <= not((layer6_outputs(1042)) xor (layer6_outputs(569)));
    outputs(602) <= not(layer6_outputs(986)) or (layer6_outputs(321));
    outputs(603) <= layer6_outputs(1544);
    outputs(604) <= layer6_outputs(1219);
    outputs(605) <= not(layer6_outputs(2228));
    outputs(606) <= not(layer6_outputs(1134));
    outputs(607) <= (layer6_outputs(339)) and not (layer6_outputs(545));
    outputs(608) <= not((layer6_outputs(400)) or (layer6_outputs(334)));
    outputs(609) <= layer6_outputs(2086);
    outputs(610) <= (layer6_outputs(197)) xor (layer6_outputs(1655));
    outputs(611) <= not((layer6_outputs(844)) or (layer6_outputs(2460)));
    outputs(612) <= not(layer6_outputs(1341));
    outputs(613) <= (layer6_outputs(2537)) and not (layer6_outputs(448));
    outputs(614) <= layer6_outputs(2531);
    outputs(615) <= layer6_outputs(61);
    outputs(616) <= layer6_outputs(2350);
    outputs(617) <= layer6_outputs(1430);
    outputs(618) <= (layer6_outputs(1721)) and (layer6_outputs(598));
    outputs(619) <= (layer6_outputs(1463)) xor (layer6_outputs(1738));
    outputs(620) <= not(layer6_outputs(2353));
    outputs(621) <= (layer6_outputs(803)) and not (layer6_outputs(1697));
    outputs(622) <= not((layer6_outputs(1096)) xor (layer6_outputs(2148)));
    outputs(623) <= layer6_outputs(1524);
    outputs(624) <= not(layer6_outputs(2133));
    outputs(625) <= not((layer6_outputs(1028)) or (layer6_outputs(671)));
    outputs(626) <= layer6_outputs(237);
    outputs(627) <= not((layer6_outputs(1275)) and (layer6_outputs(817)));
    outputs(628) <= layer6_outputs(755);
    outputs(629) <= not(layer6_outputs(1891));
    outputs(630) <= not(layer6_outputs(2294));
    outputs(631) <= not(layer6_outputs(2057));
    outputs(632) <= (layer6_outputs(2195)) and (layer6_outputs(556));
    outputs(633) <= (layer6_outputs(21)) xor (layer6_outputs(1310));
    outputs(634) <= not(layer6_outputs(1857));
    outputs(635) <= layer6_outputs(1940);
    outputs(636) <= not((layer6_outputs(1362)) xor (layer6_outputs(2030)));
    outputs(637) <= layer6_outputs(2328);
    outputs(638) <= not(layer6_outputs(154));
    outputs(639) <= layer6_outputs(2504);
    outputs(640) <= layer6_outputs(1574);
    outputs(641) <= layer6_outputs(1771);
    outputs(642) <= layer6_outputs(1278);
    outputs(643) <= layer6_outputs(1580);
    outputs(644) <= layer6_outputs(2546);
    outputs(645) <= layer6_outputs(974);
    outputs(646) <= not(layer6_outputs(1111));
    outputs(647) <= not((layer6_outputs(403)) xor (layer6_outputs(1259)));
    outputs(648) <= not(layer6_outputs(2485));
    outputs(649) <= (layer6_outputs(962)) or (layer6_outputs(1351));
    outputs(650) <= layer6_outputs(129);
    outputs(651) <= layer6_outputs(1936);
    outputs(652) <= not((layer6_outputs(629)) xor (layer6_outputs(218)));
    outputs(653) <= (layer6_outputs(354)) xor (layer6_outputs(2376));
    outputs(654) <= layer6_outputs(806);
    outputs(655) <= not((layer6_outputs(2206)) or (layer6_outputs(1570)));
    outputs(656) <= not(layer6_outputs(2175));
    outputs(657) <= not((layer6_outputs(630)) or (layer6_outputs(1955)));
    outputs(658) <= not(layer6_outputs(1482));
    outputs(659) <= not(layer6_outputs(1320));
    outputs(660) <= not(layer6_outputs(443));
    outputs(661) <= layer6_outputs(170);
    outputs(662) <= not(layer6_outputs(1778));
    outputs(663) <= layer6_outputs(1444);
    outputs(664) <= not(layer6_outputs(2479));
    outputs(665) <= (layer6_outputs(2343)) and not (layer6_outputs(93));
    outputs(666) <= layer6_outputs(2187);
    outputs(667) <= not(layer6_outputs(1057));
    outputs(668) <= layer6_outputs(1233);
    outputs(669) <= (layer6_outputs(2514)) xor (layer6_outputs(482));
    outputs(670) <= (layer6_outputs(369)) xor (layer6_outputs(1412));
    outputs(671) <= layer6_outputs(1554);
    outputs(672) <= not(layer6_outputs(305));
    outputs(673) <= not(layer6_outputs(1804));
    outputs(674) <= not(layer6_outputs(948));
    outputs(675) <= not((layer6_outputs(2322)) xor (layer6_outputs(1941)));
    outputs(676) <= layer6_outputs(644);
    outputs(677) <= not((layer6_outputs(1016)) or (layer6_outputs(2252)));
    outputs(678) <= not(layer6_outputs(1184));
    outputs(679) <= (layer6_outputs(2021)) xor (layer6_outputs(1073));
    outputs(680) <= layer6_outputs(164);
    outputs(681) <= not((layer6_outputs(574)) xor (layer6_outputs(2070)));
    outputs(682) <= not((layer6_outputs(1914)) or (layer6_outputs(1550)));
    outputs(683) <= (layer6_outputs(679)) xor (layer6_outputs(1926));
    outputs(684) <= layer6_outputs(1532);
    outputs(685) <= layer6_outputs(1547);
    outputs(686) <= layer6_outputs(1654);
    outputs(687) <= layer6_outputs(2083);
    outputs(688) <= not(layer6_outputs(307));
    outputs(689) <= layer6_outputs(267);
    outputs(690) <= layer6_outputs(961);
    outputs(691) <= not(layer6_outputs(258));
    outputs(692) <= layer6_outputs(841);
    outputs(693) <= (layer6_outputs(167)) xor (layer6_outputs(43));
    outputs(694) <= not(layer6_outputs(2206));
    outputs(695) <= (layer6_outputs(2459)) and not (layer6_outputs(9));
    outputs(696) <= layer6_outputs(1748);
    outputs(697) <= not((layer6_outputs(732)) xor (layer6_outputs(307)));
    outputs(698) <= not(layer6_outputs(1150));
    outputs(699) <= not(layer6_outputs(2075));
    outputs(700) <= layer6_outputs(509);
    outputs(701) <= layer6_outputs(970);
    outputs(702) <= layer6_outputs(898);
    outputs(703) <= not(layer6_outputs(1053));
    outputs(704) <= (layer6_outputs(1746)) or (layer6_outputs(414));
    outputs(705) <= not(layer6_outputs(2296));
    outputs(706) <= not((layer6_outputs(1181)) and (layer6_outputs(306)));
    outputs(707) <= not(layer6_outputs(2271)) or (layer6_outputs(740));
    outputs(708) <= not((layer6_outputs(2509)) xor (layer6_outputs(2246)));
    outputs(709) <= layer6_outputs(1108);
    outputs(710) <= not(layer6_outputs(1321));
    outputs(711) <= layer6_outputs(1825);
    outputs(712) <= (layer6_outputs(360)) xor (layer6_outputs(670));
    outputs(713) <= layer6_outputs(1959);
    outputs(714) <= (layer6_outputs(1219)) xor (layer6_outputs(2464));
    outputs(715) <= layer6_outputs(2446);
    outputs(716) <= (layer6_outputs(1453)) and not (layer6_outputs(1044));
    outputs(717) <= not(layer6_outputs(787));
    outputs(718) <= not(layer6_outputs(779));
    outputs(719) <= (layer6_outputs(1893)) xor (layer6_outputs(1043));
    outputs(720) <= not(layer6_outputs(335));
    outputs(721) <= (layer6_outputs(1556)) xor (layer6_outputs(567));
    outputs(722) <= layer6_outputs(1625);
    outputs(723) <= not(layer6_outputs(268));
    outputs(724) <= layer6_outputs(1351);
    outputs(725) <= (layer6_outputs(75)) xor (layer6_outputs(2387));
    outputs(726) <= layer6_outputs(2418);
    outputs(727) <= not(layer6_outputs(1238));
    outputs(728) <= not((layer6_outputs(1363)) xor (layer6_outputs(2355)));
    outputs(729) <= (layer6_outputs(2547)) and (layer6_outputs(1795));
    outputs(730) <= layer6_outputs(780);
    outputs(731) <= layer6_outputs(182);
    outputs(732) <= not(layer6_outputs(2336));
    outputs(733) <= layer6_outputs(2178);
    outputs(734) <= not((layer6_outputs(58)) xor (layer6_outputs(1928)));
    outputs(735) <= not(layer6_outputs(72));
    outputs(736) <= layer6_outputs(250);
    outputs(737) <= not(layer6_outputs(286));
    outputs(738) <= not(layer6_outputs(916));
    outputs(739) <= not(layer6_outputs(1419));
    outputs(740) <= layer6_outputs(941);
    outputs(741) <= not(layer6_outputs(1200));
    outputs(742) <= not(layer6_outputs(520));
    outputs(743) <= not(layer6_outputs(2186));
    outputs(744) <= layer6_outputs(2054);
    outputs(745) <= (layer6_outputs(2493)) xor (layer6_outputs(1941));
    outputs(746) <= not(layer6_outputs(769));
    outputs(747) <= not((layer6_outputs(2352)) xor (layer6_outputs(1452)));
    outputs(748) <= not((layer6_outputs(1745)) xor (layer6_outputs(171)));
    outputs(749) <= (layer6_outputs(970)) and not (layer6_outputs(222));
    outputs(750) <= layer6_outputs(2549);
    outputs(751) <= layer6_outputs(1129);
    outputs(752) <= not(layer6_outputs(570)) or (layer6_outputs(2191));
    outputs(753) <= not(layer6_outputs(1039));
    outputs(754) <= layer6_outputs(2055);
    outputs(755) <= layer6_outputs(1308);
    outputs(756) <= not((layer6_outputs(2535)) xor (layer6_outputs(1682)));
    outputs(757) <= not(layer6_outputs(1767));
    outputs(758) <= layer6_outputs(964);
    outputs(759) <= (layer6_outputs(1781)) and (layer6_outputs(1735));
    outputs(760) <= not(layer6_outputs(786));
    outputs(761) <= layer6_outputs(1124);
    outputs(762) <= not(layer6_outputs(1589));
    outputs(763) <= (layer6_outputs(198)) xor (layer6_outputs(1323));
    outputs(764) <= not(layer6_outputs(1094));
    outputs(765) <= layer6_outputs(2159);
    outputs(766) <= not(layer6_outputs(1703));
    outputs(767) <= not(layer6_outputs(2390));
    outputs(768) <= not((layer6_outputs(2233)) xor (layer6_outputs(949)));
    outputs(769) <= layer6_outputs(2181);
    outputs(770) <= layer6_outputs(1515);
    outputs(771) <= not(layer6_outputs(1156));
    outputs(772) <= '1';
    outputs(773) <= not(layer6_outputs(1433));
    outputs(774) <= layer6_outputs(919);
    outputs(775) <= not((layer6_outputs(1099)) xor (layer6_outputs(200)));
    outputs(776) <= not(layer6_outputs(566));
    outputs(777) <= not(layer6_outputs(1169));
    outputs(778) <= layer6_outputs(73);
    outputs(779) <= layer6_outputs(2401);
    outputs(780) <= (layer6_outputs(1698)) xor (layer6_outputs(1047));
    outputs(781) <= not(layer6_outputs(714));
    outputs(782) <= (layer6_outputs(365)) xor (layer6_outputs(1447));
    outputs(783) <= not((layer6_outputs(858)) xor (layer6_outputs(2253)));
    outputs(784) <= (layer6_outputs(2524)) xor (layer6_outputs(129));
    outputs(785) <= (layer6_outputs(847)) and (layer6_outputs(782));
    outputs(786) <= (layer6_outputs(1456)) xor (layer6_outputs(1506));
    outputs(787) <= layer6_outputs(83);
    outputs(788) <= layer6_outputs(2430);
    outputs(789) <= layer6_outputs(2128);
    outputs(790) <= (layer6_outputs(548)) xor (layer6_outputs(2302));
    outputs(791) <= not(layer6_outputs(1900));
    outputs(792) <= layer6_outputs(2532);
    outputs(793) <= not(layer6_outputs(785));
    outputs(794) <= layer6_outputs(1478);
    outputs(795) <= layer6_outputs(85);
    outputs(796) <= (layer6_outputs(1559)) xor (layer6_outputs(1407));
    outputs(797) <= (layer6_outputs(1147)) xor (layer6_outputs(505));
    outputs(798) <= layer6_outputs(1706);
    outputs(799) <= not(layer6_outputs(104));
    outputs(800) <= not(layer6_outputs(798));
    outputs(801) <= not(layer6_outputs(89));
    outputs(802) <= not(layer6_outputs(2531));
    outputs(803) <= not((layer6_outputs(488)) xor (layer6_outputs(1932)));
    outputs(804) <= not(layer6_outputs(1274));
    outputs(805) <= not((layer6_outputs(1776)) or (layer6_outputs(210)));
    outputs(806) <= layer6_outputs(1060);
    outputs(807) <= layer6_outputs(932);
    outputs(808) <= not(layer6_outputs(143));
    outputs(809) <= not(layer6_outputs(2252));
    outputs(810) <= (layer6_outputs(2415)) and not (layer6_outputs(2530));
    outputs(811) <= not(layer6_outputs(783));
    outputs(812) <= not((layer6_outputs(2130)) xor (layer6_outputs(357)));
    outputs(813) <= (layer6_outputs(434)) and (layer6_outputs(597));
    outputs(814) <= layer6_outputs(1746);
    outputs(815) <= not((layer6_outputs(266)) and (layer6_outputs(95)));
    outputs(816) <= layer6_outputs(755);
    outputs(817) <= layer6_outputs(796);
    outputs(818) <= not((layer6_outputs(2199)) xor (layer6_outputs(1736)));
    outputs(819) <= not(layer6_outputs(1246));
    outputs(820) <= (layer6_outputs(667)) xor (layer6_outputs(2155));
    outputs(821) <= not((layer6_outputs(1715)) and (layer6_outputs(1517)));
    outputs(822) <= not((layer6_outputs(1705)) xor (layer6_outputs(556)));
    outputs(823) <= layer6_outputs(927);
    outputs(824) <= not((layer6_outputs(1955)) or (layer6_outputs(1918)));
    outputs(825) <= layer6_outputs(2405);
    outputs(826) <= (layer6_outputs(166)) and (layer6_outputs(1346));
    outputs(827) <= not(layer6_outputs(1153));
    outputs(828) <= (layer6_outputs(387)) and (layer6_outputs(2441));
    outputs(829) <= (layer6_outputs(2516)) and not (layer6_outputs(2431));
    outputs(830) <= (layer6_outputs(2491)) xor (layer6_outputs(2199));
    outputs(831) <= not(layer6_outputs(2511));
    outputs(832) <= not(layer6_outputs(105));
    outputs(833) <= (layer6_outputs(1312)) xor (layer6_outputs(2149));
    outputs(834) <= (layer6_outputs(753)) and not (layer6_outputs(2481));
    outputs(835) <= layer6_outputs(1237);
    outputs(836) <= (layer6_outputs(2250)) xor (layer6_outputs(1862));
    outputs(837) <= not((layer6_outputs(1571)) xor (layer6_outputs(1059)));
    outputs(838) <= (layer6_outputs(767)) and not (layer6_outputs(2457));
    outputs(839) <= not((layer6_outputs(2046)) xor (layer6_outputs(1584)));
    outputs(840) <= (layer6_outputs(1091)) and (layer6_outputs(1369));
    outputs(841) <= layer6_outputs(1293);
    outputs(842) <= not(layer6_outputs(1747));
    outputs(843) <= not((layer6_outputs(1868)) xor (layer6_outputs(2190)));
    outputs(844) <= not(layer6_outputs(188));
    outputs(845) <= (layer6_outputs(399)) xor (layer6_outputs(2268));
    outputs(846) <= layer6_outputs(1828);
    outputs(847) <= layer6_outputs(190);
    outputs(848) <= (layer6_outputs(2147)) and not (layer6_outputs(2233));
    outputs(849) <= layer6_outputs(1582);
    outputs(850) <= (layer6_outputs(2116)) xor (layer6_outputs(1843));
    outputs(851) <= not((layer6_outputs(1328)) or (layer6_outputs(1328)));
    outputs(852) <= (layer6_outputs(1107)) and not (layer6_outputs(1049));
    outputs(853) <= (layer6_outputs(1247)) xor (layer6_outputs(2129));
    outputs(854) <= (layer6_outputs(1019)) xor (layer6_outputs(165));
    outputs(855) <= not(layer6_outputs(1195));
    outputs(856) <= not(layer6_outputs(1639));
    outputs(857) <= not(layer6_outputs(444));
    outputs(858) <= (layer6_outputs(1300)) xor (layer6_outputs(2026));
    outputs(859) <= not((layer6_outputs(833)) xor (layer6_outputs(1198)));
    outputs(860) <= not(layer6_outputs(756));
    outputs(861) <= layer6_outputs(595);
    outputs(862) <= layer6_outputs(2151);
    outputs(863) <= not(layer6_outputs(898));
    outputs(864) <= (layer6_outputs(896)) and (layer6_outputs(220));
    outputs(865) <= not((layer6_outputs(793)) xor (layer6_outputs(27)));
    outputs(866) <= layer6_outputs(1136);
    outputs(867) <= layer6_outputs(834);
    outputs(868) <= not(layer6_outputs(1966));
    outputs(869) <= layer6_outputs(2521);
    outputs(870) <= not((layer6_outputs(957)) or (layer6_outputs(1634)));
    outputs(871) <= layer6_outputs(1172);
    outputs(872) <= not(layer6_outputs(409));
    outputs(873) <= (layer6_outputs(629)) and (layer6_outputs(603));
    outputs(874) <= not((layer6_outputs(2483)) or (layer6_outputs(407)));
    outputs(875) <= layer6_outputs(1037);
    outputs(876) <= (layer6_outputs(202)) xor (layer6_outputs(397));
    outputs(877) <= not(layer6_outputs(2316));
    outputs(878) <= layer6_outputs(627);
    outputs(879) <= not(layer6_outputs(173));
    outputs(880) <= not((layer6_outputs(1051)) xor (layer6_outputs(924)));
    outputs(881) <= not((layer6_outputs(2068)) xor (layer6_outputs(6)));
    outputs(882) <= (layer6_outputs(465)) and (layer6_outputs(2214));
    outputs(883) <= not(layer6_outputs(328));
    outputs(884) <= not(layer6_outputs(1317));
    outputs(885) <= layer6_outputs(1510);
    outputs(886) <= layer6_outputs(542);
    outputs(887) <= layer6_outputs(1897);
    outputs(888) <= (layer6_outputs(2182)) xor (layer6_outputs(398));
    outputs(889) <= not(layer6_outputs(42));
    outputs(890) <= layer6_outputs(435);
    outputs(891) <= not(layer6_outputs(809));
    outputs(892) <= not(layer6_outputs(2433));
    outputs(893) <= not(layer6_outputs(318));
    outputs(894) <= layer6_outputs(675);
    outputs(895) <= layer6_outputs(192);
    outputs(896) <= not(layer6_outputs(2490));
    outputs(897) <= layer6_outputs(1417);
    outputs(898) <= (layer6_outputs(1744)) xor (layer6_outputs(1947));
    outputs(899) <= (layer6_outputs(1407)) xor (layer6_outputs(1397));
    outputs(900) <= layer6_outputs(343);
    outputs(901) <= not((layer6_outputs(1910)) xor (layer6_outputs(100)));
    outputs(902) <= layer6_outputs(2213);
    outputs(903) <= layer6_outputs(1845);
    outputs(904) <= not((layer6_outputs(567)) xor (layer6_outputs(2278)));
    outputs(905) <= not(layer6_outputs(200));
    outputs(906) <= not(layer6_outputs(67));
    outputs(907) <= not(layer6_outputs(2092));
    outputs(908) <= layer6_outputs(1027);
    outputs(909) <= not(layer6_outputs(2329));
    outputs(910) <= not((layer6_outputs(2510)) xor (layer6_outputs(810)));
    outputs(911) <= not((layer6_outputs(2185)) or (layer6_outputs(637)));
    outputs(912) <= not((layer6_outputs(1743)) xor (layer6_outputs(2077)));
    outputs(913) <= layer6_outputs(1830);
    outputs(914) <= layer6_outputs(1004);
    outputs(915) <= layer6_outputs(254);
    outputs(916) <= (layer6_outputs(209)) xor (layer6_outputs(725));
    outputs(917) <= layer6_outputs(2005);
    outputs(918) <= layer6_outputs(1971);
    outputs(919) <= (layer6_outputs(1823)) and (layer6_outputs(933));
    outputs(920) <= not(layer6_outputs(1814));
    outputs(921) <= not(layer6_outputs(1020));
    outputs(922) <= layer6_outputs(1390);
    outputs(923) <= not(layer6_outputs(360));
    outputs(924) <= (layer6_outputs(2539)) and not (layer6_outputs(2113));
    outputs(925) <= not(layer6_outputs(155));
    outputs(926) <= not((layer6_outputs(480)) xor (layer6_outputs(296)));
    outputs(927) <= layer6_outputs(80);
    outputs(928) <= not((layer6_outputs(2515)) xor (layer6_outputs(2374)));
    outputs(929) <= layer6_outputs(1521);
    outputs(930) <= layer6_outputs(1408);
    outputs(931) <= layer6_outputs(1925);
    outputs(932) <= not(layer6_outputs(1166));
    outputs(933) <= not(layer6_outputs(528));
    outputs(934) <= (layer6_outputs(1829)) xor (layer6_outputs(1000));
    outputs(935) <= (layer6_outputs(1653)) xor (layer6_outputs(2408));
    outputs(936) <= not(layer6_outputs(1826));
    outputs(937) <= not((layer6_outputs(1307)) xor (layer6_outputs(1760)));
    outputs(938) <= layer6_outputs(2345);
    outputs(939) <= layer6_outputs(2143);
    outputs(940) <= layer6_outputs(1651);
    outputs(941) <= not(layer6_outputs(2306));
    outputs(942) <= not(layer6_outputs(1470));
    outputs(943) <= (layer6_outputs(2040)) xor (layer6_outputs(2359));
    outputs(944) <= (layer6_outputs(1624)) and (layer6_outputs(704));
    outputs(945) <= not(layer6_outputs(2380));
    outputs(946) <= not((layer6_outputs(2235)) xor (layer6_outputs(1291)));
    outputs(947) <= (layer6_outputs(1865)) and not (layer6_outputs(633));
    outputs(948) <= not(layer6_outputs(1744));
    outputs(949) <= not(layer6_outputs(2197));
    outputs(950) <= (layer6_outputs(1368)) xor (layer6_outputs(1889));
    outputs(951) <= layer6_outputs(1755);
    outputs(952) <= layer6_outputs(2269);
    outputs(953) <= (layer6_outputs(1360)) and not (layer6_outputs(1389));
    outputs(954) <= not(layer6_outputs(289));
    outputs(955) <= layer6_outputs(1134);
    outputs(956) <= layer6_outputs(1214);
    outputs(957) <= not(layer6_outputs(1256));
    outputs(958) <= layer6_outputs(1980);
    outputs(959) <= not(layer6_outputs(1757));
    outputs(960) <= (layer6_outputs(2351)) xor (layer6_outputs(1074));
    outputs(961) <= not(layer6_outputs(1578));
    outputs(962) <= not((layer6_outputs(837)) and (layer6_outputs(1919)));
    outputs(963) <= (layer6_outputs(2407)) xor (layer6_outputs(1583));
    outputs(964) <= (layer6_outputs(536)) and not (layer6_outputs(260));
    outputs(965) <= not(layer6_outputs(2242));
    outputs(966) <= not(layer6_outputs(2012));
    outputs(967) <= not(layer6_outputs(424));
    outputs(968) <= not(layer6_outputs(2169));
    outputs(969) <= not(layer6_outputs(1894));
    outputs(970) <= layer6_outputs(1029);
    outputs(971) <= not(layer6_outputs(819));
    outputs(972) <= not((layer6_outputs(664)) and (layer6_outputs(304)));
    outputs(973) <= not((layer6_outputs(118)) xor (layer6_outputs(593)));
    outputs(974) <= (layer6_outputs(2030)) xor (layer6_outputs(342));
    outputs(975) <= layer6_outputs(1732);
    outputs(976) <= not(layer6_outputs(408));
    outputs(977) <= not(layer6_outputs(2483));
    outputs(978) <= not(layer6_outputs(1142));
    outputs(979) <= not((layer6_outputs(1503)) xor (layer6_outputs(2267)));
    outputs(980) <= not(layer6_outputs(2109));
    outputs(981) <= not((layer6_outputs(2550)) xor (layer6_outputs(1010)));
    outputs(982) <= (layer6_outputs(32)) or (layer6_outputs(2330));
    outputs(983) <= not(layer6_outputs(2012)) or (layer6_outputs(1988));
    outputs(984) <= not(layer6_outputs(1148));
    outputs(985) <= layer6_outputs(406);
    outputs(986) <= not(layer6_outputs(1909));
    outputs(987) <= (layer6_outputs(2090)) and not (layer6_outputs(2176));
    outputs(988) <= not((layer6_outputs(1254)) or (layer6_outputs(568)));
    outputs(989) <= layer6_outputs(174);
    outputs(990) <= not(layer6_outputs(744));
    outputs(991) <= layer6_outputs(2126);
    outputs(992) <= layer6_outputs(2474);
    outputs(993) <= layer6_outputs(402);
    outputs(994) <= layer6_outputs(648);
    outputs(995) <= layer6_outputs(481);
    outputs(996) <= not(layer6_outputs(1912));
    outputs(997) <= layer6_outputs(31);
    outputs(998) <= layer6_outputs(2193);
    outputs(999) <= not(layer6_outputs(1394));
    outputs(1000) <= not(layer6_outputs(273));
    outputs(1001) <= not(layer6_outputs(12));
    outputs(1002) <= (layer6_outputs(2360)) and not (layer6_outputs(1109));
    outputs(1003) <= not(layer6_outputs(94));
    outputs(1004) <= (layer6_outputs(2484)) xor (layer6_outputs(389));
    outputs(1005) <= (layer6_outputs(2336)) and not (layer6_outputs(2452));
    outputs(1006) <= layer6_outputs(1540);
    outputs(1007) <= layer6_outputs(501);
    outputs(1008) <= not(layer6_outputs(866));
    outputs(1009) <= not((layer6_outputs(2423)) and (layer6_outputs(2275)));
    outputs(1010) <= not((layer6_outputs(2528)) xor (layer6_outputs(145)));
    outputs(1011) <= layer6_outputs(1340);
    outputs(1012) <= layer6_outputs(208);
    outputs(1013) <= layer6_outputs(1694);
    outputs(1014) <= not(layer6_outputs(1797));
    outputs(1015) <= not((layer6_outputs(2220)) xor (layer6_outputs(1137)));
    outputs(1016) <= not(layer6_outputs(759)) or (layer6_outputs(285));
    outputs(1017) <= (layer6_outputs(1238)) and not (layer6_outputs(141));
    outputs(1018) <= (layer6_outputs(1)) xor (layer6_outputs(2326));
    outputs(1019) <= not(layer6_outputs(1045));
    outputs(1020) <= not(layer6_outputs(1154));
    outputs(1021) <= not(layer6_outputs(1072));
    outputs(1022) <= not((layer6_outputs(1687)) and (layer6_outputs(843)));
    outputs(1023) <= not(layer6_outputs(1982));
    outputs(1024) <= not(layer6_outputs(128));
    outputs(1025) <= not(layer6_outputs(2507));
    outputs(1026) <= layer6_outputs(1799);
    outputs(1027) <= not(layer6_outputs(81));
    outputs(1028) <= not(layer6_outputs(2552));
    outputs(1029) <= layer6_outputs(326);
    outputs(1030) <= (layer6_outputs(1490)) and not (layer6_outputs(521));
    outputs(1031) <= layer6_outputs(394);
    outputs(1032) <= (layer6_outputs(751)) or (layer6_outputs(2519));
    outputs(1033) <= not((layer6_outputs(1577)) or (layer6_outputs(1033)));
    outputs(1034) <= (layer6_outputs(2203)) and not (layer6_outputs(1956));
    outputs(1035) <= layer6_outputs(2281);
    outputs(1036) <= (layer6_outputs(1850)) and not (layer6_outputs(1113));
    outputs(1037) <= not(layer6_outputs(1999));
    outputs(1038) <= not(layer6_outputs(104));
    outputs(1039) <= not(layer6_outputs(2382));
    outputs(1040) <= (layer6_outputs(1647)) and not (layer6_outputs(1933));
    outputs(1041) <= not((layer6_outputs(2279)) xor (layer6_outputs(1538)));
    outputs(1042) <= layer6_outputs(780);
    outputs(1043) <= (layer6_outputs(1292)) xor (layer6_outputs(1298));
    outputs(1044) <= layer6_outputs(2038);
    outputs(1045) <= not(layer6_outputs(747));
    outputs(1046) <= not(layer6_outputs(880));
    outputs(1047) <= layer6_outputs(1553);
    outputs(1048) <= layer6_outputs(238);
    outputs(1049) <= (layer6_outputs(51)) xor (layer6_outputs(2357));
    outputs(1050) <= layer6_outputs(2448);
    outputs(1051) <= not(layer6_outputs(2398));
    outputs(1052) <= not(layer6_outputs(2377));
    outputs(1053) <= not(layer6_outputs(2065));
    outputs(1054) <= not((layer6_outputs(1287)) xor (layer6_outputs(987)));
    outputs(1055) <= '0';
    outputs(1056) <= layer6_outputs(1976);
    outputs(1057) <= not(layer6_outputs(16));
    outputs(1058) <= not((layer6_outputs(1987)) or (layer6_outputs(1298)));
    outputs(1059) <= not(layer6_outputs(1377));
    outputs(1060) <= not(layer6_outputs(227));
    outputs(1061) <= not(layer6_outputs(2135));
    outputs(1062) <= layer6_outputs(1832);
    outputs(1063) <= (layer6_outputs(358)) and (layer6_outputs(2447));
    outputs(1064) <= not((layer6_outputs(309)) xor (layer6_outputs(1535)));
    outputs(1065) <= not((layer6_outputs(2137)) xor (layer6_outputs(730)));
    outputs(1066) <= layer6_outputs(1396);
    outputs(1067) <= layer6_outputs(1215);
    outputs(1068) <= not(layer6_outputs(2264));
    outputs(1069) <= layer6_outputs(2288);
    outputs(1070) <= (layer6_outputs(2477)) xor (layer6_outputs(1858));
    outputs(1071) <= not(layer6_outputs(145)) or (layer6_outputs(1593));
    outputs(1072) <= (layer6_outputs(1003)) xor (layer6_outputs(2489));
    outputs(1073) <= not(layer6_outputs(975));
    outputs(1074) <= not((layer6_outputs(610)) xor (layer6_outputs(396)));
    outputs(1075) <= layer6_outputs(2063);
    outputs(1076) <= not((layer6_outputs(2111)) or (layer6_outputs(2208)));
    outputs(1077) <= (layer6_outputs(2056)) xor (layer6_outputs(784));
    outputs(1078) <= (layer6_outputs(966)) xor (layer6_outputs(996));
    outputs(1079) <= not((layer6_outputs(581)) xor (layer6_outputs(1923)));
    outputs(1080) <= layer6_outputs(1952);
    outputs(1081) <= not((layer6_outputs(1656)) xor (layer6_outputs(1405)));
    outputs(1082) <= not(layer6_outputs(2358));
    outputs(1083) <= layer6_outputs(606);
    outputs(1084) <= (layer6_outputs(737)) and (layer6_outputs(1494));
    outputs(1085) <= not(layer6_outputs(1543));
    outputs(1086) <= not((layer6_outputs(799)) xor (layer6_outputs(4)));
    outputs(1087) <= not(layer6_outputs(982));
    outputs(1088) <= (layer6_outputs(331)) and (layer6_outputs(264));
    outputs(1089) <= layer6_outputs(299);
    outputs(1090) <= layer6_outputs(753);
    outputs(1091) <= layer6_outputs(994);
    outputs(1092) <= (layer6_outputs(139)) xor (layer6_outputs(1147));
    outputs(1093) <= not(layer6_outputs(2196));
    outputs(1094) <= not(layer6_outputs(467)) or (layer6_outputs(1258));
    outputs(1095) <= layer6_outputs(2385);
    outputs(1096) <= (layer6_outputs(648)) and not (layer6_outputs(419));
    outputs(1097) <= layer6_outputs(1098);
    outputs(1098) <= layer6_outputs(405);
    outputs(1099) <= not(layer6_outputs(624));
    outputs(1100) <= not(layer6_outputs(380));
    outputs(1101) <= layer6_outputs(994);
    outputs(1102) <= layer6_outputs(745);
    outputs(1103) <= not((layer6_outputs(742)) xor (layer6_outputs(2293)));
    outputs(1104) <= not(layer6_outputs(517));
    outputs(1105) <= layer6_outputs(717);
    outputs(1106) <= layer6_outputs(1037);
    outputs(1107) <= (layer6_outputs(1567)) and not (layer6_outputs(2170));
    outputs(1108) <= (layer6_outputs(1121)) xor (layer6_outputs(224));
    outputs(1109) <= not(layer6_outputs(1945));
    outputs(1110) <= layer6_outputs(310);
    outputs(1111) <= (layer6_outputs(2334)) xor (layer6_outputs(826));
    outputs(1112) <= layer6_outputs(2469);
    outputs(1113) <= not((layer6_outputs(1157)) or (layer6_outputs(1221)));
    outputs(1114) <= not(layer6_outputs(290));
    outputs(1115) <= layer6_outputs(923);
    outputs(1116) <= not((layer6_outputs(2482)) or (layer6_outputs(1720)));
    outputs(1117) <= layer6_outputs(807);
    outputs(1118) <= (layer6_outputs(913)) and (layer6_outputs(807));
    outputs(1119) <= not((layer6_outputs(294)) xor (layer6_outputs(39)));
    outputs(1120) <= layer6_outputs(271);
    outputs(1121) <= not((layer6_outputs(740)) xor (layer6_outputs(332)));
    outputs(1122) <= not((layer6_outputs(263)) xor (layer6_outputs(718)));
    outputs(1123) <= layer6_outputs(1277);
    outputs(1124) <= not((layer6_outputs(975)) and (layer6_outputs(1579)));
    outputs(1125) <= not(layer6_outputs(1206));
    outputs(1126) <= not(layer6_outputs(1348));
    outputs(1127) <= not(layer6_outputs(186));
    outputs(1128) <= not(layer6_outputs(1425));
    outputs(1129) <= not(layer6_outputs(0));
    outputs(1130) <= layer6_outputs(2424);
    outputs(1131) <= layer6_outputs(263);
    outputs(1132) <= layer6_outputs(1635);
    outputs(1133) <= layer6_outputs(2341);
    outputs(1134) <= layer6_outputs(1128);
    outputs(1135) <= not(layer6_outputs(1083));
    outputs(1136) <= layer6_outputs(1481);
    outputs(1137) <= not(layer6_outputs(1026));
    outputs(1138) <= not(layer6_outputs(1790));
    outputs(1139) <= not(layer6_outputs(1234));
    outputs(1140) <= layer6_outputs(1449);
    outputs(1141) <= not(layer6_outputs(1117));
    outputs(1142) <= not((layer6_outputs(1629)) and (layer6_outputs(2379)));
    outputs(1143) <= not(layer6_outputs(1706));
    outputs(1144) <= not(layer6_outputs(161));
    outputs(1145) <= layer6_outputs(1560);
    outputs(1146) <= layer6_outputs(2506);
    outputs(1147) <= not(layer6_outputs(1901));
    outputs(1148) <= not((layer6_outputs(1360)) xor (layer6_outputs(1235)));
    outputs(1149) <= not(layer6_outputs(1443));
    outputs(1150) <= not(layer6_outputs(1688));
    outputs(1151) <= not(layer6_outputs(1678));
    outputs(1152) <= not((layer6_outputs(78)) xor (layer6_outputs(2530)));
    outputs(1153) <= not(layer6_outputs(1491));
    outputs(1154) <= not(layer6_outputs(724));
    outputs(1155) <= not(layer6_outputs(368));
    outputs(1156) <= layer6_outputs(2424);
    outputs(1157) <= layer6_outputs(133);
    outputs(1158) <= (layer6_outputs(113)) and (layer6_outputs(1190));
    outputs(1159) <= layer6_outputs(2203);
    outputs(1160) <= layer6_outputs(35);
    outputs(1161) <= not(layer6_outputs(854));
    outputs(1162) <= not(layer6_outputs(2171));
    outputs(1163) <= (layer6_outputs(680)) xor (layer6_outputs(1299));
    outputs(1164) <= (layer6_outputs(1531)) and (layer6_outputs(1868));
    outputs(1165) <= (layer6_outputs(293)) xor (layer6_outputs(1588));
    outputs(1166) <= not(layer6_outputs(678));
    outputs(1167) <= layer6_outputs(2144);
    outputs(1168) <= not(layer6_outputs(1434));
    outputs(1169) <= not((layer6_outputs(2363)) xor (layer6_outputs(2145)));
    outputs(1170) <= not((layer6_outputs(1168)) xor (layer6_outputs(444)));
    outputs(1171) <= layer6_outputs(2437);
    outputs(1172) <= layer6_outputs(671);
    outputs(1173) <= not(layer6_outputs(2089));
    outputs(1174) <= not(layer6_outputs(16));
    outputs(1175) <= not((layer6_outputs(1925)) xor (layer6_outputs(1018)));
    outputs(1176) <= layer6_outputs(1768);
    outputs(1177) <= not(layer6_outputs(232));
    outputs(1178) <= (layer6_outputs(433)) and (layer6_outputs(64));
    outputs(1179) <= not((layer6_outputs(210)) xor (layer6_outputs(884)));
    outputs(1180) <= not((layer6_outputs(665)) xor (layer6_outputs(204)));
    outputs(1181) <= not((layer6_outputs(2204)) xor (layer6_outputs(2352)));
    outputs(1182) <= not(layer6_outputs(641));
    outputs(1183) <= not(layer6_outputs(853));
    outputs(1184) <= not(layer6_outputs(2307));
    outputs(1185) <= not((layer6_outputs(2378)) xor (layer6_outputs(2503)));
    outputs(1186) <= not(layer6_outputs(1289));
    outputs(1187) <= (layer6_outputs(1082)) xor (layer6_outputs(1690));
    outputs(1188) <= (layer6_outputs(778)) xor (layer6_outputs(361));
    outputs(1189) <= not(layer6_outputs(2125));
    outputs(1190) <= (layer6_outputs(1252)) xor (layer6_outputs(938));
    outputs(1191) <= layer6_outputs(2371);
    outputs(1192) <= not(layer6_outputs(1036));
    outputs(1193) <= layer6_outputs(141);
    outputs(1194) <= not(layer6_outputs(2123));
    outputs(1195) <= not(layer6_outputs(791));
    outputs(1196) <= not(layer6_outputs(623));
    outputs(1197) <= not((layer6_outputs(1353)) or (layer6_outputs(73)));
    outputs(1198) <= not(layer6_outputs(1657));
    outputs(1199) <= layer6_outputs(466);
    outputs(1200) <= layer6_outputs(1431);
    outputs(1201) <= (layer6_outputs(1687)) xor (layer6_outputs(2034));
    outputs(1202) <= not(layer6_outputs(2311));
    outputs(1203) <= not((layer6_outputs(2270)) xor (layer6_outputs(1337)));
    outputs(1204) <= not(layer6_outputs(1091));
    outputs(1205) <= (layer6_outputs(524)) and not (layer6_outputs(2257));
    outputs(1206) <= not(layer6_outputs(854));
    outputs(1207) <= (layer6_outputs(2334)) or (layer6_outputs(2131));
    outputs(1208) <= (layer6_outputs(730)) xor (layer6_outputs(108));
    outputs(1209) <= not(layer6_outputs(359));
    outputs(1210) <= (layer6_outputs(2370)) xor (layer6_outputs(1569));
    outputs(1211) <= layer6_outputs(1860);
    outputs(1212) <= layer6_outputs(2025);
    outputs(1213) <= not((layer6_outputs(2354)) xor (layer6_outputs(897)));
    outputs(1214) <= (layer6_outputs(1843)) xor (layer6_outputs(1402));
    outputs(1215) <= not((layer6_outputs(2255)) xor (layer6_outputs(1590)));
    outputs(1216) <= layer6_outputs(2059);
    outputs(1217) <= (layer6_outputs(2048)) and (layer6_outputs(2173));
    outputs(1218) <= layer6_outputs(213);
    outputs(1219) <= (layer6_outputs(1567)) and not (layer6_outputs(470));
    outputs(1220) <= (layer6_outputs(692)) xor (layer6_outputs(982));
    outputs(1221) <= layer6_outputs(1595);
    outputs(1222) <= not(layer6_outputs(2043));
    outputs(1223) <= (layer6_outputs(1130)) and (layer6_outputs(1269));
    outputs(1224) <= not(layer6_outputs(424));
    outputs(1225) <= not((layer6_outputs(193)) xor (layer6_outputs(663)));
    outputs(1226) <= not(layer6_outputs(2029));
    outputs(1227) <= not(layer6_outputs(440));
    outputs(1228) <= (layer6_outputs(426)) and not (layer6_outputs(2132));
    outputs(1229) <= (layer6_outputs(1226)) xor (layer6_outputs(908));
    outputs(1230) <= not(layer6_outputs(1646));
    outputs(1231) <= layer6_outputs(926);
    outputs(1232) <= not(layer6_outputs(1403));
    outputs(1233) <= not(layer6_outputs(2308));
    outputs(1234) <= not(layer6_outputs(419));
    outputs(1235) <= not(layer6_outputs(1562));
    outputs(1236) <= not(layer6_outputs(1132));
    outputs(1237) <= not((layer6_outputs(485)) and (layer6_outputs(658)));
    outputs(1238) <= not(layer6_outputs(15));
    outputs(1239) <= (layer6_outputs(2218)) xor (layer6_outputs(1006));
    outputs(1240) <= not(layer6_outputs(2557));
    outputs(1241) <= (layer6_outputs(772)) xor (layer6_outputs(1671));
    outputs(1242) <= layer6_outputs(1908);
    outputs(1243) <= not(layer6_outputs(2091));
    outputs(1244) <= not(layer6_outputs(12));
    outputs(1245) <= layer6_outputs(1344);
    outputs(1246) <= layer6_outputs(288);
    outputs(1247) <= not(layer6_outputs(1763));
    outputs(1248) <= not(layer6_outputs(641));
    outputs(1249) <= layer6_outputs(1972);
    outputs(1250) <= layer6_outputs(1483);
    outputs(1251) <= layer6_outputs(2537);
    outputs(1252) <= layer6_outputs(2468);
    outputs(1253) <= not(layer6_outputs(443));
    outputs(1254) <= not((layer6_outputs(1077)) or (layer6_outputs(110)));
    outputs(1255) <= (layer6_outputs(1893)) and not (layer6_outputs(931));
    outputs(1256) <= not(layer6_outputs(1663));
    outputs(1257) <= (layer6_outputs(2244)) and not (layer6_outputs(2433));
    outputs(1258) <= (layer6_outputs(74)) and (layer6_outputs(2254));
    outputs(1259) <= not((layer6_outputs(573)) xor (layer6_outputs(849)));
    outputs(1260) <= not(layer6_outputs(468));
    outputs(1261) <= not(layer6_outputs(647));
    outputs(1262) <= not(layer6_outputs(183));
    outputs(1263) <= not((layer6_outputs(500)) and (layer6_outputs(1530)));
    outputs(1264) <= layer6_outputs(1575);
    outputs(1265) <= not(layer6_outputs(1379));
    outputs(1266) <= not(layer6_outputs(333));
    outputs(1267) <= not(layer6_outputs(2168));
    outputs(1268) <= layer6_outputs(1887);
    outputs(1269) <= not(layer6_outputs(1162));
    outputs(1270) <= layer6_outputs(566);
    outputs(1271) <= not(layer6_outputs(2465));
    outputs(1272) <= layer6_outputs(1907);
    outputs(1273) <= layer6_outputs(1370);
    outputs(1274) <= not(layer6_outputs(2088));
    outputs(1275) <= not(layer6_outputs(1336));
    outputs(1276) <= not(layer6_outputs(2470));
    outputs(1277) <= (layer6_outputs(80)) and (layer6_outputs(552));
    outputs(1278) <= (layer6_outputs(611)) xor (layer6_outputs(63));
    outputs(1279) <= not(layer6_outputs(250));
    outputs(1280) <= layer6_outputs(756);
    outputs(1281) <= not(layer6_outputs(420));
    outputs(1282) <= layer6_outputs(1116);
    outputs(1283) <= layer6_outputs(2368);
    outputs(1284) <= not((layer6_outputs(243)) or (layer6_outputs(2129)));
    outputs(1285) <= (layer6_outputs(1300)) xor (layer6_outputs(239));
    outputs(1286) <= (layer6_outputs(1180)) xor (layer6_outputs(1250));
    outputs(1287) <= not((layer6_outputs(109)) and (layer6_outputs(839)));
    outputs(1288) <= (layer6_outputs(1918)) xor (layer6_outputs(2214));
    outputs(1289) <= not(layer6_outputs(347));
    outputs(1290) <= layer6_outputs(752);
    outputs(1291) <= not(layer6_outputs(82)) or (layer6_outputs(245));
    outputs(1292) <= (layer6_outputs(152)) and not (layer6_outputs(2137));
    outputs(1293) <= (layer6_outputs(62)) xor (layer6_outputs(2045));
    outputs(1294) <= not(layer6_outputs(1699));
    outputs(1295) <= not((layer6_outputs(1571)) and (layer6_outputs(1860)));
    outputs(1296) <= not(layer6_outputs(662));
    outputs(1297) <= layer6_outputs(1516);
    outputs(1298) <= layer6_outputs(2525);
    outputs(1299) <= not(layer6_outputs(2458));
    outputs(1300) <= layer6_outputs(1963);
    outputs(1301) <= layer6_outputs(1937);
    outputs(1302) <= (layer6_outputs(927)) and not (layer6_outputs(2366));
    outputs(1303) <= not(layer6_outputs(689));
    outputs(1304) <= (layer6_outputs(1454)) xor (layer6_outputs(1888));
    outputs(1305) <= not((layer6_outputs(1920)) xor (layer6_outputs(1177)));
    outputs(1306) <= layer6_outputs(2338);
    outputs(1307) <= layer6_outputs(471);
    outputs(1308) <= not(layer6_outputs(1334));
    outputs(1309) <= layer6_outputs(1031);
    outputs(1310) <= not(layer6_outputs(269));
    outputs(1311) <= not(layer6_outputs(1833));
    outputs(1312) <= (layer6_outputs(737)) xor (layer6_outputs(1581));
    outputs(1313) <= layer6_outputs(1164);
    outputs(1314) <= not(layer6_outputs(1640));
    outputs(1315) <= not(layer6_outputs(707));
    outputs(1316) <= not((layer6_outputs(1222)) xor (layer6_outputs(1923)));
    outputs(1317) <= (layer6_outputs(2431)) xor (layer6_outputs(741));
    outputs(1318) <= not((layer6_outputs(1044)) xor (layer6_outputs(526)));
    outputs(1319) <= not((layer6_outputs(260)) xor (layer6_outputs(184)));
    outputs(1320) <= layer6_outputs(682);
    outputs(1321) <= layer6_outputs(576);
    outputs(1322) <= (layer6_outputs(1542)) and not (layer6_outputs(2092));
    outputs(1323) <= (layer6_outputs(1822)) xor (layer6_outputs(1285));
    outputs(1324) <= layer6_outputs(1643);
    outputs(1325) <= not(layer6_outputs(2110));
    outputs(1326) <= not(layer6_outputs(1366));
    outputs(1327) <= layer6_outputs(1714);
    outputs(1328) <= not(layer6_outputs(1733));
    outputs(1329) <= layer6_outputs(608);
    outputs(1330) <= not((layer6_outputs(842)) and (layer6_outputs(1784)));
    outputs(1331) <= layer6_outputs(493);
    outputs(1332) <= not((layer6_outputs(1771)) or (layer6_outputs(553)));
    outputs(1333) <= (layer6_outputs(1881)) xor (layer6_outputs(1400));
    outputs(1334) <= not((layer6_outputs(1827)) or (layer6_outputs(2520)));
    outputs(1335) <= not((layer6_outputs(1396)) xor (layer6_outputs(1536)));
    outputs(1336) <= not(layer6_outputs(2051));
    outputs(1337) <= not(layer6_outputs(2238));
    outputs(1338) <= not(layer6_outputs(1703));
    outputs(1339) <= not(layer6_outputs(1524));
    outputs(1340) <= layer6_outputs(2114);
    outputs(1341) <= (layer6_outputs(1342)) or (layer6_outputs(2239));
    outputs(1342) <= not((layer6_outputs(1052)) xor (layer6_outputs(1642)));
    outputs(1343) <= (layer6_outputs(976)) and not (layer6_outputs(1718));
    outputs(1344) <= layer6_outputs(677);
    outputs(1345) <= not((layer6_outputs(2000)) xor (layer6_outputs(1496)));
    outputs(1346) <= not((layer6_outputs(1221)) xor (layer6_outputs(2306)));
    outputs(1347) <= layer6_outputs(508);
    outputs(1348) <= (layer6_outputs(1187)) and not (layer6_outputs(626));
    outputs(1349) <= (layer6_outputs(1821)) xor (layer6_outputs(2277));
    outputs(1350) <= not((layer6_outputs(1340)) or (layer6_outputs(1241)));
    outputs(1351) <= layer6_outputs(1752);
    outputs(1352) <= not(layer6_outputs(1313));
    outputs(1353) <= layer6_outputs(1383);
    outputs(1354) <= (layer6_outputs(1001)) xor (layer6_outputs(115));
    outputs(1355) <= (layer6_outputs(1759)) xor (layer6_outputs(2535));
    outputs(1356) <= (layer6_outputs(10)) xor (layer6_outputs(1580));
    outputs(1357) <= layer6_outputs(802);
    outputs(1358) <= not((layer6_outputs(1118)) or (layer6_outputs(2047)));
    outputs(1359) <= layer6_outputs(2144);
    outputs(1360) <= not((layer6_outputs(2378)) xor (layer6_outputs(2251)));
    outputs(1361) <= (layer6_outputs(416)) and not (layer6_outputs(2064));
    outputs(1362) <= (layer6_outputs(2379)) xor (layer6_outputs(1724));
    outputs(1363) <= not(layer6_outputs(449));
    outputs(1364) <= not(layer6_outputs(2177));
    outputs(1365) <= layer6_outputs(1326);
    outputs(1366) <= layer6_outputs(1495);
    outputs(1367) <= (layer6_outputs(38)) or (layer6_outputs(992));
    outputs(1368) <= not((layer6_outputs(710)) or (layer6_outputs(2291)));
    outputs(1369) <= layer6_outputs(831);
    outputs(1370) <= layer6_outputs(750);
    outputs(1371) <= not(layer6_outputs(1095));
    outputs(1372) <= (layer6_outputs(776)) xor (layer6_outputs(2426));
    outputs(1373) <= not(layer6_outputs(2410));
    outputs(1374) <= not((layer6_outputs(1890)) xor (layer6_outputs(1283)));
    outputs(1375) <= not((layer6_outputs(1329)) and (layer6_outputs(441)));
    outputs(1376) <= not((layer6_outputs(2259)) xor (layer6_outputs(479)));
    outputs(1377) <= not(layer6_outputs(1502)) or (layer6_outputs(1194));
    outputs(1378) <= layer6_outputs(1414);
    outputs(1379) <= layer6_outputs(282);
    outputs(1380) <= not(layer6_outputs(469));
    outputs(1381) <= not(layer6_outputs(1712));
    outputs(1382) <= (layer6_outputs(571)) xor (layer6_outputs(591));
    outputs(1383) <= (layer6_outputs(667)) xor (layer6_outputs(1453));
    outputs(1384) <= (layer6_outputs(609)) and not (layer6_outputs(2548));
    outputs(1385) <= layer6_outputs(2258);
    outputs(1386) <= layer6_outputs(2223);
    outputs(1387) <= layer6_outputs(1251);
    outputs(1388) <= not((layer6_outputs(816)) xor (layer6_outputs(832)));
    outputs(1389) <= not(layer6_outputs(139)) or (layer6_outputs(659));
    outputs(1390) <= not(layer6_outputs(1400));
    outputs(1391) <= layer6_outputs(2100);
    outputs(1392) <= (layer6_outputs(473)) and not (layer6_outputs(1485));
    outputs(1393) <= layer6_outputs(1813);
    outputs(1394) <= (layer6_outputs(1315)) xor (layer6_outputs(1025));
    outputs(1395) <= layer6_outputs(1949);
    outputs(1396) <= not(layer6_outputs(691));
    outputs(1397) <= not(layer6_outputs(2422));
    outputs(1398) <= not(layer6_outputs(1437)) or (layer6_outputs(2215));
    outputs(1399) <= not(layer6_outputs(1928)) or (layer6_outputs(2331));
    outputs(1400) <= not((layer6_outputs(352)) xor (layer6_outputs(324)));
    outputs(1401) <= not(layer6_outputs(1173)) or (layer6_outputs(893));
    outputs(1402) <= not(layer6_outputs(842));
    outputs(1403) <= (layer6_outputs(266)) and not (layer6_outputs(1223));
    outputs(1404) <= not(layer6_outputs(487));
    outputs(1405) <= not((layer6_outputs(940)) or (layer6_outputs(2473)));
    outputs(1406) <= not(layer6_outputs(431));
    outputs(1407) <= (layer6_outputs(1863)) and (layer6_outputs(1240));
    outputs(1408) <= layer6_outputs(1087);
    outputs(1409) <= not(layer6_outputs(692));
    outputs(1410) <= not(layer6_outputs(2409));
    outputs(1411) <= not(layer6_outputs(1046));
    outputs(1412) <= (layer6_outputs(766)) and not (layer6_outputs(163));
    outputs(1413) <= not((layer6_outputs(1565)) xor (layer6_outputs(1177)));
    outputs(1414) <= layer6_outputs(751);
    outputs(1415) <= (layer6_outputs(0)) xor (layer6_outputs(848));
    outputs(1416) <= layer6_outputs(1184);
    outputs(1417) <= (layer6_outputs(1827)) xor (layer6_outputs(1619));
    outputs(1418) <= not(layer6_outputs(635));
    outputs(1419) <= not((layer6_outputs(118)) or (layer6_outputs(1541)));
    outputs(1420) <= layer6_outputs(2260);
    outputs(1421) <= (layer6_outputs(1062)) and not (layer6_outputs(1254));
    outputs(1422) <= (layer6_outputs(1469)) xor (layer6_outputs(1373));
    outputs(1423) <= (layer6_outputs(2112)) xor (layer6_outputs(295));
    outputs(1424) <= not(layer6_outputs(1357));
    outputs(1425) <= layer6_outputs(1163);
    outputs(1426) <= not(layer6_outputs(1692));
    outputs(1427) <= layer6_outputs(1050);
    outputs(1428) <= layer6_outputs(1464);
    outputs(1429) <= (layer6_outputs(1871)) and (layer6_outputs(1004));
    outputs(1430) <= layer6_outputs(771);
    outputs(1431) <= layer6_outputs(2065);
    outputs(1432) <= layer6_outputs(1622);
    outputs(1433) <= (layer6_outputs(2297)) xor (layer6_outputs(2465));
    outputs(1434) <= layer6_outputs(180);
    outputs(1435) <= (layer6_outputs(1816)) xor (layer6_outputs(2397));
    outputs(1436) <= not((layer6_outputs(1782)) xor (layer6_outputs(1355)));
    outputs(1437) <= not((layer6_outputs(1138)) xor (layer6_outputs(2462)));
    outputs(1438) <= (layer6_outputs(183)) xor (layer6_outputs(2372));
    outputs(1439) <= layer6_outputs(555);
    outputs(1440) <= not(layer6_outputs(770));
    outputs(1441) <= not((layer6_outputs(111)) xor (layer6_outputs(2165)));
    outputs(1442) <= not((layer6_outputs(1875)) xor (layer6_outputs(1820)));
    outputs(1443) <= layer6_outputs(206);
    outputs(1444) <= layer6_outputs(2009);
    outputs(1445) <= (layer6_outputs(412)) xor (layer6_outputs(1741));
    outputs(1446) <= not((layer6_outputs(699)) xor (layer6_outputs(909)));
    outputs(1447) <= (layer6_outputs(1192)) xor (layer6_outputs(867));
    outputs(1448) <= layer6_outputs(231);
    outputs(1449) <= not(layer6_outputs(1792));
    outputs(1450) <= (layer6_outputs(1545)) xor (layer6_outputs(2128));
    outputs(1451) <= (layer6_outputs(386)) and not (layer6_outputs(2348));
    outputs(1452) <= layer6_outputs(333);
    outputs(1453) <= layer6_outputs(559);
    outputs(1454) <= not(layer6_outputs(1927));
    outputs(1455) <= not((layer6_outputs(1605)) and (layer6_outputs(937)));
    outputs(1456) <= layer6_outputs(373);
    outputs(1457) <= not(layer6_outputs(1578));
    outputs(1458) <= not((layer6_outputs(1824)) xor (layer6_outputs(2146)));
    outputs(1459) <= not(layer6_outputs(2470));
    outputs(1460) <= not((layer6_outputs(815)) xor (layer6_outputs(1610)));
    outputs(1461) <= not(layer6_outputs(1513));
    outputs(1462) <= (layer6_outputs(48)) and not (layer6_outputs(1665));
    outputs(1463) <= not((layer6_outputs(1711)) or (layer6_outputs(1984)));
    outputs(1464) <= not(layer6_outputs(1723));
    outputs(1465) <= not(layer6_outputs(691));
    outputs(1466) <= not((layer6_outputs(1989)) xor (layer6_outputs(2084)));
    outputs(1467) <= (layer6_outputs(215)) xor (layer6_outputs(2526));
    outputs(1468) <= layer6_outputs(2365);
    outputs(1469) <= (layer6_outputs(1170)) xor (layer6_outputs(742));
    outputs(1470) <= layer6_outputs(1444);
    outputs(1471) <= layer6_outputs(2193);
    outputs(1472) <= not(layer6_outputs(1488));
    outputs(1473) <= not(layer6_outputs(1780));
    outputs(1474) <= layer6_outputs(645);
    outputs(1475) <= not(layer6_outputs(487));
    outputs(1476) <= not(layer6_outputs(1347));
    outputs(1477) <= not(layer6_outputs(2448));
    outputs(1478) <= not((layer6_outputs(2048)) xor (layer6_outputs(939)));
    outputs(1479) <= layer6_outputs(219);
    outputs(1480) <= layer6_outputs(1878);
    outputs(1481) <= layer6_outputs(278);
    outputs(1482) <= layer6_outputs(194);
    outputs(1483) <= not(layer6_outputs(2173)) or (layer6_outputs(1954));
    outputs(1484) <= not((layer6_outputs(1739)) xor (layer6_outputs(1896)));
    outputs(1485) <= layer6_outputs(326);
    outputs(1486) <= not(layer6_outputs(314));
    outputs(1487) <= not((layer6_outputs(1751)) xor (layer6_outputs(87)));
    outputs(1488) <= not(layer6_outputs(661));
    outputs(1489) <= not(layer6_outputs(2273));
    outputs(1490) <= not(layer6_outputs(1392));
    outputs(1491) <= layer6_outputs(453);
    outputs(1492) <= not(layer6_outputs(1794));
    outputs(1493) <= layer6_outputs(2506);
    outputs(1494) <= layer6_outputs(2018);
    outputs(1495) <= (layer6_outputs(1759)) and not (layer6_outputs(1018));
    outputs(1496) <= (layer6_outputs(2432)) xor (layer6_outputs(2132));
    outputs(1497) <= (layer6_outputs(1257)) xor (layer6_outputs(1212));
    outputs(1498) <= layer6_outputs(336);
    outputs(1499) <= not(layer6_outputs(1733));
    outputs(1500) <= not((layer6_outputs(579)) xor (layer6_outputs(928)));
    outputs(1501) <= not(layer6_outputs(1510));
    outputs(1502) <= layer6_outputs(1151);
    outputs(1503) <= layer6_outputs(2105);
    outputs(1504) <= not((layer6_outputs(1942)) xor (layer6_outputs(1632)));
    outputs(1505) <= layer6_outputs(763);
    outputs(1506) <= layer6_outputs(1609);
    outputs(1507) <= (layer6_outputs(1758)) xor (layer6_outputs(969));
    outputs(1508) <= not(layer6_outputs(205));
    outputs(1509) <= layer6_outputs(1015);
    outputs(1510) <= not((layer6_outputs(961)) xor (layer6_outputs(1769)));
    outputs(1511) <= not((layer6_outputs(1205)) xor (layer6_outputs(1142)));
    outputs(1512) <= layer6_outputs(653);
    outputs(1513) <= layer6_outputs(1297);
    outputs(1514) <= not(layer6_outputs(492));
    outputs(1515) <= (layer6_outputs(1981)) xor (layer6_outputs(2240));
    outputs(1516) <= (layer6_outputs(2498)) xor (layer6_outputs(1010));
    outputs(1517) <= (layer6_outputs(1338)) xor (layer6_outputs(1953));
    outputs(1518) <= not((layer6_outputs(1305)) xor (layer6_outputs(2130)));
    outputs(1519) <= (layer6_outputs(1793)) xor (layer6_outputs(1338));
    outputs(1520) <= not((layer6_outputs(664)) xor (layer6_outputs(2556)));
    outputs(1521) <= layer6_outputs(345);
    outputs(1522) <= not(layer6_outputs(635));
    outputs(1523) <= layer6_outputs(829);
    outputs(1524) <= layer6_outputs(2061);
    outputs(1525) <= not((layer6_outputs(746)) xor (layer6_outputs(2543)));
    outputs(1526) <= not(layer6_outputs(1258));
    outputs(1527) <= layer6_outputs(1841);
    outputs(1528) <= (layer6_outputs(125)) or (layer6_outputs(2119));
    outputs(1529) <= not(layer6_outputs(331));
    outputs(1530) <= layer6_outputs(676);
    outputs(1531) <= not((layer6_outputs(721)) xor (layer6_outputs(1069)));
    outputs(1532) <= not(layer6_outputs(214));
    outputs(1533) <= not(layer6_outputs(2421));
    outputs(1534) <= layer6_outputs(1566);
    outputs(1535) <= not(layer6_outputs(370));
    outputs(1536) <= layer6_outputs(1183);
    outputs(1537) <= layer6_outputs(1505);
    outputs(1538) <= layer6_outputs(1648);
    outputs(1539) <= layer6_outputs(1550);
    outputs(1540) <= layer6_outputs(2023);
    outputs(1541) <= not(layer6_outputs(1014));
    outputs(1542) <= not(layer6_outputs(196));
    outputs(1543) <= not(layer6_outputs(1877));
    outputs(1544) <= not(layer6_outputs(2313));
    outputs(1545) <= not(layer6_outputs(774));
    outputs(1546) <= not((layer6_outputs(13)) and (layer6_outputs(98)));
    outputs(1547) <= not((layer6_outputs(2117)) xor (layer6_outputs(2289)));
    outputs(1548) <= (layer6_outputs(1862)) and (layer6_outputs(2183));
    outputs(1549) <= (layer6_outputs(978)) xor (layer6_outputs(670));
    outputs(1550) <= not(layer6_outputs(119));
    outputs(1551) <= not((layer6_outputs(713)) xor (layer6_outputs(614)));
    outputs(1552) <= not(layer6_outputs(2317));
    outputs(1553) <= layer6_outputs(541);
    outputs(1554) <= layer6_outputs(1904);
    outputs(1555) <= layer6_outputs(49);
    outputs(1556) <= (layer6_outputs(754)) xor (layer6_outputs(1560));
    outputs(1557) <= not((layer6_outputs(788)) xor (layer6_outputs(951)));
    outputs(1558) <= not(layer6_outputs(152));
    outputs(1559) <= not(layer6_outputs(358));
    outputs(1560) <= not(layer6_outputs(1865));
    outputs(1561) <= layer6_outputs(2014);
    outputs(1562) <= (layer6_outputs(1647)) xor (layer6_outputs(1886));
    outputs(1563) <= not(layer6_outputs(874));
    outputs(1564) <= layer6_outputs(1883);
    outputs(1565) <= (layer6_outputs(1092)) xor (layer6_outputs(775));
    outputs(1566) <= layer6_outputs(2369);
    outputs(1567) <= layer6_outputs(1404);
    outputs(1568) <= not((layer6_outputs(1426)) xor (layer6_outputs(1922)));
    outputs(1569) <= not(layer6_outputs(2359));
    outputs(1570) <= not(layer6_outputs(476));
    outputs(1571) <= (layer6_outputs(2384)) and not (layer6_outputs(2459));
    outputs(1572) <= (layer6_outputs(1146)) and (layer6_outputs(669));
    outputs(1573) <= not((layer6_outputs(1572)) and (layer6_outputs(767)));
    outputs(1574) <= layer6_outputs(582);
    outputs(1575) <= not((layer6_outputs(570)) xor (layer6_outputs(1455)));
    outputs(1576) <= not(layer6_outputs(540)) or (layer6_outputs(1344));
    outputs(1577) <= not(layer6_outputs(2264));
    outputs(1578) <= not(layer6_outputs(1838));
    outputs(1579) <= layer6_outputs(840);
    outputs(1580) <= layer6_outputs(1552);
    outputs(1581) <= not((layer6_outputs(524)) or (layer6_outputs(858)));
    outputs(1582) <= not(layer6_outputs(110));
    outputs(1583) <= (layer6_outputs(1564)) xor (layer6_outputs(657));
    outputs(1584) <= (layer6_outputs(1189)) xor (layer6_outputs(2419));
    outputs(1585) <= (layer6_outputs(1391)) xor (layer6_outputs(2288));
    outputs(1586) <= (layer6_outputs(2311)) xor (layer6_outputs(535));
    outputs(1587) <= not(layer6_outputs(244));
    outputs(1588) <= not((layer6_outputs(1541)) xor (layer6_outputs(1054)));
    outputs(1589) <= (layer6_outputs(1413)) and (layer6_outputs(68));
    outputs(1590) <= layer6_outputs(1833);
    outputs(1591) <= layer6_outputs(1905);
    outputs(1592) <= layer6_outputs(2043);
    outputs(1593) <= not((layer6_outputs(2180)) xor (layer6_outputs(1149)));
    outputs(1594) <= layer6_outputs(1684);
    outputs(1595) <= not(layer6_outputs(598));
    outputs(1596) <= layer6_outputs(2414);
    outputs(1597) <= not((layer6_outputs(922)) xor (layer6_outputs(646)));
    outputs(1598) <= (layer6_outputs(986)) xor (layer6_outputs(1406));
    outputs(1599) <= layer6_outputs(2280);
    outputs(1600) <= not(layer6_outputs(1669));
    outputs(1601) <= not(layer6_outputs(436));
    outputs(1602) <= not(layer6_outputs(1308));
    outputs(1603) <= not(layer6_outputs(1914));
    outputs(1604) <= (layer6_outputs(1539)) and not (layer6_outputs(896));
    outputs(1605) <= (layer6_outputs(124)) xor (layer6_outputs(4));
    outputs(1606) <= layer6_outputs(1297);
    outputs(1607) <= not((layer6_outputs(778)) or (layer6_outputs(2294)));
    outputs(1608) <= not(layer6_outputs(2490)) or (layer6_outputs(1632));
    outputs(1609) <= layer6_outputs(2243);
    outputs(1610) <= not(layer6_outputs(1650));
    outputs(1611) <= layer6_outputs(112);
    outputs(1612) <= not((layer6_outputs(1075)) and (layer6_outputs(2512)));
    outputs(1613) <= not(layer6_outputs(1354));
    outputs(1614) <= not((layer6_outputs(599)) or (layer6_outputs(2415)));
    outputs(1615) <= not(layer6_outputs(857));
    outputs(1616) <= not((layer6_outputs(769)) and (layer6_outputs(1662)));
    outputs(1617) <= (layer6_outputs(1027)) xor (layer6_outputs(1834));
    outputs(1618) <= not((layer6_outputs(1798)) or (layer6_outputs(199)));
    outputs(1619) <= (layer6_outputs(1160)) xor (layer6_outputs(1604));
    outputs(1620) <= layer6_outputs(2417);
    outputs(1621) <= layer6_outputs(1539);
    outputs(1622) <= not((layer6_outputs(1470)) or (layer6_outputs(1474)));
    outputs(1623) <= layer6_outputs(2401);
    outputs(1624) <= not(layer6_outputs(308));
    outputs(1625) <= not((layer6_outputs(1748)) and (layer6_outputs(1306)));
    outputs(1626) <= not((layer6_outputs(1638)) or (layer6_outputs(1167)));
    outputs(1627) <= not(layer6_outputs(1131));
    outputs(1628) <= layer6_outputs(124);
    outputs(1629) <= not(layer6_outputs(639));
    outputs(1630) <= not(layer6_outputs(319));
    outputs(1631) <= not((layer6_outputs(793)) or (layer6_outputs(1058)));
    outputs(1632) <= (layer6_outputs(1001)) and (layer6_outputs(371));
    outputs(1633) <= layer6_outputs(1716);
    outputs(1634) <= not(layer6_outputs(379));
    outputs(1635) <= not((layer6_outputs(590)) xor (layer6_outputs(2404)));
    outputs(1636) <= layer6_outputs(614);
    outputs(1637) <= (layer6_outputs(1437)) and not (layer6_outputs(1377));
    outputs(1638) <= (layer6_outputs(651)) and (layer6_outputs(2133));
    outputs(1639) <= layer6_outputs(906);
    outputs(1640) <= layer6_outputs(2232);
    outputs(1641) <= not(layer6_outputs(1090));
    outputs(1642) <= layer6_outputs(1239);
    outputs(1643) <= not((layer6_outputs(489)) or (layer6_outputs(1663)));
    outputs(1644) <= not((layer6_outputs(900)) and (layer6_outputs(2083)));
    outputs(1645) <= layer6_outputs(242);
    outputs(1646) <= not(layer6_outputs(187));
    outputs(1647) <= (layer6_outputs(2275)) and (layer6_outputs(1637));
    outputs(1648) <= not(layer6_outputs(1913));
    outputs(1649) <= not(layer6_outputs(2526));
    outputs(1650) <= not(layer6_outputs(1498));
    outputs(1651) <= not((layer6_outputs(551)) xor (layer6_outputs(727)));
    outputs(1652) <= layer6_outputs(582);
    outputs(1653) <= not((layer6_outputs(979)) xor (layer6_outputs(1399)));
    outputs(1654) <= layer6_outputs(2234);
    outputs(1655) <= layer6_outputs(1387);
    outputs(1656) <= (layer6_outputs(1263)) xor (layer6_outputs(869));
    outputs(1657) <= layer6_outputs(2248);
    outputs(1658) <= layer6_outputs(1832);
    outputs(1659) <= not(layer6_outputs(1615));
    outputs(1660) <= not((layer6_outputs(441)) or (layer6_outputs(2550)));
    outputs(1661) <= not((layer6_outputs(591)) xor (layer6_outputs(2513)));
    outputs(1662) <= (layer6_outputs(1186)) and not (layer6_outputs(1382));
    outputs(1663) <= (layer6_outputs(1316)) and (layer6_outputs(2476));
    outputs(1664) <= layer6_outputs(906);
    outputs(1665) <= (layer6_outputs(142)) xor (layer6_outputs(947));
    outputs(1666) <= not(layer6_outputs(1275));
    outputs(1667) <= layer6_outputs(1432);
    outputs(1668) <= (layer6_outputs(804)) xor (layer6_outputs(1873));
    outputs(1669) <= not(layer6_outputs(2261));
    outputs(1670) <= (layer6_outputs(2541)) xor (layer6_outputs(2370));
    outputs(1671) <= not(layer6_outputs(1636));
    outputs(1672) <= (layer6_outputs(2207)) xor (layer6_outputs(45));
    outputs(1673) <= not(layer6_outputs(1729));
    outputs(1674) <= layer6_outputs(138);
    outputs(1675) <= not(layer6_outputs(134));
    outputs(1676) <= (layer6_outputs(1911)) and (layer6_outputs(965));
    outputs(1677) <= not(layer6_outputs(2108));
    outputs(1678) <= not(layer6_outputs(1488));
    outputs(1679) <= layer6_outputs(2321);
    outputs(1680) <= (layer6_outputs(1174)) and not (layer6_outputs(1198));
    outputs(1681) <= layer6_outputs(221);
    outputs(1682) <= not(layer6_outputs(1089));
    outputs(1683) <= not((layer6_outputs(1848)) xor (layer6_outputs(1090)));
    outputs(1684) <= layer6_outputs(669);
    outputs(1685) <= not(layer6_outputs(2087));
    outputs(1686) <= (layer6_outputs(429)) and not (layer6_outputs(953));
    outputs(1687) <= not(layer6_outputs(2451));
    outputs(1688) <= (layer6_outputs(228)) and (layer6_outputs(594));
    outputs(1689) <= not((layer6_outputs(311)) xor (layer6_outputs(1202)));
    outputs(1690) <= layer6_outputs(646);
    outputs(1691) <= not(layer6_outputs(2108));
    outputs(1692) <= not(layer6_outputs(2494));
    outputs(1693) <= not(layer6_outputs(18));
    outputs(1694) <= layer6_outputs(534);
    outputs(1695) <= (layer6_outputs(2042)) and not (layer6_outputs(2029));
    outputs(1696) <= not((layer6_outputs(703)) xor (layer6_outputs(2387)));
    outputs(1697) <= (layer6_outputs(2005)) or (layer6_outputs(1474));
    outputs(1698) <= layer6_outputs(491);
    outputs(1699) <= layer6_outputs(1691);
    outputs(1700) <= layer6_outputs(2315);
    outputs(1701) <= (layer6_outputs(2393)) and not (layer6_outputs(1366));
    outputs(1702) <= (layer6_outputs(733)) xor (layer6_outputs(900));
    outputs(1703) <= (layer6_outputs(1725)) xor (layer6_outputs(915));
    outputs(1704) <= not(layer6_outputs(372));
    outputs(1705) <= not(layer6_outputs(563));
    outputs(1706) <= not((layer6_outputs(1040)) xor (layer6_outputs(1456)));
    outputs(1707) <= not(layer6_outputs(1487));
    outputs(1708) <= layer6_outputs(1186);
    outputs(1709) <= layer6_outputs(1203);
    outputs(1710) <= not(layer6_outputs(1762));
    outputs(1711) <= not(layer6_outputs(1284)) or (layer6_outputs(1693));
    outputs(1712) <= layer6_outputs(722);
    outputs(1713) <= not(layer6_outputs(126));
    outputs(1714) <= layer6_outputs(2416);
    outputs(1715) <= (layer6_outputs(276)) xor (layer6_outputs(1702));
    outputs(1716) <= (layer6_outputs(2315)) and not (layer6_outputs(2273));
    outputs(1717) <= not((layer6_outputs(792)) xor (layer6_outputs(608)));
    outputs(1718) <= layer6_outputs(246);
    outputs(1719) <= (layer6_outputs(748)) xor (layer6_outputs(142));
    outputs(1720) <= not(layer6_outputs(1236));
    outputs(1721) <= layer6_outputs(2344);
    outputs(1722) <= not((layer6_outputs(1486)) xor (layer6_outputs(726)));
    outputs(1723) <= not(layer6_outputs(2182));
    outputs(1724) <= (layer6_outputs(1628)) xor (layer6_outputs(1707));
    outputs(1725) <= (layer6_outputs(237)) and (layer6_outputs(207));
    outputs(1726) <= not(layer6_outputs(248));
    outputs(1727) <= (layer6_outputs(1084)) or (layer6_outputs(1446));
    outputs(1728) <= (layer6_outputs(456)) and (layer6_outputs(34));
    outputs(1729) <= (layer6_outputs(1543)) xor (layer6_outputs(1053));
    outputs(1730) <= layer6_outputs(829);
    outputs(1731) <= not((layer6_outputs(128)) and (layer6_outputs(1097)));
    outputs(1732) <= (layer6_outputs(786)) and (layer6_outputs(1727));
    outputs(1733) <= (layer6_outputs(318)) and (layer6_outputs(1196));
    outputs(1734) <= layer6_outputs(879);
    outputs(1735) <= layer6_outputs(741);
    outputs(1736) <= not((layer6_outputs(634)) xor (layer6_outputs(1075)));
    outputs(1737) <= layer6_outputs(1529);
    outputs(1738) <= layer6_outputs(114);
    outputs(1739) <= not(layer6_outputs(581));
    outputs(1740) <= (layer6_outputs(2103)) and not (layer6_outputs(259));
    outputs(1741) <= not(layer6_outputs(1831));
    outputs(1742) <= layer6_outputs(1617);
    outputs(1743) <= (layer6_outputs(1879)) and not (layer6_outputs(117));
    outputs(1744) <= not(layer6_outputs(683)) or (layer6_outputs(1248));
    outputs(1745) <= (layer6_outputs(743)) and not (layer6_outputs(2300));
    outputs(1746) <= (layer6_outputs(2290)) and not (layer6_outputs(211));
    outputs(1747) <= not(layer6_outputs(1430));
    outputs(1748) <= layer6_outputs(2402);
    outputs(1749) <= not(layer6_outputs(26));
    outputs(1750) <= (layer6_outputs(977)) xor (layer6_outputs(1842));
    outputs(1751) <= not(layer6_outputs(134));
    outputs(1752) <= layer6_outputs(1270);
    outputs(1753) <= (layer6_outputs(261)) xor (layer6_outputs(1458));
    outputs(1754) <= (layer6_outputs(1652)) and not (layer6_outputs(734));
    outputs(1755) <= not(layer6_outputs(984));
    outputs(1756) <= layer6_outputs(2138);
    outputs(1757) <= layer6_outputs(457);
    outputs(1758) <= not((layer6_outputs(851)) xor (layer6_outputs(153)));
    outputs(1759) <= (layer6_outputs(1349)) and not (layer6_outputs(279));
    outputs(1760) <= layer6_outputs(2036);
    outputs(1761) <= not(layer6_outputs(2179));
    outputs(1762) <= not(layer6_outputs(2265));
    outputs(1763) <= (layer6_outputs(2351)) xor (layer6_outputs(1591));
    outputs(1764) <= not(layer6_outputs(1285)) or (layer6_outputs(1852));
    outputs(1765) <= not(layer6_outputs(1675));
    outputs(1766) <= layer6_outputs(2115);
    outputs(1767) <= layer6_outputs(952);
    outputs(1768) <= layer6_outputs(1253);
    outputs(1769) <= not(layer6_outputs(1132));
    outputs(1770) <= not(layer6_outputs(2162));
    outputs(1771) <= not(layer6_outputs(2546));
    outputs(1772) <= not(layer6_outputs(1869));
    outputs(1773) <= not(layer6_outputs(484));
    outputs(1774) <= not(layer6_outputs(2096));
    outputs(1775) <= layer6_outputs(596);
    outputs(1776) <= layer6_outputs(2);
    outputs(1777) <= layer6_outputs(946);
    outputs(1778) <= not(layer6_outputs(1421));
    outputs(1779) <= not((layer6_outputs(754)) xor (layer6_outputs(872)));
    outputs(1780) <= not((layer6_outputs(1881)) xor (layer6_outputs(1505)));
    outputs(1781) <= layer6_outputs(300);
    outputs(1782) <= layer6_outputs(412);
    outputs(1783) <= not(layer6_outputs(1130));
    outputs(1784) <= not(layer6_outputs(510));
    outputs(1785) <= not(layer6_outputs(960));
    outputs(1786) <= layer6_outputs(1974);
    outputs(1787) <= layer6_outputs(1696);
    outputs(1788) <= not(layer6_outputs(113));
    outputs(1789) <= not(layer6_outputs(1806));
    outputs(1790) <= layer6_outputs(157);
    outputs(1791) <= not((layer6_outputs(1836)) xor (layer6_outputs(2026)));
    outputs(1792) <= layer6_outputs(1783);
    outputs(1793) <= not(layer6_outputs(668));
    outputs(1794) <= layer6_outputs(1641);
    outputs(1795) <= (layer6_outputs(120)) and (layer6_outputs(1420));
    outputs(1796) <= (layer6_outputs(1563)) and (layer6_outputs(2466));
    outputs(1797) <= not(layer6_outputs(904));
    outputs(1798) <= layer6_outputs(777);
    outputs(1799) <= not((layer6_outputs(1935)) xor (layer6_outputs(212)));
    outputs(1800) <= layer6_outputs(2376);
    outputs(1801) <= not((layer6_outputs(2122)) and (layer6_outputs(54)));
    outputs(1802) <= (layer6_outputs(35)) and not (layer6_outputs(539));
    outputs(1803) <= (layer6_outputs(2226)) and not (layer6_outputs(870));
    outputs(1804) <= not((layer6_outputs(1146)) xor (layer6_outputs(1197)));
    outputs(1805) <= layer6_outputs(2032);
    outputs(1806) <= not((layer6_outputs(1017)) xor (layer6_outputs(84)));
    outputs(1807) <= not(layer6_outputs(1516));
    outputs(1808) <= not(layer6_outputs(1204));
    outputs(1809) <= not((layer6_outputs(1715)) xor (layer6_outputs(85)));
    outputs(1810) <= layer6_outputs(1171);
    outputs(1811) <= (layer6_outputs(1008)) xor (layer6_outputs(1846));
    outputs(1812) <= not(layer6_outputs(538));
    outputs(1813) <= not((layer6_outputs(157)) or (layer6_outputs(285)));
    outputs(1814) <= not((layer6_outputs(92)) xor (layer6_outputs(489)));
    outputs(1815) <= not(layer6_outputs(2396));
    outputs(1816) <= not(layer6_outputs(1255));
    outputs(1817) <= not(layer6_outputs(1853));
    outputs(1818) <= layer6_outputs(852);
    outputs(1819) <= not(layer6_outputs(511));
    outputs(1820) <= not(layer6_outputs(1973));
    outputs(1821) <= not(layer6_outputs(607));
    outputs(1822) <= (layer6_outputs(2002)) and not (layer6_outputs(998));
    outputs(1823) <= layer6_outputs(1440);
    outputs(1824) <= (layer6_outputs(2153)) and not (layer6_outputs(229));
    outputs(1825) <= (layer6_outputs(1665)) and (layer6_outputs(1927));
    outputs(1826) <= layer6_outputs(2500);
    outputs(1827) <= layer6_outputs(1838);
    outputs(1828) <= not((layer6_outputs(2042)) and (layer6_outputs(272)));
    outputs(1829) <= layer6_outputs(390);
    outputs(1830) <= not((layer6_outputs(177)) xor (layer6_outputs(617)));
    outputs(1831) <= (layer6_outputs(1002)) xor (layer6_outputs(158));
    outputs(1832) <= not((layer6_outputs(1943)) xor (layer6_outputs(1435)));
    outputs(1833) <= layer6_outputs(280);
    outputs(1834) <= not(layer6_outputs(1740));
    outputs(1835) <= layer6_outputs(464);
    outputs(1836) <= not(layer6_outputs(2335));
    outputs(1837) <= layer6_outputs(499);
    outputs(1838) <= not(layer6_outputs(1804));
    outputs(1839) <= not(layer6_outputs(899));
    outputs(1840) <= not(layer6_outputs(1335));
    outputs(1841) <= layer6_outputs(469);
    outputs(1842) <= (layer6_outputs(226)) and not (layer6_outputs(1917));
    outputs(1843) <= layer6_outputs(1765);
    outputs(1844) <= layer6_outputs(1597);
    outputs(1845) <= layer6_outputs(402);
    outputs(1846) <= not(layer6_outputs(132));
    outputs(1847) <= layer6_outputs(779);
    outputs(1848) <= not(layer6_outputs(1268));
    outputs(1849) <= layer6_outputs(125);
    outputs(1850) <= (layer6_outputs(918)) and not (layer6_outputs(2532));
    outputs(1851) <= layer6_outputs(1770);
    outputs(1852) <= layer6_outputs(2147);
    outputs(1853) <= not(layer6_outputs(1837));
    outputs(1854) <= layer6_outputs(1630);
    outputs(1855) <= (layer6_outputs(1640)) xor (layer6_outputs(1272));
    outputs(1856) <= layer6_outputs(26);
    outputs(1857) <= layer6_outputs(2353);
    outputs(1858) <= not((layer6_outputs(920)) xor (layer6_outputs(2511)));
    outputs(1859) <= not(layer6_outputs(1063));
    outputs(1860) <= layer6_outputs(968);
    outputs(1861) <= not(layer6_outputs(1728)) or (layer6_outputs(2142));
    outputs(1862) <= layer6_outputs(1777);
    outputs(1863) <= not(layer6_outputs(1659));
    outputs(1864) <= (layer6_outputs(2064)) and (layer6_outputs(632));
    outputs(1865) <= layer6_outputs(916);
    outputs(1866) <= not((layer6_outputs(1003)) xor (layer6_outputs(624)));
    outputs(1867) <= not((layer6_outputs(430)) or (layer6_outputs(1393)));
    outputs(1868) <= layer6_outputs(588);
    outputs(1869) <= (layer6_outputs(1900)) xor (layer6_outputs(795));
    outputs(1870) <= layer6_outputs(2534);
    outputs(1871) <= not(layer6_outputs(2365));
    outputs(1872) <= layer6_outputs(586);
    outputs(1873) <= layer6_outputs(1633);
    outputs(1874) <= (layer6_outputs(1305)) xor (layer6_outputs(1809));
    outputs(1875) <= not(layer6_outputs(1333));
    outputs(1876) <= layer6_outputs(2124);
    outputs(1877) <= not((layer6_outputs(613)) or (layer6_outputs(2139)));
    outputs(1878) <= (layer6_outputs(2076)) xor (layer6_outputs(19));
    outputs(1879) <= not(layer6_outputs(2253));
    outputs(1880) <= (layer6_outputs(1112)) xor (layer6_outputs(1484));
    outputs(1881) <= not((layer6_outputs(744)) xor (layer6_outputs(2304)));
    outputs(1882) <= (layer6_outputs(1125)) and not (layer6_outputs(1064));
    outputs(1883) <= layer6_outputs(2358);
    outputs(1884) <= not(layer6_outputs(1672));
    outputs(1885) <= not((layer6_outputs(437)) or (layer6_outputs(1391)));
    outputs(1886) <= not(layer6_outputs(1393));
    outputs(1887) <= not((layer6_outputs(304)) xor (layer6_outputs(1068)));
    outputs(1888) <= (layer6_outputs(654)) xor (layer6_outputs(370));
    outputs(1889) <= layer6_outputs(201);
    outputs(1890) <= not(layer6_outputs(1178));
    outputs(1891) <= layer6_outputs(6);
    outputs(1892) <= layer6_outputs(2292);
    outputs(1893) <= layer6_outputs(1210);
    outputs(1894) <= (layer6_outputs(855)) xor (layer6_outputs(1345));
    outputs(1895) <= layer6_outputs(768);
    outputs(1896) <= not(layer6_outputs(340));
    outputs(1897) <= layer6_outputs(1461);
    outputs(1898) <= layer6_outputs(832);
    outputs(1899) <= (layer6_outputs(2488)) and (layer6_outputs(421));
    outputs(1900) <= not(layer6_outputs(2269));
    outputs(1901) <= not(layer6_outputs(1661));
    outputs(1902) <= (layer6_outputs(1326)) and not (layer6_outputs(47));
    outputs(1903) <= not(layer6_outputs(2188));
    outputs(1904) <= not((layer6_outputs(221)) or (layer6_outputs(2303)));
    outputs(1905) <= (layer6_outputs(168)) and (layer6_outputs(945));
    outputs(1906) <= not((layer6_outputs(981)) xor (layer6_outputs(558)));
    outputs(1907) <= layer6_outputs(2310);
    outputs(1908) <= layer6_outputs(2340);
    outputs(1909) <= not((layer6_outputs(1653)) or (layer6_outputs(1232)));
    outputs(1910) <= layer6_outputs(23);
    outputs(1911) <= (layer6_outputs(720)) and (layer6_outputs(519));
    outputs(1912) <= not(layer6_outputs(1791));
    outputs(1913) <= not((layer6_outputs(209)) or (layer6_outputs(60)));
    outputs(1914) <= layer6_outputs(1056);
    outputs(1915) <= not((layer6_outputs(1429)) xor (layer6_outputs(2117)));
    outputs(1916) <= layer6_outputs(1587);
    outputs(1917) <= not(layer6_outputs(236)) or (layer6_outputs(2162));
    outputs(1918) <= not(layer6_outputs(202));
    outputs(1919) <= not((layer6_outputs(2369)) or (layer6_outputs(1070)));
    outputs(1920) <= layer6_outputs(1644);
    outputs(1921) <= layer6_outputs(589);
    outputs(1922) <= not(layer6_outputs(2202));
    outputs(1923) <= not((layer6_outputs(341)) or (layer6_outputs(1202)));
    outputs(1924) <= not(layer6_outputs(1752));
    outputs(1925) <= not(layer6_outputs(2201));
    outputs(1926) <= (layer6_outputs(1846)) and not (layer6_outputs(604));
    outputs(1927) <= layer6_outputs(1961);
    outputs(1928) <= not(layer6_outputs(1078));
    outputs(1929) <= not(layer6_outputs(1096)) or (layer6_outputs(30));
    outputs(1930) <= not((layer6_outputs(2037)) or (layer6_outputs(1512)));
    outputs(1931) <= not((layer6_outputs(2015)) or (layer6_outputs(395)));
    outputs(1932) <= (layer6_outputs(969)) or (layer6_outputs(1491));
    outputs(1933) <= (layer6_outputs(1339)) xor (layer6_outputs(1686));
    outputs(1934) <= not(layer6_outputs(462));
    outputs(1935) <= not(layer6_outputs(1864));
    outputs(1936) <= layer6_outputs(2478);
    outputs(1937) <= not((layer6_outputs(1120)) or (layer6_outputs(425)));
    outputs(1938) <= not((layer6_outputs(1072)) or (layer6_outputs(835)));
    outputs(1939) <= not(layer6_outputs(1622));
    outputs(1940) <= not(layer6_outputs(1534));
    outputs(1941) <= not((layer6_outputs(167)) xor (layer6_outputs(1246)));
    outputs(1942) <= layer6_outputs(2210);
    outputs(1943) <= layer6_outputs(1352);
    outputs(1944) <= (layer6_outputs(1938)) xor (layer6_outputs(401));
    outputs(1945) <= layer6_outputs(1160);
    outputs(1946) <= layer6_outputs(1013);
    outputs(1947) <= layer6_outputs(760);
    outputs(1948) <= (layer6_outputs(329)) xor (layer6_outputs(1721));
    outputs(1949) <= layer6_outputs(187);
    outputs(1950) <= (layer6_outputs(801)) xor (layer6_outputs(1369));
    outputs(1951) <= not(layer6_outputs(940));
    outputs(1952) <= layer6_outputs(640);
    outputs(1953) <= (layer6_outputs(540)) and not (layer6_outputs(2461));
    outputs(1954) <= (layer6_outputs(2227)) xor (layer6_outputs(870));
    outputs(1955) <= (layer6_outputs(180)) and (layer6_outputs(2385));
    outputs(1956) <= not((layer6_outputs(2131)) xor (layer6_outputs(150)));
    outputs(1957) <= (layer6_outputs(745)) and (layer6_outputs(2002));
    outputs(1958) <= layer6_outputs(1869);
    outputs(1959) <= layer6_outputs(1697);
    outputs(1960) <= (layer6_outputs(2390)) and not (layer6_outputs(2001));
    outputs(1961) <= not((layer6_outputs(249)) or (layer6_outputs(382)));
    outputs(1962) <= not(layer6_outputs(1211));
    outputs(1963) <= (layer6_outputs(1638)) xor (layer6_outputs(500));
    outputs(1964) <= not((layer6_outputs(599)) xor (layer6_outputs(2420)));
    outputs(1965) <= not((layer6_outputs(2374)) xor (layer6_outputs(601)));
    outputs(1966) <= layer6_outputs(950);
    outputs(1967) <= (layer6_outputs(201)) xor (layer6_outputs(883));
    outputs(1968) <= not(layer6_outputs(853));
    outputs(1969) <= not((layer6_outputs(1768)) xor (layer6_outputs(150)));
    outputs(1970) <= (layer6_outputs(1909)) and not (layer6_outputs(1115));
    outputs(1971) <= (layer6_outputs(2523)) and (layer6_outputs(1382));
    outputs(1972) <= (layer6_outputs(711)) xor (layer6_outputs(1374));
    outputs(1973) <= (layer6_outputs(855)) xor (layer6_outputs(109));
    outputs(1974) <= not(layer6_outputs(1672));
    outputs(1975) <= layer6_outputs(1000);
    outputs(1976) <= layer6_outputs(1438);
    outputs(1977) <= (layer6_outputs(429)) and (layer6_outputs(1798));
    outputs(1978) <= layer6_outputs(836);
    outputs(1979) <= not((layer6_outputs(2016)) xor (layer6_outputs(2310)));
    outputs(1980) <= not(layer6_outputs(835));
    outputs(1981) <= layer6_outputs(406);
    outputs(1982) <= (layer6_outputs(1997)) and not (layer6_outputs(1493));
    outputs(1983) <= layer6_outputs(355);
    outputs(1984) <= not(layer6_outputs(2175));
    outputs(1985) <= (layer6_outputs(1743)) and not (layer6_outputs(1576));
    outputs(1986) <= (layer6_outputs(651)) and not (layer6_outputs(1816));
    outputs(1987) <= not(layer6_outputs(2262));
    outputs(1988) <= not(layer6_outputs(592)) or (layer6_outputs(2314));
    outputs(1989) <= layer6_outputs(27);
    outputs(1990) <= (layer6_outputs(1465)) and not (layer6_outputs(1107));
    outputs(1991) <= (layer6_outputs(1831)) and not (layer6_outputs(813));
    outputs(1992) <= not(layer6_outputs(2438));
    outputs(1993) <= (layer6_outputs(1807)) xor (layer6_outputs(799));
    outputs(1994) <= not((layer6_outputs(1283)) or (layer6_outputs(2318)));
    outputs(1995) <= layer6_outputs(550);
    outputs(1996) <= not((layer6_outputs(1731)) xor (layer6_outputs(1822)));
    outputs(1997) <= layer6_outputs(1829);
    outputs(1998) <= not(layer6_outputs(2313));
    outputs(1999) <= layer6_outputs(421);
    outputs(2000) <= not(layer6_outputs(1323));
    outputs(2001) <= not(layer6_outputs(2104));
    outputs(2002) <= (layer6_outputs(992)) xor (layer6_outputs(1451));
    outputs(2003) <= (layer6_outputs(894)) and not (layer6_outputs(175));
    outputs(2004) <= not(layer6_outputs(826));
    outputs(2005) <= (layer6_outputs(2456)) and not (layer6_outputs(1385));
    outputs(2006) <= layer6_outputs(1170);
    outputs(2007) <= layer6_outputs(1669);
    outputs(2008) <= not(layer6_outputs(2192));
    outputs(2009) <= layer6_outputs(2229);
    outputs(2010) <= not(layer6_outputs(1024)) or (layer6_outputs(1890));
    outputs(2011) <= (layer6_outputs(1347)) and not (layer6_outputs(2136));
    outputs(2012) <= (layer6_outputs(1664)) and not (layer6_outputs(1839));
    outputs(2013) <= not((layer6_outputs(1598)) or (layer6_outputs(1666)));
    outputs(2014) <= (layer6_outputs(1671)) or (layer6_outputs(2028));
    outputs(2015) <= not((layer6_outputs(1022)) xor (layer6_outputs(849)));
    outputs(2016) <= not(layer6_outputs(919));
    outputs(2017) <= layer6_outputs(1514);
    outputs(2018) <= layer6_outputs(1032);
    outputs(2019) <= not(layer6_outputs(1416));
    outputs(2020) <= not(layer6_outputs(687));
    outputs(2021) <= not(layer6_outputs(144));
    outputs(2022) <= (layer6_outputs(534)) xor (layer6_outputs(2399));
    outputs(2023) <= (layer6_outputs(1127)) and not (layer6_outputs(2338));
    outputs(2024) <= not(layer6_outputs(1178));
    outputs(2025) <= not(layer6_outputs(1552));
    outputs(2026) <= not(layer6_outputs(1652));
    outputs(2027) <= not(layer6_outputs(420));
    outputs(2028) <= layer6_outputs(1365);
    outputs(2029) <= not((layer6_outputs(1679)) or (layer6_outputs(1168)));
    outputs(2030) <= not((layer6_outputs(2460)) or (layer6_outputs(249)));
    outputs(2031) <= not(layer6_outputs(905));
    outputs(2032) <= layer6_outputs(665);
    outputs(2033) <= not(layer6_outputs(2049));
    outputs(2034) <= (layer6_outputs(2022)) and (layer6_outputs(379));
    outputs(2035) <= not(layer6_outputs(148));
    outputs(2036) <= not((layer6_outputs(1967)) or (layer6_outputs(174)));
    outputs(2037) <= not((layer6_outputs(1086)) xor (layer6_outputs(2154)));
    outputs(2038) <= not((layer6_outputs(1151)) xor (layer6_outputs(1161)));
    outputs(2039) <= not(layer6_outputs(426));
    outputs(2040) <= not(layer6_outputs(1735));
    outputs(2041) <= not((layer6_outputs(2237)) xor (layer6_outputs(58)));
    outputs(2042) <= not(layer6_outputs(8));
    outputs(2043) <= (layer6_outputs(28)) and not (layer6_outputs(1253));
    outputs(2044) <= not((layer6_outputs(746)) xor (layer6_outputs(643)));
    outputs(2045) <= (layer6_outputs(2230)) and not (layer6_outputs(1779));
    outputs(2046) <= not((layer6_outputs(2020)) xor (layer6_outputs(890)));
    outputs(2047) <= layer6_outputs(381);
    outputs(2048) <= not((layer6_outputs(1761)) and (layer6_outputs(1365)));
    outputs(2049) <= not((layer6_outputs(485)) and (layer6_outputs(1155)));
    outputs(2050) <= layer6_outputs(818);
    outputs(2051) <= not(layer6_outputs(2268)) or (layer6_outputs(2405));
    outputs(2052) <= layer6_outputs(1120);
    outputs(2053) <= not((layer6_outputs(696)) xor (layer6_outputs(1467)));
    outputs(2054) <= (layer6_outputs(270)) xor (layer6_outputs(1383));
    outputs(2055) <= (layer6_outputs(1592)) xor (layer6_outputs(2257));
    outputs(2056) <= layer6_outputs(1067);
    outputs(2057) <= layer6_outputs(1685);
    outputs(2058) <= layer6_outputs(2513);
    outputs(2059) <= not(layer6_outputs(291));
    outputs(2060) <= (layer6_outputs(2454)) and not (layer6_outputs(1110));
    outputs(2061) <= not(layer6_outputs(1921));
    outputs(2062) <= layer6_outputs(1675);
    outputs(2063) <= not(layer6_outputs(616));
    outputs(2064) <= not((layer6_outputs(2093)) or (layer6_outputs(1538)));
    outputs(2065) <= not(layer6_outputs(2503));
    outputs(2066) <= layer6_outputs(70);
    outputs(2067) <= (layer6_outputs(1473)) or (layer6_outputs(1175));
    outputs(2068) <= (layer6_outputs(2259)) xor (layer6_outputs(1920));
    outputs(2069) <= (layer6_outputs(290)) xor (layer6_outputs(2545));
    outputs(2070) <= layer6_outputs(723);
    outputs(2071) <= layer6_outputs(1380);
    outputs(2072) <= not((layer6_outputs(1348)) xor (layer6_outputs(140)));
    outputs(2073) <= layer6_outputs(715);
    outputs(2074) <= not(layer6_outputs(2024)) or (layer6_outputs(1395));
    outputs(2075) <= not(layer6_outputs(2018));
    outputs(2076) <= not((layer6_outputs(2126)) and (layer6_outputs(2200)));
    outputs(2077) <= not(layer6_outputs(573));
    outputs(2078) <= layer6_outputs(2189);
    outputs(2079) <= (layer6_outputs(1361)) xor (layer6_outputs(386));
    outputs(2080) <= layer6_outputs(2);
    outputs(2081) <= not((layer6_outputs(495)) and (layer6_outputs(1533)));
    outputs(2082) <= layer6_outputs(2453);
    outputs(2083) <= (layer6_outputs(955)) xor (layer6_outputs(1128));
    outputs(2084) <= not(layer6_outputs(1749));
    outputs(2085) <= layer6_outputs(750);
    outputs(2086) <= (layer6_outputs(1288)) or (layer6_outputs(1071));
    outputs(2087) <= (layer6_outputs(1623)) or (layer6_outputs(97));
    outputs(2088) <= layer6_outputs(2036);
    outputs(2089) <= (layer6_outputs(1030)) or (layer6_outputs(223));
    outputs(2090) <= not(layer6_outputs(440)) or (layer6_outputs(734));
    outputs(2091) <= not(layer6_outputs(1585));
    outputs(2092) <= not(layer6_outputs(1154));
    outputs(2093) <= layer6_outputs(1041);
    outputs(2094) <= layer6_outputs(1279);
    outputs(2095) <= not((layer6_outputs(135)) xor (layer6_outputs(416)));
    outputs(2096) <= (layer6_outputs(2341)) and not (layer6_outputs(338));
    outputs(2097) <= not(layer6_outputs(1566));
    outputs(2098) <= not(layer6_outputs(2109));
    outputs(2099) <= layer6_outputs(682);
    outputs(2100) <= layer6_outputs(878);
    outputs(2101) <= (layer6_outputs(2453)) and not (layer6_outputs(862));
    outputs(2102) <= layer6_outputs(1409);
    outputs(2103) <= (layer6_outputs(618)) xor (layer6_outputs(1441));
    outputs(2104) <= (layer6_outputs(365)) xor (layer6_outputs(2444));
    outputs(2105) <= not(layer6_outputs(20));
    outputs(2106) <= (layer6_outputs(316)) xor (layer6_outputs(1874));
    outputs(2107) <= (layer6_outputs(705)) xor (layer6_outputs(2073));
    outputs(2108) <= (layer6_outputs(2279)) and not (layer6_outputs(578));
    outputs(2109) <= (layer6_outputs(1345)) and (layer6_outputs(1317));
    outputs(2110) <= not(layer6_outputs(972));
    outputs(2111) <= not((layer6_outputs(1408)) and (layer6_outputs(418)));
    outputs(2112) <= layer6_outputs(2371);
    outputs(2113) <= layer6_outputs(92);
    outputs(2114) <= (layer6_outputs(446)) and (layer6_outputs(1063));
    outputs(2115) <= not((layer6_outputs(1772)) and (layer6_outputs(2167)));
    outputs(2116) <= not(layer6_outputs(23));
    outputs(2117) <= not(layer6_outputs(439));
    outputs(2118) <= not((layer6_outputs(2361)) and (layer6_outputs(859)));
    outputs(2119) <= layer6_outputs(322);
    outputs(2120) <= not((layer6_outputs(507)) or (layer6_outputs(1201)));
    outputs(2121) <= (layer6_outputs(850)) xor (layer6_outputs(1848));
    outputs(2122) <= not(layer6_outputs(383));
    outputs(2123) <= not((layer6_outputs(1803)) xor (layer6_outputs(843)));
    outputs(2124) <= not(layer6_outputs(391)) or (layer6_outputs(1477));
    outputs(2125) <= layer6_outputs(1083);
    outputs(2126) <= (layer6_outputs(2372)) xor (layer6_outputs(1779));
    outputs(2127) <= not((layer6_outputs(314)) or (layer6_outputs(914)));
    outputs(2128) <= not(layer6_outputs(2362));
    outputs(2129) <= layer6_outputs(103);
    outputs(2130) <= (layer6_outputs(1719)) and (layer6_outputs(2078));
    outputs(2131) <= layer6_outputs(2305);
    outputs(2132) <= layer6_outputs(2078);
    outputs(2133) <= not(layer6_outputs(1667));
    outputs(2134) <= layer6_outputs(1419);
    outputs(2135) <= layer6_outputs(154);
    outputs(2136) <= (layer6_outputs(1251)) xor (layer6_outputs(719));
    outputs(2137) <= (layer6_outputs(216)) and not (layer6_outputs(2508));
    outputs(2138) <= not(layer6_outputs(1601));
    outputs(2139) <= layer6_outputs(1066);
    outputs(2140) <= layer6_outputs(1314);
    outputs(2141) <= layer6_outputs(634);
    outputs(2142) <= not(layer6_outputs(2010));
    outputs(2143) <= layer6_outputs(2289);
    outputs(2144) <= not(layer6_outputs(2110));
    outputs(2145) <= layer6_outputs(1891);
    outputs(2146) <= (layer6_outputs(543)) or (layer6_outputs(1023));
    outputs(2147) <= not(layer6_outputs(946));
    outputs(2148) <= layer6_outputs(2394);
    outputs(2149) <= (layer6_outputs(1384)) xor (layer6_outputs(1188));
    outputs(2150) <= (layer6_outputs(1738)) and not (layer6_outputs(2027));
    outputs(2151) <= layer6_outputs(91);
    outputs(2152) <= (layer6_outputs(819)) and not (layer6_outputs(374));
    outputs(2153) <= layer6_outputs(638);
    outputs(2154) <= not((layer6_outputs(687)) xor (layer6_outputs(178)));
    outputs(2155) <= layer6_outputs(2013);
    outputs(2156) <= layer6_outputs(2542);
    outputs(2157) <= layer6_outputs(2295);
    outputs(2158) <= not((layer6_outputs(1127)) xor (layer6_outputs(51)));
    outputs(2159) <= (layer6_outputs(1594)) xor (layer6_outputs(1964));
    outputs(2160) <= not((layer6_outputs(1052)) or (layer6_outputs(724)));
    outputs(2161) <= not(layer6_outputs(1375)) or (layer6_outputs(643));
    outputs(2162) <= not(layer6_outputs(1123));
    outputs(2163) <= (layer6_outputs(1262)) and not (layer6_outputs(1394));
    outputs(2164) <= not(layer6_outputs(1745));
    outputs(2165) <= not(layer6_outputs(1956)) or (layer6_outputs(1778));
    outputs(2166) <= (layer6_outputs(172)) xor (layer6_outputs(1944));
    outputs(2167) <= (layer6_outputs(1231)) xor (layer6_outputs(1477));
    outputs(2168) <= not(layer6_outputs(1646));
    outputs(2169) <= not(layer6_outputs(904));
    outputs(2170) <= not(layer6_outputs(494));
    outputs(2171) <= not(layer6_outputs(310));
    outputs(2172) <= (layer6_outputs(1756)) and not (layer6_outputs(343));
    outputs(2173) <= not(layer6_outputs(578));
    outputs(2174) <= not(layer6_outputs(1114));
    outputs(2175) <= layer6_outputs(2406);
    outputs(2176) <= not(layer6_outputs(2011));
    outputs(2177) <= layer6_outputs(1754);
    outputs(2178) <= '1';
    outputs(2179) <= (layer6_outputs(668)) xor (layer6_outputs(425));
    outputs(2180) <= layer6_outputs(1568);
    outputs(2181) <= layer6_outputs(1562);
    outputs(2182) <= layer6_outputs(102);
    outputs(2183) <= layer6_outputs(1603);
    outputs(2184) <= layer6_outputs(1996);
    outputs(2185) <= layer6_outputs(837);
    outputs(2186) <= not(layer6_outputs(2038)) or (layer6_outputs(1445));
    outputs(2187) <= (layer6_outputs(2258)) and not (layer6_outputs(1942));
    outputs(2188) <= (layer6_outputs(89)) and not (layer6_outputs(1349));
    outputs(2189) <= not(layer6_outputs(281));
    outputs(2190) <= (layer6_outputs(1579)) xor (layer6_outputs(1261));
    outputs(2191) <= layer6_outputs(1152);
    outputs(2192) <= not(layer6_outputs(827));
    outputs(2193) <= layer6_outputs(2332);
    outputs(2194) <= layer6_outputs(729);
    outputs(2195) <= layer6_outputs(1969);
    outputs(2196) <= (layer6_outputs(1987)) and not (layer6_outputs(2116));
    outputs(2197) <= (layer6_outputs(407)) and not (layer6_outputs(1401));
    outputs(2198) <= layer6_outputs(1162);
    outputs(2199) <= not(layer6_outputs(90));
    outputs(2200) <= not(layer6_outputs(1810));
    outputs(2201) <= (layer6_outputs(2167)) xor (layer6_outputs(2285));
    outputs(2202) <= not(layer6_outputs(2373)) or (layer6_outputs(2237));
    outputs(2203) <= not((layer6_outputs(1773)) and (layer6_outputs(2177)));
    outputs(2204) <= layer6_outputs(775);
    outputs(2205) <= (layer6_outputs(1080)) and (layer6_outputs(866));
    outputs(2206) <= not((layer6_outputs(1135)) or (layer6_outputs(943)));
    outputs(2207) <= not((layer6_outputs(1788)) xor (layer6_outputs(1655)));
    outputs(2208) <= not(layer6_outputs(848));
    outputs(2209) <= layer6_outputs(1093);
    outputs(2210) <= layer6_outputs(577);
    outputs(2211) <= (layer6_outputs(1262)) and not (layer6_outputs(2478));
    outputs(2212) <= (layer6_outputs(615)) and (layer6_outputs(2305));
    outputs(2213) <= layer6_outputs(1573);
    outputs(2214) <= layer6_outputs(2348);
    outputs(2215) <= layer6_outputs(19);
    outputs(2216) <= (layer6_outputs(156)) xor (layer6_outputs(1599));
    outputs(2217) <= not((layer6_outputs(321)) or (layer6_outputs(1511)));
    outputs(2218) <= not(layer6_outputs(2000)) or (layer6_outputs(2256));
    outputs(2219) <= layer6_outputs(1397);
    outputs(2220) <= not(layer6_outputs(2489));
    outputs(2221) <= not(layer6_outputs(2105));
    outputs(2222) <= not(layer6_outputs(720));
    outputs(2223) <= (layer6_outputs(633)) xor (layer6_outputs(2244));
    outputs(2224) <= (layer6_outputs(1441)) xor (layer6_outputs(1021));
    outputs(2225) <= layer6_outputs(388);
    outputs(2226) <= not(layer6_outputs(597));
    outputs(2227) <= not((layer6_outputs(787)) or (layer6_outputs(2160)));
    outputs(2228) <= not((layer6_outputs(1173)) and (layer6_outputs(1196)));
    outputs(2229) <= not(layer6_outputs(1574));
    outputs(2230) <= not(layer6_outputs(164));
    outputs(2231) <= not(layer6_outputs(595));
    outputs(2232) <= not(layer6_outputs(460));
    outputs(2233) <= layer6_outputs(2475);
    outputs(2234) <= layer6_outputs(2085);
    outputs(2235) <= not(layer6_outputs(62)) or (layer6_outputs(1065));
    outputs(2236) <= layer6_outputs(151);
    outputs(2237) <= not(layer6_outputs(292));
    outputs(2238) <= not((layer6_outputs(642)) and (layer6_outputs(2285)));
    outputs(2239) <= layer6_outputs(2044);
    outputs(2240) <= not(layer6_outputs(616));
    outputs(2241) <= not((layer6_outputs(1870)) xor (layer6_outputs(1100)));
    outputs(2242) <= layer6_outputs(770);
    outputs(2243) <= layer6_outputs(1259);
    outputs(2244) <= (layer6_outputs(57)) and not (layer6_outputs(2165));
    outputs(2245) <= not(layer6_outputs(225));
    outputs(2246) <= not((layer6_outputs(2350)) xor (layer6_outputs(52)));
    outputs(2247) <= not(layer6_outputs(1085));
    outputs(2248) <= (layer6_outputs(337)) xor (layer6_outputs(60));
    outputs(2249) <= layer6_outputs(2403);
    outputs(2250) <= not(layer6_outputs(30));
    outputs(2251) <= not(layer6_outputs(1216));
    outputs(2252) <= not(layer6_outputs(544));
    outputs(2253) <= not(layer6_outputs(936));
    outputs(2254) <= layer6_outputs(2425);
    outputs(2255) <= layer6_outputs(1199);
    outputs(2256) <= not(layer6_outputs(605));
    outputs(2257) <= (layer6_outputs(463)) and not (layer6_outputs(2011));
    outputs(2258) <= layer6_outputs(675);
    outputs(2259) <= (layer6_outputs(2542)) or (layer6_outputs(1885));
    outputs(2260) <= layer6_outputs(831);
    outputs(2261) <= layer6_outputs(993);
    outputs(2262) <= layer6_outputs(1792);
    outputs(2263) <= not(layer6_outputs(2449));
    outputs(2264) <= not(layer6_outputs(768));
    outputs(2265) <= not((layer6_outputs(1467)) and (layer6_outputs(1050)));
    outputs(2266) <= (layer6_outputs(2480)) and not (layer6_outputs(1520));
    outputs(2267) <= not(layer6_outputs(317));
    outputs(2268) <= layer6_outputs(2251);
    outputs(2269) <= not((layer6_outputs(1339)) xor (layer6_outputs(1493)));
    outputs(2270) <= layer6_outputs(2085);
    outputs(2271) <= layer6_outputs(1229);
    outputs(2272) <= layer6_outputs(2119);
    outputs(2273) <= not(layer6_outputs(1429)) or (layer6_outputs(308));
    outputs(2274) <= not(layer6_outputs(1828));
    outputs(2275) <= (layer6_outputs(872)) and not (layer6_outputs(2337));
    outputs(2276) <= layer6_outputs(1973);
    outputs(2277) <= layer6_outputs(979);
    outputs(2278) <= (layer6_outputs(1046)) xor (layer6_outputs(814));
    outputs(2279) <= layer6_outputs(1569);
    outputs(2280) <= layer6_outputs(1888);
    outputs(2281) <= layer6_outputs(1026);
    outputs(2282) <= layer6_outputs(36);
    outputs(2283) <= not(layer6_outputs(1635));
    outputs(2284) <= layer6_outputs(1291);
    outputs(2285) <= not((layer6_outputs(1006)) and (layer6_outputs(1529)));
    outputs(2286) <= not(layer6_outputs(1948));
    outputs(2287) <= not(layer6_outputs(300));
    outputs(2288) <= not(layer6_outputs(43));
    outputs(2289) <= layer6_outputs(2205);
    outputs(2290) <= not(layer6_outputs(2055));
    outputs(2291) <= not((layer6_outputs(430)) or (layer6_outputs(234)));
    outputs(2292) <= layer6_outputs(2098);
    outputs(2293) <= layer6_outputs(2507);
    outputs(2294) <= not(layer6_outputs(1994));
    outputs(2295) <= not(layer6_outputs(2361));
    outputs(2296) <= not(layer6_outputs(1819));
    outputs(2297) <= not(layer6_outputs(415));
    outputs(2298) <= layer6_outputs(1299);
    outputs(2299) <= layer6_outputs(2303);
    outputs(2300) <= layer6_outputs(1614);
    outputs(2301) <= not(layer6_outputs(1811));
    outputs(2302) <= (layer6_outputs(1610)) and not (layer6_outputs(1045));
    outputs(2303) <= (layer6_outputs(579)) and not (layer6_outputs(1711));
    outputs(2304) <= (layer6_outputs(1971)) xor (layer6_outputs(1915));
    outputs(2305) <= layer6_outputs(1596);
    outputs(2306) <= not(layer6_outputs(2088));
    outputs(2307) <= layer6_outputs(241);
    outputs(2308) <= (layer6_outputs(620)) and not (layer6_outputs(2188));
    outputs(2309) <= not(layer6_outputs(956));
    outputs(2310) <= not((layer6_outputs(2224)) and (layer6_outputs(2093)));
    outputs(2311) <= not(layer6_outputs(1734));
    outputs(2312) <= layer6_outputs(490);
    outputs(2313) <= layer6_outputs(393);
    outputs(2314) <= layer6_outputs(1790);
    outputs(2315) <= layer6_outputs(2466);
    outputs(2316) <= not(layer6_outputs(1773));
    outputs(2317) <= layer6_outputs(46);
    outputs(2318) <= not(layer6_outputs(2467));
    outputs(2319) <= not(layer6_outputs(1076));
    outputs(2320) <= layer6_outputs(2554);
    outputs(2321) <= layer6_outputs(1950);
    outputs(2322) <= layer6_outputs(1889);
    outputs(2323) <= not((layer6_outputs(1294)) and (layer6_outputs(1884)));
    outputs(2324) <= not(layer6_outputs(1353));
    outputs(2325) <= layer6_outputs(1796);
    outputs(2326) <= not(layer6_outputs(2318));
    outputs(2327) <= not(layer6_outputs(1229));
    outputs(2328) <= not((layer6_outputs(2349)) or (layer6_outputs(1708)));
    outputs(2329) <= (layer6_outputs(972)) and not (layer6_outputs(1081));
    outputs(2330) <= (layer6_outputs(1039)) and not (layer6_outputs(936));
    outputs(2331) <= layer6_outputs(330);
    outputs(2332) <= not(layer6_outputs(2014));
    outputs(2333) <= not(layer6_outputs(748));
    outputs(2334) <= layer6_outputs(322);
    outputs(2335) <= not(layer6_outputs(1439));
    outputs(2336) <= (layer6_outputs(2497)) xor (layer6_outputs(392));
    outputs(2337) <= layer6_outputs(2425);
    outputs(2338) <= not(layer6_outputs(1716));
    outputs(2339) <= (layer6_outputs(1378)) and (layer6_outputs(1240));
    outputs(2340) <= (layer6_outputs(1404)) xor (layer6_outputs(1179));
    outputs(2341) <= (layer6_outputs(942)) xor (layer6_outputs(1818));
    outputs(2342) <= (layer6_outputs(271)) and (layer6_outputs(1002));
    outputs(2343) <= (layer6_outputs(171)) xor (layer6_outputs(1422));
    outputs(2344) <= (layer6_outputs(278)) and not (layer6_outputs(860));
    outputs(2345) <= not(layer6_outputs(1203));
    outputs(2346) <= not(layer6_outputs(694));
    outputs(2347) <= (layer6_outputs(357)) and not (layer6_outputs(1842));
    outputs(2348) <= layer6_outputs(738);
    outputs(2349) <= not(layer6_outputs(2071));
    outputs(2350) <= (layer6_outputs(653)) xor (layer6_outputs(887));
    outputs(2351) <= (layer6_outputs(233)) xor (layer6_outputs(395));
    outputs(2352) <= not((layer6_outputs(583)) and (layer6_outputs(1722)));
    outputs(2353) <= not(layer6_outputs(820));
    outputs(2354) <= not(layer6_outputs(14));
    outputs(2355) <= (layer6_outputs(1598)) xor (layer6_outputs(1325));
    outputs(2356) <= not(layer6_outputs(2168));
    outputs(2357) <= not(layer6_outputs(2281));
    outputs(2358) <= not(layer6_outputs(815));
    outputs(2359) <= (layer6_outputs(915)) xor (layer6_outputs(1315));
    outputs(2360) <= not((layer6_outputs(2150)) or (layer6_outputs(1885)));
    outputs(2361) <= not((layer6_outputs(934)) xor (layer6_outputs(301)));
    outputs(2362) <= not(layer6_outputs(2017));
    outputs(2363) <= not(layer6_outputs(830));
    outputs(2364) <= not(layer6_outputs(1722));
    outputs(2365) <= not(layer6_outputs(2471));
    outputs(2366) <= layer6_outputs(2442);
    outputs(2367) <= not(layer6_outputs(2482));
    outputs(2368) <= layer6_outputs(188);
    outputs(2369) <= layer6_outputs(1327);
    outputs(2370) <= not((layer6_outputs(2447)) xor (layer6_outputs(2392)));
    outputs(2371) <= layer6_outputs(1901);
    outputs(2372) <= not(layer6_outputs(1211));
    outputs(2373) <= not(layer6_outputs(2161));
    outputs(2374) <= not(layer6_outputs(1912));
    outputs(2375) <= not(layer6_outputs(294));
    outputs(2376) <= (layer6_outputs(1850)) and not (layer6_outputs(1084));
    outputs(2377) <= not((layer6_outputs(2204)) xor (layer6_outputs(2007)));
    outputs(2378) <= (layer6_outputs(2099)) and (layer6_outputs(461));
    outputs(2379) <= not(layer6_outputs(2487));
    outputs(2380) <= layer6_outputs(1014);
    outputs(2381) <= layer6_outputs(280);
    outputs(2382) <= not(layer6_outputs(1708));
    outputs(2383) <= not(layer6_outputs(1854));
    outputs(2384) <= not(layer6_outputs(762));
    outputs(2385) <= layer6_outputs(1156);
    outputs(2386) <= (layer6_outputs(423)) and (layer6_outputs(2025));
    outputs(2387) <= (layer6_outputs(2505)) and not (layer6_outputs(1411));
    outputs(2388) <= layer6_outputs(1520);
    outputs(2389) <= not(layer6_outputs(1683));
    outputs(2390) <= not(layer6_outputs(2178));
    outputs(2391) <= not(layer6_outputs(1583));
    outputs(2392) <= layer6_outputs(1952);
    outputs(2393) <= not((layer6_outputs(1809)) xor (layer6_outputs(966)));
    outputs(2394) <= not(layer6_outputs(1606));
    outputs(2395) <= not(layer6_outputs(891));
    outputs(2396) <= not(layer6_outputs(728));
    outputs(2397) <= not(layer6_outputs(789));
    outputs(2398) <= not(layer6_outputs(1676));
    outputs(2399) <= not(layer6_outputs(1443));
    outputs(2400) <= not((layer6_outputs(275)) xor (layer6_outputs(123)));
    outputs(2401) <= not(layer6_outputs(1899));
    outputs(2402) <= not((layer6_outputs(1005)) xor (layer6_outputs(1140)));
    outputs(2403) <= layer6_outputs(2309);
    outputs(2404) <= layer6_outputs(477);
    outputs(2405) <= not(layer6_outputs(1521));
    outputs(2406) <= layer6_outputs(381);
    outputs(2407) <= not((layer6_outputs(2152)) xor (layer6_outputs(869)));
    outputs(2408) <= not(layer6_outputs(585));
    outputs(2409) <= not(layer6_outputs(2123));
    outputs(2410) <= (layer6_outputs(825)) and not (layer6_outputs(1228));
    outputs(2411) <= (layer6_outputs(1944)) and not (layer6_outputs(345));
    outputs(2412) <= not(layer6_outputs(216));
    outputs(2413) <= layer6_outputs(2003);
    outputs(2414) <= (layer6_outputs(2455)) and (layer6_outputs(1494));
    outputs(2415) <= (layer6_outputs(1724)) xor (layer6_outputs(1536));
    outputs(2416) <= not(layer6_outputs(943));
    outputs(2417) <= (layer6_outputs(1161)) and (layer6_outputs(580));
    outputs(2418) <= not((layer6_outputs(1507)) xor (layer6_outputs(226)));
    outputs(2419) <= layer6_outputs(565);
    outputs(2420) <= not((layer6_outputs(1986)) xor (layer6_outputs(887)));
    outputs(2421) <= not((layer6_outputs(1501)) or (layer6_outputs(1428)));
    outputs(2422) <= (layer6_outputs(2101)) and not (layer6_outputs(568));
    outputs(2423) <= not(layer6_outputs(1417));
    outputs(2424) <= not(layer6_outputs(385));
    outputs(2425) <= not((layer6_outputs(168)) xor (layer6_outputs(606)));
    outputs(2426) <= (layer6_outputs(1814)) xor (layer6_outputs(301));
    outputs(2427) <= not(layer6_outputs(899));
    outputs(2428) <= (layer6_outputs(587)) and not (layer6_outputs(2274));
    outputs(2429) <= not(layer6_outputs(376));
    outputs(2430) <= not(layer6_outputs(917));
    outputs(2431) <= (layer6_outputs(1984)) and (layer6_outputs(2082));
    outputs(2432) <= not(layer6_outputs(1634));
    outputs(2433) <= not(layer6_outputs(179));
    outputs(2434) <= not(layer6_outputs(516));
    outputs(2435) <= not((layer6_outputs(2391)) or (layer6_outputs(1509)));
    outputs(2436) <= layer6_outputs(239);
    outputs(2437) <= layer6_outputs(451);
    outputs(2438) <= not((layer6_outputs(2492)) xor (layer6_outputs(82)));
    outputs(2439) <= not(layer6_outputs(1660));
    outputs(2440) <= layer6_outputs(245);
    outputs(2441) <= (layer6_outputs(2111)) xor (layer6_outputs(650));
    outputs(2442) <= (layer6_outputs(1551)) and (layer6_outputs(990));
    outputs(2443) <= not((layer6_outputs(1766)) xor (layer6_outputs(615)));
    outputs(2444) <= (layer6_outputs(2389)) xor (layer6_outputs(2436));
    outputs(2445) <= (layer6_outputs(2342)) and not (layer6_outputs(1518));
    outputs(2446) <= not(layer6_outputs(2380));
    outputs(2447) <= (layer6_outputs(219)) or (layer6_outputs(1668));
    outputs(2448) <= not(layer6_outputs(1511));
    outputs(2449) <= not(layer6_outputs(717));
    outputs(2450) <= not((layer6_outputs(1301)) xor (layer6_outputs(1599)));
    outputs(2451) <= layer6_outputs(2004);
    outputs(2452) <= not(layer6_outputs(503));
    outputs(2453) <= layer6_outputs(1841);
    outputs(2454) <= (layer6_outputs(33)) and not (layer6_outputs(686));
    outputs(2455) <= (layer6_outputs(1992)) and (layer6_outputs(736));
    outputs(2456) <= not(layer6_outputs(2240)) or (layer6_outputs(555));
    outputs(2457) <= layer6_outputs(2441);
    outputs(2458) <= not(layer6_outputs(53));
    outputs(2459) <= layer6_outputs(2079);
    outputs(2460) <= not(layer6_outputs(2070));
    outputs(2461) <= layer6_outputs(282);
    outputs(2462) <= (layer6_outputs(380)) and not (layer6_outputs(2265));
    outputs(2463) <= layer6_outputs(930);
    outputs(2464) <= layer6_outputs(1016);
    outputs(2465) <= not(layer6_outputs(1244));
    outputs(2466) <= layer6_outputs(2205);
    outputs(2467) <= layer6_outputs(852);
    outputs(2468) <= (layer6_outputs(1327)) and not (layer6_outputs(1674));
    outputs(2469) <= (layer6_outputs(1730)) and not (layer6_outputs(2487));
    outputs(2470) <= layer6_outputs(1398);
    outputs(2471) <= not(layer6_outputs(948));
    outputs(2472) <= (layer6_outputs(2539)) xor (layer6_outputs(2444));
    outputs(2473) <= not(layer6_outputs(2024));
    outputs(2474) <= (layer6_outputs(2006)) xor (layer6_outputs(1392));
    outputs(2475) <= layer6_outputs(510);
    outputs(2476) <= not(layer6_outputs(503));
    outputs(2477) <= not((layer6_outputs(2501)) or (layer6_outputs(1959)));
    outputs(2478) <= layer6_outputs(712);
    outputs(2479) <= layer6_outputs(2013);
    outputs(2480) <= not(layer6_outputs(1892));
    outputs(2481) <= layer6_outputs(1062);
    outputs(2482) <= not((layer6_outputs(1753)) xor (layer6_outputs(895)));
    outputs(2483) <= (layer6_outputs(161)) xor (layer6_outputs(983));
    outputs(2484) <= not(layer6_outputs(2467)) or (layer6_outputs(1519));
    outputs(2485) <= (layer6_outputs(399)) xor (layer6_outputs(1386));
    outputs(2486) <= layer6_outputs(1627);
    outputs(2487) <= not((layer6_outputs(2227)) and (layer6_outputs(1153)));
    outputs(2488) <= layer6_outputs(55);
    outputs(2489) <= layer6_outputs(1786);
    outputs(2490) <= layer6_outputs(729);
    outputs(2491) <= not(layer6_outputs(432));
    outputs(2492) <= not((layer6_outputs(13)) or (layer6_outputs(1256)));
    outputs(2493) <= layer6_outputs(312);
    outputs(2494) <= not(layer6_outputs(1606));
    outputs(2495) <= (layer6_outputs(630)) and not (layer6_outputs(1823));
    outputs(2496) <= layer6_outputs(1575);
    outputs(2497) <= layer6_outputs(1386);
    outputs(2498) <= layer6_outputs(22);
    outputs(2499) <= (layer6_outputs(2366)) or (layer6_outputs(607));
    outputs(2500) <= not((layer6_outputs(2263)) xor (layer6_outputs(1077)));
    outputs(2501) <= not(layer6_outputs(2449));
    outputs(2502) <= not((layer6_outputs(2080)) xor (layer6_outputs(1701)));
    outputs(2503) <= not(layer6_outputs(2218));
    outputs(2504) <= not((layer6_outputs(478)) xor (layer6_outputs(888)));
    outputs(2505) <= not(layer6_outputs(49));
    outputs(2506) <= (layer6_outputs(389)) xor (layer6_outputs(2399));
    outputs(2507) <= not(layer6_outputs(144));
    outputs(2508) <= not(layer6_outputs(465));
    outputs(2509) <= not(layer6_outputs(998));
    outputs(2510) <= not(layer6_outputs(1295));
    outputs(2511) <= layer6_outputs(476);
    outputs(2512) <= not(layer6_outputs(875));
    outputs(2513) <= layer6_outputs(137);
    outputs(2514) <= not((layer6_outputs(878)) xor (layer6_outputs(2037)));
    outputs(2515) <= not(layer6_outputs(2035));
    outputs(2516) <= not((layer6_outputs(116)) xor (layer6_outputs(1817)));
    outputs(2517) <= (layer6_outputs(2533)) xor (layer6_outputs(1175));
    outputs(2518) <= layer6_outputs(930);
    outputs(2519) <= layer6_outputs(1225);
    outputs(2520) <= not((layer6_outputs(1245)) xor (layer6_outputs(977)));
    outputs(2521) <= (layer6_outputs(1806)) xor (layer6_outputs(530));
    outputs(2522) <= (layer6_outputs(901)) and (layer6_outputs(2266));
    outputs(2523) <= not(layer6_outputs(851));
    outputs(2524) <= not(layer6_outputs(1445));
    outputs(2525) <= not(layer6_outputs(1215));
    outputs(2526) <= not((layer6_outputs(2140)) xor (layer6_outputs(69)));
    outputs(2527) <= not((layer6_outputs(1159)) and (layer6_outputs(1602)));
    outputs(2528) <= not((layer6_outputs(2495)) xor (layer6_outputs(106)));
    outputs(2529) <= not(layer6_outputs(374));
    outputs(2530) <= (layer6_outputs(1061)) and not (layer6_outputs(2388));
    outputs(2531) <= not((layer6_outputs(2301)) and (layer6_outputs(2552)));
    outputs(2532) <= layer6_outputs(255);
    outputs(2533) <= (layer6_outputs(364)) and not (layer6_outputs(1977));
    outputs(2534) <= (layer6_outputs(1431)) or (layer6_outputs(203));
    outputs(2535) <= (layer6_outputs(1803)) xor (layer6_outputs(1847));
    outputs(2536) <= layer6_outputs(460);
    outputs(2537) <= layer6_outputs(2329);
    outputs(2538) <= (layer6_outputs(2006)) and not (layer6_outputs(2391));
    outputs(2539) <= (layer6_outputs(821)) and (layer6_outputs(1612));
    outputs(2540) <= (layer6_outputs(1455)) or (layer6_outputs(1272));
    outputs(2541) <= (layer6_outputs(1689)) and (layer6_outputs(1427));
    outputs(2542) <= (layer6_outputs(1414)) xor (layer6_outputs(811));
    outputs(2543) <= layer6_outputs(656);
    outputs(2544) <= not(layer6_outputs(2373));
    outputs(2545) <= not(layer6_outputs(2320));
    outputs(2546) <= not(layer6_outputs(1435));
    outputs(2547) <= not(layer6_outputs(2339));
    outputs(2548) <= (layer6_outputs(1985)) and (layer6_outputs(1884));
    outputs(2549) <= (layer6_outputs(2184)) and (layer6_outputs(1450));
    outputs(2550) <= layer6_outputs(2400);
    outputs(2551) <= layer6_outputs(1009);
    outputs(2552) <= layer6_outputs(1858);
    outputs(2553) <= not(layer6_outputs(2343));
    outputs(2554) <= not(layer6_outputs(1380)) or (layer6_outputs(857));
    outputs(2555) <= (layer6_outputs(2081)) xor (layer6_outputs(618));
    outputs(2556) <= not(layer6_outputs(2540));
    outputs(2557) <= not(layer6_outputs(1767));
    outputs(2558) <= layer6_outputs(1608);
    outputs(2559) <= not(layer6_outputs(2196));

end Behavioral;
