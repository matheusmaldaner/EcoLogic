library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs: in std_logic_vector(1023 downto 0);
        outputs: out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs: std_logic_vector(10239 downto 0);

begin
    layer0_outputs(0) <= not (a xor b);
    layer0_outputs(1) <= not (a or b);
    layer0_outputs(2) <= not (a or b);
    layer0_outputs(3) <= not (a or b);
    layer0_outputs(4) <= not b or a;
    layer0_outputs(5) <= a or b;
    layer0_outputs(6) <= not (a or b);
    layer0_outputs(7) <= a xor b;
    layer0_outputs(8) <= a xor b;
    layer0_outputs(9) <= a or b;
    layer0_outputs(10) <= not b;
    layer0_outputs(11) <= not (a and b);
    layer0_outputs(12) <= not b or a;
    layer0_outputs(13) <= not b;
    layer0_outputs(14) <= not a;
    layer0_outputs(15) <= not (a or b);
    layer0_outputs(16) <= b and not a;
    layer0_outputs(17) <= a or b;
    layer0_outputs(18) <= not (a and b);
    layer0_outputs(19) <= a;
    layer0_outputs(20) <= a xor b;
    layer0_outputs(21) <= not (a or b);
    layer0_outputs(22) <= a and not b;
    layer0_outputs(23) <= not a or b;
    layer0_outputs(24) <= a or b;
    layer0_outputs(25) <= not a;
    layer0_outputs(26) <= not b or a;
    layer0_outputs(27) <= a and b;
    layer0_outputs(28) <= b;
    layer0_outputs(29) <= b;
    layer0_outputs(30) <= a or b;
    layer0_outputs(31) <= a and not b;
    layer0_outputs(32) <= a and b;
    layer0_outputs(33) <= a or b;
    layer0_outputs(34) <= not (a or b);
    layer0_outputs(35) <= b;
    layer0_outputs(36) <= a and not b;
    layer0_outputs(37) <= not a;
    layer0_outputs(38) <= b and not a;
    layer0_outputs(39) <= b;
    layer0_outputs(40) <= '0';
    layer0_outputs(41) <= b and not a;
    layer0_outputs(42) <= b;
    layer0_outputs(43) <= not (a xor b);
    layer0_outputs(44) <= not (a or b);
    layer0_outputs(45) <= not b;
    layer0_outputs(46) <= a and not b;
    layer0_outputs(47) <= not (a xor b);
    layer0_outputs(48) <= b;
    layer0_outputs(49) <= a and b;
    layer0_outputs(50) <= a;
    layer0_outputs(51) <= not (a xor b);
    layer0_outputs(52) <= b and not a;
    layer0_outputs(53) <= not (a xor b);
    layer0_outputs(54) <= a xor b;
    layer0_outputs(55) <= b and not a;
    layer0_outputs(56) <= not (a or b);
    layer0_outputs(57) <= not (a xor b);
    layer0_outputs(58) <= not (a and b);
    layer0_outputs(59) <= a or b;
    layer0_outputs(60) <= a or b;
    layer0_outputs(61) <= a or b;
    layer0_outputs(62) <= a or b;
    layer0_outputs(63) <= a;
    layer0_outputs(64) <= not (a xor b);
    layer0_outputs(65) <= a or b;
    layer0_outputs(66) <= a;
    layer0_outputs(67) <= '1';
    layer0_outputs(68) <= not a;
    layer0_outputs(69) <= not (a xor b);
    layer0_outputs(70) <= not (a xor b);
    layer0_outputs(71) <= not a;
    layer0_outputs(72) <= a;
    layer0_outputs(73) <= not (a xor b);
    layer0_outputs(74) <= a xor b;
    layer0_outputs(75) <= a or b;
    layer0_outputs(76) <= b;
    layer0_outputs(77) <= not (a or b);
    layer0_outputs(78) <= not (a or b);
    layer0_outputs(79) <= not a;
    layer0_outputs(80) <= b and not a;
    layer0_outputs(81) <= not b or a;
    layer0_outputs(82) <= not b;
    layer0_outputs(83) <= b;
    layer0_outputs(84) <= not a or b;
    layer0_outputs(85) <= b;
    layer0_outputs(86) <= b;
    layer0_outputs(87) <= not b;
    layer0_outputs(88) <= not (a or b);
    layer0_outputs(89) <= a and not b;
    layer0_outputs(90) <= a xor b;
    layer0_outputs(91) <= a and b;
    layer0_outputs(92) <= not b or a;
    layer0_outputs(93) <= not (a or b);
    layer0_outputs(94) <= a or b;
    layer0_outputs(95) <= a or b;
    layer0_outputs(96) <= not (a xor b);
    layer0_outputs(97) <= not a or b;
    layer0_outputs(98) <= not (a xor b);
    layer0_outputs(99) <= not (a xor b);
    layer0_outputs(100) <= not a or b;
    layer0_outputs(101) <= a xor b;
    layer0_outputs(102) <= a xor b;
    layer0_outputs(103) <= not b;
    layer0_outputs(104) <= a or b;
    layer0_outputs(105) <= not (a or b);
    layer0_outputs(106) <= not (a or b);
    layer0_outputs(107) <= a and not b;
    layer0_outputs(108) <= b and not a;
    layer0_outputs(109) <= a xor b;
    layer0_outputs(110) <= not (a xor b);
    layer0_outputs(111) <= b and not a;
    layer0_outputs(112) <= not a or b;
    layer0_outputs(113) <= a;
    layer0_outputs(114) <= not a or b;
    layer0_outputs(115) <= not (a xor b);
    layer0_outputs(116) <= not b;
    layer0_outputs(117) <= a;
    layer0_outputs(118) <= not a;
    layer0_outputs(119) <= not b;
    layer0_outputs(120) <= not (a or b);
    layer0_outputs(121) <= not (a or b);
    layer0_outputs(122) <= not b;
    layer0_outputs(123) <= not (a or b);
    layer0_outputs(124) <= not (a or b);
    layer0_outputs(125) <= a or b;
    layer0_outputs(126) <= '0';
    layer0_outputs(127) <= b and not a;
    layer0_outputs(128) <= b and not a;
    layer0_outputs(129) <= not (a or b);
    layer0_outputs(130) <= not (a xor b);
    layer0_outputs(131) <= not b or a;
    layer0_outputs(132) <= not a;
    layer0_outputs(133) <= '0';
    layer0_outputs(134) <= not (a xor b);
    layer0_outputs(135) <= a xor b;
    layer0_outputs(136) <= b and not a;
    layer0_outputs(137) <= b and not a;
    layer0_outputs(138) <= not (a xor b);
    layer0_outputs(139) <= '0';
    layer0_outputs(140) <= b;
    layer0_outputs(141) <= a xor b;
    layer0_outputs(142) <= not b;
    layer0_outputs(143) <= not (a or b);
    layer0_outputs(144) <= not (a and b);
    layer0_outputs(145) <= a and not b;
    layer0_outputs(146) <= a or b;
    layer0_outputs(147) <= not b;
    layer0_outputs(148) <= a or b;
    layer0_outputs(149) <= not b or a;
    layer0_outputs(150) <= b and not a;
    layer0_outputs(151) <= not a or b;
    layer0_outputs(152) <= not b or a;
    layer0_outputs(153) <= b;
    layer0_outputs(154) <= not (a or b);
    layer0_outputs(155) <= not a or b;
    layer0_outputs(156) <= not (a xor b);
    layer0_outputs(157) <= a xor b;
    layer0_outputs(158) <= b and not a;
    layer0_outputs(159) <= not (a xor b);
    layer0_outputs(160) <= '1';
    layer0_outputs(161) <= not b or a;
    layer0_outputs(162) <= not (a or b);
    layer0_outputs(163) <= a or b;
    layer0_outputs(164) <= not (a xor b);
    layer0_outputs(165) <= not b;
    layer0_outputs(166) <= not b;
    layer0_outputs(167) <= a or b;
    layer0_outputs(168) <= a and not b;
    layer0_outputs(169) <= a xor b;
    layer0_outputs(170) <= b;
    layer0_outputs(171) <= a or b;
    layer0_outputs(172) <= not (a or b);
    layer0_outputs(173) <= not (a and b);
    layer0_outputs(174) <= not (a or b);
    layer0_outputs(175) <= not (a or b);
    layer0_outputs(176) <= '1';
    layer0_outputs(177) <= not (a xor b);
    layer0_outputs(178) <= b;
    layer0_outputs(179) <= a xor b;
    layer0_outputs(180) <= a or b;
    layer0_outputs(181) <= not b;
    layer0_outputs(182) <= not (a xor b);
    layer0_outputs(183) <= a and not b;
    layer0_outputs(184) <= a and not b;
    layer0_outputs(185) <= a;
    layer0_outputs(186) <= not a or b;
    layer0_outputs(187) <= '1';
    layer0_outputs(188) <= a;
    layer0_outputs(189) <= b and not a;
    layer0_outputs(190) <= a xor b;
    layer0_outputs(191) <= a or b;
    layer0_outputs(192) <= a;
    layer0_outputs(193) <= a or b;
    layer0_outputs(194) <= not b;
    layer0_outputs(195) <= not (a or b);
    layer0_outputs(196) <= not b;
    layer0_outputs(197) <= not b or a;
    layer0_outputs(198) <= a xor b;
    layer0_outputs(199) <= not (a xor b);
    layer0_outputs(200) <= not a;
    layer0_outputs(201) <= a and not b;
    layer0_outputs(202) <= b and not a;
    layer0_outputs(203) <= not b;
    layer0_outputs(204) <= not b;
    layer0_outputs(205) <= not a or b;
    layer0_outputs(206) <= a or b;
    layer0_outputs(207) <= not (a xor b);
    layer0_outputs(208) <= a xor b;
    layer0_outputs(209) <= b and not a;
    layer0_outputs(210) <= a xor b;
    layer0_outputs(211) <= b and not a;
    layer0_outputs(212) <= a;
    layer0_outputs(213) <= a or b;
    layer0_outputs(214) <= not (a xor b);
    layer0_outputs(215) <= not (a or b);
    layer0_outputs(216) <= a xor b;
    layer0_outputs(217) <= not a or b;
    layer0_outputs(218) <= not (a or b);
    layer0_outputs(219) <= a xor b;
    layer0_outputs(220) <= not a or b;
    layer0_outputs(221) <= b and not a;
    layer0_outputs(222) <= b and not a;
    layer0_outputs(223) <= a or b;
    layer0_outputs(224) <= not (a and b);
    layer0_outputs(225) <= not (a xor b);
    layer0_outputs(226) <= not a;
    layer0_outputs(227) <= not (a xor b);
    layer0_outputs(228) <= not (a or b);
    layer0_outputs(229) <= not b;
    layer0_outputs(230) <= not (a xor b);
    layer0_outputs(231) <= b and not a;
    layer0_outputs(232) <= a or b;
    layer0_outputs(233) <= not (a or b);
    layer0_outputs(234) <= '0';
    layer0_outputs(235) <= not b;
    layer0_outputs(236) <= b and not a;
    layer0_outputs(237) <= not a or b;
    layer0_outputs(238) <= not a;
    layer0_outputs(239) <= not (a or b);
    layer0_outputs(240) <= a or b;
    layer0_outputs(241) <= '1';
    layer0_outputs(242) <= not (a xor b);
    layer0_outputs(243) <= b;
    layer0_outputs(244) <= a and b;
    layer0_outputs(245) <= a and not b;
    layer0_outputs(246) <= not b;
    layer0_outputs(247) <= a and not b;
    layer0_outputs(248) <= not (a or b);
    layer0_outputs(249) <= not b;
    layer0_outputs(250) <= a or b;
    layer0_outputs(251) <= a xor b;
    layer0_outputs(252) <= not b;
    layer0_outputs(253) <= b;
    layer0_outputs(254) <= '0';
    layer0_outputs(255) <= a xor b;
    layer0_outputs(256) <= a or b;
    layer0_outputs(257) <= a xor b;
    layer0_outputs(258) <= not a;
    layer0_outputs(259) <= not (a or b);
    layer0_outputs(260) <= not (a or b);
    layer0_outputs(261) <= not a or b;
    layer0_outputs(262) <= not (a xor b);
    layer0_outputs(263) <= not a or b;
    layer0_outputs(264) <= a or b;
    layer0_outputs(265) <= not a;
    layer0_outputs(266) <= not (a or b);
    layer0_outputs(267) <= a and not b;
    layer0_outputs(268) <= a;
    layer0_outputs(269) <= b;
    layer0_outputs(270) <= a xor b;
    layer0_outputs(271) <= a;
    layer0_outputs(272) <= a and b;
    layer0_outputs(273) <= b and not a;
    layer0_outputs(274) <= not b;
    layer0_outputs(275) <= b and not a;
    layer0_outputs(276) <= not a or b;
    layer0_outputs(277) <= a or b;
    layer0_outputs(278) <= a or b;
    layer0_outputs(279) <= not a;
    layer0_outputs(280) <= a and b;
    layer0_outputs(281) <= not a or b;
    layer0_outputs(282) <= not b;
    layer0_outputs(283) <= not (a or b);
    layer0_outputs(284) <= not (a xor b);
    layer0_outputs(285) <= a or b;
    layer0_outputs(286) <= not b;
    layer0_outputs(287) <= not (a and b);
    layer0_outputs(288) <= not b;
    layer0_outputs(289) <= '0';
    layer0_outputs(290) <= a xor b;
    layer0_outputs(291) <= not a;
    layer0_outputs(292) <= a or b;
    layer0_outputs(293) <= a or b;
    layer0_outputs(294) <= not (a and b);
    layer0_outputs(295) <= not (a or b);
    layer0_outputs(296) <= a;
    layer0_outputs(297) <= b;
    layer0_outputs(298) <= not b or a;
    layer0_outputs(299) <= not a;
    layer0_outputs(300) <= not b or a;
    layer0_outputs(301) <= a and b;
    layer0_outputs(302) <= '0';
    layer0_outputs(303) <= a xor b;
    layer0_outputs(304) <= a or b;
    layer0_outputs(305) <= not (a and b);
    layer0_outputs(306) <= not b;
    layer0_outputs(307) <= b and not a;
    layer0_outputs(308) <= not a or b;
    layer0_outputs(309) <= not (a and b);
    layer0_outputs(310) <= a and b;
    layer0_outputs(311) <= not b or a;
    layer0_outputs(312) <= a or b;
    layer0_outputs(313) <= not (a xor b);
    layer0_outputs(314) <= a and not b;
    layer0_outputs(315) <= a xor b;
    layer0_outputs(316) <= b;
    layer0_outputs(317) <= not (a and b);
    layer0_outputs(318) <= b and not a;
    layer0_outputs(319) <= not b;
    layer0_outputs(320) <= not (a xor b);
    layer0_outputs(321) <= a or b;
    layer0_outputs(322) <= not b or a;
    layer0_outputs(323) <= b;
    layer0_outputs(324) <= a or b;
    layer0_outputs(325) <= a and not b;
    layer0_outputs(326) <= b;
    layer0_outputs(327) <= a or b;
    layer0_outputs(328) <= a;
    layer0_outputs(329) <= a or b;
    layer0_outputs(330) <= not (a and b);
    layer0_outputs(331) <= not (a or b);
    layer0_outputs(332) <= not (a and b);
    layer0_outputs(333) <= not a or b;
    layer0_outputs(334) <= not (a xor b);
    layer0_outputs(335) <= not b or a;
    layer0_outputs(336) <= a xor b;
    layer0_outputs(337) <= not (a xor b);
    layer0_outputs(338) <= not (a and b);
    layer0_outputs(339) <= not (a or b);
    layer0_outputs(340) <= a or b;
    layer0_outputs(341) <= not (a xor b);
    layer0_outputs(342) <= not (a or b);
    layer0_outputs(343) <= not b or a;
    layer0_outputs(344) <= not (a or b);
    layer0_outputs(345) <= not (a xor b);
    layer0_outputs(346) <= a xor b;
    layer0_outputs(347) <= a or b;
    layer0_outputs(348) <= a or b;
    layer0_outputs(349) <= not (a xor b);
    layer0_outputs(350) <= a or b;
    layer0_outputs(351) <= not b;
    layer0_outputs(352) <= a;
    layer0_outputs(353) <= a xor b;
    layer0_outputs(354) <= b and not a;
    layer0_outputs(355) <= a or b;
    layer0_outputs(356) <= not (a xor b);
    layer0_outputs(357) <= a xor b;
    layer0_outputs(358) <= not a or b;
    layer0_outputs(359) <= a;
    layer0_outputs(360) <= not (a xor b);
    layer0_outputs(361) <= not a;
    layer0_outputs(362) <= not (a or b);
    layer0_outputs(363) <= not (a xor b);
    layer0_outputs(364) <= a xor b;
    layer0_outputs(365) <= not b;
    layer0_outputs(366) <= a and not b;
    layer0_outputs(367) <= not (a or b);
    layer0_outputs(368) <= not a;
    layer0_outputs(369) <= a or b;
    layer0_outputs(370) <= a and b;
    layer0_outputs(371) <= not (a or b);
    layer0_outputs(372) <= a or b;
    layer0_outputs(373) <= not (a or b);
    layer0_outputs(374) <= not (a and b);
    layer0_outputs(375) <= a or b;
    layer0_outputs(376) <= a and not b;
    layer0_outputs(377) <= not (a or b);
    layer0_outputs(378) <= not (a xor b);
    layer0_outputs(379) <= a or b;
    layer0_outputs(380) <= b;
    layer0_outputs(381) <= not b or a;
    layer0_outputs(382) <= a xor b;
    layer0_outputs(383) <= not (a xor b);
    layer0_outputs(384) <= not b or a;
    layer0_outputs(385) <= a xor b;
    layer0_outputs(386) <= not b or a;
    layer0_outputs(387) <= b;
    layer0_outputs(388) <= a and b;
    layer0_outputs(389) <= not (a xor b);
    layer0_outputs(390) <= not (a xor b);
    layer0_outputs(391) <= not a;
    layer0_outputs(392) <= not b or a;
    layer0_outputs(393) <= b;
    layer0_outputs(394) <= b and not a;
    layer0_outputs(395) <= a xor b;
    layer0_outputs(396) <= not a;
    layer0_outputs(397) <= not a;
    layer0_outputs(398) <= b;
    layer0_outputs(399) <= a xor b;
    layer0_outputs(400) <= a and not b;
    layer0_outputs(401) <= not b;
    layer0_outputs(402) <= a and not b;
    layer0_outputs(403) <= not b or a;
    layer0_outputs(404) <= not a;
    layer0_outputs(405) <= not (a or b);
    layer0_outputs(406) <= not a;
    layer0_outputs(407) <= not (a or b);
    layer0_outputs(408) <= not (a or b);
    layer0_outputs(409) <= not (a xor b);
    layer0_outputs(410) <= not (a and b);
    layer0_outputs(411) <= not b;
    layer0_outputs(412) <= not (a or b);
    layer0_outputs(413) <= a or b;
    layer0_outputs(414) <= b and not a;
    layer0_outputs(415) <= b and not a;
    layer0_outputs(416) <= not (a or b);
    layer0_outputs(417) <= '0';
    layer0_outputs(418) <= not a;
    layer0_outputs(419) <= not a or b;
    layer0_outputs(420) <= not (a or b);
    layer0_outputs(421) <= not b or a;
    layer0_outputs(422) <= a and b;
    layer0_outputs(423) <= not a or b;
    layer0_outputs(424) <= not (a xor b);
    layer0_outputs(425) <= not (a and b);
    layer0_outputs(426) <= not (a or b);
    layer0_outputs(427) <= not (a or b);
    layer0_outputs(428) <= not a;
    layer0_outputs(429) <= not (a or b);
    layer0_outputs(430) <= not b or a;
    layer0_outputs(431) <= not (a xor b);
    layer0_outputs(432) <= '0';
    layer0_outputs(433) <= a or b;
    layer0_outputs(434) <= a xor b;
    layer0_outputs(435) <= not (a or b);
    layer0_outputs(436) <= not (a xor b);
    layer0_outputs(437) <= not b or a;
    layer0_outputs(438) <= b and not a;
    layer0_outputs(439) <= a;
    layer0_outputs(440) <= b;
    layer0_outputs(441) <= a xor b;
    layer0_outputs(442) <= not b;
    layer0_outputs(443) <= not (a or b);
    layer0_outputs(444) <= a and b;
    layer0_outputs(445) <= a or b;
    layer0_outputs(446) <= not b or a;
    layer0_outputs(447) <= not (a or b);
    layer0_outputs(448) <= not (a or b);
    layer0_outputs(449) <= a;
    layer0_outputs(450) <= a xor b;
    layer0_outputs(451) <= b;
    layer0_outputs(452) <= not b;
    layer0_outputs(453) <= not b or a;
    layer0_outputs(454) <= a xor b;
    layer0_outputs(455) <= '0';
    layer0_outputs(456) <= not a or b;
    layer0_outputs(457) <= not (a xor b);
    layer0_outputs(458) <= not a or b;
    layer0_outputs(459) <= not a;
    layer0_outputs(460) <= a and b;
    layer0_outputs(461) <= not (a or b);
    layer0_outputs(462) <= not (a or b);
    layer0_outputs(463) <= b and not a;
    layer0_outputs(464) <= not (a xor b);
    layer0_outputs(465) <= a xor b;
    layer0_outputs(466) <= a and not b;
    layer0_outputs(467) <= b;
    layer0_outputs(468) <= a;
    layer0_outputs(469) <= b and not a;
    layer0_outputs(470) <= a or b;
    layer0_outputs(471) <= b;
    layer0_outputs(472) <= b and not a;
    layer0_outputs(473) <= a and not b;
    layer0_outputs(474) <= not (a xor b);
    layer0_outputs(475) <= not (a or b);
    layer0_outputs(476) <= not (a or b);
    layer0_outputs(477) <= a xor b;
    layer0_outputs(478) <= '0';
    layer0_outputs(479) <= not (a and b);
    layer0_outputs(480) <= not a;
    layer0_outputs(481) <= not (a or b);
    layer0_outputs(482) <= a or b;
    layer0_outputs(483) <= a;
    layer0_outputs(484) <= not (a or b);
    layer0_outputs(485) <= a xor b;
    layer0_outputs(486) <= not (a or b);
    layer0_outputs(487) <= a and not b;
    layer0_outputs(488) <= a or b;
    layer0_outputs(489) <= a xor b;
    layer0_outputs(490) <= a and b;
    layer0_outputs(491) <= a or b;
    layer0_outputs(492) <= not b;
    layer0_outputs(493) <= a xor b;
    layer0_outputs(494) <= not (a xor b);
    layer0_outputs(495) <= not b;
    layer0_outputs(496) <= not a or b;
    layer0_outputs(497) <= not a;
    layer0_outputs(498) <= a xor b;
    layer0_outputs(499) <= not (a or b);
    layer0_outputs(500) <= a and not b;
    layer0_outputs(501) <= not (a xor b);
    layer0_outputs(502) <= not b or a;
    layer0_outputs(503) <= not a;
    layer0_outputs(504) <= not (a xor b);
    layer0_outputs(505) <= not a;
    layer0_outputs(506) <= '1';
    layer0_outputs(507) <= not a;
    layer0_outputs(508) <= a and not b;
    layer0_outputs(509) <= a and not b;
    layer0_outputs(510) <= a or b;
    layer0_outputs(511) <= not b;
    layer0_outputs(512) <= not (a or b);
    layer0_outputs(513) <= not a or b;
    layer0_outputs(514) <= not (a xor b);
    layer0_outputs(515) <= not a or b;
    layer0_outputs(516) <= '1';
    layer0_outputs(517) <= a xor b;
    layer0_outputs(518) <= a and not b;
    layer0_outputs(519) <= not a or b;
    layer0_outputs(520) <= b and not a;
    layer0_outputs(521) <= a xor b;
    layer0_outputs(522) <= a;
    layer0_outputs(523) <= a and not b;
    layer0_outputs(524) <= not a;
    layer0_outputs(525) <= a or b;
    layer0_outputs(526) <= not (a or b);
    layer0_outputs(527) <= not (a and b);
    layer0_outputs(528) <= a;
    layer0_outputs(529) <= not (a or b);
    layer0_outputs(530) <= not b or a;
    layer0_outputs(531) <= a or b;
    layer0_outputs(532) <= a or b;
    layer0_outputs(533) <= not (a or b);
    layer0_outputs(534) <= b;
    layer0_outputs(535) <= not (a or b);
    layer0_outputs(536) <= not (a xor b);
    layer0_outputs(537) <= not (a or b);
    layer0_outputs(538) <= not a;
    layer0_outputs(539) <= not b or a;
    layer0_outputs(540) <= not b;
    layer0_outputs(541) <= a and not b;
    layer0_outputs(542) <= not (a or b);
    layer0_outputs(543) <= not (a or b);
    layer0_outputs(544) <= not b;
    layer0_outputs(545) <= a or b;
    layer0_outputs(546) <= not (a xor b);
    layer0_outputs(547) <= not (a or b);
    layer0_outputs(548) <= not b or a;
    layer0_outputs(549) <= a or b;
    layer0_outputs(550) <= b;
    layer0_outputs(551) <= b;
    layer0_outputs(552) <= not a or b;
    layer0_outputs(553) <= not (a xor b);
    layer0_outputs(554) <= not b;
    layer0_outputs(555) <= not b or a;
    layer0_outputs(556) <= not b;
    layer0_outputs(557) <= not (a or b);
    layer0_outputs(558) <= a;
    layer0_outputs(559) <= not a or b;
    layer0_outputs(560) <= a or b;
    layer0_outputs(561) <= a xor b;
    layer0_outputs(562) <= not a;
    layer0_outputs(563) <= a or b;
    layer0_outputs(564) <= '0';
    layer0_outputs(565) <= not b;
    layer0_outputs(566) <= not a or b;
    layer0_outputs(567) <= a or b;
    layer0_outputs(568) <= b and not a;
    layer0_outputs(569) <= a and b;
    layer0_outputs(570) <= b;
    layer0_outputs(571) <= not (a xor b);
    layer0_outputs(572) <= '0';
    layer0_outputs(573) <= not (a or b);
    layer0_outputs(574) <= not a;
    layer0_outputs(575) <= not (a or b);
    layer0_outputs(576) <= not (a xor b);
    layer0_outputs(577) <= '0';
    layer0_outputs(578) <= not a or b;
    layer0_outputs(579) <= b;
    layer0_outputs(580) <= '1';
    layer0_outputs(581) <= b and not a;
    layer0_outputs(582) <= '0';
    layer0_outputs(583) <= not a;
    layer0_outputs(584) <= not b;
    layer0_outputs(585) <= b and not a;
    layer0_outputs(586) <= a xor b;
    layer0_outputs(587) <= not (a or b);
    layer0_outputs(588) <= a or b;
    layer0_outputs(589) <= a and not b;
    layer0_outputs(590) <= a or b;
    layer0_outputs(591) <= '0';
    layer0_outputs(592) <= a or b;
    layer0_outputs(593) <= b;
    layer0_outputs(594) <= b;
    layer0_outputs(595) <= not a;
    layer0_outputs(596) <= not (a xor b);
    layer0_outputs(597) <= a xor b;
    layer0_outputs(598) <= not (a or b);
    layer0_outputs(599) <= a or b;
    layer0_outputs(600) <= a;
    layer0_outputs(601) <= not a;
    layer0_outputs(602) <= b;
    layer0_outputs(603) <= a xor b;
    layer0_outputs(604) <= b;
    layer0_outputs(605) <= not a or b;
    layer0_outputs(606) <= not (a xor b);
    layer0_outputs(607) <= a xor b;
    layer0_outputs(608) <= a or b;
    layer0_outputs(609) <= b;
    layer0_outputs(610) <= b and not a;
    layer0_outputs(611) <= not (a or b);
    layer0_outputs(612) <= a or b;
    layer0_outputs(613) <= '1';
    layer0_outputs(614) <= a and not b;
    layer0_outputs(615) <= a or b;
    layer0_outputs(616) <= a or b;
    layer0_outputs(617) <= a or b;
    layer0_outputs(618) <= a and not b;
    layer0_outputs(619) <= not (a and b);
    layer0_outputs(620) <= b;
    layer0_outputs(621) <= a xor b;
    layer0_outputs(622) <= '0';
    layer0_outputs(623) <= '0';
    layer0_outputs(624) <= not (a xor b);
    layer0_outputs(625) <= not (a xor b);
    layer0_outputs(626) <= a or b;
    layer0_outputs(627) <= not b;
    layer0_outputs(628) <= a and not b;
    layer0_outputs(629) <= b;
    layer0_outputs(630) <= not (a or b);
    layer0_outputs(631) <= not (a or b);
    layer0_outputs(632) <= a;
    layer0_outputs(633) <= not b or a;
    layer0_outputs(634) <= a and not b;
    layer0_outputs(635) <= '1';
    layer0_outputs(636) <= b;
    layer0_outputs(637) <= a or b;
    layer0_outputs(638) <= b and not a;
    layer0_outputs(639) <= a or b;
    layer0_outputs(640) <= b and not a;
    layer0_outputs(641) <= a xor b;
    layer0_outputs(642) <= a xor b;
    layer0_outputs(643) <= a and not b;
    layer0_outputs(644) <= not a or b;
    layer0_outputs(645) <= not (a or b);
    layer0_outputs(646) <= a or b;
    layer0_outputs(647) <= not (a or b);
    layer0_outputs(648) <= a;
    layer0_outputs(649) <= b and not a;
    layer0_outputs(650) <= b and not a;
    layer0_outputs(651) <= b and not a;
    layer0_outputs(652) <= a xor b;
    layer0_outputs(653) <= not (a or b);
    layer0_outputs(654) <= a xor b;
    layer0_outputs(655) <= not a or b;
    layer0_outputs(656) <= a;
    layer0_outputs(657) <= not (a or b);
    layer0_outputs(658) <= b and not a;
    layer0_outputs(659) <= not a or b;
    layer0_outputs(660) <= a;
    layer0_outputs(661) <= a and not b;
    layer0_outputs(662) <= not b;
    layer0_outputs(663) <= b and not a;
    layer0_outputs(664) <= not (a xor b);
    layer0_outputs(665) <= b and not a;
    layer0_outputs(666) <= b;
    layer0_outputs(667) <= not a;
    layer0_outputs(668) <= '1';
    layer0_outputs(669) <= not b or a;
    layer0_outputs(670) <= a or b;
    layer0_outputs(671) <= not (a and b);
    layer0_outputs(672) <= a;
    layer0_outputs(673) <= a or b;
    layer0_outputs(674) <= not a or b;
    layer0_outputs(675) <= b and not a;
    layer0_outputs(676) <= not b;
    layer0_outputs(677) <= not (a xor b);
    layer0_outputs(678) <= a;
    layer0_outputs(679) <= a xor b;
    layer0_outputs(680) <= not (a xor b);
    layer0_outputs(681) <= a xor b;
    layer0_outputs(682) <= a or b;
    layer0_outputs(683) <= not (a xor b);
    layer0_outputs(684) <= not b or a;
    layer0_outputs(685) <= b;
    layer0_outputs(686) <= a;
    layer0_outputs(687) <= not (a xor b);
    layer0_outputs(688) <= a or b;
    layer0_outputs(689) <= a xor b;
    layer0_outputs(690) <= a xor b;
    layer0_outputs(691) <= a or b;
    layer0_outputs(692) <= a xor b;
    layer0_outputs(693) <= a xor b;
    layer0_outputs(694) <= a xor b;
    layer0_outputs(695) <= b and not a;
    layer0_outputs(696) <= not (a xor b);
    layer0_outputs(697) <= not (a or b);
    layer0_outputs(698) <= a and b;
    layer0_outputs(699) <= not (a or b);
    layer0_outputs(700) <= not b;
    layer0_outputs(701) <= a and not b;
    layer0_outputs(702) <= not a;
    layer0_outputs(703) <= a;
    layer0_outputs(704) <= a;
    layer0_outputs(705) <= not a;
    layer0_outputs(706) <= not (a or b);
    layer0_outputs(707) <= not (a or b);
    layer0_outputs(708) <= not a or b;
    layer0_outputs(709) <= not (a xor b);
    layer0_outputs(710) <= not b;
    layer0_outputs(711) <= a or b;
    layer0_outputs(712) <= a and not b;
    layer0_outputs(713) <= not a or b;
    layer0_outputs(714) <= not a;
    layer0_outputs(715) <= not (a or b);
    layer0_outputs(716) <= a xor b;
    layer0_outputs(717) <= a or b;
    layer0_outputs(718) <= a or b;
    layer0_outputs(719) <= not (a or b);
    layer0_outputs(720) <= a or b;
    layer0_outputs(721) <= b and not a;
    layer0_outputs(722) <= not b;
    layer0_outputs(723) <= a or b;
    layer0_outputs(724) <= a or b;
    layer0_outputs(725) <= not a or b;
    layer0_outputs(726) <= a and not b;
    layer0_outputs(727) <= b;
    layer0_outputs(728) <= not (a xor b);
    layer0_outputs(729) <= not (a or b);
    layer0_outputs(730) <= not a or b;
    layer0_outputs(731) <= a and b;
    layer0_outputs(732) <= not b;
    layer0_outputs(733) <= b;
    layer0_outputs(734) <= a xor b;
    layer0_outputs(735) <= a or b;
    layer0_outputs(736) <= not b;
    layer0_outputs(737) <= not (a or b);
    layer0_outputs(738) <= not (a or b);
    layer0_outputs(739) <= not a or b;
    layer0_outputs(740) <= b and not a;
    layer0_outputs(741) <= not a;
    layer0_outputs(742) <= not a;
    layer0_outputs(743) <= a or b;
    layer0_outputs(744) <= a;
    layer0_outputs(745) <= a or b;
    layer0_outputs(746) <= '0';
    layer0_outputs(747) <= not (a xor b);
    layer0_outputs(748) <= a and not b;
    layer0_outputs(749) <= '0';
    layer0_outputs(750) <= not (a xor b);
    layer0_outputs(751) <= not a;
    layer0_outputs(752) <= not (a or b);
    layer0_outputs(753) <= not (a xor b);
    layer0_outputs(754) <= a or b;
    layer0_outputs(755) <= not (a or b);
    layer0_outputs(756) <= a;
    layer0_outputs(757) <= b;
    layer0_outputs(758) <= not a;
    layer0_outputs(759) <= not (a or b);
    layer0_outputs(760) <= a;
    layer0_outputs(761) <= b and not a;
    layer0_outputs(762) <= a;
    layer0_outputs(763) <= not (a xor b);
    layer0_outputs(764) <= not (a or b);
    layer0_outputs(765) <= a or b;
    layer0_outputs(766) <= not (a or b);
    layer0_outputs(767) <= a;
    layer0_outputs(768) <= not (a or b);
    layer0_outputs(769) <= b and not a;
    layer0_outputs(770) <= not (a xor b);
    layer0_outputs(771) <= b;
    layer0_outputs(772) <= not (a or b);
    layer0_outputs(773) <= a xor b;
    layer0_outputs(774) <= a xor b;
    layer0_outputs(775) <= a;
    layer0_outputs(776) <= b and not a;
    layer0_outputs(777) <= b;
    layer0_outputs(778) <= not (a or b);
    layer0_outputs(779) <= not (a or b);
    layer0_outputs(780) <= not a or b;
    layer0_outputs(781) <= not a or b;
    layer0_outputs(782) <= not (a or b);
    layer0_outputs(783) <= not (a or b);
    layer0_outputs(784) <= not (a xor b);
    layer0_outputs(785) <= a xor b;
    layer0_outputs(786) <= a xor b;
    layer0_outputs(787) <= not (a xor b);
    layer0_outputs(788) <= not a;
    layer0_outputs(789) <= not b;
    layer0_outputs(790) <= not a or b;
    layer0_outputs(791) <= a or b;
    layer0_outputs(792) <= b and not a;
    layer0_outputs(793) <= not (a xor b);
    layer0_outputs(794) <= a and not b;
    layer0_outputs(795) <= a xor b;
    layer0_outputs(796) <= a xor b;
    layer0_outputs(797) <= not (a or b);
    layer0_outputs(798) <= not (a xor b);
    layer0_outputs(799) <= not a;
    layer0_outputs(800) <= not a or b;
    layer0_outputs(801) <= not (a or b);
    layer0_outputs(802) <= not b;
    layer0_outputs(803) <= a and not b;
    layer0_outputs(804) <= not (a xor b);
    layer0_outputs(805) <= not (a and b);
    layer0_outputs(806) <= not (a or b);
    layer0_outputs(807) <= not (a or b);
    layer0_outputs(808) <= not b;
    layer0_outputs(809) <= a xor b;
    layer0_outputs(810) <= a xor b;
    layer0_outputs(811) <= '0';
    layer0_outputs(812) <= b and not a;
    layer0_outputs(813) <= '0';
    layer0_outputs(814) <= a or b;
    layer0_outputs(815) <= a or b;
    layer0_outputs(816) <= not (a or b);
    layer0_outputs(817) <= b;
    layer0_outputs(818) <= not (a xor b);
    layer0_outputs(819) <= a;
    layer0_outputs(820) <= b;
    layer0_outputs(821) <= a;
    layer0_outputs(822) <= not (a or b);
    layer0_outputs(823) <= b;
    layer0_outputs(824) <= not (a or b);
    layer0_outputs(825) <= not (a and b);
    layer0_outputs(826) <= not (a or b);
    layer0_outputs(827) <= not (a or b);
    layer0_outputs(828) <= not a or b;
    layer0_outputs(829) <= not (a or b);
    layer0_outputs(830) <= not (a xor b);
    layer0_outputs(831) <= b and not a;
    layer0_outputs(832) <= '0';
    layer0_outputs(833) <= not (a xor b);
    layer0_outputs(834) <= b and not a;
    layer0_outputs(835) <= a or b;
    layer0_outputs(836) <= a and not b;
    layer0_outputs(837) <= b and not a;
    layer0_outputs(838) <= not (a xor b);
    layer0_outputs(839) <= not (a xor b);
    layer0_outputs(840) <= not (a and b);
    layer0_outputs(841) <= not (a xor b);
    layer0_outputs(842) <= not b or a;
    layer0_outputs(843) <= '1';
    layer0_outputs(844) <= b and not a;
    layer0_outputs(845) <= not (a or b);
    layer0_outputs(846) <= not (a or b);
    layer0_outputs(847) <= not (a xor b);
    layer0_outputs(848) <= a;
    layer0_outputs(849) <= not (a and b);
    layer0_outputs(850) <= a or b;
    layer0_outputs(851) <= not (a xor b);
    layer0_outputs(852) <= not a;
    layer0_outputs(853) <= not b;
    layer0_outputs(854) <= not b;
    layer0_outputs(855) <= a or b;
    layer0_outputs(856) <= a and not b;
    layer0_outputs(857) <= not (a or b);
    layer0_outputs(858) <= a or b;
    layer0_outputs(859) <= b;
    layer0_outputs(860) <= a or b;
    layer0_outputs(861) <= not b;
    layer0_outputs(862) <= a;
    layer0_outputs(863) <= not (a or b);
    layer0_outputs(864) <= not (a or b);
    layer0_outputs(865) <= not (a and b);
    layer0_outputs(866) <= not (a or b);
    layer0_outputs(867) <= b and not a;
    layer0_outputs(868) <= b;
    layer0_outputs(869) <= a or b;
    layer0_outputs(870) <= a or b;
    layer0_outputs(871) <= a and not b;
    layer0_outputs(872) <= a;
    layer0_outputs(873) <= a and not b;
    layer0_outputs(874) <= a xor b;
    layer0_outputs(875) <= not b;
    layer0_outputs(876) <= a xor b;
    layer0_outputs(877) <= a and not b;
    layer0_outputs(878) <= not b or a;
    layer0_outputs(879) <= not a;
    layer0_outputs(880) <= a xor b;
    layer0_outputs(881) <= a or b;
    layer0_outputs(882) <= a;
    layer0_outputs(883) <= not (a or b);
    layer0_outputs(884) <= a xor b;
    layer0_outputs(885) <= a or b;
    layer0_outputs(886) <= b and not a;
    layer0_outputs(887) <= not a or b;
    layer0_outputs(888) <= a;
    layer0_outputs(889) <= b;
    layer0_outputs(890) <= not b or a;
    layer0_outputs(891) <= not (a xor b);
    layer0_outputs(892) <= a;
    layer0_outputs(893) <= '1';
    layer0_outputs(894) <= a or b;
    layer0_outputs(895) <= a or b;
    layer0_outputs(896) <= a;
    layer0_outputs(897) <= not b or a;
    layer0_outputs(898) <= a and b;
    layer0_outputs(899) <= a or b;
    layer0_outputs(900) <= not (a or b);
    layer0_outputs(901) <= a or b;
    layer0_outputs(902) <= not a;
    layer0_outputs(903) <= a and not b;
    layer0_outputs(904) <= '0';
    layer0_outputs(905) <= not (a or b);
    layer0_outputs(906) <= a and b;
    layer0_outputs(907) <= not a or b;
    layer0_outputs(908) <= not (a or b);
    layer0_outputs(909) <= not (a xor b);
    layer0_outputs(910) <= not (a xor b);
    layer0_outputs(911) <= b;
    layer0_outputs(912) <= not a or b;
    layer0_outputs(913) <= not (a xor b);
    layer0_outputs(914) <= a or b;
    layer0_outputs(915) <= b and not a;
    layer0_outputs(916) <= not (a or b);
    layer0_outputs(917) <= not (a xor b);
    layer0_outputs(918) <= a or b;
    layer0_outputs(919) <= a or b;
    layer0_outputs(920) <= not (a xor b);
    layer0_outputs(921) <= b;
    layer0_outputs(922) <= b and not a;
    layer0_outputs(923) <= a xor b;
    layer0_outputs(924) <= not (a or b);
    layer0_outputs(925) <= not (a or b);
    layer0_outputs(926) <= not b or a;
    layer0_outputs(927) <= not (a xor b);
    layer0_outputs(928) <= not (a or b);
    layer0_outputs(929) <= a;
    layer0_outputs(930) <= b and not a;
    layer0_outputs(931) <= not b or a;
    layer0_outputs(932) <= not (a xor b);
    layer0_outputs(933) <= a and b;
    layer0_outputs(934) <= b;
    layer0_outputs(935) <= a;
    layer0_outputs(936) <= a;
    layer0_outputs(937) <= not (a or b);
    layer0_outputs(938) <= a or b;
    layer0_outputs(939) <= not b or a;
    layer0_outputs(940) <= not b;
    layer0_outputs(941) <= b;
    layer0_outputs(942) <= a xor b;
    layer0_outputs(943) <= a or b;
    layer0_outputs(944) <= not (a or b);
    layer0_outputs(945) <= a xor b;
    layer0_outputs(946) <= '1';
    layer0_outputs(947) <= not b;
    layer0_outputs(948) <= not a or b;
    layer0_outputs(949) <= a or b;
    layer0_outputs(950) <= not a;
    layer0_outputs(951) <= a and not b;
    layer0_outputs(952) <= not a;
    layer0_outputs(953) <= b and not a;
    layer0_outputs(954) <= not (a and b);
    layer0_outputs(955) <= not (a xor b);
    layer0_outputs(956) <= a or b;
    layer0_outputs(957) <= not (a or b);
    layer0_outputs(958) <= not a;
    layer0_outputs(959) <= a or b;
    layer0_outputs(960) <= not a;
    layer0_outputs(961) <= not (a and b);
    layer0_outputs(962) <= not (a or b);
    layer0_outputs(963) <= a or b;
    layer0_outputs(964) <= not a;
    layer0_outputs(965) <= b and not a;
    layer0_outputs(966) <= a;
    layer0_outputs(967) <= a and b;
    layer0_outputs(968) <= not (a or b);
    layer0_outputs(969) <= not b or a;
    layer0_outputs(970) <= not b or a;
    layer0_outputs(971) <= a or b;
    layer0_outputs(972) <= not (a and b);
    layer0_outputs(973) <= not a;
    layer0_outputs(974) <= not b;
    layer0_outputs(975) <= not a;
    layer0_outputs(976) <= not b;
    layer0_outputs(977) <= a or b;
    layer0_outputs(978) <= not b or a;
    layer0_outputs(979) <= not a or b;
    layer0_outputs(980) <= a;
    layer0_outputs(981) <= a xor b;
    layer0_outputs(982) <= b;
    layer0_outputs(983) <= a and not b;
    layer0_outputs(984) <= b and not a;
    layer0_outputs(985) <= a or b;
    layer0_outputs(986) <= a and not b;
    layer0_outputs(987) <= not (a or b);
    layer0_outputs(988) <= a;
    layer0_outputs(989) <= a or b;
    layer0_outputs(990) <= b;
    layer0_outputs(991) <= b;
    layer0_outputs(992) <= not (a or b);
    layer0_outputs(993) <= b;
    layer0_outputs(994) <= not a;
    layer0_outputs(995) <= b;
    layer0_outputs(996) <= not (a and b);
    layer0_outputs(997) <= not b;
    layer0_outputs(998) <= '1';
    layer0_outputs(999) <= a and b;
    layer0_outputs(1000) <= a;
    layer0_outputs(1001) <= not (a or b);
    layer0_outputs(1002) <= '1';
    layer0_outputs(1003) <= not (a or b);
    layer0_outputs(1004) <= a or b;
    layer0_outputs(1005) <= not b;
    layer0_outputs(1006) <= not b or a;
    layer0_outputs(1007) <= a;
    layer0_outputs(1008) <= a or b;
    layer0_outputs(1009) <= not a;
    layer0_outputs(1010) <= a or b;
    layer0_outputs(1011) <= a;
    layer0_outputs(1012) <= not (a or b);
    layer0_outputs(1013) <= not (a xor b);
    layer0_outputs(1014) <= b and not a;
    layer0_outputs(1015) <= not (a and b);
    layer0_outputs(1016) <= a or b;
    layer0_outputs(1017) <= not a or b;
    layer0_outputs(1018) <= not (a or b);
    layer0_outputs(1019) <= not b;
    layer0_outputs(1020) <= a and not b;
    layer0_outputs(1021) <= a;
    layer0_outputs(1022) <= a and not b;
    layer0_outputs(1023) <= not (a or b);
    layer0_outputs(1024) <= not b;
    layer0_outputs(1025) <= a and not b;
    layer0_outputs(1026) <= a;
    layer0_outputs(1027) <= not a or b;
    layer0_outputs(1028) <= a and not b;
    layer0_outputs(1029) <= not b;
    layer0_outputs(1030) <= not a;
    layer0_outputs(1031) <= not a;
    layer0_outputs(1032) <= not (a xor b);
    layer0_outputs(1033) <= a xor b;
    layer0_outputs(1034) <= a or b;
    layer0_outputs(1035) <= a;
    layer0_outputs(1036) <= a or b;
    layer0_outputs(1037) <= a xor b;
    layer0_outputs(1038) <= not (a or b);
    layer0_outputs(1039) <= a or b;
    layer0_outputs(1040) <= b;
    layer0_outputs(1041) <= not (a xor b);
    layer0_outputs(1042) <= a;
    layer0_outputs(1043) <= not (a and b);
    layer0_outputs(1044) <= b;
    layer0_outputs(1045) <= a and not b;
    layer0_outputs(1046) <= not b;
    layer0_outputs(1047) <= a xor b;
    layer0_outputs(1048) <= a and not b;
    layer0_outputs(1049) <= a and not b;
    layer0_outputs(1050) <= '1';
    layer0_outputs(1051) <= not (a xor b);
    layer0_outputs(1052) <= not (a or b);
    layer0_outputs(1053) <= b;
    layer0_outputs(1054) <= b;
    layer0_outputs(1055) <= a and b;
    layer0_outputs(1056) <= not (a or b);
    layer0_outputs(1057) <= not a or b;
    layer0_outputs(1058) <= not (a or b);
    layer0_outputs(1059) <= not a or b;
    layer0_outputs(1060) <= a xor b;
    layer0_outputs(1061) <= a or b;
    layer0_outputs(1062) <= not (a xor b);
    layer0_outputs(1063) <= not (a or b);
    layer0_outputs(1064) <= not (a xor b);
    layer0_outputs(1065) <= not b or a;
    layer0_outputs(1066) <= a and not b;
    layer0_outputs(1067) <= not a or b;
    layer0_outputs(1068) <= a or b;
    layer0_outputs(1069) <= b and not a;
    layer0_outputs(1070) <= a and not b;
    layer0_outputs(1071) <= not b;
    layer0_outputs(1072) <= b and not a;
    layer0_outputs(1073) <= not b or a;
    layer0_outputs(1074) <= a;
    layer0_outputs(1075) <= not (a xor b);
    layer0_outputs(1076) <= not (a or b);
    layer0_outputs(1077) <= a or b;
    layer0_outputs(1078) <= a or b;
    layer0_outputs(1079) <= b and not a;
    layer0_outputs(1080) <= a xor b;
    layer0_outputs(1081) <= not a;
    layer0_outputs(1082) <= not (a or b);
    layer0_outputs(1083) <= b;
    layer0_outputs(1084) <= not (a xor b);
    layer0_outputs(1085) <= not b or a;
    layer0_outputs(1086) <= a;
    layer0_outputs(1087) <= not (a and b);
    layer0_outputs(1088) <= b and not a;
    layer0_outputs(1089) <= not (a and b);
    layer0_outputs(1090) <= '0';
    layer0_outputs(1091) <= not (a xor b);
    layer0_outputs(1092) <= not b or a;
    layer0_outputs(1093) <= b;
    layer0_outputs(1094) <= not (a xor b);
    layer0_outputs(1095) <= a and not b;
    layer0_outputs(1096) <= a xor b;
    layer0_outputs(1097) <= a or b;
    layer0_outputs(1098) <= a or b;
    layer0_outputs(1099) <= not (a or b);
    layer0_outputs(1100) <= not b;
    layer0_outputs(1101) <= a or b;
    layer0_outputs(1102) <= not b;
    layer0_outputs(1103) <= not a or b;
    layer0_outputs(1104) <= a or b;
    layer0_outputs(1105) <= b and not a;
    layer0_outputs(1106) <= not (a xor b);
    layer0_outputs(1107) <= a or b;
    layer0_outputs(1108) <= a xor b;
    layer0_outputs(1109) <= not a;
    layer0_outputs(1110) <= b;
    layer0_outputs(1111) <= not a or b;
    layer0_outputs(1112) <= not a;
    layer0_outputs(1113) <= b;
    layer0_outputs(1114) <= not (a xor b);
    layer0_outputs(1115) <= not a or b;
    layer0_outputs(1116) <= a or b;
    layer0_outputs(1117) <= b;
    layer0_outputs(1118) <= a xor b;
    layer0_outputs(1119) <= not a;
    layer0_outputs(1120) <= b;
    layer0_outputs(1121) <= a and not b;
    layer0_outputs(1122) <= not (a or b);
    layer0_outputs(1123) <= not a or b;
    layer0_outputs(1124) <= not a;
    layer0_outputs(1125) <= a and not b;
    layer0_outputs(1126) <= not b;
    layer0_outputs(1127) <= not (a xor b);
    layer0_outputs(1128) <= not a or b;
    layer0_outputs(1129) <= b and not a;
    layer0_outputs(1130) <= not a;
    layer0_outputs(1131) <= not (a or b);
    layer0_outputs(1132) <= not (a xor b);
    layer0_outputs(1133) <= a or b;
    layer0_outputs(1134) <= b;
    layer0_outputs(1135) <= not b or a;
    layer0_outputs(1136) <= not (a or b);
    layer0_outputs(1137) <= a xor b;
    layer0_outputs(1138) <= a or b;
    layer0_outputs(1139) <= a xor b;
    layer0_outputs(1140) <= not a or b;
    layer0_outputs(1141) <= not (a xor b);
    layer0_outputs(1142) <= a or b;
    layer0_outputs(1143) <= '1';
    layer0_outputs(1144) <= a;
    layer0_outputs(1145) <= b;
    layer0_outputs(1146) <= a or b;
    layer0_outputs(1147) <= a;
    layer0_outputs(1148) <= a xor b;
    layer0_outputs(1149) <= a and b;
    layer0_outputs(1150) <= a and not b;
    layer0_outputs(1151) <= not (a xor b);
    layer0_outputs(1152) <= not (a or b);
    layer0_outputs(1153) <= '0';
    layer0_outputs(1154) <= a or b;
    layer0_outputs(1155) <= not a;
    layer0_outputs(1156) <= a xor b;
    layer0_outputs(1157) <= a or b;
    layer0_outputs(1158) <= not (a or b);
    layer0_outputs(1159) <= not (a xor b);
    layer0_outputs(1160) <= not a;
    layer0_outputs(1161) <= not (a xor b);
    layer0_outputs(1162) <= a and not b;
    layer0_outputs(1163) <= a and not b;
    layer0_outputs(1164) <= b;
    layer0_outputs(1165) <= not (a xor b);
    layer0_outputs(1166) <= not b or a;
    layer0_outputs(1167) <= not a or b;
    layer0_outputs(1168) <= a xor b;
    layer0_outputs(1169) <= not b or a;
    layer0_outputs(1170) <= a;
    layer0_outputs(1171) <= not a;
    layer0_outputs(1172) <= a xor b;
    layer0_outputs(1173) <= a xor b;
    layer0_outputs(1174) <= not b;
    layer0_outputs(1175) <= not (a and b);
    layer0_outputs(1176) <= a or b;
    layer0_outputs(1177) <= not (a or b);
    layer0_outputs(1178) <= a or b;
    layer0_outputs(1179) <= a or b;
    layer0_outputs(1180) <= not b or a;
    layer0_outputs(1181) <= a;
    layer0_outputs(1182) <= not b;
    layer0_outputs(1183) <= not b;
    layer0_outputs(1184) <= not (a or b);
    layer0_outputs(1185) <= b;
    layer0_outputs(1186) <= '0';
    layer0_outputs(1187) <= not b;
    layer0_outputs(1188) <= b and not a;
    layer0_outputs(1189) <= a or b;
    layer0_outputs(1190) <= not (a xor b);
    layer0_outputs(1191) <= a;
    layer0_outputs(1192) <= not a or b;
    layer0_outputs(1193) <= not b;
    layer0_outputs(1194) <= not (a or b);
    layer0_outputs(1195) <= a or b;
    layer0_outputs(1196) <= not b;
    layer0_outputs(1197) <= b;
    layer0_outputs(1198) <= a;
    layer0_outputs(1199) <= a;
    layer0_outputs(1200) <= b;
    layer0_outputs(1201) <= '1';
    layer0_outputs(1202) <= not a or b;
    layer0_outputs(1203) <= not (a xor b);
    layer0_outputs(1204) <= a and b;
    layer0_outputs(1205) <= not a;
    layer0_outputs(1206) <= not (a or b);
    layer0_outputs(1207) <= a and b;
    layer0_outputs(1208) <= a;
    layer0_outputs(1209) <= not (a or b);
    layer0_outputs(1210) <= not b;
    layer0_outputs(1211) <= b and not a;
    layer0_outputs(1212) <= a xor b;
    layer0_outputs(1213) <= not (a or b);
    layer0_outputs(1214) <= b and not a;
    layer0_outputs(1215) <= b;
    layer0_outputs(1216) <= not b;
    layer0_outputs(1217) <= a and b;
    layer0_outputs(1218) <= not (a or b);
    layer0_outputs(1219) <= a xor b;
    layer0_outputs(1220) <= b;
    layer0_outputs(1221) <= b and not a;
    layer0_outputs(1222) <= not (a xor b);
    layer0_outputs(1223) <= not (a or b);
    layer0_outputs(1224) <= not (a or b);
    layer0_outputs(1225) <= not (a and b);
    layer0_outputs(1226) <= not b or a;
    layer0_outputs(1227) <= b;
    layer0_outputs(1228) <= not (a xor b);
    layer0_outputs(1229) <= a and not b;
    layer0_outputs(1230) <= not a;
    layer0_outputs(1231) <= not (a xor b);
    layer0_outputs(1232) <= not (a xor b);
    layer0_outputs(1233) <= not a or b;
    layer0_outputs(1234) <= a or b;
    layer0_outputs(1235) <= not (a xor b);
    layer0_outputs(1236) <= not (a or b);
    layer0_outputs(1237) <= a xor b;
    layer0_outputs(1238) <= a;
    layer0_outputs(1239) <= a and not b;
    layer0_outputs(1240) <= not b or a;
    layer0_outputs(1241) <= a or b;
    layer0_outputs(1242) <= a or b;
    layer0_outputs(1243) <= '1';
    layer0_outputs(1244) <= a xor b;
    layer0_outputs(1245) <= not b;
    layer0_outputs(1246) <= not (a xor b);
    layer0_outputs(1247) <= b;
    layer0_outputs(1248) <= not (a or b);
    layer0_outputs(1249) <= a;
    layer0_outputs(1250) <= not a;
    layer0_outputs(1251) <= a;
    layer0_outputs(1252) <= a;
    layer0_outputs(1253) <= a or b;
    layer0_outputs(1254) <= not (a or b);
    layer0_outputs(1255) <= a;
    layer0_outputs(1256) <= not b or a;
    layer0_outputs(1257) <= '0';
    layer0_outputs(1258) <= not a;
    layer0_outputs(1259) <= not (a or b);
    layer0_outputs(1260) <= a;
    layer0_outputs(1261) <= a;
    layer0_outputs(1262) <= not a;
    layer0_outputs(1263) <= a and b;
    layer0_outputs(1264) <= a xor b;
    layer0_outputs(1265) <= a or b;
    layer0_outputs(1266) <= not a;
    layer0_outputs(1267) <= not a or b;
    layer0_outputs(1268) <= not (a xor b);
    layer0_outputs(1269) <= not b or a;
    layer0_outputs(1270) <= b and not a;
    layer0_outputs(1271) <= not (a xor b);
    layer0_outputs(1272) <= not b or a;
    layer0_outputs(1273) <= not a;
    layer0_outputs(1274) <= not b or a;
    layer0_outputs(1275) <= a;
    layer0_outputs(1276) <= not (a or b);
    layer0_outputs(1277) <= not a;
    layer0_outputs(1278) <= a;
    layer0_outputs(1279) <= not (a and b);
    layer0_outputs(1280) <= not a;
    layer0_outputs(1281) <= not (a xor b);
    layer0_outputs(1282) <= not (a or b);
    layer0_outputs(1283) <= a xor b;
    layer0_outputs(1284) <= a;
    layer0_outputs(1285) <= a or b;
    layer0_outputs(1286) <= not b;
    layer0_outputs(1287) <= not (a and b);
    layer0_outputs(1288) <= not a or b;
    layer0_outputs(1289) <= a xor b;
    layer0_outputs(1290) <= not (a xor b);
    layer0_outputs(1291) <= b and not a;
    layer0_outputs(1292) <= not b;
    layer0_outputs(1293) <= a;
    layer0_outputs(1294) <= b;
    layer0_outputs(1295) <= a or b;
    layer0_outputs(1296) <= not a or b;
    layer0_outputs(1297) <= not a;
    layer0_outputs(1298) <= not a;
    layer0_outputs(1299) <= a and not b;
    layer0_outputs(1300) <= b;
    layer0_outputs(1301) <= not b or a;
    layer0_outputs(1302) <= not (a and b);
    layer0_outputs(1303) <= '0';
    layer0_outputs(1304) <= not (a xor b);
    layer0_outputs(1305) <= b and not a;
    layer0_outputs(1306) <= not (a or b);
    layer0_outputs(1307) <= a or b;
    layer0_outputs(1308) <= b and not a;
    layer0_outputs(1309) <= b and not a;
    layer0_outputs(1310) <= a xor b;
    layer0_outputs(1311) <= not (a and b);
    layer0_outputs(1312) <= a xor b;
    layer0_outputs(1313) <= b and not a;
    layer0_outputs(1314) <= not (a xor b);
    layer0_outputs(1315) <= b;
    layer0_outputs(1316) <= b and not a;
    layer0_outputs(1317) <= not a;
    layer0_outputs(1318) <= a or b;
    layer0_outputs(1319) <= a or b;
    layer0_outputs(1320) <= a or b;
    layer0_outputs(1321) <= not (a xor b);
    layer0_outputs(1322) <= not b or a;
    layer0_outputs(1323) <= b and not a;
    layer0_outputs(1324) <= a or b;
    layer0_outputs(1325) <= a;
    layer0_outputs(1326) <= a and not b;
    layer0_outputs(1327) <= not (a xor b);
    layer0_outputs(1328) <= a xor b;
    layer0_outputs(1329) <= not a or b;
    layer0_outputs(1330) <= a or b;
    layer0_outputs(1331) <= a and not b;
    layer0_outputs(1332) <= not a;
    layer0_outputs(1333) <= b;
    layer0_outputs(1334) <= not (a xor b);
    layer0_outputs(1335) <= a xor b;
    layer0_outputs(1336) <= not (a xor b);
    layer0_outputs(1337) <= a xor b;
    layer0_outputs(1338) <= a and not b;
    layer0_outputs(1339) <= not (a xor b);
    layer0_outputs(1340) <= a or b;
    layer0_outputs(1341) <= not (a or b);
    layer0_outputs(1342) <= a xor b;
    layer0_outputs(1343) <= a and not b;
    layer0_outputs(1344) <= '1';
    layer0_outputs(1345) <= a and not b;
    layer0_outputs(1346) <= a xor b;
    layer0_outputs(1347) <= not b or a;
    layer0_outputs(1348) <= not (a xor b);
    layer0_outputs(1349) <= a;
    layer0_outputs(1350) <= a and not b;
    layer0_outputs(1351) <= a or b;
    layer0_outputs(1352) <= a;
    layer0_outputs(1353) <= not (a xor b);
    layer0_outputs(1354) <= not b;
    layer0_outputs(1355) <= a;
    layer0_outputs(1356) <= not (a xor b);
    layer0_outputs(1357) <= a and b;
    layer0_outputs(1358) <= not b or a;
    layer0_outputs(1359) <= a xor b;
    layer0_outputs(1360) <= not a or b;
    layer0_outputs(1361) <= a xor b;
    layer0_outputs(1362) <= b and not a;
    layer0_outputs(1363) <= a and not b;
    layer0_outputs(1364) <= b and not a;
    layer0_outputs(1365) <= a or b;
    layer0_outputs(1366) <= b and not a;
    layer0_outputs(1367) <= not b;
    layer0_outputs(1368) <= a or b;
    layer0_outputs(1369) <= a xor b;
    layer0_outputs(1370) <= b and not a;
    layer0_outputs(1371) <= not a or b;
    layer0_outputs(1372) <= not b or a;
    layer0_outputs(1373) <= a and not b;
    layer0_outputs(1374) <= a;
    layer0_outputs(1375) <= not (a xor b);
    layer0_outputs(1376) <= not (a or b);
    layer0_outputs(1377) <= a or b;
    layer0_outputs(1378) <= not (a xor b);
    layer0_outputs(1379) <= not (a and b);
    layer0_outputs(1380) <= a or b;
    layer0_outputs(1381) <= a;
    layer0_outputs(1382) <= not b or a;
    layer0_outputs(1383) <= not (a and b);
    layer0_outputs(1384) <= a;
    layer0_outputs(1385) <= a;
    layer0_outputs(1386) <= a or b;
    layer0_outputs(1387) <= a or b;
    layer0_outputs(1388) <= '1';
    layer0_outputs(1389) <= not (a or b);
    layer0_outputs(1390) <= not (a or b);
    layer0_outputs(1391) <= a or b;
    layer0_outputs(1392) <= a;
    layer0_outputs(1393) <= not a or b;
    layer0_outputs(1394) <= a or b;
    layer0_outputs(1395) <= a or b;
    layer0_outputs(1396) <= a or b;
    layer0_outputs(1397) <= not a or b;
    layer0_outputs(1398) <= b and not a;
    layer0_outputs(1399) <= not (a or b);
    layer0_outputs(1400) <= not (a or b);
    layer0_outputs(1401) <= a or b;
    layer0_outputs(1402) <= not (a xor b);
    layer0_outputs(1403) <= not b;
    layer0_outputs(1404) <= a or b;
    layer0_outputs(1405) <= a and not b;
    layer0_outputs(1406) <= a and not b;
    layer0_outputs(1407) <= not (a xor b);
    layer0_outputs(1408) <= not (a or b);
    layer0_outputs(1409) <= not a;
    layer0_outputs(1410) <= a xor b;
    layer0_outputs(1411) <= not b or a;
    layer0_outputs(1412) <= a xor b;
    layer0_outputs(1413) <= not a;
    layer0_outputs(1414) <= '1';
    layer0_outputs(1415) <= a xor b;
    layer0_outputs(1416) <= not b;
    layer0_outputs(1417) <= b;
    layer0_outputs(1418) <= not a or b;
    layer0_outputs(1419) <= not b;
    layer0_outputs(1420) <= not b or a;
    layer0_outputs(1421) <= a and not b;
    layer0_outputs(1422) <= not a or b;
    layer0_outputs(1423) <= not (a or b);
    layer0_outputs(1424) <= a xor b;
    layer0_outputs(1425) <= not (a xor b);
    layer0_outputs(1426) <= b;
    layer0_outputs(1427) <= a xor b;
    layer0_outputs(1428) <= '0';
    layer0_outputs(1429) <= a and b;
    layer0_outputs(1430) <= not (a or b);
    layer0_outputs(1431) <= not b;
    layer0_outputs(1432) <= not b or a;
    layer0_outputs(1433) <= a or b;
    layer0_outputs(1434) <= not (a or b);
    layer0_outputs(1435) <= not a;
    layer0_outputs(1436) <= not (a and b);
    layer0_outputs(1437) <= a or b;
    layer0_outputs(1438) <= b;
    layer0_outputs(1439) <= not a;
    layer0_outputs(1440) <= not a;
    layer0_outputs(1441) <= not (a or b);
    layer0_outputs(1442) <= not b;
    layer0_outputs(1443) <= not a;
    layer0_outputs(1444) <= not a or b;
    layer0_outputs(1445) <= a;
    layer0_outputs(1446) <= a or b;
    layer0_outputs(1447) <= b and not a;
    layer0_outputs(1448) <= not (a and b);
    layer0_outputs(1449) <= not a;
    layer0_outputs(1450) <= not (a xor b);
    layer0_outputs(1451) <= b and not a;
    layer0_outputs(1452) <= a and not b;
    layer0_outputs(1453) <= not b;
    layer0_outputs(1454) <= not b;
    layer0_outputs(1455) <= not (a or b);
    layer0_outputs(1456) <= a xor b;
    layer0_outputs(1457) <= b and not a;
    layer0_outputs(1458) <= not (a or b);
    layer0_outputs(1459) <= b and not a;
    layer0_outputs(1460) <= a and not b;
    layer0_outputs(1461) <= b and not a;
    layer0_outputs(1462) <= a or b;
    layer0_outputs(1463) <= a xor b;
    layer0_outputs(1464) <= not a;
    layer0_outputs(1465) <= not (a xor b);
    layer0_outputs(1466) <= not a;
    layer0_outputs(1467) <= a xor b;
    layer0_outputs(1468) <= a or b;
    layer0_outputs(1469) <= a and not b;
    layer0_outputs(1470) <= a xor b;
    layer0_outputs(1471) <= not a;
    layer0_outputs(1472) <= b and not a;
    layer0_outputs(1473) <= a;
    layer0_outputs(1474) <= '0';
    layer0_outputs(1475) <= not b;
    layer0_outputs(1476) <= a;
    layer0_outputs(1477) <= a or b;
    layer0_outputs(1478) <= a xor b;
    layer0_outputs(1479) <= a or b;
    layer0_outputs(1480) <= a xor b;
    layer0_outputs(1481) <= not a or b;
    layer0_outputs(1482) <= not a or b;
    layer0_outputs(1483) <= not b or a;
    layer0_outputs(1484) <= not (a xor b);
    layer0_outputs(1485) <= a and not b;
    layer0_outputs(1486) <= a;
    layer0_outputs(1487) <= not b or a;
    layer0_outputs(1488) <= not b;
    layer0_outputs(1489) <= not b or a;
    layer0_outputs(1490) <= not b;
    layer0_outputs(1491) <= not b;
    layer0_outputs(1492) <= b and not a;
    layer0_outputs(1493) <= not (a or b);
    layer0_outputs(1494) <= not a or b;
    layer0_outputs(1495) <= b and not a;
    layer0_outputs(1496) <= b;
    layer0_outputs(1497) <= a;
    layer0_outputs(1498) <= b;
    layer0_outputs(1499) <= not (a xor b);
    layer0_outputs(1500) <= a or b;
    layer0_outputs(1501) <= not (a xor b);
    layer0_outputs(1502) <= not (a xor b);
    layer0_outputs(1503) <= b and not a;
    layer0_outputs(1504) <= b and not a;
    layer0_outputs(1505) <= not (a or b);
    layer0_outputs(1506) <= a or b;
    layer0_outputs(1507) <= a xor b;
    layer0_outputs(1508) <= a or b;
    layer0_outputs(1509) <= not b or a;
    layer0_outputs(1510) <= not (a xor b);
    layer0_outputs(1511) <= not b or a;
    layer0_outputs(1512) <= b;
    layer0_outputs(1513) <= a;
    layer0_outputs(1514) <= not (a or b);
    layer0_outputs(1515) <= not (a xor b);
    layer0_outputs(1516) <= not b;
    layer0_outputs(1517) <= not a;
    layer0_outputs(1518) <= not a;
    layer0_outputs(1519) <= a;
    layer0_outputs(1520) <= not b or a;
    layer0_outputs(1521) <= a xor b;
    layer0_outputs(1522) <= not a;
    layer0_outputs(1523) <= a;
    layer0_outputs(1524) <= not a;
    layer0_outputs(1525) <= not b or a;
    layer0_outputs(1526) <= not a;
    layer0_outputs(1527) <= a or b;
    layer0_outputs(1528) <= a;
    layer0_outputs(1529) <= a or b;
    layer0_outputs(1530) <= a or b;
    layer0_outputs(1531) <= not b or a;
    layer0_outputs(1532) <= not (a and b);
    layer0_outputs(1533) <= '0';
    layer0_outputs(1534) <= a and not b;
    layer0_outputs(1535) <= b and not a;
    layer0_outputs(1536) <= not a or b;
    layer0_outputs(1537) <= not b or a;
    layer0_outputs(1538) <= a or b;
    layer0_outputs(1539) <= a or b;
    layer0_outputs(1540) <= not (a or b);
    layer0_outputs(1541) <= not (a or b);
    layer0_outputs(1542) <= not b;
    layer0_outputs(1543) <= a or b;
    layer0_outputs(1544) <= a or b;
    layer0_outputs(1545) <= a or b;
    layer0_outputs(1546) <= a;
    layer0_outputs(1547) <= a and b;
    layer0_outputs(1548) <= '1';
    layer0_outputs(1549) <= a xor b;
    layer0_outputs(1550) <= a and b;
    layer0_outputs(1551) <= a xor b;
    layer0_outputs(1552) <= not (a or b);
    layer0_outputs(1553) <= a xor b;
    layer0_outputs(1554) <= a or b;
    layer0_outputs(1555) <= a and not b;
    layer0_outputs(1556) <= not (a or b);
    layer0_outputs(1557) <= not (a and b);
    layer0_outputs(1558) <= a and not b;
    layer0_outputs(1559) <= not b;
    layer0_outputs(1560) <= a and not b;
    layer0_outputs(1561) <= a or b;
    layer0_outputs(1562) <= a or b;
    layer0_outputs(1563) <= b;
    layer0_outputs(1564) <= a xor b;
    layer0_outputs(1565) <= a xor b;
    layer0_outputs(1566) <= not b or a;
    layer0_outputs(1567) <= '1';
    layer0_outputs(1568) <= not (a or b);
    layer0_outputs(1569) <= a xor b;
    layer0_outputs(1570) <= not (a xor b);
    layer0_outputs(1571) <= not (a or b);
    layer0_outputs(1572) <= not a;
    layer0_outputs(1573) <= not (a or b);
    layer0_outputs(1574) <= b and not a;
    layer0_outputs(1575) <= a or b;
    layer0_outputs(1576) <= a xor b;
    layer0_outputs(1577) <= not (a xor b);
    layer0_outputs(1578) <= not b or a;
    layer0_outputs(1579) <= a;
    layer0_outputs(1580) <= b and not a;
    layer0_outputs(1581) <= a xor b;
    layer0_outputs(1582) <= not a or b;
    layer0_outputs(1583) <= a or b;
    layer0_outputs(1584) <= not (a xor b);
    layer0_outputs(1585) <= a and not b;
    layer0_outputs(1586) <= not b;
    layer0_outputs(1587) <= not a or b;
    layer0_outputs(1588) <= b and not a;
    layer0_outputs(1589) <= a or b;
    layer0_outputs(1590) <= not b;
    layer0_outputs(1591) <= b and not a;
    layer0_outputs(1592) <= '0';
    layer0_outputs(1593) <= not (a or b);
    layer0_outputs(1594) <= not a or b;
    layer0_outputs(1595) <= not b;
    layer0_outputs(1596) <= not a;
    layer0_outputs(1597) <= not (a xor b);
    layer0_outputs(1598) <= a or b;
    layer0_outputs(1599) <= a;
    layer0_outputs(1600) <= a or b;
    layer0_outputs(1601) <= not (a and b);
    layer0_outputs(1602) <= a and not b;
    layer0_outputs(1603) <= a and not b;
    layer0_outputs(1604) <= not (a or b);
    layer0_outputs(1605) <= '1';
    layer0_outputs(1606) <= not b;
    layer0_outputs(1607) <= not b;
    layer0_outputs(1608) <= not (a xor b);
    layer0_outputs(1609) <= a or b;
    layer0_outputs(1610) <= a and b;
    layer0_outputs(1611) <= not a;
    layer0_outputs(1612) <= '1';
    layer0_outputs(1613) <= a and b;
    layer0_outputs(1614) <= not (a xor b);
    layer0_outputs(1615) <= not a or b;
    layer0_outputs(1616) <= not b;
    layer0_outputs(1617) <= a xor b;
    layer0_outputs(1618) <= a;
    layer0_outputs(1619) <= a;
    layer0_outputs(1620) <= not b;
    layer0_outputs(1621) <= not (a or b);
    layer0_outputs(1622) <= not b or a;
    layer0_outputs(1623) <= b;
    layer0_outputs(1624) <= a and b;
    layer0_outputs(1625) <= not (a or b);
    layer0_outputs(1626) <= not a;
    layer0_outputs(1627) <= a;
    layer0_outputs(1628) <= not (a xor b);
    layer0_outputs(1629) <= a and b;
    layer0_outputs(1630) <= b and not a;
    layer0_outputs(1631) <= not (a xor b);
    layer0_outputs(1632) <= a xor b;
    layer0_outputs(1633) <= a xor b;
    layer0_outputs(1634) <= a xor b;
    layer0_outputs(1635) <= a;
    layer0_outputs(1636) <= not b;
    layer0_outputs(1637) <= not (a or b);
    layer0_outputs(1638) <= not b or a;
    layer0_outputs(1639) <= not b;
    layer0_outputs(1640) <= a xor b;
    layer0_outputs(1641) <= not b or a;
    layer0_outputs(1642) <= a and not b;
    layer0_outputs(1643) <= not a or b;
    layer0_outputs(1644) <= a and not b;
    layer0_outputs(1645) <= a xor b;
    layer0_outputs(1646) <= a or b;
    layer0_outputs(1647) <= not (a or b);
    layer0_outputs(1648) <= a xor b;
    layer0_outputs(1649) <= not (a xor b);
    layer0_outputs(1650) <= not b or a;
    layer0_outputs(1651) <= not (a xor b);
    layer0_outputs(1652) <= not (a xor b);
    layer0_outputs(1653) <= a;
    layer0_outputs(1654) <= not (a or b);
    layer0_outputs(1655) <= '1';
    layer0_outputs(1656) <= a;
    layer0_outputs(1657) <= not b or a;
    layer0_outputs(1658) <= b and not a;
    layer0_outputs(1659) <= b and not a;
    layer0_outputs(1660) <= a or b;
    layer0_outputs(1661) <= a or b;
    layer0_outputs(1662) <= a xor b;
    layer0_outputs(1663) <= not (a or b);
    layer0_outputs(1664) <= a xor b;
    layer0_outputs(1665) <= not (a or b);
    layer0_outputs(1666) <= not a;
    layer0_outputs(1667) <= not (a or b);
    layer0_outputs(1668) <= not (a and b);
    layer0_outputs(1669) <= not (a xor b);
    layer0_outputs(1670) <= a or b;
    layer0_outputs(1671) <= a or b;
    layer0_outputs(1672) <= a or b;
    layer0_outputs(1673) <= not (a or b);
    layer0_outputs(1674) <= not (a or b);
    layer0_outputs(1675) <= not (a xor b);
    layer0_outputs(1676) <= not (a or b);
    layer0_outputs(1677) <= b;
    layer0_outputs(1678) <= a;
    layer0_outputs(1679) <= not (a xor b);
    layer0_outputs(1680) <= a and not b;
    layer0_outputs(1681) <= '1';
    layer0_outputs(1682) <= b and not a;
    layer0_outputs(1683) <= not (a and b);
    layer0_outputs(1684) <= a or b;
    layer0_outputs(1685) <= not b or a;
    layer0_outputs(1686) <= not (a xor b);
    layer0_outputs(1687) <= a or b;
    layer0_outputs(1688) <= a xor b;
    layer0_outputs(1689) <= a or b;
    layer0_outputs(1690) <= not b;
    layer0_outputs(1691) <= a or b;
    layer0_outputs(1692) <= b and not a;
    layer0_outputs(1693) <= a and not b;
    layer0_outputs(1694) <= a and not b;
    layer0_outputs(1695) <= b and not a;
    layer0_outputs(1696) <= a;
    layer0_outputs(1697) <= not a or b;
    layer0_outputs(1698) <= a or b;
    layer0_outputs(1699) <= not (a xor b);
    layer0_outputs(1700) <= b and not a;
    layer0_outputs(1701) <= not b;
    layer0_outputs(1702) <= b;
    layer0_outputs(1703) <= not b or a;
    layer0_outputs(1704) <= b and not a;
    layer0_outputs(1705) <= a and not b;
    layer0_outputs(1706) <= a or b;
    layer0_outputs(1707) <= b and not a;
    layer0_outputs(1708) <= not (a xor b);
    layer0_outputs(1709) <= b and not a;
    layer0_outputs(1710) <= not a or b;
    layer0_outputs(1711) <= not a or b;
    layer0_outputs(1712) <= a and not b;
    layer0_outputs(1713) <= a;
    layer0_outputs(1714) <= not (a or b);
    layer0_outputs(1715) <= not a or b;
    layer0_outputs(1716) <= a and not b;
    layer0_outputs(1717) <= not (a or b);
    layer0_outputs(1718) <= a xor b;
    layer0_outputs(1719) <= not a or b;
    layer0_outputs(1720) <= not (a xor b);
    layer0_outputs(1721) <= not (a and b);
    layer0_outputs(1722) <= b and not a;
    layer0_outputs(1723) <= a and not b;
    layer0_outputs(1724) <= b and not a;
    layer0_outputs(1725) <= a;
    layer0_outputs(1726) <= a;
    layer0_outputs(1727) <= b;
    layer0_outputs(1728) <= not (a or b);
    layer0_outputs(1729) <= not a;
    layer0_outputs(1730) <= not a;
    layer0_outputs(1731) <= a xor b;
    layer0_outputs(1732) <= not a;
    layer0_outputs(1733) <= not b or a;
    layer0_outputs(1734) <= a xor b;
    layer0_outputs(1735) <= not (a xor b);
    layer0_outputs(1736) <= not (a xor b);
    layer0_outputs(1737) <= a;
    layer0_outputs(1738) <= not b or a;
    layer0_outputs(1739) <= not (a and b);
    layer0_outputs(1740) <= a or b;
    layer0_outputs(1741) <= not (a or b);
    layer0_outputs(1742) <= a or b;
    layer0_outputs(1743) <= not (a or b);
    layer0_outputs(1744) <= '1';
    layer0_outputs(1745) <= not a;
    layer0_outputs(1746) <= a xor b;
    layer0_outputs(1747) <= a or b;
    layer0_outputs(1748) <= b and not a;
    layer0_outputs(1749) <= a or b;
    layer0_outputs(1750) <= a xor b;
    layer0_outputs(1751) <= b and not a;
    layer0_outputs(1752) <= b and not a;
    layer0_outputs(1753) <= not (a or b);
    layer0_outputs(1754) <= not (a or b);
    layer0_outputs(1755) <= a and not b;
    layer0_outputs(1756) <= not b or a;
    layer0_outputs(1757) <= not (a or b);
    layer0_outputs(1758) <= b;
    layer0_outputs(1759) <= b;
    layer0_outputs(1760) <= not (a xor b);
    layer0_outputs(1761) <= not (a or b);
    layer0_outputs(1762) <= b and not a;
    layer0_outputs(1763) <= a xor b;
    layer0_outputs(1764) <= b;
    layer0_outputs(1765) <= not a;
    layer0_outputs(1766) <= not (a xor b);
    layer0_outputs(1767) <= not b or a;
    layer0_outputs(1768) <= not b or a;
    layer0_outputs(1769) <= not a or b;
    layer0_outputs(1770) <= a and not b;
    layer0_outputs(1771) <= a and b;
    layer0_outputs(1772) <= not (a xor b);
    layer0_outputs(1773) <= not (a or b);
    layer0_outputs(1774) <= not (a or b);
    layer0_outputs(1775) <= b and not a;
    layer0_outputs(1776) <= b and not a;
    layer0_outputs(1777) <= a xor b;
    layer0_outputs(1778) <= not (a or b);
    layer0_outputs(1779) <= not (a xor b);
    layer0_outputs(1780) <= not (a or b);
    layer0_outputs(1781) <= not a;
    layer0_outputs(1782) <= not a or b;
    layer0_outputs(1783) <= not (a xor b);
    layer0_outputs(1784) <= a or b;
    layer0_outputs(1785) <= not a;
    layer0_outputs(1786) <= not (a or b);
    layer0_outputs(1787) <= not (a xor b);
    layer0_outputs(1788) <= a;
    layer0_outputs(1789) <= a and b;
    layer0_outputs(1790) <= not a;
    layer0_outputs(1791) <= not b or a;
    layer0_outputs(1792) <= '1';
    layer0_outputs(1793) <= a;
    layer0_outputs(1794) <= not (a xor b);
    layer0_outputs(1795) <= b and not a;
    layer0_outputs(1796) <= a;
    layer0_outputs(1797) <= a or b;
    layer0_outputs(1798) <= a or b;
    layer0_outputs(1799) <= not b or a;
    layer0_outputs(1800) <= b;
    layer0_outputs(1801) <= a xor b;
    layer0_outputs(1802) <= not a;
    layer0_outputs(1803) <= b;
    layer0_outputs(1804) <= '1';
    layer0_outputs(1805) <= not (a and b);
    layer0_outputs(1806) <= not (a xor b);
    layer0_outputs(1807) <= a;
    layer0_outputs(1808) <= not b;
    layer0_outputs(1809) <= not b or a;
    layer0_outputs(1810) <= a xor b;
    layer0_outputs(1811) <= not b or a;
    layer0_outputs(1812) <= a or b;
    layer0_outputs(1813) <= not (a or b);
    layer0_outputs(1814) <= a xor b;
    layer0_outputs(1815) <= not b;
    layer0_outputs(1816) <= not a;
    layer0_outputs(1817) <= not (a or b);
    layer0_outputs(1818) <= a;
    layer0_outputs(1819) <= not (a xor b);
    layer0_outputs(1820) <= not (a xor b);
    layer0_outputs(1821) <= a xor b;
    layer0_outputs(1822) <= b;
    layer0_outputs(1823) <= b;
    layer0_outputs(1824) <= not b or a;
    layer0_outputs(1825) <= not (a or b);
    layer0_outputs(1826) <= a and not b;
    layer0_outputs(1827) <= a or b;
    layer0_outputs(1828) <= not (a xor b);
    layer0_outputs(1829) <= not (a xor b);
    layer0_outputs(1830) <= not b;
    layer0_outputs(1831) <= not a or b;
    layer0_outputs(1832) <= a xor b;
    layer0_outputs(1833) <= a or b;
    layer0_outputs(1834) <= not (a or b);
    layer0_outputs(1835) <= b;
    layer0_outputs(1836) <= b and not a;
    layer0_outputs(1837) <= a xor b;
    layer0_outputs(1838) <= b and not a;
    layer0_outputs(1839) <= not (a and b);
    layer0_outputs(1840) <= not b;
    layer0_outputs(1841) <= a or b;
    layer0_outputs(1842) <= not (a or b);
    layer0_outputs(1843) <= a or b;
    layer0_outputs(1844) <= b and not a;
    layer0_outputs(1845) <= a xor b;
    layer0_outputs(1846) <= not a;
    layer0_outputs(1847) <= a xor b;
    layer0_outputs(1848) <= a;
    layer0_outputs(1849) <= a;
    layer0_outputs(1850) <= a or b;
    layer0_outputs(1851) <= b;
    layer0_outputs(1852) <= a xor b;
    layer0_outputs(1853) <= a and not b;
    layer0_outputs(1854) <= b;
    layer0_outputs(1855) <= a or b;
    layer0_outputs(1856) <= not b or a;
    layer0_outputs(1857) <= a and not b;
    layer0_outputs(1858) <= b and not a;
    layer0_outputs(1859) <= not (a or b);
    layer0_outputs(1860) <= not b or a;
    layer0_outputs(1861) <= a or b;
    layer0_outputs(1862) <= not a;
    layer0_outputs(1863) <= not b;
    layer0_outputs(1864) <= not a or b;
    layer0_outputs(1865) <= not (a xor b);
    layer0_outputs(1866) <= not a;
    layer0_outputs(1867) <= a xor b;
    layer0_outputs(1868) <= a and not b;
    layer0_outputs(1869) <= not (a xor b);
    layer0_outputs(1870) <= not b;
    layer0_outputs(1871) <= not (a xor b);
    layer0_outputs(1872) <= a;
    layer0_outputs(1873) <= a xor b;
    layer0_outputs(1874) <= not b;
    layer0_outputs(1875) <= not b;
    layer0_outputs(1876) <= b;
    layer0_outputs(1877) <= not (a or b);
    layer0_outputs(1878) <= a xor b;
    layer0_outputs(1879) <= not b;
    layer0_outputs(1880) <= a and not b;
    layer0_outputs(1881) <= a or b;
    layer0_outputs(1882) <= a;
    layer0_outputs(1883) <= b;
    layer0_outputs(1884) <= not b or a;
    layer0_outputs(1885) <= not (a xor b);
    layer0_outputs(1886) <= '0';
    layer0_outputs(1887) <= not a or b;
    layer0_outputs(1888) <= not a;
    layer0_outputs(1889) <= a xor b;
    layer0_outputs(1890) <= a xor b;
    layer0_outputs(1891) <= not b or a;
    layer0_outputs(1892) <= not (a or b);
    layer0_outputs(1893) <= a or b;
    layer0_outputs(1894) <= '1';
    layer0_outputs(1895) <= not b;
    layer0_outputs(1896) <= a xor b;
    layer0_outputs(1897) <= not b;
    layer0_outputs(1898) <= a or b;
    layer0_outputs(1899) <= not a;
    layer0_outputs(1900) <= b;
    layer0_outputs(1901) <= b;
    layer0_outputs(1902) <= a or b;
    layer0_outputs(1903) <= not (a or b);
    layer0_outputs(1904) <= not (a and b);
    layer0_outputs(1905) <= not (a and b);
    layer0_outputs(1906) <= b and not a;
    layer0_outputs(1907) <= a and not b;
    layer0_outputs(1908) <= a xor b;
    layer0_outputs(1909) <= b and not a;
    layer0_outputs(1910) <= b;
    layer0_outputs(1911) <= not (a or b);
    layer0_outputs(1912) <= not b;
    layer0_outputs(1913) <= a;
    layer0_outputs(1914) <= b;
    layer0_outputs(1915) <= not (a or b);
    layer0_outputs(1916) <= a and not b;
    layer0_outputs(1917) <= not (a or b);
    layer0_outputs(1918) <= b;
    layer0_outputs(1919) <= b and not a;
    layer0_outputs(1920) <= not b or a;
    layer0_outputs(1921) <= not b or a;
    layer0_outputs(1922) <= a xor b;
    layer0_outputs(1923) <= not (a xor b);
    layer0_outputs(1924) <= not b or a;
    layer0_outputs(1925) <= not b;
    layer0_outputs(1926) <= b and not a;
    layer0_outputs(1927) <= a and b;
    layer0_outputs(1928) <= a xor b;
    layer0_outputs(1929) <= a and not b;
    layer0_outputs(1930) <= not (a xor b);
    layer0_outputs(1931) <= b;
    layer0_outputs(1932) <= a xor b;
    layer0_outputs(1933) <= a or b;
    layer0_outputs(1934) <= not (a or b);
    layer0_outputs(1935) <= not (a xor b);
    layer0_outputs(1936) <= a or b;
    layer0_outputs(1937) <= a or b;
    layer0_outputs(1938) <= not (a xor b);
    layer0_outputs(1939) <= not b;
    layer0_outputs(1940) <= b;
    layer0_outputs(1941) <= not b;
    layer0_outputs(1942) <= not b or a;
    layer0_outputs(1943) <= not a or b;
    layer0_outputs(1944) <= not (a or b);
    layer0_outputs(1945) <= not a or b;
    layer0_outputs(1946) <= not b;
    layer0_outputs(1947) <= a or b;
    layer0_outputs(1948) <= not (a or b);
    layer0_outputs(1949) <= not a or b;
    layer0_outputs(1950) <= a and b;
    layer0_outputs(1951) <= not (a or b);
    layer0_outputs(1952) <= a;
    layer0_outputs(1953) <= a xor b;
    layer0_outputs(1954) <= not a;
    layer0_outputs(1955) <= not b;
    layer0_outputs(1956) <= not (a and b);
    layer0_outputs(1957) <= a and not b;
    layer0_outputs(1958) <= a and not b;
    layer0_outputs(1959) <= a;
    layer0_outputs(1960) <= '0';
    layer0_outputs(1961) <= a or b;
    layer0_outputs(1962) <= a or b;
    layer0_outputs(1963) <= not (a or b);
    layer0_outputs(1964) <= not b;
    layer0_outputs(1965) <= a;
    layer0_outputs(1966) <= not (a xor b);
    layer0_outputs(1967) <= not b or a;
    layer0_outputs(1968) <= not a or b;
    layer0_outputs(1969) <= '1';
    layer0_outputs(1970) <= not b or a;
    layer0_outputs(1971) <= a;
    layer0_outputs(1972) <= not (a xor b);
    layer0_outputs(1973) <= a xor b;
    layer0_outputs(1974) <= not (a xor b);
    layer0_outputs(1975) <= not b or a;
    layer0_outputs(1976) <= a xor b;
    layer0_outputs(1977) <= a or b;
    layer0_outputs(1978) <= a and not b;
    layer0_outputs(1979) <= not a or b;
    layer0_outputs(1980) <= a xor b;
    layer0_outputs(1981) <= not a or b;
    layer0_outputs(1982) <= not (a or b);
    layer0_outputs(1983) <= a xor b;
    layer0_outputs(1984) <= '1';
    layer0_outputs(1985) <= not (a and b);
    layer0_outputs(1986) <= a and not b;
    layer0_outputs(1987) <= not b or a;
    layer0_outputs(1988) <= b and not a;
    layer0_outputs(1989) <= not (a or b);
    layer0_outputs(1990) <= '1';
    layer0_outputs(1991) <= a;
    layer0_outputs(1992) <= b;
    layer0_outputs(1993) <= not (a xor b);
    layer0_outputs(1994) <= not a or b;
    layer0_outputs(1995) <= not b or a;
    layer0_outputs(1996) <= b;
    layer0_outputs(1997) <= a or b;
    layer0_outputs(1998) <= not (a or b);
    layer0_outputs(1999) <= b;
    layer0_outputs(2000) <= not b;
    layer0_outputs(2001) <= a or b;
    layer0_outputs(2002) <= not (a xor b);
    layer0_outputs(2003) <= not a or b;
    layer0_outputs(2004) <= a or b;
    layer0_outputs(2005) <= not b or a;
    layer0_outputs(2006) <= not b or a;
    layer0_outputs(2007) <= not (a and b);
    layer0_outputs(2008) <= a or b;
    layer0_outputs(2009) <= a or b;
    layer0_outputs(2010) <= a and b;
    layer0_outputs(2011) <= b and not a;
    layer0_outputs(2012) <= not (a or b);
    layer0_outputs(2013) <= not (a xor b);
    layer0_outputs(2014) <= a xor b;
    layer0_outputs(2015) <= '0';
    layer0_outputs(2016) <= not (a xor b);
    layer0_outputs(2017) <= b and not a;
    layer0_outputs(2018) <= a and not b;
    layer0_outputs(2019) <= not b;
    layer0_outputs(2020) <= a or b;
    layer0_outputs(2021) <= a;
    layer0_outputs(2022) <= not (a or b);
    layer0_outputs(2023) <= a and not b;
    layer0_outputs(2024) <= not (a xor b);
    layer0_outputs(2025) <= not a;
    layer0_outputs(2026) <= not a or b;
    layer0_outputs(2027) <= b and not a;
    layer0_outputs(2028) <= not b;
    layer0_outputs(2029) <= a xor b;
    layer0_outputs(2030) <= a and not b;
    layer0_outputs(2031) <= not (a or b);
    layer0_outputs(2032) <= a;
    layer0_outputs(2033) <= a and b;
    layer0_outputs(2034) <= not (a or b);
    layer0_outputs(2035) <= not a;
    layer0_outputs(2036) <= b and not a;
    layer0_outputs(2037) <= b;
    layer0_outputs(2038) <= a or b;
    layer0_outputs(2039) <= a;
    layer0_outputs(2040) <= not a or b;
    layer0_outputs(2041) <= not (a xor b);
    layer0_outputs(2042) <= not (a xor b);
    layer0_outputs(2043) <= not (a or b);
    layer0_outputs(2044) <= a;
    layer0_outputs(2045) <= not (a xor b);
    layer0_outputs(2046) <= b and not a;
    layer0_outputs(2047) <= not b or a;
    layer0_outputs(2048) <= not (a or b);
    layer0_outputs(2049) <= not (a xor b);
    layer0_outputs(2050) <= not (a xor b);
    layer0_outputs(2051) <= not b;
    layer0_outputs(2052) <= a;
    layer0_outputs(2053) <= a and not b;
    layer0_outputs(2054) <= not (a or b);
    layer0_outputs(2055) <= b;
    layer0_outputs(2056) <= not (a or b);
    layer0_outputs(2057) <= a and not b;
    layer0_outputs(2058) <= b and not a;
    layer0_outputs(2059) <= a;
    layer0_outputs(2060) <= not a;
    layer0_outputs(2061) <= a;
    layer0_outputs(2062) <= a and not b;
    layer0_outputs(2063) <= b and not a;
    layer0_outputs(2064) <= b and not a;
    layer0_outputs(2065) <= b;
    layer0_outputs(2066) <= a xor b;
    layer0_outputs(2067) <= a or b;
    layer0_outputs(2068) <= a and not b;
    layer0_outputs(2069) <= not a or b;
    layer0_outputs(2070) <= not (a xor b);
    layer0_outputs(2071) <= not a or b;
    layer0_outputs(2072) <= a xor b;
    layer0_outputs(2073) <= b;
    layer0_outputs(2074) <= a or b;
    layer0_outputs(2075) <= not (a or b);
    layer0_outputs(2076) <= not (a xor b);
    layer0_outputs(2077) <= a and not b;
    layer0_outputs(2078) <= a xor b;
    layer0_outputs(2079) <= b and not a;
    layer0_outputs(2080) <= b;
    layer0_outputs(2081) <= not (a or b);
    layer0_outputs(2082) <= a or b;
    layer0_outputs(2083) <= a and not b;
    layer0_outputs(2084) <= a and not b;
    layer0_outputs(2085) <= not (a or b);
    layer0_outputs(2086) <= not (a or b);
    layer0_outputs(2087) <= b and not a;
    layer0_outputs(2088) <= not a;
    layer0_outputs(2089) <= not (a xor b);
    layer0_outputs(2090) <= not a;
    layer0_outputs(2091) <= a;
    layer0_outputs(2092) <= a or b;
    layer0_outputs(2093) <= b and not a;
    layer0_outputs(2094) <= not (a xor b);
    layer0_outputs(2095) <= not a or b;
    layer0_outputs(2096) <= a or b;
    layer0_outputs(2097) <= b and not a;
    layer0_outputs(2098) <= a;
    layer0_outputs(2099) <= not (a or b);
    layer0_outputs(2100) <= not a or b;
    layer0_outputs(2101) <= not (a or b);
    layer0_outputs(2102) <= a xor b;
    layer0_outputs(2103) <= not a;
    layer0_outputs(2104) <= a or b;
    layer0_outputs(2105) <= a and not b;
    layer0_outputs(2106) <= not a or b;
    layer0_outputs(2107) <= a and not b;
    layer0_outputs(2108) <= a xor b;
    layer0_outputs(2109) <= not a;
    layer0_outputs(2110) <= a and not b;
    layer0_outputs(2111) <= not b or a;
    layer0_outputs(2112) <= a xor b;
    layer0_outputs(2113) <= '0';
    layer0_outputs(2114) <= not b;
    layer0_outputs(2115) <= not (a or b);
    layer0_outputs(2116) <= a or b;
    layer0_outputs(2117) <= a xor b;
    layer0_outputs(2118) <= a or b;
    layer0_outputs(2119) <= not a or b;
    layer0_outputs(2120) <= a xor b;
    layer0_outputs(2121) <= a;
    layer0_outputs(2122) <= a;
    layer0_outputs(2123) <= not (a and b);
    layer0_outputs(2124) <= a;
    layer0_outputs(2125) <= a and not b;
    layer0_outputs(2126) <= a or b;
    layer0_outputs(2127) <= not (a xor b);
    layer0_outputs(2128) <= b;
    layer0_outputs(2129) <= a or b;
    layer0_outputs(2130) <= b and not a;
    layer0_outputs(2131) <= b;
    layer0_outputs(2132) <= not (a xor b);
    layer0_outputs(2133) <= not a or b;
    layer0_outputs(2134) <= a or b;
    layer0_outputs(2135) <= not b or a;
    layer0_outputs(2136) <= b and not a;
    layer0_outputs(2137) <= not (a or b);
    layer0_outputs(2138) <= not (a or b);
    layer0_outputs(2139) <= a and not b;
    layer0_outputs(2140) <= b;
    layer0_outputs(2141) <= a xor b;
    layer0_outputs(2142) <= a and not b;
    layer0_outputs(2143) <= a or b;
    layer0_outputs(2144) <= a and b;
    layer0_outputs(2145) <= not (a xor b);
    layer0_outputs(2146) <= b and not a;
    layer0_outputs(2147) <= not a;
    layer0_outputs(2148) <= a or b;
    layer0_outputs(2149) <= a and not b;
    layer0_outputs(2150) <= a;
    layer0_outputs(2151) <= a or b;
    layer0_outputs(2152) <= a and b;
    layer0_outputs(2153) <= not b or a;
    layer0_outputs(2154) <= a and not b;
    layer0_outputs(2155) <= a;
    layer0_outputs(2156) <= not b or a;
    layer0_outputs(2157) <= not a;
    layer0_outputs(2158) <= not a or b;
    layer0_outputs(2159) <= not (a or b);
    layer0_outputs(2160) <= not a or b;
    layer0_outputs(2161) <= not a;
    layer0_outputs(2162) <= a or b;
    layer0_outputs(2163) <= not (a xor b);
    layer0_outputs(2164) <= a;
    layer0_outputs(2165) <= a or b;
    layer0_outputs(2166) <= not (a xor b);
    layer0_outputs(2167) <= not b or a;
    layer0_outputs(2168) <= not (a xor b);
    layer0_outputs(2169) <= a or b;
    layer0_outputs(2170) <= a;
    layer0_outputs(2171) <= a or b;
    layer0_outputs(2172) <= b and not a;
    layer0_outputs(2173) <= a or b;
    layer0_outputs(2174) <= not (a xor b);
    layer0_outputs(2175) <= not (a or b);
    layer0_outputs(2176) <= a or b;
    layer0_outputs(2177) <= a;
    layer0_outputs(2178) <= a xor b;
    layer0_outputs(2179) <= not (a and b);
    layer0_outputs(2180) <= a;
    layer0_outputs(2181) <= b and not a;
    layer0_outputs(2182) <= not (a xor b);
    layer0_outputs(2183) <= '1';
    layer0_outputs(2184) <= not (a xor b);
    layer0_outputs(2185) <= not b or a;
    layer0_outputs(2186) <= a and b;
    layer0_outputs(2187) <= a;
    layer0_outputs(2188) <= b and not a;
    layer0_outputs(2189) <= a and not b;
    layer0_outputs(2190) <= a xor b;
    layer0_outputs(2191) <= not b or a;
    layer0_outputs(2192) <= a or b;
    layer0_outputs(2193) <= not a or b;
    layer0_outputs(2194) <= not (a or b);
    layer0_outputs(2195) <= a xor b;
    layer0_outputs(2196) <= not (a xor b);
    layer0_outputs(2197) <= not a or b;
    layer0_outputs(2198) <= b;
    layer0_outputs(2199) <= a or b;
    layer0_outputs(2200) <= a and b;
    layer0_outputs(2201) <= not (a xor b);
    layer0_outputs(2202) <= a xor b;
    layer0_outputs(2203) <= a xor b;
    layer0_outputs(2204) <= a or b;
    layer0_outputs(2205) <= '1';
    layer0_outputs(2206) <= a xor b;
    layer0_outputs(2207) <= a or b;
    layer0_outputs(2208) <= not a or b;
    layer0_outputs(2209) <= a;
    layer0_outputs(2210) <= not (a or b);
    layer0_outputs(2211) <= b;
    layer0_outputs(2212) <= a xor b;
    layer0_outputs(2213) <= not (a xor b);
    layer0_outputs(2214) <= not (a or b);
    layer0_outputs(2215) <= a or b;
    layer0_outputs(2216) <= not (a xor b);
    layer0_outputs(2217) <= not (a or b);
    layer0_outputs(2218) <= not (a xor b);
    layer0_outputs(2219) <= a and not b;
    layer0_outputs(2220) <= not b or a;
    layer0_outputs(2221) <= not (a xor b);
    layer0_outputs(2222) <= a;
    layer0_outputs(2223) <= not (a or b);
    layer0_outputs(2224) <= a or b;
    layer0_outputs(2225) <= b;
    layer0_outputs(2226) <= a xor b;
    layer0_outputs(2227) <= not (a or b);
    layer0_outputs(2228) <= not (a or b);
    layer0_outputs(2229) <= a xor b;
    layer0_outputs(2230) <= a xor b;
    layer0_outputs(2231) <= a and not b;
    layer0_outputs(2232) <= not (a or b);
    layer0_outputs(2233) <= a and not b;
    layer0_outputs(2234) <= not b or a;
    layer0_outputs(2235) <= not (a xor b);
    layer0_outputs(2236) <= not (a or b);
    layer0_outputs(2237) <= not b or a;
    layer0_outputs(2238) <= not a or b;
    layer0_outputs(2239) <= a or b;
    layer0_outputs(2240) <= a;
    layer0_outputs(2241) <= a or b;
    layer0_outputs(2242) <= not a or b;
    layer0_outputs(2243) <= not (a xor b);
    layer0_outputs(2244) <= a or b;
    layer0_outputs(2245) <= not (a xor b);
    layer0_outputs(2246) <= not b or a;
    layer0_outputs(2247) <= b;
    layer0_outputs(2248) <= not (a or b);
    layer0_outputs(2249) <= b and not a;
    layer0_outputs(2250) <= not (a or b);
    layer0_outputs(2251) <= not (a and b);
    layer0_outputs(2252) <= a xor b;
    layer0_outputs(2253) <= a;
    layer0_outputs(2254) <= not b;
    layer0_outputs(2255) <= a or b;
    layer0_outputs(2256) <= not (a and b);
    layer0_outputs(2257) <= not a or b;
    layer0_outputs(2258) <= b and not a;
    layer0_outputs(2259) <= not (a xor b);
    layer0_outputs(2260) <= not b;
    layer0_outputs(2261) <= not (a and b);
    layer0_outputs(2262) <= not a;
    layer0_outputs(2263) <= b and not a;
    layer0_outputs(2264) <= not b;
    layer0_outputs(2265) <= a or b;
    layer0_outputs(2266) <= not (a xor b);
    layer0_outputs(2267) <= a xor b;
    layer0_outputs(2268) <= not a or b;
    layer0_outputs(2269) <= a xor b;
    layer0_outputs(2270) <= not b;
    layer0_outputs(2271) <= a xor b;
    layer0_outputs(2272) <= not (a xor b);
    layer0_outputs(2273) <= not a;
    layer0_outputs(2274) <= b and not a;
    layer0_outputs(2275) <= a xor b;
    layer0_outputs(2276) <= not b or a;
    layer0_outputs(2277) <= '0';
    layer0_outputs(2278) <= b;
    layer0_outputs(2279) <= not (a or b);
    layer0_outputs(2280) <= a xor b;
    layer0_outputs(2281) <= not a or b;
    layer0_outputs(2282) <= not (a or b);
    layer0_outputs(2283) <= not a;
    layer0_outputs(2284) <= a or b;
    layer0_outputs(2285) <= not (a xor b);
    layer0_outputs(2286) <= not a;
    layer0_outputs(2287) <= not a;
    layer0_outputs(2288) <= a or b;
    layer0_outputs(2289) <= not a;
    layer0_outputs(2290) <= not b;
    layer0_outputs(2291) <= a;
    layer0_outputs(2292) <= not (a xor b);
    layer0_outputs(2293) <= not b or a;
    layer0_outputs(2294) <= a or b;
    layer0_outputs(2295) <= a or b;
    layer0_outputs(2296) <= '0';
    layer0_outputs(2297) <= a;
    layer0_outputs(2298) <= a or b;
    layer0_outputs(2299) <= a and not b;
    layer0_outputs(2300) <= not a;
    layer0_outputs(2301) <= b;
    layer0_outputs(2302) <= a or b;
    layer0_outputs(2303) <= not b or a;
    layer0_outputs(2304) <= not a;
    layer0_outputs(2305) <= b and not a;
    layer0_outputs(2306) <= a xor b;
    layer0_outputs(2307) <= not a;
    layer0_outputs(2308) <= not a or b;
    layer0_outputs(2309) <= '1';
    layer0_outputs(2310) <= not (a or b);
    layer0_outputs(2311) <= not (a xor b);
    layer0_outputs(2312) <= a or b;
    layer0_outputs(2313) <= b;
    layer0_outputs(2314) <= a and not b;
    layer0_outputs(2315) <= not a;
    layer0_outputs(2316) <= a and b;
    layer0_outputs(2317) <= a and not b;
    layer0_outputs(2318) <= not (a or b);
    layer0_outputs(2319) <= not (a xor b);
    layer0_outputs(2320) <= not b or a;
    layer0_outputs(2321) <= not b or a;
    layer0_outputs(2322) <= b and not a;
    layer0_outputs(2323) <= not (a xor b);
    layer0_outputs(2324) <= a;
    layer0_outputs(2325) <= a xor b;
    layer0_outputs(2326) <= b;
    layer0_outputs(2327) <= not (a or b);
    layer0_outputs(2328) <= not (a or b);
    layer0_outputs(2329) <= not a;
    layer0_outputs(2330) <= not a or b;
    layer0_outputs(2331) <= not (a or b);
    layer0_outputs(2332) <= b and not a;
    layer0_outputs(2333) <= not a or b;
    layer0_outputs(2334) <= not (a xor b);
    layer0_outputs(2335) <= a xor b;
    layer0_outputs(2336) <= not (a or b);
    layer0_outputs(2337) <= not a;
    layer0_outputs(2338) <= a and not b;
    layer0_outputs(2339) <= not (a or b);
    layer0_outputs(2340) <= not a or b;
    layer0_outputs(2341) <= a;
    layer0_outputs(2342) <= '0';
    layer0_outputs(2343) <= a or b;
    layer0_outputs(2344) <= not a;
    layer0_outputs(2345) <= not b;
    layer0_outputs(2346) <= not a or b;
    layer0_outputs(2347) <= a xor b;
    layer0_outputs(2348) <= b and not a;
    layer0_outputs(2349) <= a xor b;
    layer0_outputs(2350) <= b;
    layer0_outputs(2351) <= a or b;
    layer0_outputs(2352) <= not a;
    layer0_outputs(2353) <= '1';
    layer0_outputs(2354) <= not (a xor b);
    layer0_outputs(2355) <= a or b;
    layer0_outputs(2356) <= b;
    layer0_outputs(2357) <= a and not b;
    layer0_outputs(2358) <= not a;
    layer0_outputs(2359) <= a xor b;
    layer0_outputs(2360) <= a;
    layer0_outputs(2361) <= not a or b;
    layer0_outputs(2362) <= not a;
    layer0_outputs(2363) <= a;
    layer0_outputs(2364) <= a;
    layer0_outputs(2365) <= a and not b;
    layer0_outputs(2366) <= not a;
    layer0_outputs(2367) <= b;
    layer0_outputs(2368) <= not (a and b);
    layer0_outputs(2369) <= not b or a;
    layer0_outputs(2370) <= not (a or b);
    layer0_outputs(2371) <= not b;
    layer0_outputs(2372) <= b;
    layer0_outputs(2373) <= a or b;
    layer0_outputs(2374) <= a xor b;
    layer0_outputs(2375) <= '0';
    layer0_outputs(2376) <= a or b;
    layer0_outputs(2377) <= a;
    layer0_outputs(2378) <= a or b;
    layer0_outputs(2379) <= not (a or b);
    layer0_outputs(2380) <= b;
    layer0_outputs(2381) <= b and not a;
    layer0_outputs(2382) <= not a or b;
    layer0_outputs(2383) <= not b;
    layer0_outputs(2384) <= b;
    layer0_outputs(2385) <= a;
    layer0_outputs(2386) <= not a;
    layer0_outputs(2387) <= a or b;
    layer0_outputs(2388) <= a or b;
    layer0_outputs(2389) <= a xor b;
    layer0_outputs(2390) <= not a;
    layer0_outputs(2391) <= not a;
    layer0_outputs(2392) <= b and not a;
    layer0_outputs(2393) <= a or b;
    layer0_outputs(2394) <= a and not b;
    layer0_outputs(2395) <= not (a or b);
    layer0_outputs(2396) <= not a or b;
    layer0_outputs(2397) <= a xor b;
    layer0_outputs(2398) <= a or b;
    layer0_outputs(2399) <= a and b;
    layer0_outputs(2400) <= not (a xor b);
    layer0_outputs(2401) <= b and not a;
    layer0_outputs(2402) <= '0';
    layer0_outputs(2403) <= not (a xor b);
    layer0_outputs(2404) <= not b;
    layer0_outputs(2405) <= not a;
    layer0_outputs(2406) <= not (a or b);
    layer0_outputs(2407) <= a xor b;
    layer0_outputs(2408) <= not (a xor b);
    layer0_outputs(2409) <= b and not a;
    layer0_outputs(2410) <= a xor b;
    layer0_outputs(2411) <= a and b;
    layer0_outputs(2412) <= a or b;
    layer0_outputs(2413) <= not (a or b);
    layer0_outputs(2414) <= a or b;
    layer0_outputs(2415) <= a or b;
    layer0_outputs(2416) <= a;
    layer0_outputs(2417) <= not (a xor b);
    layer0_outputs(2418) <= a or b;
    layer0_outputs(2419) <= not b or a;
    layer0_outputs(2420) <= a xor b;
    layer0_outputs(2421) <= a xor b;
    layer0_outputs(2422) <= not (a or b);
    layer0_outputs(2423) <= not b or a;
    layer0_outputs(2424) <= not a;
    layer0_outputs(2425) <= a or b;
    layer0_outputs(2426) <= not (a or b);
    layer0_outputs(2427) <= b;
    layer0_outputs(2428) <= a and not b;
    layer0_outputs(2429) <= not (a xor b);
    layer0_outputs(2430) <= not (a xor b);
    layer0_outputs(2431) <= a xor b;
    layer0_outputs(2432) <= not b;
    layer0_outputs(2433) <= b;
    layer0_outputs(2434) <= not (a or b);
    layer0_outputs(2435) <= not (a xor b);
    layer0_outputs(2436) <= not (a or b);
    layer0_outputs(2437) <= not b;
    layer0_outputs(2438) <= not (a xor b);
    layer0_outputs(2439) <= not (a or b);
    layer0_outputs(2440) <= not (a or b);
    layer0_outputs(2441) <= b;
    layer0_outputs(2442) <= not a or b;
    layer0_outputs(2443) <= not b;
    layer0_outputs(2444) <= b;
    layer0_outputs(2445) <= '0';
    layer0_outputs(2446) <= b;
    layer0_outputs(2447) <= not (a xor b);
    layer0_outputs(2448) <= b;
    layer0_outputs(2449) <= not b or a;
    layer0_outputs(2450) <= a xor b;
    layer0_outputs(2451) <= not b or a;
    layer0_outputs(2452) <= not a or b;
    layer0_outputs(2453) <= not b or a;
    layer0_outputs(2454) <= a and not b;
    layer0_outputs(2455) <= not (a and b);
    layer0_outputs(2456) <= not (a and b);
    layer0_outputs(2457) <= not (a or b);
    layer0_outputs(2458) <= a or b;
    layer0_outputs(2459) <= a and not b;
    layer0_outputs(2460) <= not (a xor b);
    layer0_outputs(2461) <= not (a or b);
    layer0_outputs(2462) <= not (a or b);
    layer0_outputs(2463) <= not a;
    layer0_outputs(2464) <= '1';
    layer0_outputs(2465) <= a or b;
    layer0_outputs(2466) <= b and not a;
    layer0_outputs(2467) <= a or b;
    layer0_outputs(2468) <= a or b;
    layer0_outputs(2469) <= not a or b;
    layer0_outputs(2470) <= not a;
    layer0_outputs(2471) <= a xor b;
    layer0_outputs(2472) <= not b or a;
    layer0_outputs(2473) <= a or b;
    layer0_outputs(2474) <= not (a or b);
    layer0_outputs(2475) <= not b;
    layer0_outputs(2476) <= a or b;
    layer0_outputs(2477) <= not (a or b);
    layer0_outputs(2478) <= a or b;
    layer0_outputs(2479) <= a or b;
    layer0_outputs(2480) <= a xor b;
    layer0_outputs(2481) <= b and not a;
    layer0_outputs(2482) <= not (a xor b);
    layer0_outputs(2483) <= not a;
    layer0_outputs(2484) <= not (a or b);
    layer0_outputs(2485) <= a or b;
    layer0_outputs(2486) <= not (a or b);
    layer0_outputs(2487) <= not a or b;
    layer0_outputs(2488) <= not a or b;
    layer0_outputs(2489) <= not (a or b);
    layer0_outputs(2490) <= not (a xor b);
    layer0_outputs(2491) <= a or b;
    layer0_outputs(2492) <= '1';
    layer0_outputs(2493) <= not (a or b);
    layer0_outputs(2494) <= not b or a;
    layer0_outputs(2495) <= not a or b;
    layer0_outputs(2496) <= not (a xor b);
    layer0_outputs(2497) <= a and not b;
    layer0_outputs(2498) <= a xor b;
    layer0_outputs(2499) <= not (a or b);
    layer0_outputs(2500) <= not b;
    layer0_outputs(2501) <= not b;
    layer0_outputs(2502) <= b;
    layer0_outputs(2503) <= b;
    layer0_outputs(2504) <= '0';
    layer0_outputs(2505) <= not (a xor b);
    layer0_outputs(2506) <= a or b;
    layer0_outputs(2507) <= not b;
    layer0_outputs(2508) <= not (a or b);
    layer0_outputs(2509) <= not (a xor b);
    layer0_outputs(2510) <= b;
    layer0_outputs(2511) <= not a;
    layer0_outputs(2512) <= a or b;
    layer0_outputs(2513) <= not b or a;
    layer0_outputs(2514) <= a xor b;
    layer0_outputs(2515) <= not b;
    layer0_outputs(2516) <= not (a or b);
    layer0_outputs(2517) <= a or b;
    layer0_outputs(2518) <= not (a or b);
    layer0_outputs(2519) <= a xor b;
    layer0_outputs(2520) <= a or b;
    layer0_outputs(2521) <= not a;
    layer0_outputs(2522) <= not a;
    layer0_outputs(2523) <= a and b;
    layer0_outputs(2524) <= not b;
    layer0_outputs(2525) <= a and not b;
    layer0_outputs(2526) <= not (a or b);
    layer0_outputs(2527) <= not a;
    layer0_outputs(2528) <= not b or a;
    layer0_outputs(2529) <= a;
    layer0_outputs(2530) <= a xor b;
    layer0_outputs(2531) <= a xor b;
    layer0_outputs(2532) <= a xor b;
    layer0_outputs(2533) <= b and not a;
    layer0_outputs(2534) <= not a;
    layer0_outputs(2535) <= not b or a;
    layer0_outputs(2536) <= not (a or b);
    layer0_outputs(2537) <= not b or a;
    layer0_outputs(2538) <= a or b;
    layer0_outputs(2539) <= a xor b;
    layer0_outputs(2540) <= a or b;
    layer0_outputs(2541) <= not b;
    layer0_outputs(2542) <= not (a or b);
    layer0_outputs(2543) <= not a;
    layer0_outputs(2544) <= a and not b;
    layer0_outputs(2545) <= a xor b;
    layer0_outputs(2546) <= a xor b;
    layer0_outputs(2547) <= a xor b;
    layer0_outputs(2548) <= not a;
    layer0_outputs(2549) <= not b;
    layer0_outputs(2550) <= not a;
    layer0_outputs(2551) <= a and not b;
    layer0_outputs(2552) <= b;
    layer0_outputs(2553) <= not b;
    layer0_outputs(2554) <= not (a or b);
    layer0_outputs(2555) <= not (a or b);
    layer0_outputs(2556) <= b and not a;
    layer0_outputs(2557) <= a and not b;
    layer0_outputs(2558) <= not (a or b);
    layer0_outputs(2559) <= b;
    layer0_outputs(2560) <= a and b;
    layer0_outputs(2561) <= not (a or b);
    layer0_outputs(2562) <= not (a or b);
    layer0_outputs(2563) <= not b;
    layer0_outputs(2564) <= not (a xor b);
    layer0_outputs(2565) <= a or b;
    layer0_outputs(2566) <= a xor b;
    layer0_outputs(2567) <= a or b;
    layer0_outputs(2568) <= a or b;
    layer0_outputs(2569) <= a xor b;
    layer0_outputs(2570) <= a xor b;
    layer0_outputs(2571) <= a or b;
    layer0_outputs(2572) <= not a;
    layer0_outputs(2573) <= a or b;
    layer0_outputs(2574) <= b;
    layer0_outputs(2575) <= a and not b;
    layer0_outputs(2576) <= a xor b;
    layer0_outputs(2577) <= a xor b;
    layer0_outputs(2578) <= a;
    layer0_outputs(2579) <= not a or b;
    layer0_outputs(2580) <= not a;
    layer0_outputs(2581) <= b;
    layer0_outputs(2582) <= b and not a;
    layer0_outputs(2583) <= a xor b;
    layer0_outputs(2584) <= a xor b;
    layer0_outputs(2585) <= not b or a;
    layer0_outputs(2586) <= a or b;
    layer0_outputs(2587) <= not a or b;
    layer0_outputs(2588) <= a;
    layer0_outputs(2589) <= a xor b;
    layer0_outputs(2590) <= a or b;
    layer0_outputs(2591) <= not (a xor b);
    layer0_outputs(2592) <= not (a xor b);
    layer0_outputs(2593) <= a;
    layer0_outputs(2594) <= a or b;
    layer0_outputs(2595) <= a and not b;
    layer0_outputs(2596) <= b;
    layer0_outputs(2597) <= a;
    layer0_outputs(2598) <= a;
    layer0_outputs(2599) <= a xor b;
    layer0_outputs(2600) <= a or b;
    layer0_outputs(2601) <= not (a or b);
    layer0_outputs(2602) <= not a or b;
    layer0_outputs(2603) <= not b or a;
    layer0_outputs(2604) <= not b or a;
    layer0_outputs(2605) <= a and not b;
    layer0_outputs(2606) <= not b;
    layer0_outputs(2607) <= a or b;
    layer0_outputs(2608) <= not (a or b);
    layer0_outputs(2609) <= b and not a;
    layer0_outputs(2610) <= not (a or b);
    layer0_outputs(2611) <= not (a or b);
    layer0_outputs(2612) <= a or b;
    layer0_outputs(2613) <= not b;
    layer0_outputs(2614) <= a and not b;
    layer0_outputs(2615) <= a;
    layer0_outputs(2616) <= a xor b;
    layer0_outputs(2617) <= b;
    layer0_outputs(2618) <= a or b;
    layer0_outputs(2619) <= a xor b;
    layer0_outputs(2620) <= a xor b;
    layer0_outputs(2621) <= not (a or b);
    layer0_outputs(2622) <= b and not a;
    layer0_outputs(2623) <= a and not b;
    layer0_outputs(2624) <= a xor b;
    layer0_outputs(2625) <= not (a or b);
    layer0_outputs(2626) <= not b or a;
    layer0_outputs(2627) <= not a;
    layer0_outputs(2628) <= a or b;
    layer0_outputs(2629) <= not (a or b);
    layer0_outputs(2630) <= b and not a;
    layer0_outputs(2631) <= a xor b;
    layer0_outputs(2632) <= not (a xor b);
    layer0_outputs(2633) <= not (a or b);
    layer0_outputs(2634) <= b;
    layer0_outputs(2635) <= not b;
    layer0_outputs(2636) <= a or b;
    layer0_outputs(2637) <= a or b;
    layer0_outputs(2638) <= a or b;
    layer0_outputs(2639) <= a;
    layer0_outputs(2640) <= not a;
    layer0_outputs(2641) <= a;
    layer0_outputs(2642) <= not b;
    layer0_outputs(2643) <= not b;
    layer0_outputs(2644) <= not b;
    layer0_outputs(2645) <= a;
    layer0_outputs(2646) <= not (a or b);
    layer0_outputs(2647) <= not (a and b);
    layer0_outputs(2648) <= not a or b;
    layer0_outputs(2649) <= not a;
    layer0_outputs(2650) <= a xor b;
    layer0_outputs(2651) <= a or b;
    layer0_outputs(2652) <= a and not b;
    layer0_outputs(2653) <= not a;
    layer0_outputs(2654) <= not (a or b);
    layer0_outputs(2655) <= a and not b;
    layer0_outputs(2656) <= not b or a;
    layer0_outputs(2657) <= not b or a;
    layer0_outputs(2658) <= not b or a;
    layer0_outputs(2659) <= a xor b;
    layer0_outputs(2660) <= b;
    layer0_outputs(2661) <= not b;
    layer0_outputs(2662) <= not a;
    layer0_outputs(2663) <= not a or b;
    layer0_outputs(2664) <= not b or a;
    layer0_outputs(2665) <= a and not b;
    layer0_outputs(2666) <= not (a or b);
    layer0_outputs(2667) <= b and not a;
    layer0_outputs(2668) <= not a;
    layer0_outputs(2669) <= b;
    layer0_outputs(2670) <= not a;
    layer0_outputs(2671) <= not a or b;
    layer0_outputs(2672) <= not a or b;
    layer0_outputs(2673) <= not (a or b);
    layer0_outputs(2674) <= a and not b;
    layer0_outputs(2675) <= a or b;
    layer0_outputs(2676) <= b and not a;
    layer0_outputs(2677) <= b;
    layer0_outputs(2678) <= not b or a;
    layer0_outputs(2679) <= a xor b;
    layer0_outputs(2680) <= not (a xor b);
    layer0_outputs(2681) <= b and not a;
    layer0_outputs(2682) <= not (a or b);
    layer0_outputs(2683) <= '1';
    layer0_outputs(2684) <= a and b;
    layer0_outputs(2685) <= not b;
    layer0_outputs(2686) <= not (a or b);
    layer0_outputs(2687) <= a and not b;
    layer0_outputs(2688) <= not b;
    layer0_outputs(2689) <= not (a xor b);
    layer0_outputs(2690) <= not b or a;
    layer0_outputs(2691) <= a xor b;
    layer0_outputs(2692) <= not (a and b);
    layer0_outputs(2693) <= a xor b;
    layer0_outputs(2694) <= a or b;
    layer0_outputs(2695) <= not b;
    layer0_outputs(2696) <= a xor b;
    layer0_outputs(2697) <= not b;
    layer0_outputs(2698) <= a or b;
    layer0_outputs(2699) <= a or b;
    layer0_outputs(2700) <= not (a or b);
    layer0_outputs(2701) <= not (a or b);
    layer0_outputs(2702) <= not a or b;
    layer0_outputs(2703) <= b and not a;
    layer0_outputs(2704) <= not a or b;
    layer0_outputs(2705) <= not a or b;
    layer0_outputs(2706) <= not a;
    layer0_outputs(2707) <= b and not a;
    layer0_outputs(2708) <= a or b;
    layer0_outputs(2709) <= b and not a;
    layer0_outputs(2710) <= b;
    layer0_outputs(2711) <= not (a or b);
    layer0_outputs(2712) <= a or b;
    layer0_outputs(2713) <= not a or b;
    layer0_outputs(2714) <= not (a or b);
    layer0_outputs(2715) <= a xor b;
    layer0_outputs(2716) <= not b;
    layer0_outputs(2717) <= a xor b;
    layer0_outputs(2718) <= not b;
    layer0_outputs(2719) <= not a or b;
    layer0_outputs(2720) <= not (a or b);
    layer0_outputs(2721) <= b;
    layer0_outputs(2722) <= '1';
    layer0_outputs(2723) <= a;
    layer0_outputs(2724) <= not (a or b);
    layer0_outputs(2725) <= b and not a;
    layer0_outputs(2726) <= a xor b;
    layer0_outputs(2727) <= b;
    layer0_outputs(2728) <= a or b;
    layer0_outputs(2729) <= a and not b;
    layer0_outputs(2730) <= not (a xor b);
    layer0_outputs(2731) <= not (a xor b);
    layer0_outputs(2732) <= '1';
    layer0_outputs(2733) <= not a or b;
    layer0_outputs(2734) <= not (a xor b);
    layer0_outputs(2735) <= not b or a;
    layer0_outputs(2736) <= not a;
    layer0_outputs(2737) <= not b or a;
    layer0_outputs(2738) <= not (a xor b);
    layer0_outputs(2739) <= not (a or b);
    layer0_outputs(2740) <= not (a or b);
    layer0_outputs(2741) <= a xor b;
    layer0_outputs(2742) <= not a or b;
    layer0_outputs(2743) <= not (a or b);
    layer0_outputs(2744) <= not a;
    layer0_outputs(2745) <= a xor b;
    layer0_outputs(2746) <= not (a or b);
    layer0_outputs(2747) <= b;
    layer0_outputs(2748) <= a;
    layer0_outputs(2749) <= not (a xor b);
    layer0_outputs(2750) <= not (a xor b);
    layer0_outputs(2751) <= not (a and b);
    layer0_outputs(2752) <= not (a xor b);
    layer0_outputs(2753) <= a and not b;
    layer0_outputs(2754) <= not b or a;
    layer0_outputs(2755) <= not b or a;
    layer0_outputs(2756) <= not b or a;
    layer0_outputs(2757) <= a or b;
    layer0_outputs(2758) <= a or b;
    layer0_outputs(2759) <= a or b;
    layer0_outputs(2760) <= a or b;
    layer0_outputs(2761) <= not (a or b);
    layer0_outputs(2762) <= not (a xor b);
    layer0_outputs(2763) <= not (a or b);
    layer0_outputs(2764) <= not a or b;
    layer0_outputs(2765) <= not (a or b);
    layer0_outputs(2766) <= not b or a;
    layer0_outputs(2767) <= b and not a;
    layer0_outputs(2768) <= a;
    layer0_outputs(2769) <= b and not a;
    layer0_outputs(2770) <= a or b;
    layer0_outputs(2771) <= not (a or b);
    layer0_outputs(2772) <= a xor b;
    layer0_outputs(2773) <= a or b;
    layer0_outputs(2774) <= a and not b;
    layer0_outputs(2775) <= a;
    layer0_outputs(2776) <= a and not b;
    layer0_outputs(2777) <= a and not b;
    layer0_outputs(2778) <= a and not b;
    layer0_outputs(2779) <= b;
    layer0_outputs(2780) <= not b or a;
    layer0_outputs(2781) <= not (a or b);
    layer0_outputs(2782) <= b and not a;
    layer0_outputs(2783) <= a or b;
    layer0_outputs(2784) <= not (a or b);
    layer0_outputs(2785) <= not (a or b);
    layer0_outputs(2786) <= not (a and b);
    layer0_outputs(2787) <= b and not a;
    layer0_outputs(2788) <= not (a or b);
    layer0_outputs(2789) <= not b;
    layer0_outputs(2790) <= b;
    layer0_outputs(2791) <= not a or b;
    layer0_outputs(2792) <= not a;
    layer0_outputs(2793) <= not (a or b);
    layer0_outputs(2794) <= not (a or b);
    layer0_outputs(2795) <= a or b;
    layer0_outputs(2796) <= not b;
    layer0_outputs(2797) <= a and not b;
    layer0_outputs(2798) <= not (a and b);
    layer0_outputs(2799) <= '1';
    layer0_outputs(2800) <= not (a or b);
    layer0_outputs(2801) <= a or b;
    layer0_outputs(2802) <= a xor b;
    layer0_outputs(2803) <= not a;
    layer0_outputs(2804) <= not b or a;
    layer0_outputs(2805) <= a or b;
    layer0_outputs(2806) <= not (a and b);
    layer0_outputs(2807) <= not a or b;
    layer0_outputs(2808) <= b;
    layer0_outputs(2809) <= not b or a;
    layer0_outputs(2810) <= b;
    layer0_outputs(2811) <= a or b;
    layer0_outputs(2812) <= not (a and b);
    layer0_outputs(2813) <= not b;
    layer0_outputs(2814) <= not (a and b);
    layer0_outputs(2815) <= b and not a;
    layer0_outputs(2816) <= not b or a;
    layer0_outputs(2817) <= '0';
    layer0_outputs(2818) <= a and not b;
    layer0_outputs(2819) <= not (a or b);
    layer0_outputs(2820) <= not b;
    layer0_outputs(2821) <= not b or a;
    layer0_outputs(2822) <= '1';
    layer0_outputs(2823) <= not (a xor b);
    layer0_outputs(2824) <= a xor b;
    layer0_outputs(2825) <= b;
    layer0_outputs(2826) <= a or b;
    layer0_outputs(2827) <= not (a or b);
    layer0_outputs(2828) <= not b or a;
    layer0_outputs(2829) <= a xor b;
    layer0_outputs(2830) <= not b;
    layer0_outputs(2831) <= a xor b;
    layer0_outputs(2832) <= a xor b;
    layer0_outputs(2833) <= a and not b;
    layer0_outputs(2834) <= not (a or b);
    layer0_outputs(2835) <= not (a or b);
    layer0_outputs(2836) <= not b;
    layer0_outputs(2837) <= a xor b;
    layer0_outputs(2838) <= not b;
    layer0_outputs(2839) <= b;
    layer0_outputs(2840) <= a;
    layer0_outputs(2841) <= a or b;
    layer0_outputs(2842) <= a or b;
    layer0_outputs(2843) <= not a;
    layer0_outputs(2844) <= not b or a;
    layer0_outputs(2845) <= not (a or b);
    layer0_outputs(2846) <= a or b;
    layer0_outputs(2847) <= not a;
    layer0_outputs(2848) <= not (a xor b);
    layer0_outputs(2849) <= not a or b;
    layer0_outputs(2850) <= b;
    layer0_outputs(2851) <= not (a or b);
    layer0_outputs(2852) <= a and b;
    layer0_outputs(2853) <= not a or b;
    layer0_outputs(2854) <= a xor b;
    layer0_outputs(2855) <= not a or b;
    layer0_outputs(2856) <= '0';
    layer0_outputs(2857) <= a;
    layer0_outputs(2858) <= not (a xor b);
    layer0_outputs(2859) <= not (a or b);
    layer0_outputs(2860) <= a xor b;
    layer0_outputs(2861) <= not (a xor b);
    layer0_outputs(2862) <= not (a or b);
    layer0_outputs(2863) <= not (a xor b);
    layer0_outputs(2864) <= not (a xor b);
    layer0_outputs(2865) <= a or b;
    layer0_outputs(2866) <= not (a xor b);
    layer0_outputs(2867) <= a and not b;
    layer0_outputs(2868) <= not (a xor b);
    layer0_outputs(2869) <= not b;
    layer0_outputs(2870) <= a xor b;
    layer0_outputs(2871) <= not b;
    layer0_outputs(2872) <= a and not b;
    layer0_outputs(2873) <= a or b;
    layer0_outputs(2874) <= a;
    layer0_outputs(2875) <= a xor b;
    layer0_outputs(2876) <= b;
    layer0_outputs(2877) <= b and not a;
    layer0_outputs(2878) <= a;
    layer0_outputs(2879) <= a or b;
    layer0_outputs(2880) <= not (a xor b);
    layer0_outputs(2881) <= a and b;
    layer0_outputs(2882) <= a and not b;
    layer0_outputs(2883) <= a or b;
    layer0_outputs(2884) <= b;
    layer0_outputs(2885) <= a and not b;
    layer0_outputs(2886) <= not b;
    layer0_outputs(2887) <= b and not a;
    layer0_outputs(2888) <= not b;
    layer0_outputs(2889) <= b;
    layer0_outputs(2890) <= not (a and b);
    layer0_outputs(2891) <= a or b;
    layer0_outputs(2892) <= not a;
    layer0_outputs(2893) <= a and b;
    layer0_outputs(2894) <= b;
    layer0_outputs(2895) <= a xor b;
    layer0_outputs(2896) <= a and not b;
    layer0_outputs(2897) <= b;
    layer0_outputs(2898) <= not (a or b);
    layer0_outputs(2899) <= not a or b;
    layer0_outputs(2900) <= a and not b;
    layer0_outputs(2901) <= a or b;
    layer0_outputs(2902) <= not (a or b);
    layer0_outputs(2903) <= not (a xor b);
    layer0_outputs(2904) <= a and not b;
    layer0_outputs(2905) <= not (a or b);
    layer0_outputs(2906) <= not (a xor b);
    layer0_outputs(2907) <= b;
    layer0_outputs(2908) <= b;
    layer0_outputs(2909) <= a;
    layer0_outputs(2910) <= not b;
    layer0_outputs(2911) <= not (a xor b);
    layer0_outputs(2912) <= a and not b;
    layer0_outputs(2913) <= not a;
    layer0_outputs(2914) <= a or b;
    layer0_outputs(2915) <= not b;
    layer0_outputs(2916) <= '0';
    layer0_outputs(2917) <= not a or b;
    layer0_outputs(2918) <= not a or b;
    layer0_outputs(2919) <= not (a xor b);
    layer0_outputs(2920) <= not a;
    layer0_outputs(2921) <= a and not b;
    layer0_outputs(2922) <= a xor b;
    layer0_outputs(2923) <= not (a xor b);
    layer0_outputs(2924) <= b and not a;
    layer0_outputs(2925) <= a xor b;
    layer0_outputs(2926) <= not a or b;
    layer0_outputs(2927) <= b;
    layer0_outputs(2928) <= a and not b;
    layer0_outputs(2929) <= not (a or b);
    layer0_outputs(2930) <= a or b;
    layer0_outputs(2931) <= a or b;
    layer0_outputs(2932) <= not (a or b);
    layer0_outputs(2933) <= not (a xor b);
    layer0_outputs(2934) <= not a;
    layer0_outputs(2935) <= b and not a;
    layer0_outputs(2936) <= b and not a;
    layer0_outputs(2937) <= a xor b;
    layer0_outputs(2938) <= b;
    layer0_outputs(2939) <= a xor b;
    layer0_outputs(2940) <= b;
    layer0_outputs(2941) <= not (a or b);
    layer0_outputs(2942) <= not a or b;
    layer0_outputs(2943) <= not b;
    layer0_outputs(2944) <= not a;
    layer0_outputs(2945) <= a or b;
    layer0_outputs(2946) <= a and not b;
    layer0_outputs(2947) <= not (a xor b);
    layer0_outputs(2948) <= a or b;
    layer0_outputs(2949) <= b and not a;
    layer0_outputs(2950) <= a xor b;
    layer0_outputs(2951) <= b;
    layer0_outputs(2952) <= b and not a;
    layer0_outputs(2953) <= a;
    layer0_outputs(2954) <= not b or a;
    layer0_outputs(2955) <= not (a xor b);
    layer0_outputs(2956) <= a;
    layer0_outputs(2957) <= a and not b;
    layer0_outputs(2958) <= a xor b;
    layer0_outputs(2959) <= a and b;
    layer0_outputs(2960) <= not (a xor b);
    layer0_outputs(2961) <= a;
    layer0_outputs(2962) <= not (a or b);
    layer0_outputs(2963) <= not (a xor b);
    layer0_outputs(2964) <= not (a or b);
    layer0_outputs(2965) <= not a or b;
    layer0_outputs(2966) <= a and not b;
    layer0_outputs(2967) <= a or b;
    layer0_outputs(2968) <= a xor b;
    layer0_outputs(2969) <= not a;
    layer0_outputs(2970) <= a xor b;
    layer0_outputs(2971) <= not a;
    layer0_outputs(2972) <= not a;
    layer0_outputs(2973) <= b and not a;
    layer0_outputs(2974) <= not (a xor b);
    layer0_outputs(2975) <= a and not b;
    layer0_outputs(2976) <= a or b;
    layer0_outputs(2977) <= not b;
    layer0_outputs(2978) <= a xor b;
    layer0_outputs(2979) <= '0';
    layer0_outputs(2980) <= not (a or b);
    layer0_outputs(2981) <= b;
    layer0_outputs(2982) <= '1';
    layer0_outputs(2983) <= not (a or b);
    layer0_outputs(2984) <= b and not a;
    layer0_outputs(2985) <= a or b;
    layer0_outputs(2986) <= a or b;
    layer0_outputs(2987) <= b;
    layer0_outputs(2988) <= not a or b;
    layer0_outputs(2989) <= '0';
    layer0_outputs(2990) <= a or b;
    layer0_outputs(2991) <= a;
    layer0_outputs(2992) <= a or b;
    layer0_outputs(2993) <= not (a or b);
    layer0_outputs(2994) <= not b;
    layer0_outputs(2995) <= a;
    layer0_outputs(2996) <= not a or b;
    layer0_outputs(2997) <= not (a or b);
    layer0_outputs(2998) <= b;
    layer0_outputs(2999) <= '0';
    layer0_outputs(3000) <= '1';
    layer0_outputs(3001) <= not b;
    layer0_outputs(3002) <= not (a xor b);
    layer0_outputs(3003) <= '0';
    layer0_outputs(3004) <= a or b;
    layer0_outputs(3005) <= '0';
    layer0_outputs(3006) <= not a;
    layer0_outputs(3007) <= not b;
    layer0_outputs(3008) <= not (a or b);
    layer0_outputs(3009) <= a;
    layer0_outputs(3010) <= not (a or b);
    layer0_outputs(3011) <= not (a or b);
    layer0_outputs(3012) <= b;
    layer0_outputs(3013) <= a or b;
    layer0_outputs(3014) <= a or b;
    layer0_outputs(3015) <= not (a or b);
    layer0_outputs(3016) <= not (a xor b);
    layer0_outputs(3017) <= a and not b;
    layer0_outputs(3018) <= '0';
    layer0_outputs(3019) <= a and not b;
    layer0_outputs(3020) <= not (a xor b);
    layer0_outputs(3021) <= not (a xor b);
    layer0_outputs(3022) <= not a or b;
    layer0_outputs(3023) <= not (a xor b);
    layer0_outputs(3024) <= a;
    layer0_outputs(3025) <= not b;
    layer0_outputs(3026) <= not (a xor b);
    layer0_outputs(3027) <= not (a xor b);
    layer0_outputs(3028) <= not b;
    layer0_outputs(3029) <= not (a or b);
    layer0_outputs(3030) <= b;
    layer0_outputs(3031) <= not a or b;
    layer0_outputs(3032) <= '0';
    layer0_outputs(3033) <= not (a xor b);
    layer0_outputs(3034) <= not a;
    layer0_outputs(3035) <= not b or a;
    layer0_outputs(3036) <= a and not b;
    layer0_outputs(3037) <= not a;
    layer0_outputs(3038) <= not b;
    layer0_outputs(3039) <= not (a or b);
    layer0_outputs(3040) <= not b or a;
    layer0_outputs(3041) <= not (a xor b);
    layer0_outputs(3042) <= not a or b;
    layer0_outputs(3043) <= a or b;
    layer0_outputs(3044) <= b and not a;
    layer0_outputs(3045) <= not (a xor b);
    layer0_outputs(3046) <= not a or b;
    layer0_outputs(3047) <= a or b;
    layer0_outputs(3048) <= b;
    layer0_outputs(3049) <= not b or a;
    layer0_outputs(3050) <= a or b;
    layer0_outputs(3051) <= b and not a;
    layer0_outputs(3052) <= b and not a;
    layer0_outputs(3053) <= a and b;
    layer0_outputs(3054) <= not (a xor b);
    layer0_outputs(3055) <= b and not a;
    layer0_outputs(3056) <= not b or a;
    layer0_outputs(3057) <= a xor b;
    layer0_outputs(3058) <= not (a or b);
    layer0_outputs(3059) <= a xor b;
    layer0_outputs(3060) <= not (a xor b);
    layer0_outputs(3061) <= not a;
    layer0_outputs(3062) <= not (a xor b);
    layer0_outputs(3063) <= not b or a;
    layer0_outputs(3064) <= a and not b;
    layer0_outputs(3065) <= not (a or b);
    layer0_outputs(3066) <= not (a xor b);
    layer0_outputs(3067) <= a xor b;
    layer0_outputs(3068) <= a or b;
    layer0_outputs(3069) <= a;
    layer0_outputs(3070) <= a;
    layer0_outputs(3071) <= a xor b;
    layer0_outputs(3072) <= a;
    layer0_outputs(3073) <= not (a or b);
    layer0_outputs(3074) <= not (a or b);
    layer0_outputs(3075) <= a xor b;
    layer0_outputs(3076) <= not (a xor b);
    layer0_outputs(3077) <= not a or b;
    layer0_outputs(3078) <= not (a or b);
    layer0_outputs(3079) <= a xor b;
    layer0_outputs(3080) <= a or b;
    layer0_outputs(3081) <= not b or a;
    layer0_outputs(3082) <= a and not b;
    layer0_outputs(3083) <= not (a xor b);
    layer0_outputs(3084) <= not b or a;
    layer0_outputs(3085) <= b and not a;
    layer0_outputs(3086) <= not b;
    layer0_outputs(3087) <= a;
    layer0_outputs(3088) <= b;
    layer0_outputs(3089) <= a;
    layer0_outputs(3090) <= b and not a;
    layer0_outputs(3091) <= not (a or b);
    layer0_outputs(3092) <= not b;
    layer0_outputs(3093) <= not a;
    layer0_outputs(3094) <= a xor b;
    layer0_outputs(3095) <= b and not a;
    layer0_outputs(3096) <= not b;
    layer0_outputs(3097) <= not (a xor b);
    layer0_outputs(3098) <= b and not a;
    layer0_outputs(3099) <= a and b;
    layer0_outputs(3100) <= not b or a;
    layer0_outputs(3101) <= b and not a;
    layer0_outputs(3102) <= a or b;
    layer0_outputs(3103) <= b and not a;
    layer0_outputs(3104) <= not (a xor b);
    layer0_outputs(3105) <= not (a xor b);
    layer0_outputs(3106) <= not b;
    layer0_outputs(3107) <= '1';
    layer0_outputs(3108) <= not b;
    layer0_outputs(3109) <= a and b;
    layer0_outputs(3110) <= b and not a;
    layer0_outputs(3111) <= a xor b;
    layer0_outputs(3112) <= not a or b;
    layer0_outputs(3113) <= not b;
    layer0_outputs(3114) <= not a;
    layer0_outputs(3115) <= not a;
    layer0_outputs(3116) <= b and not a;
    layer0_outputs(3117) <= not (a or b);
    layer0_outputs(3118) <= not (a or b);
    layer0_outputs(3119) <= a and not b;
    layer0_outputs(3120) <= not b;
    layer0_outputs(3121) <= a or b;
    layer0_outputs(3122) <= not b or a;
    layer0_outputs(3123) <= b and not a;
    layer0_outputs(3124) <= not (a or b);
    layer0_outputs(3125) <= not (a or b);
    layer0_outputs(3126) <= not (a xor b);
    layer0_outputs(3127) <= not (a or b);
    layer0_outputs(3128) <= a or b;
    layer0_outputs(3129) <= a or b;
    layer0_outputs(3130) <= not b or a;
    layer0_outputs(3131) <= not a;
    layer0_outputs(3132) <= b and not a;
    layer0_outputs(3133) <= not a or b;
    layer0_outputs(3134) <= not (a and b);
    layer0_outputs(3135) <= not (a or b);
    layer0_outputs(3136) <= a or b;
    layer0_outputs(3137) <= not a or b;
    layer0_outputs(3138) <= b;
    layer0_outputs(3139) <= b;
    layer0_outputs(3140) <= '1';
    layer0_outputs(3141) <= a;
    layer0_outputs(3142) <= b;
    layer0_outputs(3143) <= not b or a;
    layer0_outputs(3144) <= not a;
    layer0_outputs(3145) <= not b;
    layer0_outputs(3146) <= a and not b;
    layer0_outputs(3147) <= a or b;
    layer0_outputs(3148) <= not (a xor b);
    layer0_outputs(3149) <= not a;
    layer0_outputs(3150) <= not (a xor b);
    layer0_outputs(3151) <= not a or b;
    layer0_outputs(3152) <= not a or b;
    layer0_outputs(3153) <= not a or b;
    layer0_outputs(3154) <= not a;
    layer0_outputs(3155) <= b and not a;
    layer0_outputs(3156) <= b;
    layer0_outputs(3157) <= not (a or b);
    layer0_outputs(3158) <= not b;
    layer0_outputs(3159) <= not a or b;
    layer0_outputs(3160) <= a or b;
    layer0_outputs(3161) <= b and not a;
    layer0_outputs(3162) <= not b;
    layer0_outputs(3163) <= not (a xor b);
    layer0_outputs(3164) <= a xor b;
    layer0_outputs(3165) <= not (a and b);
    layer0_outputs(3166) <= not b;
    layer0_outputs(3167) <= not (a or b);
    layer0_outputs(3168) <= a;
    layer0_outputs(3169) <= a or b;
    layer0_outputs(3170) <= '0';
    layer0_outputs(3171) <= not (a xor b);
    layer0_outputs(3172) <= not a or b;
    layer0_outputs(3173) <= not b;
    layer0_outputs(3174) <= a and b;
    layer0_outputs(3175) <= a and not b;
    layer0_outputs(3176) <= not b or a;
    layer0_outputs(3177) <= a or b;
    layer0_outputs(3178) <= not b;
    layer0_outputs(3179) <= not a;
    layer0_outputs(3180) <= a xor b;
    layer0_outputs(3181) <= b;
    layer0_outputs(3182) <= a or b;
    layer0_outputs(3183) <= b and not a;
    layer0_outputs(3184) <= not a or b;
    layer0_outputs(3185) <= not (a xor b);
    layer0_outputs(3186) <= a;
    layer0_outputs(3187) <= not b;
    layer0_outputs(3188) <= not a;
    layer0_outputs(3189) <= b;
    layer0_outputs(3190) <= not a or b;
    layer0_outputs(3191) <= not a;
    layer0_outputs(3192) <= a xor b;
    layer0_outputs(3193) <= not a or b;
    layer0_outputs(3194) <= not a;
    layer0_outputs(3195) <= not a or b;
    layer0_outputs(3196) <= not (a xor b);
    layer0_outputs(3197) <= not b or a;
    layer0_outputs(3198) <= a xor b;
    layer0_outputs(3199) <= b;
    layer0_outputs(3200) <= not a;
    layer0_outputs(3201) <= not a;
    layer0_outputs(3202) <= not a;
    layer0_outputs(3203) <= a and not b;
    layer0_outputs(3204) <= not b;
    layer0_outputs(3205) <= a xor b;
    layer0_outputs(3206) <= a and not b;
    layer0_outputs(3207) <= not b;
    layer0_outputs(3208) <= not b or a;
    layer0_outputs(3209) <= not a;
    layer0_outputs(3210) <= a or b;
    layer0_outputs(3211) <= not a or b;
    layer0_outputs(3212) <= '1';
    layer0_outputs(3213) <= a xor b;
    layer0_outputs(3214) <= not (a xor b);
    layer0_outputs(3215) <= a or b;
    layer0_outputs(3216) <= not a or b;
    layer0_outputs(3217) <= not a or b;
    layer0_outputs(3218) <= a and not b;
    layer0_outputs(3219) <= a xor b;
    layer0_outputs(3220) <= a or b;
    layer0_outputs(3221) <= not a;
    layer0_outputs(3222) <= a xor b;
    layer0_outputs(3223) <= a or b;
    layer0_outputs(3224) <= not (a xor b);
    layer0_outputs(3225) <= b;
    layer0_outputs(3226) <= a xor b;
    layer0_outputs(3227) <= not a or b;
    layer0_outputs(3228) <= a and not b;
    layer0_outputs(3229) <= not b or a;
    layer0_outputs(3230) <= not a;
    layer0_outputs(3231) <= not b;
    layer0_outputs(3232) <= a or b;
    layer0_outputs(3233) <= a or b;
    layer0_outputs(3234) <= not (a or b);
    layer0_outputs(3235) <= a xor b;
    layer0_outputs(3236) <= not (a or b);
    layer0_outputs(3237) <= a and not b;
    layer0_outputs(3238) <= not a or b;
    layer0_outputs(3239) <= b;
    layer0_outputs(3240) <= a and not b;
    layer0_outputs(3241) <= not (a xor b);
    layer0_outputs(3242) <= b and not a;
    layer0_outputs(3243) <= not b;
    layer0_outputs(3244) <= a or b;
    layer0_outputs(3245) <= not b;
    layer0_outputs(3246) <= a or b;
    layer0_outputs(3247) <= not a or b;
    layer0_outputs(3248) <= not (a xor b);
    layer0_outputs(3249) <= not (a xor b);
    layer0_outputs(3250) <= not a or b;
    layer0_outputs(3251) <= a;
    layer0_outputs(3252) <= a or b;
    layer0_outputs(3253) <= not a or b;
    layer0_outputs(3254) <= not (a xor b);
    layer0_outputs(3255) <= not (a xor b);
    layer0_outputs(3256) <= a and not b;
    layer0_outputs(3257) <= not (a xor b);
    layer0_outputs(3258) <= a or b;
    layer0_outputs(3259) <= b and not a;
    layer0_outputs(3260) <= not b or a;
    layer0_outputs(3261) <= a xor b;
    layer0_outputs(3262) <= not b or a;
    layer0_outputs(3263) <= a or b;
    layer0_outputs(3264) <= not a or b;
    layer0_outputs(3265) <= not b;
    layer0_outputs(3266) <= b;
    layer0_outputs(3267) <= b;
    layer0_outputs(3268) <= b and not a;
    layer0_outputs(3269) <= not (a xor b);
    layer0_outputs(3270) <= b and not a;
    layer0_outputs(3271) <= not (a and b);
    layer0_outputs(3272) <= a and b;
    layer0_outputs(3273) <= not a or b;
    layer0_outputs(3274) <= '1';
    layer0_outputs(3275) <= a or b;
    layer0_outputs(3276) <= a or b;
    layer0_outputs(3277) <= not a;
    layer0_outputs(3278) <= a and b;
    layer0_outputs(3279) <= a or b;
    layer0_outputs(3280) <= not b;
    layer0_outputs(3281) <= not (a xor b);
    layer0_outputs(3282) <= a;
    layer0_outputs(3283) <= not (a or b);
    layer0_outputs(3284) <= b;
    layer0_outputs(3285) <= not (a xor b);
    layer0_outputs(3286) <= not b or a;
    layer0_outputs(3287) <= a xor b;
    layer0_outputs(3288) <= not a;
    layer0_outputs(3289) <= not a or b;
    layer0_outputs(3290) <= not (a xor b);
    layer0_outputs(3291) <= not (a or b);
    layer0_outputs(3292) <= a and not b;
    layer0_outputs(3293) <= b;
    layer0_outputs(3294) <= not b or a;
    layer0_outputs(3295) <= not b or a;
    layer0_outputs(3296) <= b and not a;
    layer0_outputs(3297) <= not (a or b);
    layer0_outputs(3298) <= a or b;
    layer0_outputs(3299) <= not (a xor b);
    layer0_outputs(3300) <= a or b;
    layer0_outputs(3301) <= a xor b;
    layer0_outputs(3302) <= not b;
    layer0_outputs(3303) <= not b or a;
    layer0_outputs(3304) <= not b or a;
    layer0_outputs(3305) <= a;
    layer0_outputs(3306) <= not (a or b);
    layer0_outputs(3307) <= a xor b;
    layer0_outputs(3308) <= b and not a;
    layer0_outputs(3309) <= not (a xor b);
    layer0_outputs(3310) <= not (a and b);
    layer0_outputs(3311) <= a or b;
    layer0_outputs(3312) <= not (a xor b);
    layer0_outputs(3313) <= not a or b;
    layer0_outputs(3314) <= not (a and b);
    layer0_outputs(3315) <= not (a xor b);
    layer0_outputs(3316) <= not (a xor b);
    layer0_outputs(3317) <= a or b;
    layer0_outputs(3318) <= not (a or b);
    layer0_outputs(3319) <= not (a xor b);
    layer0_outputs(3320) <= '0';
    layer0_outputs(3321) <= a;
    layer0_outputs(3322) <= a and not b;
    layer0_outputs(3323) <= b and not a;
    layer0_outputs(3324) <= a or b;
    layer0_outputs(3325) <= not (a xor b);
    layer0_outputs(3326) <= not a;
    layer0_outputs(3327) <= not a;
    layer0_outputs(3328) <= not (a xor b);
    layer0_outputs(3329) <= a;
    layer0_outputs(3330) <= a xor b;
    layer0_outputs(3331) <= a xor b;
    layer0_outputs(3332) <= a;
    layer0_outputs(3333) <= not b or a;
    layer0_outputs(3334) <= a and not b;
    layer0_outputs(3335) <= a xor b;
    layer0_outputs(3336) <= not (a xor b);
    layer0_outputs(3337) <= a xor b;
    layer0_outputs(3338) <= not b or a;
    layer0_outputs(3339) <= b and not a;
    layer0_outputs(3340) <= a or b;
    layer0_outputs(3341) <= not (a xor b);
    layer0_outputs(3342) <= not (a or b);
    layer0_outputs(3343) <= a or b;
    layer0_outputs(3344) <= a and not b;
    layer0_outputs(3345) <= not b;
    layer0_outputs(3346) <= b;
    layer0_outputs(3347) <= b;
    layer0_outputs(3348) <= not b;
    layer0_outputs(3349) <= a and b;
    layer0_outputs(3350) <= a or b;
    layer0_outputs(3351) <= not b;
    layer0_outputs(3352) <= a;
    layer0_outputs(3353) <= not b;
    layer0_outputs(3354) <= not b;
    layer0_outputs(3355) <= a;
    layer0_outputs(3356) <= a and not b;
    layer0_outputs(3357) <= a or b;
    layer0_outputs(3358) <= not b or a;
    layer0_outputs(3359) <= not a;
    layer0_outputs(3360) <= not a;
    layer0_outputs(3361) <= not a or b;
    layer0_outputs(3362) <= not a or b;
    layer0_outputs(3363) <= not b or a;
    layer0_outputs(3364) <= not b or a;
    layer0_outputs(3365) <= not a or b;
    layer0_outputs(3366) <= not (a or b);
    layer0_outputs(3367) <= not b or a;
    layer0_outputs(3368) <= a;
    layer0_outputs(3369) <= b;
    layer0_outputs(3370) <= not b or a;
    layer0_outputs(3371) <= not (a and b);
    layer0_outputs(3372) <= a or b;
    layer0_outputs(3373) <= not b or a;
    layer0_outputs(3374) <= not (a or b);
    layer0_outputs(3375) <= not a;
    layer0_outputs(3376) <= not (a xor b);
    layer0_outputs(3377) <= b;
    layer0_outputs(3378) <= not a or b;
    layer0_outputs(3379) <= not (a or b);
    layer0_outputs(3380) <= a or b;
    layer0_outputs(3381) <= a and not b;
    layer0_outputs(3382) <= a xor b;
    layer0_outputs(3383) <= a or b;
    layer0_outputs(3384) <= not a;
    layer0_outputs(3385) <= b and not a;
    layer0_outputs(3386) <= not b or a;
    layer0_outputs(3387) <= not b or a;
    layer0_outputs(3388) <= not (a or b);
    layer0_outputs(3389) <= not a;
    layer0_outputs(3390) <= not a;
    layer0_outputs(3391) <= a or b;
    layer0_outputs(3392) <= '1';
    layer0_outputs(3393) <= not (a or b);
    layer0_outputs(3394) <= a xor b;
    layer0_outputs(3395) <= not (a or b);
    layer0_outputs(3396) <= not (a xor b);
    layer0_outputs(3397) <= not (a and b);
    layer0_outputs(3398) <= not a;
    layer0_outputs(3399) <= b and not a;
    layer0_outputs(3400) <= not (a or b);
    layer0_outputs(3401) <= not (a xor b);
    layer0_outputs(3402) <= not a or b;
    layer0_outputs(3403) <= a xor b;
    layer0_outputs(3404) <= b and not a;
    layer0_outputs(3405) <= not (a or b);
    layer0_outputs(3406) <= not (a xor b);
    layer0_outputs(3407) <= a;
    layer0_outputs(3408) <= not b or a;
    layer0_outputs(3409) <= not b or a;
    layer0_outputs(3410) <= a or b;
    layer0_outputs(3411) <= a and not b;
    layer0_outputs(3412) <= not (a or b);
    layer0_outputs(3413) <= not (a xor b);
    layer0_outputs(3414) <= not a or b;
    layer0_outputs(3415) <= not a or b;
    layer0_outputs(3416) <= a xor b;
    layer0_outputs(3417) <= not (a or b);
    layer0_outputs(3418) <= '0';
    layer0_outputs(3419) <= not (a xor b);
    layer0_outputs(3420) <= not a or b;
    layer0_outputs(3421) <= not a;
    layer0_outputs(3422) <= a;
    layer0_outputs(3423) <= b and not a;
    layer0_outputs(3424) <= not b;
    layer0_outputs(3425) <= not (a and b);
    layer0_outputs(3426) <= not b;
    layer0_outputs(3427) <= a and not b;
    layer0_outputs(3428) <= b and not a;
    layer0_outputs(3429) <= not b;
    layer0_outputs(3430) <= not (a or b);
    layer0_outputs(3431) <= a;
    layer0_outputs(3432) <= not b;
    layer0_outputs(3433) <= not (a or b);
    layer0_outputs(3434) <= not a or b;
    layer0_outputs(3435) <= not a;
    layer0_outputs(3436) <= not a or b;
    layer0_outputs(3437) <= not (a or b);
    layer0_outputs(3438) <= not b or a;
    layer0_outputs(3439) <= a or b;
    layer0_outputs(3440) <= not (a or b);
    layer0_outputs(3441) <= b and not a;
    layer0_outputs(3442) <= not a or b;
    layer0_outputs(3443) <= not (a xor b);
    layer0_outputs(3444) <= a;
    layer0_outputs(3445) <= a or b;
    layer0_outputs(3446) <= not (a or b);
    layer0_outputs(3447) <= '0';
    layer0_outputs(3448) <= not b;
    layer0_outputs(3449) <= not (a or b);
    layer0_outputs(3450) <= not a;
    layer0_outputs(3451) <= not b or a;
    layer0_outputs(3452) <= a xor b;
    layer0_outputs(3453) <= not b or a;
    layer0_outputs(3454) <= not a;
    layer0_outputs(3455) <= not (a or b);
    layer0_outputs(3456) <= a;
    layer0_outputs(3457) <= not b;
    layer0_outputs(3458) <= a or b;
    layer0_outputs(3459) <= not b;
    layer0_outputs(3460) <= not b or a;
    layer0_outputs(3461) <= '0';
    layer0_outputs(3462) <= a xor b;
    layer0_outputs(3463) <= b and not a;
    layer0_outputs(3464) <= a and not b;
    layer0_outputs(3465) <= not (a or b);
    layer0_outputs(3466) <= not b or a;
    layer0_outputs(3467) <= a or b;
    layer0_outputs(3468) <= a;
    layer0_outputs(3469) <= b and not a;
    layer0_outputs(3470) <= b and not a;
    layer0_outputs(3471) <= a xor b;
    layer0_outputs(3472) <= a and not b;
    layer0_outputs(3473) <= not (a or b);
    layer0_outputs(3474) <= a and not b;
    layer0_outputs(3475) <= a or b;
    layer0_outputs(3476) <= not a or b;
    layer0_outputs(3477) <= not a;
    layer0_outputs(3478) <= a and not b;
    layer0_outputs(3479) <= b;
    layer0_outputs(3480) <= not b or a;
    layer0_outputs(3481) <= not (a xor b);
    layer0_outputs(3482) <= not (a or b);
    layer0_outputs(3483) <= not a;
    layer0_outputs(3484) <= a xor b;
    layer0_outputs(3485) <= not (a or b);
    layer0_outputs(3486) <= not b or a;
    layer0_outputs(3487) <= not b;
    layer0_outputs(3488) <= a or b;
    layer0_outputs(3489) <= not (a xor b);
    layer0_outputs(3490) <= '0';
    layer0_outputs(3491) <= a;
    layer0_outputs(3492) <= not a or b;
    layer0_outputs(3493) <= not a or b;
    layer0_outputs(3494) <= a or b;
    layer0_outputs(3495) <= not a or b;
    layer0_outputs(3496) <= not (a or b);
    layer0_outputs(3497) <= a and b;
    layer0_outputs(3498) <= not (a or b);
    layer0_outputs(3499) <= a;
    layer0_outputs(3500) <= not (a xor b);
    layer0_outputs(3501) <= a xor b;
    layer0_outputs(3502) <= not (a or b);
    layer0_outputs(3503) <= not (a xor b);
    layer0_outputs(3504) <= not (a xor b);
    layer0_outputs(3505) <= not (a or b);
    layer0_outputs(3506) <= not (a and b);
    layer0_outputs(3507) <= b and not a;
    layer0_outputs(3508) <= not (a and b);
    layer0_outputs(3509) <= a or b;
    layer0_outputs(3510) <= not (a or b);
    layer0_outputs(3511) <= not (a or b);
    layer0_outputs(3512) <= not b or a;
    layer0_outputs(3513) <= not b;
    layer0_outputs(3514) <= not (a xor b);
    layer0_outputs(3515) <= not (a xor b);
    layer0_outputs(3516) <= not b;
    layer0_outputs(3517) <= '0';
    layer0_outputs(3518) <= not a or b;
    layer0_outputs(3519) <= not a or b;
    layer0_outputs(3520) <= not b or a;
    layer0_outputs(3521) <= not a;
    layer0_outputs(3522) <= a and not b;
    layer0_outputs(3523) <= '1';
    layer0_outputs(3524) <= b and not a;
    layer0_outputs(3525) <= not a;
    layer0_outputs(3526) <= a and b;
    layer0_outputs(3527) <= a and b;
    layer0_outputs(3528) <= not b or a;
    layer0_outputs(3529) <= a xor b;
    layer0_outputs(3530) <= not (a xor b);
    layer0_outputs(3531) <= not (a or b);
    layer0_outputs(3532) <= b and not a;
    layer0_outputs(3533) <= a;
    layer0_outputs(3534) <= a or b;
    layer0_outputs(3535) <= not a;
    layer0_outputs(3536) <= not b or a;
    layer0_outputs(3537) <= a and not b;
    layer0_outputs(3538) <= not b;
    layer0_outputs(3539) <= not (a or b);
    layer0_outputs(3540) <= a or b;
    layer0_outputs(3541) <= not a;
    layer0_outputs(3542) <= a xor b;
    layer0_outputs(3543) <= a or b;
    layer0_outputs(3544) <= '1';
    layer0_outputs(3545) <= a or b;
    layer0_outputs(3546) <= a xor b;
    layer0_outputs(3547) <= a and not b;
    layer0_outputs(3548) <= '1';
    layer0_outputs(3549) <= not b or a;
    layer0_outputs(3550) <= b;
    layer0_outputs(3551) <= not (a xor b);
    layer0_outputs(3552) <= b and not a;
    layer0_outputs(3553) <= a xor b;
    layer0_outputs(3554) <= not a;
    layer0_outputs(3555) <= a xor b;
    layer0_outputs(3556) <= not a;
    layer0_outputs(3557) <= b and not a;
    layer0_outputs(3558) <= not b;
    layer0_outputs(3559) <= not a or b;
    layer0_outputs(3560) <= a;
    layer0_outputs(3561) <= not b;
    layer0_outputs(3562) <= a or b;
    layer0_outputs(3563) <= a xor b;
    layer0_outputs(3564) <= a;
    layer0_outputs(3565) <= b;
    layer0_outputs(3566) <= not a or b;
    layer0_outputs(3567) <= a and b;
    layer0_outputs(3568) <= not (a or b);
    layer0_outputs(3569) <= not (a or b);
    layer0_outputs(3570) <= b;
    layer0_outputs(3571) <= not (a xor b);
    layer0_outputs(3572) <= not a or b;
    layer0_outputs(3573) <= not (a or b);
    layer0_outputs(3574) <= a or b;
    layer0_outputs(3575) <= not b;
    layer0_outputs(3576) <= not a;
    layer0_outputs(3577) <= a and not b;
    layer0_outputs(3578) <= not (a or b);
    layer0_outputs(3579) <= not (a or b);
    layer0_outputs(3580) <= not b;
    layer0_outputs(3581) <= b;
    layer0_outputs(3582) <= not (a or b);
    layer0_outputs(3583) <= not (a or b);
    layer0_outputs(3584) <= a;
    layer0_outputs(3585) <= a and not b;
    layer0_outputs(3586) <= a or b;
    layer0_outputs(3587) <= not b;
    layer0_outputs(3588) <= a xor b;
    layer0_outputs(3589) <= not a;
    layer0_outputs(3590) <= not b;
    layer0_outputs(3591) <= not (a or b);
    layer0_outputs(3592) <= a and not b;
    layer0_outputs(3593) <= not b or a;
    layer0_outputs(3594) <= a or b;
    layer0_outputs(3595) <= not b or a;
    layer0_outputs(3596) <= a or b;
    layer0_outputs(3597) <= a or b;
    layer0_outputs(3598) <= not (a or b);
    layer0_outputs(3599) <= not b or a;
    layer0_outputs(3600) <= a xor b;
    layer0_outputs(3601) <= not (a xor b);
    layer0_outputs(3602) <= not a;
    layer0_outputs(3603) <= not b or a;
    layer0_outputs(3604) <= b;
    layer0_outputs(3605) <= b;
    layer0_outputs(3606) <= not (a and b);
    layer0_outputs(3607) <= not a;
    layer0_outputs(3608) <= not (a xor b);
    layer0_outputs(3609) <= not b or a;
    layer0_outputs(3610) <= not b;
    layer0_outputs(3611) <= a or b;
    layer0_outputs(3612) <= a;
    layer0_outputs(3613) <= a or b;
    layer0_outputs(3614) <= not b or a;
    layer0_outputs(3615) <= not (a or b);
    layer0_outputs(3616) <= not a;
    layer0_outputs(3617) <= b and not a;
    layer0_outputs(3618) <= a or b;
    layer0_outputs(3619) <= not b or a;
    layer0_outputs(3620) <= not (a or b);
    layer0_outputs(3621) <= a or b;
    layer0_outputs(3622) <= a and not b;
    layer0_outputs(3623) <= b;
    layer0_outputs(3624) <= not a or b;
    layer0_outputs(3625) <= a or b;
    layer0_outputs(3626) <= not (a or b);
    layer0_outputs(3627) <= a;
    layer0_outputs(3628) <= a xor b;
    layer0_outputs(3629) <= a xor b;
    layer0_outputs(3630) <= a xor b;
    layer0_outputs(3631) <= not b or a;
    layer0_outputs(3632) <= b and not a;
    layer0_outputs(3633) <= not a;
    layer0_outputs(3634) <= not (a or b);
    layer0_outputs(3635) <= not b or a;
    layer0_outputs(3636) <= not (a or b);
    layer0_outputs(3637) <= a and not b;
    layer0_outputs(3638) <= b and not a;
    layer0_outputs(3639) <= a xor b;
    layer0_outputs(3640) <= not (a xor b);
    layer0_outputs(3641) <= not (a or b);
    layer0_outputs(3642) <= b;
    layer0_outputs(3643) <= not b;
    layer0_outputs(3644) <= not b;
    layer0_outputs(3645) <= not (a xor b);
    layer0_outputs(3646) <= a or b;
    layer0_outputs(3647) <= '0';
    layer0_outputs(3648) <= a or b;
    layer0_outputs(3649) <= not a;
    layer0_outputs(3650) <= a xor b;
    layer0_outputs(3651) <= b and not a;
    layer0_outputs(3652) <= a;
    layer0_outputs(3653) <= a xor b;
    layer0_outputs(3654) <= a and not b;
    layer0_outputs(3655) <= not b;
    layer0_outputs(3656) <= not (a or b);
    layer0_outputs(3657) <= not (a or b);
    layer0_outputs(3658) <= not (a or b);
    layer0_outputs(3659) <= a and b;
    layer0_outputs(3660) <= not a or b;
    layer0_outputs(3661) <= a xor b;
    layer0_outputs(3662) <= not a;
    layer0_outputs(3663) <= not a or b;
    layer0_outputs(3664) <= a xor b;
    layer0_outputs(3665) <= b;
    layer0_outputs(3666) <= not a or b;
    layer0_outputs(3667) <= not b or a;
    layer0_outputs(3668) <= not a or b;
    layer0_outputs(3669) <= not (a xor b);
    layer0_outputs(3670) <= a xor b;
    layer0_outputs(3671) <= not a or b;
    layer0_outputs(3672) <= not a;
    layer0_outputs(3673) <= a xor b;
    layer0_outputs(3674) <= a or b;
    layer0_outputs(3675) <= not (a xor b);
    layer0_outputs(3676) <= b;
    layer0_outputs(3677) <= a or b;
    layer0_outputs(3678) <= not a;
    layer0_outputs(3679) <= not b or a;
    layer0_outputs(3680) <= a xor b;
    layer0_outputs(3681) <= a and b;
    layer0_outputs(3682) <= not (a or b);
    layer0_outputs(3683) <= a;
    layer0_outputs(3684) <= not a;
    layer0_outputs(3685) <= not a;
    layer0_outputs(3686) <= a;
    layer0_outputs(3687) <= a xor b;
    layer0_outputs(3688) <= a;
    layer0_outputs(3689) <= not (a or b);
    layer0_outputs(3690) <= a and not b;
    layer0_outputs(3691) <= not (a or b);
    layer0_outputs(3692) <= not (a or b);
    layer0_outputs(3693) <= a;
    layer0_outputs(3694) <= b;
    layer0_outputs(3695) <= '1';
    layer0_outputs(3696) <= not b;
    layer0_outputs(3697) <= '1';
    layer0_outputs(3698) <= not b;
    layer0_outputs(3699) <= b;
    layer0_outputs(3700) <= a and b;
    layer0_outputs(3701) <= not a or b;
    layer0_outputs(3702) <= b and not a;
    layer0_outputs(3703) <= not (a or b);
    layer0_outputs(3704) <= not (a or b);
    layer0_outputs(3705) <= not (a xor b);
    layer0_outputs(3706) <= not b;
    layer0_outputs(3707) <= a or b;
    layer0_outputs(3708) <= a or b;
    layer0_outputs(3709) <= b and not a;
    layer0_outputs(3710) <= a or b;
    layer0_outputs(3711) <= not (a and b);
    layer0_outputs(3712) <= a and not b;
    layer0_outputs(3713) <= a xor b;
    layer0_outputs(3714) <= not (a or b);
    layer0_outputs(3715) <= not b or a;
    layer0_outputs(3716) <= a xor b;
    layer0_outputs(3717) <= b and not a;
    layer0_outputs(3718) <= not a or b;
    layer0_outputs(3719) <= a or b;
    layer0_outputs(3720) <= b and not a;
    layer0_outputs(3721) <= a;
    layer0_outputs(3722) <= not (a xor b);
    layer0_outputs(3723) <= a or b;
    layer0_outputs(3724) <= '1';
    layer0_outputs(3725) <= a xor b;
    layer0_outputs(3726) <= not (a or b);
    layer0_outputs(3727) <= not (a or b);
    layer0_outputs(3728) <= not (a or b);
    layer0_outputs(3729) <= a or b;
    layer0_outputs(3730) <= not (a or b);
    layer0_outputs(3731) <= a or b;
    layer0_outputs(3732) <= a and not b;
    layer0_outputs(3733) <= a or b;
    layer0_outputs(3734) <= not (a xor b);
    layer0_outputs(3735) <= '0';
    layer0_outputs(3736) <= a;
    layer0_outputs(3737) <= not a;
    layer0_outputs(3738) <= b;
    layer0_outputs(3739) <= b and not a;
    layer0_outputs(3740) <= a xor b;
    layer0_outputs(3741) <= not a or b;
    layer0_outputs(3742) <= not a;
    layer0_outputs(3743) <= a or b;
    layer0_outputs(3744) <= a or b;
    layer0_outputs(3745) <= a and not b;
    layer0_outputs(3746) <= b and not a;
    layer0_outputs(3747) <= not (a or b);
    layer0_outputs(3748) <= not (a or b);
    layer0_outputs(3749) <= not b or a;
    layer0_outputs(3750) <= a xor b;
    layer0_outputs(3751) <= not a;
    layer0_outputs(3752) <= not (a or b);
    layer0_outputs(3753) <= not (a and b);
    layer0_outputs(3754) <= a;
    layer0_outputs(3755) <= a;
    layer0_outputs(3756) <= a and not b;
    layer0_outputs(3757) <= not b or a;
    layer0_outputs(3758) <= not b;
    layer0_outputs(3759) <= a or b;
    layer0_outputs(3760) <= not a;
    layer0_outputs(3761) <= b and not a;
    layer0_outputs(3762) <= not (a or b);
    layer0_outputs(3763) <= a and not b;
    layer0_outputs(3764) <= not (a and b);
    layer0_outputs(3765) <= a or b;
    layer0_outputs(3766) <= not (a xor b);
    layer0_outputs(3767) <= not b;
    layer0_outputs(3768) <= not a;
    layer0_outputs(3769) <= b and not a;
    layer0_outputs(3770) <= not (a xor b);
    layer0_outputs(3771) <= a and not b;
    layer0_outputs(3772) <= b and not a;
    layer0_outputs(3773) <= a and b;
    layer0_outputs(3774) <= not (a or b);
    layer0_outputs(3775) <= b;
    layer0_outputs(3776) <= not (a xor b);
    layer0_outputs(3777) <= b;
    layer0_outputs(3778) <= not (a or b);
    layer0_outputs(3779) <= a xor b;
    layer0_outputs(3780) <= not (a xor b);
    layer0_outputs(3781) <= a;
    layer0_outputs(3782) <= a xor b;
    layer0_outputs(3783) <= b and not a;
    layer0_outputs(3784) <= '1';
    layer0_outputs(3785) <= a;
    layer0_outputs(3786) <= a;
    layer0_outputs(3787) <= a or b;
    layer0_outputs(3788) <= '1';
    layer0_outputs(3789) <= '1';
    layer0_outputs(3790) <= a xor b;
    layer0_outputs(3791) <= b and not a;
    layer0_outputs(3792) <= a or b;
    layer0_outputs(3793) <= a xor b;
    layer0_outputs(3794) <= not b;
    layer0_outputs(3795) <= not b;
    layer0_outputs(3796) <= not a;
    layer0_outputs(3797) <= a or b;
    layer0_outputs(3798) <= not (a xor b);
    layer0_outputs(3799) <= a or b;
    layer0_outputs(3800) <= a or b;
    layer0_outputs(3801) <= '1';
    layer0_outputs(3802) <= a xor b;
    layer0_outputs(3803) <= not a;
    layer0_outputs(3804) <= not b or a;
    layer0_outputs(3805) <= a xor b;
    layer0_outputs(3806) <= a xor b;
    layer0_outputs(3807) <= b;
    layer0_outputs(3808) <= a;
    layer0_outputs(3809) <= not (a xor b);
    layer0_outputs(3810) <= not b or a;
    layer0_outputs(3811) <= b and not a;
    layer0_outputs(3812) <= not (a and b);
    layer0_outputs(3813) <= not a or b;
    layer0_outputs(3814) <= a xor b;
    layer0_outputs(3815) <= not (a xor b);
    layer0_outputs(3816) <= a xor b;
    layer0_outputs(3817) <= not (a or b);
    layer0_outputs(3818) <= not (a or b);
    layer0_outputs(3819) <= a or b;
    layer0_outputs(3820) <= not (a xor b);
    layer0_outputs(3821) <= a and not b;
    layer0_outputs(3822) <= a and not b;
    layer0_outputs(3823) <= not (a or b);
    layer0_outputs(3824) <= not (a or b);
    layer0_outputs(3825) <= not a or b;
    layer0_outputs(3826) <= not a;
    layer0_outputs(3827) <= b;
    layer0_outputs(3828) <= '0';
    layer0_outputs(3829) <= a or b;
    layer0_outputs(3830) <= a and not b;
    layer0_outputs(3831) <= not b;
    layer0_outputs(3832) <= a xor b;
    layer0_outputs(3833) <= not (a or b);
    layer0_outputs(3834) <= b and not a;
    layer0_outputs(3835) <= not a;
    layer0_outputs(3836) <= not (a or b);
    layer0_outputs(3837) <= a xor b;
    layer0_outputs(3838) <= not (a xor b);
    layer0_outputs(3839) <= a or b;
    layer0_outputs(3840) <= not (a or b);
    layer0_outputs(3841) <= b and not a;
    layer0_outputs(3842) <= a xor b;
    layer0_outputs(3843) <= not (a or b);
    layer0_outputs(3844) <= not a;
    layer0_outputs(3845) <= not (a or b);
    layer0_outputs(3846) <= '0';
    layer0_outputs(3847) <= a and not b;
    layer0_outputs(3848) <= not (a or b);
    layer0_outputs(3849) <= a xor b;
    layer0_outputs(3850) <= not b;
    layer0_outputs(3851) <= b;
    layer0_outputs(3852) <= a or b;
    layer0_outputs(3853) <= not (a xor b);
    layer0_outputs(3854) <= not (a or b);
    layer0_outputs(3855) <= not a or b;
    layer0_outputs(3856) <= not (a and b);
    layer0_outputs(3857) <= not a;
    layer0_outputs(3858) <= not (a or b);
    layer0_outputs(3859) <= b;
    layer0_outputs(3860) <= b;
    layer0_outputs(3861) <= a and not b;
    layer0_outputs(3862) <= not b;
    layer0_outputs(3863) <= a or b;
    layer0_outputs(3864) <= not b;
    layer0_outputs(3865) <= not b;
    layer0_outputs(3866) <= not (a xor b);
    layer0_outputs(3867) <= not (a or b);
    layer0_outputs(3868) <= not (a or b);
    layer0_outputs(3869) <= b;
    layer0_outputs(3870) <= '1';
    layer0_outputs(3871) <= not (a xor b);
    layer0_outputs(3872) <= a;
    layer0_outputs(3873) <= a xor b;
    layer0_outputs(3874) <= not b or a;
    layer0_outputs(3875) <= a or b;
    layer0_outputs(3876) <= b and not a;
    layer0_outputs(3877) <= not (a and b);
    layer0_outputs(3878) <= not (a or b);
    layer0_outputs(3879) <= not (a xor b);
    layer0_outputs(3880) <= a xor b;
    layer0_outputs(3881) <= a;
    layer0_outputs(3882) <= not a;
    layer0_outputs(3883) <= not b;
    layer0_outputs(3884) <= not (a or b);
    layer0_outputs(3885) <= a or b;
    layer0_outputs(3886) <= a or b;
    layer0_outputs(3887) <= b;
    layer0_outputs(3888) <= not b;
    layer0_outputs(3889) <= a and not b;
    layer0_outputs(3890) <= not a or b;
    layer0_outputs(3891) <= not a or b;
    layer0_outputs(3892) <= not a or b;
    layer0_outputs(3893) <= not b;
    layer0_outputs(3894) <= not a or b;
    layer0_outputs(3895) <= a xor b;
    layer0_outputs(3896) <= not a or b;
    layer0_outputs(3897) <= not a;
    layer0_outputs(3898) <= a and b;
    layer0_outputs(3899) <= b and not a;
    layer0_outputs(3900) <= a;
    layer0_outputs(3901) <= not b or a;
    layer0_outputs(3902) <= not a or b;
    layer0_outputs(3903) <= not a or b;
    layer0_outputs(3904) <= not b;
    layer0_outputs(3905) <= not (a or b);
    layer0_outputs(3906) <= not b;
    layer0_outputs(3907) <= a and not b;
    layer0_outputs(3908) <= '0';
    layer0_outputs(3909) <= not a;
    layer0_outputs(3910) <= not (a or b);
    layer0_outputs(3911) <= not b;
    layer0_outputs(3912) <= a;
    layer0_outputs(3913) <= b;
    layer0_outputs(3914) <= a and not b;
    layer0_outputs(3915) <= not (a xor b);
    layer0_outputs(3916) <= not b;
    layer0_outputs(3917) <= a;
    layer0_outputs(3918) <= a or b;
    layer0_outputs(3919) <= not b or a;
    layer0_outputs(3920) <= a or b;
    layer0_outputs(3921) <= not a or b;
    layer0_outputs(3922) <= not (a and b);
    layer0_outputs(3923) <= not (a or b);
    layer0_outputs(3924) <= not b;
    layer0_outputs(3925) <= a and b;
    layer0_outputs(3926) <= not b or a;
    layer0_outputs(3927) <= not (a xor b);
    layer0_outputs(3928) <= not b;
    layer0_outputs(3929) <= not (a or b);
    layer0_outputs(3930) <= b and not a;
    layer0_outputs(3931) <= b and not a;
    layer0_outputs(3932) <= not (a or b);
    layer0_outputs(3933) <= a or b;
    layer0_outputs(3934) <= not a or b;
    layer0_outputs(3935) <= not (a xor b);
    layer0_outputs(3936) <= a or b;
    layer0_outputs(3937) <= a and not b;
    layer0_outputs(3938) <= not a or b;
    layer0_outputs(3939) <= '1';
    layer0_outputs(3940) <= a xor b;
    layer0_outputs(3941) <= not b;
    layer0_outputs(3942) <= not b or a;
    layer0_outputs(3943) <= a or b;
    layer0_outputs(3944) <= b;
    layer0_outputs(3945) <= a and not b;
    layer0_outputs(3946) <= a;
    layer0_outputs(3947) <= a and b;
    layer0_outputs(3948) <= not a;
    layer0_outputs(3949) <= not (a or b);
    layer0_outputs(3950) <= not (a xor b);
    layer0_outputs(3951) <= a or b;
    layer0_outputs(3952) <= not (a or b);
    layer0_outputs(3953) <= not (a xor b);
    layer0_outputs(3954) <= a;
    layer0_outputs(3955) <= a or b;
    layer0_outputs(3956) <= a xor b;
    layer0_outputs(3957) <= a or b;
    layer0_outputs(3958) <= not (a xor b);
    layer0_outputs(3959) <= not b;
    layer0_outputs(3960) <= not a or b;
    layer0_outputs(3961) <= a;
    layer0_outputs(3962) <= not a;
    layer0_outputs(3963) <= not (a or b);
    layer0_outputs(3964) <= a or b;
    layer0_outputs(3965) <= not a or b;
    layer0_outputs(3966) <= a xor b;
    layer0_outputs(3967) <= a;
    layer0_outputs(3968) <= not (a or b);
    layer0_outputs(3969) <= not (a xor b);
    layer0_outputs(3970) <= b and not a;
    layer0_outputs(3971) <= not a;
    layer0_outputs(3972) <= a xor b;
    layer0_outputs(3973) <= b and not a;
    layer0_outputs(3974) <= a xor b;
    layer0_outputs(3975) <= b and not a;
    layer0_outputs(3976) <= a;
    layer0_outputs(3977) <= not b or a;
    layer0_outputs(3978) <= a xor b;
    layer0_outputs(3979) <= not (a xor b);
    layer0_outputs(3980) <= not b or a;
    layer0_outputs(3981) <= not a or b;
    layer0_outputs(3982) <= not a or b;
    layer0_outputs(3983) <= b;
    layer0_outputs(3984) <= b and not a;
    layer0_outputs(3985) <= b and not a;
    layer0_outputs(3986) <= not a;
    layer0_outputs(3987) <= a and b;
    layer0_outputs(3988) <= not (a xor b);
    layer0_outputs(3989) <= a or b;
    layer0_outputs(3990) <= a xor b;
    layer0_outputs(3991) <= not b;
    layer0_outputs(3992) <= not (a or b);
    layer0_outputs(3993) <= a xor b;
    layer0_outputs(3994) <= not a or b;
    layer0_outputs(3995) <= b;
    layer0_outputs(3996) <= a or b;
    layer0_outputs(3997) <= not b;
    layer0_outputs(3998) <= a and not b;
    layer0_outputs(3999) <= b and not a;
    layer0_outputs(4000) <= b and not a;
    layer0_outputs(4001) <= a;
    layer0_outputs(4002) <= not (a xor b);
    layer0_outputs(4003) <= a xor b;
    layer0_outputs(4004) <= a;
    layer0_outputs(4005) <= a or b;
    layer0_outputs(4006) <= b;
    layer0_outputs(4007) <= not a or b;
    layer0_outputs(4008) <= not a;
    layer0_outputs(4009) <= a;
    layer0_outputs(4010) <= a and b;
    layer0_outputs(4011) <= not a;
    layer0_outputs(4012) <= a and not b;
    layer0_outputs(4013) <= a and not b;
    layer0_outputs(4014) <= not a;
    layer0_outputs(4015) <= a xor b;
    layer0_outputs(4016) <= not (a and b);
    layer0_outputs(4017) <= not a;
    layer0_outputs(4018) <= not b;
    layer0_outputs(4019) <= not (a and b);
    layer0_outputs(4020) <= not (a or b);
    layer0_outputs(4021) <= not b;
    layer0_outputs(4022) <= '1';
    layer0_outputs(4023) <= not b or a;
    layer0_outputs(4024) <= b;
    layer0_outputs(4025) <= not b or a;
    layer0_outputs(4026) <= not (a or b);
    layer0_outputs(4027) <= not (a or b);
    layer0_outputs(4028) <= a and not b;
    layer0_outputs(4029) <= not (a or b);
    layer0_outputs(4030) <= not (a or b);
    layer0_outputs(4031) <= not (a or b);
    layer0_outputs(4032) <= not (a and b);
    layer0_outputs(4033) <= not a or b;
    layer0_outputs(4034) <= a or b;
    layer0_outputs(4035) <= not (a xor b);
    layer0_outputs(4036) <= not a or b;
    layer0_outputs(4037) <= not a;
    layer0_outputs(4038) <= a xor b;
    layer0_outputs(4039) <= a or b;
    layer0_outputs(4040) <= b;
    layer0_outputs(4041) <= a and not b;
    layer0_outputs(4042) <= b;
    layer0_outputs(4043) <= a xor b;
    layer0_outputs(4044) <= a or b;
    layer0_outputs(4045) <= a and b;
    layer0_outputs(4046) <= a or b;
    layer0_outputs(4047) <= a or b;
    layer0_outputs(4048) <= not (a xor b);
    layer0_outputs(4049) <= not (a xor b);
    layer0_outputs(4050) <= a xor b;
    layer0_outputs(4051) <= not (a xor b);
    layer0_outputs(4052) <= b;
    layer0_outputs(4053) <= not a or b;
    layer0_outputs(4054) <= a xor b;
    layer0_outputs(4055) <= '0';
    layer0_outputs(4056) <= b;
    layer0_outputs(4057) <= a xor b;
    layer0_outputs(4058) <= not a or b;
    layer0_outputs(4059) <= not (a or b);
    layer0_outputs(4060) <= a or b;
    layer0_outputs(4061) <= not a or b;
    layer0_outputs(4062) <= a xor b;
    layer0_outputs(4063) <= not a;
    layer0_outputs(4064) <= a and not b;
    layer0_outputs(4065) <= not (a xor b);
    layer0_outputs(4066) <= not a;
    layer0_outputs(4067) <= '1';
    layer0_outputs(4068) <= a or b;
    layer0_outputs(4069) <= b;
    layer0_outputs(4070) <= a and b;
    layer0_outputs(4071) <= not (a or b);
    layer0_outputs(4072) <= a;
    layer0_outputs(4073) <= not (a or b);
    layer0_outputs(4074) <= a xor b;
    layer0_outputs(4075) <= a;
    layer0_outputs(4076) <= not (a or b);
    layer0_outputs(4077) <= a or b;
    layer0_outputs(4078) <= b;
    layer0_outputs(4079) <= not (a or b);
    layer0_outputs(4080) <= not (a or b);
    layer0_outputs(4081) <= a xor b;
    layer0_outputs(4082) <= b and not a;
    layer0_outputs(4083) <= not a;
    layer0_outputs(4084) <= not (a xor b);
    layer0_outputs(4085) <= not (a and b);
    layer0_outputs(4086) <= a;
    layer0_outputs(4087) <= '1';
    layer0_outputs(4088) <= not b or a;
    layer0_outputs(4089) <= not (a xor b);
    layer0_outputs(4090) <= not (a xor b);
    layer0_outputs(4091) <= not (a xor b);
    layer0_outputs(4092) <= not (a or b);
    layer0_outputs(4093) <= not b;
    layer0_outputs(4094) <= a;
    layer0_outputs(4095) <= not b;
    layer0_outputs(4096) <= '0';
    layer0_outputs(4097) <= a and not b;
    layer0_outputs(4098) <= not a or b;
    layer0_outputs(4099) <= b and not a;
    layer0_outputs(4100) <= not b;
    layer0_outputs(4101) <= '0';
    layer0_outputs(4102) <= a;
    layer0_outputs(4103) <= not a or b;
    layer0_outputs(4104) <= a;
    layer0_outputs(4105) <= not (a xor b);
    layer0_outputs(4106) <= not a or b;
    layer0_outputs(4107) <= not b;
    layer0_outputs(4108) <= a;
    layer0_outputs(4109) <= a and not b;
    layer0_outputs(4110) <= not (a xor b);
    layer0_outputs(4111) <= a xor b;
    layer0_outputs(4112) <= b;
    layer0_outputs(4113) <= a xor b;
    layer0_outputs(4114) <= not a;
    layer0_outputs(4115) <= not b or a;
    layer0_outputs(4116) <= b and not a;
    layer0_outputs(4117) <= a or b;
    layer0_outputs(4118) <= not (a or b);
    layer0_outputs(4119) <= a and not b;
    layer0_outputs(4120) <= a xor b;
    layer0_outputs(4121) <= a and b;
    layer0_outputs(4122) <= not a or b;
    layer0_outputs(4123) <= a xor b;
    layer0_outputs(4124) <= not a or b;
    layer0_outputs(4125) <= a and b;
    layer0_outputs(4126) <= not b;
    layer0_outputs(4127) <= b and not a;
    layer0_outputs(4128) <= not a;
    layer0_outputs(4129) <= b and not a;
    layer0_outputs(4130) <= b and not a;
    layer0_outputs(4131) <= a or b;
    layer0_outputs(4132) <= a and b;
    layer0_outputs(4133) <= not (a and b);
    layer0_outputs(4134) <= b and not a;
    layer0_outputs(4135) <= b;
    layer0_outputs(4136) <= b and not a;
    layer0_outputs(4137) <= b and not a;
    layer0_outputs(4138) <= not a or b;
    layer0_outputs(4139) <= not (a xor b);
    layer0_outputs(4140) <= a and not b;
    layer0_outputs(4141) <= not b or a;
    layer0_outputs(4142) <= not b or a;
    layer0_outputs(4143) <= a;
    layer0_outputs(4144) <= not b or a;
    layer0_outputs(4145) <= not (a or b);
    layer0_outputs(4146) <= a;
    layer0_outputs(4147) <= a;
    layer0_outputs(4148) <= a and b;
    layer0_outputs(4149) <= not a;
    layer0_outputs(4150) <= a and not b;
    layer0_outputs(4151) <= not a or b;
    layer0_outputs(4152) <= not b;
    layer0_outputs(4153) <= not (a xor b);
    layer0_outputs(4154) <= a;
    layer0_outputs(4155) <= not (a xor b);
    layer0_outputs(4156) <= a xor b;
    layer0_outputs(4157) <= a;
    layer0_outputs(4158) <= not (a or b);
    layer0_outputs(4159) <= a;
    layer0_outputs(4160) <= not a or b;
    layer0_outputs(4161) <= a;
    layer0_outputs(4162) <= not b or a;
    layer0_outputs(4163) <= not a;
    layer0_outputs(4164) <= not b;
    layer0_outputs(4165) <= not (a and b);
    layer0_outputs(4166) <= not b;
    layer0_outputs(4167) <= not (a or b);
    layer0_outputs(4168) <= not (a xor b);
    layer0_outputs(4169) <= not a or b;
    layer0_outputs(4170) <= not b or a;
    layer0_outputs(4171) <= a or b;
    layer0_outputs(4172) <= a or b;
    layer0_outputs(4173) <= not a or b;
    layer0_outputs(4174) <= not (a or b);
    layer0_outputs(4175) <= a or b;
    layer0_outputs(4176) <= '0';
    layer0_outputs(4177) <= not (a xor b);
    layer0_outputs(4178) <= not a;
    layer0_outputs(4179) <= not a or b;
    layer0_outputs(4180) <= not (a or b);
    layer0_outputs(4181) <= not (a xor b);
    layer0_outputs(4182) <= not b or a;
    layer0_outputs(4183) <= a xor b;
    layer0_outputs(4184) <= not b or a;
    layer0_outputs(4185) <= a or b;
    layer0_outputs(4186) <= '0';
    layer0_outputs(4187) <= a and not b;
    layer0_outputs(4188) <= not (a xor b);
    layer0_outputs(4189) <= not a or b;
    layer0_outputs(4190) <= a or b;
    layer0_outputs(4191) <= a or b;
    layer0_outputs(4192) <= not (a xor b);
    layer0_outputs(4193) <= a;
    layer0_outputs(4194) <= not (a or b);
    layer0_outputs(4195) <= a;
    layer0_outputs(4196) <= a xor b;
    layer0_outputs(4197) <= a xor b;
    layer0_outputs(4198) <= not (a xor b);
    layer0_outputs(4199) <= a;
    layer0_outputs(4200) <= a or b;
    layer0_outputs(4201) <= not a;
    layer0_outputs(4202) <= '0';
    layer0_outputs(4203) <= '0';
    layer0_outputs(4204) <= b;
    layer0_outputs(4205) <= a;
    layer0_outputs(4206) <= not (a xor b);
    layer0_outputs(4207) <= a or b;
    layer0_outputs(4208) <= b;
    layer0_outputs(4209) <= a or b;
    layer0_outputs(4210) <= not (a xor b);
    layer0_outputs(4211) <= not (a or b);
    layer0_outputs(4212) <= not (a or b);
    layer0_outputs(4213) <= not a;
    layer0_outputs(4214) <= a and not b;
    layer0_outputs(4215) <= a or b;
    layer0_outputs(4216) <= a and not b;
    layer0_outputs(4217) <= b;
    layer0_outputs(4218) <= not (a or b);
    layer0_outputs(4219) <= not (a or b);
    layer0_outputs(4220) <= not a or b;
    layer0_outputs(4221) <= not b;
    layer0_outputs(4222) <= a xor b;
    layer0_outputs(4223) <= not b;
    layer0_outputs(4224) <= not (a or b);
    layer0_outputs(4225) <= not b;
    layer0_outputs(4226) <= a and not b;
    layer0_outputs(4227) <= not (a or b);
    layer0_outputs(4228) <= not (a or b);
    layer0_outputs(4229) <= b;
    layer0_outputs(4230) <= not (a or b);
    layer0_outputs(4231) <= a xor b;
    layer0_outputs(4232) <= a or b;
    layer0_outputs(4233) <= a or b;
    layer0_outputs(4234) <= not (a or b);
    layer0_outputs(4235) <= not a;
    layer0_outputs(4236) <= '1';
    layer0_outputs(4237) <= not (a or b);
    layer0_outputs(4238) <= '1';
    layer0_outputs(4239) <= a;
    layer0_outputs(4240) <= a and not b;
    layer0_outputs(4241) <= a or b;
    layer0_outputs(4242) <= not b or a;
    layer0_outputs(4243) <= a or b;
    layer0_outputs(4244) <= not b or a;
    layer0_outputs(4245) <= a xor b;
    layer0_outputs(4246) <= not b;
    layer0_outputs(4247) <= not a;
    layer0_outputs(4248) <= b;
    layer0_outputs(4249) <= not a;
    layer0_outputs(4250) <= a and not b;
    layer0_outputs(4251) <= b;
    layer0_outputs(4252) <= not b;
    layer0_outputs(4253) <= not (a or b);
    layer0_outputs(4254) <= not b;
    layer0_outputs(4255) <= not (a or b);
    layer0_outputs(4256) <= not (a xor b);
    layer0_outputs(4257) <= not (a xor b);
    layer0_outputs(4258) <= a and not b;
    layer0_outputs(4259) <= a and b;
    layer0_outputs(4260) <= not a or b;
    layer0_outputs(4261) <= not (a or b);
    layer0_outputs(4262) <= a and not b;
    layer0_outputs(4263) <= not a;
    layer0_outputs(4264) <= a xor b;
    layer0_outputs(4265) <= a or b;
    layer0_outputs(4266) <= a xor b;
    layer0_outputs(4267) <= a or b;
    layer0_outputs(4268) <= a xor b;
    layer0_outputs(4269) <= not (a xor b);
    layer0_outputs(4270) <= not (a xor b);
    layer0_outputs(4271) <= '1';
    layer0_outputs(4272) <= not b or a;
    layer0_outputs(4273) <= a and not b;
    layer0_outputs(4274) <= not a;
    layer0_outputs(4275) <= b and not a;
    layer0_outputs(4276) <= not (a or b);
    layer0_outputs(4277) <= a or b;
    layer0_outputs(4278) <= a;
    layer0_outputs(4279) <= not b or a;
    layer0_outputs(4280) <= not (a or b);
    layer0_outputs(4281) <= a;
    layer0_outputs(4282) <= not a;
    layer0_outputs(4283) <= not (a or b);
    layer0_outputs(4284) <= not b or a;
    layer0_outputs(4285) <= '1';
    layer0_outputs(4286) <= a and b;
    layer0_outputs(4287) <= a or b;
    layer0_outputs(4288) <= not b or a;
    layer0_outputs(4289) <= a;
    layer0_outputs(4290) <= not (a and b);
    layer0_outputs(4291) <= '0';
    layer0_outputs(4292) <= a xor b;
    layer0_outputs(4293) <= not b or a;
    layer0_outputs(4294) <= not a or b;
    layer0_outputs(4295) <= a and not b;
    layer0_outputs(4296) <= a or b;
    layer0_outputs(4297) <= a and b;
    layer0_outputs(4298) <= not b;
    layer0_outputs(4299) <= b;
    layer0_outputs(4300) <= a or b;
    layer0_outputs(4301) <= not a;
    layer0_outputs(4302) <= a xor b;
    layer0_outputs(4303) <= a and not b;
    layer0_outputs(4304) <= a or b;
    layer0_outputs(4305) <= not (a or b);
    layer0_outputs(4306) <= not (a or b);
    layer0_outputs(4307) <= a or b;
    layer0_outputs(4308) <= b;
    layer0_outputs(4309) <= not b;
    layer0_outputs(4310) <= not b or a;
    layer0_outputs(4311) <= not (a xor b);
    layer0_outputs(4312) <= not (a or b);
    layer0_outputs(4313) <= not b or a;
    layer0_outputs(4314) <= not (a xor b);
    layer0_outputs(4315) <= a and not b;
    layer0_outputs(4316) <= not (a xor b);
    layer0_outputs(4317) <= not (a or b);
    layer0_outputs(4318) <= not a or b;
    layer0_outputs(4319) <= not a or b;
    layer0_outputs(4320) <= not (a xor b);
    layer0_outputs(4321) <= not a;
    layer0_outputs(4322) <= not (a or b);
    layer0_outputs(4323) <= not a;
    layer0_outputs(4324) <= not (a xor b);
    layer0_outputs(4325) <= not a or b;
    layer0_outputs(4326) <= b;
    layer0_outputs(4327) <= not a;
    layer0_outputs(4328) <= not (a or b);
    layer0_outputs(4329) <= '0';
    layer0_outputs(4330) <= b and not a;
    layer0_outputs(4331) <= a xor b;
    layer0_outputs(4332) <= a and not b;
    layer0_outputs(4333) <= not (a xor b);
    layer0_outputs(4334) <= not a;
    layer0_outputs(4335) <= b;
    layer0_outputs(4336) <= a and not b;
    layer0_outputs(4337) <= b and not a;
    layer0_outputs(4338) <= a or b;
    layer0_outputs(4339) <= not a or b;
    layer0_outputs(4340) <= a;
    layer0_outputs(4341) <= not a;
    layer0_outputs(4342) <= a or b;
    layer0_outputs(4343) <= a or b;
    layer0_outputs(4344) <= b and not a;
    layer0_outputs(4345) <= not (a or b);
    layer0_outputs(4346) <= not b;
    layer0_outputs(4347) <= a or b;
    layer0_outputs(4348) <= not (a or b);
    layer0_outputs(4349) <= a or b;
    layer0_outputs(4350) <= not a or b;
    layer0_outputs(4351) <= a or b;
    layer0_outputs(4352) <= a;
    layer0_outputs(4353) <= b and not a;
    layer0_outputs(4354) <= not b;
    layer0_outputs(4355) <= not a;
    layer0_outputs(4356) <= '0';
    layer0_outputs(4357) <= a xor b;
    layer0_outputs(4358) <= not b or a;
    layer0_outputs(4359) <= not b;
    layer0_outputs(4360) <= not (a or b);
    layer0_outputs(4361) <= a;
    layer0_outputs(4362) <= a or b;
    layer0_outputs(4363) <= not a;
    layer0_outputs(4364) <= a;
    layer0_outputs(4365) <= a xor b;
    layer0_outputs(4366) <= a xor b;
    layer0_outputs(4367) <= not (a or b);
    layer0_outputs(4368) <= not (a or b);
    layer0_outputs(4369) <= '0';
    layer0_outputs(4370) <= a or b;
    layer0_outputs(4371) <= b;
    layer0_outputs(4372) <= a;
    layer0_outputs(4373) <= not (a xor b);
    layer0_outputs(4374) <= not (a or b);
    layer0_outputs(4375) <= not (a xor b);
    layer0_outputs(4376) <= not (a or b);
    layer0_outputs(4377) <= b;
    layer0_outputs(4378) <= not (a xor b);
    layer0_outputs(4379) <= not (a or b);
    layer0_outputs(4380) <= b and not a;
    layer0_outputs(4381) <= not b or a;
    layer0_outputs(4382) <= not b;
    layer0_outputs(4383) <= not b;
    layer0_outputs(4384) <= not a;
    layer0_outputs(4385) <= not b or a;
    layer0_outputs(4386) <= not b or a;
    layer0_outputs(4387) <= not b;
    layer0_outputs(4388) <= a or b;
    layer0_outputs(4389) <= a and not b;
    layer0_outputs(4390) <= a xor b;
    layer0_outputs(4391) <= b and not a;
    layer0_outputs(4392) <= not b;
    layer0_outputs(4393) <= a;
    layer0_outputs(4394) <= a xor b;
    layer0_outputs(4395) <= not a or b;
    layer0_outputs(4396) <= not a or b;
    layer0_outputs(4397) <= a or b;
    layer0_outputs(4398) <= not a or b;
    layer0_outputs(4399) <= not a or b;
    layer0_outputs(4400) <= b;
    layer0_outputs(4401) <= a xor b;
    layer0_outputs(4402) <= not a;
    layer0_outputs(4403) <= not a or b;
    layer0_outputs(4404) <= b and not a;
    layer0_outputs(4405) <= a xor b;
    layer0_outputs(4406) <= a;
    layer0_outputs(4407) <= not a;
    layer0_outputs(4408) <= a;
    layer0_outputs(4409) <= a xor b;
    layer0_outputs(4410) <= not (a xor b);
    layer0_outputs(4411) <= a or b;
    layer0_outputs(4412) <= not a;
    layer0_outputs(4413) <= not (a xor b);
    layer0_outputs(4414) <= not b or a;
    layer0_outputs(4415) <= not b or a;
    layer0_outputs(4416) <= a xor b;
    layer0_outputs(4417) <= not a;
    layer0_outputs(4418) <= a or b;
    layer0_outputs(4419) <= not b or a;
    layer0_outputs(4420) <= not (a xor b);
    layer0_outputs(4421) <= b and not a;
    layer0_outputs(4422) <= a;
    layer0_outputs(4423) <= a xor b;
    layer0_outputs(4424) <= a or b;
    layer0_outputs(4425) <= b and not a;
    layer0_outputs(4426) <= not a;
    layer0_outputs(4427) <= not (a or b);
    layer0_outputs(4428) <= b;
    layer0_outputs(4429) <= a or b;
    layer0_outputs(4430) <= not (a xor b);
    layer0_outputs(4431) <= not (a xor b);
    layer0_outputs(4432) <= b and not a;
    layer0_outputs(4433) <= not b or a;
    layer0_outputs(4434) <= not a;
    layer0_outputs(4435) <= a or b;
    layer0_outputs(4436) <= a xor b;
    layer0_outputs(4437) <= not (a or b);
    layer0_outputs(4438) <= not (a or b);
    layer0_outputs(4439) <= not b or a;
    layer0_outputs(4440) <= not a;
    layer0_outputs(4441) <= not a or b;
    layer0_outputs(4442) <= not a or b;
    layer0_outputs(4443) <= not (a xor b);
    layer0_outputs(4444) <= a and not b;
    layer0_outputs(4445) <= a xor b;
    layer0_outputs(4446) <= not b;
    layer0_outputs(4447) <= a xor b;
    layer0_outputs(4448) <= not b;
    layer0_outputs(4449) <= a xor b;
    layer0_outputs(4450) <= a and not b;
    layer0_outputs(4451) <= not b or a;
    layer0_outputs(4452) <= b;
    layer0_outputs(4453) <= a xor b;
    layer0_outputs(4454) <= a and not b;
    layer0_outputs(4455) <= b;
    layer0_outputs(4456) <= not (a xor b);
    layer0_outputs(4457) <= a and not b;
    layer0_outputs(4458) <= not (a or b);
    layer0_outputs(4459) <= not b or a;
    layer0_outputs(4460) <= b;
    layer0_outputs(4461) <= a and b;
    layer0_outputs(4462) <= not a or b;
    layer0_outputs(4463) <= not b or a;
    layer0_outputs(4464) <= a xor b;
    layer0_outputs(4465) <= a and b;
    layer0_outputs(4466) <= not a;
    layer0_outputs(4467) <= a;
    layer0_outputs(4468) <= b;
    layer0_outputs(4469) <= a and not b;
    layer0_outputs(4470) <= not a;
    layer0_outputs(4471) <= a or b;
    layer0_outputs(4472) <= a and not b;
    layer0_outputs(4473) <= not (a or b);
    layer0_outputs(4474) <= a or b;
    layer0_outputs(4475) <= a xor b;
    layer0_outputs(4476) <= a;
    layer0_outputs(4477) <= a or b;
    layer0_outputs(4478) <= a or b;
    layer0_outputs(4479) <= a xor b;
    layer0_outputs(4480) <= not b or a;
    layer0_outputs(4481) <= not a;
    layer0_outputs(4482) <= not (a xor b);
    layer0_outputs(4483) <= '0';
    layer0_outputs(4484) <= a and not b;
    layer0_outputs(4485) <= not b;
    layer0_outputs(4486) <= a and not b;
    layer0_outputs(4487) <= not (a or b);
    layer0_outputs(4488) <= not (a and b);
    layer0_outputs(4489) <= a or b;
    layer0_outputs(4490) <= '0';
    layer0_outputs(4491) <= not (a or b);
    layer0_outputs(4492) <= a and not b;
    layer0_outputs(4493) <= a or b;
    layer0_outputs(4494) <= a and not b;
    layer0_outputs(4495) <= '0';
    layer0_outputs(4496) <= a;
    layer0_outputs(4497) <= a and not b;
    layer0_outputs(4498) <= a or b;
    layer0_outputs(4499) <= not (a or b);
    layer0_outputs(4500) <= not (a or b);
    layer0_outputs(4501) <= not (a xor b);
    layer0_outputs(4502) <= a;
    layer0_outputs(4503) <= a or b;
    layer0_outputs(4504) <= not (a and b);
    layer0_outputs(4505) <= not (a and b);
    layer0_outputs(4506) <= not (a or b);
    layer0_outputs(4507) <= not (a and b);
    layer0_outputs(4508) <= b;
    layer0_outputs(4509) <= b;
    layer0_outputs(4510) <= a xor b;
    layer0_outputs(4511) <= a;
    layer0_outputs(4512) <= not b;
    layer0_outputs(4513) <= not a or b;
    layer0_outputs(4514) <= a and not b;
    layer0_outputs(4515) <= a xor b;
    layer0_outputs(4516) <= not (a xor b);
    layer0_outputs(4517) <= not b or a;
    layer0_outputs(4518) <= not (a xor b);
    layer0_outputs(4519) <= a;
    layer0_outputs(4520) <= not a or b;
    layer0_outputs(4521) <= b and not a;
    layer0_outputs(4522) <= not (a or b);
    layer0_outputs(4523) <= not b;
    layer0_outputs(4524) <= not (a and b);
    layer0_outputs(4525) <= a;
    layer0_outputs(4526) <= not a;
    layer0_outputs(4527) <= a or b;
    layer0_outputs(4528) <= b;
    layer0_outputs(4529) <= not b or a;
    layer0_outputs(4530) <= not b;
    layer0_outputs(4531) <= a xor b;
    layer0_outputs(4532) <= b;
    layer0_outputs(4533) <= a and not b;
    layer0_outputs(4534) <= not (a or b);
    layer0_outputs(4535) <= not (a or b);
    layer0_outputs(4536) <= not (a or b);
    layer0_outputs(4537) <= a and not b;
    layer0_outputs(4538) <= a or b;
    layer0_outputs(4539) <= not (a or b);
    layer0_outputs(4540) <= not b or a;
    layer0_outputs(4541) <= not (a or b);
    layer0_outputs(4542) <= a or b;
    layer0_outputs(4543) <= not b or a;
    layer0_outputs(4544) <= '0';
    layer0_outputs(4545) <= a;
    layer0_outputs(4546) <= b and not a;
    layer0_outputs(4547) <= not (a xor b);
    layer0_outputs(4548) <= a xor b;
    layer0_outputs(4549) <= a or b;
    layer0_outputs(4550) <= a and not b;
    layer0_outputs(4551) <= not b;
    layer0_outputs(4552) <= b;
    layer0_outputs(4553) <= a and b;
    layer0_outputs(4554) <= not b or a;
    layer0_outputs(4555) <= not (a xor b);
    layer0_outputs(4556) <= a or b;
    layer0_outputs(4557) <= not b or a;
    layer0_outputs(4558) <= not (a or b);
    layer0_outputs(4559) <= not a;
    layer0_outputs(4560) <= not b or a;
    layer0_outputs(4561) <= not a;
    layer0_outputs(4562) <= a xor b;
    layer0_outputs(4563) <= not b or a;
    layer0_outputs(4564) <= not b;
    layer0_outputs(4565) <= not (a or b);
    layer0_outputs(4566) <= b;
    layer0_outputs(4567) <= a xor b;
    layer0_outputs(4568) <= not (a or b);
    layer0_outputs(4569) <= b;
    layer0_outputs(4570) <= not a;
    layer0_outputs(4571) <= a and not b;
    layer0_outputs(4572) <= b;
    layer0_outputs(4573) <= b and not a;
    layer0_outputs(4574) <= '0';
    layer0_outputs(4575) <= not b or a;
    layer0_outputs(4576) <= a xor b;
    layer0_outputs(4577) <= b;
    layer0_outputs(4578) <= not a;
    layer0_outputs(4579) <= not (a or b);
    layer0_outputs(4580) <= not a or b;
    layer0_outputs(4581) <= not (a xor b);
    layer0_outputs(4582) <= not a or b;
    layer0_outputs(4583) <= a and not b;
    layer0_outputs(4584) <= a and b;
    layer0_outputs(4585) <= a;
    layer0_outputs(4586) <= a xor b;
    layer0_outputs(4587) <= a xor b;
    layer0_outputs(4588) <= not b;
    layer0_outputs(4589) <= a xor b;
    layer0_outputs(4590) <= not b or a;
    layer0_outputs(4591) <= not b or a;
    layer0_outputs(4592) <= not a or b;
    layer0_outputs(4593) <= a xor b;
    layer0_outputs(4594) <= not b or a;
    layer0_outputs(4595) <= a or b;
    layer0_outputs(4596) <= a and not b;
    layer0_outputs(4597) <= not b or a;
    layer0_outputs(4598) <= a and not b;
    layer0_outputs(4599) <= b;
    layer0_outputs(4600) <= not a or b;
    layer0_outputs(4601) <= not (a xor b);
    layer0_outputs(4602) <= a xor b;
    layer0_outputs(4603) <= a or b;
    layer0_outputs(4604) <= not a or b;
    layer0_outputs(4605) <= a or b;
    layer0_outputs(4606) <= not b;
    layer0_outputs(4607) <= not (a or b);
    layer0_outputs(4608) <= not (a or b);
    layer0_outputs(4609) <= b and not a;
    layer0_outputs(4610) <= b and not a;
    layer0_outputs(4611) <= b;
    layer0_outputs(4612) <= not (a xor b);
    layer0_outputs(4613) <= '1';
    layer0_outputs(4614) <= a or b;
    layer0_outputs(4615) <= not a;
    layer0_outputs(4616) <= not (a or b);
    layer0_outputs(4617) <= not a or b;
    layer0_outputs(4618) <= b;
    layer0_outputs(4619) <= b and not a;
    layer0_outputs(4620) <= a xor b;
    layer0_outputs(4621) <= b and not a;
    layer0_outputs(4622) <= not b or a;
    layer0_outputs(4623) <= not a or b;
    layer0_outputs(4624) <= not b;
    layer0_outputs(4625) <= not b;
    layer0_outputs(4626) <= a;
    layer0_outputs(4627) <= b and not a;
    layer0_outputs(4628) <= a and not b;
    layer0_outputs(4629) <= not a or b;
    layer0_outputs(4630) <= a;
    layer0_outputs(4631) <= not b;
    layer0_outputs(4632) <= not a;
    layer0_outputs(4633) <= b and not a;
    layer0_outputs(4634) <= not (a xor b);
    layer0_outputs(4635) <= not (a or b);
    layer0_outputs(4636) <= not (a xor b);
    layer0_outputs(4637) <= a;
    layer0_outputs(4638) <= '1';
    layer0_outputs(4639) <= not b or a;
    layer0_outputs(4640) <= a or b;
    layer0_outputs(4641) <= a or b;
    layer0_outputs(4642) <= b;
    layer0_outputs(4643) <= not a or b;
    layer0_outputs(4644) <= a and b;
    layer0_outputs(4645) <= '0';
    layer0_outputs(4646) <= not (a xor b);
    layer0_outputs(4647) <= b;
    layer0_outputs(4648) <= a and not b;
    layer0_outputs(4649) <= b;
    layer0_outputs(4650) <= a or b;
    layer0_outputs(4651) <= not (a xor b);
    layer0_outputs(4652) <= '0';
    layer0_outputs(4653) <= a and not b;
    layer0_outputs(4654) <= a;
    layer0_outputs(4655) <= not (a xor b);
    layer0_outputs(4656) <= a xor b;
    layer0_outputs(4657) <= a and not b;
    layer0_outputs(4658) <= not (a xor b);
    layer0_outputs(4659) <= not (a xor b);
    layer0_outputs(4660) <= a and b;
    layer0_outputs(4661) <= '1';
    layer0_outputs(4662) <= a xor b;
    layer0_outputs(4663) <= not (a xor b);
    layer0_outputs(4664) <= not (a or b);
    layer0_outputs(4665) <= a xor b;
    layer0_outputs(4666) <= not b;
    layer0_outputs(4667) <= a or b;
    layer0_outputs(4668) <= a;
    layer0_outputs(4669) <= '1';
    layer0_outputs(4670) <= b;
    layer0_outputs(4671) <= a and not b;
    layer0_outputs(4672) <= not a or b;
    layer0_outputs(4673) <= a and b;
    layer0_outputs(4674) <= a;
    layer0_outputs(4675) <= b;
    layer0_outputs(4676) <= b and not a;
    layer0_outputs(4677) <= not a;
    layer0_outputs(4678) <= not a or b;
    layer0_outputs(4679) <= a or b;
    layer0_outputs(4680) <= not a;
    layer0_outputs(4681) <= a and not b;
    layer0_outputs(4682) <= a or b;
    layer0_outputs(4683) <= not a;
    layer0_outputs(4684) <= not (a or b);
    layer0_outputs(4685) <= a and not b;
    layer0_outputs(4686) <= a or b;
    layer0_outputs(4687) <= not b;
    layer0_outputs(4688) <= a or b;
    layer0_outputs(4689) <= not b or a;
    layer0_outputs(4690) <= not b;
    layer0_outputs(4691) <= not (a or b);
    layer0_outputs(4692) <= not a;
    layer0_outputs(4693) <= not a;
    layer0_outputs(4694) <= not (a xor b);
    layer0_outputs(4695) <= a or b;
    layer0_outputs(4696) <= a or b;
    layer0_outputs(4697) <= a and not b;
    layer0_outputs(4698) <= a or b;
    layer0_outputs(4699) <= not (a xor b);
    layer0_outputs(4700) <= not b;
    layer0_outputs(4701) <= a and not b;
    layer0_outputs(4702) <= not (a and b);
    layer0_outputs(4703) <= a xor b;
    layer0_outputs(4704) <= not b or a;
    layer0_outputs(4705) <= a and not b;
    layer0_outputs(4706) <= a or b;
    layer0_outputs(4707) <= not (a or b);
    layer0_outputs(4708) <= b;
    layer0_outputs(4709) <= a or b;
    layer0_outputs(4710) <= not (a or b);
    layer0_outputs(4711) <= a and not b;
    layer0_outputs(4712) <= b;
    layer0_outputs(4713) <= not (a xor b);
    layer0_outputs(4714) <= not a;
    layer0_outputs(4715) <= not b;
    layer0_outputs(4716) <= b;
    layer0_outputs(4717) <= '0';
    layer0_outputs(4718) <= a and not b;
    layer0_outputs(4719) <= not (a or b);
    layer0_outputs(4720) <= a and not b;
    layer0_outputs(4721) <= a xor b;
    layer0_outputs(4722) <= a or b;
    layer0_outputs(4723) <= '0';
    layer0_outputs(4724) <= not a or b;
    layer0_outputs(4725) <= not b or a;
    layer0_outputs(4726) <= a xor b;
    layer0_outputs(4727) <= not b or a;
    layer0_outputs(4728) <= b;
    layer0_outputs(4729) <= b;
    layer0_outputs(4730) <= not (a xor b);
    layer0_outputs(4731) <= a xor b;
    layer0_outputs(4732) <= a xor b;
    layer0_outputs(4733) <= not a or b;
    layer0_outputs(4734) <= b and not a;
    layer0_outputs(4735) <= not a;
    layer0_outputs(4736) <= not (a xor b);
    layer0_outputs(4737) <= a or b;
    layer0_outputs(4738) <= a xor b;
    layer0_outputs(4739) <= a;
    layer0_outputs(4740) <= a and b;
    layer0_outputs(4741) <= a;
    layer0_outputs(4742) <= not (a xor b);
    layer0_outputs(4743) <= b and not a;
    layer0_outputs(4744) <= not b;
    layer0_outputs(4745) <= not a or b;
    layer0_outputs(4746) <= not (a or b);
    layer0_outputs(4747) <= a xor b;
    layer0_outputs(4748) <= a;
    layer0_outputs(4749) <= b;
    layer0_outputs(4750) <= '0';
    layer0_outputs(4751) <= a xor b;
    layer0_outputs(4752) <= not (a or b);
    layer0_outputs(4753) <= not (a or b);
    layer0_outputs(4754) <= a or b;
    layer0_outputs(4755) <= a;
    layer0_outputs(4756) <= not (a xor b);
    layer0_outputs(4757) <= not (a or b);
    layer0_outputs(4758) <= not a;
    layer0_outputs(4759) <= not (a xor b);
    layer0_outputs(4760) <= a xor b;
    layer0_outputs(4761) <= b;
    layer0_outputs(4762) <= a or b;
    layer0_outputs(4763) <= a or b;
    layer0_outputs(4764) <= not (a or b);
    layer0_outputs(4765) <= a or b;
    layer0_outputs(4766) <= not a;
    layer0_outputs(4767) <= not (a or b);
    layer0_outputs(4768) <= a or b;
    layer0_outputs(4769) <= a xor b;
    layer0_outputs(4770) <= a xor b;
    layer0_outputs(4771) <= not (a or b);
    layer0_outputs(4772) <= not a;
    layer0_outputs(4773) <= not a;
    layer0_outputs(4774) <= a or b;
    layer0_outputs(4775) <= b and not a;
    layer0_outputs(4776) <= not a or b;
    layer0_outputs(4777) <= a and not b;
    layer0_outputs(4778) <= a xor b;
    layer0_outputs(4779) <= a or b;
    layer0_outputs(4780) <= b;
    layer0_outputs(4781) <= not b or a;
    layer0_outputs(4782) <= not b or a;
    layer0_outputs(4783) <= a xor b;
    layer0_outputs(4784) <= not (a xor b);
    layer0_outputs(4785) <= not (a xor b);
    layer0_outputs(4786) <= not a;
    layer0_outputs(4787) <= not (a xor b);
    layer0_outputs(4788) <= a xor b;
    layer0_outputs(4789) <= a xor b;
    layer0_outputs(4790) <= not b or a;
    layer0_outputs(4791) <= a;
    layer0_outputs(4792) <= not b;
    layer0_outputs(4793) <= not (a or b);
    layer0_outputs(4794) <= a;
    layer0_outputs(4795) <= a xor b;
    layer0_outputs(4796) <= a or b;
    layer0_outputs(4797) <= not a or b;
    layer0_outputs(4798) <= not a;
    layer0_outputs(4799) <= a and not b;
    layer0_outputs(4800) <= a;
    layer0_outputs(4801) <= a or b;
    layer0_outputs(4802) <= a and not b;
    layer0_outputs(4803) <= not (a or b);
    layer0_outputs(4804) <= not (a xor b);
    layer0_outputs(4805) <= a or b;
    layer0_outputs(4806) <= '0';
    layer0_outputs(4807) <= b;
    layer0_outputs(4808) <= a xor b;
    layer0_outputs(4809) <= b;
    layer0_outputs(4810) <= b;
    layer0_outputs(4811) <= a and not b;
    layer0_outputs(4812) <= not a or b;
    layer0_outputs(4813) <= not b;
    layer0_outputs(4814) <= b;
    layer0_outputs(4815) <= b and not a;
    layer0_outputs(4816) <= b;
    layer0_outputs(4817) <= not (a xor b);
    layer0_outputs(4818) <= not a;
    layer0_outputs(4819) <= a and not b;
    layer0_outputs(4820) <= a and not b;
    layer0_outputs(4821) <= not b or a;
    layer0_outputs(4822) <= a and b;
    layer0_outputs(4823) <= a;
    layer0_outputs(4824) <= not (a or b);
    layer0_outputs(4825) <= not (a xor b);
    layer0_outputs(4826) <= b;
    layer0_outputs(4827) <= not a or b;
    layer0_outputs(4828) <= not (a xor b);
    layer0_outputs(4829) <= not a;
    layer0_outputs(4830) <= a or b;
    layer0_outputs(4831) <= not (a or b);
    layer0_outputs(4832) <= not (a or b);
    layer0_outputs(4833) <= a or b;
    layer0_outputs(4834) <= a or b;
    layer0_outputs(4835) <= not (a or b);
    layer0_outputs(4836) <= '1';
    layer0_outputs(4837) <= a xor b;
    layer0_outputs(4838) <= not b or a;
    layer0_outputs(4839) <= not a;
    layer0_outputs(4840) <= a;
    layer0_outputs(4841) <= not a;
    layer0_outputs(4842) <= a and not b;
    layer0_outputs(4843) <= not (a or b);
    layer0_outputs(4844) <= not a or b;
    layer0_outputs(4845) <= not (a xor b);
    layer0_outputs(4846) <= b and not a;
    layer0_outputs(4847) <= a xor b;
    layer0_outputs(4848) <= b;
    layer0_outputs(4849) <= a and not b;
    layer0_outputs(4850) <= a or b;
    layer0_outputs(4851) <= a and b;
    layer0_outputs(4852) <= not (a or b);
    layer0_outputs(4853) <= not b or a;
    layer0_outputs(4854) <= not (a or b);
    layer0_outputs(4855) <= a xor b;
    layer0_outputs(4856) <= b and not a;
    layer0_outputs(4857) <= not (a and b);
    layer0_outputs(4858) <= not a or b;
    layer0_outputs(4859) <= a xor b;
    layer0_outputs(4860) <= b;
    layer0_outputs(4861) <= not (a or b);
    layer0_outputs(4862) <= not (a and b);
    layer0_outputs(4863) <= not (a xor b);
    layer0_outputs(4864) <= not (a or b);
    layer0_outputs(4865) <= not b or a;
    layer0_outputs(4866) <= a xor b;
    layer0_outputs(4867) <= not b or a;
    layer0_outputs(4868) <= a or b;
    layer0_outputs(4869) <= '1';
    layer0_outputs(4870) <= a and not b;
    layer0_outputs(4871) <= not b;
    layer0_outputs(4872) <= a xor b;
    layer0_outputs(4873) <= b;
    layer0_outputs(4874) <= b and not a;
    layer0_outputs(4875) <= b and not a;
    layer0_outputs(4876) <= a or b;
    layer0_outputs(4877) <= a;
    layer0_outputs(4878) <= b and not a;
    layer0_outputs(4879) <= '1';
    layer0_outputs(4880) <= not (a or b);
    layer0_outputs(4881) <= '0';
    layer0_outputs(4882) <= b and not a;
    layer0_outputs(4883) <= a xor b;
    layer0_outputs(4884) <= a xor b;
    layer0_outputs(4885) <= a and not b;
    layer0_outputs(4886) <= a or b;
    layer0_outputs(4887) <= not b;
    layer0_outputs(4888) <= b;
    layer0_outputs(4889) <= not (a xor b);
    layer0_outputs(4890) <= not (a xor b);
    layer0_outputs(4891) <= not b;
    layer0_outputs(4892) <= a and not b;
    layer0_outputs(4893) <= not (a or b);
    layer0_outputs(4894) <= not (a or b);
    layer0_outputs(4895) <= not (a or b);
    layer0_outputs(4896) <= not (a or b);
    layer0_outputs(4897) <= a and not b;
    layer0_outputs(4898) <= a and not b;
    layer0_outputs(4899) <= a xor b;
    layer0_outputs(4900) <= not (a xor b);
    layer0_outputs(4901) <= not (a or b);
    layer0_outputs(4902) <= not (a or b);
    layer0_outputs(4903) <= not (a xor b);
    layer0_outputs(4904) <= b and not a;
    layer0_outputs(4905) <= a and b;
    layer0_outputs(4906) <= not b;
    layer0_outputs(4907) <= a xor b;
    layer0_outputs(4908) <= b and not a;
    layer0_outputs(4909) <= not (a xor b);
    layer0_outputs(4910) <= a xor b;
    layer0_outputs(4911) <= not b or a;
    layer0_outputs(4912) <= not (a or b);
    layer0_outputs(4913) <= a;
    layer0_outputs(4914) <= not (a or b);
    layer0_outputs(4915) <= not (a or b);
    layer0_outputs(4916) <= a or b;
    layer0_outputs(4917) <= not a;
    layer0_outputs(4918) <= a or b;
    layer0_outputs(4919) <= not (a or b);
    layer0_outputs(4920) <= not (a xor b);
    layer0_outputs(4921) <= not (a xor b);
    layer0_outputs(4922) <= a;
    layer0_outputs(4923) <= a and b;
    layer0_outputs(4924) <= not (a or b);
    layer0_outputs(4925) <= a;
    layer0_outputs(4926) <= not (a or b);
    layer0_outputs(4927) <= not (a xor b);
    layer0_outputs(4928) <= not b;
    layer0_outputs(4929) <= not b or a;
    layer0_outputs(4930) <= a;
    layer0_outputs(4931) <= b;
    layer0_outputs(4932) <= a xor b;
    layer0_outputs(4933) <= not (a or b);
    layer0_outputs(4934) <= a;
    layer0_outputs(4935) <= not a or b;
    layer0_outputs(4936) <= not b or a;
    layer0_outputs(4937) <= not (a or b);
    layer0_outputs(4938) <= not (a or b);
    layer0_outputs(4939) <= b and not a;
    layer0_outputs(4940) <= not (a xor b);
    layer0_outputs(4941) <= a or b;
    layer0_outputs(4942) <= a xor b;
    layer0_outputs(4943) <= a xor b;
    layer0_outputs(4944) <= not b;
    layer0_outputs(4945) <= a and not b;
    layer0_outputs(4946) <= not (a or b);
    layer0_outputs(4947) <= not (a xor b);
    layer0_outputs(4948) <= not a or b;
    layer0_outputs(4949) <= not (a or b);
    layer0_outputs(4950) <= b;
    layer0_outputs(4951) <= not a;
    layer0_outputs(4952) <= not (a xor b);
    layer0_outputs(4953) <= a;
    layer0_outputs(4954) <= a xor b;
    layer0_outputs(4955) <= not (a or b);
    layer0_outputs(4956) <= not b or a;
    layer0_outputs(4957) <= not (a or b);
    layer0_outputs(4958) <= a xor b;
    layer0_outputs(4959) <= not (a or b);
    layer0_outputs(4960) <= not (a or b);
    layer0_outputs(4961) <= b and not a;
    layer0_outputs(4962) <= a and not b;
    layer0_outputs(4963) <= not (a xor b);
    layer0_outputs(4964) <= not a;
    layer0_outputs(4965) <= not (a xor b);
    layer0_outputs(4966) <= a;
    layer0_outputs(4967) <= not a or b;
    layer0_outputs(4968) <= not b or a;
    layer0_outputs(4969) <= not (a xor b);
    layer0_outputs(4970) <= not b or a;
    layer0_outputs(4971) <= not b;
    layer0_outputs(4972) <= a or b;
    layer0_outputs(4973) <= a or b;
    layer0_outputs(4974) <= a xor b;
    layer0_outputs(4975) <= a and not b;
    layer0_outputs(4976) <= not b;
    layer0_outputs(4977) <= a and not b;
    layer0_outputs(4978) <= b;
    layer0_outputs(4979) <= not b or a;
    layer0_outputs(4980) <= not b or a;
    layer0_outputs(4981) <= a xor b;
    layer0_outputs(4982) <= b and not a;
    layer0_outputs(4983) <= not a or b;
    layer0_outputs(4984) <= '1';
    layer0_outputs(4985) <= not a or b;
    layer0_outputs(4986) <= a and not b;
    layer0_outputs(4987) <= '1';
    layer0_outputs(4988) <= a xor b;
    layer0_outputs(4989) <= not b;
    layer0_outputs(4990) <= b and not a;
    layer0_outputs(4991) <= a xor b;
    layer0_outputs(4992) <= a and not b;
    layer0_outputs(4993) <= not (a or b);
    layer0_outputs(4994) <= not a or b;
    layer0_outputs(4995) <= '1';
    layer0_outputs(4996) <= a and not b;
    layer0_outputs(4997) <= not (a or b);
    layer0_outputs(4998) <= a or b;
    layer0_outputs(4999) <= not (a xor b);
    layer0_outputs(5000) <= not b or a;
    layer0_outputs(5001) <= a or b;
    layer0_outputs(5002) <= b;
    layer0_outputs(5003) <= not b;
    layer0_outputs(5004) <= not (a or b);
    layer0_outputs(5005) <= not b;
    layer0_outputs(5006) <= b;
    layer0_outputs(5007) <= a and b;
    layer0_outputs(5008) <= not a;
    layer0_outputs(5009) <= a xor b;
    layer0_outputs(5010) <= not (a or b);
    layer0_outputs(5011) <= not b or a;
    layer0_outputs(5012) <= not (a or b);
    layer0_outputs(5013) <= not b or a;
    layer0_outputs(5014) <= a or b;
    layer0_outputs(5015) <= a xor b;
    layer0_outputs(5016) <= a xor b;
    layer0_outputs(5017) <= a xor b;
    layer0_outputs(5018) <= not (a or b);
    layer0_outputs(5019) <= not b or a;
    layer0_outputs(5020) <= a and not b;
    layer0_outputs(5021) <= a xor b;
    layer0_outputs(5022) <= a or b;
    layer0_outputs(5023) <= a;
    layer0_outputs(5024) <= a and not b;
    layer0_outputs(5025) <= not (a xor b);
    layer0_outputs(5026) <= not (a or b);
    layer0_outputs(5027) <= not (a and b);
    layer0_outputs(5028) <= not b;
    layer0_outputs(5029) <= a;
    layer0_outputs(5030) <= not a;
    layer0_outputs(5031) <= not (a xor b);
    layer0_outputs(5032) <= a;
    layer0_outputs(5033) <= b;
    layer0_outputs(5034) <= not (a or b);
    layer0_outputs(5035) <= a;
    layer0_outputs(5036) <= b;
    layer0_outputs(5037) <= not (a or b);
    layer0_outputs(5038) <= not b;
    layer0_outputs(5039) <= a and not b;
    layer0_outputs(5040) <= not (a or b);
    layer0_outputs(5041) <= not b or a;
    layer0_outputs(5042) <= b;
    layer0_outputs(5043) <= a and b;
    layer0_outputs(5044) <= not (a xor b);
    layer0_outputs(5045) <= a xor b;
    layer0_outputs(5046) <= a and not b;
    layer0_outputs(5047) <= b and not a;
    layer0_outputs(5048) <= not (a xor b);
    layer0_outputs(5049) <= not (a and b);
    layer0_outputs(5050) <= not (a or b);
    layer0_outputs(5051) <= not (a xor b);
    layer0_outputs(5052) <= not b;
    layer0_outputs(5053) <= not b or a;
    layer0_outputs(5054) <= '1';
    layer0_outputs(5055) <= not (a or b);
    layer0_outputs(5056) <= a and b;
    layer0_outputs(5057) <= not (a or b);
    layer0_outputs(5058) <= not (a or b);
    layer0_outputs(5059) <= a xor b;
    layer0_outputs(5060) <= a xor b;
    layer0_outputs(5061) <= a;
    layer0_outputs(5062) <= not (a and b);
    layer0_outputs(5063) <= not a;
    layer0_outputs(5064) <= not a or b;
    layer0_outputs(5065) <= not (a or b);
    layer0_outputs(5066) <= a xor b;
    layer0_outputs(5067) <= not a;
    layer0_outputs(5068) <= not (a or b);
    layer0_outputs(5069) <= a;
    layer0_outputs(5070) <= b;
    layer0_outputs(5071) <= a;
    layer0_outputs(5072) <= not a;
    layer0_outputs(5073) <= not a;
    layer0_outputs(5074) <= a xor b;
    layer0_outputs(5075) <= not (a xor b);
    layer0_outputs(5076) <= a and not b;
    layer0_outputs(5077) <= not (a xor b);
    layer0_outputs(5078) <= a xor b;
    layer0_outputs(5079) <= a;
    layer0_outputs(5080) <= not a;
    layer0_outputs(5081) <= a or b;
    layer0_outputs(5082) <= b;
    layer0_outputs(5083) <= not (a or b);
    layer0_outputs(5084) <= b and not a;
    layer0_outputs(5085) <= not (a xor b);
    layer0_outputs(5086) <= a or b;
    layer0_outputs(5087) <= not b;
    layer0_outputs(5088) <= a or b;
    layer0_outputs(5089) <= not b or a;
    layer0_outputs(5090) <= a xor b;
    layer0_outputs(5091) <= not a or b;
    layer0_outputs(5092) <= a or b;
    layer0_outputs(5093) <= a and not b;
    layer0_outputs(5094) <= not b or a;
    layer0_outputs(5095) <= a xor b;
    layer0_outputs(5096) <= not a or b;
    layer0_outputs(5097) <= a;
    layer0_outputs(5098) <= b and not a;
    layer0_outputs(5099) <= not a or b;
    layer0_outputs(5100) <= a or b;
    layer0_outputs(5101) <= '1';
    layer0_outputs(5102) <= a xor b;
    layer0_outputs(5103) <= a or b;
    layer0_outputs(5104) <= a xor b;
    layer0_outputs(5105) <= a xor b;
    layer0_outputs(5106) <= a and not b;
    layer0_outputs(5107) <= a xor b;
    layer0_outputs(5108) <= not (a or b);
    layer0_outputs(5109) <= not a or b;
    layer0_outputs(5110) <= not a or b;
    layer0_outputs(5111) <= '1';
    layer0_outputs(5112) <= a xor b;
    layer0_outputs(5113) <= a or b;
    layer0_outputs(5114) <= a;
    layer0_outputs(5115) <= not a;
    layer0_outputs(5116) <= not b;
    layer0_outputs(5117) <= a;
    layer0_outputs(5118) <= a or b;
    layer0_outputs(5119) <= not b or a;
    layer0_outputs(5120) <= a and b;
    layer0_outputs(5121) <= a;
    layer0_outputs(5122) <= a or b;
    layer0_outputs(5123) <= a or b;
    layer0_outputs(5124) <= not (a or b);
    layer0_outputs(5125) <= not b or a;
    layer0_outputs(5126) <= not a;
    layer0_outputs(5127) <= a and b;
    layer0_outputs(5128) <= not (a xor b);
    layer0_outputs(5129) <= not a;
    layer0_outputs(5130) <= b;
    layer0_outputs(5131) <= b and not a;
    layer0_outputs(5132) <= not (a xor b);
    layer0_outputs(5133) <= a;
    layer0_outputs(5134) <= '0';
    layer0_outputs(5135) <= not a or b;
    layer0_outputs(5136) <= not b or a;
    layer0_outputs(5137) <= a xor b;
    layer0_outputs(5138) <= not (a or b);
    layer0_outputs(5139) <= b and not a;
    layer0_outputs(5140) <= not b;
    layer0_outputs(5141) <= a xor b;
    layer0_outputs(5142) <= not b or a;
    layer0_outputs(5143) <= not b or a;
    layer0_outputs(5144) <= '1';
    layer0_outputs(5145) <= not b;
    layer0_outputs(5146) <= not (a xor b);
    layer0_outputs(5147) <= not (a xor b);
    layer0_outputs(5148) <= a or b;
    layer0_outputs(5149) <= b and not a;
    layer0_outputs(5150) <= a or b;
    layer0_outputs(5151) <= a or b;
    layer0_outputs(5152) <= not b;
    layer0_outputs(5153) <= not (a xor b);
    layer0_outputs(5154) <= a or b;
    layer0_outputs(5155) <= not b;
    layer0_outputs(5156) <= not (a or b);
    layer0_outputs(5157) <= not a or b;
    layer0_outputs(5158) <= a;
    layer0_outputs(5159) <= b and not a;
    layer0_outputs(5160) <= not (a or b);
    layer0_outputs(5161) <= b and not a;
    layer0_outputs(5162) <= not (a and b);
    layer0_outputs(5163) <= a;
    layer0_outputs(5164) <= not (a or b);
    layer0_outputs(5165) <= not b;
    layer0_outputs(5166) <= a or b;
    layer0_outputs(5167) <= a or b;
    layer0_outputs(5168) <= a xor b;
    layer0_outputs(5169) <= b;
    layer0_outputs(5170) <= a or b;
    layer0_outputs(5171) <= not a or b;
    layer0_outputs(5172) <= a or b;
    layer0_outputs(5173) <= b;
    layer0_outputs(5174) <= not a;
    layer0_outputs(5175) <= b and not a;
    layer0_outputs(5176) <= not b;
    layer0_outputs(5177) <= a or b;
    layer0_outputs(5178) <= not (a or b);
    layer0_outputs(5179) <= b;
    layer0_outputs(5180) <= not (a xor b);
    layer0_outputs(5181) <= not (a or b);
    layer0_outputs(5182) <= b and not a;
    layer0_outputs(5183) <= a xor b;
    layer0_outputs(5184) <= a and not b;
    layer0_outputs(5185) <= a;
    layer0_outputs(5186) <= a and not b;
    layer0_outputs(5187) <= not b or a;
    layer0_outputs(5188) <= b;
    layer0_outputs(5189) <= a or b;
    layer0_outputs(5190) <= b and not a;
    layer0_outputs(5191) <= '1';
    layer0_outputs(5192) <= '1';
    layer0_outputs(5193) <= a or b;
    layer0_outputs(5194) <= not (a or b);
    layer0_outputs(5195) <= not (a or b);
    layer0_outputs(5196) <= b and not a;
    layer0_outputs(5197) <= a and b;
    layer0_outputs(5198) <= a;
    layer0_outputs(5199) <= a;
    layer0_outputs(5200) <= b;
    layer0_outputs(5201) <= not (a xor b);
    layer0_outputs(5202) <= b;
    layer0_outputs(5203) <= a or b;
    layer0_outputs(5204) <= a or b;
    layer0_outputs(5205) <= not b;
    layer0_outputs(5206) <= a or b;
    layer0_outputs(5207) <= not a;
    layer0_outputs(5208) <= '1';
    layer0_outputs(5209) <= not b or a;
    layer0_outputs(5210) <= not a;
    layer0_outputs(5211) <= a or b;
    layer0_outputs(5212) <= not (a or b);
    layer0_outputs(5213) <= not a or b;
    layer0_outputs(5214) <= not b or a;
    layer0_outputs(5215) <= a or b;
    layer0_outputs(5216) <= not (a or b);
    layer0_outputs(5217) <= a and not b;
    layer0_outputs(5218) <= not b;
    layer0_outputs(5219) <= not (a or b);
    layer0_outputs(5220) <= a xor b;
    layer0_outputs(5221) <= a or b;
    layer0_outputs(5222) <= a and b;
    layer0_outputs(5223) <= a or b;
    layer0_outputs(5224) <= a xor b;
    layer0_outputs(5225) <= a and not b;
    layer0_outputs(5226) <= not b;
    layer0_outputs(5227) <= not (a xor b);
    layer0_outputs(5228) <= not (a xor b);
    layer0_outputs(5229) <= a;
    layer0_outputs(5230) <= not a;
    layer0_outputs(5231) <= not (a or b);
    layer0_outputs(5232) <= not (a or b);
    layer0_outputs(5233) <= not a or b;
    layer0_outputs(5234) <= not a;
    layer0_outputs(5235) <= a;
    layer0_outputs(5236) <= not a or b;
    layer0_outputs(5237) <= not (a xor b);
    layer0_outputs(5238) <= not b or a;
    layer0_outputs(5239) <= b and not a;
    layer0_outputs(5240) <= a or b;
    layer0_outputs(5241) <= a and b;
    layer0_outputs(5242) <= not (a or b);
    layer0_outputs(5243) <= b;
    layer0_outputs(5244) <= not (a or b);
    layer0_outputs(5245) <= a and b;
    layer0_outputs(5246) <= '1';
    layer0_outputs(5247) <= not b or a;
    layer0_outputs(5248) <= a or b;
    layer0_outputs(5249) <= a;
    layer0_outputs(5250) <= b;
    layer0_outputs(5251) <= not b or a;
    layer0_outputs(5252) <= not a;
    layer0_outputs(5253) <= a xor b;
    layer0_outputs(5254) <= b;
    layer0_outputs(5255) <= a or b;
    layer0_outputs(5256) <= a xor b;
    layer0_outputs(5257) <= not a;
    layer0_outputs(5258) <= a xor b;
    layer0_outputs(5259) <= not (a or b);
    layer0_outputs(5260) <= a or b;
    layer0_outputs(5261) <= not (a xor b);
    layer0_outputs(5262) <= b;
    layer0_outputs(5263) <= not (a or b);
    layer0_outputs(5264) <= a xor b;
    layer0_outputs(5265) <= not b or a;
    layer0_outputs(5266) <= not b;
    layer0_outputs(5267) <= not a or b;
    layer0_outputs(5268) <= a xor b;
    layer0_outputs(5269) <= a xor b;
    layer0_outputs(5270) <= b;
    layer0_outputs(5271) <= not (a or b);
    layer0_outputs(5272) <= b;
    layer0_outputs(5273) <= a;
    layer0_outputs(5274) <= not (a xor b);
    layer0_outputs(5275) <= a;
    layer0_outputs(5276) <= not a;
    layer0_outputs(5277) <= a or b;
    layer0_outputs(5278) <= not (a xor b);
    layer0_outputs(5279) <= not b or a;
    layer0_outputs(5280) <= not b or a;
    layer0_outputs(5281) <= a;
    layer0_outputs(5282) <= a or b;
    layer0_outputs(5283) <= a xor b;
    layer0_outputs(5284) <= a or b;
    layer0_outputs(5285) <= a or b;
    layer0_outputs(5286) <= not b or a;
    layer0_outputs(5287) <= b and not a;
    layer0_outputs(5288) <= not a;
    layer0_outputs(5289) <= a;
    layer0_outputs(5290) <= a and not b;
    layer0_outputs(5291) <= b and not a;
    layer0_outputs(5292) <= b;
    layer0_outputs(5293) <= a or b;
    layer0_outputs(5294) <= a xor b;
    layer0_outputs(5295) <= not (a xor b);
    layer0_outputs(5296) <= not (a xor b);
    layer0_outputs(5297) <= a and not b;
    layer0_outputs(5298) <= not a or b;
    layer0_outputs(5299) <= a xor b;
    layer0_outputs(5300) <= not a;
    layer0_outputs(5301) <= a and not b;
    layer0_outputs(5302) <= a;
    layer0_outputs(5303) <= not a or b;
    layer0_outputs(5304) <= a;
    layer0_outputs(5305) <= not a or b;
    layer0_outputs(5306) <= '1';
    layer0_outputs(5307) <= not b;
    layer0_outputs(5308) <= a or b;
    layer0_outputs(5309) <= not b;
    layer0_outputs(5310) <= a or b;
    layer0_outputs(5311) <= a xor b;
    layer0_outputs(5312) <= not (a xor b);
    layer0_outputs(5313) <= '1';
    layer0_outputs(5314) <= a xor b;
    layer0_outputs(5315) <= not a or b;
    layer0_outputs(5316) <= not (a or b);
    layer0_outputs(5317) <= not (a or b);
    layer0_outputs(5318) <= a and not b;
    layer0_outputs(5319) <= a xor b;
    layer0_outputs(5320) <= a and not b;
    layer0_outputs(5321) <= b;
    layer0_outputs(5322) <= a or b;
    layer0_outputs(5323) <= not b;
    layer0_outputs(5324) <= not (a and b);
    layer0_outputs(5325) <= not b or a;
    layer0_outputs(5326) <= not (a or b);
    layer0_outputs(5327) <= not b or a;
    layer0_outputs(5328) <= not (a or b);
    layer0_outputs(5329) <= a and not b;
    layer0_outputs(5330) <= a xor b;
    layer0_outputs(5331) <= not (a and b);
    layer0_outputs(5332) <= not (a or b);
    layer0_outputs(5333) <= not (a or b);
    layer0_outputs(5334) <= not a;
    layer0_outputs(5335) <= not b or a;
    layer0_outputs(5336) <= not a;
    layer0_outputs(5337) <= b;
    layer0_outputs(5338) <= b;
    layer0_outputs(5339) <= a xor b;
    layer0_outputs(5340) <= not (a xor b);
    layer0_outputs(5341) <= b and not a;
    layer0_outputs(5342) <= b and not a;
    layer0_outputs(5343) <= not b;
    layer0_outputs(5344) <= not b or a;
    layer0_outputs(5345) <= not b;
    layer0_outputs(5346) <= not (a xor b);
    layer0_outputs(5347) <= '0';
    layer0_outputs(5348) <= a or b;
    layer0_outputs(5349) <= not (a xor b);
    layer0_outputs(5350) <= not (a xor b);
    layer0_outputs(5351) <= not (a xor b);
    layer0_outputs(5352) <= a xor b;
    layer0_outputs(5353) <= not a or b;
    layer0_outputs(5354) <= a or b;
    layer0_outputs(5355) <= b;
    layer0_outputs(5356) <= not a or b;
    layer0_outputs(5357) <= not (a xor b);
    layer0_outputs(5358) <= b and not a;
    layer0_outputs(5359) <= a or b;
    layer0_outputs(5360) <= a xor b;
    layer0_outputs(5361) <= a;
    layer0_outputs(5362) <= a or b;
    layer0_outputs(5363) <= not b;
    layer0_outputs(5364) <= a or b;
    layer0_outputs(5365) <= '1';
    layer0_outputs(5366) <= b and not a;
    layer0_outputs(5367) <= not a;
    layer0_outputs(5368) <= a;
    layer0_outputs(5369) <= b;
    layer0_outputs(5370) <= b;
    layer0_outputs(5371) <= not (a or b);
    layer0_outputs(5372) <= not (a xor b);
    layer0_outputs(5373) <= a;
    layer0_outputs(5374) <= not a or b;
    layer0_outputs(5375) <= a or b;
    layer0_outputs(5376) <= not a or b;
    layer0_outputs(5377) <= a or b;
    layer0_outputs(5378) <= not (a xor b);
    layer0_outputs(5379) <= not (a or b);
    layer0_outputs(5380) <= a and not b;
    layer0_outputs(5381) <= not (a xor b);
    layer0_outputs(5382) <= not (a or b);
    layer0_outputs(5383) <= '1';
    layer0_outputs(5384) <= not (a xor b);
    layer0_outputs(5385) <= a or b;
    layer0_outputs(5386) <= not (a or b);
    layer0_outputs(5387) <= not (a or b);
    layer0_outputs(5388) <= a or b;
    layer0_outputs(5389) <= b;
    layer0_outputs(5390) <= b;
    layer0_outputs(5391) <= not (a or b);
    layer0_outputs(5392) <= not (a and b);
    layer0_outputs(5393) <= a or b;
    layer0_outputs(5394) <= not a or b;
    layer0_outputs(5395) <= not a;
    layer0_outputs(5396) <= a;
    layer0_outputs(5397) <= b and not a;
    layer0_outputs(5398) <= not (a or b);
    layer0_outputs(5399) <= not a or b;
    layer0_outputs(5400) <= not a or b;
    layer0_outputs(5401) <= a and not b;
    layer0_outputs(5402) <= a;
    layer0_outputs(5403) <= not (a xor b);
    layer0_outputs(5404) <= not (a or b);
    layer0_outputs(5405) <= not (a xor b);
    layer0_outputs(5406) <= not b;
    layer0_outputs(5407) <= a;
    layer0_outputs(5408) <= a or b;
    layer0_outputs(5409) <= a and not b;
    layer0_outputs(5410) <= b;
    layer0_outputs(5411) <= a or b;
    layer0_outputs(5412) <= not a;
    layer0_outputs(5413) <= b;
    layer0_outputs(5414) <= '0';
    layer0_outputs(5415) <= a and not b;
    layer0_outputs(5416) <= not (a or b);
    layer0_outputs(5417) <= not b or a;
    layer0_outputs(5418) <= not (a xor b);
    layer0_outputs(5419) <= not a or b;
    layer0_outputs(5420) <= b;
    layer0_outputs(5421) <= not a or b;
    layer0_outputs(5422) <= not (a or b);
    layer0_outputs(5423) <= b and not a;
    layer0_outputs(5424) <= not (a or b);
    layer0_outputs(5425) <= b and not a;
    layer0_outputs(5426) <= a and b;
    layer0_outputs(5427) <= not a or b;
    layer0_outputs(5428) <= b and not a;
    layer0_outputs(5429) <= b;
    layer0_outputs(5430) <= not (a xor b);
    layer0_outputs(5431) <= a and b;
    layer0_outputs(5432) <= not (a xor b);
    layer0_outputs(5433) <= not a;
    layer0_outputs(5434) <= not a or b;
    layer0_outputs(5435) <= not (a xor b);
    layer0_outputs(5436) <= a or b;
    layer0_outputs(5437) <= not a;
    layer0_outputs(5438) <= a;
    layer0_outputs(5439) <= a;
    layer0_outputs(5440) <= not a or b;
    layer0_outputs(5441) <= a;
    layer0_outputs(5442) <= not b;
    layer0_outputs(5443) <= a or b;
    layer0_outputs(5444) <= '1';
    layer0_outputs(5445) <= not (a or b);
    layer0_outputs(5446) <= not a;
    layer0_outputs(5447) <= not a or b;
    layer0_outputs(5448) <= not a or b;
    layer0_outputs(5449) <= not (a or b);
    layer0_outputs(5450) <= a;
    layer0_outputs(5451) <= not (a or b);
    layer0_outputs(5452) <= not (a or b);
    layer0_outputs(5453) <= a or b;
    layer0_outputs(5454) <= a xor b;
    layer0_outputs(5455) <= not (a or b);
    layer0_outputs(5456) <= not (a xor b);
    layer0_outputs(5457) <= a;
    layer0_outputs(5458) <= a or b;
    layer0_outputs(5459) <= a xor b;
    layer0_outputs(5460) <= not (a or b);
    layer0_outputs(5461) <= not (a and b);
    layer0_outputs(5462) <= a or b;
    layer0_outputs(5463) <= a and not b;
    layer0_outputs(5464) <= a;
    layer0_outputs(5465) <= not (a or b);
    layer0_outputs(5466) <= not (a xor b);
    layer0_outputs(5467) <= a xor b;
    layer0_outputs(5468) <= a or b;
    layer0_outputs(5469) <= a or b;
    layer0_outputs(5470) <= not a;
    layer0_outputs(5471) <= a or b;
    layer0_outputs(5472) <= not a;
    layer0_outputs(5473) <= not b;
    layer0_outputs(5474) <= not a or b;
    layer0_outputs(5475) <= not b;
    layer0_outputs(5476) <= not (a or b);
    layer0_outputs(5477) <= b and not a;
    layer0_outputs(5478) <= '1';
    layer0_outputs(5479) <= not (a or b);
    layer0_outputs(5480) <= not b;
    layer0_outputs(5481) <= b and not a;
    layer0_outputs(5482) <= a and not b;
    layer0_outputs(5483) <= not b;
    layer0_outputs(5484) <= b and not a;
    layer0_outputs(5485) <= not b or a;
    layer0_outputs(5486) <= b and not a;
    layer0_outputs(5487) <= not (a xor b);
    layer0_outputs(5488) <= a or b;
    layer0_outputs(5489) <= not (a xor b);
    layer0_outputs(5490) <= a and not b;
    layer0_outputs(5491) <= not (a xor b);
    layer0_outputs(5492) <= a xor b;
    layer0_outputs(5493) <= a or b;
    layer0_outputs(5494) <= a or b;
    layer0_outputs(5495) <= not (a xor b);
    layer0_outputs(5496) <= a;
    layer0_outputs(5497) <= a;
    layer0_outputs(5498) <= a or b;
    layer0_outputs(5499) <= not b;
    layer0_outputs(5500) <= not (a or b);
    layer0_outputs(5501) <= b;
    layer0_outputs(5502) <= not (a or b);
    layer0_outputs(5503) <= b;
    layer0_outputs(5504) <= a;
    layer0_outputs(5505) <= '0';
    layer0_outputs(5506) <= a;
    layer0_outputs(5507) <= a or b;
    layer0_outputs(5508) <= a xor b;
    layer0_outputs(5509) <= not (a or b);
    layer0_outputs(5510) <= a or b;
    layer0_outputs(5511) <= '1';
    layer0_outputs(5512) <= not (a xor b);
    layer0_outputs(5513) <= b;
    layer0_outputs(5514) <= not a;
    layer0_outputs(5515) <= a or b;
    layer0_outputs(5516) <= not (a or b);
    layer0_outputs(5517) <= a xor b;
    layer0_outputs(5518) <= not b or a;
    layer0_outputs(5519) <= a or b;
    layer0_outputs(5520) <= not (a or b);
    layer0_outputs(5521) <= a xor b;
    layer0_outputs(5522) <= not a;
    layer0_outputs(5523) <= not (a or b);
    layer0_outputs(5524) <= not (a or b);
    layer0_outputs(5525) <= a or b;
    layer0_outputs(5526) <= a xor b;
    layer0_outputs(5527) <= not (a and b);
    layer0_outputs(5528) <= b;
    layer0_outputs(5529) <= a;
    layer0_outputs(5530) <= not (a xor b);
    layer0_outputs(5531) <= not b or a;
    layer0_outputs(5532) <= not b;
    layer0_outputs(5533) <= a and b;
    layer0_outputs(5534) <= a or b;
    layer0_outputs(5535) <= not b;
    layer0_outputs(5536) <= b;
    layer0_outputs(5537) <= a or b;
    layer0_outputs(5538) <= a and not b;
    layer0_outputs(5539) <= a or b;
    layer0_outputs(5540) <= not b or a;
    layer0_outputs(5541) <= not (a xor b);
    layer0_outputs(5542) <= a xor b;
    layer0_outputs(5543) <= a xor b;
    layer0_outputs(5544) <= a;
    layer0_outputs(5545) <= a xor b;
    layer0_outputs(5546) <= not a or b;
    layer0_outputs(5547) <= not (a or b);
    layer0_outputs(5548) <= a or b;
    layer0_outputs(5549) <= not (a or b);
    layer0_outputs(5550) <= not b or a;
    layer0_outputs(5551) <= b;
    layer0_outputs(5552) <= not (a or b);
    layer0_outputs(5553) <= not (a xor b);
    layer0_outputs(5554) <= a or b;
    layer0_outputs(5555) <= not b;
    layer0_outputs(5556) <= a and b;
    layer0_outputs(5557) <= a or b;
    layer0_outputs(5558) <= a or b;
    layer0_outputs(5559) <= not a;
    layer0_outputs(5560) <= a or b;
    layer0_outputs(5561) <= a or b;
    layer0_outputs(5562) <= not a;
    layer0_outputs(5563) <= a or b;
    layer0_outputs(5564) <= a or b;
    layer0_outputs(5565) <= not (a or b);
    layer0_outputs(5566) <= not a;
    layer0_outputs(5567) <= not (a xor b);
    layer0_outputs(5568) <= a;
    layer0_outputs(5569) <= not (a or b);
    layer0_outputs(5570) <= a or b;
    layer0_outputs(5571) <= not b or a;
    layer0_outputs(5572) <= not b;
    layer0_outputs(5573) <= a or b;
    layer0_outputs(5574) <= b and not a;
    layer0_outputs(5575) <= b and not a;
    layer0_outputs(5576) <= a xor b;
    layer0_outputs(5577) <= a or b;
    layer0_outputs(5578) <= not b;
    layer0_outputs(5579) <= not (a xor b);
    layer0_outputs(5580) <= a and not b;
    layer0_outputs(5581) <= a and not b;
    layer0_outputs(5582) <= not (a xor b);
    layer0_outputs(5583) <= not (a xor b);
    layer0_outputs(5584) <= not b or a;
    layer0_outputs(5585) <= not b or a;
    layer0_outputs(5586) <= '1';
    layer0_outputs(5587) <= a or b;
    layer0_outputs(5588) <= not (a xor b);
    layer0_outputs(5589) <= not a or b;
    layer0_outputs(5590) <= not (a xor b);
    layer0_outputs(5591) <= not a or b;
    layer0_outputs(5592) <= a and b;
    layer0_outputs(5593) <= a xor b;
    layer0_outputs(5594) <= '0';
    layer0_outputs(5595) <= '0';
    layer0_outputs(5596) <= not a or b;
    layer0_outputs(5597) <= b and not a;
    layer0_outputs(5598) <= not (a xor b);
    layer0_outputs(5599) <= not (a xor b);
    layer0_outputs(5600) <= a and not b;
    layer0_outputs(5601) <= a or b;
    layer0_outputs(5602) <= a xor b;
    layer0_outputs(5603) <= not b or a;
    layer0_outputs(5604) <= b;
    layer0_outputs(5605) <= not (a or b);
    layer0_outputs(5606) <= a and b;
    layer0_outputs(5607) <= a or b;
    layer0_outputs(5608) <= a and not b;
    layer0_outputs(5609) <= not (a xor b);
    layer0_outputs(5610) <= a or b;
    layer0_outputs(5611) <= not b or a;
    layer0_outputs(5612) <= a xor b;
    layer0_outputs(5613) <= b and not a;
    layer0_outputs(5614) <= not b or a;
    layer0_outputs(5615) <= a and not b;
    layer0_outputs(5616) <= not (a or b);
    layer0_outputs(5617) <= a or b;
    layer0_outputs(5618) <= not (a or b);
    layer0_outputs(5619) <= b;
    layer0_outputs(5620) <= a and not b;
    layer0_outputs(5621) <= a or b;
    layer0_outputs(5622) <= not b or a;
    layer0_outputs(5623) <= a or b;
    layer0_outputs(5624) <= a or b;
    layer0_outputs(5625) <= a xor b;
    layer0_outputs(5626) <= a xor b;
    layer0_outputs(5627) <= a;
    layer0_outputs(5628) <= not b;
    layer0_outputs(5629) <= not (a or b);
    layer0_outputs(5630) <= not a;
    layer0_outputs(5631) <= not (a xor b);
    layer0_outputs(5632) <= not (a xor b);
    layer0_outputs(5633) <= not (a xor b);
    layer0_outputs(5634) <= a xor b;
    layer0_outputs(5635) <= b;
    layer0_outputs(5636) <= b;
    layer0_outputs(5637) <= a xor b;
    layer0_outputs(5638) <= not (a or b);
    layer0_outputs(5639) <= not a;
    layer0_outputs(5640) <= a and not b;
    layer0_outputs(5641) <= b;
    layer0_outputs(5642) <= not (a or b);
    layer0_outputs(5643) <= a or b;
    layer0_outputs(5644) <= not a;
    layer0_outputs(5645) <= a;
    layer0_outputs(5646) <= not (a xor b);
    layer0_outputs(5647) <= not (a and b);
    layer0_outputs(5648) <= not a or b;
    layer0_outputs(5649) <= not (a or b);
    layer0_outputs(5650) <= b and not a;
    layer0_outputs(5651) <= not a or b;
    layer0_outputs(5652) <= b;
    layer0_outputs(5653) <= b;
    layer0_outputs(5654) <= not (a or b);
    layer0_outputs(5655) <= not a;
    layer0_outputs(5656) <= a;
    layer0_outputs(5657) <= a xor b;
    layer0_outputs(5658) <= not (a xor b);
    layer0_outputs(5659) <= not (a or b);
    layer0_outputs(5660) <= b and not a;
    layer0_outputs(5661) <= not (a and b);
    layer0_outputs(5662) <= b;
    layer0_outputs(5663) <= a;
    layer0_outputs(5664) <= not (a xor b);
    layer0_outputs(5665) <= b and not a;
    layer0_outputs(5666) <= a or b;
    layer0_outputs(5667) <= not a or b;
    layer0_outputs(5668) <= not (a or b);
    layer0_outputs(5669) <= not a or b;
    layer0_outputs(5670) <= b and not a;
    layer0_outputs(5671) <= not (a or b);
    layer0_outputs(5672) <= a or b;
    layer0_outputs(5673) <= not (a xor b);
    layer0_outputs(5674) <= a or b;
    layer0_outputs(5675) <= not (a and b);
    layer0_outputs(5676) <= a or b;
    layer0_outputs(5677) <= not b;
    layer0_outputs(5678) <= not (a or b);
    layer0_outputs(5679) <= '1';
    layer0_outputs(5680) <= a and not b;
    layer0_outputs(5681) <= not (a and b);
    layer0_outputs(5682) <= not b;
    layer0_outputs(5683) <= not (a or b);
    layer0_outputs(5684) <= b and not a;
    layer0_outputs(5685) <= b and not a;
    layer0_outputs(5686) <= not (a xor b);
    layer0_outputs(5687) <= '1';
    layer0_outputs(5688) <= not a;
    layer0_outputs(5689) <= '1';
    layer0_outputs(5690) <= a and not b;
    layer0_outputs(5691) <= a xor b;
    layer0_outputs(5692) <= b and not a;
    layer0_outputs(5693) <= a xor b;
    layer0_outputs(5694) <= not b;
    layer0_outputs(5695) <= b;
    layer0_outputs(5696) <= b;
    layer0_outputs(5697) <= a and not b;
    layer0_outputs(5698) <= b;
    layer0_outputs(5699) <= b;
    layer0_outputs(5700) <= a or b;
    layer0_outputs(5701) <= a;
    layer0_outputs(5702) <= b;
    layer0_outputs(5703) <= '0';
    layer0_outputs(5704) <= b and not a;
    layer0_outputs(5705) <= not (a or b);
    layer0_outputs(5706) <= a and not b;
    layer0_outputs(5707) <= a and not b;
    layer0_outputs(5708) <= not (a or b);
    layer0_outputs(5709) <= not (a xor b);
    layer0_outputs(5710) <= not b;
    layer0_outputs(5711) <= not a or b;
    layer0_outputs(5712) <= b;
    layer0_outputs(5713) <= a xor b;
    layer0_outputs(5714) <= b and not a;
    layer0_outputs(5715) <= b;
    layer0_outputs(5716) <= not b;
    layer0_outputs(5717) <= not (a xor b);
    layer0_outputs(5718) <= not (a or b);
    layer0_outputs(5719) <= not b;
    layer0_outputs(5720) <= '0';
    layer0_outputs(5721) <= not (a or b);
    layer0_outputs(5722) <= not a;
    layer0_outputs(5723) <= a or b;
    layer0_outputs(5724) <= a and b;
    layer0_outputs(5725) <= a;
    layer0_outputs(5726) <= b;
    layer0_outputs(5727) <= a;
    layer0_outputs(5728) <= a;
    layer0_outputs(5729) <= b and not a;
    layer0_outputs(5730) <= not (a or b);
    layer0_outputs(5731) <= b;
    layer0_outputs(5732) <= a and not b;
    layer0_outputs(5733) <= not (a and b);
    layer0_outputs(5734) <= a xor b;
    layer0_outputs(5735) <= not b or a;
    layer0_outputs(5736) <= not (a or b);
    layer0_outputs(5737) <= a or b;
    layer0_outputs(5738) <= a and not b;
    layer0_outputs(5739) <= a and b;
    layer0_outputs(5740) <= not (a or b);
    layer0_outputs(5741) <= not a or b;
    layer0_outputs(5742) <= b and not a;
    layer0_outputs(5743) <= b and not a;
    layer0_outputs(5744) <= not (a xor b);
    layer0_outputs(5745) <= not (a xor b);
    layer0_outputs(5746) <= b and not a;
    layer0_outputs(5747) <= not (a and b);
    layer0_outputs(5748) <= a or b;
    layer0_outputs(5749) <= a or b;
    layer0_outputs(5750) <= a or b;
    layer0_outputs(5751) <= not a or b;
    layer0_outputs(5752) <= not (a and b);
    layer0_outputs(5753) <= a;
    layer0_outputs(5754) <= a;
    layer0_outputs(5755) <= not b or a;
    layer0_outputs(5756) <= not b or a;
    layer0_outputs(5757) <= not (a xor b);
    layer0_outputs(5758) <= not a;
    layer0_outputs(5759) <= a or b;
    layer0_outputs(5760) <= not b;
    layer0_outputs(5761) <= a or b;
    layer0_outputs(5762) <= b;
    layer0_outputs(5763) <= a;
    layer0_outputs(5764) <= not a or b;
    layer0_outputs(5765) <= a or b;
    layer0_outputs(5766) <= not (a or b);
    layer0_outputs(5767) <= not (a xor b);
    layer0_outputs(5768) <= not a;
    layer0_outputs(5769) <= not b;
    layer0_outputs(5770) <= not (a and b);
    layer0_outputs(5771) <= not a;
    layer0_outputs(5772) <= a;
    layer0_outputs(5773) <= '1';
    layer0_outputs(5774) <= b;
    layer0_outputs(5775) <= not (a or b);
    layer0_outputs(5776) <= a;
    layer0_outputs(5777) <= not a;
    layer0_outputs(5778) <= a or b;
    layer0_outputs(5779) <= a or b;
    layer0_outputs(5780) <= a;
    layer0_outputs(5781) <= a;
    layer0_outputs(5782) <= not b or a;
    layer0_outputs(5783) <= a and b;
    layer0_outputs(5784) <= a xor b;
    layer0_outputs(5785) <= a;
    layer0_outputs(5786) <= a and not b;
    layer0_outputs(5787) <= a xor b;
    layer0_outputs(5788) <= not (a xor b);
    layer0_outputs(5789) <= b and not a;
    layer0_outputs(5790) <= a or b;
    layer0_outputs(5791) <= not (a xor b);
    layer0_outputs(5792) <= not b;
    layer0_outputs(5793) <= '0';
    layer0_outputs(5794) <= not a or b;
    layer0_outputs(5795) <= b;
    layer0_outputs(5796) <= not (a or b);
    layer0_outputs(5797) <= not (a or b);
    layer0_outputs(5798) <= not a;
    layer0_outputs(5799) <= a xor b;
    layer0_outputs(5800) <= not (a or b);
    layer0_outputs(5801) <= not (a or b);
    layer0_outputs(5802) <= not (a or b);
    layer0_outputs(5803) <= a and not b;
    layer0_outputs(5804) <= a or b;
    layer0_outputs(5805) <= not a;
    layer0_outputs(5806) <= not (a or b);
    layer0_outputs(5807) <= b;
    layer0_outputs(5808) <= b;
    layer0_outputs(5809) <= b and not a;
    layer0_outputs(5810) <= a or b;
    layer0_outputs(5811) <= not (a or b);
    layer0_outputs(5812) <= a or b;
    layer0_outputs(5813) <= a;
    layer0_outputs(5814) <= b and not a;
    layer0_outputs(5815) <= a and b;
    layer0_outputs(5816) <= not b;
    layer0_outputs(5817) <= b;
    layer0_outputs(5818) <= a or b;
    layer0_outputs(5819) <= not a;
    layer0_outputs(5820) <= not (a or b);
    layer0_outputs(5821) <= not (a xor b);
    layer0_outputs(5822) <= not a or b;
    layer0_outputs(5823) <= a and not b;
    layer0_outputs(5824) <= b and not a;
    layer0_outputs(5825) <= not a or b;
    layer0_outputs(5826) <= a and not b;
    layer0_outputs(5827) <= a xor b;
    layer0_outputs(5828) <= not (a or b);
    layer0_outputs(5829) <= a or b;
    layer0_outputs(5830) <= b;
    layer0_outputs(5831) <= not (a or b);
    layer0_outputs(5832) <= not (a or b);
    layer0_outputs(5833) <= a or b;
    layer0_outputs(5834) <= a and not b;
    layer0_outputs(5835) <= a xor b;
    layer0_outputs(5836) <= a xor b;
    layer0_outputs(5837) <= b;
    layer0_outputs(5838) <= b;
    layer0_outputs(5839) <= not b or a;
    layer0_outputs(5840) <= not b;
    layer0_outputs(5841) <= not b or a;
    layer0_outputs(5842) <= not b;
    layer0_outputs(5843) <= not (a or b);
    layer0_outputs(5844) <= a xor b;
    layer0_outputs(5845) <= '1';
    layer0_outputs(5846) <= a xor b;
    layer0_outputs(5847) <= not b or a;
    layer0_outputs(5848) <= a;
    layer0_outputs(5849) <= a;
    layer0_outputs(5850) <= a and not b;
    layer0_outputs(5851) <= a xor b;
    layer0_outputs(5852) <= not b or a;
    layer0_outputs(5853) <= a and not b;
    layer0_outputs(5854) <= not (a or b);
    layer0_outputs(5855) <= not (a xor b);
    layer0_outputs(5856) <= not a;
    layer0_outputs(5857) <= b;
    layer0_outputs(5858) <= not (a and b);
    layer0_outputs(5859) <= not a;
    layer0_outputs(5860) <= a or b;
    layer0_outputs(5861) <= not (a xor b);
    layer0_outputs(5862) <= not (a or b);
    layer0_outputs(5863) <= a xor b;
    layer0_outputs(5864) <= not b or a;
    layer0_outputs(5865) <= a or b;
    layer0_outputs(5866) <= a;
    layer0_outputs(5867) <= a or b;
    layer0_outputs(5868) <= a;
    layer0_outputs(5869) <= not b;
    layer0_outputs(5870) <= not (a xor b);
    layer0_outputs(5871) <= a or b;
    layer0_outputs(5872) <= a and b;
    layer0_outputs(5873) <= b and not a;
    layer0_outputs(5874) <= a and not b;
    layer0_outputs(5875) <= b;
    layer0_outputs(5876) <= not (a and b);
    layer0_outputs(5877) <= not b or a;
    layer0_outputs(5878) <= a and not b;
    layer0_outputs(5879) <= not (a or b);
    layer0_outputs(5880) <= b;
    layer0_outputs(5881) <= not b;
    layer0_outputs(5882) <= '1';
    layer0_outputs(5883) <= '0';
    layer0_outputs(5884) <= not (a and b);
    layer0_outputs(5885) <= b;
    layer0_outputs(5886) <= a xor b;
    layer0_outputs(5887) <= not (a or b);
    layer0_outputs(5888) <= not b or a;
    layer0_outputs(5889) <= b and not a;
    layer0_outputs(5890) <= not (a or b);
    layer0_outputs(5891) <= b and not a;
    layer0_outputs(5892) <= a or b;
    layer0_outputs(5893) <= a xor b;
    layer0_outputs(5894) <= '1';
    layer0_outputs(5895) <= not (a or b);
    layer0_outputs(5896) <= not a;
    layer0_outputs(5897) <= not (a xor b);
    layer0_outputs(5898) <= b and not a;
    layer0_outputs(5899) <= b and not a;
    layer0_outputs(5900) <= a;
    layer0_outputs(5901) <= a;
    layer0_outputs(5902) <= not b or a;
    layer0_outputs(5903) <= not a;
    layer0_outputs(5904) <= b;
    layer0_outputs(5905) <= not (a xor b);
    layer0_outputs(5906) <= a;
    layer0_outputs(5907) <= a or b;
    layer0_outputs(5908) <= not (a or b);
    layer0_outputs(5909) <= a or b;
    layer0_outputs(5910) <= a;
    layer0_outputs(5911) <= not a;
    layer0_outputs(5912) <= b;
    layer0_outputs(5913) <= a and b;
    layer0_outputs(5914) <= not a;
    layer0_outputs(5915) <= a and b;
    layer0_outputs(5916) <= a;
    layer0_outputs(5917) <= not b or a;
    layer0_outputs(5918) <= a or b;
    layer0_outputs(5919) <= not a or b;
    layer0_outputs(5920) <= a xor b;
    layer0_outputs(5921) <= a and not b;
    layer0_outputs(5922) <= not (a or b);
    layer0_outputs(5923) <= a and b;
    layer0_outputs(5924) <= not (a xor b);
    layer0_outputs(5925) <= not (a or b);
    layer0_outputs(5926) <= a;
    layer0_outputs(5927) <= a and not b;
    layer0_outputs(5928) <= a;
    layer0_outputs(5929) <= a or b;
    layer0_outputs(5930) <= b;
    layer0_outputs(5931) <= not (a xor b);
    layer0_outputs(5932) <= not (a xor b);
    layer0_outputs(5933) <= a or b;
    layer0_outputs(5934) <= '1';
    layer0_outputs(5935) <= a xor b;
    layer0_outputs(5936) <= a;
    layer0_outputs(5937) <= '0';
    layer0_outputs(5938) <= b;
    layer0_outputs(5939) <= a and not b;
    layer0_outputs(5940) <= not (a xor b);
    layer0_outputs(5941) <= not b;
    layer0_outputs(5942) <= a and not b;
    layer0_outputs(5943) <= not a;
    layer0_outputs(5944) <= not (a or b);
    layer0_outputs(5945) <= not (a xor b);
    layer0_outputs(5946) <= not a or b;
    layer0_outputs(5947) <= b;
    layer0_outputs(5948) <= a;
    layer0_outputs(5949) <= not (a or b);
    layer0_outputs(5950) <= b;
    layer0_outputs(5951) <= not (a or b);
    layer0_outputs(5952) <= a and not b;
    layer0_outputs(5953) <= a xor b;
    layer0_outputs(5954) <= '1';
    layer0_outputs(5955) <= a;
    layer0_outputs(5956) <= not (a xor b);
    layer0_outputs(5957) <= not a;
    layer0_outputs(5958) <= '0';
    layer0_outputs(5959) <= not a;
    layer0_outputs(5960) <= not b or a;
    layer0_outputs(5961) <= b;
    layer0_outputs(5962) <= not (a or b);
    layer0_outputs(5963) <= not (a or b);
    layer0_outputs(5964) <= b and not a;
    layer0_outputs(5965) <= not a;
    layer0_outputs(5966) <= a xor b;
    layer0_outputs(5967) <= a;
    layer0_outputs(5968) <= a xor b;
    layer0_outputs(5969) <= a or b;
    layer0_outputs(5970) <= not (a and b);
    layer0_outputs(5971) <= not (a xor b);
    layer0_outputs(5972) <= not a or b;
    layer0_outputs(5973) <= not b or a;
    layer0_outputs(5974) <= a or b;
    layer0_outputs(5975) <= not a;
    layer0_outputs(5976) <= not b or a;
    layer0_outputs(5977) <= a and b;
    layer0_outputs(5978) <= a or b;
    layer0_outputs(5979) <= not a or b;
    layer0_outputs(5980) <= '0';
    layer0_outputs(5981) <= b;
    layer0_outputs(5982) <= a and not b;
    layer0_outputs(5983) <= not (a or b);
    layer0_outputs(5984) <= b;
    layer0_outputs(5985) <= a or b;
    layer0_outputs(5986) <= a xor b;
    layer0_outputs(5987) <= a and not b;
    layer0_outputs(5988) <= not (a or b);
    layer0_outputs(5989) <= b;
    layer0_outputs(5990) <= a or b;
    layer0_outputs(5991) <= not (a or b);
    layer0_outputs(5992) <= not b or a;
    layer0_outputs(5993) <= not a or b;
    layer0_outputs(5994) <= not (a and b);
    layer0_outputs(5995) <= not a;
    layer0_outputs(5996) <= not a or b;
    layer0_outputs(5997) <= b and not a;
    layer0_outputs(5998) <= a xor b;
    layer0_outputs(5999) <= not (a or b);
    layer0_outputs(6000) <= not a;
    layer0_outputs(6001) <= not (a or b);
    layer0_outputs(6002) <= not b or a;
    layer0_outputs(6003) <= b and not a;
    layer0_outputs(6004) <= a or b;
    layer0_outputs(6005) <= a;
    layer0_outputs(6006) <= not (a xor b);
    layer0_outputs(6007) <= not a or b;
    layer0_outputs(6008) <= a or b;
    layer0_outputs(6009) <= not a;
    layer0_outputs(6010) <= a or b;
    layer0_outputs(6011) <= not a;
    layer0_outputs(6012) <= not b or a;
    layer0_outputs(6013) <= a xor b;
    layer0_outputs(6014) <= a xor b;
    layer0_outputs(6015) <= b and not a;
    layer0_outputs(6016) <= a;
    layer0_outputs(6017) <= a and not b;
    layer0_outputs(6018) <= b and not a;
    layer0_outputs(6019) <= not b or a;
    layer0_outputs(6020) <= b and not a;
    layer0_outputs(6021) <= not a or b;
    layer0_outputs(6022) <= not a;
    layer0_outputs(6023) <= a xor b;
    layer0_outputs(6024) <= b and not a;
    layer0_outputs(6025) <= not (a and b);
    layer0_outputs(6026) <= b and not a;
    layer0_outputs(6027) <= b;
    layer0_outputs(6028) <= a or b;
    layer0_outputs(6029) <= not (a or b);
    layer0_outputs(6030) <= not (a or b);
    layer0_outputs(6031) <= b and not a;
    layer0_outputs(6032) <= a or b;
    layer0_outputs(6033) <= not a;
    layer0_outputs(6034) <= a xor b;
    layer0_outputs(6035) <= not b or a;
    layer0_outputs(6036) <= not a;
    layer0_outputs(6037) <= not (a or b);
    layer0_outputs(6038) <= not b;
    layer0_outputs(6039) <= not b;
    layer0_outputs(6040) <= a;
    layer0_outputs(6041) <= a xor b;
    layer0_outputs(6042) <= not b or a;
    layer0_outputs(6043) <= a and b;
    layer0_outputs(6044) <= not (a xor b);
    layer0_outputs(6045) <= not b;
    layer0_outputs(6046) <= a;
    layer0_outputs(6047) <= not a or b;
    layer0_outputs(6048) <= not (a xor b);
    layer0_outputs(6049) <= a and not b;
    layer0_outputs(6050) <= a and not b;
    layer0_outputs(6051) <= not b;
    layer0_outputs(6052) <= a;
    layer0_outputs(6053) <= not (a or b);
    layer0_outputs(6054) <= not b or a;
    layer0_outputs(6055) <= a or b;
    layer0_outputs(6056) <= not (a xor b);
    layer0_outputs(6057) <= a and not b;
    layer0_outputs(6058) <= a and not b;
    layer0_outputs(6059) <= not (a and b);
    layer0_outputs(6060) <= not (a and b);
    layer0_outputs(6061) <= not (a and b);
    layer0_outputs(6062) <= a or b;
    layer0_outputs(6063) <= not b or a;
    layer0_outputs(6064) <= not (a or b);
    layer0_outputs(6065) <= a and not b;
    layer0_outputs(6066) <= a or b;
    layer0_outputs(6067) <= a xor b;
    layer0_outputs(6068) <= b;
    layer0_outputs(6069) <= a or b;
    layer0_outputs(6070) <= a xor b;
    layer0_outputs(6071) <= a and not b;
    layer0_outputs(6072) <= not (a or b);
    layer0_outputs(6073) <= not (a or b);
    layer0_outputs(6074) <= a;
    layer0_outputs(6075) <= not a or b;
    layer0_outputs(6076) <= not a or b;
    layer0_outputs(6077) <= a or b;
    layer0_outputs(6078) <= not b or a;
    layer0_outputs(6079) <= a or b;
    layer0_outputs(6080) <= a or b;
    layer0_outputs(6081) <= not (a or b);
    layer0_outputs(6082) <= a xor b;
    layer0_outputs(6083) <= a xor b;
    layer0_outputs(6084) <= b and not a;
    layer0_outputs(6085) <= not (a xor b);
    layer0_outputs(6086) <= not (a xor b);
    layer0_outputs(6087) <= '0';
    layer0_outputs(6088) <= not (a or b);
    layer0_outputs(6089) <= not (a or b);
    layer0_outputs(6090) <= a;
    layer0_outputs(6091) <= a or b;
    layer0_outputs(6092) <= a or b;
    layer0_outputs(6093) <= a xor b;
    layer0_outputs(6094) <= a and b;
    layer0_outputs(6095) <= not (a or b);
    layer0_outputs(6096) <= not b;
    layer0_outputs(6097) <= b and not a;
    layer0_outputs(6098) <= not a or b;
    layer0_outputs(6099) <= a xor b;
    layer0_outputs(6100) <= b;
    layer0_outputs(6101) <= b and not a;
    layer0_outputs(6102) <= not b or a;
    layer0_outputs(6103) <= not b or a;
    layer0_outputs(6104) <= a and not b;
    layer0_outputs(6105) <= a xor b;
    layer0_outputs(6106) <= not a or b;
    layer0_outputs(6107) <= not a or b;
    layer0_outputs(6108) <= a or b;
    layer0_outputs(6109) <= not b;
    layer0_outputs(6110) <= a or b;
    layer0_outputs(6111) <= a or b;
    layer0_outputs(6112) <= not (a xor b);
    layer0_outputs(6113) <= not b;
    layer0_outputs(6114) <= b;
    layer0_outputs(6115) <= a or b;
    layer0_outputs(6116) <= not a;
    layer0_outputs(6117) <= not b or a;
    layer0_outputs(6118) <= a xor b;
    layer0_outputs(6119) <= a xor b;
    layer0_outputs(6120) <= b and not a;
    layer0_outputs(6121) <= a;
    layer0_outputs(6122) <= a and not b;
    layer0_outputs(6123) <= not (a and b);
    layer0_outputs(6124) <= '1';
    layer0_outputs(6125) <= a xor b;
    layer0_outputs(6126) <= not a or b;
    layer0_outputs(6127) <= not a or b;
    layer0_outputs(6128) <= a or b;
    layer0_outputs(6129) <= not (a xor b);
    layer0_outputs(6130) <= not b or a;
    layer0_outputs(6131) <= not b;
    layer0_outputs(6132) <= a and b;
    layer0_outputs(6133) <= not a;
    layer0_outputs(6134) <= not a;
    layer0_outputs(6135) <= not (a or b);
    layer0_outputs(6136) <= a xor b;
    layer0_outputs(6137) <= not (a and b);
    layer0_outputs(6138) <= b;
    layer0_outputs(6139) <= not (a xor b);
    layer0_outputs(6140) <= not (a xor b);
    layer0_outputs(6141) <= a or b;
    layer0_outputs(6142) <= a and not b;
    layer0_outputs(6143) <= a or b;
    layer0_outputs(6144) <= a xor b;
    layer0_outputs(6145) <= a and not b;
    layer0_outputs(6146) <= a xor b;
    layer0_outputs(6147) <= b;
    layer0_outputs(6148) <= not b;
    layer0_outputs(6149) <= a or b;
    layer0_outputs(6150) <= a xor b;
    layer0_outputs(6151) <= not b or a;
    layer0_outputs(6152) <= not (a or b);
    layer0_outputs(6153) <= a or b;
    layer0_outputs(6154) <= a or b;
    layer0_outputs(6155) <= not (a and b);
    layer0_outputs(6156) <= '0';
    layer0_outputs(6157) <= not a or b;
    layer0_outputs(6158) <= a and b;
    layer0_outputs(6159) <= a or b;
    layer0_outputs(6160) <= not a or b;
    layer0_outputs(6161) <= a or b;
    layer0_outputs(6162) <= a or b;
    layer0_outputs(6163) <= a xor b;
    layer0_outputs(6164) <= a or b;
    layer0_outputs(6165) <= a and not b;
    layer0_outputs(6166) <= a and not b;
    layer0_outputs(6167) <= '1';
    layer0_outputs(6168) <= a;
    layer0_outputs(6169) <= not (a or b);
    layer0_outputs(6170) <= not a;
    layer0_outputs(6171) <= a or b;
    layer0_outputs(6172) <= not (a xor b);
    layer0_outputs(6173) <= a xor b;
    layer0_outputs(6174) <= not a or b;
    layer0_outputs(6175) <= not b or a;
    layer0_outputs(6176) <= not b;
    layer0_outputs(6177) <= not (a or b);
    layer0_outputs(6178) <= b;
    layer0_outputs(6179) <= not (a or b);
    layer0_outputs(6180) <= a and not b;
    layer0_outputs(6181) <= not a or b;
    layer0_outputs(6182) <= not a;
    layer0_outputs(6183) <= not (a xor b);
    layer0_outputs(6184) <= not (a or b);
    layer0_outputs(6185) <= not (a or b);
    layer0_outputs(6186) <= a;
    layer0_outputs(6187) <= not (a xor b);
    layer0_outputs(6188) <= a;
    layer0_outputs(6189) <= a xor b;
    layer0_outputs(6190) <= not (a or b);
    layer0_outputs(6191) <= a;
    layer0_outputs(6192) <= not (a and b);
    layer0_outputs(6193) <= a or b;
    layer0_outputs(6194) <= a or b;
    layer0_outputs(6195) <= not a or b;
    layer0_outputs(6196) <= not a or b;
    layer0_outputs(6197) <= a and not b;
    layer0_outputs(6198) <= a or b;
    layer0_outputs(6199) <= b and not a;
    layer0_outputs(6200) <= not a;
    layer0_outputs(6201) <= a and not b;
    layer0_outputs(6202) <= a and b;
    layer0_outputs(6203) <= a xor b;
    layer0_outputs(6204) <= not a;
    layer0_outputs(6205) <= a and not b;
    layer0_outputs(6206) <= not (a or b);
    layer0_outputs(6207) <= b;
    layer0_outputs(6208) <= '0';
    layer0_outputs(6209) <= b and not a;
    layer0_outputs(6210) <= a;
    layer0_outputs(6211) <= not (a or b);
    layer0_outputs(6212) <= not (a or b);
    layer0_outputs(6213) <= not (a or b);
    layer0_outputs(6214) <= not b;
    layer0_outputs(6215) <= a or b;
    layer0_outputs(6216) <= a or b;
    layer0_outputs(6217) <= a xor b;
    layer0_outputs(6218) <= a xor b;
    layer0_outputs(6219) <= a xor b;
    layer0_outputs(6220) <= not (a or b);
    layer0_outputs(6221) <= not (a or b);
    layer0_outputs(6222) <= a and not b;
    layer0_outputs(6223) <= a and not b;
    layer0_outputs(6224) <= not (a and b);
    layer0_outputs(6225) <= not (a and b);
    layer0_outputs(6226) <= not (a or b);
    layer0_outputs(6227) <= not b or a;
    layer0_outputs(6228) <= b and not a;
    layer0_outputs(6229) <= a xor b;
    layer0_outputs(6230) <= a and not b;
    layer0_outputs(6231) <= a;
    layer0_outputs(6232) <= not b;
    layer0_outputs(6233) <= a;
    layer0_outputs(6234) <= a;
    layer0_outputs(6235) <= not (a xor b);
    layer0_outputs(6236) <= a;
    layer0_outputs(6237) <= a or b;
    layer0_outputs(6238) <= not (a xor b);
    layer0_outputs(6239) <= not (a xor b);
    layer0_outputs(6240) <= '1';
    layer0_outputs(6241) <= a or b;
    layer0_outputs(6242) <= not a;
    layer0_outputs(6243) <= '1';
    layer0_outputs(6244) <= not (a or b);
    layer0_outputs(6245) <= a or b;
    layer0_outputs(6246) <= not a or b;
    layer0_outputs(6247) <= not b or a;
    layer0_outputs(6248) <= not (a xor b);
    layer0_outputs(6249) <= not (a xor b);
    layer0_outputs(6250) <= not b or a;
    layer0_outputs(6251) <= a or b;
    layer0_outputs(6252) <= not b;
    layer0_outputs(6253) <= not (a or b);
    layer0_outputs(6254) <= not a or b;
    layer0_outputs(6255) <= a and not b;
    layer0_outputs(6256) <= not (a and b);
    layer0_outputs(6257) <= not (a or b);
    layer0_outputs(6258) <= not (a and b);
    layer0_outputs(6259) <= not (a xor b);
    layer0_outputs(6260) <= a xor b;
    layer0_outputs(6261) <= not (a or b);
    layer0_outputs(6262) <= a;
    layer0_outputs(6263) <= '1';
    layer0_outputs(6264) <= not a or b;
    layer0_outputs(6265) <= not (a xor b);
    layer0_outputs(6266) <= a xor b;
    layer0_outputs(6267) <= not (a xor b);
    layer0_outputs(6268) <= not b;
    layer0_outputs(6269) <= not (a or b);
    layer0_outputs(6270) <= b;
    layer0_outputs(6271) <= a xor b;
    layer0_outputs(6272) <= not a;
    layer0_outputs(6273) <= a;
    layer0_outputs(6274) <= a and not b;
    layer0_outputs(6275) <= b and not a;
    layer0_outputs(6276) <= a or b;
    layer0_outputs(6277) <= not (a xor b);
    layer0_outputs(6278) <= a or b;
    layer0_outputs(6279) <= a;
    layer0_outputs(6280) <= a xor b;
    layer0_outputs(6281) <= b and not a;
    layer0_outputs(6282) <= not a or b;
    layer0_outputs(6283) <= not b or a;
    layer0_outputs(6284) <= b;
    layer0_outputs(6285) <= b and not a;
    layer0_outputs(6286) <= a and not b;
    layer0_outputs(6287) <= not b;
    layer0_outputs(6288) <= not b or a;
    layer0_outputs(6289) <= b;
    layer0_outputs(6290) <= not a or b;
    layer0_outputs(6291) <= not (a xor b);
    layer0_outputs(6292) <= a and not b;
    layer0_outputs(6293) <= not a or b;
    layer0_outputs(6294) <= not (a or b);
    layer0_outputs(6295) <= not (a or b);
    layer0_outputs(6296) <= b;
    layer0_outputs(6297) <= a xor b;
    layer0_outputs(6298) <= not a or b;
    layer0_outputs(6299) <= not a;
    layer0_outputs(6300) <= a;
    layer0_outputs(6301) <= a xor b;
    layer0_outputs(6302) <= a or b;
    layer0_outputs(6303) <= not (a xor b);
    layer0_outputs(6304) <= b;
    layer0_outputs(6305) <= not (a or b);
    layer0_outputs(6306) <= a xor b;
    layer0_outputs(6307) <= b;
    layer0_outputs(6308) <= not a or b;
    layer0_outputs(6309) <= a and not b;
    layer0_outputs(6310) <= not a or b;
    layer0_outputs(6311) <= not (a xor b);
    layer0_outputs(6312) <= not (a xor b);
    layer0_outputs(6313) <= a or b;
    layer0_outputs(6314) <= a and b;
    layer0_outputs(6315) <= a or b;
    layer0_outputs(6316) <= not (a and b);
    layer0_outputs(6317) <= a xor b;
    layer0_outputs(6318) <= a or b;
    layer0_outputs(6319) <= b;
    layer0_outputs(6320) <= not a or b;
    layer0_outputs(6321) <= not a or b;
    layer0_outputs(6322) <= a or b;
    layer0_outputs(6323) <= not (a xor b);
    layer0_outputs(6324) <= not b or a;
    layer0_outputs(6325) <= b;
    layer0_outputs(6326) <= not (a or b);
    layer0_outputs(6327) <= a;
    layer0_outputs(6328) <= not (a xor b);
    layer0_outputs(6329) <= a or b;
    layer0_outputs(6330) <= not (a or b);
    layer0_outputs(6331) <= '1';
    layer0_outputs(6332) <= a and not b;
    layer0_outputs(6333) <= a xor b;
    layer0_outputs(6334) <= not a or b;
    layer0_outputs(6335) <= a and not b;
    layer0_outputs(6336) <= not a or b;
    layer0_outputs(6337) <= not (a or b);
    layer0_outputs(6338) <= not (a xor b);
    layer0_outputs(6339) <= not (a xor b);
    layer0_outputs(6340) <= a;
    layer0_outputs(6341) <= b;
    layer0_outputs(6342) <= a or b;
    layer0_outputs(6343) <= b and not a;
    layer0_outputs(6344) <= not b or a;
    layer0_outputs(6345) <= b and not a;
    layer0_outputs(6346) <= not b;
    layer0_outputs(6347) <= not b;
    layer0_outputs(6348) <= '1';
    layer0_outputs(6349) <= not a;
    layer0_outputs(6350) <= a;
    layer0_outputs(6351) <= a or b;
    layer0_outputs(6352) <= not a;
    layer0_outputs(6353) <= b;
    layer0_outputs(6354) <= a or b;
    layer0_outputs(6355) <= not b;
    layer0_outputs(6356) <= a and not b;
    layer0_outputs(6357) <= not (a or b);
    layer0_outputs(6358) <= not (a xor b);
    layer0_outputs(6359) <= a or b;
    layer0_outputs(6360) <= a or b;
    layer0_outputs(6361) <= not (a or b);
    layer0_outputs(6362) <= not a or b;
    layer0_outputs(6363) <= not b or a;
    layer0_outputs(6364) <= not a;
    layer0_outputs(6365) <= '0';
    layer0_outputs(6366) <= not b or a;
    layer0_outputs(6367) <= not a;
    layer0_outputs(6368) <= not a or b;
    layer0_outputs(6369) <= not (a or b);
    layer0_outputs(6370) <= not (a and b);
    layer0_outputs(6371) <= not (a or b);
    layer0_outputs(6372) <= b;
    layer0_outputs(6373) <= not a or b;
    layer0_outputs(6374) <= b and not a;
    layer0_outputs(6375) <= not b;
    layer0_outputs(6376) <= b;
    layer0_outputs(6377) <= not a;
    layer0_outputs(6378) <= not (a or b);
    layer0_outputs(6379) <= not b or a;
    layer0_outputs(6380) <= not b;
    layer0_outputs(6381) <= a or b;
    layer0_outputs(6382) <= not (a xor b);
    layer0_outputs(6383) <= '0';
    layer0_outputs(6384) <= a xor b;
    layer0_outputs(6385) <= a xor b;
    layer0_outputs(6386) <= not (a xor b);
    layer0_outputs(6387) <= a and not b;
    layer0_outputs(6388) <= a xor b;
    layer0_outputs(6389) <= not (a or b);
    layer0_outputs(6390) <= not (a xor b);
    layer0_outputs(6391) <= '0';
    layer0_outputs(6392) <= a or b;
    layer0_outputs(6393) <= a xor b;
    layer0_outputs(6394) <= a or b;
    layer0_outputs(6395) <= b and not a;
    layer0_outputs(6396) <= not a or b;
    layer0_outputs(6397) <= '0';
    layer0_outputs(6398) <= a or b;
    layer0_outputs(6399) <= not (a or b);
    layer0_outputs(6400) <= a xor b;
    layer0_outputs(6401) <= b and not a;
    layer0_outputs(6402) <= not b;
    layer0_outputs(6403) <= '1';
    layer0_outputs(6404) <= not b;
    layer0_outputs(6405) <= a or b;
    layer0_outputs(6406) <= not b or a;
    layer0_outputs(6407) <= not b;
    layer0_outputs(6408) <= not (a and b);
    layer0_outputs(6409) <= a;
    layer0_outputs(6410) <= a;
    layer0_outputs(6411) <= a or b;
    layer0_outputs(6412) <= not a;
    layer0_outputs(6413) <= not a or b;
    layer0_outputs(6414) <= not b or a;
    layer0_outputs(6415) <= a;
    layer0_outputs(6416) <= not b or a;
    layer0_outputs(6417) <= '1';
    layer0_outputs(6418) <= a xor b;
    layer0_outputs(6419) <= a xor b;
    layer0_outputs(6420) <= b and not a;
    layer0_outputs(6421) <= not a;
    layer0_outputs(6422) <= b;
    layer0_outputs(6423) <= a or b;
    layer0_outputs(6424) <= a or b;
    layer0_outputs(6425) <= a;
    layer0_outputs(6426) <= not a;
    layer0_outputs(6427) <= b;
    layer0_outputs(6428) <= not (a and b);
    layer0_outputs(6429) <= a xor b;
    layer0_outputs(6430) <= a;
    layer0_outputs(6431) <= a or b;
    layer0_outputs(6432) <= a xor b;
    layer0_outputs(6433) <= b;
    layer0_outputs(6434) <= not a;
    layer0_outputs(6435) <= a or b;
    layer0_outputs(6436) <= a or b;
    layer0_outputs(6437) <= not (a or b);
    layer0_outputs(6438) <= not (a xor b);
    layer0_outputs(6439) <= not (a xor b);
    layer0_outputs(6440) <= not b;
    layer0_outputs(6441) <= b and not a;
    layer0_outputs(6442) <= not (a or b);
    layer0_outputs(6443) <= a;
    layer0_outputs(6444) <= not (a or b);
    layer0_outputs(6445) <= a;
    layer0_outputs(6446) <= b and not a;
    layer0_outputs(6447) <= not b;
    layer0_outputs(6448) <= a and not b;
    layer0_outputs(6449) <= not (a or b);
    layer0_outputs(6450) <= not (a or b);
    layer0_outputs(6451) <= a or b;
    layer0_outputs(6452) <= b;
    layer0_outputs(6453) <= a;
    layer0_outputs(6454) <= a and not b;
    layer0_outputs(6455) <= a;
    layer0_outputs(6456) <= not (a or b);
    layer0_outputs(6457) <= b;
    layer0_outputs(6458) <= not (a xor b);
    layer0_outputs(6459) <= not b;
    layer0_outputs(6460) <= not (a or b);
    layer0_outputs(6461) <= a xor b;
    layer0_outputs(6462) <= not (a or b);
    layer0_outputs(6463) <= a and b;
    layer0_outputs(6464) <= not (a or b);
    layer0_outputs(6465) <= b;
    layer0_outputs(6466) <= not b;
    layer0_outputs(6467) <= not a;
    layer0_outputs(6468) <= a and b;
    layer0_outputs(6469) <= a;
    layer0_outputs(6470) <= not (a xor b);
    layer0_outputs(6471) <= not b;
    layer0_outputs(6472) <= a and not b;
    layer0_outputs(6473) <= a xor b;
    layer0_outputs(6474) <= not (a or b);
    layer0_outputs(6475) <= b and not a;
    layer0_outputs(6476) <= b and not a;
    layer0_outputs(6477) <= a and not b;
    layer0_outputs(6478) <= '1';
    layer0_outputs(6479) <= not b;
    layer0_outputs(6480) <= a or b;
    layer0_outputs(6481) <= a or b;
    layer0_outputs(6482) <= a xor b;
    layer0_outputs(6483) <= a and b;
    layer0_outputs(6484) <= a;
    layer0_outputs(6485) <= a and not b;
    layer0_outputs(6486) <= not a or b;
    layer0_outputs(6487) <= b and not a;
    layer0_outputs(6488) <= a and not b;
    layer0_outputs(6489) <= b;
    layer0_outputs(6490) <= b;
    layer0_outputs(6491) <= '1';
    layer0_outputs(6492) <= '1';
    layer0_outputs(6493) <= a or b;
    layer0_outputs(6494) <= a and not b;
    layer0_outputs(6495) <= a and not b;
    layer0_outputs(6496) <= a or b;
    layer0_outputs(6497) <= not a;
    layer0_outputs(6498) <= a or b;
    layer0_outputs(6499) <= a or b;
    layer0_outputs(6500) <= a xor b;
    layer0_outputs(6501) <= b;
    layer0_outputs(6502) <= not a;
    layer0_outputs(6503) <= not b;
    layer0_outputs(6504) <= a or b;
    layer0_outputs(6505) <= not a;
    layer0_outputs(6506) <= not a or b;
    layer0_outputs(6507) <= not (a and b);
    layer0_outputs(6508) <= a xor b;
    layer0_outputs(6509) <= b;
    layer0_outputs(6510) <= a and not b;
    layer0_outputs(6511) <= not b;
    layer0_outputs(6512) <= b and not a;
    layer0_outputs(6513) <= a;
    layer0_outputs(6514) <= not a;
    layer0_outputs(6515) <= not (a xor b);
    layer0_outputs(6516) <= b and not a;
    layer0_outputs(6517) <= a xor b;
    layer0_outputs(6518) <= not a;
    layer0_outputs(6519) <= a xor b;
    layer0_outputs(6520) <= not (a or b);
    layer0_outputs(6521) <= a or b;
    layer0_outputs(6522) <= not a;
    layer0_outputs(6523) <= a and b;
    layer0_outputs(6524) <= not (a xor b);
    layer0_outputs(6525) <= not (a and b);
    layer0_outputs(6526) <= not a;
    layer0_outputs(6527) <= a or b;
    layer0_outputs(6528) <= b;
    layer0_outputs(6529) <= not a or b;
    layer0_outputs(6530) <= not (a xor b);
    layer0_outputs(6531) <= not a or b;
    layer0_outputs(6532) <= not a or b;
    layer0_outputs(6533) <= not a;
    layer0_outputs(6534) <= a or b;
    layer0_outputs(6535) <= not b;
    layer0_outputs(6536) <= not (a xor b);
    layer0_outputs(6537) <= not b or a;
    layer0_outputs(6538) <= not b or a;
    layer0_outputs(6539) <= b and not a;
    layer0_outputs(6540) <= b;
    layer0_outputs(6541) <= not b;
    layer0_outputs(6542) <= a;
    layer0_outputs(6543) <= a or b;
    layer0_outputs(6544) <= not a;
    layer0_outputs(6545) <= a or b;
    layer0_outputs(6546) <= a or b;
    layer0_outputs(6547) <= not b;
    layer0_outputs(6548) <= not (a xor b);
    layer0_outputs(6549) <= a or b;
    layer0_outputs(6550) <= a or b;
    layer0_outputs(6551) <= not (a xor b);
    layer0_outputs(6552) <= a and not b;
    layer0_outputs(6553) <= not b;
    layer0_outputs(6554) <= not (a or b);
    layer0_outputs(6555) <= not a or b;
    layer0_outputs(6556) <= a and not b;
    layer0_outputs(6557) <= a;
    layer0_outputs(6558) <= a or b;
    layer0_outputs(6559) <= not (a or b);
    layer0_outputs(6560) <= not (a or b);
    layer0_outputs(6561) <= not a or b;
    layer0_outputs(6562) <= not (a xor b);
    layer0_outputs(6563) <= '0';
    layer0_outputs(6564) <= not (a or b);
    layer0_outputs(6565) <= not a;
    layer0_outputs(6566) <= a xor b;
    layer0_outputs(6567) <= a or b;
    layer0_outputs(6568) <= not b or a;
    layer0_outputs(6569) <= not (a xor b);
    layer0_outputs(6570) <= a and not b;
    layer0_outputs(6571) <= not b;
    layer0_outputs(6572) <= not b;
    layer0_outputs(6573) <= not (a or b);
    layer0_outputs(6574) <= a;
    layer0_outputs(6575) <= not b;
    layer0_outputs(6576) <= a xor b;
    layer0_outputs(6577) <= a xor b;
    layer0_outputs(6578) <= a and b;
    layer0_outputs(6579) <= not b;
    layer0_outputs(6580) <= not a;
    layer0_outputs(6581) <= not a;
    layer0_outputs(6582) <= not b or a;
    layer0_outputs(6583) <= not b;
    layer0_outputs(6584) <= not b;
    layer0_outputs(6585) <= not (a xor b);
    layer0_outputs(6586) <= not (a or b);
    layer0_outputs(6587) <= a;
    layer0_outputs(6588) <= not (a or b);
    layer0_outputs(6589) <= b and not a;
    layer0_outputs(6590) <= a or b;
    layer0_outputs(6591) <= a xor b;
    layer0_outputs(6592) <= not (a xor b);
    layer0_outputs(6593) <= '0';
    layer0_outputs(6594) <= not (a or b);
    layer0_outputs(6595) <= '0';
    layer0_outputs(6596) <= not (a xor b);
    layer0_outputs(6597) <= a;
    layer0_outputs(6598) <= not (a or b);
    layer0_outputs(6599) <= not a;
    layer0_outputs(6600) <= not (a or b);
    layer0_outputs(6601) <= a and not b;
    layer0_outputs(6602) <= not a;
    layer0_outputs(6603) <= not (a xor b);
    layer0_outputs(6604) <= a;
    layer0_outputs(6605) <= a and not b;
    layer0_outputs(6606) <= a or b;
    layer0_outputs(6607) <= not a or b;
    layer0_outputs(6608) <= a or b;
    layer0_outputs(6609) <= a and b;
    layer0_outputs(6610) <= a xor b;
    layer0_outputs(6611) <= b and not a;
    layer0_outputs(6612) <= not (a or b);
    layer0_outputs(6613) <= not a;
    layer0_outputs(6614) <= not b or a;
    layer0_outputs(6615) <= not a;
    layer0_outputs(6616) <= not b;
    layer0_outputs(6617) <= a or b;
    layer0_outputs(6618) <= not (a or b);
    layer0_outputs(6619) <= a or b;
    layer0_outputs(6620) <= not (a or b);
    layer0_outputs(6621) <= not b or a;
    layer0_outputs(6622) <= not b;
    layer0_outputs(6623) <= a and not b;
    layer0_outputs(6624) <= not (a xor b);
    layer0_outputs(6625) <= a and not b;
    layer0_outputs(6626) <= b;
    layer0_outputs(6627) <= not (a or b);
    layer0_outputs(6628) <= not (a xor b);
    layer0_outputs(6629) <= a or b;
    layer0_outputs(6630) <= not (a or b);
    layer0_outputs(6631) <= not a;
    layer0_outputs(6632) <= a or b;
    layer0_outputs(6633) <= not (a xor b);
    layer0_outputs(6634) <= a and not b;
    layer0_outputs(6635) <= a or b;
    layer0_outputs(6636) <= not (a xor b);
    layer0_outputs(6637) <= a and not b;
    layer0_outputs(6638) <= a;
    layer0_outputs(6639) <= not (a or b);
    layer0_outputs(6640) <= not b;
    layer0_outputs(6641) <= a;
    layer0_outputs(6642) <= b and not a;
    layer0_outputs(6643) <= not (a xor b);
    layer0_outputs(6644) <= b;
    layer0_outputs(6645) <= b;
    layer0_outputs(6646) <= b and not a;
    layer0_outputs(6647) <= not (a or b);
    layer0_outputs(6648) <= a or b;
    layer0_outputs(6649) <= not a or b;
    layer0_outputs(6650) <= b and not a;
    layer0_outputs(6651) <= not b or a;
    layer0_outputs(6652) <= not b;
    layer0_outputs(6653) <= a xor b;
    layer0_outputs(6654) <= b;
    layer0_outputs(6655) <= not b or a;
    layer0_outputs(6656) <= a;
    layer0_outputs(6657) <= not a or b;
    layer0_outputs(6658) <= not b or a;
    layer0_outputs(6659) <= not a or b;
    layer0_outputs(6660) <= a;
    layer0_outputs(6661) <= not b or a;
    layer0_outputs(6662) <= not (a or b);
    layer0_outputs(6663) <= not a or b;
    layer0_outputs(6664) <= b;
    layer0_outputs(6665) <= not a;
    layer0_outputs(6666) <= not b;
    layer0_outputs(6667) <= not a or b;
    layer0_outputs(6668) <= a or b;
    layer0_outputs(6669) <= a or b;
    layer0_outputs(6670) <= a xor b;
    layer0_outputs(6671) <= '0';
    layer0_outputs(6672) <= not b;
    layer0_outputs(6673) <= b and not a;
    layer0_outputs(6674) <= b and not a;
    layer0_outputs(6675) <= not (a and b);
    layer0_outputs(6676) <= not (a or b);
    layer0_outputs(6677) <= a xor b;
    layer0_outputs(6678) <= not a;
    layer0_outputs(6679) <= a xor b;
    layer0_outputs(6680) <= not (a and b);
    layer0_outputs(6681) <= a and not b;
    layer0_outputs(6682) <= not (a or b);
    layer0_outputs(6683) <= not (a xor b);
    layer0_outputs(6684) <= b;
    layer0_outputs(6685) <= not b;
    layer0_outputs(6686) <= '0';
    layer0_outputs(6687) <= a and not b;
    layer0_outputs(6688) <= a xor b;
    layer0_outputs(6689) <= a;
    layer0_outputs(6690) <= '0';
    layer0_outputs(6691) <= b and not a;
    layer0_outputs(6692) <= b and not a;
    layer0_outputs(6693) <= a or b;
    layer0_outputs(6694) <= a or b;
    layer0_outputs(6695) <= not (a or b);
    layer0_outputs(6696) <= b and not a;
    layer0_outputs(6697) <= not b or a;
    layer0_outputs(6698) <= not b;
    layer0_outputs(6699) <= a xor b;
    layer0_outputs(6700) <= a;
    layer0_outputs(6701) <= not (a xor b);
    layer0_outputs(6702) <= '1';
    layer0_outputs(6703) <= a xor b;
    layer0_outputs(6704) <= not (a or b);
    layer0_outputs(6705) <= b;
    layer0_outputs(6706) <= a and not b;
    layer0_outputs(6707) <= a and not b;
    layer0_outputs(6708) <= a xor b;
    layer0_outputs(6709) <= a xor b;
    layer0_outputs(6710) <= not (a or b);
    layer0_outputs(6711) <= not b or a;
    layer0_outputs(6712) <= a or b;
    layer0_outputs(6713) <= a;
    layer0_outputs(6714) <= not (a or b);
    layer0_outputs(6715) <= a or b;
    layer0_outputs(6716) <= not b;
    layer0_outputs(6717) <= not (a xor b);
    layer0_outputs(6718) <= not (a xor b);
    layer0_outputs(6719) <= b;
    layer0_outputs(6720) <= not (a xor b);
    layer0_outputs(6721) <= a and not b;
    layer0_outputs(6722) <= '0';
    layer0_outputs(6723) <= not (a or b);
    layer0_outputs(6724) <= b and not a;
    layer0_outputs(6725) <= not b or a;
    layer0_outputs(6726) <= not b or a;
    layer0_outputs(6727) <= not (a xor b);
    layer0_outputs(6728) <= '1';
    layer0_outputs(6729) <= not (a xor b);
    layer0_outputs(6730) <= a xor b;
    layer0_outputs(6731) <= a or b;
    layer0_outputs(6732) <= a or b;
    layer0_outputs(6733) <= not a or b;
    layer0_outputs(6734) <= a or b;
    layer0_outputs(6735) <= a or b;
    layer0_outputs(6736) <= not b or a;
    layer0_outputs(6737) <= a or b;
    layer0_outputs(6738) <= a or b;
    layer0_outputs(6739) <= a;
    layer0_outputs(6740) <= not (a or b);
    layer0_outputs(6741) <= b;
    layer0_outputs(6742) <= a;
    layer0_outputs(6743) <= not (a xor b);
    layer0_outputs(6744) <= not (a or b);
    layer0_outputs(6745) <= b;
    layer0_outputs(6746) <= not b or a;
    layer0_outputs(6747) <= not (a or b);
    layer0_outputs(6748) <= not (a xor b);
    layer0_outputs(6749) <= a;
    layer0_outputs(6750) <= b;
    layer0_outputs(6751) <= not (a or b);
    layer0_outputs(6752) <= a;
    layer0_outputs(6753) <= not (a xor b);
    layer0_outputs(6754) <= not a;
    layer0_outputs(6755) <= not (a and b);
    layer0_outputs(6756) <= a xor b;
    layer0_outputs(6757) <= not (a or b);
    layer0_outputs(6758) <= not a or b;
    layer0_outputs(6759) <= a or b;
    layer0_outputs(6760) <= not b or a;
    layer0_outputs(6761) <= '1';
    layer0_outputs(6762) <= b and not a;
    layer0_outputs(6763) <= not (a xor b);
    layer0_outputs(6764) <= not (a xor b);
    layer0_outputs(6765) <= not a;
    layer0_outputs(6766) <= not b;
    layer0_outputs(6767) <= not (a or b);
    layer0_outputs(6768) <= not b or a;
    layer0_outputs(6769) <= not a;
    layer0_outputs(6770) <= not a or b;
    layer0_outputs(6771) <= not (a or b);
    layer0_outputs(6772) <= not (a xor b);
    layer0_outputs(6773) <= a and b;
    layer0_outputs(6774) <= b and not a;
    layer0_outputs(6775) <= '1';
    layer0_outputs(6776) <= not a;
    layer0_outputs(6777) <= not b or a;
    layer0_outputs(6778) <= a;
    layer0_outputs(6779) <= b and not a;
    layer0_outputs(6780) <= not a;
    layer0_outputs(6781) <= a and not b;
    layer0_outputs(6782) <= not b or a;
    layer0_outputs(6783) <= not a;
    layer0_outputs(6784) <= b;
    layer0_outputs(6785) <= not a;
    layer0_outputs(6786) <= not (a or b);
    layer0_outputs(6787) <= a;
    layer0_outputs(6788) <= a or b;
    layer0_outputs(6789) <= '0';
    layer0_outputs(6790) <= not (a xor b);
    layer0_outputs(6791) <= not b or a;
    layer0_outputs(6792) <= not b or a;
    layer0_outputs(6793) <= a or b;
    layer0_outputs(6794) <= '1';
    layer0_outputs(6795) <= '0';
    layer0_outputs(6796) <= not a or b;
    layer0_outputs(6797) <= a xor b;
    layer0_outputs(6798) <= a;
    layer0_outputs(6799) <= not b or a;
    layer0_outputs(6800) <= not b;
    layer0_outputs(6801) <= a or b;
    layer0_outputs(6802) <= a or b;
    layer0_outputs(6803) <= a and not b;
    layer0_outputs(6804) <= a or b;
    layer0_outputs(6805) <= not a;
    layer0_outputs(6806) <= a xor b;
    layer0_outputs(6807) <= '1';
    layer0_outputs(6808) <= a xor b;
    layer0_outputs(6809) <= not (a or b);
    layer0_outputs(6810) <= a or b;
    layer0_outputs(6811) <= a and not b;
    layer0_outputs(6812) <= not (a or b);
    layer0_outputs(6813) <= a xor b;
    layer0_outputs(6814) <= not a or b;
    layer0_outputs(6815) <= not a or b;
    layer0_outputs(6816) <= not b;
    layer0_outputs(6817) <= not a or b;
    layer0_outputs(6818) <= not (a or b);
    layer0_outputs(6819) <= not b;
    layer0_outputs(6820) <= not b;
    layer0_outputs(6821) <= '1';
    layer0_outputs(6822) <= b and not a;
    layer0_outputs(6823) <= b;
    layer0_outputs(6824) <= a and b;
    layer0_outputs(6825) <= not b or a;
    layer0_outputs(6826) <= b;
    layer0_outputs(6827) <= not (a xor b);
    layer0_outputs(6828) <= not a;
    layer0_outputs(6829) <= a or b;
    layer0_outputs(6830) <= a xor b;
    layer0_outputs(6831) <= not (a or b);
    layer0_outputs(6832) <= a;
    layer0_outputs(6833) <= not (a or b);
    layer0_outputs(6834) <= a or b;
    layer0_outputs(6835) <= b and not a;
    layer0_outputs(6836) <= '1';
    layer0_outputs(6837) <= b and not a;
    layer0_outputs(6838) <= '0';
    layer0_outputs(6839) <= not (a xor b);
    layer0_outputs(6840) <= a and b;
    layer0_outputs(6841) <= not b;
    layer0_outputs(6842) <= '1';
    layer0_outputs(6843) <= b;
    layer0_outputs(6844) <= a or b;
    layer0_outputs(6845) <= a and not b;
    layer0_outputs(6846) <= b;
    layer0_outputs(6847) <= not b;
    layer0_outputs(6848) <= a xor b;
    layer0_outputs(6849) <= a xor b;
    layer0_outputs(6850) <= not (a xor b);
    layer0_outputs(6851) <= not b;
    layer0_outputs(6852) <= not (a and b);
    layer0_outputs(6853) <= a or b;
    layer0_outputs(6854) <= '0';
    layer0_outputs(6855) <= not (a or b);
    layer0_outputs(6856) <= a and not b;
    layer0_outputs(6857) <= not a or b;
    layer0_outputs(6858) <= '1';
    layer0_outputs(6859) <= a xor b;
    layer0_outputs(6860) <= b;
    layer0_outputs(6861) <= a xor b;
    layer0_outputs(6862) <= not a;
    layer0_outputs(6863) <= a and not b;
    layer0_outputs(6864) <= not a or b;
    layer0_outputs(6865) <= a or b;
    layer0_outputs(6866) <= a xor b;
    layer0_outputs(6867) <= b;
    layer0_outputs(6868) <= b;
    layer0_outputs(6869) <= b;
    layer0_outputs(6870) <= a or b;
    layer0_outputs(6871) <= a xor b;
    layer0_outputs(6872) <= b and not a;
    layer0_outputs(6873) <= a or b;
    layer0_outputs(6874) <= not (a xor b);
    layer0_outputs(6875) <= not a;
    layer0_outputs(6876) <= a xor b;
    layer0_outputs(6877) <= b and not a;
    layer0_outputs(6878) <= not (a xor b);
    layer0_outputs(6879) <= a xor b;
    layer0_outputs(6880) <= not b or a;
    layer0_outputs(6881) <= a xor b;
    layer0_outputs(6882) <= not (a or b);
    layer0_outputs(6883) <= not b;
    layer0_outputs(6884) <= not a or b;
    layer0_outputs(6885) <= '0';
    layer0_outputs(6886) <= not b or a;
    layer0_outputs(6887) <= a xor b;
    layer0_outputs(6888) <= not b;
    layer0_outputs(6889) <= not (a xor b);
    layer0_outputs(6890) <= not b;
    layer0_outputs(6891) <= not (a or b);
    layer0_outputs(6892) <= not (a or b);
    layer0_outputs(6893) <= not (a and b);
    layer0_outputs(6894) <= not a or b;
    layer0_outputs(6895) <= a;
    layer0_outputs(6896) <= '1';
    layer0_outputs(6897) <= not (a or b);
    layer0_outputs(6898) <= a xor b;
    layer0_outputs(6899) <= not (a xor b);
    layer0_outputs(6900) <= not a or b;
    layer0_outputs(6901) <= not (a xor b);
    layer0_outputs(6902) <= a or b;
    layer0_outputs(6903) <= not (a xor b);
    layer0_outputs(6904) <= b;
    layer0_outputs(6905) <= not a or b;
    layer0_outputs(6906) <= not b;
    layer0_outputs(6907) <= not (a xor b);
    layer0_outputs(6908) <= not (a or b);
    layer0_outputs(6909) <= a;
    layer0_outputs(6910) <= not (a xor b);
    layer0_outputs(6911) <= not (a or b);
    layer0_outputs(6912) <= not (a or b);
    layer0_outputs(6913) <= not (a xor b);
    layer0_outputs(6914) <= a and not b;
    layer0_outputs(6915) <= not a or b;
    layer0_outputs(6916) <= not b;
    layer0_outputs(6917) <= a xor b;
    layer0_outputs(6918) <= not (a or b);
    layer0_outputs(6919) <= not a or b;
    layer0_outputs(6920) <= a;
    layer0_outputs(6921) <= a and not b;
    layer0_outputs(6922) <= not (a or b);
    layer0_outputs(6923) <= not b or a;
    layer0_outputs(6924) <= not (a xor b);
    layer0_outputs(6925) <= not a or b;
    layer0_outputs(6926) <= a xor b;
    layer0_outputs(6927) <= a xor b;
    layer0_outputs(6928) <= a or b;
    layer0_outputs(6929) <= not (a xor b);
    layer0_outputs(6930) <= not b;
    layer0_outputs(6931) <= not (a or b);
    layer0_outputs(6932) <= a or b;
    layer0_outputs(6933) <= a xor b;
    layer0_outputs(6934) <= not (a or b);
    layer0_outputs(6935) <= a xor b;
    layer0_outputs(6936) <= '0';
    layer0_outputs(6937) <= b and not a;
    layer0_outputs(6938) <= not a;
    layer0_outputs(6939) <= not a or b;
    layer0_outputs(6940) <= a and b;
    layer0_outputs(6941) <= '0';
    layer0_outputs(6942) <= not (a xor b);
    layer0_outputs(6943) <= a or b;
    layer0_outputs(6944) <= not b or a;
    layer0_outputs(6945) <= not a;
    layer0_outputs(6946) <= b;
    layer0_outputs(6947) <= not a;
    layer0_outputs(6948) <= not (a or b);
    layer0_outputs(6949) <= b;
    layer0_outputs(6950) <= b and not a;
    layer0_outputs(6951) <= a or b;
    layer0_outputs(6952) <= not b or a;
    layer0_outputs(6953) <= not a;
    layer0_outputs(6954) <= not b or a;
    layer0_outputs(6955) <= a or b;
    layer0_outputs(6956) <= not b;
    layer0_outputs(6957) <= not b;
    layer0_outputs(6958) <= a or b;
    layer0_outputs(6959) <= a or b;
    layer0_outputs(6960) <= a xor b;
    layer0_outputs(6961) <= a xor b;
    layer0_outputs(6962) <= b and not a;
    layer0_outputs(6963) <= not (a or b);
    layer0_outputs(6964) <= not a or b;
    layer0_outputs(6965) <= not a or b;
    layer0_outputs(6966) <= not a;
    layer0_outputs(6967) <= not (a xor b);
    layer0_outputs(6968) <= a;
    layer0_outputs(6969) <= a xor b;
    layer0_outputs(6970) <= not b;
    layer0_outputs(6971) <= not b or a;
    layer0_outputs(6972) <= not (a xor b);
    layer0_outputs(6973) <= a;
    layer0_outputs(6974) <= not a or b;
    layer0_outputs(6975) <= not (a or b);
    layer0_outputs(6976) <= a;
    layer0_outputs(6977) <= a and b;
    layer0_outputs(6978) <= b and not a;
    layer0_outputs(6979) <= a xor b;
    layer0_outputs(6980) <= a or b;
    layer0_outputs(6981) <= a or b;
    layer0_outputs(6982) <= a xor b;
    layer0_outputs(6983) <= not (a or b);
    layer0_outputs(6984) <= a and not b;
    layer0_outputs(6985) <= not (a xor b);
    layer0_outputs(6986) <= '1';
    layer0_outputs(6987) <= not (a or b);
    layer0_outputs(6988) <= not (a xor b);
    layer0_outputs(6989) <= a or b;
    layer0_outputs(6990) <= not a or b;
    layer0_outputs(6991) <= not (a or b);
    layer0_outputs(6992) <= b and not a;
    layer0_outputs(6993) <= not a;
    layer0_outputs(6994) <= a or b;
    layer0_outputs(6995) <= b;
    layer0_outputs(6996) <= a or b;
    layer0_outputs(6997) <= not (a or b);
    layer0_outputs(6998) <= '0';
    layer0_outputs(6999) <= not a or b;
    layer0_outputs(7000) <= a;
    layer0_outputs(7001) <= not b or a;
    layer0_outputs(7002) <= not b or a;
    layer0_outputs(7003) <= not (a or b);
    layer0_outputs(7004) <= '0';
    layer0_outputs(7005) <= not (a and b);
    layer0_outputs(7006) <= a;
    layer0_outputs(7007) <= a or b;
    layer0_outputs(7008) <= a or b;
    layer0_outputs(7009) <= not (a or b);
    layer0_outputs(7010) <= not b;
    layer0_outputs(7011) <= not (a or b);
    layer0_outputs(7012) <= not (a or b);
    layer0_outputs(7013) <= b and not a;
    layer0_outputs(7014) <= not (a xor b);
    layer0_outputs(7015) <= not (a xor b);
    layer0_outputs(7016) <= not (a or b);
    layer0_outputs(7017) <= a xor b;
    layer0_outputs(7018) <= a or b;
    layer0_outputs(7019) <= not (a xor b);
    layer0_outputs(7020) <= b and not a;
    layer0_outputs(7021) <= not (a or b);
    layer0_outputs(7022) <= not (a and b);
    layer0_outputs(7023) <= b;
    layer0_outputs(7024) <= a or b;
    layer0_outputs(7025) <= not b;
    layer0_outputs(7026) <= not (a or b);
    layer0_outputs(7027) <= a and not b;
    layer0_outputs(7028) <= b and not a;
    layer0_outputs(7029) <= b and not a;
    layer0_outputs(7030) <= not b;
    layer0_outputs(7031) <= a or b;
    layer0_outputs(7032) <= not (a or b);
    layer0_outputs(7033) <= not b;
    layer0_outputs(7034) <= a xor b;
    layer0_outputs(7035) <= not a or b;
    layer0_outputs(7036) <= b;
    layer0_outputs(7037) <= not b;
    layer0_outputs(7038) <= a and not b;
    layer0_outputs(7039) <= a and not b;
    layer0_outputs(7040) <= b and not a;
    layer0_outputs(7041) <= not (a xor b);
    layer0_outputs(7042) <= not b;
    layer0_outputs(7043) <= a or b;
    layer0_outputs(7044) <= a xor b;
    layer0_outputs(7045) <= not b;
    layer0_outputs(7046) <= not (a xor b);
    layer0_outputs(7047) <= a or b;
    layer0_outputs(7048) <= a or b;
    layer0_outputs(7049) <= a or b;
    layer0_outputs(7050) <= a or b;
    layer0_outputs(7051) <= not a;
    layer0_outputs(7052) <= b;
    layer0_outputs(7053) <= not (a xor b);
    layer0_outputs(7054) <= not (a or b);
    layer0_outputs(7055) <= not a or b;
    layer0_outputs(7056) <= '0';
    layer0_outputs(7057) <= b;
    layer0_outputs(7058) <= a or b;
    layer0_outputs(7059) <= not (a or b);
    layer0_outputs(7060) <= not a;
    layer0_outputs(7061) <= a or b;
    layer0_outputs(7062) <= not b;
    layer0_outputs(7063) <= not b or a;
    layer0_outputs(7064) <= not (a xor b);
    layer0_outputs(7065) <= '0';
    layer0_outputs(7066) <= not (a xor b);
    layer0_outputs(7067) <= b;
    layer0_outputs(7068) <= not a or b;
    layer0_outputs(7069) <= b and not a;
    layer0_outputs(7070) <= not (a xor b);
    layer0_outputs(7071) <= not b;
    layer0_outputs(7072) <= not (a and b);
    layer0_outputs(7073) <= not (a or b);
    layer0_outputs(7074) <= not (a or b);
    layer0_outputs(7075) <= not (a xor b);
    layer0_outputs(7076) <= b and not a;
    layer0_outputs(7077) <= not (a xor b);
    layer0_outputs(7078) <= not a or b;
    layer0_outputs(7079) <= a or b;
    layer0_outputs(7080) <= not (a xor b);
    layer0_outputs(7081) <= a xor b;
    layer0_outputs(7082) <= b;
    layer0_outputs(7083) <= a or b;
    layer0_outputs(7084) <= '1';
    layer0_outputs(7085) <= b and not a;
    layer0_outputs(7086) <= a or b;
    layer0_outputs(7087) <= a and not b;
    layer0_outputs(7088) <= not a or b;
    layer0_outputs(7089) <= b and not a;
    layer0_outputs(7090) <= a or b;
    layer0_outputs(7091) <= '1';
    layer0_outputs(7092) <= not (a xor b);
    layer0_outputs(7093) <= a and not b;
    layer0_outputs(7094) <= not b or a;
    layer0_outputs(7095) <= a or b;
    layer0_outputs(7096) <= '1';
    layer0_outputs(7097) <= b;
    layer0_outputs(7098) <= a xor b;
    layer0_outputs(7099) <= a or b;
    layer0_outputs(7100) <= a and not b;
    layer0_outputs(7101) <= a or b;
    layer0_outputs(7102) <= '1';
    layer0_outputs(7103) <= not b;
    layer0_outputs(7104) <= b and not a;
    layer0_outputs(7105) <= a xor b;
    layer0_outputs(7106) <= a;
    layer0_outputs(7107) <= not (a or b);
    layer0_outputs(7108) <= not a;
    layer0_outputs(7109) <= not b;
    layer0_outputs(7110) <= a or b;
    layer0_outputs(7111) <= b and not a;
    layer0_outputs(7112) <= not (a or b);
    layer0_outputs(7113) <= not b or a;
    layer0_outputs(7114) <= a or b;
    layer0_outputs(7115) <= a;
    layer0_outputs(7116) <= a;
    layer0_outputs(7117) <= not a;
    layer0_outputs(7118) <= not b or a;
    layer0_outputs(7119) <= not a;
    layer0_outputs(7120) <= b;
    layer0_outputs(7121) <= not a;
    layer0_outputs(7122) <= b;
    layer0_outputs(7123) <= a xor b;
    layer0_outputs(7124) <= not (a xor b);
    layer0_outputs(7125) <= not b;
    layer0_outputs(7126) <= b and not a;
    layer0_outputs(7127) <= not a or b;
    layer0_outputs(7128) <= a or b;
    layer0_outputs(7129) <= not b;
    layer0_outputs(7130) <= not (a or b);
    layer0_outputs(7131) <= not (a or b);
    layer0_outputs(7132) <= a or b;
    layer0_outputs(7133) <= a or b;
    layer0_outputs(7134) <= a;
    layer0_outputs(7135) <= not (a xor b);
    layer0_outputs(7136) <= not (a or b);
    layer0_outputs(7137) <= b and not a;
    layer0_outputs(7138) <= not b or a;
    layer0_outputs(7139) <= b;
    layer0_outputs(7140) <= not (a or b);
    layer0_outputs(7141) <= a or b;
    layer0_outputs(7142) <= not a;
    layer0_outputs(7143) <= a and not b;
    layer0_outputs(7144) <= not (a xor b);
    layer0_outputs(7145) <= not (a or b);
    layer0_outputs(7146) <= not b;
    layer0_outputs(7147) <= a and not b;
    layer0_outputs(7148) <= not a or b;
    layer0_outputs(7149) <= a xor b;
    layer0_outputs(7150) <= not (a xor b);
    layer0_outputs(7151) <= not a or b;
    layer0_outputs(7152) <= not (a or b);
    layer0_outputs(7153) <= not b or a;
    layer0_outputs(7154) <= a xor b;
    layer0_outputs(7155) <= not (a or b);
    layer0_outputs(7156) <= a or b;
    layer0_outputs(7157) <= not (a or b);
    layer0_outputs(7158) <= not a;
    layer0_outputs(7159) <= not (a or b);
    layer0_outputs(7160) <= b;
    layer0_outputs(7161) <= a or b;
    layer0_outputs(7162) <= a;
    layer0_outputs(7163) <= a and not b;
    layer0_outputs(7164) <= not a;
    layer0_outputs(7165) <= not b;
    layer0_outputs(7166) <= not b;
    layer0_outputs(7167) <= a or b;
    layer0_outputs(7168) <= not b or a;
    layer0_outputs(7169) <= a or b;
    layer0_outputs(7170) <= a and not b;
    layer0_outputs(7171) <= not b;
    layer0_outputs(7172) <= not a;
    layer0_outputs(7173) <= not (a or b);
    layer0_outputs(7174) <= not a or b;
    layer0_outputs(7175) <= not (a or b);
    layer0_outputs(7176) <= not b;
    layer0_outputs(7177) <= a or b;
    layer0_outputs(7178) <= not a or b;
    layer0_outputs(7179) <= a and b;
    layer0_outputs(7180) <= '1';
    layer0_outputs(7181) <= not b;
    layer0_outputs(7182) <= not (a or b);
    layer0_outputs(7183) <= a or b;
    layer0_outputs(7184) <= a and not b;
    layer0_outputs(7185) <= not a or b;
    layer0_outputs(7186) <= not b;
    layer0_outputs(7187) <= not (a xor b);
    layer0_outputs(7188) <= a;
    layer0_outputs(7189) <= not (a xor b);
    layer0_outputs(7190) <= a and not b;
    layer0_outputs(7191) <= '0';
    layer0_outputs(7192) <= a and not b;
    layer0_outputs(7193) <= not a or b;
    layer0_outputs(7194) <= not (a or b);
    layer0_outputs(7195) <= not b;
    layer0_outputs(7196) <= not (a or b);
    layer0_outputs(7197) <= b and not a;
    layer0_outputs(7198) <= b and not a;
    layer0_outputs(7199) <= b;
    layer0_outputs(7200) <= not (a xor b);
    layer0_outputs(7201) <= a xor b;
    layer0_outputs(7202) <= a or b;
    layer0_outputs(7203) <= not (a or b);
    layer0_outputs(7204) <= a xor b;
    layer0_outputs(7205) <= not (a and b);
    layer0_outputs(7206) <= not b or a;
    layer0_outputs(7207) <= not a or b;
    layer0_outputs(7208) <= a xor b;
    layer0_outputs(7209) <= b;
    layer0_outputs(7210) <= not (a xor b);
    layer0_outputs(7211) <= b;
    layer0_outputs(7212) <= not (a or b);
    layer0_outputs(7213) <= a;
    layer0_outputs(7214) <= not b;
    layer0_outputs(7215) <= b and not a;
    layer0_outputs(7216) <= a or b;
    layer0_outputs(7217) <= a;
    layer0_outputs(7218) <= a and not b;
    layer0_outputs(7219) <= not a or b;
    layer0_outputs(7220) <= a xor b;
    layer0_outputs(7221) <= not (a or b);
    layer0_outputs(7222) <= b;
    layer0_outputs(7223) <= a;
    layer0_outputs(7224) <= not (a or b);
    layer0_outputs(7225) <= not b or a;
    layer0_outputs(7226) <= a or b;
    layer0_outputs(7227) <= not (a or b);
    layer0_outputs(7228) <= not (a xor b);
    layer0_outputs(7229) <= not (a xor b);
    layer0_outputs(7230) <= a or b;
    layer0_outputs(7231) <= b;
    layer0_outputs(7232) <= a and not b;
    layer0_outputs(7233) <= not (a or b);
    layer0_outputs(7234) <= a or b;
    layer0_outputs(7235) <= a;
    layer0_outputs(7236) <= not (a xor b);
    layer0_outputs(7237) <= a;
    layer0_outputs(7238) <= a and not b;
    layer0_outputs(7239) <= not (a or b);
    layer0_outputs(7240) <= not b;
    layer0_outputs(7241) <= a or b;
    layer0_outputs(7242) <= not (a or b);
    layer0_outputs(7243) <= not (a or b);
    layer0_outputs(7244) <= a or b;
    layer0_outputs(7245) <= b and not a;
    layer0_outputs(7246) <= not (a xor b);
    layer0_outputs(7247) <= a or b;
    layer0_outputs(7248) <= not (a and b);
    layer0_outputs(7249) <= not (a xor b);
    layer0_outputs(7250) <= not a;
    layer0_outputs(7251) <= a and not b;
    layer0_outputs(7252) <= not (a xor b);
    layer0_outputs(7253) <= b;
    layer0_outputs(7254) <= not (a and b);
    layer0_outputs(7255) <= not (a xor b);
    layer0_outputs(7256) <= '0';
    layer0_outputs(7257) <= a;
    layer0_outputs(7258) <= a or b;
    layer0_outputs(7259) <= not (a or b);
    layer0_outputs(7260) <= b and not a;
    layer0_outputs(7261) <= a;
    layer0_outputs(7262) <= b;
    layer0_outputs(7263) <= a;
    layer0_outputs(7264) <= not a;
    layer0_outputs(7265) <= not (a xor b);
    layer0_outputs(7266) <= a or b;
    layer0_outputs(7267) <= a;
    layer0_outputs(7268) <= not b;
    layer0_outputs(7269) <= not a;
    layer0_outputs(7270) <= not b;
    layer0_outputs(7271) <= not (a or b);
    layer0_outputs(7272) <= a or b;
    layer0_outputs(7273) <= not (a or b);
    layer0_outputs(7274) <= a or b;
    layer0_outputs(7275) <= a and b;
    layer0_outputs(7276) <= not (a or b);
    layer0_outputs(7277) <= not b;
    layer0_outputs(7278) <= not (a or b);
    layer0_outputs(7279) <= not (a and b);
    layer0_outputs(7280) <= not (a xor b);
    layer0_outputs(7281) <= not b;
    layer0_outputs(7282) <= a;
    layer0_outputs(7283) <= not a;
    layer0_outputs(7284) <= not a or b;
    layer0_outputs(7285) <= not b;
    layer0_outputs(7286) <= a;
    layer0_outputs(7287) <= not (a or b);
    layer0_outputs(7288) <= a xor b;
    layer0_outputs(7289) <= not (a xor b);
    layer0_outputs(7290) <= not (a xor b);
    layer0_outputs(7291) <= not b;
    layer0_outputs(7292) <= not b or a;
    layer0_outputs(7293) <= not (a or b);
    layer0_outputs(7294) <= not a;
    layer0_outputs(7295) <= b and not a;
    layer0_outputs(7296) <= a xor b;
    layer0_outputs(7297) <= b;
    layer0_outputs(7298) <= not (a or b);
    layer0_outputs(7299) <= not a;
    layer0_outputs(7300) <= not (a and b);
    layer0_outputs(7301) <= a or b;
    layer0_outputs(7302) <= a or b;
    layer0_outputs(7303) <= not (a or b);
    layer0_outputs(7304) <= not (a or b);
    layer0_outputs(7305) <= not b or a;
    layer0_outputs(7306) <= a or b;
    layer0_outputs(7307) <= a and not b;
    layer0_outputs(7308) <= not b;
    layer0_outputs(7309) <= not (a xor b);
    layer0_outputs(7310) <= a;
    layer0_outputs(7311) <= not a or b;
    layer0_outputs(7312) <= b and not a;
    layer0_outputs(7313) <= not a;
    layer0_outputs(7314) <= '1';
    layer0_outputs(7315) <= a;
    layer0_outputs(7316) <= not (a or b);
    layer0_outputs(7317) <= not (a xor b);
    layer0_outputs(7318) <= b;
    layer0_outputs(7319) <= a;
    layer0_outputs(7320) <= not (a xor b);
    layer0_outputs(7321) <= not b or a;
    layer0_outputs(7322) <= not a or b;
    layer0_outputs(7323) <= not a or b;
    layer0_outputs(7324) <= not b;
    layer0_outputs(7325) <= b;
    layer0_outputs(7326) <= a xor b;
    layer0_outputs(7327) <= not (a or b);
    layer0_outputs(7328) <= not b;
    layer0_outputs(7329) <= not (a xor b);
    layer0_outputs(7330) <= not (a or b);
    layer0_outputs(7331) <= not (a or b);
    layer0_outputs(7332) <= not (a or b);
    layer0_outputs(7333) <= a and not b;
    layer0_outputs(7334) <= not (a or b);
    layer0_outputs(7335) <= not b;
    layer0_outputs(7336) <= b and not a;
    layer0_outputs(7337) <= a;
    layer0_outputs(7338) <= not (a xor b);
    layer0_outputs(7339) <= a and b;
    layer0_outputs(7340) <= b and not a;
    layer0_outputs(7341) <= not (a or b);
    layer0_outputs(7342) <= not a;
    layer0_outputs(7343) <= a;
    layer0_outputs(7344) <= a or b;
    layer0_outputs(7345) <= b and not a;
    layer0_outputs(7346) <= not (a xor b);
    layer0_outputs(7347) <= '1';
    layer0_outputs(7348) <= '0';
    layer0_outputs(7349) <= not (a or b);
    layer0_outputs(7350) <= a or b;
    layer0_outputs(7351) <= a;
    layer0_outputs(7352) <= not b;
    layer0_outputs(7353) <= a or b;
    layer0_outputs(7354) <= b;
    layer0_outputs(7355) <= a or b;
    layer0_outputs(7356) <= not (a xor b);
    layer0_outputs(7357) <= a and not b;
    layer0_outputs(7358) <= not a;
    layer0_outputs(7359) <= b and not a;
    layer0_outputs(7360) <= not a or b;
    layer0_outputs(7361) <= a xor b;
    layer0_outputs(7362) <= not (a xor b);
    layer0_outputs(7363) <= b;
    layer0_outputs(7364) <= not (a or b);
    layer0_outputs(7365) <= a xor b;
    layer0_outputs(7366) <= not a;
    layer0_outputs(7367) <= not a;
    layer0_outputs(7368) <= not a or b;
    layer0_outputs(7369) <= not (a xor b);
    layer0_outputs(7370) <= b and not a;
    layer0_outputs(7371) <= a or b;
    layer0_outputs(7372) <= not (a xor b);
    layer0_outputs(7373) <= a or b;
    layer0_outputs(7374) <= a or b;
    layer0_outputs(7375) <= a and not b;
    layer0_outputs(7376) <= not a;
    layer0_outputs(7377) <= a or b;
    layer0_outputs(7378) <= b and not a;
    layer0_outputs(7379) <= not a or b;
    layer0_outputs(7380) <= not (a or b);
    layer0_outputs(7381) <= b and not a;
    layer0_outputs(7382) <= not b;
    layer0_outputs(7383) <= a xor b;
    layer0_outputs(7384) <= a xor b;
    layer0_outputs(7385) <= '0';
    layer0_outputs(7386) <= not (a or b);
    layer0_outputs(7387) <= a or b;
    layer0_outputs(7388) <= a and not b;
    layer0_outputs(7389) <= a and not b;
    layer0_outputs(7390) <= a or b;
    layer0_outputs(7391) <= not a or b;
    layer0_outputs(7392) <= not (a xor b);
    layer0_outputs(7393) <= not a or b;
    layer0_outputs(7394) <= not b or a;
    layer0_outputs(7395) <= not (a xor b);
    layer0_outputs(7396) <= not (a xor b);
    layer0_outputs(7397) <= not (a or b);
    layer0_outputs(7398) <= not b or a;
    layer0_outputs(7399) <= b;
    layer0_outputs(7400) <= not (a and b);
    layer0_outputs(7401) <= a or b;
    layer0_outputs(7402) <= not a or b;
    layer0_outputs(7403) <= not (a or b);
    layer0_outputs(7404) <= a or b;
    layer0_outputs(7405) <= a or b;
    layer0_outputs(7406) <= a;
    layer0_outputs(7407) <= a xor b;
    layer0_outputs(7408) <= a xor b;
    layer0_outputs(7409) <= a or b;
    layer0_outputs(7410) <= a or b;
    layer0_outputs(7411) <= not (a or b);
    layer0_outputs(7412) <= not b;
    layer0_outputs(7413) <= a;
    layer0_outputs(7414) <= not a;
    layer0_outputs(7415) <= not (a xor b);
    layer0_outputs(7416) <= not (a xor b);
    layer0_outputs(7417) <= not b;
    layer0_outputs(7418) <= a or b;
    layer0_outputs(7419) <= not (a xor b);
    layer0_outputs(7420) <= a or b;
    layer0_outputs(7421) <= a;
    layer0_outputs(7422) <= a and not b;
    layer0_outputs(7423) <= not (a xor b);
    layer0_outputs(7424) <= not (a or b);
    layer0_outputs(7425) <= not b or a;
    layer0_outputs(7426) <= b;
    layer0_outputs(7427) <= not b;
    layer0_outputs(7428) <= b;
    layer0_outputs(7429) <= not a or b;
    layer0_outputs(7430) <= a xor b;
    layer0_outputs(7431) <= not (a xor b);
    layer0_outputs(7432) <= not (a or b);
    layer0_outputs(7433) <= not a or b;
    layer0_outputs(7434) <= a and b;
    layer0_outputs(7435) <= not (a xor b);
    layer0_outputs(7436) <= a xor b;
    layer0_outputs(7437) <= not (a xor b);
    layer0_outputs(7438) <= b;
    layer0_outputs(7439) <= a and not b;
    layer0_outputs(7440) <= not (a or b);
    layer0_outputs(7441) <= a xor b;
    layer0_outputs(7442) <= not (a or b);
    layer0_outputs(7443) <= a or b;
    layer0_outputs(7444) <= not b;
    layer0_outputs(7445) <= a and b;
    layer0_outputs(7446) <= not a;
    layer0_outputs(7447) <= not b;
    layer0_outputs(7448) <= not (a and b);
    layer0_outputs(7449) <= a and b;
    layer0_outputs(7450) <= a xor b;
    layer0_outputs(7451) <= not b;
    layer0_outputs(7452) <= a xor b;
    layer0_outputs(7453) <= not b;
    layer0_outputs(7454) <= '0';
    layer0_outputs(7455) <= b and not a;
    layer0_outputs(7456) <= not (a xor b);
    layer0_outputs(7457) <= b and not a;
    layer0_outputs(7458) <= b and not a;
    layer0_outputs(7459) <= '1';
    layer0_outputs(7460) <= not (a and b);
    layer0_outputs(7461) <= not (a or b);
    layer0_outputs(7462) <= not (a or b);
    layer0_outputs(7463) <= a and b;
    layer0_outputs(7464) <= not a or b;
    layer0_outputs(7465) <= not (a xor b);
    layer0_outputs(7466) <= a xor b;
    layer0_outputs(7467) <= b;
    layer0_outputs(7468) <= a and not b;
    layer0_outputs(7469) <= not a or b;
    layer0_outputs(7470) <= b and not a;
    layer0_outputs(7471) <= not (a or b);
    layer0_outputs(7472) <= not a;
    layer0_outputs(7473) <= not (a or b);
    layer0_outputs(7474) <= not (a xor b);
    layer0_outputs(7475) <= a and b;
    layer0_outputs(7476) <= not b;
    layer0_outputs(7477) <= not a or b;
    layer0_outputs(7478) <= not (a or b);
    layer0_outputs(7479) <= not (a xor b);
    layer0_outputs(7480) <= not b or a;
    layer0_outputs(7481) <= a;
    layer0_outputs(7482) <= a;
    layer0_outputs(7483) <= b;
    layer0_outputs(7484) <= not (a xor b);
    layer0_outputs(7485) <= b and not a;
    layer0_outputs(7486) <= a xor b;
    layer0_outputs(7487) <= not a or b;
    layer0_outputs(7488) <= not b or a;
    layer0_outputs(7489) <= a xor b;
    layer0_outputs(7490) <= b;
    layer0_outputs(7491) <= a xor b;
    layer0_outputs(7492) <= not (a xor b);
    layer0_outputs(7493) <= not (a xor b);
    layer0_outputs(7494) <= not (a and b);
    layer0_outputs(7495) <= b and not a;
    layer0_outputs(7496) <= b;
    layer0_outputs(7497) <= not a or b;
    layer0_outputs(7498) <= b and not a;
    layer0_outputs(7499) <= not a or b;
    layer0_outputs(7500) <= not (a xor b);
    layer0_outputs(7501) <= not (a and b);
    layer0_outputs(7502) <= a xor b;
    layer0_outputs(7503) <= a and not b;
    layer0_outputs(7504) <= a or b;
    layer0_outputs(7505) <= a or b;
    layer0_outputs(7506) <= a or b;
    layer0_outputs(7507) <= not (a xor b);
    layer0_outputs(7508) <= not a or b;
    layer0_outputs(7509) <= not (a xor b);
    layer0_outputs(7510) <= not (a xor b);
    layer0_outputs(7511) <= a and not b;
    layer0_outputs(7512) <= a xor b;
    layer0_outputs(7513) <= b;
    layer0_outputs(7514) <= a or b;
    layer0_outputs(7515) <= not a;
    layer0_outputs(7516) <= a;
    layer0_outputs(7517) <= not a or b;
    layer0_outputs(7518) <= a and b;
    layer0_outputs(7519) <= not b;
    layer0_outputs(7520) <= a;
    layer0_outputs(7521) <= a or b;
    layer0_outputs(7522) <= b and not a;
    layer0_outputs(7523) <= not (a xor b);
    layer0_outputs(7524) <= not a;
    layer0_outputs(7525) <= a;
    layer0_outputs(7526) <= a or b;
    layer0_outputs(7527) <= not a or b;
    layer0_outputs(7528) <= b;
    layer0_outputs(7529) <= a or b;
    layer0_outputs(7530) <= not b or a;
    layer0_outputs(7531) <= a xor b;
    layer0_outputs(7532) <= a;
    layer0_outputs(7533) <= a or b;
    layer0_outputs(7534) <= not (a xor b);
    layer0_outputs(7535) <= not (a or b);
    layer0_outputs(7536) <= a and not b;
    layer0_outputs(7537) <= a or b;
    layer0_outputs(7538) <= a and b;
    layer0_outputs(7539) <= '0';
    layer0_outputs(7540) <= a;
    layer0_outputs(7541) <= not (a xor b);
    layer0_outputs(7542) <= not b or a;
    layer0_outputs(7543) <= not a or b;
    layer0_outputs(7544) <= not a or b;
    layer0_outputs(7545) <= a and b;
    layer0_outputs(7546) <= not b or a;
    layer0_outputs(7547) <= not b;
    layer0_outputs(7548) <= '1';
    layer0_outputs(7549) <= a;
    layer0_outputs(7550) <= not (a or b);
    layer0_outputs(7551) <= not b;
    layer0_outputs(7552) <= a xor b;
    layer0_outputs(7553) <= not b;
    layer0_outputs(7554) <= not (a or b);
    layer0_outputs(7555) <= not a or b;
    layer0_outputs(7556) <= a xor b;
    layer0_outputs(7557) <= not a;
    layer0_outputs(7558) <= a or b;
    layer0_outputs(7559) <= a and not b;
    layer0_outputs(7560) <= not b;
    layer0_outputs(7561) <= b and not a;
    layer0_outputs(7562) <= b;
    layer0_outputs(7563) <= not a;
    layer0_outputs(7564) <= a;
    layer0_outputs(7565) <= a or b;
    layer0_outputs(7566) <= not a or b;
    layer0_outputs(7567) <= a and not b;
    layer0_outputs(7568) <= a xor b;
    layer0_outputs(7569) <= not a or b;
    layer0_outputs(7570) <= a;
    layer0_outputs(7571) <= not b;
    layer0_outputs(7572) <= not (a or b);
    layer0_outputs(7573) <= a xor b;
    layer0_outputs(7574) <= not a;
    layer0_outputs(7575) <= not b;
    layer0_outputs(7576) <= not b or a;
    layer0_outputs(7577) <= not (a xor b);
    layer0_outputs(7578) <= a or b;
    layer0_outputs(7579) <= a or b;
    layer0_outputs(7580) <= a xor b;
    layer0_outputs(7581) <= a or b;
    layer0_outputs(7582) <= not (a or b);
    layer0_outputs(7583) <= a or b;
    layer0_outputs(7584) <= a and not b;
    layer0_outputs(7585) <= not a;
    layer0_outputs(7586) <= a or b;
    layer0_outputs(7587) <= a or b;
    layer0_outputs(7588) <= b;
    layer0_outputs(7589) <= a and not b;
    layer0_outputs(7590) <= not b;
    layer0_outputs(7591) <= a;
    layer0_outputs(7592) <= not b;
    layer0_outputs(7593) <= not (a xor b);
    layer0_outputs(7594) <= a or b;
    layer0_outputs(7595) <= not (a xor b);
    layer0_outputs(7596) <= not a;
    layer0_outputs(7597) <= not a or b;
    layer0_outputs(7598) <= not (a or b);
    layer0_outputs(7599) <= not (a xor b);
    layer0_outputs(7600) <= b and not a;
    layer0_outputs(7601) <= not (a xor b);
    layer0_outputs(7602) <= b;
    layer0_outputs(7603) <= not a;
    layer0_outputs(7604) <= not a;
    layer0_outputs(7605) <= not a or b;
    layer0_outputs(7606) <= not b;
    layer0_outputs(7607) <= a or b;
    layer0_outputs(7608) <= not a;
    layer0_outputs(7609) <= not a or b;
    layer0_outputs(7610) <= not (a or b);
    layer0_outputs(7611) <= b and not a;
    layer0_outputs(7612) <= not a or b;
    layer0_outputs(7613) <= '0';
    layer0_outputs(7614) <= a and b;
    layer0_outputs(7615) <= not (a or b);
    layer0_outputs(7616) <= not (a xor b);
    layer0_outputs(7617) <= not a;
    layer0_outputs(7618) <= not b;
    layer0_outputs(7619) <= a and b;
    layer0_outputs(7620) <= a or b;
    layer0_outputs(7621) <= not b or a;
    layer0_outputs(7622) <= not a or b;
    layer0_outputs(7623) <= not b;
    layer0_outputs(7624) <= a and not b;
    layer0_outputs(7625) <= a xor b;
    layer0_outputs(7626) <= a xor b;
    layer0_outputs(7627) <= '1';
    layer0_outputs(7628) <= a or b;
    layer0_outputs(7629) <= a and not b;
    layer0_outputs(7630) <= b;
    layer0_outputs(7631) <= not a;
    layer0_outputs(7632) <= not (a and b);
    layer0_outputs(7633) <= not b or a;
    layer0_outputs(7634) <= '1';
    layer0_outputs(7635) <= not (a or b);
    layer0_outputs(7636) <= not (a xor b);
    layer0_outputs(7637) <= not a;
    layer0_outputs(7638) <= not (a xor b);
    layer0_outputs(7639) <= not (a or b);
    layer0_outputs(7640) <= not (a or b);
    layer0_outputs(7641) <= not (a or b);
    layer0_outputs(7642) <= not (a or b);
    layer0_outputs(7643) <= a xor b;
    layer0_outputs(7644) <= a xor b;
    layer0_outputs(7645) <= not (a xor b);
    layer0_outputs(7646) <= not (a or b);
    layer0_outputs(7647) <= not (a or b);
    layer0_outputs(7648) <= b and not a;
    layer0_outputs(7649) <= not b;
    layer0_outputs(7650) <= not b or a;
    layer0_outputs(7651) <= a and b;
    layer0_outputs(7652) <= a xor b;
    layer0_outputs(7653) <= not a or b;
    layer0_outputs(7654) <= not (a or b);
    layer0_outputs(7655) <= b;
    layer0_outputs(7656) <= b and not a;
    layer0_outputs(7657) <= not (a or b);
    layer0_outputs(7658) <= not (a and b);
    layer0_outputs(7659) <= not b or a;
    layer0_outputs(7660) <= '0';
    layer0_outputs(7661) <= not (a xor b);
    layer0_outputs(7662) <= b and not a;
    layer0_outputs(7663) <= not (a xor b);
    layer0_outputs(7664) <= '0';
    layer0_outputs(7665) <= a or b;
    layer0_outputs(7666) <= '1';
    layer0_outputs(7667) <= not (a or b);
    layer0_outputs(7668) <= a or b;
    layer0_outputs(7669) <= a and b;
    layer0_outputs(7670) <= not a or b;
    layer0_outputs(7671) <= a xor b;
    layer0_outputs(7672) <= a or b;
    layer0_outputs(7673) <= not (a or b);
    layer0_outputs(7674) <= not (a or b);
    layer0_outputs(7675) <= not a or b;
    layer0_outputs(7676) <= not (a xor b);
    layer0_outputs(7677) <= a or b;
    layer0_outputs(7678) <= b;
    layer0_outputs(7679) <= b and not a;
    layer0_outputs(7680) <= a and b;
    layer0_outputs(7681) <= b;
    layer0_outputs(7682) <= not a or b;
    layer0_outputs(7683) <= not (a xor b);
    layer0_outputs(7684) <= not a or b;
    layer0_outputs(7685) <= not b or a;
    layer0_outputs(7686) <= b;
    layer0_outputs(7687) <= a and not b;
    layer0_outputs(7688) <= not b or a;
    layer0_outputs(7689) <= not (a xor b);
    layer0_outputs(7690) <= not a or b;
    layer0_outputs(7691) <= not b or a;
    layer0_outputs(7692) <= not (a or b);
    layer0_outputs(7693) <= not (a or b);
    layer0_outputs(7694) <= a and b;
    layer0_outputs(7695) <= not (a and b);
    layer0_outputs(7696) <= b and not a;
    layer0_outputs(7697) <= not a;
    layer0_outputs(7698) <= b;
    layer0_outputs(7699) <= not (a xor b);
    layer0_outputs(7700) <= not b or a;
    layer0_outputs(7701) <= b;
    layer0_outputs(7702) <= b;
    layer0_outputs(7703) <= not (a or b);
    layer0_outputs(7704) <= '0';
    layer0_outputs(7705) <= not (a or b);
    layer0_outputs(7706) <= b and not a;
    layer0_outputs(7707) <= b and not a;
    layer0_outputs(7708) <= not b or a;
    layer0_outputs(7709) <= b;
    layer0_outputs(7710) <= not (a xor b);
    layer0_outputs(7711) <= a;
    layer0_outputs(7712) <= a xor b;
    layer0_outputs(7713) <= not (a or b);
    layer0_outputs(7714) <= not (a and b);
    layer0_outputs(7715) <= not a or b;
    layer0_outputs(7716) <= not a or b;
    layer0_outputs(7717) <= not (a xor b);
    layer0_outputs(7718) <= not a;
    layer0_outputs(7719) <= not (a and b);
    layer0_outputs(7720) <= not a or b;
    layer0_outputs(7721) <= a;
    layer0_outputs(7722) <= a and not b;
    layer0_outputs(7723) <= not (a and b);
    layer0_outputs(7724) <= not a;
    layer0_outputs(7725) <= not (a or b);
    layer0_outputs(7726) <= a xor b;
    layer0_outputs(7727) <= a and not b;
    layer0_outputs(7728) <= a or b;
    layer0_outputs(7729) <= b;
    layer0_outputs(7730) <= not a;
    layer0_outputs(7731) <= a xor b;
    layer0_outputs(7732) <= not (a or b);
    layer0_outputs(7733) <= not (a xor b);
    layer0_outputs(7734) <= not a;
    layer0_outputs(7735) <= not a or b;
    layer0_outputs(7736) <= not (a or b);
    layer0_outputs(7737) <= not (a or b);
    layer0_outputs(7738) <= not a or b;
    layer0_outputs(7739) <= a;
    layer0_outputs(7740) <= a;
    layer0_outputs(7741) <= a and not b;
    layer0_outputs(7742) <= not b;
    layer0_outputs(7743) <= b and not a;
    layer0_outputs(7744) <= not (a xor b);
    layer0_outputs(7745) <= not b;
    layer0_outputs(7746) <= not (a xor b);
    layer0_outputs(7747) <= not b;
    layer0_outputs(7748) <= not a or b;
    layer0_outputs(7749) <= a or b;
    layer0_outputs(7750) <= b;
    layer0_outputs(7751) <= a xor b;
    layer0_outputs(7752) <= b and not a;
    layer0_outputs(7753) <= not a or b;
    layer0_outputs(7754) <= not a or b;
    layer0_outputs(7755) <= a or b;
    layer0_outputs(7756) <= a and not b;
    layer0_outputs(7757) <= not a or b;
    layer0_outputs(7758) <= not (a xor b);
    layer0_outputs(7759) <= a and b;
    layer0_outputs(7760) <= not (a or b);
    layer0_outputs(7761) <= a or b;
    layer0_outputs(7762) <= not (a and b);
    layer0_outputs(7763) <= b;
    layer0_outputs(7764) <= not (a xor b);
    layer0_outputs(7765) <= not (a or b);
    layer0_outputs(7766) <= a and not b;
    layer0_outputs(7767) <= a or b;
    layer0_outputs(7768) <= a and not b;
    layer0_outputs(7769) <= b and not a;
    layer0_outputs(7770) <= a xor b;
    layer0_outputs(7771) <= a xor b;
    layer0_outputs(7772) <= a xor b;
    layer0_outputs(7773) <= a and not b;
    layer0_outputs(7774) <= a and b;
    layer0_outputs(7775) <= b and not a;
    layer0_outputs(7776) <= a and b;
    layer0_outputs(7777) <= not a;
    layer0_outputs(7778) <= not b or a;
    layer0_outputs(7779) <= a xor b;
    layer0_outputs(7780) <= a and b;
    layer0_outputs(7781) <= b and not a;
    layer0_outputs(7782) <= not a or b;
    layer0_outputs(7783) <= not (a or b);
    layer0_outputs(7784) <= a and b;
    layer0_outputs(7785) <= not a;
    layer0_outputs(7786) <= b;
    layer0_outputs(7787) <= not (a or b);
    layer0_outputs(7788) <= b and not a;
    layer0_outputs(7789) <= not (a or b);
    layer0_outputs(7790) <= a and not b;
    layer0_outputs(7791) <= not (a or b);
    layer0_outputs(7792) <= not b or a;
    layer0_outputs(7793) <= b and not a;
    layer0_outputs(7794) <= not (a or b);
    layer0_outputs(7795) <= b and not a;
    layer0_outputs(7796) <= a;
    layer0_outputs(7797) <= a or b;
    layer0_outputs(7798) <= not (a xor b);
    layer0_outputs(7799) <= not (a or b);
    layer0_outputs(7800) <= a xor b;
    layer0_outputs(7801) <= b;
    layer0_outputs(7802) <= a;
    layer0_outputs(7803) <= '1';
    layer0_outputs(7804) <= a or b;
    layer0_outputs(7805) <= b and not a;
    layer0_outputs(7806) <= b and not a;
    layer0_outputs(7807) <= not a or b;
    layer0_outputs(7808) <= not (a xor b);
    layer0_outputs(7809) <= a;
    layer0_outputs(7810) <= not a;
    layer0_outputs(7811) <= not (a or b);
    layer0_outputs(7812) <= not (a or b);
    layer0_outputs(7813) <= not b;
    layer0_outputs(7814) <= not (a or b);
    layer0_outputs(7815) <= a and b;
    layer0_outputs(7816) <= a or b;
    layer0_outputs(7817) <= a and not b;
    layer0_outputs(7818) <= a xor b;
    layer0_outputs(7819) <= a or b;
    layer0_outputs(7820) <= not a or b;
    layer0_outputs(7821) <= not (a or b);
    layer0_outputs(7822) <= not (a or b);
    layer0_outputs(7823) <= b and not a;
    layer0_outputs(7824) <= '1';
    layer0_outputs(7825) <= not b or a;
    layer0_outputs(7826) <= not (a or b);
    layer0_outputs(7827) <= a or b;
    layer0_outputs(7828) <= not (a or b);
    layer0_outputs(7829) <= b;
    layer0_outputs(7830) <= not b;
    layer0_outputs(7831) <= a or b;
    layer0_outputs(7832) <= not b;
    layer0_outputs(7833) <= not (a or b);
    layer0_outputs(7834) <= not a or b;
    layer0_outputs(7835) <= b and not a;
    layer0_outputs(7836) <= a and not b;
    layer0_outputs(7837) <= not a or b;
    layer0_outputs(7838) <= a or b;
    layer0_outputs(7839) <= a and not b;
    layer0_outputs(7840) <= a and not b;
    layer0_outputs(7841) <= not (a or b);
    layer0_outputs(7842) <= '1';
    layer0_outputs(7843) <= '0';
    layer0_outputs(7844) <= b;
    layer0_outputs(7845) <= not (a or b);
    layer0_outputs(7846) <= not a or b;
    layer0_outputs(7847) <= not a or b;
    layer0_outputs(7848) <= not a;
    layer0_outputs(7849) <= a and not b;
    layer0_outputs(7850) <= a;
    layer0_outputs(7851) <= a and not b;
    layer0_outputs(7852) <= a and not b;
    layer0_outputs(7853) <= not a or b;
    layer0_outputs(7854) <= not (a xor b);
    layer0_outputs(7855) <= not (a or b);
    layer0_outputs(7856) <= a or b;
    layer0_outputs(7857) <= a and not b;
    layer0_outputs(7858) <= not a or b;
    layer0_outputs(7859) <= a or b;
    layer0_outputs(7860) <= not a or b;
    layer0_outputs(7861) <= not a;
    layer0_outputs(7862) <= a xor b;
    layer0_outputs(7863) <= a xor b;
    layer0_outputs(7864) <= not a;
    layer0_outputs(7865) <= not b or a;
    layer0_outputs(7866) <= a or b;
    layer0_outputs(7867) <= a xor b;
    layer0_outputs(7868) <= b;
    layer0_outputs(7869) <= a and b;
    layer0_outputs(7870) <= b and not a;
    layer0_outputs(7871) <= not (a or b);
    layer0_outputs(7872) <= not (a xor b);
    layer0_outputs(7873) <= a and b;
    layer0_outputs(7874) <= not (a or b);
    layer0_outputs(7875) <= not a;
    layer0_outputs(7876) <= a and not b;
    layer0_outputs(7877) <= not a or b;
    layer0_outputs(7878) <= not a;
    layer0_outputs(7879) <= not a;
    layer0_outputs(7880) <= not (a or b);
    layer0_outputs(7881) <= not (a or b);
    layer0_outputs(7882) <= a and not b;
    layer0_outputs(7883) <= not a;
    layer0_outputs(7884) <= a xor b;
    layer0_outputs(7885) <= b and not a;
    layer0_outputs(7886) <= not b or a;
    layer0_outputs(7887) <= not b;
    layer0_outputs(7888) <= b;
    layer0_outputs(7889) <= not a or b;
    layer0_outputs(7890) <= a or b;
    layer0_outputs(7891) <= a and not b;
    layer0_outputs(7892) <= a or b;
    layer0_outputs(7893) <= not (a or b);
    layer0_outputs(7894) <= not a;
    layer0_outputs(7895) <= a or b;
    layer0_outputs(7896) <= not (a and b);
    layer0_outputs(7897) <= not b or a;
    layer0_outputs(7898) <= b and not a;
    layer0_outputs(7899) <= a or b;
    layer0_outputs(7900) <= not (a xor b);
    layer0_outputs(7901) <= not a or b;
    layer0_outputs(7902) <= not (a xor b);
    layer0_outputs(7903) <= not b;
    layer0_outputs(7904) <= a and not b;
    layer0_outputs(7905) <= '0';
    layer0_outputs(7906) <= '1';
    layer0_outputs(7907) <= a and b;
    layer0_outputs(7908) <= not b;
    layer0_outputs(7909) <= b and not a;
    layer0_outputs(7910) <= a and not b;
    layer0_outputs(7911) <= not (a and b);
    layer0_outputs(7912) <= not (a or b);
    layer0_outputs(7913) <= not b or a;
    layer0_outputs(7914) <= not a;
    layer0_outputs(7915) <= b;
    layer0_outputs(7916) <= not (a or b);
    layer0_outputs(7917) <= b and not a;
    layer0_outputs(7918) <= not a;
    layer0_outputs(7919) <= not b;
    layer0_outputs(7920) <= not b;
    layer0_outputs(7921) <= a xor b;
    layer0_outputs(7922) <= not b or a;
    layer0_outputs(7923) <= a or b;
    layer0_outputs(7924) <= a or b;
    layer0_outputs(7925) <= not (a or b);
    layer0_outputs(7926) <= not a;
    layer0_outputs(7927) <= a;
    layer0_outputs(7928) <= a xor b;
    layer0_outputs(7929) <= b;
    layer0_outputs(7930) <= b and not a;
    layer0_outputs(7931) <= b and not a;
    layer0_outputs(7932) <= not b;
    layer0_outputs(7933) <= not (a and b);
    layer0_outputs(7934) <= a and not b;
    layer0_outputs(7935) <= a and not b;
    layer0_outputs(7936) <= not b;
    layer0_outputs(7937) <= not b or a;
    layer0_outputs(7938) <= a xor b;
    layer0_outputs(7939) <= '0';
    layer0_outputs(7940) <= not b;
    layer0_outputs(7941) <= b and not a;
    layer0_outputs(7942) <= a or b;
    layer0_outputs(7943) <= '1';
    layer0_outputs(7944) <= a;
    layer0_outputs(7945) <= not a or b;
    layer0_outputs(7946) <= b;
    layer0_outputs(7947) <= b;
    layer0_outputs(7948) <= '0';
    layer0_outputs(7949) <= not b;
    layer0_outputs(7950) <= not (a or b);
    layer0_outputs(7951) <= not (a or b);
    layer0_outputs(7952) <= not b;
    layer0_outputs(7953) <= b and not a;
    layer0_outputs(7954) <= not b;
    layer0_outputs(7955) <= b and not a;
    layer0_outputs(7956) <= not b;
    layer0_outputs(7957) <= a and not b;
    layer0_outputs(7958) <= not b;
    layer0_outputs(7959) <= not a or b;
    layer0_outputs(7960) <= b;
    layer0_outputs(7961) <= a and not b;
    layer0_outputs(7962) <= a xor b;
    layer0_outputs(7963) <= a;
    layer0_outputs(7964) <= not a;
    layer0_outputs(7965) <= a xor b;
    layer0_outputs(7966) <= not a;
    layer0_outputs(7967) <= not (a or b);
    layer0_outputs(7968) <= a and not b;
    layer0_outputs(7969) <= not b or a;
    layer0_outputs(7970) <= a xor b;
    layer0_outputs(7971) <= '0';
    layer0_outputs(7972) <= not a;
    layer0_outputs(7973) <= not a or b;
    layer0_outputs(7974) <= a;
    layer0_outputs(7975) <= b;
    layer0_outputs(7976) <= not (a or b);
    layer0_outputs(7977) <= a or b;
    layer0_outputs(7978) <= a xor b;
    layer0_outputs(7979) <= b and not a;
    layer0_outputs(7980) <= not b;
    layer0_outputs(7981) <= not b;
    layer0_outputs(7982) <= a or b;
    layer0_outputs(7983) <= not (a or b);
    layer0_outputs(7984) <= not a or b;
    layer0_outputs(7985) <= not (a or b);
    layer0_outputs(7986) <= not a;
    layer0_outputs(7987) <= a xor b;
    layer0_outputs(7988) <= a;
    layer0_outputs(7989) <= a or b;
    layer0_outputs(7990) <= a and not b;
    layer0_outputs(7991) <= not (a xor b);
    layer0_outputs(7992) <= a xor b;
    layer0_outputs(7993) <= a or b;
    layer0_outputs(7994) <= a xor b;
    layer0_outputs(7995) <= a or b;
    layer0_outputs(7996) <= not b;
    layer0_outputs(7997) <= a or b;
    layer0_outputs(7998) <= b;
    layer0_outputs(7999) <= '1';
    layer0_outputs(8000) <= not a;
    layer0_outputs(8001) <= a or b;
    layer0_outputs(8002) <= not (a xor b);
    layer0_outputs(8003) <= not a;
    layer0_outputs(8004) <= a xor b;
    layer0_outputs(8005) <= not (a xor b);
    layer0_outputs(8006) <= b and not a;
    layer0_outputs(8007) <= '1';
    layer0_outputs(8008) <= not b;
    layer0_outputs(8009) <= a or b;
    layer0_outputs(8010) <= a xor b;
    layer0_outputs(8011) <= not b or a;
    layer0_outputs(8012) <= not (a xor b);
    layer0_outputs(8013) <= a;
    layer0_outputs(8014) <= b and not a;
    layer0_outputs(8015) <= not (a xor b);
    layer0_outputs(8016) <= not b;
    layer0_outputs(8017) <= '0';
    layer0_outputs(8018) <= a or b;
    layer0_outputs(8019) <= a and not b;
    layer0_outputs(8020) <= b;
    layer0_outputs(8021) <= not a;
    layer0_outputs(8022) <= a or b;
    layer0_outputs(8023) <= a;
    layer0_outputs(8024) <= not (a xor b);
    layer0_outputs(8025) <= not (a or b);
    layer0_outputs(8026) <= a;
    layer0_outputs(8027) <= '0';
    layer0_outputs(8028) <= a or b;
    layer0_outputs(8029) <= not (a xor b);
    layer0_outputs(8030) <= not b;
    layer0_outputs(8031) <= not (a or b);
    layer0_outputs(8032) <= a;
    layer0_outputs(8033) <= not a or b;
    layer0_outputs(8034) <= not b;
    layer0_outputs(8035) <= b and not a;
    layer0_outputs(8036) <= a or b;
    layer0_outputs(8037) <= b;
    layer0_outputs(8038) <= not b;
    layer0_outputs(8039) <= b;
    layer0_outputs(8040) <= a or b;
    layer0_outputs(8041) <= a and b;
    layer0_outputs(8042) <= b;
    layer0_outputs(8043) <= not (a xor b);
    layer0_outputs(8044) <= not a or b;
    layer0_outputs(8045) <= not (a or b);
    layer0_outputs(8046) <= a and not b;
    layer0_outputs(8047) <= not a;
    layer0_outputs(8048) <= not (a or b);
    layer0_outputs(8049) <= not (a xor b);
    layer0_outputs(8050) <= not b;
    layer0_outputs(8051) <= b;
    layer0_outputs(8052) <= a xor b;
    layer0_outputs(8053) <= not b or a;
    layer0_outputs(8054) <= a;
    layer0_outputs(8055) <= not (a xor b);
    layer0_outputs(8056) <= '1';
    layer0_outputs(8057) <= a or b;
    layer0_outputs(8058) <= '1';
    layer0_outputs(8059) <= a;
    layer0_outputs(8060) <= not b;
    layer0_outputs(8061) <= not (a and b);
    layer0_outputs(8062) <= a and not b;
    layer0_outputs(8063) <= a xor b;
    layer0_outputs(8064) <= not b or a;
    layer0_outputs(8065) <= not (a or b);
    layer0_outputs(8066) <= b;
    layer0_outputs(8067) <= b;
    layer0_outputs(8068) <= a xor b;
    layer0_outputs(8069) <= a and not b;
    layer0_outputs(8070) <= b and not a;
    layer0_outputs(8071) <= b;
    layer0_outputs(8072) <= a xor b;
    layer0_outputs(8073) <= a and b;
    layer0_outputs(8074) <= b;
    layer0_outputs(8075) <= not a;
    layer0_outputs(8076) <= not a;
    layer0_outputs(8077) <= a xor b;
    layer0_outputs(8078) <= a or b;
    layer0_outputs(8079) <= b and not a;
    layer0_outputs(8080) <= not a;
    layer0_outputs(8081) <= a or b;
    layer0_outputs(8082) <= not a or b;
    layer0_outputs(8083) <= b and not a;
    layer0_outputs(8084) <= a or b;
    layer0_outputs(8085) <= b and not a;
    layer0_outputs(8086) <= not (a or b);
    layer0_outputs(8087) <= not (a or b);
    layer0_outputs(8088) <= a xor b;
    layer0_outputs(8089) <= a xor b;
    layer0_outputs(8090) <= a xor b;
    layer0_outputs(8091) <= not (a or b);
    layer0_outputs(8092) <= b;
    layer0_outputs(8093) <= not a;
    layer0_outputs(8094) <= not (a or b);
    layer0_outputs(8095) <= not a;
    layer0_outputs(8096) <= not b or a;
    layer0_outputs(8097) <= not b or a;
    layer0_outputs(8098) <= not (a xor b);
    layer0_outputs(8099) <= not a;
    layer0_outputs(8100) <= not b;
    layer0_outputs(8101) <= a xor b;
    layer0_outputs(8102) <= a;
    layer0_outputs(8103) <= not b;
    layer0_outputs(8104) <= a or b;
    layer0_outputs(8105) <= a or b;
    layer0_outputs(8106) <= b and not a;
    layer0_outputs(8107) <= a or b;
    layer0_outputs(8108) <= not a;
    layer0_outputs(8109) <= b;
    layer0_outputs(8110) <= not b;
    layer0_outputs(8111) <= '1';
    layer0_outputs(8112) <= a;
    layer0_outputs(8113) <= a and not b;
    layer0_outputs(8114) <= not (a or b);
    layer0_outputs(8115) <= a xor b;
    layer0_outputs(8116) <= a xor b;
    layer0_outputs(8117) <= a;
    layer0_outputs(8118) <= a and not b;
    layer0_outputs(8119) <= a;
    layer0_outputs(8120) <= not b or a;
    layer0_outputs(8121) <= not (a or b);
    layer0_outputs(8122) <= not b;
    layer0_outputs(8123) <= a;
    layer0_outputs(8124) <= a and not b;
    layer0_outputs(8125) <= a or b;
    layer0_outputs(8126) <= not (a xor b);
    layer0_outputs(8127) <= not (a or b);
    layer0_outputs(8128) <= a or b;
    layer0_outputs(8129) <= a;
    layer0_outputs(8130) <= not a or b;
    layer0_outputs(8131) <= a and not b;
    layer0_outputs(8132) <= not (a xor b);
    layer0_outputs(8133) <= not (a and b);
    layer0_outputs(8134) <= a;
    layer0_outputs(8135) <= '0';
    layer0_outputs(8136) <= a xor b;
    layer0_outputs(8137) <= not a;
    layer0_outputs(8138) <= a;
    layer0_outputs(8139) <= a xor b;
    layer0_outputs(8140) <= not (a xor b);
    layer0_outputs(8141) <= not a;
    layer0_outputs(8142) <= not (a xor b);
    layer0_outputs(8143) <= not (a or b);
    layer0_outputs(8144) <= a;
    layer0_outputs(8145) <= not b;
    layer0_outputs(8146) <= a or b;
    layer0_outputs(8147) <= not b;
    layer0_outputs(8148) <= a xor b;
    layer0_outputs(8149) <= a xor b;
    layer0_outputs(8150) <= not a;
    layer0_outputs(8151) <= not (a or b);
    layer0_outputs(8152) <= not b or a;
    layer0_outputs(8153) <= a or b;
    layer0_outputs(8154) <= not b;
    layer0_outputs(8155) <= a and b;
    layer0_outputs(8156) <= not b or a;
    layer0_outputs(8157) <= not (a xor b);
    layer0_outputs(8158) <= b;
    layer0_outputs(8159) <= not a;
    layer0_outputs(8160) <= not b or a;
    layer0_outputs(8161) <= b and not a;
    layer0_outputs(8162) <= b;
    layer0_outputs(8163) <= not a or b;
    layer0_outputs(8164) <= not (a or b);
    layer0_outputs(8165) <= not a;
    layer0_outputs(8166) <= '1';
    layer0_outputs(8167) <= not a or b;
    layer0_outputs(8168) <= not b;
    layer0_outputs(8169) <= not (a or b);
    layer0_outputs(8170) <= b and not a;
    layer0_outputs(8171) <= not (a or b);
    layer0_outputs(8172) <= a;
    layer0_outputs(8173) <= not b;
    layer0_outputs(8174) <= not b;
    layer0_outputs(8175) <= not (a or b);
    layer0_outputs(8176) <= not (a or b);
    layer0_outputs(8177) <= not (a or b);
    layer0_outputs(8178) <= a or b;
    layer0_outputs(8179) <= a xor b;
    layer0_outputs(8180) <= not (a xor b);
    layer0_outputs(8181) <= a xor b;
    layer0_outputs(8182) <= a and b;
    layer0_outputs(8183) <= not (a or b);
    layer0_outputs(8184) <= a xor b;
    layer0_outputs(8185) <= not (a xor b);
    layer0_outputs(8186) <= a or b;
    layer0_outputs(8187) <= not a;
    layer0_outputs(8188) <= a and b;
    layer0_outputs(8189) <= b and not a;
    layer0_outputs(8190) <= a;
    layer0_outputs(8191) <= a xor b;
    layer0_outputs(8192) <= not (a xor b);
    layer0_outputs(8193) <= not a or b;
    layer0_outputs(8194) <= b and not a;
    layer0_outputs(8195) <= a or b;
    layer0_outputs(8196) <= a or b;
    layer0_outputs(8197) <= not (a and b);
    layer0_outputs(8198) <= not a;
    layer0_outputs(8199) <= not (a or b);
    layer0_outputs(8200) <= not (a or b);
    layer0_outputs(8201) <= '0';
    layer0_outputs(8202) <= b and not a;
    layer0_outputs(8203) <= not (a or b);
    layer0_outputs(8204) <= not b or a;
    layer0_outputs(8205) <= not b;
    layer0_outputs(8206) <= a and not b;
    layer0_outputs(8207) <= a and not b;
    layer0_outputs(8208) <= not (a xor b);
    layer0_outputs(8209) <= not a or b;
    layer0_outputs(8210) <= a;
    layer0_outputs(8211) <= a;
    layer0_outputs(8212) <= a;
    layer0_outputs(8213) <= not a;
    layer0_outputs(8214) <= not b;
    layer0_outputs(8215) <= a xor b;
    layer0_outputs(8216) <= not (a or b);
    layer0_outputs(8217) <= a xor b;
    layer0_outputs(8218) <= not b or a;
    layer0_outputs(8219) <= a and b;
    layer0_outputs(8220) <= a or b;
    layer0_outputs(8221) <= not a or b;
    layer0_outputs(8222) <= b;
    layer0_outputs(8223) <= not (a and b);
    layer0_outputs(8224) <= a and not b;
    layer0_outputs(8225) <= a or b;
    layer0_outputs(8226) <= not a;
    layer0_outputs(8227) <= b and not a;
    layer0_outputs(8228) <= b and not a;
    layer0_outputs(8229) <= a or b;
    layer0_outputs(8230) <= not (a xor b);
    layer0_outputs(8231) <= not b;
    layer0_outputs(8232) <= not (a and b);
    layer0_outputs(8233) <= a xor b;
    layer0_outputs(8234) <= '0';
    layer0_outputs(8235) <= not a or b;
    layer0_outputs(8236) <= not b or a;
    layer0_outputs(8237) <= a or b;
    layer0_outputs(8238) <= not (a or b);
    layer0_outputs(8239) <= a and not b;
    layer0_outputs(8240) <= b and not a;
    layer0_outputs(8241) <= b;
    layer0_outputs(8242) <= not (a xor b);
    layer0_outputs(8243) <= not a;
    layer0_outputs(8244) <= not (a or b);
    layer0_outputs(8245) <= a or b;
    layer0_outputs(8246) <= not (a xor b);
    layer0_outputs(8247) <= not a or b;
    layer0_outputs(8248) <= not a;
    layer0_outputs(8249) <= not (a or b);
    layer0_outputs(8250) <= a xor b;
    layer0_outputs(8251) <= a or b;
    layer0_outputs(8252) <= b;
    layer0_outputs(8253) <= a or b;
    layer0_outputs(8254) <= not (a xor b);
    layer0_outputs(8255) <= a and b;
    layer0_outputs(8256) <= not (a or b);
    layer0_outputs(8257) <= not (a xor b);
    layer0_outputs(8258) <= '0';
    layer0_outputs(8259) <= a or b;
    layer0_outputs(8260) <= a and not b;
    layer0_outputs(8261) <= a and not b;
    layer0_outputs(8262) <= '1';
    layer0_outputs(8263) <= a or b;
    layer0_outputs(8264) <= not a or b;
    layer0_outputs(8265) <= a or b;
    layer0_outputs(8266) <= not (a xor b);
    layer0_outputs(8267) <= a;
    layer0_outputs(8268) <= not (a xor b);
    layer0_outputs(8269) <= not a or b;
    layer0_outputs(8270) <= a or b;
    layer0_outputs(8271) <= not a;
    layer0_outputs(8272) <= not a;
    layer0_outputs(8273) <= not b;
    layer0_outputs(8274) <= a or b;
    layer0_outputs(8275) <= a xor b;
    layer0_outputs(8276) <= not (a xor b);
    layer0_outputs(8277) <= b and not a;
    layer0_outputs(8278) <= '0';
    layer0_outputs(8279) <= not a;
    layer0_outputs(8280) <= b;
    layer0_outputs(8281) <= not (a xor b);
    layer0_outputs(8282) <= a and not b;
    layer0_outputs(8283) <= not a;
    layer0_outputs(8284) <= a;
    layer0_outputs(8285) <= '1';
    layer0_outputs(8286) <= a or b;
    layer0_outputs(8287) <= not b or a;
    layer0_outputs(8288) <= not a;
    layer0_outputs(8289) <= not (a and b);
    layer0_outputs(8290) <= a and not b;
    layer0_outputs(8291) <= a or b;
    layer0_outputs(8292) <= a xor b;
    layer0_outputs(8293) <= not a;
    layer0_outputs(8294) <= not a;
    layer0_outputs(8295) <= not b;
    layer0_outputs(8296) <= not b;
    layer0_outputs(8297) <= not b or a;
    layer0_outputs(8298) <= b and not a;
    layer0_outputs(8299) <= not (a xor b);
    layer0_outputs(8300) <= a;
    layer0_outputs(8301) <= not a or b;
    layer0_outputs(8302) <= a or b;
    layer0_outputs(8303) <= not (a xor b);
    layer0_outputs(8304) <= b;
    layer0_outputs(8305) <= not b or a;
    layer0_outputs(8306) <= a and b;
    layer0_outputs(8307) <= b;
    layer0_outputs(8308) <= a or b;
    layer0_outputs(8309) <= not (a xor b);
    layer0_outputs(8310) <= a or b;
    layer0_outputs(8311) <= a xor b;
    layer0_outputs(8312) <= b and not a;
    layer0_outputs(8313) <= b and not a;
    layer0_outputs(8314) <= not (a xor b);
    layer0_outputs(8315) <= a xor b;
    layer0_outputs(8316) <= a or b;
    layer0_outputs(8317) <= a or b;
    layer0_outputs(8318) <= a or b;
    layer0_outputs(8319) <= a xor b;
    layer0_outputs(8320) <= not (a or b);
    layer0_outputs(8321) <= not (a or b);
    layer0_outputs(8322) <= a or b;
    layer0_outputs(8323) <= a xor b;
    layer0_outputs(8324) <= not (a or b);
    layer0_outputs(8325) <= not a or b;
    layer0_outputs(8326) <= not (a xor b);
    layer0_outputs(8327) <= a;
    layer0_outputs(8328) <= a and not b;
    layer0_outputs(8329) <= not (a or b);
    layer0_outputs(8330) <= b and not a;
    layer0_outputs(8331) <= not (a xor b);
    layer0_outputs(8332) <= not (a xor b);
    layer0_outputs(8333) <= not (a xor b);
    layer0_outputs(8334) <= not a or b;
    layer0_outputs(8335) <= a or b;
    layer0_outputs(8336) <= b and not a;
    layer0_outputs(8337) <= a xor b;
    layer0_outputs(8338) <= a and not b;
    layer0_outputs(8339) <= a xor b;
    layer0_outputs(8340) <= a and not b;
    layer0_outputs(8341) <= not b;
    layer0_outputs(8342) <= not b or a;
    layer0_outputs(8343) <= a xor b;
    layer0_outputs(8344) <= not a;
    layer0_outputs(8345) <= a xor b;
    layer0_outputs(8346) <= not (a or b);
    layer0_outputs(8347) <= not b or a;
    layer0_outputs(8348) <= not a or b;
    layer0_outputs(8349) <= not (a and b);
    layer0_outputs(8350) <= a xor b;
    layer0_outputs(8351) <= a and b;
    layer0_outputs(8352) <= not (a xor b);
    layer0_outputs(8353) <= not b or a;
    layer0_outputs(8354) <= a and not b;
    layer0_outputs(8355) <= a xor b;
    layer0_outputs(8356) <= not (a or b);
    layer0_outputs(8357) <= not (a or b);
    layer0_outputs(8358) <= b;
    layer0_outputs(8359) <= not b or a;
    layer0_outputs(8360) <= a or b;
    layer0_outputs(8361) <= b and not a;
    layer0_outputs(8362) <= not b or a;
    layer0_outputs(8363) <= not (a xor b);
    layer0_outputs(8364) <= not a;
    layer0_outputs(8365) <= a and b;
    layer0_outputs(8366) <= a and not b;
    layer0_outputs(8367) <= not b or a;
    layer0_outputs(8368) <= b;
    layer0_outputs(8369) <= not a or b;
    layer0_outputs(8370) <= a or b;
    layer0_outputs(8371) <= a or b;
    layer0_outputs(8372) <= a or b;
    layer0_outputs(8373) <= b and not a;
    layer0_outputs(8374) <= b;
    layer0_outputs(8375) <= b;
    layer0_outputs(8376) <= not a or b;
    layer0_outputs(8377) <= not b;
    layer0_outputs(8378) <= a;
    layer0_outputs(8379) <= not (a xor b);
    layer0_outputs(8380) <= not b;
    layer0_outputs(8381) <= not (a or b);
    layer0_outputs(8382) <= b and not a;
    layer0_outputs(8383) <= not a or b;
    layer0_outputs(8384) <= not a or b;
    layer0_outputs(8385) <= a and not b;
    layer0_outputs(8386) <= not (a xor b);
    layer0_outputs(8387) <= not a;
    layer0_outputs(8388) <= a;
    layer0_outputs(8389) <= a or b;
    layer0_outputs(8390) <= a and not b;
    layer0_outputs(8391) <= not (a xor b);
    layer0_outputs(8392) <= not (a xor b);
    layer0_outputs(8393) <= '1';
    layer0_outputs(8394) <= b;
    layer0_outputs(8395) <= not (a xor b);
    layer0_outputs(8396) <= not b or a;
    layer0_outputs(8397) <= a and not b;
    layer0_outputs(8398) <= a;
    layer0_outputs(8399) <= a;
    layer0_outputs(8400) <= a xor b;
    layer0_outputs(8401) <= not (a xor b);
    layer0_outputs(8402) <= a;
    layer0_outputs(8403) <= a xor b;
    layer0_outputs(8404) <= a or b;
    layer0_outputs(8405) <= not (a or b);
    layer0_outputs(8406) <= a or b;
    layer0_outputs(8407) <= a and not b;
    layer0_outputs(8408) <= not b;
    layer0_outputs(8409) <= not b or a;
    layer0_outputs(8410) <= a and b;
    layer0_outputs(8411) <= b and not a;
    layer0_outputs(8412) <= not b;
    layer0_outputs(8413) <= a and b;
    layer0_outputs(8414) <= not (a or b);
    layer0_outputs(8415) <= b and not a;
    layer0_outputs(8416) <= not (a or b);
    layer0_outputs(8417) <= a or b;
    layer0_outputs(8418) <= b and not a;
    layer0_outputs(8419) <= not (a xor b);
    layer0_outputs(8420) <= b and not a;
    layer0_outputs(8421) <= a xor b;
    layer0_outputs(8422) <= a or b;
    layer0_outputs(8423) <= not a;
    layer0_outputs(8424) <= not a or b;
    layer0_outputs(8425) <= not a;
    layer0_outputs(8426) <= not b or a;
    layer0_outputs(8427) <= a and b;
    layer0_outputs(8428) <= not b;
    layer0_outputs(8429) <= not b or a;
    layer0_outputs(8430) <= not (a or b);
    layer0_outputs(8431) <= a or b;
    layer0_outputs(8432) <= not a;
    layer0_outputs(8433) <= a or b;
    layer0_outputs(8434) <= b;
    layer0_outputs(8435) <= a;
    layer0_outputs(8436) <= a xor b;
    layer0_outputs(8437) <= not a;
    layer0_outputs(8438) <= a or b;
    layer0_outputs(8439) <= b and not a;
    layer0_outputs(8440) <= a xor b;
    layer0_outputs(8441) <= a and not b;
    layer0_outputs(8442) <= a;
    layer0_outputs(8443) <= b;
    layer0_outputs(8444) <= a;
    layer0_outputs(8445) <= not (a or b);
    layer0_outputs(8446) <= a;
    layer0_outputs(8447) <= b and not a;
    layer0_outputs(8448) <= not a or b;
    layer0_outputs(8449) <= not (a or b);
    layer0_outputs(8450) <= not (a xor b);
    layer0_outputs(8451) <= not a or b;
    layer0_outputs(8452) <= not (a or b);
    layer0_outputs(8453) <= not a or b;
    layer0_outputs(8454) <= b and not a;
    layer0_outputs(8455) <= not (a xor b);
    layer0_outputs(8456) <= a and not b;
    layer0_outputs(8457) <= not a or b;
    layer0_outputs(8458) <= not (a or b);
    layer0_outputs(8459) <= b and not a;
    layer0_outputs(8460) <= not (a xor b);
    layer0_outputs(8461) <= not b or a;
    layer0_outputs(8462) <= not a;
    layer0_outputs(8463) <= b;
    layer0_outputs(8464) <= a or b;
    layer0_outputs(8465) <= not b;
    layer0_outputs(8466) <= a xor b;
    layer0_outputs(8467) <= a or b;
    layer0_outputs(8468) <= a;
    layer0_outputs(8469) <= not a;
    layer0_outputs(8470) <= not (a xor b);
    layer0_outputs(8471) <= a xor b;
    layer0_outputs(8472) <= a and not b;
    layer0_outputs(8473) <= b;
    layer0_outputs(8474) <= not b;
    layer0_outputs(8475) <= not b;
    layer0_outputs(8476) <= not a;
    layer0_outputs(8477) <= b and not a;
    layer0_outputs(8478) <= not a or b;
    layer0_outputs(8479) <= not a or b;
    layer0_outputs(8480) <= not b;
    layer0_outputs(8481) <= a or b;
    layer0_outputs(8482) <= not (a xor b);
    layer0_outputs(8483) <= not (a or b);
    layer0_outputs(8484) <= not (a or b);
    layer0_outputs(8485) <= a and not b;
    layer0_outputs(8486) <= not b or a;
    layer0_outputs(8487) <= not a or b;
    layer0_outputs(8488) <= a and b;
    layer0_outputs(8489) <= a;
    layer0_outputs(8490) <= not b or a;
    layer0_outputs(8491) <= not (a xor b);
    layer0_outputs(8492) <= a and not b;
    layer0_outputs(8493) <= a or b;
    layer0_outputs(8494) <= not b;
    layer0_outputs(8495) <= a;
    layer0_outputs(8496) <= not (a xor b);
    layer0_outputs(8497) <= not (a or b);
    layer0_outputs(8498) <= not (a or b);
    layer0_outputs(8499) <= not b;
    layer0_outputs(8500) <= not (a xor b);
    layer0_outputs(8501) <= a xor b;
    layer0_outputs(8502) <= not a;
    layer0_outputs(8503) <= a or b;
    layer0_outputs(8504) <= not a;
    layer0_outputs(8505) <= not (a xor b);
    layer0_outputs(8506) <= not a;
    layer0_outputs(8507) <= not b or a;
    layer0_outputs(8508) <= b and not a;
    layer0_outputs(8509) <= not b;
    layer0_outputs(8510) <= a or b;
    layer0_outputs(8511) <= not a or b;
    layer0_outputs(8512) <= not (a xor b);
    layer0_outputs(8513) <= not (a and b);
    layer0_outputs(8514) <= b;
    layer0_outputs(8515) <= not b;
    layer0_outputs(8516) <= a xor b;
    layer0_outputs(8517) <= not (a or b);
    layer0_outputs(8518) <= not (a or b);
    layer0_outputs(8519) <= not (a xor b);
    layer0_outputs(8520) <= not (a or b);
    layer0_outputs(8521) <= a and b;
    layer0_outputs(8522) <= a and b;
    layer0_outputs(8523) <= a or b;
    layer0_outputs(8524) <= a xor b;
    layer0_outputs(8525) <= a xor b;
    layer0_outputs(8526) <= a or b;
    layer0_outputs(8527) <= not b;
    layer0_outputs(8528) <= a and not b;
    layer0_outputs(8529) <= not a;
    layer0_outputs(8530) <= a or b;
    layer0_outputs(8531) <= not b;
    layer0_outputs(8532) <= a or b;
    layer0_outputs(8533) <= not (a xor b);
    layer0_outputs(8534) <= not b;
    layer0_outputs(8535) <= not (a or b);
    layer0_outputs(8536) <= not a;
    layer0_outputs(8537) <= a and b;
    layer0_outputs(8538) <= not a;
    layer0_outputs(8539) <= a;
    layer0_outputs(8540) <= a xor b;
    layer0_outputs(8541) <= '1';
    layer0_outputs(8542) <= b and not a;
    layer0_outputs(8543) <= a;
    layer0_outputs(8544) <= a and not b;
    layer0_outputs(8545) <= not (a xor b);
    layer0_outputs(8546) <= b;
    layer0_outputs(8547) <= not b;
    layer0_outputs(8548) <= not a;
    layer0_outputs(8549) <= '1';
    layer0_outputs(8550) <= not b;
    layer0_outputs(8551) <= '1';
    layer0_outputs(8552) <= a xor b;
    layer0_outputs(8553) <= not a or b;
    layer0_outputs(8554) <= b;
    layer0_outputs(8555) <= b and not a;
    layer0_outputs(8556) <= a or b;
    layer0_outputs(8557) <= not (a or b);
    layer0_outputs(8558) <= b;
    layer0_outputs(8559) <= b;
    layer0_outputs(8560) <= not a;
    layer0_outputs(8561) <= a;
    layer0_outputs(8562) <= a or b;
    layer0_outputs(8563) <= b;
    layer0_outputs(8564) <= not a or b;
    layer0_outputs(8565) <= a;
    layer0_outputs(8566) <= b;
    layer0_outputs(8567) <= not b or a;
    layer0_outputs(8568) <= a and not b;
    layer0_outputs(8569) <= not (a or b);
    layer0_outputs(8570) <= not a or b;
    layer0_outputs(8571) <= not b or a;
    layer0_outputs(8572) <= a or b;
    layer0_outputs(8573) <= a xor b;
    layer0_outputs(8574) <= b;
    layer0_outputs(8575) <= not b or a;
    layer0_outputs(8576) <= not b or a;
    layer0_outputs(8577) <= a;
    layer0_outputs(8578) <= not a;
    layer0_outputs(8579) <= not (a xor b);
    layer0_outputs(8580) <= not (a or b);
    layer0_outputs(8581) <= '0';
    layer0_outputs(8582) <= b and not a;
    layer0_outputs(8583) <= not (a or b);
    layer0_outputs(8584) <= not (a xor b);
    layer0_outputs(8585) <= not (a or b);
    layer0_outputs(8586) <= b;
    layer0_outputs(8587) <= not (a or b);
    layer0_outputs(8588) <= b and not a;
    layer0_outputs(8589) <= a and not b;
    layer0_outputs(8590) <= b;
    layer0_outputs(8591) <= not a or b;
    layer0_outputs(8592) <= not (a or b);
    layer0_outputs(8593) <= not a;
    layer0_outputs(8594) <= not a;
    layer0_outputs(8595) <= a;
    layer0_outputs(8596) <= a and b;
    layer0_outputs(8597) <= not b;
    layer0_outputs(8598) <= not (a xor b);
    layer0_outputs(8599) <= a or b;
    layer0_outputs(8600) <= a or b;
    layer0_outputs(8601) <= not (a or b);
    layer0_outputs(8602) <= not (a xor b);
    layer0_outputs(8603) <= a or b;
    layer0_outputs(8604) <= not b or a;
    layer0_outputs(8605) <= a and b;
    layer0_outputs(8606) <= a;
    layer0_outputs(8607) <= not b;
    layer0_outputs(8608) <= not (a or b);
    layer0_outputs(8609) <= b and not a;
    layer0_outputs(8610) <= not a or b;
    layer0_outputs(8611) <= not (a or b);
    layer0_outputs(8612) <= not a;
    layer0_outputs(8613) <= b and not a;
    layer0_outputs(8614) <= a xor b;
    layer0_outputs(8615) <= not (a or b);
    layer0_outputs(8616) <= b and not a;
    layer0_outputs(8617) <= b;
    layer0_outputs(8618) <= not (a or b);
    layer0_outputs(8619) <= a and b;
    layer0_outputs(8620) <= not (a xor b);
    layer0_outputs(8621) <= a;
    layer0_outputs(8622) <= a and not b;
    layer0_outputs(8623) <= not (a or b);
    layer0_outputs(8624) <= '0';
    layer0_outputs(8625) <= a and b;
    layer0_outputs(8626) <= not (a xor b);
    layer0_outputs(8627) <= not a or b;
    layer0_outputs(8628) <= a xor b;
    layer0_outputs(8629) <= not b or a;
    layer0_outputs(8630) <= b and not a;
    layer0_outputs(8631) <= not (a xor b);
    layer0_outputs(8632) <= a or b;
    layer0_outputs(8633) <= a and not b;
    layer0_outputs(8634) <= not (a xor b);
    layer0_outputs(8635) <= not a;
    layer0_outputs(8636) <= b;
    layer0_outputs(8637) <= a;
    layer0_outputs(8638) <= not a or b;
    layer0_outputs(8639) <= a or b;
    layer0_outputs(8640) <= not (a or b);
    layer0_outputs(8641) <= not (a or b);
    layer0_outputs(8642) <= b and not a;
    layer0_outputs(8643) <= not (a or b);
    layer0_outputs(8644) <= not b;
    layer0_outputs(8645) <= not (a or b);
    layer0_outputs(8646) <= not a;
    layer0_outputs(8647) <= a and b;
    layer0_outputs(8648) <= a and not b;
    layer0_outputs(8649) <= not a;
    layer0_outputs(8650) <= a xor b;
    layer0_outputs(8651) <= a or b;
    layer0_outputs(8652) <= b;
    layer0_outputs(8653) <= not (a xor b);
    layer0_outputs(8654) <= not a or b;
    layer0_outputs(8655) <= '1';
    layer0_outputs(8656) <= a or b;
    layer0_outputs(8657) <= a or b;
    layer0_outputs(8658) <= '1';
    layer0_outputs(8659) <= a;
    layer0_outputs(8660) <= b;
    layer0_outputs(8661) <= not a or b;
    layer0_outputs(8662) <= not b or a;
    layer0_outputs(8663) <= a or b;
    layer0_outputs(8664) <= not (a or b);
    layer0_outputs(8665) <= a;
    layer0_outputs(8666) <= not a;
    layer0_outputs(8667) <= b;
    layer0_outputs(8668) <= a xor b;
    layer0_outputs(8669) <= a and not b;
    layer0_outputs(8670) <= not (a xor b);
    layer0_outputs(8671) <= not (a xor b);
    layer0_outputs(8672) <= not (a and b);
    layer0_outputs(8673) <= a or b;
    layer0_outputs(8674) <= a or b;
    layer0_outputs(8675) <= a and b;
    layer0_outputs(8676) <= not a;
    layer0_outputs(8677) <= not (a or b);
    layer0_outputs(8678) <= a or b;
    layer0_outputs(8679) <= a xor b;
    layer0_outputs(8680) <= a and not b;
    layer0_outputs(8681) <= b and not a;
    layer0_outputs(8682) <= a or b;
    layer0_outputs(8683) <= '0';
    layer0_outputs(8684) <= not (a or b);
    layer0_outputs(8685) <= not (a xor b);
    layer0_outputs(8686) <= not b;
    layer0_outputs(8687) <= not (a xor b);
    layer0_outputs(8688) <= a and not b;
    layer0_outputs(8689) <= a or b;
    layer0_outputs(8690) <= not (a xor b);
    layer0_outputs(8691) <= not a;
    layer0_outputs(8692) <= a and not b;
    layer0_outputs(8693) <= not a or b;
    layer0_outputs(8694) <= a or b;
    layer0_outputs(8695) <= a and b;
    layer0_outputs(8696) <= b and not a;
    layer0_outputs(8697) <= b and not a;
    layer0_outputs(8698) <= a or b;
    layer0_outputs(8699) <= not a or b;
    layer0_outputs(8700) <= not (a xor b);
    layer0_outputs(8701) <= not (a and b);
    layer0_outputs(8702) <= a or b;
    layer0_outputs(8703) <= not (a or b);
    layer0_outputs(8704) <= not (a xor b);
    layer0_outputs(8705) <= a or b;
    layer0_outputs(8706) <= not b or a;
    layer0_outputs(8707) <= b;
    layer0_outputs(8708) <= not (a or b);
    layer0_outputs(8709) <= not (a or b);
    layer0_outputs(8710) <= a;
    layer0_outputs(8711) <= a xor b;
    layer0_outputs(8712) <= not (a or b);
    layer0_outputs(8713) <= a;
    layer0_outputs(8714) <= b and not a;
    layer0_outputs(8715) <= not (a xor b);
    layer0_outputs(8716) <= not (a or b);
    layer0_outputs(8717) <= b and not a;
    layer0_outputs(8718) <= a;
    layer0_outputs(8719) <= not a or b;
    layer0_outputs(8720) <= not (a xor b);
    layer0_outputs(8721) <= a or b;
    layer0_outputs(8722) <= a and not b;
    layer0_outputs(8723) <= a and b;
    layer0_outputs(8724) <= b and not a;
    layer0_outputs(8725) <= a xor b;
    layer0_outputs(8726) <= not (a or b);
    layer0_outputs(8727) <= not (a or b);
    layer0_outputs(8728) <= not a or b;
    layer0_outputs(8729) <= a or b;
    layer0_outputs(8730) <= not b;
    layer0_outputs(8731) <= not b or a;
    layer0_outputs(8732) <= not a or b;
    layer0_outputs(8733) <= not a or b;
    layer0_outputs(8734) <= not (a or b);
    layer0_outputs(8735) <= a or b;
    layer0_outputs(8736) <= not (a or b);
    layer0_outputs(8737) <= a xor b;
    layer0_outputs(8738) <= a or b;
    layer0_outputs(8739) <= not (a or b);
    layer0_outputs(8740) <= a or b;
    layer0_outputs(8741) <= a or b;
    layer0_outputs(8742) <= not a or b;
    layer0_outputs(8743) <= b;
    layer0_outputs(8744) <= not a;
    layer0_outputs(8745) <= a or b;
    layer0_outputs(8746) <= not a or b;
    layer0_outputs(8747) <= a and not b;
    layer0_outputs(8748) <= not (a xor b);
    layer0_outputs(8749) <= a or b;
    layer0_outputs(8750) <= not (a or b);
    layer0_outputs(8751) <= not a;
    layer0_outputs(8752) <= not b;
    layer0_outputs(8753) <= not a;
    layer0_outputs(8754) <= not (a or b);
    layer0_outputs(8755) <= '1';
    layer0_outputs(8756) <= a and not b;
    layer0_outputs(8757) <= not (a xor b);
    layer0_outputs(8758) <= a;
    layer0_outputs(8759) <= not a;
    layer0_outputs(8760) <= b;
    layer0_outputs(8761) <= not b;
    layer0_outputs(8762) <= not a or b;
    layer0_outputs(8763) <= not (a xor b);
    layer0_outputs(8764) <= b and not a;
    layer0_outputs(8765) <= not a or b;
    layer0_outputs(8766) <= b;
    layer0_outputs(8767) <= a or b;
    layer0_outputs(8768) <= a;
    layer0_outputs(8769) <= not a or b;
    layer0_outputs(8770) <= not a;
    layer0_outputs(8771) <= a or b;
    layer0_outputs(8772) <= a or b;
    layer0_outputs(8773) <= a;
    layer0_outputs(8774) <= not b or a;
    layer0_outputs(8775) <= a or b;
    layer0_outputs(8776) <= a xor b;
    layer0_outputs(8777) <= not (a or b);
    layer0_outputs(8778) <= a and not b;
    layer0_outputs(8779) <= not (a or b);
    layer0_outputs(8780) <= not (a or b);
    layer0_outputs(8781) <= not (a xor b);
    layer0_outputs(8782) <= a and not b;
    layer0_outputs(8783) <= not (a and b);
    layer0_outputs(8784) <= a xor b;
    layer0_outputs(8785) <= '1';
    layer0_outputs(8786) <= not b or a;
    layer0_outputs(8787) <= not (a xor b);
    layer0_outputs(8788) <= a and not b;
    layer0_outputs(8789) <= not (a xor b);
    layer0_outputs(8790) <= a or b;
    layer0_outputs(8791) <= b and not a;
    layer0_outputs(8792) <= not (a or b);
    layer0_outputs(8793) <= not b;
    layer0_outputs(8794) <= '1';
    layer0_outputs(8795) <= b and not a;
    layer0_outputs(8796) <= a xor b;
    layer0_outputs(8797) <= not a;
    layer0_outputs(8798) <= not a or b;
    layer0_outputs(8799) <= not (a or b);
    layer0_outputs(8800) <= a xor b;
    layer0_outputs(8801) <= a or b;
    layer0_outputs(8802) <= a xor b;
    layer0_outputs(8803) <= not a;
    layer0_outputs(8804) <= a xor b;
    layer0_outputs(8805) <= a and not b;
    layer0_outputs(8806) <= a or b;
    layer0_outputs(8807) <= b;
    layer0_outputs(8808) <= not a;
    layer0_outputs(8809) <= a;
    layer0_outputs(8810) <= '1';
    layer0_outputs(8811) <= not a;
    layer0_outputs(8812) <= not (a xor b);
    layer0_outputs(8813) <= b and not a;
    layer0_outputs(8814) <= not b;
    layer0_outputs(8815) <= a;
    layer0_outputs(8816) <= not (a or b);
    layer0_outputs(8817) <= b and not a;
    layer0_outputs(8818) <= a or b;
    layer0_outputs(8819) <= a and not b;
    layer0_outputs(8820) <= b and not a;
    layer0_outputs(8821) <= not (a or b);
    layer0_outputs(8822) <= not b;
    layer0_outputs(8823) <= not a;
    layer0_outputs(8824) <= not b;
    layer0_outputs(8825) <= not b or a;
    layer0_outputs(8826) <= a and not b;
    layer0_outputs(8827) <= not a or b;
    layer0_outputs(8828) <= not (a or b);
    layer0_outputs(8829) <= a or b;
    layer0_outputs(8830) <= a xor b;
    layer0_outputs(8831) <= not a or b;
    layer0_outputs(8832) <= not b or a;
    layer0_outputs(8833) <= not (a or b);
    layer0_outputs(8834) <= not b;
    layer0_outputs(8835) <= not (a or b);
    layer0_outputs(8836) <= not a or b;
    layer0_outputs(8837) <= not (a or b);
    layer0_outputs(8838) <= not (a or b);
    layer0_outputs(8839) <= a or b;
    layer0_outputs(8840) <= a and not b;
    layer0_outputs(8841) <= not b;
    layer0_outputs(8842) <= a or b;
    layer0_outputs(8843) <= not (a or b);
    layer0_outputs(8844) <= not (a or b);
    layer0_outputs(8845) <= not (a xor b);
    layer0_outputs(8846) <= b and not a;
    layer0_outputs(8847) <= a;
    layer0_outputs(8848) <= a and not b;
    layer0_outputs(8849) <= a xor b;
    layer0_outputs(8850) <= not (a and b);
    layer0_outputs(8851) <= not a;
    layer0_outputs(8852) <= a;
    layer0_outputs(8853) <= not b or a;
    layer0_outputs(8854) <= not (a xor b);
    layer0_outputs(8855) <= a xor b;
    layer0_outputs(8856) <= not (a and b);
    layer0_outputs(8857) <= not (a or b);
    layer0_outputs(8858) <= b and not a;
    layer0_outputs(8859) <= not (a and b);
    layer0_outputs(8860) <= not b;
    layer0_outputs(8861) <= '0';
    layer0_outputs(8862) <= a;
    layer0_outputs(8863) <= not (a or b);
    layer0_outputs(8864) <= not (a or b);
    layer0_outputs(8865) <= not (a and b);
    layer0_outputs(8866) <= a xor b;
    layer0_outputs(8867) <= a xor b;
    layer0_outputs(8868) <= not (a or b);
    layer0_outputs(8869) <= a or b;
    layer0_outputs(8870) <= a and b;
    layer0_outputs(8871) <= b;
    layer0_outputs(8872) <= not b or a;
    layer0_outputs(8873) <= not (a or b);
    layer0_outputs(8874) <= not (a xor b);
    layer0_outputs(8875) <= not a or b;
    layer0_outputs(8876) <= '0';
    layer0_outputs(8877) <= a and b;
    layer0_outputs(8878) <= a or b;
    layer0_outputs(8879) <= not b;
    layer0_outputs(8880) <= '1';
    layer0_outputs(8881) <= not (a or b);
    layer0_outputs(8882) <= b;
    layer0_outputs(8883) <= not (a xor b);
    layer0_outputs(8884) <= not a;
    layer0_outputs(8885) <= not a or b;
    layer0_outputs(8886) <= not a;
    layer0_outputs(8887) <= b;
    layer0_outputs(8888) <= a xor b;
    layer0_outputs(8889) <= a or b;
    layer0_outputs(8890) <= a or b;
    layer0_outputs(8891) <= b and not a;
    layer0_outputs(8892) <= b;
    layer0_outputs(8893) <= b;
    layer0_outputs(8894) <= not b or a;
    layer0_outputs(8895) <= a or b;
    layer0_outputs(8896) <= not a or b;
    layer0_outputs(8897) <= not b or a;
    layer0_outputs(8898) <= a and not b;
    layer0_outputs(8899) <= not b;
    layer0_outputs(8900) <= not (a or b);
    layer0_outputs(8901) <= not (a or b);
    layer0_outputs(8902) <= a;
    layer0_outputs(8903) <= a or b;
    layer0_outputs(8904) <= not (a or b);
    layer0_outputs(8905) <= b;
    layer0_outputs(8906) <= not b;
    layer0_outputs(8907) <= b and not a;
    layer0_outputs(8908) <= b;
    layer0_outputs(8909) <= not (a xor b);
    layer0_outputs(8910) <= not a or b;
    layer0_outputs(8911) <= not (a or b);
    layer0_outputs(8912) <= not (a xor b);
    layer0_outputs(8913) <= '1';
    layer0_outputs(8914) <= not (a or b);
    layer0_outputs(8915) <= b;
    layer0_outputs(8916) <= a or b;
    layer0_outputs(8917) <= b and not a;
    layer0_outputs(8918) <= not (a or b);
    layer0_outputs(8919) <= a and not b;
    layer0_outputs(8920) <= b;
    layer0_outputs(8921) <= not b or a;
    layer0_outputs(8922) <= b and not a;
    layer0_outputs(8923) <= not b or a;
    layer0_outputs(8924) <= '1';
    layer0_outputs(8925) <= a xor b;
    layer0_outputs(8926) <= not (a xor b);
    layer0_outputs(8927) <= not (a xor b);
    layer0_outputs(8928) <= not (a or b);
    layer0_outputs(8929) <= not a;
    layer0_outputs(8930) <= a xor b;
    layer0_outputs(8931) <= a or b;
    layer0_outputs(8932) <= not (a or b);
    layer0_outputs(8933) <= a xor b;
    layer0_outputs(8934) <= not b;
    layer0_outputs(8935) <= a or b;
    layer0_outputs(8936) <= a xor b;
    layer0_outputs(8937) <= not (a or b);
    layer0_outputs(8938) <= not b or a;
    layer0_outputs(8939) <= not a;
    layer0_outputs(8940) <= not b;
    layer0_outputs(8941) <= b;
    layer0_outputs(8942) <= a xor b;
    layer0_outputs(8943) <= not (a xor b);
    layer0_outputs(8944) <= not a;
    layer0_outputs(8945) <= not (a or b);
    layer0_outputs(8946) <= a xor b;
    layer0_outputs(8947) <= not b;
    layer0_outputs(8948) <= not a;
    layer0_outputs(8949) <= a or b;
    layer0_outputs(8950) <= not (a xor b);
    layer0_outputs(8951) <= not a;
    layer0_outputs(8952) <= a and not b;
    layer0_outputs(8953) <= a xor b;
    layer0_outputs(8954) <= a or b;
    layer0_outputs(8955) <= a or b;
    layer0_outputs(8956) <= a;
    layer0_outputs(8957) <= not a or b;
    layer0_outputs(8958) <= a and not b;
    layer0_outputs(8959) <= b;
    layer0_outputs(8960) <= b;
    layer0_outputs(8961) <= a xor b;
    layer0_outputs(8962) <= a or b;
    layer0_outputs(8963) <= a and not b;
    layer0_outputs(8964) <= a xor b;
    layer0_outputs(8965) <= not a;
    layer0_outputs(8966) <= not a or b;
    layer0_outputs(8967) <= not (a or b);
    layer0_outputs(8968) <= not (a xor b);
    layer0_outputs(8969) <= not (a or b);
    layer0_outputs(8970) <= b;
    layer0_outputs(8971) <= a and not b;
    layer0_outputs(8972) <= not (a or b);
    layer0_outputs(8973) <= not (a or b);
    layer0_outputs(8974) <= not a;
    layer0_outputs(8975) <= not (a and b);
    layer0_outputs(8976) <= a or b;
    layer0_outputs(8977) <= '1';
    layer0_outputs(8978) <= a xor b;
    layer0_outputs(8979) <= not a;
    layer0_outputs(8980) <= not (a xor b);
    layer0_outputs(8981) <= not a or b;
    layer0_outputs(8982) <= a or b;
    layer0_outputs(8983) <= not (a or b);
    layer0_outputs(8984) <= b and not a;
    layer0_outputs(8985) <= not (a or b);
    layer0_outputs(8986) <= a and not b;
    layer0_outputs(8987) <= not (a or b);
    layer0_outputs(8988) <= not a;
    layer0_outputs(8989) <= not (a xor b);
    layer0_outputs(8990) <= a or b;
    layer0_outputs(8991) <= a or b;
    layer0_outputs(8992) <= not (a or b);
    layer0_outputs(8993) <= b;
    layer0_outputs(8994) <= b;
    layer0_outputs(8995) <= not b or a;
    layer0_outputs(8996) <= not b;
    layer0_outputs(8997) <= not (a or b);
    layer0_outputs(8998) <= b and not a;
    layer0_outputs(8999) <= a and b;
    layer0_outputs(9000) <= a xor b;
    layer0_outputs(9001) <= b and not a;
    layer0_outputs(9002) <= a;
    layer0_outputs(9003) <= b;
    layer0_outputs(9004) <= a and b;
    layer0_outputs(9005) <= not a or b;
    layer0_outputs(9006) <= not b or a;
    layer0_outputs(9007) <= a xor b;
    layer0_outputs(9008) <= a or b;
    layer0_outputs(9009) <= b and not a;
    layer0_outputs(9010) <= a xor b;
    layer0_outputs(9011) <= a and not b;
    layer0_outputs(9012) <= not (a or b);
    layer0_outputs(9013) <= not (a or b);
    layer0_outputs(9014) <= a;
    layer0_outputs(9015) <= not (a or b);
    layer0_outputs(9016) <= not b or a;
    layer0_outputs(9017) <= b and not a;
    layer0_outputs(9018) <= not (a or b);
    layer0_outputs(9019) <= a and not b;
    layer0_outputs(9020) <= not (a xor b);
    layer0_outputs(9021) <= not (a xor b);
    layer0_outputs(9022) <= not (a or b);
    layer0_outputs(9023) <= a or b;
    layer0_outputs(9024) <= a;
    layer0_outputs(9025) <= not (a or b);
    layer0_outputs(9026) <= b and not a;
    layer0_outputs(9027) <= not (a xor b);
    layer0_outputs(9028) <= a and not b;
    layer0_outputs(9029) <= not (a or b);
    layer0_outputs(9030) <= not (a xor b);
    layer0_outputs(9031) <= a and not b;
    layer0_outputs(9032) <= a xor b;
    layer0_outputs(9033) <= b and not a;
    layer0_outputs(9034) <= a;
    layer0_outputs(9035) <= a and not b;
    layer0_outputs(9036) <= a xor b;
    layer0_outputs(9037) <= a and not b;
    layer0_outputs(9038) <= not (a or b);
    layer0_outputs(9039) <= a and not b;
    layer0_outputs(9040) <= a and b;
    layer0_outputs(9041) <= b and not a;
    layer0_outputs(9042) <= a xor b;
    layer0_outputs(9043) <= not b or a;
    layer0_outputs(9044) <= b and not a;
    layer0_outputs(9045) <= a;
    layer0_outputs(9046) <= not a or b;
    layer0_outputs(9047) <= not a or b;
    layer0_outputs(9048) <= a or b;
    layer0_outputs(9049) <= b and not a;
    layer0_outputs(9050) <= b and not a;
    layer0_outputs(9051) <= a xor b;
    layer0_outputs(9052) <= not (a or b);
    layer0_outputs(9053) <= not a;
    layer0_outputs(9054) <= not a;
    layer0_outputs(9055) <= a and not b;
    layer0_outputs(9056) <= a xor b;
    layer0_outputs(9057) <= not (a or b);
    layer0_outputs(9058) <= a or b;
    layer0_outputs(9059) <= not b or a;
    layer0_outputs(9060) <= b;
    layer0_outputs(9061) <= not (a or b);
    layer0_outputs(9062) <= a and not b;
    layer0_outputs(9063) <= not (a or b);
    layer0_outputs(9064) <= not (a xor b);
    layer0_outputs(9065) <= not b or a;
    layer0_outputs(9066) <= not b;
    layer0_outputs(9067) <= not a;
    layer0_outputs(9068) <= a and not b;
    layer0_outputs(9069) <= a or b;
    layer0_outputs(9070) <= not (a or b);
    layer0_outputs(9071) <= a or b;
    layer0_outputs(9072) <= not (a xor b);
    layer0_outputs(9073) <= '1';
    layer0_outputs(9074) <= a xor b;
    layer0_outputs(9075) <= a xor b;
    layer0_outputs(9076) <= not (a and b);
    layer0_outputs(9077) <= not (a or b);
    layer0_outputs(9078) <= a and b;
    layer0_outputs(9079) <= a;
    layer0_outputs(9080) <= not a;
    layer0_outputs(9081) <= a or b;
    layer0_outputs(9082) <= a and not b;
    layer0_outputs(9083) <= a xor b;
    layer0_outputs(9084) <= not b or a;
    layer0_outputs(9085) <= a or b;
    layer0_outputs(9086) <= not b;
    layer0_outputs(9087) <= not (a or b);
    layer0_outputs(9088) <= b and not a;
    layer0_outputs(9089) <= not a;
    layer0_outputs(9090) <= b and not a;
    layer0_outputs(9091) <= not (a or b);
    layer0_outputs(9092) <= '1';
    layer0_outputs(9093) <= not a or b;
    layer0_outputs(9094) <= b and not a;
    layer0_outputs(9095) <= '1';
    layer0_outputs(9096) <= a or b;
    layer0_outputs(9097) <= not (a or b);
    layer0_outputs(9098) <= not (a or b);
    layer0_outputs(9099) <= b and not a;
    layer0_outputs(9100) <= not (a and b);
    layer0_outputs(9101) <= not (a xor b);
    layer0_outputs(9102) <= not b or a;
    layer0_outputs(9103) <= not b or a;
    layer0_outputs(9104) <= not (a xor b);
    layer0_outputs(9105) <= b;
    layer0_outputs(9106) <= not (a or b);
    layer0_outputs(9107) <= a or b;
    layer0_outputs(9108) <= not (a xor b);
    layer0_outputs(9109) <= a;
    layer0_outputs(9110) <= b and not a;
    layer0_outputs(9111) <= a xor b;
    layer0_outputs(9112) <= a or b;
    layer0_outputs(9113) <= not (a xor b);
    layer0_outputs(9114) <= not a;
    layer0_outputs(9115) <= a xor b;
    layer0_outputs(9116) <= a and not b;
    layer0_outputs(9117) <= not b;
    layer0_outputs(9118) <= not (a xor b);
    layer0_outputs(9119) <= not a;
    layer0_outputs(9120) <= b and not a;
    layer0_outputs(9121) <= b and not a;
    layer0_outputs(9122) <= a and b;
    layer0_outputs(9123) <= a xor b;
    layer0_outputs(9124) <= not b;
    layer0_outputs(9125) <= not b or a;
    layer0_outputs(9126) <= b and not a;
    layer0_outputs(9127) <= a;
    layer0_outputs(9128) <= not (a xor b);
    layer0_outputs(9129) <= not b or a;
    layer0_outputs(9130) <= not b or a;
    layer0_outputs(9131) <= a;
    layer0_outputs(9132) <= not (a or b);
    layer0_outputs(9133) <= not (a xor b);
    layer0_outputs(9134) <= not (a or b);
    layer0_outputs(9135) <= not (a xor b);
    layer0_outputs(9136) <= not (a or b);
    layer0_outputs(9137) <= '0';
    layer0_outputs(9138) <= a or b;
    layer0_outputs(9139) <= not b or a;
    layer0_outputs(9140) <= a and not b;
    layer0_outputs(9141) <= a and not b;
    layer0_outputs(9142) <= not (a xor b);
    layer0_outputs(9143) <= not a;
    layer0_outputs(9144) <= b;
    layer0_outputs(9145) <= not a;
    layer0_outputs(9146) <= not (a or b);
    layer0_outputs(9147) <= not (a or b);
    layer0_outputs(9148) <= a and not b;
    layer0_outputs(9149) <= a and b;
    layer0_outputs(9150) <= '0';
    layer0_outputs(9151) <= not (a or b);
    layer0_outputs(9152) <= a and not b;
    layer0_outputs(9153) <= a and not b;
    layer0_outputs(9154) <= '0';
    layer0_outputs(9155) <= not a or b;
    layer0_outputs(9156) <= b;
    layer0_outputs(9157) <= not b;
    layer0_outputs(9158) <= a and not b;
    layer0_outputs(9159) <= a xor b;
    layer0_outputs(9160) <= not (a or b);
    layer0_outputs(9161) <= a xor b;
    layer0_outputs(9162) <= not b or a;
    layer0_outputs(9163) <= a or b;
    layer0_outputs(9164) <= not (a or b);
    layer0_outputs(9165) <= not a or b;
    layer0_outputs(9166) <= a xor b;
    layer0_outputs(9167) <= b;
    layer0_outputs(9168) <= not (a xor b);
    layer0_outputs(9169) <= not a or b;
    layer0_outputs(9170) <= b;
    layer0_outputs(9171) <= b and not a;
    layer0_outputs(9172) <= not (a xor b);
    layer0_outputs(9173) <= not b or a;
    layer0_outputs(9174) <= b;
    layer0_outputs(9175) <= not b or a;
    layer0_outputs(9176) <= not (a xor b);
    layer0_outputs(9177) <= not a or b;
    layer0_outputs(9178) <= not b or a;
    layer0_outputs(9179) <= a or b;
    layer0_outputs(9180) <= not (a or b);
    layer0_outputs(9181) <= not a;
    layer0_outputs(9182) <= not b;
    layer0_outputs(9183) <= not (a xor b);
    layer0_outputs(9184) <= not (a or b);
    layer0_outputs(9185) <= a or b;
    layer0_outputs(9186) <= not b or a;
    layer0_outputs(9187) <= not (a or b);
    layer0_outputs(9188) <= not (a and b);
    layer0_outputs(9189) <= not b or a;
    layer0_outputs(9190) <= b;
    layer0_outputs(9191) <= a xor b;
    layer0_outputs(9192) <= a or b;
    layer0_outputs(9193) <= not (a xor b);
    layer0_outputs(9194) <= not (a or b);
    layer0_outputs(9195) <= not a;
    layer0_outputs(9196) <= a or b;
    layer0_outputs(9197) <= a;
    layer0_outputs(9198) <= not b;
    layer0_outputs(9199) <= a;
    layer0_outputs(9200) <= a or b;
    layer0_outputs(9201) <= a or b;
    layer0_outputs(9202) <= '0';
    layer0_outputs(9203) <= not a or b;
    layer0_outputs(9204) <= '0';
    layer0_outputs(9205) <= not a;
    layer0_outputs(9206) <= not b;
    layer0_outputs(9207) <= a and not b;
    layer0_outputs(9208) <= not a or b;
    layer0_outputs(9209) <= a or b;
    layer0_outputs(9210) <= a and b;
    layer0_outputs(9211) <= a xor b;
    layer0_outputs(9212) <= not b or a;
    layer0_outputs(9213) <= a or b;
    layer0_outputs(9214) <= not (a and b);
    layer0_outputs(9215) <= not b or a;
    layer0_outputs(9216) <= b;
    layer0_outputs(9217) <= a;
    layer0_outputs(9218) <= a;
    layer0_outputs(9219) <= not (a or b);
    layer0_outputs(9220) <= a and not b;
    layer0_outputs(9221) <= b;
    layer0_outputs(9222) <= not (a xor b);
    layer0_outputs(9223) <= not (a xor b);
    layer0_outputs(9224) <= not a or b;
    layer0_outputs(9225) <= not b or a;
    layer0_outputs(9226) <= not (a or b);
    layer0_outputs(9227) <= not (a or b);
    layer0_outputs(9228) <= a;
    layer0_outputs(9229) <= not b or a;
    layer0_outputs(9230) <= a and not b;
    layer0_outputs(9231) <= a xor b;
    layer0_outputs(9232) <= b and not a;
    layer0_outputs(9233) <= a;
    layer0_outputs(9234) <= '1';
    layer0_outputs(9235) <= a xor b;
    layer0_outputs(9236) <= b and not a;
    layer0_outputs(9237) <= a or b;
    layer0_outputs(9238) <= b;
    layer0_outputs(9239) <= a or b;
    layer0_outputs(9240) <= a or b;
    layer0_outputs(9241) <= a xor b;
    layer0_outputs(9242) <= a or b;
    layer0_outputs(9243) <= not b or a;
    layer0_outputs(9244) <= b;
    layer0_outputs(9245) <= a;
    layer0_outputs(9246) <= not b or a;
    layer0_outputs(9247) <= '0';
    layer0_outputs(9248) <= not (a xor b);
    layer0_outputs(9249) <= not (a or b);
    layer0_outputs(9250) <= not (a xor b);
    layer0_outputs(9251) <= not a or b;
    layer0_outputs(9252) <= not b or a;
    layer0_outputs(9253) <= b;
    layer0_outputs(9254) <= a and not b;
    layer0_outputs(9255) <= a or b;
    layer0_outputs(9256) <= not a or b;
    layer0_outputs(9257) <= a;
    layer0_outputs(9258) <= not b;
    layer0_outputs(9259) <= a xor b;
    layer0_outputs(9260) <= b and not a;
    layer0_outputs(9261) <= not b or a;
    layer0_outputs(9262) <= not (a or b);
    layer0_outputs(9263) <= b and not a;
    layer0_outputs(9264) <= '0';
    layer0_outputs(9265) <= a xor b;
    layer0_outputs(9266) <= not a or b;
    layer0_outputs(9267) <= a xor b;
    layer0_outputs(9268) <= not a;
    layer0_outputs(9269) <= a xor b;
    layer0_outputs(9270) <= a xor b;
    layer0_outputs(9271) <= not b;
    layer0_outputs(9272) <= a and not b;
    layer0_outputs(9273) <= not (a and b);
    layer0_outputs(9274) <= not a or b;
    layer0_outputs(9275) <= b;
    layer0_outputs(9276) <= not b or a;
    layer0_outputs(9277) <= a or b;
    layer0_outputs(9278) <= not (a or b);
    layer0_outputs(9279) <= not b;
    layer0_outputs(9280) <= not b;
    layer0_outputs(9281) <= a;
    layer0_outputs(9282) <= not a;
    layer0_outputs(9283) <= a and not b;
    layer0_outputs(9284) <= a and not b;
    layer0_outputs(9285) <= a xor b;
    layer0_outputs(9286) <= not a or b;
    layer0_outputs(9287) <= not (a or b);
    layer0_outputs(9288) <= not (a xor b);
    layer0_outputs(9289) <= not a or b;
    layer0_outputs(9290) <= not a;
    layer0_outputs(9291) <= a and not b;
    layer0_outputs(9292) <= not (a or b);
    layer0_outputs(9293) <= a xor b;
    layer0_outputs(9294) <= a or b;
    layer0_outputs(9295) <= a or b;
    layer0_outputs(9296) <= a;
    layer0_outputs(9297) <= not a or b;
    layer0_outputs(9298) <= b and not a;
    layer0_outputs(9299) <= a or b;
    layer0_outputs(9300) <= a and not b;
    layer0_outputs(9301) <= a and not b;
    layer0_outputs(9302) <= not a;
    layer0_outputs(9303) <= a xor b;
    layer0_outputs(9304) <= b and not a;
    layer0_outputs(9305) <= not a;
    layer0_outputs(9306) <= not (a or b);
    layer0_outputs(9307) <= a and not b;
    layer0_outputs(9308) <= a xor b;
    layer0_outputs(9309) <= a or b;
    layer0_outputs(9310) <= a and not b;
    layer0_outputs(9311) <= not b or a;
    layer0_outputs(9312) <= not b;
    layer0_outputs(9313) <= not a;
    layer0_outputs(9314) <= not (a or b);
    layer0_outputs(9315) <= '1';
    layer0_outputs(9316) <= not (a or b);
    layer0_outputs(9317) <= not a;
    layer0_outputs(9318) <= not b or a;
    layer0_outputs(9319) <= not (a and b);
    layer0_outputs(9320) <= not b;
    layer0_outputs(9321) <= a and b;
    layer0_outputs(9322) <= not (a or b);
    layer0_outputs(9323) <= a or b;
    layer0_outputs(9324) <= a or b;
    layer0_outputs(9325) <= a;
    layer0_outputs(9326) <= '0';
    layer0_outputs(9327) <= a or b;
    layer0_outputs(9328) <= not (a and b);
    layer0_outputs(9329) <= a or b;
    layer0_outputs(9330) <= not b or a;
    layer0_outputs(9331) <= not (a or b);
    layer0_outputs(9332) <= not b or a;
    layer0_outputs(9333) <= b and not a;
    layer0_outputs(9334) <= not b;
    layer0_outputs(9335) <= not a or b;
    layer0_outputs(9336) <= not b or a;
    layer0_outputs(9337) <= b and not a;
    layer0_outputs(9338) <= not (a or b);
    layer0_outputs(9339) <= b and not a;
    layer0_outputs(9340) <= not b or a;
    layer0_outputs(9341) <= not (a xor b);
    layer0_outputs(9342) <= a xor b;
    layer0_outputs(9343) <= b;
    layer0_outputs(9344) <= not b or a;
    layer0_outputs(9345) <= not a or b;
    layer0_outputs(9346) <= a and b;
    layer0_outputs(9347) <= not b or a;
    layer0_outputs(9348) <= a or b;
    layer0_outputs(9349) <= not b or a;
    layer0_outputs(9350) <= b and not a;
    layer0_outputs(9351) <= not (a or b);
    layer0_outputs(9352) <= not (a or b);
    layer0_outputs(9353) <= not b;
    layer0_outputs(9354) <= not b or a;
    layer0_outputs(9355) <= not b;
    layer0_outputs(9356) <= b and not a;
    layer0_outputs(9357) <= b;
    layer0_outputs(9358) <= not (a and b);
    layer0_outputs(9359) <= not (a or b);
    layer0_outputs(9360) <= a;
    layer0_outputs(9361) <= not (a xor b);
    layer0_outputs(9362) <= a and not b;
    layer0_outputs(9363) <= not b;
    layer0_outputs(9364) <= not (a or b);
    layer0_outputs(9365) <= not a or b;
    layer0_outputs(9366) <= a xor b;
    layer0_outputs(9367) <= not (a xor b);
    layer0_outputs(9368) <= not (a xor b);
    layer0_outputs(9369) <= a;
    layer0_outputs(9370) <= a;
    layer0_outputs(9371) <= not b;
    layer0_outputs(9372) <= b and not a;
    layer0_outputs(9373) <= not (a xor b);
    layer0_outputs(9374) <= a xor b;
    layer0_outputs(9375) <= not a or b;
    layer0_outputs(9376) <= not (a xor b);
    layer0_outputs(9377) <= a and not b;
    layer0_outputs(9378) <= a and b;
    layer0_outputs(9379) <= a or b;
    layer0_outputs(9380) <= '1';
    layer0_outputs(9381) <= a xor b;
    layer0_outputs(9382) <= not a or b;
    layer0_outputs(9383) <= not (a or b);
    layer0_outputs(9384) <= b;
    layer0_outputs(9385) <= not a or b;
    layer0_outputs(9386) <= b;
    layer0_outputs(9387) <= not (a or b);
    layer0_outputs(9388) <= '1';
    layer0_outputs(9389) <= b and not a;
    layer0_outputs(9390) <= not b;
    layer0_outputs(9391) <= not a;
    layer0_outputs(9392) <= a or b;
    layer0_outputs(9393) <= a or b;
    layer0_outputs(9394) <= not (a xor b);
    layer0_outputs(9395) <= not (a or b);
    layer0_outputs(9396) <= not (a xor b);
    layer0_outputs(9397) <= a;
    layer0_outputs(9398) <= a or b;
    layer0_outputs(9399) <= b and not a;
    layer0_outputs(9400) <= '0';
    layer0_outputs(9401) <= b;
    layer0_outputs(9402) <= '0';
    layer0_outputs(9403) <= not (a xor b);
    layer0_outputs(9404) <= not (a xor b);
    layer0_outputs(9405) <= not (a xor b);
    layer0_outputs(9406) <= not (a or b);
    layer0_outputs(9407) <= a or b;
    layer0_outputs(9408) <= not (a and b);
    layer0_outputs(9409) <= a or b;
    layer0_outputs(9410) <= b and not a;
    layer0_outputs(9411) <= not (a or b);
    layer0_outputs(9412) <= not a or b;
    layer0_outputs(9413) <= a;
    layer0_outputs(9414) <= not b or a;
    layer0_outputs(9415) <= a and not b;
    layer0_outputs(9416) <= not b;
    layer0_outputs(9417) <= not (a xor b);
    layer0_outputs(9418) <= not a or b;
    layer0_outputs(9419) <= not a;
    layer0_outputs(9420) <= not (a xor b);
    layer0_outputs(9421) <= a or b;
    layer0_outputs(9422) <= not (a and b);
    layer0_outputs(9423) <= b;
    layer0_outputs(9424) <= a and b;
    layer0_outputs(9425) <= a or b;
    layer0_outputs(9426) <= not a or b;
    layer0_outputs(9427) <= a or b;
    layer0_outputs(9428) <= not a or b;
    layer0_outputs(9429) <= not a;
    layer0_outputs(9430) <= a or b;
    layer0_outputs(9431) <= not a;
    layer0_outputs(9432) <= not b or a;
    layer0_outputs(9433) <= a and not b;
    layer0_outputs(9434) <= a and b;
    layer0_outputs(9435) <= b;
    layer0_outputs(9436) <= a or b;
    layer0_outputs(9437) <= a or b;
    layer0_outputs(9438) <= b;
    layer0_outputs(9439) <= not a or b;
    layer0_outputs(9440) <= b;
    layer0_outputs(9441) <= '0';
    layer0_outputs(9442) <= not a or b;
    layer0_outputs(9443) <= '1';
    layer0_outputs(9444) <= not b or a;
    layer0_outputs(9445) <= a and not b;
    layer0_outputs(9446) <= not a or b;
    layer0_outputs(9447) <= a or b;
    layer0_outputs(9448) <= not b;
    layer0_outputs(9449) <= not b;
    layer0_outputs(9450) <= b;
    layer0_outputs(9451) <= a;
    layer0_outputs(9452) <= a and b;
    layer0_outputs(9453) <= b and not a;
    layer0_outputs(9454) <= a xor b;
    layer0_outputs(9455) <= not (a or b);
    layer0_outputs(9456) <= not (a or b);
    layer0_outputs(9457) <= not (a or b);
    layer0_outputs(9458) <= not a;
    layer0_outputs(9459) <= not a;
    layer0_outputs(9460) <= not (a or b);
    layer0_outputs(9461) <= not b or a;
    layer0_outputs(9462) <= b;
    layer0_outputs(9463) <= not b;
    layer0_outputs(9464) <= a xor b;
    layer0_outputs(9465) <= b and not a;
    layer0_outputs(9466) <= a and b;
    layer0_outputs(9467) <= a xor b;
    layer0_outputs(9468) <= a xor b;
    layer0_outputs(9469) <= not (a or b);
    layer0_outputs(9470) <= a and not b;
    layer0_outputs(9471) <= a and b;
    layer0_outputs(9472) <= b;
    layer0_outputs(9473) <= a or b;
    layer0_outputs(9474) <= not (a or b);
    layer0_outputs(9475) <= not a;
    layer0_outputs(9476) <= a or b;
    layer0_outputs(9477) <= not b or a;
    layer0_outputs(9478) <= not (a or b);
    layer0_outputs(9479) <= b and not a;
    layer0_outputs(9480) <= not (a or b);
    layer0_outputs(9481) <= a and not b;
    layer0_outputs(9482) <= a and not b;
    layer0_outputs(9483) <= a or b;
    layer0_outputs(9484) <= a or b;
    layer0_outputs(9485) <= not a;
    layer0_outputs(9486) <= a or b;
    layer0_outputs(9487) <= not (a or b);
    layer0_outputs(9488) <= a or b;
    layer0_outputs(9489) <= b and not a;
    layer0_outputs(9490) <= not b;
    layer0_outputs(9491) <= not a or b;
    layer0_outputs(9492) <= not (a xor b);
    layer0_outputs(9493) <= b and not a;
    layer0_outputs(9494) <= b and not a;
    layer0_outputs(9495) <= not b;
    layer0_outputs(9496) <= not (a xor b);
    layer0_outputs(9497) <= '1';
    layer0_outputs(9498) <= a or b;
    layer0_outputs(9499) <= a or b;
    layer0_outputs(9500) <= not (a xor b);
    layer0_outputs(9501) <= b and not a;
    layer0_outputs(9502) <= b;
    layer0_outputs(9503) <= b;
    layer0_outputs(9504) <= not (a or b);
    layer0_outputs(9505) <= not (a xor b);
    layer0_outputs(9506) <= not (a or b);
    layer0_outputs(9507) <= not a or b;
    layer0_outputs(9508) <= a xor b;
    layer0_outputs(9509) <= b;
    layer0_outputs(9510) <= not (a or b);
    layer0_outputs(9511) <= a or b;
    layer0_outputs(9512) <= not (a or b);
    layer0_outputs(9513) <= a or b;
    layer0_outputs(9514) <= a and not b;
    layer0_outputs(9515) <= a xor b;
    layer0_outputs(9516) <= not a;
    layer0_outputs(9517) <= not (a or b);
    layer0_outputs(9518) <= a xor b;
    layer0_outputs(9519) <= a xor b;
    layer0_outputs(9520) <= not (a xor b);
    layer0_outputs(9521) <= not a;
    layer0_outputs(9522) <= not b;
    layer0_outputs(9523) <= not (a xor b);
    layer0_outputs(9524) <= not (a xor b);
    layer0_outputs(9525) <= a or b;
    layer0_outputs(9526) <= a and b;
    layer0_outputs(9527) <= a and b;
    layer0_outputs(9528) <= not b or a;
    layer0_outputs(9529) <= a or b;
    layer0_outputs(9530) <= not (a or b);
    layer0_outputs(9531) <= a xor b;
    layer0_outputs(9532) <= not (a or b);
    layer0_outputs(9533) <= not (a xor b);
    layer0_outputs(9534) <= not (a and b);
    layer0_outputs(9535) <= a;
    layer0_outputs(9536) <= b and not a;
    layer0_outputs(9537) <= '0';
    layer0_outputs(9538) <= not (a xor b);
    layer0_outputs(9539) <= not (a or b);
    layer0_outputs(9540) <= not b;
    layer0_outputs(9541) <= a xor b;
    layer0_outputs(9542) <= not b;
    layer0_outputs(9543) <= not (a or b);
    layer0_outputs(9544) <= a xor b;
    layer0_outputs(9545) <= not b;
    layer0_outputs(9546) <= a xor b;
    layer0_outputs(9547) <= not (a xor b);
    layer0_outputs(9548) <= not (a or b);
    layer0_outputs(9549) <= a;
    layer0_outputs(9550) <= not b;
    layer0_outputs(9551) <= not (a xor b);
    layer0_outputs(9552) <= not b;
    layer0_outputs(9553) <= a xor b;
    layer0_outputs(9554) <= not (a xor b);
    layer0_outputs(9555) <= a or b;
    layer0_outputs(9556) <= not b or a;
    layer0_outputs(9557) <= not a;
    layer0_outputs(9558) <= a xor b;
    layer0_outputs(9559) <= not (a xor b);
    layer0_outputs(9560) <= not (a or b);
    layer0_outputs(9561) <= a or b;
    layer0_outputs(9562) <= a;
    layer0_outputs(9563) <= a;
    layer0_outputs(9564) <= not (a xor b);
    layer0_outputs(9565) <= '1';
    layer0_outputs(9566) <= not (a xor b);
    layer0_outputs(9567) <= not (a xor b);
    layer0_outputs(9568) <= not b;
    layer0_outputs(9569) <= a xor b;
    layer0_outputs(9570) <= not (a xor b);
    layer0_outputs(9571) <= a and not b;
    layer0_outputs(9572) <= not b or a;
    layer0_outputs(9573) <= not a;
    layer0_outputs(9574) <= not a or b;
    layer0_outputs(9575) <= not (a and b);
    layer0_outputs(9576) <= b;
    layer0_outputs(9577) <= a or b;
    layer0_outputs(9578) <= b;
    layer0_outputs(9579) <= not (a and b);
    layer0_outputs(9580) <= b;
    layer0_outputs(9581) <= not b or a;
    layer0_outputs(9582) <= a xor b;
    layer0_outputs(9583) <= not (a xor b);
    layer0_outputs(9584) <= a or b;
    layer0_outputs(9585) <= not b;
    layer0_outputs(9586) <= a or b;
    layer0_outputs(9587) <= not b or a;
    layer0_outputs(9588) <= b and not a;
    layer0_outputs(9589) <= not (a xor b);
    layer0_outputs(9590) <= a and not b;
    layer0_outputs(9591) <= not (a or b);
    layer0_outputs(9592) <= a or b;
    layer0_outputs(9593) <= not (a or b);
    layer0_outputs(9594) <= a or b;
    layer0_outputs(9595) <= not (a xor b);
    layer0_outputs(9596) <= not b;
    layer0_outputs(9597) <= '0';
    layer0_outputs(9598) <= not b;
    layer0_outputs(9599) <= not (a or b);
    layer0_outputs(9600) <= a xor b;
    layer0_outputs(9601) <= b and not a;
    layer0_outputs(9602) <= '1';
    layer0_outputs(9603) <= a xor b;
    layer0_outputs(9604) <= not (a xor b);
    layer0_outputs(9605) <= b;
    layer0_outputs(9606) <= not (a xor b);
    layer0_outputs(9607) <= b;
    layer0_outputs(9608) <= not b;
    layer0_outputs(9609) <= a or b;
    layer0_outputs(9610) <= not b or a;
    layer0_outputs(9611) <= '1';
    layer0_outputs(9612) <= not (a xor b);
    layer0_outputs(9613) <= a xor b;
    layer0_outputs(9614) <= not a;
    layer0_outputs(9615) <= a or b;
    layer0_outputs(9616) <= not a;
    layer0_outputs(9617) <= not a;
    layer0_outputs(9618) <= a or b;
    layer0_outputs(9619) <= a xor b;
    layer0_outputs(9620) <= a or b;
    layer0_outputs(9621) <= '1';
    layer0_outputs(9622) <= not a or b;
    layer0_outputs(9623) <= a or b;
    layer0_outputs(9624) <= '0';
    layer0_outputs(9625) <= a xor b;
    layer0_outputs(9626) <= '0';
    layer0_outputs(9627) <= not (a and b);
    layer0_outputs(9628) <= not b;
    layer0_outputs(9629) <= a;
    layer0_outputs(9630) <= '0';
    layer0_outputs(9631) <= a and b;
    layer0_outputs(9632) <= a or b;
    layer0_outputs(9633) <= not (a or b);
    layer0_outputs(9634) <= not a or b;
    layer0_outputs(9635) <= a xor b;
    layer0_outputs(9636) <= a xor b;
    layer0_outputs(9637) <= '1';
    layer0_outputs(9638) <= not (a xor b);
    layer0_outputs(9639) <= not (a and b);
    layer0_outputs(9640) <= not a;
    layer0_outputs(9641) <= b;
    layer0_outputs(9642) <= a and not b;
    layer0_outputs(9643) <= b and not a;
    layer0_outputs(9644) <= not (a or b);
    layer0_outputs(9645) <= a or b;
    layer0_outputs(9646) <= a or b;
    layer0_outputs(9647) <= a or b;
    layer0_outputs(9648) <= a xor b;
    layer0_outputs(9649) <= not (a and b);
    layer0_outputs(9650) <= b and not a;
    layer0_outputs(9651) <= a or b;
    layer0_outputs(9652) <= a or b;
    layer0_outputs(9653) <= a or b;
    layer0_outputs(9654) <= not a;
    layer0_outputs(9655) <= not b or a;
    layer0_outputs(9656) <= a or b;
    layer0_outputs(9657) <= not (a xor b);
    layer0_outputs(9658) <= b;
    layer0_outputs(9659) <= a xor b;
    layer0_outputs(9660) <= not (a xor b);
    layer0_outputs(9661) <= not a;
    layer0_outputs(9662) <= a or b;
    layer0_outputs(9663) <= a and b;
    layer0_outputs(9664) <= a;
    layer0_outputs(9665) <= a or b;
    layer0_outputs(9666) <= b and not a;
    layer0_outputs(9667) <= not (a xor b);
    layer0_outputs(9668) <= not (a xor b);
    layer0_outputs(9669) <= b;
    layer0_outputs(9670) <= not a or b;
    layer0_outputs(9671) <= not a or b;
    layer0_outputs(9672) <= not b;
    layer0_outputs(9673) <= not a;
    layer0_outputs(9674) <= not (a or b);
    layer0_outputs(9675) <= b;
    layer0_outputs(9676) <= not b or a;
    layer0_outputs(9677) <= a or b;
    layer0_outputs(9678) <= '0';
    layer0_outputs(9679) <= not a;
    layer0_outputs(9680) <= a and b;
    layer0_outputs(9681) <= not (a or b);
    layer0_outputs(9682) <= not a or b;
    layer0_outputs(9683) <= not a or b;
    layer0_outputs(9684) <= b and not a;
    layer0_outputs(9685) <= not a;
    layer0_outputs(9686) <= not b;
    layer0_outputs(9687) <= a xor b;
    layer0_outputs(9688) <= a and b;
    layer0_outputs(9689) <= b;
    layer0_outputs(9690) <= a and not b;
    layer0_outputs(9691) <= not (a and b);
    layer0_outputs(9692) <= a and not b;
    layer0_outputs(9693) <= not a or b;
    layer0_outputs(9694) <= not b;
    layer0_outputs(9695) <= not (a or b);
    layer0_outputs(9696) <= a or b;
    layer0_outputs(9697) <= a or b;
    layer0_outputs(9698) <= not (a or b);
    layer0_outputs(9699) <= not a or b;
    layer0_outputs(9700) <= not a;
    layer0_outputs(9701) <= not (a or b);
    layer0_outputs(9702) <= not (a xor b);
    layer0_outputs(9703) <= a;
    layer0_outputs(9704) <= a and b;
    layer0_outputs(9705) <= '1';
    layer0_outputs(9706) <= '1';
    layer0_outputs(9707) <= a xor b;
    layer0_outputs(9708) <= not (a xor b);
    layer0_outputs(9709) <= a and not b;
    layer0_outputs(9710) <= b and not a;
    layer0_outputs(9711) <= not a or b;
    layer0_outputs(9712) <= not b or a;
    layer0_outputs(9713) <= a and b;
    layer0_outputs(9714) <= not b or a;
    layer0_outputs(9715) <= a and not b;
    layer0_outputs(9716) <= a and b;
    layer0_outputs(9717) <= a;
    layer0_outputs(9718) <= not b or a;
    layer0_outputs(9719) <= a and not b;
    layer0_outputs(9720) <= a xor b;
    layer0_outputs(9721) <= a;
    layer0_outputs(9722) <= '0';
    layer0_outputs(9723) <= a or b;
    layer0_outputs(9724) <= not a or b;
    layer0_outputs(9725) <= a xor b;
    layer0_outputs(9726) <= a and not b;
    layer0_outputs(9727) <= not a or b;
    layer0_outputs(9728) <= not (a xor b);
    layer0_outputs(9729) <= a;
    layer0_outputs(9730) <= not (a xor b);
    layer0_outputs(9731) <= a or b;
    layer0_outputs(9732) <= a and not b;
    layer0_outputs(9733) <= not (a or b);
    layer0_outputs(9734) <= b;
    layer0_outputs(9735) <= not a or b;
    layer0_outputs(9736) <= not a or b;
    layer0_outputs(9737) <= not (a and b);
    layer0_outputs(9738) <= a xor b;
    layer0_outputs(9739) <= a or b;
    layer0_outputs(9740) <= a or b;
    layer0_outputs(9741) <= not (a or b);
    layer0_outputs(9742) <= not b;
    layer0_outputs(9743) <= a;
    layer0_outputs(9744) <= not (a xor b);
    layer0_outputs(9745) <= a or b;
    layer0_outputs(9746) <= not (a xor b);
    layer0_outputs(9747) <= not (a xor b);
    layer0_outputs(9748) <= not b;
    layer0_outputs(9749) <= a;
    layer0_outputs(9750) <= not a or b;
    layer0_outputs(9751) <= not b;
    layer0_outputs(9752) <= '0';
    layer0_outputs(9753) <= not (a xor b);
    layer0_outputs(9754) <= not b or a;
    layer0_outputs(9755) <= a;
    layer0_outputs(9756) <= a xor b;
    layer0_outputs(9757) <= a xor b;
    layer0_outputs(9758) <= not (a xor b);
    layer0_outputs(9759) <= not b or a;
    layer0_outputs(9760) <= not (a xor b);
    layer0_outputs(9761) <= a and b;
    layer0_outputs(9762) <= a or b;
    layer0_outputs(9763) <= a xor b;
    layer0_outputs(9764) <= b;
    layer0_outputs(9765) <= '0';
    layer0_outputs(9766) <= not b or a;
    layer0_outputs(9767) <= not a or b;
    layer0_outputs(9768) <= not b or a;
    layer0_outputs(9769) <= a or b;
    layer0_outputs(9770) <= not a or b;
    layer0_outputs(9771) <= not (a or b);
    layer0_outputs(9772) <= a and not b;
    layer0_outputs(9773) <= a xor b;
    layer0_outputs(9774) <= not (a or b);
    layer0_outputs(9775) <= not (a xor b);
    layer0_outputs(9776) <= a or b;
    layer0_outputs(9777) <= a or b;
    layer0_outputs(9778) <= b and not a;
    layer0_outputs(9779) <= '1';
    layer0_outputs(9780) <= not b or a;
    layer0_outputs(9781) <= a xor b;
    layer0_outputs(9782) <= not (a or b);
    layer0_outputs(9783) <= a xor b;
    layer0_outputs(9784) <= not (a xor b);
    layer0_outputs(9785) <= a;
    layer0_outputs(9786) <= not b or a;
    layer0_outputs(9787) <= a or b;
    layer0_outputs(9788) <= a or b;
    layer0_outputs(9789) <= a and not b;
    layer0_outputs(9790) <= a or b;
    layer0_outputs(9791) <= not b or a;
    layer0_outputs(9792) <= a and b;
    layer0_outputs(9793) <= not (a and b);
    layer0_outputs(9794) <= not b;
    layer0_outputs(9795) <= a or b;
    layer0_outputs(9796) <= not b or a;
    layer0_outputs(9797) <= b;
    layer0_outputs(9798) <= b and not a;
    layer0_outputs(9799) <= b and not a;
    layer0_outputs(9800) <= a xor b;
    layer0_outputs(9801) <= a or b;
    layer0_outputs(9802) <= a and not b;
    layer0_outputs(9803) <= not (a or b);
    layer0_outputs(9804) <= not (a or b);
    layer0_outputs(9805) <= b and not a;
    layer0_outputs(9806) <= not b;
    layer0_outputs(9807) <= not a;
    layer0_outputs(9808) <= not b;
    layer0_outputs(9809) <= a and not b;
    layer0_outputs(9810) <= a xor b;
    layer0_outputs(9811) <= a and not b;
    layer0_outputs(9812) <= not (a and b);
    layer0_outputs(9813) <= a and not b;
    layer0_outputs(9814) <= not (a xor b);
    layer0_outputs(9815) <= a xor b;
    layer0_outputs(9816) <= not (a xor b);
    layer0_outputs(9817) <= a and not b;
    layer0_outputs(9818) <= not (a xor b);
    layer0_outputs(9819) <= b;
    layer0_outputs(9820) <= b;
    layer0_outputs(9821) <= not (a or b);
    layer0_outputs(9822) <= not b;
    layer0_outputs(9823) <= b;
    layer0_outputs(9824) <= not (a xor b);
    layer0_outputs(9825) <= '1';
    layer0_outputs(9826) <= b;
    layer0_outputs(9827) <= not a or b;
    layer0_outputs(9828) <= b and not a;
    layer0_outputs(9829) <= not (a xor b);
    layer0_outputs(9830) <= not b or a;
    layer0_outputs(9831) <= not (a or b);
    layer0_outputs(9832) <= a or b;
    layer0_outputs(9833) <= b;
    layer0_outputs(9834) <= not a;
    layer0_outputs(9835) <= not a or b;
    layer0_outputs(9836) <= not a or b;
    layer0_outputs(9837) <= a;
    layer0_outputs(9838) <= b and not a;
    layer0_outputs(9839) <= a and not b;
    layer0_outputs(9840) <= a or b;
    layer0_outputs(9841) <= not (a xor b);
    layer0_outputs(9842) <= not a or b;
    layer0_outputs(9843) <= b;
    layer0_outputs(9844) <= a;
    layer0_outputs(9845) <= a xor b;
    layer0_outputs(9846) <= a xor b;
    layer0_outputs(9847) <= a xor b;
    layer0_outputs(9848) <= a;
    layer0_outputs(9849) <= not b or a;
    layer0_outputs(9850) <= not b or a;
    layer0_outputs(9851) <= a xor b;
    layer0_outputs(9852) <= not (a or b);
    layer0_outputs(9853) <= not b or a;
    layer0_outputs(9854) <= not a or b;
    layer0_outputs(9855) <= a or b;
    layer0_outputs(9856) <= not a;
    layer0_outputs(9857) <= not (a or b);
    layer0_outputs(9858) <= not b;
    layer0_outputs(9859) <= not (a xor b);
    layer0_outputs(9860) <= a;
    layer0_outputs(9861) <= a;
    layer0_outputs(9862) <= not (a xor b);
    layer0_outputs(9863) <= not a or b;
    layer0_outputs(9864) <= a xor b;
    layer0_outputs(9865) <= not (a or b);
    layer0_outputs(9866) <= not (a or b);
    layer0_outputs(9867) <= not (a or b);
    layer0_outputs(9868) <= not b;
    layer0_outputs(9869) <= a or b;
    layer0_outputs(9870) <= not b or a;
    layer0_outputs(9871) <= a xor b;
    layer0_outputs(9872) <= not b or a;
    layer0_outputs(9873) <= a and not b;
    layer0_outputs(9874) <= '0';
    layer0_outputs(9875) <= not b;
    layer0_outputs(9876) <= a xor b;
    layer0_outputs(9877) <= a or b;
    layer0_outputs(9878) <= not a or b;
    layer0_outputs(9879) <= not (a or b);
    layer0_outputs(9880) <= not (a or b);
    layer0_outputs(9881) <= a or b;
    layer0_outputs(9882) <= b;
    layer0_outputs(9883) <= not b or a;
    layer0_outputs(9884) <= not b or a;
    layer0_outputs(9885) <= not a or b;
    layer0_outputs(9886) <= not b or a;
    layer0_outputs(9887) <= not a;
    layer0_outputs(9888) <= a or b;
    layer0_outputs(9889) <= b;
    layer0_outputs(9890) <= b;
    layer0_outputs(9891) <= not (a xor b);
    layer0_outputs(9892) <= not a;
    layer0_outputs(9893) <= '1';
    layer0_outputs(9894) <= a;
    layer0_outputs(9895) <= '1';
    layer0_outputs(9896) <= not (a xor b);
    layer0_outputs(9897) <= a xor b;
    layer0_outputs(9898) <= not b or a;
    layer0_outputs(9899) <= not (a or b);
    layer0_outputs(9900) <= not b or a;
    layer0_outputs(9901) <= not a or b;
    layer0_outputs(9902) <= not a;
    layer0_outputs(9903) <= a xor b;
    layer0_outputs(9904) <= a or b;
    layer0_outputs(9905) <= a or b;
    layer0_outputs(9906) <= a or b;
    layer0_outputs(9907) <= a xor b;
    layer0_outputs(9908) <= a or b;
    layer0_outputs(9909) <= b and not a;
    layer0_outputs(9910) <= not b or a;
    layer0_outputs(9911) <= not a or b;
    layer0_outputs(9912) <= b and not a;
    layer0_outputs(9913) <= not (a xor b);
    layer0_outputs(9914) <= not (a xor b);
    layer0_outputs(9915) <= b and not a;
    layer0_outputs(9916) <= not a or b;
    layer0_outputs(9917) <= not (a or b);
    layer0_outputs(9918) <= a and b;
    layer0_outputs(9919) <= not b;
    layer0_outputs(9920) <= not (a or b);
    layer0_outputs(9921) <= a xor b;
    layer0_outputs(9922) <= a xor b;
    layer0_outputs(9923) <= not (a and b);
    layer0_outputs(9924) <= b and not a;
    layer0_outputs(9925) <= a or b;
    layer0_outputs(9926) <= a or b;
    layer0_outputs(9927) <= a or b;
    layer0_outputs(9928) <= a xor b;
    layer0_outputs(9929) <= not (a xor b);
    layer0_outputs(9930) <= b;
    layer0_outputs(9931) <= not (a or b);
    layer0_outputs(9932) <= not a or b;
    layer0_outputs(9933) <= not b or a;
    layer0_outputs(9934) <= not (a or b);
    layer0_outputs(9935) <= a xor b;
    layer0_outputs(9936) <= not (a or b);
    layer0_outputs(9937) <= a or b;
    layer0_outputs(9938) <= a;
    layer0_outputs(9939) <= not b;
    layer0_outputs(9940) <= a;
    layer0_outputs(9941) <= not a;
    layer0_outputs(9942) <= not b or a;
    layer0_outputs(9943) <= b and not a;
    layer0_outputs(9944) <= not a;
    layer0_outputs(9945) <= a or b;
    layer0_outputs(9946) <= not (a or b);
    layer0_outputs(9947) <= '1';
    layer0_outputs(9948) <= not a;
    layer0_outputs(9949) <= not a or b;
    layer0_outputs(9950) <= not (a xor b);
    layer0_outputs(9951) <= not b or a;
    layer0_outputs(9952) <= b and not a;
    layer0_outputs(9953) <= b and not a;
    layer0_outputs(9954) <= b;
    layer0_outputs(9955) <= a xor b;
    layer0_outputs(9956) <= not (a xor b);
    layer0_outputs(9957) <= b;
    layer0_outputs(9958) <= not (a or b);
    layer0_outputs(9959) <= a xor b;
    layer0_outputs(9960) <= not b;
    layer0_outputs(9961) <= a xor b;
    layer0_outputs(9962) <= not a or b;
    layer0_outputs(9963) <= a or b;
    layer0_outputs(9964) <= not a or b;
    layer0_outputs(9965) <= not (a xor b);
    layer0_outputs(9966) <= b;
    layer0_outputs(9967) <= not (a xor b);
    layer0_outputs(9968) <= not a or b;
    layer0_outputs(9969) <= not b;
    layer0_outputs(9970) <= a or b;
    layer0_outputs(9971) <= not b or a;
    layer0_outputs(9972) <= not a;
    layer0_outputs(9973) <= not a;
    layer0_outputs(9974) <= not (a or b);
    layer0_outputs(9975) <= b and not a;
    layer0_outputs(9976) <= not b;
    layer0_outputs(9977) <= a and b;
    layer0_outputs(9978) <= not a or b;
    layer0_outputs(9979) <= not (a or b);
    layer0_outputs(9980) <= a or b;
    layer0_outputs(9981) <= '0';
    layer0_outputs(9982) <= a and not b;
    layer0_outputs(9983) <= not (a and b);
    layer0_outputs(9984) <= not (a or b);
    layer0_outputs(9985) <= a and not b;
    layer0_outputs(9986) <= b and not a;
    layer0_outputs(9987) <= a and b;
    layer0_outputs(9988) <= not (a or b);
    layer0_outputs(9989) <= not b or a;
    layer0_outputs(9990) <= not a or b;
    layer0_outputs(9991) <= not (a or b);
    layer0_outputs(9992) <= b and not a;
    layer0_outputs(9993) <= '1';
    layer0_outputs(9994) <= a;
    layer0_outputs(9995) <= a xor b;
    layer0_outputs(9996) <= a or b;
    layer0_outputs(9997) <= a or b;
    layer0_outputs(9998) <= a and b;
    layer0_outputs(9999) <= not b;
    layer0_outputs(10000) <= b;
    layer0_outputs(10001) <= a and not b;
    layer0_outputs(10002) <= not a;
    layer0_outputs(10003) <= not (a xor b);
    layer0_outputs(10004) <= not (a or b);
    layer0_outputs(10005) <= not (a or b);
    layer0_outputs(10006) <= not (a or b);
    layer0_outputs(10007) <= not (a and b);
    layer0_outputs(10008) <= a or b;
    layer0_outputs(10009) <= a xor b;
    layer0_outputs(10010) <= not a;
    layer0_outputs(10011) <= not a or b;
    layer0_outputs(10012) <= not (a or b);
    layer0_outputs(10013) <= not b;
    layer0_outputs(10014) <= not (a or b);
    layer0_outputs(10015) <= not a or b;
    layer0_outputs(10016) <= not a;
    layer0_outputs(10017) <= not (a xor b);
    layer0_outputs(10018) <= a and not b;
    layer0_outputs(10019) <= b;
    layer0_outputs(10020) <= not (a or b);
    layer0_outputs(10021) <= b and not a;
    layer0_outputs(10022) <= a xor b;
    layer0_outputs(10023) <= a and b;
    layer0_outputs(10024) <= a and b;
    layer0_outputs(10025) <= a;
    layer0_outputs(10026) <= not b;
    layer0_outputs(10027) <= b and not a;
    layer0_outputs(10028) <= '0';
    layer0_outputs(10029) <= not (a xor b);
    layer0_outputs(10030) <= a xor b;
    layer0_outputs(10031) <= a or b;
    layer0_outputs(10032) <= not (a xor b);
    layer0_outputs(10033) <= not (a xor b);
    layer0_outputs(10034) <= b;
    layer0_outputs(10035) <= a or b;
    layer0_outputs(10036) <= a;
    layer0_outputs(10037) <= not (a xor b);
    layer0_outputs(10038) <= b;
    layer0_outputs(10039) <= not a or b;
    layer0_outputs(10040) <= a or b;
    layer0_outputs(10041) <= a and b;
    layer0_outputs(10042) <= b;
    layer0_outputs(10043) <= not (a xor b);
    layer0_outputs(10044) <= b and not a;
    layer0_outputs(10045) <= a xor b;
    layer0_outputs(10046) <= b and not a;
    layer0_outputs(10047) <= not a;
    layer0_outputs(10048) <= not b;
    layer0_outputs(10049) <= b;
    layer0_outputs(10050) <= a and not b;
    layer0_outputs(10051) <= a or b;
    layer0_outputs(10052) <= not (a or b);
    layer0_outputs(10053) <= a and not b;
    layer0_outputs(10054) <= not b or a;
    layer0_outputs(10055) <= b and not a;
    layer0_outputs(10056) <= a or b;
    layer0_outputs(10057) <= a xor b;
    layer0_outputs(10058) <= not b;
    layer0_outputs(10059) <= a xor b;
    layer0_outputs(10060) <= a xor b;
    layer0_outputs(10061) <= not (a or b);
    layer0_outputs(10062) <= a or b;
    layer0_outputs(10063) <= a and b;
    layer0_outputs(10064) <= b;
    layer0_outputs(10065) <= a or b;
    layer0_outputs(10066) <= a or b;
    layer0_outputs(10067) <= not (a or b);
    layer0_outputs(10068) <= not (a xor b);
    layer0_outputs(10069) <= not b or a;
    layer0_outputs(10070) <= a xor b;
    layer0_outputs(10071) <= not b or a;
    layer0_outputs(10072) <= not a or b;
    layer0_outputs(10073) <= a and not b;
    layer0_outputs(10074) <= a and not b;
    layer0_outputs(10075) <= a and b;
    layer0_outputs(10076) <= b;
    layer0_outputs(10077) <= a;
    layer0_outputs(10078) <= b;
    layer0_outputs(10079) <= a;
    layer0_outputs(10080) <= not b;
    layer0_outputs(10081) <= not a or b;
    layer0_outputs(10082) <= not (a xor b);
    layer0_outputs(10083) <= a xor b;
    layer0_outputs(10084) <= a xor b;
    layer0_outputs(10085) <= a and not b;
    layer0_outputs(10086) <= not a;
    layer0_outputs(10087) <= not b;
    layer0_outputs(10088) <= not (a xor b);
    layer0_outputs(10089) <= not (a or b);
    layer0_outputs(10090) <= b and not a;
    layer0_outputs(10091) <= not b;
    layer0_outputs(10092) <= not (a xor b);
    layer0_outputs(10093) <= a xor b;
    layer0_outputs(10094) <= a;
    layer0_outputs(10095) <= not (a xor b);
    layer0_outputs(10096) <= a xor b;
    layer0_outputs(10097) <= b;
    layer0_outputs(10098) <= a;
    layer0_outputs(10099) <= b;
    layer0_outputs(10100) <= b;
    layer0_outputs(10101) <= b;
    layer0_outputs(10102) <= a or b;
    layer0_outputs(10103) <= a or b;
    layer0_outputs(10104) <= not (a or b);
    layer0_outputs(10105) <= not a or b;
    layer0_outputs(10106) <= not (a xor b);
    layer0_outputs(10107) <= b;
    layer0_outputs(10108) <= a or b;
    layer0_outputs(10109) <= b;
    layer0_outputs(10110) <= a and b;
    layer0_outputs(10111) <= not a or b;
    layer0_outputs(10112) <= not b or a;
    layer0_outputs(10113) <= a or b;
    layer0_outputs(10114) <= not a or b;
    layer0_outputs(10115) <= b and not a;
    layer0_outputs(10116) <= a or b;
    layer0_outputs(10117) <= a or b;
    layer0_outputs(10118) <= '1';
    layer0_outputs(10119) <= '0';
    layer0_outputs(10120) <= '1';
    layer0_outputs(10121) <= b;
    layer0_outputs(10122) <= not (a xor b);
    layer0_outputs(10123) <= a and not b;
    layer0_outputs(10124) <= a or b;
    layer0_outputs(10125) <= not (a or b);
    layer0_outputs(10126) <= not (a or b);
    layer0_outputs(10127) <= not a or b;
    layer0_outputs(10128) <= not (a and b);
    layer0_outputs(10129) <= '1';
    layer0_outputs(10130) <= a and not b;
    layer0_outputs(10131) <= a and not b;
    layer0_outputs(10132) <= not (a or b);
    layer0_outputs(10133) <= '1';
    layer0_outputs(10134) <= not a or b;
    layer0_outputs(10135) <= not (a xor b);
    layer0_outputs(10136) <= a or b;
    layer0_outputs(10137) <= a or b;
    layer0_outputs(10138) <= not (a or b);
    layer0_outputs(10139) <= not b or a;
    layer0_outputs(10140) <= not (a and b);
    layer0_outputs(10141) <= a;
    layer0_outputs(10142) <= b and not a;
    layer0_outputs(10143) <= not a or b;
    layer0_outputs(10144) <= a or b;
    layer0_outputs(10145) <= a xor b;
    layer0_outputs(10146) <= b;
    layer0_outputs(10147) <= b and not a;
    layer0_outputs(10148) <= not (a or b);
    layer0_outputs(10149) <= a or b;
    layer0_outputs(10150) <= not (a xor b);
    layer0_outputs(10151) <= not a;
    layer0_outputs(10152) <= not b or a;
    layer0_outputs(10153) <= a;
    layer0_outputs(10154) <= a xor b;
    layer0_outputs(10155) <= a;
    layer0_outputs(10156) <= a or b;
    layer0_outputs(10157) <= a xor b;
    layer0_outputs(10158) <= not (a xor b);
    layer0_outputs(10159) <= not b;
    layer0_outputs(10160) <= not b or a;
    layer0_outputs(10161) <= not b or a;
    layer0_outputs(10162) <= a or b;
    layer0_outputs(10163) <= not a;
    layer0_outputs(10164) <= a;
    layer0_outputs(10165) <= a or b;
    layer0_outputs(10166) <= not (a xor b);
    layer0_outputs(10167) <= a or b;
    layer0_outputs(10168) <= not (a or b);
    layer0_outputs(10169) <= not (a xor b);
    layer0_outputs(10170) <= not (a xor b);
    layer0_outputs(10171) <= not b;
    layer0_outputs(10172) <= a;
    layer0_outputs(10173) <= not (a and b);
    layer0_outputs(10174) <= a or b;
    layer0_outputs(10175) <= a and not b;
    layer0_outputs(10176) <= not (a or b);
    layer0_outputs(10177) <= a and not b;
    layer0_outputs(10178) <= '1';
    layer0_outputs(10179) <= b;
    layer0_outputs(10180) <= b;
    layer0_outputs(10181) <= not b or a;
    layer0_outputs(10182) <= a or b;
    layer0_outputs(10183) <= a xor b;
    layer0_outputs(10184) <= not b;
    layer0_outputs(10185) <= a or b;
    layer0_outputs(10186) <= b and not a;
    layer0_outputs(10187) <= not (a or b);
    layer0_outputs(10188) <= a or b;
    layer0_outputs(10189) <= not (a xor b);
    layer0_outputs(10190) <= not a or b;
    layer0_outputs(10191) <= a xor b;
    layer0_outputs(10192) <= a or b;
    layer0_outputs(10193) <= not a or b;
    layer0_outputs(10194) <= not (a or b);
    layer0_outputs(10195) <= b;
    layer0_outputs(10196) <= a or b;
    layer0_outputs(10197) <= not b or a;
    layer0_outputs(10198) <= not (a xor b);
    layer0_outputs(10199) <= not a;
    layer0_outputs(10200) <= a;
    layer0_outputs(10201) <= '1';
    layer0_outputs(10202) <= a and not b;
    layer0_outputs(10203) <= b and not a;
    layer0_outputs(10204) <= a and b;
    layer0_outputs(10205) <= not a or b;
    layer0_outputs(10206) <= a or b;
    layer0_outputs(10207) <= a xor b;
    layer0_outputs(10208) <= not b or a;
    layer0_outputs(10209) <= not b or a;
    layer0_outputs(10210) <= b and not a;
    layer0_outputs(10211) <= a xor b;
    layer0_outputs(10212) <= '0';
    layer0_outputs(10213) <= not a;
    layer0_outputs(10214) <= not a;
    layer0_outputs(10215) <= not b or a;
    layer0_outputs(10216) <= a or b;
    layer0_outputs(10217) <= not (a or b);
    layer0_outputs(10218) <= a;
    layer0_outputs(10219) <= a xor b;
    layer0_outputs(10220) <= not a;
    layer0_outputs(10221) <= a xor b;
    layer0_outputs(10222) <= b;
    layer0_outputs(10223) <= not (a or b);
    layer0_outputs(10224) <= a or b;
    layer0_outputs(10225) <= a or b;
    layer0_outputs(10226) <= b and not a;
    layer0_outputs(10227) <= a xor b;
    layer0_outputs(10228) <= a or b;
    layer0_outputs(10229) <= a and not b;
    layer0_outputs(10230) <= not (a and b);
    layer0_outputs(10231) <= not (a xor b);
    layer0_outputs(10232) <= b;
    layer0_outputs(10233) <= not (a xor b);
    layer0_outputs(10234) <= a xor b;
    layer0_outputs(10235) <= '0';
    layer0_outputs(10236) <= not a;
    layer0_outputs(10237) <= b;
    layer0_outputs(10238) <= b and not a;
    layer0_outputs(10239) <= not (a xor b);
    outputs(0) <= a and not b;
    outputs(1) <= a;
    outputs(2) <= b;
    outputs(3) <= b and not a;
    outputs(4) <= not b;
    outputs(5) <= not (a xor b);
    outputs(6) <= not (a xor b);
    outputs(7) <= a;
    outputs(8) <= not a;
    outputs(9) <= a xor b;
    outputs(10) <= not (a xor b);
    outputs(11) <= a and not b;
    outputs(12) <= a xor b;
    outputs(13) <= b;
    outputs(14) <= b;
    outputs(15) <= b;
    outputs(16) <= a;
    outputs(17) <= a;
    outputs(18) <= not a;
    outputs(19) <= b;
    outputs(20) <= not b or a;
    outputs(21) <= b and not a;
    outputs(22) <= a xor b;
    outputs(23) <= a;
    outputs(24) <= a and b;
    outputs(25) <= b and not a;
    outputs(26) <= not a or b;
    outputs(27) <= not a or b;
    outputs(28) <= b;
    outputs(29) <= a;
    outputs(30) <= a or b;
    outputs(31) <= b and not a;
    outputs(32) <= not a;
    outputs(33) <= not (a xor b);
    outputs(34) <= a or b;
    outputs(35) <= a and not b;
    outputs(36) <= not (a xor b);
    outputs(37) <= b and not a;
    outputs(38) <= a xor b;
    outputs(39) <= not b;
    outputs(40) <= b;
    outputs(41) <= b;
    outputs(42) <= not a;
    outputs(43) <= a;
    outputs(44) <= a or b;
    outputs(45) <= a or b;
    outputs(46) <= not (a xor b);
    outputs(47) <= not b;
    outputs(48) <= not b or a;
    outputs(49) <= not (a and b);
    outputs(50) <= not a;
    outputs(51) <= not (a xor b);
    outputs(52) <= a and b;
    outputs(53) <= not (a or b);
    outputs(54) <= a and b;
    outputs(55) <= b and not a;
    outputs(56) <= b;
    outputs(57) <= not b;
    outputs(58) <= b and not a;
    outputs(59) <= b and not a;
    outputs(60) <= b and not a;
    outputs(61) <= not a;
    outputs(62) <= not (a xor b);
    outputs(63) <= a;
    outputs(64) <= a;
    outputs(65) <= not (a or b);
    outputs(66) <= not a;
    outputs(67) <= not b;
    outputs(68) <= a and not b;
    outputs(69) <= not b;
    outputs(70) <= not (a xor b);
    outputs(71) <= not (a and b);
    outputs(72) <= b;
    outputs(73) <= b and not a;
    outputs(74) <= not b;
    outputs(75) <= a;
    outputs(76) <= not a;
    outputs(77) <= not (a xor b);
    outputs(78) <= a and b;
    outputs(79) <= not a;
    outputs(80) <= not a;
    outputs(81) <= not (a xor b);
    outputs(82) <= not a;
    outputs(83) <= b;
    outputs(84) <= not b;
    outputs(85) <= a xor b;
    outputs(86) <= a xor b;
    outputs(87) <= a;
    outputs(88) <= b;
    outputs(89) <= b;
    outputs(90) <= not a;
    outputs(91) <= a xor b;
    outputs(92) <= a xor b;
    outputs(93) <= a and b;
    outputs(94) <= not (a xor b);
    outputs(95) <= not b;
    outputs(96) <= a and not b;
    outputs(97) <= not b;
    outputs(98) <= a xor b;
    outputs(99) <= not a;
    outputs(100) <= not b;
    outputs(101) <= b;
    outputs(102) <= a;
    outputs(103) <= not (a xor b);
    outputs(104) <= a and not b;
    outputs(105) <= a;
    outputs(106) <= a and b;
    outputs(107) <= not (a and b);
    outputs(108) <= a xor b;
    outputs(109) <= a xor b;
    outputs(110) <= not (a xor b);
    outputs(111) <= not (a or b);
    outputs(112) <= a or b;
    outputs(113) <= not (a xor b);
    outputs(114) <= b and not a;
    outputs(115) <= not (a xor b);
    outputs(116) <= not (a xor b);
    outputs(117) <= not b or a;
    outputs(118) <= b;
    outputs(119) <= b;
    outputs(120) <= not (a or b);
    outputs(121) <= a and not b;
    outputs(122) <= a xor b;
    outputs(123) <= a;
    outputs(124) <= a and not b;
    outputs(125) <= not (a xor b);
    outputs(126) <= a xor b;
    outputs(127) <= b and not a;
    outputs(128) <= b;
    outputs(129) <= not a;
    outputs(130) <= a xor b;
    outputs(131) <= b;
    outputs(132) <= not b;
    outputs(133) <= a;
    outputs(134) <= b;
    outputs(135) <= a xor b;
    outputs(136) <= not a;
    outputs(137) <= a;
    outputs(138) <= not a;
    outputs(139) <= not b;
    outputs(140) <= not (a xor b);
    outputs(141) <= b;
    outputs(142) <= a xor b;
    outputs(143) <= b and not a;
    outputs(144) <= not b;
    outputs(145) <= b;
    outputs(146) <= not a;
    outputs(147) <= a xor b;
    outputs(148) <= a;
    outputs(149) <= b and not a;
    outputs(150) <= not a;
    outputs(151) <= not (a xor b);
    outputs(152) <= a and b;
    outputs(153) <= not b;
    outputs(154) <= a and not b;
    outputs(155) <= not a;
    outputs(156) <= a or b;
    outputs(157) <= a;
    outputs(158) <= a xor b;
    outputs(159) <= a xor b;
    outputs(160) <= not a;
    outputs(161) <= not b or a;
    outputs(162) <= not (a and b);
    outputs(163) <= b;
    outputs(164) <= not b;
    outputs(165) <= a xor b;
    outputs(166) <= a xor b;
    outputs(167) <= not (a xor b);
    outputs(168) <= a;
    outputs(169) <= a xor b;
    outputs(170) <= not b;
    outputs(171) <= not (a xor b);
    outputs(172) <= a and not b;
    outputs(173) <= not a or b;
    outputs(174) <= not b;
    outputs(175) <= not (a xor b);
    outputs(176) <= not a;
    outputs(177) <= not a or b;
    outputs(178) <= b;
    outputs(179) <= not (a xor b);
    outputs(180) <= not b;
    outputs(181) <= a;
    outputs(182) <= not a;
    outputs(183) <= not b;
    outputs(184) <= a;
    outputs(185) <= a xor b;
    outputs(186) <= a;
    outputs(187) <= a;
    outputs(188) <= not a;
    outputs(189) <= a;
    outputs(190) <= not (a xor b);
    outputs(191) <= not b;
    outputs(192) <= b and not a;
    outputs(193) <= not a;
    outputs(194) <= a xor b;
    outputs(195) <= a xor b;
    outputs(196) <= not (a xor b);
    outputs(197) <= not b;
    outputs(198) <= b;
    outputs(199) <= not (a xor b);
    outputs(200) <= a xor b;
    outputs(201) <= a;
    outputs(202) <= not (a or b);
    outputs(203) <= a;
    outputs(204) <= b;
    outputs(205) <= not b or a;
    outputs(206) <= not (a xor b);
    outputs(207) <= b;
    outputs(208) <= not a or b;
    outputs(209) <= b;
    outputs(210) <= b;
    outputs(211) <= a;
    outputs(212) <= a;
    outputs(213) <= a xor b;
    outputs(214) <= not b;
    outputs(215) <= b;
    outputs(216) <= not a;
    outputs(217) <= b;
    outputs(218) <= not (a and b);
    outputs(219) <= not (a xor b);
    outputs(220) <= a and b;
    outputs(221) <= not b;
    outputs(222) <= a xor b;
    outputs(223) <= a and not b;
    outputs(224) <= a or b;
    outputs(225) <= b;
    outputs(226) <= a xor b;
    outputs(227) <= b;
    outputs(228) <= a or b;
    outputs(229) <= a and b;
    outputs(230) <= not b;
    outputs(231) <= not b;
    outputs(232) <= not (a xor b);
    outputs(233) <= b;
    outputs(234) <= not a;
    outputs(235) <= not b;
    outputs(236) <= not a;
    outputs(237) <= not (a xor b);
    outputs(238) <= a xor b;
    outputs(239) <= not b or a;
    outputs(240) <= a and b;
    outputs(241) <= not (a and b);
    outputs(242) <= not a;
    outputs(243) <= b;
    outputs(244) <= a;
    outputs(245) <= not (a or b);
    outputs(246) <= not b;
    outputs(247) <= b and not a;
    outputs(248) <= not a;
    outputs(249) <= b;
    outputs(250) <= b;
    outputs(251) <= not (a xor b);
    outputs(252) <= not (a or b);
    outputs(253) <= not a;
    outputs(254) <= not (a xor b);
    outputs(255) <= not b;
    outputs(256) <= a and not b;
    outputs(257) <= a xor b;
    outputs(258) <= a xor b;
    outputs(259) <= a and not b;
    outputs(260) <= not (a and b);
    outputs(261) <= not a;
    outputs(262) <= a;
    outputs(263) <= not a;
    outputs(264) <= b;
    outputs(265) <= not (a or b);
    outputs(266) <= not a;
    outputs(267) <= a or b;
    outputs(268) <= a and b;
    outputs(269) <= not b;
    outputs(270) <= not a;
    outputs(271) <= not b or a;
    outputs(272) <= not a;
    outputs(273) <= a xor b;
    outputs(274) <= a;
    outputs(275) <= not (a or b);
    outputs(276) <= not (a or b);
    outputs(277) <= not b;
    outputs(278) <= not (a and b);
    outputs(279) <= not b;
    outputs(280) <= a;
    outputs(281) <= a xor b;
    outputs(282) <= not a;
    outputs(283) <= not (a and b);
    outputs(284) <= a xor b;
    outputs(285) <= not (a xor b);
    outputs(286) <= not b;
    outputs(287) <= not (a xor b);
    outputs(288) <= not b;
    outputs(289) <= not a;
    outputs(290) <= b and not a;
    outputs(291) <= b;
    outputs(292) <= not b;
    outputs(293) <= not b;
    outputs(294) <= not b;
    outputs(295) <= b;
    outputs(296) <= a xor b;
    outputs(297) <= not a;
    outputs(298) <= not (a xor b);
    outputs(299) <= a and not b;
    outputs(300) <= a;
    outputs(301) <= not (a xor b);
    outputs(302) <= a;
    outputs(303) <= b;
    outputs(304) <= not a;
    outputs(305) <= not a;
    outputs(306) <= b;
    outputs(307) <= not a;
    outputs(308) <= not (a xor b);
    outputs(309) <= not a;
    outputs(310) <= b;
    outputs(311) <= a;
    outputs(312) <= not a;
    outputs(313) <= b;
    outputs(314) <= not b;
    outputs(315) <= not (a or b);
    outputs(316) <= not b;
    outputs(317) <= not (a and b);
    outputs(318) <= not b;
    outputs(319) <= b and not a;
    outputs(320) <= a and not b;
    outputs(321) <= b;
    outputs(322) <= b;
    outputs(323) <= a xor b;
    outputs(324) <= not a;
    outputs(325) <= a and not b;
    outputs(326) <= not a;
    outputs(327) <= not (a xor b);
    outputs(328) <= not (a and b);
    outputs(329) <= not (a and b);
    outputs(330) <= not (a xor b);
    outputs(331) <= a xor b;
    outputs(332) <= not a;
    outputs(333) <= a xor b;
    outputs(334) <= not (a xor b);
    outputs(335) <= a;
    outputs(336) <= not b;
    outputs(337) <= a xor b;
    outputs(338) <= not (a or b);
    outputs(339) <= not b;
    outputs(340) <= a xor b;
    outputs(341) <= a xor b;
    outputs(342) <= a xor b;
    outputs(343) <= a and not b;
    outputs(344) <= not b or a;
    outputs(345) <= not a;
    outputs(346) <= a xor b;
    outputs(347) <= b;
    outputs(348) <= not (a or b);
    outputs(349) <= a and not b;
    outputs(350) <= not b;
    outputs(351) <= not a;
    outputs(352) <= b;
    outputs(353) <= a xor b;
    outputs(354) <= not (a or b);
    outputs(355) <= not b;
    outputs(356) <= not b;
    outputs(357) <= b and not a;
    outputs(358) <= not (a or b);
    outputs(359) <= not b;
    outputs(360) <= a;
    outputs(361) <= a and b;
    outputs(362) <= a and not b;
    outputs(363) <= a and not b;
    outputs(364) <= not b;
    outputs(365) <= not (a and b);
    outputs(366) <= a xor b;
    outputs(367) <= b;
    outputs(368) <= not (a xor b);
    outputs(369) <= not b;
    outputs(370) <= not a or b;
    outputs(371) <= not (a xor b);
    outputs(372) <= a and not b;
    outputs(373) <= b;
    outputs(374) <= not a;
    outputs(375) <= not (a xor b);
    outputs(376) <= b;
    outputs(377) <= not b;
    outputs(378) <= not a;
    outputs(379) <= a xor b;
    outputs(380) <= not (a xor b);
    outputs(381) <= a and not b;
    outputs(382) <= a and not b;
    outputs(383) <= a and b;
    outputs(384) <= not b;
    outputs(385) <= a;
    outputs(386) <= a xor b;
    outputs(387) <= a xor b;
    outputs(388) <= not b;
    outputs(389) <= not (a xor b);
    outputs(390) <= a;
    outputs(391) <= not (a xor b);
    outputs(392) <= a xor b;
    outputs(393) <= b;
    outputs(394) <= a;
    outputs(395) <= a xor b;
    outputs(396) <= not (a xor b);
    outputs(397) <= b;
    outputs(398) <= not b;
    outputs(399) <= b;
    outputs(400) <= not (a xor b);
    outputs(401) <= not (a xor b);
    outputs(402) <= not (a xor b);
    outputs(403) <= not (a or b);
    outputs(404) <= b;
    outputs(405) <= not (a or b);
    outputs(406) <= a and b;
    outputs(407) <= not a or b;
    outputs(408) <= a;
    outputs(409) <= a;
    outputs(410) <= b;
    outputs(411) <= not a or b;
    outputs(412) <= not (a or b);
    outputs(413) <= a;
    outputs(414) <= not a;
    outputs(415) <= a;
    outputs(416) <= not (a xor b);
    outputs(417) <= b;
    outputs(418) <= a xor b;
    outputs(419) <= not b;
    outputs(420) <= not (a xor b);
    outputs(421) <= b and not a;
    outputs(422) <= not a;
    outputs(423) <= a;
    outputs(424) <= not b;
    outputs(425) <= a and b;
    outputs(426) <= a xor b;
    outputs(427) <= not (a xor b);
    outputs(428) <= not b;
    outputs(429) <= a and b;
    outputs(430) <= a xor b;
    outputs(431) <= not (a or b);
    outputs(432) <= a and not b;
    outputs(433) <= not (a xor b);
    outputs(434) <= b;
    outputs(435) <= not a;
    outputs(436) <= not (a or b);
    outputs(437) <= a or b;
    outputs(438) <= b and not a;
    outputs(439) <= not a;
    outputs(440) <= not b;
    outputs(441) <= a;
    outputs(442) <= a;
    outputs(443) <= b and not a;
    outputs(444) <= a xor b;
    outputs(445) <= a xor b;
    outputs(446) <= b and not a;
    outputs(447) <= a and not b;
    outputs(448) <= a xor b;
    outputs(449) <= not (a xor b);
    outputs(450) <= b;
    outputs(451) <= a and b;
    outputs(452) <= a and not b;
    outputs(453) <= not (a or b);
    outputs(454) <= b;
    outputs(455) <= not (a xor b);
    outputs(456) <= a and not b;
    outputs(457) <= not a;
    outputs(458) <= a;
    outputs(459) <= not a;
    outputs(460) <= a and not b;
    outputs(461) <= not b;
    outputs(462) <= not b;
    outputs(463) <= a or b;
    outputs(464) <= b;
    outputs(465) <= not (a xor b);
    outputs(466) <= a and b;
    outputs(467) <= not (a xor b);
    outputs(468) <= b;
    outputs(469) <= not (a xor b);
    outputs(470) <= not b;
    outputs(471) <= not (a xor b);
    outputs(472) <= not (a and b);
    outputs(473) <= a;
    outputs(474) <= a;
    outputs(475) <= a xor b;
    outputs(476) <= a;
    outputs(477) <= a;
    outputs(478) <= not b;
    outputs(479) <= a xor b;
    outputs(480) <= b and not a;
    outputs(481) <= a or b;
    outputs(482) <= not (a xor b);
    outputs(483) <= not a;
    outputs(484) <= a;
    outputs(485) <= a and b;
    outputs(486) <= b;
    outputs(487) <= a or b;
    outputs(488) <= a;
    outputs(489) <= a and not b;
    outputs(490) <= not b;
    outputs(491) <= a or b;
    outputs(492) <= a xor b;
    outputs(493) <= not b or a;
    outputs(494) <= not a;
    outputs(495) <= a and b;
    outputs(496) <= a and not b;
    outputs(497) <= a and b;
    outputs(498) <= not a;
    outputs(499) <= a;
    outputs(500) <= a;
    outputs(501) <= not (a or b);
    outputs(502) <= a xor b;
    outputs(503) <= not a;
    outputs(504) <= not (a or b);
    outputs(505) <= not (a xor b);
    outputs(506) <= b;
    outputs(507) <= a xor b;
    outputs(508) <= a xor b;
    outputs(509) <= not b;
    outputs(510) <= not (a xor b);
    outputs(511) <= a and b;
    outputs(512) <= a and b;
    outputs(513) <= not a;
    outputs(514) <= a xor b;
    outputs(515) <= a;
    outputs(516) <= a xor b;
    outputs(517) <= not b;
    outputs(518) <= a;
    outputs(519) <= not a;
    outputs(520) <= not (a and b);
    outputs(521) <= not a;
    outputs(522) <= not b;
    outputs(523) <= not b;
    outputs(524) <= not (a or b);
    outputs(525) <= not a or b;
    outputs(526) <= not a;
    outputs(527) <= a or b;
    outputs(528) <= not b;
    outputs(529) <= not b;
    outputs(530) <= b;
    outputs(531) <= a and b;
    outputs(532) <= b and not a;
    outputs(533) <= b;
    outputs(534) <= not (a xor b);
    outputs(535) <= a xor b;
    outputs(536) <= a;
    outputs(537) <= a xor b;
    outputs(538) <= a xor b;
    outputs(539) <= not a;
    outputs(540) <= b;
    outputs(541) <= a or b;
    outputs(542) <= not (a xor b);
    outputs(543) <= a and not b;
    outputs(544) <= b;
    outputs(545) <= not b;
    outputs(546) <= not a;
    outputs(547) <= b;
    outputs(548) <= a;
    outputs(549) <= a;
    outputs(550) <= not (a xor b);
    outputs(551) <= not (a xor b);
    outputs(552) <= not a;
    outputs(553) <= not (a xor b);
    outputs(554) <= a;
    outputs(555) <= not b;
    outputs(556) <= not a;
    outputs(557) <= not a or b;
    outputs(558) <= not (a and b);
    outputs(559) <= not (a xor b);
    outputs(560) <= not a;
    outputs(561) <= not (a or b);
    outputs(562) <= b;
    outputs(563) <= b and not a;
    outputs(564) <= not (a xor b);
    outputs(565) <= not (a xor b);
    outputs(566) <= not a or b;
    outputs(567) <= a;
    outputs(568) <= not (a xor b);
    outputs(569) <= not (a xor b);
    outputs(570) <= not a;
    outputs(571) <= not (a xor b);
    outputs(572) <= not a;
    outputs(573) <= a;
    outputs(574) <= not a;
    outputs(575) <= a;
    outputs(576) <= not a;
    outputs(577) <= a;
    outputs(578) <= not (a xor b);
    outputs(579) <= not (a xor b);
    outputs(580) <= b and not a;
    outputs(581) <= not b;
    outputs(582) <= not b;
    outputs(583) <= a and b;
    outputs(584) <= a and b;
    outputs(585) <= not (a xor b);
    outputs(586) <= a and b;
    outputs(587) <= not b;
    outputs(588) <= not b;
    outputs(589) <= a or b;
    outputs(590) <= not a;
    outputs(591) <= not b;
    outputs(592) <= a xor b;
    outputs(593) <= not (a xor b);
    outputs(594) <= not a;
    outputs(595) <= a xor b;
    outputs(596) <= a xor b;
    outputs(597) <= not b;
    outputs(598) <= b;
    outputs(599) <= a and not b;
    outputs(600) <= not a;
    outputs(601) <= not b or a;
    outputs(602) <= not b or a;
    outputs(603) <= not b;
    outputs(604) <= b and not a;
    outputs(605) <= not (a xor b);
    outputs(606) <= not (a or b);
    outputs(607) <= a;
    outputs(608) <= b;
    outputs(609) <= a;
    outputs(610) <= b;
    outputs(611) <= not a;
    outputs(612) <= a;
    outputs(613) <= b;
    outputs(614) <= not a;
    outputs(615) <= a and not b;
    outputs(616) <= a xor b;
    outputs(617) <= not a;
    outputs(618) <= not (a xor b);
    outputs(619) <= not a;
    outputs(620) <= b;
    outputs(621) <= not b;
    outputs(622) <= b;
    outputs(623) <= b and not a;
    outputs(624) <= not b;
    outputs(625) <= not a;
    outputs(626) <= a xor b;
    outputs(627) <= a or b;
    outputs(628) <= b;
    outputs(629) <= not b;
    outputs(630) <= a;
    outputs(631) <= a;
    outputs(632) <= not a;
    outputs(633) <= a xor b;
    outputs(634) <= not (a xor b);
    outputs(635) <= a and b;
    outputs(636) <= not (a xor b);
    outputs(637) <= a and b;
    outputs(638) <= a;
    outputs(639) <= not a;
    outputs(640) <= a and not b;
    outputs(641) <= not (a xor b);
    outputs(642) <= not b;
    outputs(643) <= not a or b;
    outputs(644) <= a;
    outputs(645) <= a and b;
    outputs(646) <= a xor b;
    outputs(647) <= not a or b;
    outputs(648) <= b;
    outputs(649) <= a and not b;
    outputs(650) <= a and not b;
    outputs(651) <= not b;
    outputs(652) <= not b;
    outputs(653) <= a xor b;
    outputs(654) <= a;
    outputs(655) <= not (a xor b);
    outputs(656) <= a and not b;
    outputs(657) <= b and not a;
    outputs(658) <= not (a and b);
    outputs(659) <= b;
    outputs(660) <= b and not a;
    outputs(661) <= not a or b;
    outputs(662) <= a and b;
    outputs(663) <= not a;
    outputs(664) <= not b;
    outputs(665) <= a;
    outputs(666) <= a and b;
    outputs(667) <= not (a xor b);
    outputs(668) <= not (a or b);
    outputs(669) <= a;
    outputs(670) <= not (a xor b);
    outputs(671) <= not b;
    outputs(672) <= not b;
    outputs(673) <= a xor b;
    outputs(674) <= a and b;
    outputs(675) <= not a;
    outputs(676) <= a;
    outputs(677) <= b;
    outputs(678) <= b;
    outputs(679) <= not a;
    outputs(680) <= not (a or b);
    outputs(681) <= b;
    outputs(682) <= a;
    outputs(683) <= not a;
    outputs(684) <= a;
    outputs(685) <= not (a xor b);
    outputs(686) <= a xor b;
    outputs(687) <= a or b;
    outputs(688) <= a xor b;
    outputs(689) <= b and not a;
    outputs(690) <= a xor b;
    outputs(691) <= not (a and b);
    outputs(692) <= a xor b;
    outputs(693) <= not a;
    outputs(694) <= not b or a;
    outputs(695) <= not (a or b);
    outputs(696) <= not (a xor b);
    outputs(697) <= a;
    outputs(698) <= b;
    outputs(699) <= a;
    outputs(700) <= not b;
    outputs(701) <= b and not a;
    outputs(702) <= not b;
    outputs(703) <= a or b;
    outputs(704) <= b and not a;
    outputs(705) <= a or b;
    outputs(706) <= not a;
    outputs(707) <= not (a or b);
    outputs(708) <= not (a xor b);
    outputs(709) <= a;
    outputs(710) <= b;
    outputs(711) <= not b or a;
    outputs(712) <= b;
    outputs(713) <= not (a or b);
    outputs(714) <= a and not b;
    outputs(715) <= not (a xor b);
    outputs(716) <= a xor b;
    outputs(717) <= b;
    outputs(718) <= not (a xor b);
    outputs(719) <= not a or b;
    outputs(720) <= a xor b;
    outputs(721) <= a or b;
    outputs(722) <= not b;
    outputs(723) <= not a;
    outputs(724) <= b and not a;
    outputs(725) <= a;
    outputs(726) <= b;
    outputs(727) <= a and b;
    outputs(728) <= a xor b;
    outputs(729) <= not a;
    outputs(730) <= not (a xor b);
    outputs(731) <= not a;
    outputs(732) <= a xor b;
    outputs(733) <= not b;
    outputs(734) <= not (a xor b);
    outputs(735) <= b;
    outputs(736) <= not (a xor b);
    outputs(737) <= a xor b;
    outputs(738) <= a and b;
    outputs(739) <= not (a xor b);
    outputs(740) <= a and not b;
    outputs(741) <= not (a xor b);
    outputs(742) <= not (a xor b);
    outputs(743) <= not (a or b);
    outputs(744) <= not (a xor b);
    outputs(745) <= not (a xor b);
    outputs(746) <= b;
    outputs(747) <= not (a xor b);
    outputs(748) <= not (a or b);
    outputs(749) <= b and not a;
    outputs(750) <= a xor b;
    outputs(751) <= a;
    outputs(752) <= not b;
    outputs(753) <= not a;
    outputs(754) <= not b;
    outputs(755) <= not b or a;
    outputs(756) <= not a;
    outputs(757) <= not (a and b);
    outputs(758) <= not (a xor b);
    outputs(759) <= a and not b;
    outputs(760) <= a xor b;
    outputs(761) <= not (a and b);
    outputs(762) <= not (a and b);
    outputs(763) <= a and b;
    outputs(764) <= not b;
    outputs(765) <= not b;
    outputs(766) <= a and not b;
    outputs(767) <= a;
    outputs(768) <= not (a or b);
    outputs(769) <= a and not b;
    outputs(770) <= a;
    outputs(771) <= a;
    outputs(772) <= a or b;
    outputs(773) <= not (a xor b);
    outputs(774) <= not a or b;
    outputs(775) <= b;
    outputs(776) <= a xor b;
    outputs(777) <= not a or b;
    outputs(778) <= a or b;
    outputs(779) <= a;
    outputs(780) <= a or b;
    outputs(781) <= not b;
    outputs(782) <= a xor b;
    outputs(783) <= a;
    outputs(784) <= a xor b;
    outputs(785) <= a xor b;
    outputs(786) <= a and not b;
    outputs(787) <= a;
    outputs(788) <= not b;
    outputs(789) <= not (a xor b);
    outputs(790) <= a xor b;
    outputs(791) <= not (a xor b);
    outputs(792) <= not b;
    outputs(793) <= a xor b;
    outputs(794) <= not b;
    outputs(795) <= not b;
    outputs(796) <= a and b;
    outputs(797) <= not b;
    outputs(798) <= a and not b;
    outputs(799) <= b and not a;
    outputs(800) <= not a;
    outputs(801) <= a and not b;
    outputs(802) <= not a;
    outputs(803) <= not a;
    outputs(804) <= a xor b;
    outputs(805) <= not b;
    outputs(806) <= not (a and b);
    outputs(807) <= not (a xor b);
    outputs(808) <= b;
    outputs(809) <= a and b;
    outputs(810) <= a;
    outputs(811) <= not (a xor b);
    outputs(812) <= a;
    outputs(813) <= not a;
    outputs(814) <= not (a xor b);
    outputs(815) <= not (a and b);
    outputs(816) <= not b;
    outputs(817) <= not (a xor b);
    outputs(818) <= a xor b;
    outputs(819) <= not b;
    outputs(820) <= not (a xor b);
    outputs(821) <= a and not b;
    outputs(822) <= a;
    outputs(823) <= not b;
    outputs(824) <= not (a xor b);
    outputs(825) <= not (a xor b);
    outputs(826) <= a or b;
    outputs(827) <= a;
    outputs(828) <= a and b;
    outputs(829) <= a and not b;
    outputs(830) <= not (a xor b);
    outputs(831) <= not a;
    outputs(832) <= b and not a;
    outputs(833) <= not (a xor b);
    outputs(834) <= a and not b;
    outputs(835) <= a and b;
    outputs(836) <= a and not b;
    outputs(837) <= a;
    outputs(838) <= a and b;
    outputs(839) <= a;
    outputs(840) <= a xor b;
    outputs(841) <= not b;
    outputs(842) <= a and not b;
    outputs(843) <= not b;
    outputs(844) <= a xor b;
    outputs(845) <= a;
    outputs(846) <= not (a xor b);
    outputs(847) <= a xor b;
    outputs(848) <= not (a or b);
    outputs(849) <= a and not b;
    outputs(850) <= a;
    outputs(851) <= a;
    outputs(852) <= not (a or b);
    outputs(853) <= not b;
    outputs(854) <= b;
    outputs(855) <= b and not a;
    outputs(856) <= b;
    outputs(857) <= a;
    outputs(858) <= a;
    outputs(859) <= a and not b;
    outputs(860) <= b;
    outputs(861) <= not b or a;
    outputs(862) <= a and b;
    outputs(863) <= not b or a;
    outputs(864) <= not (a xor b);
    outputs(865) <= not (a xor b);
    outputs(866) <= a and not b;
    outputs(867) <= a;
    outputs(868) <= a xor b;
    outputs(869) <= a and not b;
    outputs(870) <= not (a xor b);
    outputs(871) <= a;
    outputs(872) <= a xor b;
    outputs(873) <= a xor b;
    outputs(874) <= a;
    outputs(875) <= not a or b;
    outputs(876) <= not b;
    outputs(877) <= b and not a;
    outputs(878) <= not b;
    outputs(879) <= b;
    outputs(880) <= not b;
    outputs(881) <= not (a xor b);
    outputs(882) <= not (a or b);
    outputs(883) <= not (a xor b);
    outputs(884) <= a xor b;
    outputs(885) <= a and b;
    outputs(886) <= not (a xor b);
    outputs(887) <= b;
    outputs(888) <= b;
    outputs(889) <= a xor b;
    outputs(890) <= a;
    outputs(891) <= a or b;
    outputs(892) <= not (a xor b);
    outputs(893) <= not (a xor b);
    outputs(894) <= not (a xor b);
    outputs(895) <= not a;
    outputs(896) <= not a or b;
    outputs(897) <= a and b;
    outputs(898) <= not a;
    outputs(899) <= not (a xor b);
    outputs(900) <= not b;
    outputs(901) <= not (a or b);
    outputs(902) <= a;
    outputs(903) <= not (a or b);
    outputs(904) <= not (a xor b);
    outputs(905) <= a xor b;
    outputs(906) <= not (a xor b);
    outputs(907) <= not (a or b);
    outputs(908) <= not b;
    outputs(909) <= not (a and b);
    outputs(910) <= not (a xor b);
    outputs(911) <= b;
    outputs(912) <= a xor b;
    outputs(913) <= not a or b;
    outputs(914) <= b;
    outputs(915) <= a;
    outputs(916) <= not b;
    outputs(917) <= a;
    outputs(918) <= not a;
    outputs(919) <= a xor b;
    outputs(920) <= not (a xor b);
    outputs(921) <= a and not b;
    outputs(922) <= not (a xor b);
    outputs(923) <= b;
    outputs(924) <= a xor b;
    outputs(925) <= a xor b;
    outputs(926) <= not b;
    outputs(927) <= a xor b;
    outputs(928) <= b;
    outputs(929) <= a xor b;
    outputs(930) <= not b;
    outputs(931) <= not (a xor b);
    outputs(932) <= not b;
    outputs(933) <= b;
    outputs(934) <= not (a and b);
    outputs(935) <= not b;
    outputs(936) <= a xor b;
    outputs(937) <= b and not a;
    outputs(938) <= b;
    outputs(939) <= not b;
    outputs(940) <= a xor b;
    outputs(941) <= a and not b;
    outputs(942) <= not a or b;
    outputs(943) <= a;
    outputs(944) <= not b or a;
    outputs(945) <= not (a or b);
    outputs(946) <= b and not a;
    outputs(947) <= b;
    outputs(948) <= a and b;
    outputs(949) <= a;
    outputs(950) <= not b or a;
    outputs(951) <= not a;
    outputs(952) <= not (a xor b);
    outputs(953) <= a;
    outputs(954) <= a and b;
    outputs(955) <= not (a and b);
    outputs(956) <= not (a xor b);
    outputs(957) <= b;
    outputs(958) <= a;
    outputs(959) <= a xor b;
    outputs(960) <= not a or b;
    outputs(961) <= a;
    outputs(962) <= not (a xor b);
    outputs(963) <= not b;
    outputs(964) <= b;
    outputs(965) <= a;
    outputs(966) <= a and not b;
    outputs(967) <= not (a and b);
    outputs(968) <= a and b;
    outputs(969) <= a xor b;
    outputs(970) <= a xor b;
    outputs(971) <= not a;
    outputs(972) <= not (a xor b);
    outputs(973) <= a and not b;
    outputs(974) <= a xor b;
    outputs(975) <= not (a and b);
    outputs(976) <= not a;
    outputs(977) <= not (a xor b);
    outputs(978) <= a;
    outputs(979) <= a;
    outputs(980) <= a and not b;
    outputs(981) <= not (a xor b);
    outputs(982) <= not (a or b);
    outputs(983) <= a and not b;
    outputs(984) <= not (a xor b);
    outputs(985) <= b;
    outputs(986) <= b;
    outputs(987) <= not a;
    outputs(988) <= a;
    outputs(989) <= not (a xor b);
    outputs(990) <= not a;
    outputs(991) <= not (a xor b);
    outputs(992) <= not (a and b);
    outputs(993) <= a;
    outputs(994) <= a xor b;
    outputs(995) <= not a;
    outputs(996) <= a;
    outputs(997) <= not (a or b);
    outputs(998) <= not b;
    outputs(999) <= a;
    outputs(1000) <= not b;
    outputs(1001) <= b;
    outputs(1002) <= b;
    outputs(1003) <= not a;
    outputs(1004) <= a and b;
    outputs(1005) <= a;
    outputs(1006) <= not b;
    outputs(1007) <= not (a and b);
    outputs(1008) <= a xor b;
    outputs(1009) <= not b or a;
    outputs(1010) <= a and not b;
    outputs(1011) <= a xor b;
    outputs(1012) <= not (a xor b);
    outputs(1013) <= b;
    outputs(1014) <= a;
    outputs(1015) <= a;
    outputs(1016) <= a and not b;
    outputs(1017) <= a xor b;
    outputs(1018) <= not (a or b);
    outputs(1019) <= not (a xor b);
    outputs(1020) <= b;
    outputs(1021) <= not (a or b);
    outputs(1022) <= a xor b;
    outputs(1023) <= a xor b;
    outputs(1024) <= a and b;
    outputs(1025) <= a xor b;
    outputs(1026) <= b and not a;
    outputs(1027) <= b and not a;
    outputs(1028) <= not (a xor b);
    outputs(1029) <= not (a xor b);
    outputs(1030) <= b and not a;
    outputs(1031) <= b and not a;
    outputs(1032) <= b and not a;
    outputs(1033) <= a and b;
    outputs(1034) <= not b or a;
    outputs(1035) <= a;
    outputs(1036) <= b;
    outputs(1037) <= not (a xor b);
    outputs(1038) <= a and b;
    outputs(1039) <= not a;
    outputs(1040) <= not (a or b);
    outputs(1041) <= a and not b;
    outputs(1042) <= not (a or b);
    outputs(1043) <= a;
    outputs(1044) <= not (a xor b);
    outputs(1045) <= not b;
    outputs(1046) <= a xor b;
    outputs(1047) <= not (a or b);
    outputs(1048) <= a and not b;
    outputs(1049) <= b;
    outputs(1050) <= a and not b;
    outputs(1051) <= a and not b;
    outputs(1052) <= a;
    outputs(1053) <= not (a xor b);
    outputs(1054) <= a;
    outputs(1055) <= b and not a;
    outputs(1056) <= a and b;
    outputs(1057) <= a;
    outputs(1058) <= not (a or b);
    outputs(1059) <= a;
    outputs(1060) <= a and not b;
    outputs(1061) <= a and not b;
    outputs(1062) <= a xor b;
    outputs(1063) <= a and not b;
    outputs(1064) <= not b;
    outputs(1065) <= not a or b;
    outputs(1066) <= a xor b;
    outputs(1067) <= not a;
    outputs(1068) <= b and not a;
    outputs(1069) <= b;
    outputs(1070) <= a and not b;
    outputs(1071) <= b and not a;
    outputs(1072) <= a xor b;
    outputs(1073) <= b;
    outputs(1074) <= a and b;
    outputs(1075) <= a;
    outputs(1076) <= a and b;
    outputs(1077) <= not (a or b);
    outputs(1078) <= not (a xor b);
    outputs(1079) <= b and not a;
    outputs(1080) <= a and not b;
    outputs(1081) <= not (a or b);
    outputs(1082) <= b and not a;
    outputs(1083) <= not a;
    outputs(1084) <= a and b;
    outputs(1085) <= not a;
    outputs(1086) <= b and not a;
    outputs(1087) <= b and not a;
    outputs(1088) <= not (a or b);
    outputs(1089) <= b and not a;
    outputs(1090) <= b and not a;
    outputs(1091) <= a xor b;
    outputs(1092) <= not a;
    outputs(1093) <= b and not a;
    outputs(1094) <= not b;
    outputs(1095) <= b and not a;
    outputs(1096) <= not (a or b);
    outputs(1097) <= '0';
    outputs(1098) <= a and b;
    outputs(1099) <= b and not a;
    outputs(1100) <= a and b;
    outputs(1101) <= a and not b;
    outputs(1102) <= b and not a;
    outputs(1103) <= not a;
    outputs(1104) <= a and not b;
    outputs(1105) <= a xor b;
    outputs(1106) <= b and not a;
    outputs(1107) <= a and not b;
    outputs(1108) <= not a;
    outputs(1109) <= b and not a;
    outputs(1110) <= b and not a;
    outputs(1111) <= a and not b;
    outputs(1112) <= not (a or b);
    outputs(1113) <= b and not a;
    outputs(1114) <= b and not a;
    outputs(1115) <= a;
    outputs(1116) <= a and b;
    outputs(1117) <= b and not a;
    outputs(1118) <= not a;
    outputs(1119) <= a xor b;
    outputs(1120) <= b and not a;
    outputs(1121) <= a and not b;
    outputs(1122) <= b and not a;
    outputs(1123) <= b and not a;
    outputs(1124) <= a and not b;
    outputs(1125) <= a and not b;
    outputs(1126) <= b and not a;
    outputs(1127) <= b and not a;
    outputs(1128) <= a and not b;
    outputs(1129) <= a xor b;
    outputs(1130) <= not b;
    outputs(1131) <= not a;
    outputs(1132) <= a and b;
    outputs(1133) <= a xor b;
    outputs(1134) <= a and not b;
    outputs(1135) <= a xor b;
    outputs(1136) <= not b;
    outputs(1137) <= '0';
    outputs(1138) <= not (a xor b);
    outputs(1139) <= b and not a;
    outputs(1140) <= b and not a;
    outputs(1141) <= '0';
    outputs(1142) <= not a;
    outputs(1143) <= a and not b;
    outputs(1144) <= b;
    outputs(1145) <= not a;
    outputs(1146) <= a xor b;
    outputs(1147) <= not (a or b);
    outputs(1148) <= a and not b;
    outputs(1149) <= not (a or b);
    outputs(1150) <= not (a xor b);
    outputs(1151) <= a xor b;
    outputs(1152) <= a and not b;
    outputs(1153) <= a and not b;
    outputs(1154) <= a xor b;
    outputs(1155) <= b;
    outputs(1156) <= b;
    outputs(1157) <= not (a xor b);
    outputs(1158) <= a and not b;
    outputs(1159) <= a and not b;
    outputs(1160) <= b;
    outputs(1161) <= b and not a;
    outputs(1162) <= b;
    outputs(1163) <= a and not b;
    outputs(1164) <= b and not a;
    outputs(1165) <= a xor b;
    outputs(1166) <= a xor b;
    outputs(1167) <= a and not b;
    outputs(1168) <= not (a or b);
    outputs(1169) <= a and not b;
    outputs(1170) <= b;
    outputs(1171) <= not (a xor b);
    outputs(1172) <= not (a or b);
    outputs(1173) <= '0';
    outputs(1174) <= a and b;
    outputs(1175) <= a xor b;
    outputs(1176) <= not a or b;
    outputs(1177) <= b and not a;
    outputs(1178) <= not (a or b);
    outputs(1179) <= a and not b;
    outputs(1180) <= a and b;
    outputs(1181) <= a and b;
    outputs(1182) <= b and not a;
    outputs(1183) <= a and b;
    outputs(1184) <= a xor b;
    outputs(1185) <= not (a or b);
    outputs(1186) <= not (a xor b);
    outputs(1187) <= '0';
    outputs(1188) <= not (a xor b);
    outputs(1189) <= a and b;
    outputs(1190) <= not (a or b);
    outputs(1191) <= not a or b;
    outputs(1192) <= not b;
    outputs(1193) <= not (a xor b);
    outputs(1194) <= not (a or b);
    outputs(1195) <= a and b;
    outputs(1196) <= not b;
    outputs(1197) <= a;
    outputs(1198) <= not b;
    outputs(1199) <= '0';
    outputs(1200) <= b;
    outputs(1201) <= a xor b;
    outputs(1202) <= not b;
    outputs(1203) <= not (a xor b);
    outputs(1204) <= b;
    outputs(1205) <= a and b;
    outputs(1206) <= not (a and b);
    outputs(1207) <= a and not b;
    outputs(1208) <= a xor b;
    outputs(1209) <= b;
    outputs(1210) <= a and not b;
    outputs(1211) <= a xor b;
    outputs(1212) <= '0';
    outputs(1213) <= not (a or b);
    outputs(1214) <= a and not b;
    outputs(1215) <= a and b;
    outputs(1216) <= not (a xor b);
    outputs(1217) <= a and not b;
    outputs(1218) <= a and b;
    outputs(1219) <= b;
    outputs(1220) <= b and not a;
    outputs(1221) <= not a;
    outputs(1222) <= not b;
    outputs(1223) <= not (a or b);
    outputs(1224) <= a xor b;
    outputs(1225) <= a and b;
    outputs(1226) <= not (a or b);
    outputs(1227) <= b;
    outputs(1228) <= a;
    outputs(1229) <= not (a or b);
    outputs(1230) <= not (a or b);
    outputs(1231) <= a xor b;
    outputs(1232) <= a and not b;
    outputs(1233) <= a and b;
    outputs(1234) <= a and not b;
    outputs(1235) <= a and b;
    outputs(1236) <= not a;
    outputs(1237) <= a and b;
    outputs(1238) <= b and not a;
    outputs(1239) <= not (a xor b);
    outputs(1240) <= not a;
    outputs(1241) <= not (a or b);
    outputs(1242) <= a and b;
    outputs(1243) <= not b;
    outputs(1244) <= not a;
    outputs(1245) <= a;
    outputs(1246) <= '0';
    outputs(1247) <= a;
    outputs(1248) <= a;
    outputs(1249) <= a and b;
    outputs(1250) <= a;
    outputs(1251) <= b and not a;
    outputs(1252) <= a xor b;
    outputs(1253) <= a and not b;
    outputs(1254) <= b and not a;
    outputs(1255) <= a and b;
    outputs(1256) <= not b;
    outputs(1257) <= b;
    outputs(1258) <= not (a and b);
    outputs(1259) <= not a;
    outputs(1260) <= a xor b;
    outputs(1261) <= not (a or b);
    outputs(1262) <= b and not a;
    outputs(1263) <= not (a or b);
    outputs(1264) <= not b;
    outputs(1265) <= a and not b;
    outputs(1266) <= not b;
    outputs(1267) <= a;
    outputs(1268) <= not b;
    outputs(1269) <= b;
    outputs(1270) <= not (a or b);
    outputs(1271) <= b and not a;
    outputs(1272) <= b and not a;
    outputs(1273) <= a and not b;
    outputs(1274) <= a and b;
    outputs(1275) <= not b;
    outputs(1276) <= b;
    outputs(1277) <= not a;
    outputs(1278) <= a and not b;
    outputs(1279) <= not b;
    outputs(1280) <= b and not a;
    outputs(1281) <= not (a xor b);
    outputs(1282) <= '0';
    outputs(1283) <= a and b;
    outputs(1284) <= a and b;
    outputs(1285) <= a and not b;
    outputs(1286) <= not a;
    outputs(1287) <= a and b;
    outputs(1288) <= a;
    outputs(1289) <= a and not b;
    outputs(1290) <= a and b;
    outputs(1291) <= not (a or b);
    outputs(1292) <= not (a xor b);
    outputs(1293) <= a and b;
    outputs(1294) <= not (a or b);
    outputs(1295) <= a;
    outputs(1296) <= not (a xor b);
    outputs(1297) <= not (a xor b);
    outputs(1298) <= a;
    outputs(1299) <= a and not b;
    outputs(1300) <= not a;
    outputs(1301) <= not b;
    outputs(1302) <= a and b;
    outputs(1303) <= a and not b;
    outputs(1304) <= not (a or b);
    outputs(1305) <= b and not a;
    outputs(1306) <= not b;
    outputs(1307) <= not b;
    outputs(1308) <= not a;
    outputs(1309) <= b and not a;
    outputs(1310) <= '0';
    outputs(1311) <= a and not b;
    outputs(1312) <= not (a or b);
    outputs(1313) <= a xor b;
    outputs(1314) <= not a;
    outputs(1315) <= a and not b;
    outputs(1316) <= b;
    outputs(1317) <= b and not a;
    outputs(1318) <= a and b;
    outputs(1319) <= not a;
    outputs(1320) <= b and not a;
    outputs(1321) <= not a;
    outputs(1322) <= not b;
    outputs(1323) <= not b;
    outputs(1324) <= b;
    outputs(1325) <= a and not b;
    outputs(1326) <= not (a or b);
    outputs(1327) <= b;
    outputs(1328) <= not (a or b);
    outputs(1329) <= b and not a;
    outputs(1330) <= a or b;
    outputs(1331) <= not a;
    outputs(1332) <= a and b;
    outputs(1333) <= a;
    outputs(1334) <= not a;
    outputs(1335) <= b and not a;
    outputs(1336) <= '0';
    outputs(1337) <= a;
    outputs(1338) <= a and b;
    outputs(1339) <= not a;
    outputs(1340) <= not b;
    outputs(1341) <= a and b;
    outputs(1342) <= a and not b;
    outputs(1343) <= a and not b;
    outputs(1344) <= a;
    outputs(1345) <= b and not a;
    outputs(1346) <= b;
    outputs(1347) <= not (a or b);
    outputs(1348) <= a and not b;
    outputs(1349) <= a and b;
    outputs(1350) <= b;
    outputs(1351) <= not (a or b);
    outputs(1352) <= not (a or b);
    outputs(1353) <= not (a or b);
    outputs(1354) <= a and not b;
    outputs(1355) <= a and b;
    outputs(1356) <= not a;
    outputs(1357) <= a and b;
    outputs(1358) <= b;
    outputs(1359) <= b;
    outputs(1360) <= not b;
    outputs(1361) <= a;
    outputs(1362) <= b and not a;
    outputs(1363) <= a xor b;
    outputs(1364) <= not (a or b);
    outputs(1365) <= a xor b;
    outputs(1366) <= a and not b;
    outputs(1367) <= b and not a;
    outputs(1368) <= not a;
    outputs(1369) <= a;
    outputs(1370) <= b and not a;
    outputs(1371) <= a xor b;
    outputs(1372) <= not (a xor b);
    outputs(1373) <= b and not a;
    outputs(1374) <= a;
    outputs(1375) <= b;
    outputs(1376) <= b and not a;
    outputs(1377) <= b and not a;
    outputs(1378) <= b and not a;
    outputs(1379) <= b and not a;
    outputs(1380) <= a xor b;
    outputs(1381) <= b and not a;
    outputs(1382) <= not (a or b);
    outputs(1383) <= not (a and b);
    outputs(1384) <= a xor b;
    outputs(1385) <= a and not b;
    outputs(1386) <= a and b;
    outputs(1387) <= a and b;
    outputs(1388) <= b and not a;
    outputs(1389) <= '0';
    outputs(1390) <= b;
    outputs(1391) <= a xor b;
    outputs(1392) <= a and b;
    outputs(1393) <= a and not b;
    outputs(1394) <= a and b;
    outputs(1395) <= not (a or b);
    outputs(1396) <= a and b;
    outputs(1397) <= b and not a;
    outputs(1398) <= a xor b;
    outputs(1399) <= a and not b;
    outputs(1400) <= not (a xor b);
    outputs(1401) <= not (a or b);
    outputs(1402) <= a xor b;
    outputs(1403) <= a and b;
    outputs(1404) <= a and b;
    outputs(1405) <= '0';
    outputs(1406) <= a and b;
    outputs(1407) <= a and not b;
    outputs(1408) <= not (a xor b);
    outputs(1409) <= a;
    outputs(1410) <= not a;
    outputs(1411) <= b;
    outputs(1412) <= a and not b;
    outputs(1413) <= not (a xor b);
    outputs(1414) <= not (a or b);
    outputs(1415) <= b;
    outputs(1416) <= not a;
    outputs(1417) <= a and not b;
    outputs(1418) <= not (a or b);
    outputs(1419) <= a and not b;
    outputs(1420) <= a and b;
    outputs(1421) <= a and not b;
    outputs(1422) <= b;
    outputs(1423) <= b and not a;
    outputs(1424) <= a xor b;
    outputs(1425) <= b;
    outputs(1426) <= b and not a;
    outputs(1427) <= b and not a;
    outputs(1428) <= a and b;
    outputs(1429) <= b and not a;
    outputs(1430) <= a and b;
    outputs(1431) <= not (a or b);
    outputs(1432) <= not b;
    outputs(1433) <= a xor b;
    outputs(1434) <= b and not a;
    outputs(1435) <= a and b;
    outputs(1436) <= not (a or b);
    outputs(1437) <= a xor b;
    outputs(1438) <= not a;
    outputs(1439) <= a xor b;
    outputs(1440) <= '0';
    outputs(1441) <= not a;
    outputs(1442) <= a;
    outputs(1443) <= not (a or b);
    outputs(1444) <= a;
    outputs(1445) <= a and not b;
    outputs(1446) <= not (a xor b);
    outputs(1447) <= a or b;
    outputs(1448) <= b and not a;
    outputs(1449) <= a and b;
    outputs(1450) <= not a;
    outputs(1451) <= not (a xor b);
    outputs(1452) <= a xor b;
    outputs(1453) <= not (a or b);
    outputs(1454) <= b;
    outputs(1455) <= a;
    outputs(1456) <= not (a or b);
    outputs(1457) <= b and not a;
    outputs(1458) <= b and not a;
    outputs(1459) <= b and not a;
    outputs(1460) <= not b;
    outputs(1461) <= b;
    outputs(1462) <= not (a or b);
    outputs(1463) <= not (a or b);
    outputs(1464) <= b and not a;
    outputs(1465) <= a;
    outputs(1466) <= a and b;
    outputs(1467) <= a and not b;
    outputs(1468) <= not (a xor b);
    outputs(1469) <= a and b;
    outputs(1470) <= a xor b;
    outputs(1471) <= not a;
    outputs(1472) <= a and not b;
    outputs(1473) <= a and not b;
    outputs(1474) <= b;
    outputs(1475) <= not a;
    outputs(1476) <= not b;
    outputs(1477) <= not (a xor b);
    outputs(1478) <= not a;
    outputs(1479) <= a and b;
    outputs(1480) <= not b;
    outputs(1481) <= a and not b;
    outputs(1482) <= not (a xor b);
    outputs(1483) <= b;
    outputs(1484) <= not (a or b);
    outputs(1485) <= a;
    outputs(1486) <= a and b;
    outputs(1487) <= '0';
    outputs(1488) <= a and not b;
    outputs(1489) <= not a;
    outputs(1490) <= not a;
    outputs(1491) <= a xor b;
    outputs(1492) <= not (a or b);
    outputs(1493) <= not (a xor b);
    outputs(1494) <= a and b;
    outputs(1495) <= not b;
    outputs(1496) <= a and not b;
    outputs(1497) <= a and not b;
    outputs(1498) <= '0';
    outputs(1499) <= a;
    outputs(1500) <= b and not a;
    outputs(1501) <= b and not a;
    outputs(1502) <= a and not b;
    outputs(1503) <= a and b;
    outputs(1504) <= b and not a;
    outputs(1505) <= a xor b;
    outputs(1506) <= a and not b;
    outputs(1507) <= not b;
    outputs(1508) <= a xor b;
    outputs(1509) <= b and not a;
    outputs(1510) <= a;
    outputs(1511) <= a and b;
    outputs(1512) <= not (a xor b);
    outputs(1513) <= a and b;
    outputs(1514) <= b and not a;
    outputs(1515) <= b and not a;
    outputs(1516) <= b;
    outputs(1517) <= b and not a;
    outputs(1518) <= a xor b;
    outputs(1519) <= not a or b;
    outputs(1520) <= not (a or b);
    outputs(1521) <= a;
    outputs(1522) <= a and not b;
    outputs(1523) <= '0';
    outputs(1524) <= a xor b;
    outputs(1525) <= not a or b;
    outputs(1526) <= b and not a;
    outputs(1527) <= '0';
    outputs(1528) <= not (a or b);
    outputs(1529) <= not (a xor b);
    outputs(1530) <= not (a xor b);
    outputs(1531) <= not (a xor b);
    outputs(1532) <= not (a xor b);
    outputs(1533) <= not b;
    outputs(1534) <= b and not a;
    outputs(1535) <= b and not a;
    outputs(1536) <= a;
    outputs(1537) <= a and b;
    outputs(1538) <= a and b;
    outputs(1539) <= a;
    outputs(1540) <= not (a xor b);
    outputs(1541) <= not (a or b);
    outputs(1542) <= not a;
    outputs(1543) <= '0';
    outputs(1544) <= a xor b;
    outputs(1545) <= not (a xor b);
    outputs(1546) <= not b;
    outputs(1547) <= a;
    outputs(1548) <= a and not b;
    outputs(1549) <= a and b;
    outputs(1550) <= not (a or b);
    outputs(1551) <= a and not b;
    outputs(1552) <= not (a xor b);
    outputs(1553) <= a;
    outputs(1554) <= b and not a;
    outputs(1555) <= a and not b;
    outputs(1556) <= not a;
    outputs(1557) <= b and not a;
    outputs(1558) <= a and b;
    outputs(1559) <= not (a or b);
    outputs(1560) <= a and not b;
    outputs(1561) <= b and not a;
    outputs(1562) <= a xor b;
    outputs(1563) <= b and not a;
    outputs(1564) <= not a;
    outputs(1565) <= not (a or b);
    outputs(1566) <= b and not a;
    outputs(1567) <= not (a or b);
    outputs(1568) <= not a;
    outputs(1569) <= a and not b;
    outputs(1570) <= a and not b;
    outputs(1571) <= not (a xor b);
    outputs(1572) <= a xor b;
    outputs(1573) <= not b;
    outputs(1574) <= not a;
    outputs(1575) <= a and b;
    outputs(1576) <= a and not b;
    outputs(1577) <= a xor b;
    outputs(1578) <= not a;
    outputs(1579) <= not (a xor b);
    outputs(1580) <= not (a xor b);
    outputs(1581) <= b;
    outputs(1582) <= a and b;
    outputs(1583) <= b and not a;
    outputs(1584) <= b and not a;
    outputs(1585) <= a xor b;
    outputs(1586) <= a and not b;
    outputs(1587) <= a and not b;
    outputs(1588) <= b;
    outputs(1589) <= a and b;
    outputs(1590) <= not (a or b);
    outputs(1591) <= not (a or b);
    outputs(1592) <= a xor b;
    outputs(1593) <= b and not a;
    outputs(1594) <= not b;
    outputs(1595) <= not a;
    outputs(1596) <= not b;
    outputs(1597) <= a and not b;
    outputs(1598) <= '0';
    outputs(1599) <= b;
    outputs(1600) <= a and not b;
    outputs(1601) <= not (a or b);
    outputs(1602) <= a and not b;
    outputs(1603) <= not a;
    outputs(1604) <= a and b;
    outputs(1605) <= '0';
    outputs(1606) <= a xor b;
    outputs(1607) <= not a;
    outputs(1608) <= a xor b;
    outputs(1609) <= not (a xor b);
    outputs(1610) <= not a;
    outputs(1611) <= not (a or b);
    outputs(1612) <= b;
    outputs(1613) <= a and not b;
    outputs(1614) <= b and not a;
    outputs(1615) <= a and b;
    outputs(1616) <= a;
    outputs(1617) <= not (a xor b);
    outputs(1618) <= not (a or b);
    outputs(1619) <= a and b;
    outputs(1620) <= not b or a;
    outputs(1621) <= not (a xor b);
    outputs(1622) <= a and b;
    outputs(1623) <= '0';
    outputs(1624) <= not (a xor b);
    outputs(1625) <= a and b;
    outputs(1626) <= a and not b;
    outputs(1627) <= b and not a;
    outputs(1628) <= not a;
    outputs(1629) <= not a;
    outputs(1630) <= a and b;
    outputs(1631) <= a and b;
    outputs(1632) <= b;
    outputs(1633) <= b;
    outputs(1634) <= not (a xor b);
    outputs(1635) <= not b;
    outputs(1636) <= not a;
    outputs(1637) <= a;
    outputs(1638) <= not b;
    outputs(1639) <= a and not b;
    outputs(1640) <= not (a xor b);
    outputs(1641) <= a;
    outputs(1642) <= a xor b;
    outputs(1643) <= not (a or b);
    outputs(1644) <= a xor b;
    outputs(1645) <= '0';
    outputs(1646) <= not (a xor b);
    outputs(1647) <= '0';
    outputs(1648) <= b;
    outputs(1649) <= not (a or b);
    outputs(1650) <= not (a or b);
    outputs(1651) <= a and b;
    outputs(1652) <= a xor b;
    outputs(1653) <= not (a xor b);
    outputs(1654) <= not (a or b);
    outputs(1655) <= not b;
    outputs(1656) <= a;
    outputs(1657) <= b and not a;
    outputs(1658) <= not a;
    outputs(1659) <= a and b;
    outputs(1660) <= not a;
    outputs(1661) <= b and not a;
    outputs(1662) <= a xor b;
    outputs(1663) <= a and b;
    outputs(1664) <= a xor b;
    outputs(1665) <= b;
    outputs(1666) <= a xor b;
    outputs(1667) <= b and not a;
    outputs(1668) <= '0';
    outputs(1669) <= a and not b;
    outputs(1670) <= a and not b;
    outputs(1671) <= not (a xor b);
    outputs(1672) <= a and b;
    outputs(1673) <= a xor b;
    outputs(1674) <= not a;
    outputs(1675) <= b and not a;
    outputs(1676) <= not b;
    outputs(1677) <= not b;
    outputs(1678) <= not (a or b);
    outputs(1679) <= a and b;
    outputs(1680) <= a;
    outputs(1681) <= a and b;
    outputs(1682) <= a and b;
    outputs(1683) <= a and not b;
    outputs(1684) <= a xor b;
    outputs(1685) <= a and b;
    outputs(1686) <= b and not a;
    outputs(1687) <= a and not b;
    outputs(1688) <= a;
    outputs(1689) <= a and not b;
    outputs(1690) <= a and not b;
    outputs(1691) <= b and not a;
    outputs(1692) <= not (a xor b);
    outputs(1693) <= not (a or b);
    outputs(1694) <= a and b;
    outputs(1695) <= not b or a;
    outputs(1696) <= not (a or b);
    outputs(1697) <= not (a or b);
    outputs(1698) <= b;
    outputs(1699) <= b;
    outputs(1700) <= a xor b;
    outputs(1701) <= a xor b;
    outputs(1702) <= a and b;
    outputs(1703) <= a and not b;
    outputs(1704) <= not (a or b);
    outputs(1705) <= not (a or b);
    outputs(1706) <= not b;
    outputs(1707) <= a xor b;
    outputs(1708) <= a xor b;
    outputs(1709) <= a and b;
    outputs(1710) <= a and b;
    outputs(1711) <= not a or b;
    outputs(1712) <= not (a or b);
    outputs(1713) <= b and not a;
    outputs(1714) <= not (a xor b);
    outputs(1715) <= not (a or b);
    outputs(1716) <= not b;
    outputs(1717) <= a and b;
    outputs(1718) <= not b;
    outputs(1719) <= b and not a;
    outputs(1720) <= a xor b;
    outputs(1721) <= not a;
    outputs(1722) <= not b;
    outputs(1723) <= not a;
    outputs(1724) <= not a;
    outputs(1725) <= not b;
    outputs(1726) <= not b;
    outputs(1727) <= a and not b;
    outputs(1728) <= a;
    outputs(1729) <= a xor b;
    outputs(1730) <= not a;
    outputs(1731) <= b and not a;
    outputs(1732) <= a and b;
    outputs(1733) <= not (a xor b);
    outputs(1734) <= a and not b;
    outputs(1735) <= a and not b;
    outputs(1736) <= b and not a;
    outputs(1737) <= a and not b;
    outputs(1738) <= '0';
    outputs(1739) <= not b;
    outputs(1740) <= not (a xor b);
    outputs(1741) <= b and not a;
    outputs(1742) <= '0';
    outputs(1743) <= not (a or b);
    outputs(1744) <= not (a or b);
    outputs(1745) <= a and b;
    outputs(1746) <= not b;
    outputs(1747) <= not a or b;
    outputs(1748) <= b and not a;
    outputs(1749) <= '0';
    outputs(1750) <= not (a or b);
    outputs(1751) <= not (a xor b);
    outputs(1752) <= not a;
    outputs(1753) <= b and not a;
    outputs(1754) <= a xor b;
    outputs(1755) <= a and b;
    outputs(1756) <= a;
    outputs(1757) <= b and not a;
    outputs(1758) <= not (a or b);
    outputs(1759) <= not (a or b);
    outputs(1760) <= b and not a;
    outputs(1761) <= a and not b;
    outputs(1762) <= a xor b;
    outputs(1763) <= b and not a;
    outputs(1764) <= not a;
    outputs(1765) <= not (a xor b);
    outputs(1766) <= not (a or b);
    outputs(1767) <= a;
    outputs(1768) <= a and not b;
    outputs(1769) <= b;
    outputs(1770) <= a and b;
    outputs(1771) <= a;
    outputs(1772) <= b and not a;
    outputs(1773) <= b and not a;
    outputs(1774) <= not (a or b);
    outputs(1775) <= a;
    outputs(1776) <= a;
    outputs(1777) <= not (a or b);
    outputs(1778) <= a and b;
    outputs(1779) <= a;
    outputs(1780) <= not (a xor b);
    outputs(1781) <= not (a xor b);
    outputs(1782) <= b and not a;
    outputs(1783) <= not (a xor b);
    outputs(1784) <= b and not a;
    outputs(1785) <= a and b;
    outputs(1786) <= a and b;
    outputs(1787) <= not b;
    outputs(1788) <= a;
    outputs(1789) <= b;
    outputs(1790) <= a and not b;
    outputs(1791) <= not (a or b);
    outputs(1792) <= not b;
    outputs(1793) <= not (a or b);
    outputs(1794) <= a and not b;
    outputs(1795) <= a;
    outputs(1796) <= a and not b;
    outputs(1797) <= b and not a;
    outputs(1798) <= '0';
    outputs(1799) <= a;
    outputs(1800) <= a xor b;
    outputs(1801) <= b;
    outputs(1802) <= b;
    outputs(1803) <= not (a or b);
    outputs(1804) <= b and not a;
    outputs(1805) <= a and not b;
    outputs(1806) <= not (a xor b);
    outputs(1807) <= not (a or b);
    outputs(1808) <= a and b;
    outputs(1809) <= a xor b;
    outputs(1810) <= not (a xor b);
    outputs(1811) <= a and not b;
    outputs(1812) <= not (a or b);
    outputs(1813) <= a and b;
    outputs(1814) <= b and not a;
    outputs(1815) <= a and b;
    outputs(1816) <= not b;
    outputs(1817) <= not a;
    outputs(1818) <= b and not a;
    outputs(1819) <= b and not a;
    outputs(1820) <= a and b;
    outputs(1821) <= not b;
    outputs(1822) <= not a;
    outputs(1823) <= b and not a;
    outputs(1824) <= not (a or b);
    outputs(1825) <= a xor b;
    outputs(1826) <= a and b;
    outputs(1827) <= not a;
    outputs(1828) <= not (a or b);
    outputs(1829) <= a and b;
    outputs(1830) <= a and b;
    outputs(1831) <= b and not a;
    outputs(1832) <= not (a or b);
    outputs(1833) <= a and b;
    outputs(1834) <= b and not a;
    outputs(1835) <= not a;
    outputs(1836) <= a and not b;
    outputs(1837) <= b and not a;
    outputs(1838) <= b and not a;
    outputs(1839) <= not (a and b);
    outputs(1840) <= a or b;
    outputs(1841) <= not (a xor b);
    outputs(1842) <= a;
    outputs(1843) <= '0';
    outputs(1844) <= a and not b;
    outputs(1845) <= a and b;
    outputs(1846) <= not b;
    outputs(1847) <= not b;
    outputs(1848) <= not (a or b);
    outputs(1849) <= not (a xor b);
    outputs(1850) <= a xor b;
    outputs(1851) <= b;
    outputs(1852) <= a;
    outputs(1853) <= not (a xor b);
    outputs(1854) <= not (a xor b);
    outputs(1855) <= not (a or b);
    outputs(1856) <= not a;
    outputs(1857) <= not b;
    outputs(1858) <= a and b;
    outputs(1859) <= a and b;
    outputs(1860) <= a and b;
    outputs(1861) <= not a;
    outputs(1862) <= a xor b;
    outputs(1863) <= a and b;
    outputs(1864) <= b and not a;
    outputs(1865) <= not (a xor b);
    outputs(1866) <= not (a xor b);
    outputs(1867) <= a and b;
    outputs(1868) <= a and b;
    outputs(1869) <= not (a or b);
    outputs(1870) <= '0';
    outputs(1871) <= not b;
    outputs(1872) <= a and not b;
    outputs(1873) <= a xor b;
    outputs(1874) <= '0';
    outputs(1875) <= not (a or b);
    outputs(1876) <= not (a or b);
    outputs(1877) <= b;
    outputs(1878) <= not b;
    outputs(1879) <= b and not a;
    outputs(1880) <= a and not b;
    outputs(1881) <= a and not b;
    outputs(1882) <= a and b;
    outputs(1883) <= a and b;
    outputs(1884) <= b and not a;
    outputs(1885) <= b;
    outputs(1886) <= not (a or b);
    outputs(1887) <= not a or b;
    outputs(1888) <= not (a xor b);
    outputs(1889) <= not a;
    outputs(1890) <= a;
    outputs(1891) <= a and not b;
    outputs(1892) <= a and not b;
    outputs(1893) <= not (a or b);
    outputs(1894) <= a and b;
    outputs(1895) <= not a;
    outputs(1896) <= a and b;
    outputs(1897) <= a;
    outputs(1898) <= not b;
    outputs(1899) <= b;
    outputs(1900) <= a xor b;
    outputs(1901) <= not (a or b);
    outputs(1902) <= a and not b;
    outputs(1903) <= a and not b;
    outputs(1904) <= not b;
    outputs(1905) <= not (a or b);
    outputs(1906) <= b and not a;
    outputs(1907) <= a and not b;
    outputs(1908) <= a and not b;
    outputs(1909) <= not (a or b);
    outputs(1910) <= '0';
    outputs(1911) <= not (a xor b);
    outputs(1912) <= b and not a;
    outputs(1913) <= not a;
    outputs(1914) <= a and b;
    outputs(1915) <= b and not a;
    outputs(1916) <= a and b;
    outputs(1917) <= a xor b;
    outputs(1918) <= a;
    outputs(1919) <= a and b;
    outputs(1920) <= a and b;
    outputs(1921) <= b and not a;
    outputs(1922) <= b;
    outputs(1923) <= a and not b;
    outputs(1924) <= b and not a;
    outputs(1925) <= b and not a;
    outputs(1926) <= a and b;
    outputs(1927) <= a xor b;
    outputs(1928) <= a;
    outputs(1929) <= a;
    outputs(1930) <= a and not b;
    outputs(1931) <= '0';
    outputs(1932) <= a and not b;
    outputs(1933) <= not (a or b);
    outputs(1934) <= a xor b;
    outputs(1935) <= not b;
    outputs(1936) <= a xor b;
    outputs(1937) <= not a;
    outputs(1938) <= b and not a;
    outputs(1939) <= not a;
    outputs(1940) <= b;
    outputs(1941) <= a;
    outputs(1942) <= a and b;
    outputs(1943) <= a and not b;
    outputs(1944) <= a and not b;
    outputs(1945) <= not (a or b);
    outputs(1946) <= a and not b;
    outputs(1947) <= a and b;
    outputs(1948) <= a and not b;
    outputs(1949) <= not a;
    outputs(1950) <= b and not a;
    outputs(1951) <= b and not a;
    outputs(1952) <= not (a or b);
    outputs(1953) <= a;
    outputs(1954) <= b;
    outputs(1955) <= not (a or b);
    outputs(1956) <= not (a or b);
    outputs(1957) <= not b;
    outputs(1958) <= a and not b;
    outputs(1959) <= b and not a;
    outputs(1960) <= a and not b;
    outputs(1961) <= a and not b;
    outputs(1962) <= not (a or b);
    outputs(1963) <= b;
    outputs(1964) <= not b;
    outputs(1965) <= b and not a;
    outputs(1966) <= a and not b;
    outputs(1967) <= not (a or b);
    outputs(1968) <= a or b;
    outputs(1969) <= not b;
    outputs(1970) <= a xor b;
    outputs(1971) <= b and not a;
    outputs(1972) <= not a;
    outputs(1973) <= not (a or b);
    outputs(1974) <= b and not a;
    outputs(1975) <= b;
    outputs(1976) <= a xor b;
    outputs(1977) <= a;
    outputs(1978) <= not (a xor b);
    outputs(1979) <= b;
    outputs(1980) <= not (a or b);
    outputs(1981) <= b and not a;
    outputs(1982) <= a xor b;
    outputs(1983) <= b and not a;
    outputs(1984) <= a and b;
    outputs(1985) <= not (a or b);
    outputs(1986) <= a xor b;
    outputs(1987) <= a xor b;
    outputs(1988) <= not (a or b);
    outputs(1989) <= not (a xor b);
    outputs(1990) <= not (a or b);
    outputs(1991) <= not b;
    outputs(1992) <= not (a xor b);
    outputs(1993) <= not (a xor b);
    outputs(1994) <= a and not b;
    outputs(1995) <= a;
    outputs(1996) <= not (a and b);
    outputs(1997) <= not (a or b);
    outputs(1998) <= not (a xor b);
    outputs(1999) <= not (a or b);
    outputs(2000) <= '0';
    outputs(2001) <= b and not a;
    outputs(2002) <= b;
    outputs(2003) <= a and not b;
    outputs(2004) <= not (a or b);
    outputs(2005) <= b;
    outputs(2006) <= not (a xor b);
    outputs(2007) <= not (a xor b);
    outputs(2008) <= '0';
    outputs(2009) <= a;
    outputs(2010) <= a and not b;
    outputs(2011) <= a and b;
    outputs(2012) <= a xor b;
    outputs(2013) <= a;
    outputs(2014) <= a and not b;
    outputs(2015) <= a and not b;
    outputs(2016) <= '0';
    outputs(2017) <= not a;
    outputs(2018) <= b;
    outputs(2019) <= '0';
    outputs(2020) <= not (a or b);
    outputs(2021) <= not (a xor b);
    outputs(2022) <= a and not b;
    outputs(2023) <= not (a or b);
    outputs(2024) <= not (a xor b);
    outputs(2025) <= not b;
    outputs(2026) <= not a;
    outputs(2027) <= a or b;
    outputs(2028) <= not a;
    outputs(2029) <= not (a or b);
    outputs(2030) <= a and not b;
    outputs(2031) <= b and not a;
    outputs(2032) <= a and b;
    outputs(2033) <= b;
    outputs(2034) <= not a;
    outputs(2035) <= a xor b;
    outputs(2036) <= a and not b;
    outputs(2037) <= not a;
    outputs(2038) <= not (a or b);
    outputs(2039) <= a xor b;
    outputs(2040) <= not b;
    outputs(2041) <= not a;
    outputs(2042) <= not b;
    outputs(2043) <= a and not b;
    outputs(2044) <= a and not b;
    outputs(2045) <= a and b;
    outputs(2046) <= b and not a;
    outputs(2047) <= b and not a;
    outputs(2048) <= not a;
    outputs(2049) <= b;
    outputs(2050) <= a xor b;
    outputs(2051) <= not (a xor b);
    outputs(2052) <= a xor b;
    outputs(2053) <= b;
    outputs(2054) <= not (a xor b);
    outputs(2055) <= not (a xor b);
    outputs(2056) <= a or b;
    outputs(2057) <= not (a xor b);
    outputs(2058) <= a xor b;
    outputs(2059) <= not (a or b);
    outputs(2060) <= a and not b;
    outputs(2061) <= not (a xor b);
    outputs(2062) <= a or b;
    outputs(2063) <= a and not b;
    outputs(2064) <= not (a or b);
    outputs(2065) <= a xor b;
    outputs(2066) <= not a or b;
    outputs(2067) <= a and b;
    outputs(2068) <= not (a xor b);
    outputs(2069) <= a and not b;
    outputs(2070) <= not (a and b);
    outputs(2071) <= not (a and b);
    outputs(2072) <= b and not a;
    outputs(2073) <= not a;
    outputs(2074) <= a;
    outputs(2075) <= not (a or b);
    outputs(2076) <= a xor b;
    outputs(2077) <= a xor b;
    outputs(2078) <= a;
    outputs(2079) <= a;
    outputs(2080) <= not a or b;
    outputs(2081) <= a xor b;
    outputs(2082) <= not a;
    outputs(2083) <= a xor b;
    outputs(2084) <= not (a and b);
    outputs(2085) <= a;
    outputs(2086) <= not (a xor b);
    outputs(2087) <= b;
    outputs(2088) <= not (a xor b);
    outputs(2089) <= b;
    outputs(2090) <= a or b;
    outputs(2091) <= not a or b;
    outputs(2092) <= not (a xor b);
    outputs(2093) <= a and not b;
    outputs(2094) <= not b;
    outputs(2095) <= not (a xor b);
    outputs(2096) <= not a or b;
    outputs(2097) <= not (a or b);
    outputs(2098) <= a;
    outputs(2099) <= b and not a;
    outputs(2100) <= a;
    outputs(2101) <= not (a and b);
    outputs(2102) <= a xor b;
    outputs(2103) <= not (a or b);
    outputs(2104) <= not (a and b);
    outputs(2105) <= not (a and b);
    outputs(2106) <= not a;
    outputs(2107) <= a;
    outputs(2108) <= b;
    outputs(2109) <= not (a xor b);
    outputs(2110) <= a;
    outputs(2111) <= a;
    outputs(2112) <= not a or b;
    outputs(2113) <= not b;
    outputs(2114) <= b;
    outputs(2115) <= b;
    outputs(2116) <= not b;
    outputs(2117) <= a;
    outputs(2118) <= b;
    outputs(2119) <= a or b;
    outputs(2120) <= not (a xor b);
    outputs(2121) <= not (a xor b);
    outputs(2122) <= a and b;
    outputs(2123) <= b;
    outputs(2124) <= not b;
    outputs(2125) <= not b;
    outputs(2126) <= b and not a;
    outputs(2127) <= not b;
    outputs(2128) <= a xor b;
    outputs(2129) <= not b;
    outputs(2130) <= a xor b;
    outputs(2131) <= a and b;
    outputs(2132) <= a;
    outputs(2133) <= b and not a;
    outputs(2134) <= not (a and b);
    outputs(2135) <= b and not a;
    outputs(2136) <= not a;
    outputs(2137) <= a;
    outputs(2138) <= a or b;
    outputs(2139) <= a and b;
    outputs(2140) <= not b;
    outputs(2141) <= a xor b;
    outputs(2142) <= not (a and b);
    outputs(2143) <= not (a xor b);
    outputs(2144) <= a xor b;
    outputs(2145) <= a xor b;
    outputs(2146) <= not (a and b);
    outputs(2147) <= not a;
    outputs(2148) <= not (a xor b);
    outputs(2149) <= b;
    outputs(2150) <= not a;
    outputs(2151) <= not b or a;
    outputs(2152) <= not (a xor b);
    outputs(2153) <= a xor b;
    outputs(2154) <= b and not a;
    outputs(2155) <= not (a xor b);
    outputs(2156) <= not (a and b);
    outputs(2157) <= not (a xor b);
    outputs(2158) <= not a;
    outputs(2159) <= not a;
    outputs(2160) <= not b;
    outputs(2161) <= not b or a;
    outputs(2162) <= b;
    outputs(2163) <= not a;
    outputs(2164) <= a or b;
    outputs(2165) <= not a or b;
    outputs(2166) <= a xor b;
    outputs(2167) <= not b or a;
    outputs(2168) <= not (a xor b);
    outputs(2169) <= b;
    outputs(2170) <= not b;
    outputs(2171) <= a and b;
    outputs(2172) <= a xor b;
    outputs(2173) <= not a;
    outputs(2174) <= not (a xor b);
    outputs(2175) <= not a or b;
    outputs(2176) <= a;
    outputs(2177) <= not (a and b);
    outputs(2178) <= a xor b;
    outputs(2179) <= not (a xor b);
    outputs(2180) <= b and not a;
    outputs(2181) <= a xor b;
    outputs(2182) <= a xor b;
    outputs(2183) <= not b or a;
    outputs(2184) <= a xor b;
    outputs(2185) <= not (a xor b);
    outputs(2186) <= a xor b;
    outputs(2187) <= a;
    outputs(2188) <= a xor b;
    outputs(2189) <= a and not b;
    outputs(2190) <= not b;
    outputs(2191) <= not b;
    outputs(2192) <= a and b;
    outputs(2193) <= b;
    outputs(2194) <= a;
    outputs(2195) <= not b;
    outputs(2196) <= not b;
    outputs(2197) <= not (a or b);
    outputs(2198) <= not (a xor b);
    outputs(2199) <= a xor b;
    outputs(2200) <= a xor b;
    outputs(2201) <= not (a xor b);
    outputs(2202) <= not a;
    outputs(2203) <= not (a xor b);
    outputs(2204) <= not (a and b);
    outputs(2205) <= a;
    outputs(2206) <= not (a and b);
    outputs(2207) <= not a or b;
    outputs(2208) <= a;
    outputs(2209) <= not a;
    outputs(2210) <= a;
    outputs(2211) <= a xor b;
    outputs(2212) <= b;
    outputs(2213) <= b;
    outputs(2214) <= a xor b;
    outputs(2215) <= not a or b;
    outputs(2216) <= not a;
    outputs(2217) <= a and not b;
    outputs(2218) <= not b or a;
    outputs(2219) <= not (a xor b);
    outputs(2220) <= not b;
    outputs(2221) <= not a;
    outputs(2222) <= not (a xor b);
    outputs(2223) <= a xor b;
    outputs(2224) <= a;
    outputs(2225) <= a and not b;
    outputs(2226) <= not (a xor b);
    outputs(2227) <= b;
    outputs(2228) <= b;
    outputs(2229) <= not b;
    outputs(2230) <= '1';
    outputs(2231) <= not b;
    outputs(2232) <= a xor b;
    outputs(2233) <= not (a xor b);
    outputs(2234) <= a and b;
    outputs(2235) <= not (a xor b);
    outputs(2236) <= not (a xor b);
    outputs(2237) <= a and not b;
    outputs(2238) <= a and not b;
    outputs(2239) <= a;
    outputs(2240) <= not b or a;
    outputs(2241) <= not b or a;
    outputs(2242) <= a xor b;
    outputs(2243) <= a xor b;
    outputs(2244) <= not (a xor b);
    outputs(2245) <= not (a and b);
    outputs(2246) <= not (a xor b);
    outputs(2247) <= b;
    outputs(2248) <= not a;
    outputs(2249) <= a and not b;
    outputs(2250) <= a;
    outputs(2251) <= not (a xor b);
    outputs(2252) <= b;
    outputs(2253) <= a xor b;
    outputs(2254) <= not a;
    outputs(2255) <= not (a xor b);
    outputs(2256) <= not b or a;
    outputs(2257) <= a or b;
    outputs(2258) <= not (a xor b);
    outputs(2259) <= a and not b;
    outputs(2260) <= not b;
    outputs(2261) <= a and not b;
    outputs(2262) <= not (a xor b);
    outputs(2263) <= not b;
    outputs(2264) <= not (a xor b);
    outputs(2265) <= not (a xor b);
    outputs(2266) <= b;
    outputs(2267) <= not a;
    outputs(2268) <= not b;
    outputs(2269) <= not (a and b);
    outputs(2270) <= a;
    outputs(2271) <= not b;
    outputs(2272) <= not b or a;
    outputs(2273) <= a xor b;
    outputs(2274) <= not (a xor b);
    outputs(2275) <= b;
    outputs(2276) <= not a or b;
    outputs(2277) <= a;
    outputs(2278) <= a xor b;
    outputs(2279) <= not (a and b);
    outputs(2280) <= a and not b;
    outputs(2281) <= not (a xor b);
    outputs(2282) <= not b or a;
    outputs(2283) <= b;
    outputs(2284) <= not b;
    outputs(2285) <= b;
    outputs(2286) <= not b;
    outputs(2287) <= not a or b;
    outputs(2288) <= b and not a;
    outputs(2289) <= not b;
    outputs(2290) <= a xor b;
    outputs(2291) <= a and b;
    outputs(2292) <= not a;
    outputs(2293) <= not b;
    outputs(2294) <= not a or b;
    outputs(2295) <= not (a or b);
    outputs(2296) <= a;
    outputs(2297) <= not b;
    outputs(2298) <= not (a xor b);
    outputs(2299) <= not a or b;
    outputs(2300) <= a;
    outputs(2301) <= not (a and b);
    outputs(2302) <= a xor b;
    outputs(2303) <= not b;
    outputs(2304) <= not b or a;
    outputs(2305) <= not a;
    outputs(2306) <= not (a xor b);
    outputs(2307) <= not (a xor b);
    outputs(2308) <= a xor b;
    outputs(2309) <= b;
    outputs(2310) <= not (a xor b);
    outputs(2311) <= not a or b;
    outputs(2312) <= a and not b;
    outputs(2313) <= not b;
    outputs(2314) <= b;
    outputs(2315) <= not b;
    outputs(2316) <= b and not a;
    outputs(2317) <= not a;
    outputs(2318) <= not a;
    outputs(2319) <= b;
    outputs(2320) <= not (a xor b);
    outputs(2321) <= b;
    outputs(2322) <= a;
    outputs(2323) <= not a;
    outputs(2324) <= not (a or b);
    outputs(2325) <= not b or a;
    outputs(2326) <= not a or b;
    outputs(2327) <= not (a xor b);
    outputs(2328) <= a;
    outputs(2329) <= a xor b;
    outputs(2330) <= a;
    outputs(2331) <= a or b;
    outputs(2332) <= not b or a;
    outputs(2333) <= not (a and b);
    outputs(2334) <= not (a xor b);
    outputs(2335) <= b and not a;
    outputs(2336) <= a;
    outputs(2337) <= not a;
    outputs(2338) <= not (a xor b);
    outputs(2339) <= a and not b;
    outputs(2340) <= not a;
    outputs(2341) <= a or b;
    outputs(2342) <= not a;
    outputs(2343) <= not (a xor b);
    outputs(2344) <= not (a xor b);
    outputs(2345) <= a;
    outputs(2346) <= b and not a;
    outputs(2347) <= b and not a;
    outputs(2348) <= a xor b;
    outputs(2349) <= b;
    outputs(2350) <= not (a xor b);
    outputs(2351) <= b;
    outputs(2352) <= a and b;
    outputs(2353) <= b;
    outputs(2354) <= a and not b;
    outputs(2355) <= not a;
    outputs(2356) <= a;
    outputs(2357) <= not (a xor b);
    outputs(2358) <= a;
    outputs(2359) <= a;
    outputs(2360) <= not a or b;
    outputs(2361) <= a and b;
    outputs(2362) <= b;
    outputs(2363) <= b;
    outputs(2364) <= a or b;
    outputs(2365) <= b;
    outputs(2366) <= a xor b;
    outputs(2367) <= not (a or b);
    outputs(2368) <= b;
    outputs(2369) <= a xor b;
    outputs(2370) <= not (a and b);
    outputs(2371) <= a xor b;
    outputs(2372) <= not b;
    outputs(2373) <= not (a xor b);
    outputs(2374) <= not a or b;
    outputs(2375) <= not b;
    outputs(2376) <= a xor b;
    outputs(2377) <= a;
    outputs(2378) <= not b;
    outputs(2379) <= b;
    outputs(2380) <= b;
    outputs(2381) <= a xor b;
    outputs(2382) <= a xor b;
    outputs(2383) <= not a;
    outputs(2384) <= not (a xor b);
    outputs(2385) <= not (a and b);
    outputs(2386) <= not b or a;
    outputs(2387) <= not (a xor b);
    outputs(2388) <= a xor b;
    outputs(2389) <= b;
    outputs(2390) <= b and not a;
    outputs(2391) <= a xor b;
    outputs(2392) <= not (a xor b);
    outputs(2393) <= not a or b;
    outputs(2394) <= a;
    outputs(2395) <= not b;
    outputs(2396) <= a;
    outputs(2397) <= not (a and b);
    outputs(2398) <= not (a xor b);
    outputs(2399) <= not a;
    outputs(2400) <= not a;
    outputs(2401) <= not b or a;
    outputs(2402) <= not b;
    outputs(2403) <= not (a or b);
    outputs(2404) <= a xor b;
    outputs(2405) <= not (a and b);
    outputs(2406) <= a xor b;
    outputs(2407) <= a xor b;
    outputs(2408) <= a xor b;
    outputs(2409) <= a or b;
    outputs(2410) <= not (a xor b);
    outputs(2411) <= b and not a;
    outputs(2412) <= a xor b;
    outputs(2413) <= not a;
    outputs(2414) <= a xor b;
    outputs(2415) <= a or b;
    outputs(2416) <= a xor b;
    outputs(2417) <= not b;
    outputs(2418) <= not (a xor b);
    outputs(2419) <= a xor b;
    outputs(2420) <= not a or b;
    outputs(2421) <= not (a or b);
    outputs(2422) <= a or b;
    outputs(2423) <= not (a and b);
    outputs(2424) <= a;
    outputs(2425) <= not (a and b);
    outputs(2426) <= not b or a;
    outputs(2427) <= not (a and b);
    outputs(2428) <= not (a xor b);
    outputs(2429) <= not a;
    outputs(2430) <= a and b;
    outputs(2431) <= a or b;
    outputs(2432) <= a xor b;
    outputs(2433) <= not (a xor b);
    outputs(2434) <= a xor b;
    outputs(2435) <= a or b;
    outputs(2436) <= a;
    outputs(2437) <= not b;
    outputs(2438) <= a xor b;
    outputs(2439) <= b;
    outputs(2440) <= not (a and b);
    outputs(2441) <= a xor b;
    outputs(2442) <= a;
    outputs(2443) <= not (a xor b);
    outputs(2444) <= a or b;
    outputs(2445) <= a and not b;
    outputs(2446) <= not (a xor b);
    outputs(2447) <= not (a xor b);
    outputs(2448) <= not a;
    outputs(2449) <= not a;
    outputs(2450) <= not b;
    outputs(2451) <= not (a and b);
    outputs(2452) <= not b or a;
    outputs(2453) <= not b or a;
    outputs(2454) <= a;
    outputs(2455) <= not b or a;
    outputs(2456) <= not a;
    outputs(2457) <= not a;
    outputs(2458) <= b;
    outputs(2459) <= not a;
    outputs(2460) <= a and not b;
    outputs(2461) <= a xor b;
    outputs(2462) <= not (a xor b);
    outputs(2463) <= not (a or b);
    outputs(2464) <= b;
    outputs(2465) <= not (a xor b);
    outputs(2466) <= a xor b;
    outputs(2467) <= a and b;
    outputs(2468) <= not (a or b);
    outputs(2469) <= not (a xor b);
    outputs(2470) <= not (a and b);
    outputs(2471) <= a;
    outputs(2472) <= not a or b;
    outputs(2473) <= not (a xor b);
    outputs(2474) <= not (a xor b);
    outputs(2475) <= not a;
    outputs(2476) <= b;
    outputs(2477) <= not (a and b);
    outputs(2478) <= a;
    outputs(2479) <= not a or b;
    outputs(2480) <= b and not a;
    outputs(2481) <= a;
    outputs(2482) <= b and not a;
    outputs(2483) <= a;
    outputs(2484) <= not (a xor b);
    outputs(2485) <= not (a and b);
    outputs(2486) <= not (a xor b);
    outputs(2487) <= not (a xor b);
    outputs(2488) <= not (a and b);
    outputs(2489) <= not b;
    outputs(2490) <= not (a xor b);
    outputs(2491) <= a xor b;
    outputs(2492) <= a and b;
    outputs(2493) <= a or b;
    outputs(2494) <= a and not b;
    outputs(2495) <= not b;
    outputs(2496) <= not (a xor b);
    outputs(2497) <= not b or a;
    outputs(2498) <= a xor b;
    outputs(2499) <= a and b;
    outputs(2500) <= a and not b;
    outputs(2501) <= not (a and b);
    outputs(2502) <= not (a xor b);
    outputs(2503) <= not a;
    outputs(2504) <= not b;
    outputs(2505) <= a and b;
    outputs(2506) <= not b;
    outputs(2507) <= a or b;
    outputs(2508) <= not (a xor b);
    outputs(2509) <= a xor b;
    outputs(2510) <= not b;
    outputs(2511) <= b;
    outputs(2512) <= not a;
    outputs(2513) <= not b;
    outputs(2514) <= b;
    outputs(2515) <= not b;
    outputs(2516) <= b;
    outputs(2517) <= a xor b;
    outputs(2518) <= not a;
    outputs(2519) <= not b;
    outputs(2520) <= a xor b;
    outputs(2521) <= not (a xor b);
    outputs(2522) <= not b;
    outputs(2523) <= a or b;
    outputs(2524) <= a xor b;
    outputs(2525) <= not (a xor b);
    outputs(2526) <= a;
    outputs(2527) <= not b or a;
    outputs(2528) <= a;
    outputs(2529) <= not b;
    outputs(2530) <= a xor b;
    outputs(2531) <= not b or a;
    outputs(2532) <= a and not b;
    outputs(2533) <= not a or b;
    outputs(2534) <= not b;
    outputs(2535) <= a and not b;
    outputs(2536) <= a;
    outputs(2537) <= b;
    outputs(2538) <= a and b;
    outputs(2539) <= b;
    outputs(2540) <= not (a and b);
    outputs(2541) <= b and not a;
    outputs(2542) <= not (a and b);
    outputs(2543) <= not (a xor b);
    outputs(2544) <= b;
    outputs(2545) <= a and b;
    outputs(2546) <= a;
    outputs(2547) <= b;
    outputs(2548) <= b and not a;
    outputs(2549) <= not (a and b);
    outputs(2550) <= a;
    outputs(2551) <= not b or a;
    outputs(2552) <= a;
    outputs(2553) <= a xor b;
    outputs(2554) <= not (a xor b);
    outputs(2555) <= not (a and b);
    outputs(2556) <= not (a xor b);
    outputs(2557) <= a;
    outputs(2558) <= a or b;
    outputs(2559) <= not (a and b);
    outputs(2560) <= a;
    outputs(2561) <= a or b;
    outputs(2562) <= a xor b;
    outputs(2563) <= not b;
    outputs(2564) <= not (a xor b);
    outputs(2565) <= not b;
    outputs(2566) <= not a or b;
    outputs(2567) <= a and b;
    outputs(2568) <= a;
    outputs(2569) <= not (a xor b);
    outputs(2570) <= not (a or b);
    outputs(2571) <= a;
    outputs(2572) <= a xor b;
    outputs(2573) <= not b;
    outputs(2574) <= not b;
    outputs(2575) <= not (a or b);
    outputs(2576) <= a;
    outputs(2577) <= b;
    outputs(2578) <= not (a xor b);
    outputs(2579) <= b;
    outputs(2580) <= not (a and b);
    outputs(2581) <= not (a xor b);
    outputs(2582) <= a xor b;
    outputs(2583) <= b;
    outputs(2584) <= not a;
    outputs(2585) <= not (a or b);
    outputs(2586) <= a xor b;
    outputs(2587) <= not b;
    outputs(2588) <= a;
    outputs(2589) <= not b or a;
    outputs(2590) <= not (a and b);
    outputs(2591) <= a;
    outputs(2592) <= not a;
    outputs(2593) <= b;
    outputs(2594) <= not b;
    outputs(2595) <= not a;
    outputs(2596) <= not b or a;
    outputs(2597) <= b;
    outputs(2598) <= not b;
    outputs(2599) <= not (a xor b);
    outputs(2600) <= not a;
    outputs(2601) <= a;
    outputs(2602) <= a or b;
    outputs(2603) <= a;
    outputs(2604) <= a or b;
    outputs(2605) <= not b or a;
    outputs(2606) <= not (a and b);
    outputs(2607) <= a xor b;
    outputs(2608) <= not b;
    outputs(2609) <= not b or a;
    outputs(2610) <= not b;
    outputs(2611) <= not (a xor b);
    outputs(2612) <= not b;
    outputs(2613) <= not b;
    outputs(2614) <= not b;
    outputs(2615) <= not (a and b);
    outputs(2616) <= not b;
    outputs(2617) <= not b or a;
    outputs(2618) <= not a;
    outputs(2619) <= not b;
    outputs(2620) <= a or b;
    outputs(2621) <= a;
    outputs(2622) <= not (a and b);
    outputs(2623) <= a or b;
    outputs(2624) <= not a;
    outputs(2625) <= a;
    outputs(2626) <= not b or a;
    outputs(2627) <= b;
    outputs(2628) <= not (a or b);
    outputs(2629) <= a;
    outputs(2630) <= not (a xor b);
    outputs(2631) <= a xor b;
    outputs(2632) <= not b;
    outputs(2633) <= a xor b;
    outputs(2634) <= a;
    outputs(2635) <= not b;
    outputs(2636) <= not b;
    outputs(2637) <= not (a or b);
    outputs(2638) <= not b;
    outputs(2639) <= b;
    outputs(2640) <= a xor b;
    outputs(2641) <= a xor b;
    outputs(2642) <= not b or a;
    outputs(2643) <= b;
    outputs(2644) <= not b;
    outputs(2645) <= not (a xor b);
    outputs(2646) <= not (a and b);
    outputs(2647) <= not (a xor b);
    outputs(2648) <= a xor b;
    outputs(2649) <= b and not a;
    outputs(2650) <= a;
    outputs(2651) <= not b;
    outputs(2652) <= not (a xor b);
    outputs(2653) <= '1';
    outputs(2654) <= not a or b;
    outputs(2655) <= a;
    outputs(2656) <= not a;
    outputs(2657) <= a or b;
    outputs(2658) <= a xor b;
    outputs(2659) <= a and b;
    outputs(2660) <= a or b;
    outputs(2661) <= not b;
    outputs(2662) <= not (a and b);
    outputs(2663) <= not a;
    outputs(2664) <= a xor b;
    outputs(2665) <= not (a xor b);
    outputs(2666) <= not b or a;
    outputs(2667) <= b;
    outputs(2668) <= a and b;
    outputs(2669) <= not (a and b);
    outputs(2670) <= a and not b;
    outputs(2671) <= not b;
    outputs(2672) <= not a;
    outputs(2673) <= b;
    outputs(2674) <= not (a xor b);
    outputs(2675) <= a;
    outputs(2676) <= not (a xor b);
    outputs(2677) <= not a or b;
    outputs(2678) <= b;
    outputs(2679) <= a or b;
    outputs(2680) <= a or b;
    outputs(2681) <= not a;
    outputs(2682) <= a;
    outputs(2683) <= not a;
    outputs(2684) <= not (a xor b);
    outputs(2685) <= not b;
    outputs(2686) <= a xor b;
    outputs(2687) <= not (a xor b);
    outputs(2688) <= b and not a;
    outputs(2689) <= not a or b;
    outputs(2690) <= not b;
    outputs(2691) <= b;
    outputs(2692) <= not b or a;
    outputs(2693) <= b;
    outputs(2694) <= b;
    outputs(2695) <= not b;
    outputs(2696) <= a xor b;
    outputs(2697) <= not (a xor b);
    outputs(2698) <= not b or a;
    outputs(2699) <= b and not a;
    outputs(2700) <= a xor b;
    outputs(2701) <= not b;
    outputs(2702) <= not (a xor b);
    outputs(2703) <= not b or a;
    outputs(2704) <= not (a xor b);
    outputs(2705) <= not a or b;
    outputs(2706) <= not (a and b);
    outputs(2707) <= not b;
    outputs(2708) <= not (a xor b);
    outputs(2709) <= a;
    outputs(2710) <= not (a xor b);
    outputs(2711) <= b;
    outputs(2712) <= a and not b;
    outputs(2713) <= b and not a;
    outputs(2714) <= not b;
    outputs(2715) <= not (a xor b);
    outputs(2716) <= a xor b;
    outputs(2717) <= not (a xor b);
    outputs(2718) <= a;
    outputs(2719) <= a xor b;
    outputs(2720) <= a;
    outputs(2721) <= not (a xor b);
    outputs(2722) <= not a;
    outputs(2723) <= a xor b;
    outputs(2724) <= a or b;
    outputs(2725) <= b;
    outputs(2726) <= not (a xor b);
    outputs(2727) <= not a;
    outputs(2728) <= not a;
    outputs(2729) <= a;
    outputs(2730) <= a;
    outputs(2731) <= b and not a;
    outputs(2732) <= not a;
    outputs(2733) <= not b;
    outputs(2734) <= b;
    outputs(2735) <= not b;
    outputs(2736) <= a xor b;
    outputs(2737) <= a;
    outputs(2738) <= a xor b;
    outputs(2739) <= not (a xor b);
    outputs(2740) <= not a or b;
    outputs(2741) <= a;
    outputs(2742) <= a xor b;
    outputs(2743) <= not a or b;
    outputs(2744) <= not (a xor b);
    outputs(2745) <= not b or a;
    outputs(2746) <= b and not a;
    outputs(2747) <= b;
    outputs(2748) <= a and b;
    outputs(2749) <= not b;
    outputs(2750) <= not a;
    outputs(2751) <= not (a and b);
    outputs(2752) <= b and not a;
    outputs(2753) <= a;
    outputs(2754) <= not b;
    outputs(2755) <= not a;
    outputs(2756) <= b and not a;
    outputs(2757) <= not (a xor b);
    outputs(2758) <= a xor b;
    outputs(2759) <= not a or b;
    outputs(2760) <= a or b;
    outputs(2761) <= not b or a;
    outputs(2762) <= not (a xor b);
    outputs(2763) <= a xor b;
    outputs(2764) <= not a;
    outputs(2765) <= not b;
    outputs(2766) <= a xor b;
    outputs(2767) <= not (a xor b);
    outputs(2768) <= not (a xor b);
    outputs(2769) <= a xor b;
    outputs(2770) <= a and not b;
    outputs(2771) <= a xor b;
    outputs(2772) <= not a;
    outputs(2773) <= not (a xor b);
    outputs(2774) <= b;
    outputs(2775) <= not (a and b);
    outputs(2776) <= a xor b;
    outputs(2777) <= not a;
    outputs(2778) <= b;
    outputs(2779) <= b;
    outputs(2780) <= a;
    outputs(2781) <= a;
    outputs(2782) <= a;
    outputs(2783) <= not (a or b);
    outputs(2784) <= a;
    outputs(2785) <= not b;
    outputs(2786) <= not (a or b);
    outputs(2787) <= not (a xor b);
    outputs(2788) <= not b;
    outputs(2789) <= not b;
    outputs(2790) <= a or b;
    outputs(2791) <= not (a xor b);
    outputs(2792) <= not (a and b);
    outputs(2793) <= not (a and b);
    outputs(2794) <= not (a or b);
    outputs(2795) <= a and b;
    outputs(2796) <= b;
    outputs(2797) <= not a;
    outputs(2798) <= a or b;
    outputs(2799) <= a;
    outputs(2800) <= b;
    outputs(2801) <= b;
    outputs(2802) <= not (a xor b);
    outputs(2803) <= a;
    outputs(2804) <= not (a xor b);
    outputs(2805) <= not b;
    outputs(2806) <= b;
    outputs(2807) <= a xor b;
    outputs(2808) <= not b;
    outputs(2809) <= a;
    outputs(2810) <= a;
    outputs(2811) <= a xor b;
    outputs(2812) <= b;
    outputs(2813) <= a;
    outputs(2814) <= not b;
    outputs(2815) <= not a;
    outputs(2816) <= not a;
    outputs(2817) <= a xor b;
    outputs(2818) <= not a;
    outputs(2819) <= a;
    outputs(2820) <= not b;
    outputs(2821) <= a;
    outputs(2822) <= not b;
    outputs(2823) <= b;
    outputs(2824) <= not a;
    outputs(2825) <= not a;
    outputs(2826) <= not (a xor b);
    outputs(2827) <= a or b;
    outputs(2828) <= not (a xor b);
    outputs(2829) <= not b;
    outputs(2830) <= not (a xor b);
    outputs(2831) <= not (a xor b);
    outputs(2832) <= a xor b;
    outputs(2833) <= a;
    outputs(2834) <= a xor b;
    outputs(2835) <= b and not a;
    outputs(2836) <= a xor b;
    outputs(2837) <= not (a xor b);
    outputs(2838) <= not b or a;
    outputs(2839) <= b and not a;
    outputs(2840) <= not (a or b);
    outputs(2841) <= a and not b;
    outputs(2842) <= not (a xor b);
    outputs(2843) <= not b;
    outputs(2844) <= b;
    outputs(2845) <= a;
    outputs(2846) <= a and b;
    outputs(2847) <= a or b;
    outputs(2848) <= a and not b;
    outputs(2849) <= b;
    outputs(2850) <= a xor b;
    outputs(2851) <= not a;
    outputs(2852) <= not b;
    outputs(2853) <= not (a and b);
    outputs(2854) <= not b or a;
    outputs(2855) <= b;
    outputs(2856) <= not a;
    outputs(2857) <= not (a xor b);
    outputs(2858) <= b;
    outputs(2859) <= not a;
    outputs(2860) <= not a;
    outputs(2861) <= a xor b;
    outputs(2862) <= not b;
    outputs(2863) <= a;
    outputs(2864) <= b;
    outputs(2865) <= a and not b;
    outputs(2866) <= not b;
    outputs(2867) <= a xor b;
    outputs(2868) <= not (a or b);
    outputs(2869) <= a and b;
    outputs(2870) <= not (a xor b);
    outputs(2871) <= not b or a;
    outputs(2872) <= not a;
    outputs(2873) <= a or b;
    outputs(2874) <= not (a and b);
    outputs(2875) <= b;
    outputs(2876) <= not a;
    outputs(2877) <= not (a xor b);
    outputs(2878) <= a;
    outputs(2879) <= a and not b;
    outputs(2880) <= not (a xor b);
    outputs(2881) <= a or b;
    outputs(2882) <= not b or a;
    outputs(2883) <= not a;
    outputs(2884) <= a and not b;
    outputs(2885) <= a and not b;
    outputs(2886) <= not a;
    outputs(2887) <= not a;
    outputs(2888) <= not (a xor b);
    outputs(2889) <= '0';
    outputs(2890) <= b;
    outputs(2891) <= b;
    outputs(2892) <= b;
    outputs(2893) <= a;
    outputs(2894) <= a xor b;
    outputs(2895) <= not b;
    outputs(2896) <= b;
    outputs(2897) <= not (a xor b);
    outputs(2898) <= not a;
    outputs(2899) <= a;
    outputs(2900) <= b and not a;
    outputs(2901) <= b;
    outputs(2902) <= not (a and b);
    outputs(2903) <= not b;
    outputs(2904) <= a;
    outputs(2905) <= not (a xor b);
    outputs(2906) <= not b;
    outputs(2907) <= not b;
    outputs(2908) <= not a;
    outputs(2909) <= not (a and b);
    outputs(2910) <= a and b;
    outputs(2911) <= a;
    outputs(2912) <= b and not a;
    outputs(2913) <= b and not a;
    outputs(2914) <= b;
    outputs(2915) <= not b or a;
    outputs(2916) <= not a;
    outputs(2917) <= not b;
    outputs(2918) <= not b;
    outputs(2919) <= a xor b;
    outputs(2920) <= not a or b;
    outputs(2921) <= a;
    outputs(2922) <= not a;
    outputs(2923) <= not a;
    outputs(2924) <= not a;
    outputs(2925) <= a or b;
    outputs(2926) <= a;
    outputs(2927) <= not (a xor b);
    outputs(2928) <= b;
    outputs(2929) <= a or b;
    outputs(2930) <= a;
    outputs(2931) <= a or b;
    outputs(2932) <= not a or b;
    outputs(2933) <= not (a xor b);
    outputs(2934) <= not (a xor b);
    outputs(2935) <= not (a xor b);
    outputs(2936) <= not (a xor b);
    outputs(2937) <= not a;
    outputs(2938) <= a xor b;
    outputs(2939) <= not a;
    outputs(2940) <= not b;
    outputs(2941) <= not a;
    outputs(2942) <= b;
    outputs(2943) <= a xor b;
    outputs(2944) <= a;
    outputs(2945) <= a or b;
    outputs(2946) <= a;
    outputs(2947) <= not a;
    outputs(2948) <= a;
    outputs(2949) <= not a or b;
    outputs(2950) <= a and not b;
    outputs(2951) <= a xor b;
    outputs(2952) <= a xor b;
    outputs(2953) <= not (a or b);
    outputs(2954) <= not a;
    outputs(2955) <= not (a or b);
    outputs(2956) <= a;
    outputs(2957) <= not b;
    outputs(2958) <= b;
    outputs(2959) <= not b;
    outputs(2960) <= not a;
    outputs(2961) <= a;
    outputs(2962) <= a xor b;
    outputs(2963) <= a xor b;
    outputs(2964) <= not a;
    outputs(2965) <= a;
    outputs(2966) <= a;
    outputs(2967) <= not (a and b);
    outputs(2968) <= a or b;
    outputs(2969) <= b;
    outputs(2970) <= a;
    outputs(2971) <= not (a and b);
    outputs(2972) <= not b;
    outputs(2973) <= not (a or b);
    outputs(2974) <= a or b;
    outputs(2975) <= not (a xor b);
    outputs(2976) <= a xor b;
    outputs(2977) <= not (a xor b);
    outputs(2978) <= a;
    outputs(2979) <= not b or a;
    outputs(2980) <= b and not a;
    outputs(2981) <= b;
    outputs(2982) <= not a;
    outputs(2983) <= not (a xor b);
    outputs(2984) <= a;
    outputs(2985) <= a xor b;
    outputs(2986) <= not b or a;
    outputs(2987) <= a or b;
    outputs(2988) <= b;
    outputs(2989) <= b and not a;
    outputs(2990) <= not (a xor b);
    outputs(2991) <= not b;
    outputs(2992) <= a or b;
    outputs(2993) <= a and b;
    outputs(2994) <= a xor b;
    outputs(2995) <= not a;
    outputs(2996) <= not (a xor b);
    outputs(2997) <= a;
    outputs(2998) <= b;
    outputs(2999) <= a or b;
    outputs(3000) <= not b;
    outputs(3001) <= a;
    outputs(3002) <= not a;
    outputs(3003) <= not (a or b);
    outputs(3004) <= a;
    outputs(3005) <= not (a xor b);
    outputs(3006) <= not (a xor b);
    outputs(3007) <= a;
    outputs(3008) <= b and not a;
    outputs(3009) <= a and b;
    outputs(3010) <= b and not a;
    outputs(3011) <= a or b;
    outputs(3012) <= b and not a;
    outputs(3013) <= a xor b;
    outputs(3014) <= not b;
    outputs(3015) <= a and b;
    outputs(3016) <= a;
    outputs(3017) <= a xor b;
    outputs(3018) <= a or b;
    outputs(3019) <= a;
    outputs(3020) <= not b;
    outputs(3021) <= not a;
    outputs(3022) <= not b;
    outputs(3023) <= a and not b;
    outputs(3024) <= not b;
    outputs(3025) <= not a;
    outputs(3026) <= not b;
    outputs(3027) <= a and not b;
    outputs(3028) <= not (a and b);
    outputs(3029) <= not b;
    outputs(3030) <= b and not a;
    outputs(3031) <= not b;
    outputs(3032) <= b;
    outputs(3033) <= not a or b;
    outputs(3034) <= a;
    outputs(3035) <= a;
    outputs(3036) <= not (a and b);
    outputs(3037) <= not b;
    outputs(3038) <= not b;
    outputs(3039) <= a;
    outputs(3040) <= not b;
    outputs(3041) <= not (a or b);
    outputs(3042) <= b;
    outputs(3043) <= a or b;
    outputs(3044) <= a and b;
    outputs(3045) <= not (a xor b);
    outputs(3046) <= not b;
    outputs(3047) <= not a;
    outputs(3048) <= not b;
    outputs(3049) <= a;
    outputs(3050) <= not b;
    outputs(3051) <= not b;
    outputs(3052) <= not b;
    outputs(3053) <= not (a xor b);
    outputs(3054) <= not (a xor b);
    outputs(3055) <= not (a and b);
    outputs(3056) <= not b;
    outputs(3057) <= b;
    outputs(3058) <= not a or b;
    outputs(3059) <= not b;
    outputs(3060) <= a or b;
    outputs(3061) <= b;
    outputs(3062) <= not a;
    outputs(3063) <= not (a and b);
    outputs(3064) <= not a;
    outputs(3065) <= a and not b;
    outputs(3066) <= a xor b;
    outputs(3067) <= a and b;
    outputs(3068) <= b and not a;
    outputs(3069) <= not (a xor b);
    outputs(3070) <= b;
    outputs(3071) <= not a;
    outputs(3072) <= not b or a;
    outputs(3073) <= not (a or b);
    outputs(3074) <= not (a xor b);
    outputs(3075) <= not a;
    outputs(3076) <= a and not b;
    outputs(3077) <= b;
    outputs(3078) <= not (a and b);
    outputs(3079) <= a xor b;
    outputs(3080) <= b and not a;
    outputs(3081) <= not (a or b);
    outputs(3082) <= not a;
    outputs(3083) <= a;
    outputs(3084) <= not a;
    outputs(3085) <= a;
    outputs(3086) <= b and not a;
    outputs(3087) <= a;
    outputs(3088) <= a and not b;
    outputs(3089) <= a or b;
    outputs(3090) <= b;
    outputs(3091) <= a xor b;
    outputs(3092) <= not (a or b);
    outputs(3093) <= a xor b;
    outputs(3094) <= b and not a;
    outputs(3095) <= b;
    outputs(3096) <= not (a xor b);
    outputs(3097) <= not (a xor b);
    outputs(3098) <= a;
    outputs(3099) <= not a or b;
    outputs(3100) <= not b or a;
    outputs(3101) <= not a or b;
    outputs(3102) <= not (a xor b);
    outputs(3103) <= not a or b;
    outputs(3104) <= a xor b;
    outputs(3105) <= not b;
    outputs(3106) <= not (a xor b);
    outputs(3107) <= not b;
    outputs(3108) <= not b;
    outputs(3109) <= a xor b;
    outputs(3110) <= a and not b;
    outputs(3111) <= not b;
    outputs(3112) <= not a;
    outputs(3113) <= a and b;
    outputs(3114) <= not b or a;
    outputs(3115) <= a xor b;
    outputs(3116) <= not (a and b);
    outputs(3117) <= not a;
    outputs(3118) <= a and b;
    outputs(3119) <= a xor b;
    outputs(3120) <= not (a and b);
    outputs(3121) <= not (a xor b);
    outputs(3122) <= not (a xor b);
    outputs(3123) <= b;
    outputs(3124) <= b;
    outputs(3125) <= b;
    outputs(3126) <= a;
    outputs(3127) <= b and not a;
    outputs(3128) <= not b or a;
    outputs(3129) <= a;
    outputs(3130) <= b and not a;
    outputs(3131) <= not (a xor b);
    outputs(3132) <= b;
    outputs(3133) <= a xor b;
    outputs(3134) <= not a;
    outputs(3135) <= a or b;
    outputs(3136) <= not (a or b);
    outputs(3137) <= a xor b;
    outputs(3138) <= not b;
    outputs(3139) <= not b;
    outputs(3140) <= b;
    outputs(3141) <= not (a xor b);
    outputs(3142) <= not b;
    outputs(3143) <= not a;
    outputs(3144) <= not (a xor b);
    outputs(3145) <= not b or a;
    outputs(3146) <= b;
    outputs(3147) <= not a or b;
    outputs(3148) <= not (a and b);
    outputs(3149) <= a;
    outputs(3150) <= b;
    outputs(3151) <= not (a xor b);
    outputs(3152) <= not a;
    outputs(3153) <= not (a xor b);
    outputs(3154) <= not (a and b);
    outputs(3155) <= not a;
    outputs(3156) <= b;
    outputs(3157) <= not b;
    outputs(3158) <= not b;
    outputs(3159) <= a xor b;
    outputs(3160) <= not b;
    outputs(3161) <= a xor b;
    outputs(3162) <= not b or a;
    outputs(3163) <= a or b;
    outputs(3164) <= not b or a;
    outputs(3165) <= a or b;
    outputs(3166) <= b;
    outputs(3167) <= not a;
    outputs(3168) <= b and not a;
    outputs(3169) <= b and not a;
    outputs(3170) <= a or b;
    outputs(3171) <= a and not b;
    outputs(3172) <= not b or a;
    outputs(3173) <= not b or a;
    outputs(3174) <= a xor b;
    outputs(3175) <= not b;
    outputs(3176) <= a and not b;
    outputs(3177) <= not (a and b);
    outputs(3178) <= not (a xor b);
    outputs(3179) <= not a;
    outputs(3180) <= a or b;
    outputs(3181) <= a or b;
    outputs(3182) <= not b;
    outputs(3183) <= not (a xor b);
    outputs(3184) <= a or b;
    outputs(3185) <= not b;
    outputs(3186) <= a xor b;
    outputs(3187) <= a or b;
    outputs(3188) <= a and b;
    outputs(3189) <= a;
    outputs(3190) <= a;
    outputs(3191) <= a;
    outputs(3192) <= not a;
    outputs(3193) <= a xor b;
    outputs(3194) <= b;
    outputs(3195) <= not b;
    outputs(3196) <= b;
    outputs(3197) <= not (a and b);
    outputs(3198) <= a and not b;
    outputs(3199) <= not (a xor b);
    outputs(3200) <= a;
    outputs(3201) <= not b;
    outputs(3202) <= b and not a;
    outputs(3203) <= not (a xor b);
    outputs(3204) <= a and not b;
    outputs(3205) <= not a;
    outputs(3206) <= a xor b;
    outputs(3207) <= not (a or b);
    outputs(3208) <= b and not a;
    outputs(3209) <= not a;
    outputs(3210) <= not a;
    outputs(3211) <= not (a xor b);
    outputs(3212) <= a;
    outputs(3213) <= a xor b;
    outputs(3214) <= a xor b;
    outputs(3215) <= not b;
    outputs(3216) <= a xor b;
    outputs(3217) <= a;
    outputs(3218) <= b;
    outputs(3219) <= not b;
    outputs(3220) <= b;
    outputs(3221) <= a and b;
    outputs(3222) <= not b or a;
    outputs(3223) <= not a;
    outputs(3224) <= not a;
    outputs(3225) <= not (a or b);
    outputs(3226) <= not (a xor b);
    outputs(3227) <= not b;
    outputs(3228) <= not b or a;
    outputs(3229) <= not (a xor b);
    outputs(3230) <= not (a and b);
    outputs(3231) <= not a or b;
    outputs(3232) <= a;
    outputs(3233) <= not b;
    outputs(3234) <= a xor b;
    outputs(3235) <= not b;
    outputs(3236) <= not b;
    outputs(3237) <= a and not b;
    outputs(3238) <= a and b;
    outputs(3239) <= a and not b;
    outputs(3240) <= not b;
    outputs(3241) <= a;
    outputs(3242) <= a and b;
    outputs(3243) <= not b;
    outputs(3244) <= not a;
    outputs(3245) <= b;
    outputs(3246) <= b and not a;
    outputs(3247) <= a;
    outputs(3248) <= not a or b;
    outputs(3249) <= not (a and b);
    outputs(3250) <= not b or a;
    outputs(3251) <= a xor b;
    outputs(3252) <= not a;
    outputs(3253) <= b;
    outputs(3254) <= not a;
    outputs(3255) <= a;
    outputs(3256) <= a;
    outputs(3257) <= b;
    outputs(3258) <= not a or b;
    outputs(3259) <= not (a or b);
    outputs(3260) <= a xor b;
    outputs(3261) <= not (a xor b);
    outputs(3262) <= a and b;
    outputs(3263) <= not b or a;
    outputs(3264) <= not (a xor b);
    outputs(3265) <= a;
    outputs(3266) <= not (a or b);
    outputs(3267) <= not a;
    outputs(3268) <= b;
    outputs(3269) <= not a or b;
    outputs(3270) <= a and b;
    outputs(3271) <= not (a xor b);
    outputs(3272) <= not (a and b);
    outputs(3273) <= not (a xor b);
    outputs(3274) <= not (a and b);
    outputs(3275) <= not (a and b);
    outputs(3276) <= not (a and b);
    outputs(3277) <= a and b;
    outputs(3278) <= not (a xor b);
    outputs(3279) <= b;
    outputs(3280) <= not a;
    outputs(3281) <= b and not a;
    outputs(3282) <= not (a xor b);
    outputs(3283) <= a and b;
    outputs(3284) <= not b;
    outputs(3285) <= not b;
    outputs(3286) <= not b;
    outputs(3287) <= not a or b;
    outputs(3288) <= a and not b;
    outputs(3289) <= a;
    outputs(3290) <= a;
    outputs(3291) <= not a;
    outputs(3292) <= a xor b;
    outputs(3293) <= not a;
    outputs(3294) <= not b or a;
    outputs(3295) <= not a;
    outputs(3296) <= a and b;
    outputs(3297) <= a;
    outputs(3298) <= not (a and b);
    outputs(3299) <= a xor b;
    outputs(3300) <= not (a or b);
    outputs(3301) <= not a;
    outputs(3302) <= a and not b;
    outputs(3303) <= a;
    outputs(3304) <= b;
    outputs(3305) <= not (a and b);
    outputs(3306) <= not (a and b);
    outputs(3307) <= a;
    outputs(3308) <= not a;
    outputs(3309) <= not a;
    outputs(3310) <= not a;
    outputs(3311) <= b;
    outputs(3312) <= a or b;
    outputs(3313) <= a and not b;
    outputs(3314) <= b and not a;
    outputs(3315) <= a and b;
    outputs(3316) <= not a;
    outputs(3317) <= b;
    outputs(3318) <= b and not a;
    outputs(3319) <= a;
    outputs(3320) <= not b;
    outputs(3321) <= a or b;
    outputs(3322) <= not b or a;
    outputs(3323) <= not (a and b);
    outputs(3324) <= not a;
    outputs(3325) <= a;
    outputs(3326) <= not (a xor b);
    outputs(3327) <= b;
    outputs(3328) <= not (a and b);
    outputs(3329) <= not (a and b);
    outputs(3330) <= b;
    outputs(3331) <= a or b;
    outputs(3332) <= not (a xor b);
    outputs(3333) <= not b or a;
    outputs(3334) <= not b or a;
    outputs(3335) <= not b;
    outputs(3336) <= not b;
    outputs(3337) <= a;
    outputs(3338) <= a and not b;
    outputs(3339) <= a xor b;
    outputs(3340) <= a xor b;
    outputs(3341) <= not b or a;
    outputs(3342) <= not (a xor b);
    outputs(3343) <= not b;
    outputs(3344) <= not (a xor b);
    outputs(3345) <= not a or b;
    outputs(3346) <= not a;
    outputs(3347) <= a xor b;
    outputs(3348) <= a xor b;
    outputs(3349) <= a or b;
    outputs(3350) <= not b or a;
    outputs(3351) <= not (a xor b);
    outputs(3352) <= b;
    outputs(3353) <= a xor b;
    outputs(3354) <= not a;
    outputs(3355) <= not b;
    outputs(3356) <= not a;
    outputs(3357) <= a;
    outputs(3358) <= a xor b;
    outputs(3359) <= not b;
    outputs(3360) <= not b;
    outputs(3361) <= not (a or b);
    outputs(3362) <= a;
    outputs(3363) <= not (a and b);
    outputs(3364) <= not (a xor b);
    outputs(3365) <= a xor b;
    outputs(3366) <= not (a xor b);
    outputs(3367) <= not b;
    outputs(3368) <= not a or b;
    outputs(3369) <= b;
    outputs(3370) <= not a;
    outputs(3371) <= not (a xor b);
    outputs(3372) <= a and b;
    outputs(3373) <= not (a xor b);
    outputs(3374) <= a and not b;
    outputs(3375) <= a;
    outputs(3376) <= a and b;
    outputs(3377) <= not (a or b);
    outputs(3378) <= not (a xor b);
    outputs(3379) <= b;
    outputs(3380) <= not (a and b);
    outputs(3381) <= a xor b;
    outputs(3382) <= a xor b;
    outputs(3383) <= a xor b;
    outputs(3384) <= a;
    outputs(3385) <= a;
    outputs(3386) <= a and b;
    outputs(3387) <= a and not b;
    outputs(3388) <= not a;
    outputs(3389) <= not b or a;
    outputs(3390) <= not b;
    outputs(3391) <= a;
    outputs(3392) <= b;
    outputs(3393) <= a and not b;
    outputs(3394) <= not (a xor b);
    outputs(3395) <= not (a or b);
    outputs(3396) <= not a;
    outputs(3397) <= not b or a;
    outputs(3398) <= not (a xor b);
    outputs(3399) <= a;
    outputs(3400) <= not (a xor b);
    outputs(3401) <= not a;
    outputs(3402) <= not a;
    outputs(3403) <= a and b;
    outputs(3404) <= a;
    outputs(3405) <= not b or a;
    outputs(3406) <= not (a xor b);
    outputs(3407) <= a xor b;
    outputs(3408) <= a or b;
    outputs(3409) <= not a;
    outputs(3410) <= b;
    outputs(3411) <= a and b;
    outputs(3412) <= a xor b;
    outputs(3413) <= not (a xor b);
    outputs(3414) <= b;
    outputs(3415) <= a or b;
    outputs(3416) <= a;
    outputs(3417) <= b and not a;
    outputs(3418) <= not a;
    outputs(3419) <= b and not a;
    outputs(3420) <= a and b;
    outputs(3421) <= not (a or b);
    outputs(3422) <= a xor b;
    outputs(3423) <= not b or a;
    outputs(3424) <= not (a and b);
    outputs(3425) <= not b;
    outputs(3426) <= a xor b;
    outputs(3427) <= a or b;
    outputs(3428) <= b;
    outputs(3429) <= not a;
    outputs(3430) <= not (a xor b);
    outputs(3431) <= a xor b;
    outputs(3432) <= not a or b;
    outputs(3433) <= not a;
    outputs(3434) <= b;
    outputs(3435) <= not a;
    outputs(3436) <= a or b;
    outputs(3437) <= a xor b;
    outputs(3438) <= not a;
    outputs(3439) <= not (a xor b);
    outputs(3440) <= a;
    outputs(3441) <= a and b;
    outputs(3442) <= not a or b;
    outputs(3443) <= a;
    outputs(3444) <= a;
    outputs(3445) <= a xor b;
    outputs(3446) <= a xor b;
    outputs(3447) <= not (a xor b);
    outputs(3448) <= a xor b;
    outputs(3449) <= a;
    outputs(3450) <= not a;
    outputs(3451) <= a xor b;
    outputs(3452) <= not (a and b);
    outputs(3453) <= not (a xor b);
    outputs(3454) <= a xor b;
    outputs(3455) <= not b or a;
    outputs(3456) <= a xor b;
    outputs(3457) <= a xor b;
    outputs(3458) <= not b;
    outputs(3459) <= not a or b;
    outputs(3460) <= b;
    outputs(3461) <= a;
    outputs(3462) <= not (a xor b);
    outputs(3463) <= not (a or b);
    outputs(3464) <= not b or a;
    outputs(3465) <= a and b;
    outputs(3466) <= not (a xor b);
    outputs(3467) <= b;
    outputs(3468) <= b;
    outputs(3469) <= not a;
    outputs(3470) <= a xor b;
    outputs(3471) <= not a;
    outputs(3472) <= b and not a;
    outputs(3473) <= a xor b;
    outputs(3474) <= not (a xor b);
    outputs(3475) <= a;
    outputs(3476) <= not a;
    outputs(3477) <= not a or b;
    outputs(3478) <= a xor b;
    outputs(3479) <= not b;
    outputs(3480) <= not (a xor b);
    outputs(3481) <= a and b;
    outputs(3482) <= a;
    outputs(3483) <= a;
    outputs(3484) <= b and not a;
    outputs(3485) <= not a or b;
    outputs(3486) <= not b;
    outputs(3487) <= a;
    outputs(3488) <= not (a xor b);
    outputs(3489) <= not (a xor b);
    outputs(3490) <= a;
    outputs(3491) <= b and not a;
    outputs(3492) <= not b or a;
    outputs(3493) <= not a or b;
    outputs(3494) <= a or b;
    outputs(3495) <= not (a xor b);
    outputs(3496) <= b;
    outputs(3497) <= a xor b;
    outputs(3498) <= not b;
    outputs(3499) <= not (a xor b);
    outputs(3500) <= not (a and b);
    outputs(3501) <= a xor b;
    outputs(3502) <= a and not b;
    outputs(3503) <= not b;
    outputs(3504) <= a and not b;
    outputs(3505) <= not a or b;
    outputs(3506) <= not (a xor b);
    outputs(3507) <= not (a and b);
    outputs(3508) <= a or b;
    outputs(3509) <= a and b;
    outputs(3510) <= not b;
    outputs(3511) <= a xor b;
    outputs(3512) <= not a or b;
    outputs(3513) <= a;
    outputs(3514) <= not b or a;
    outputs(3515) <= a or b;
    outputs(3516) <= not a;
    outputs(3517) <= not a or b;
    outputs(3518) <= a and not b;
    outputs(3519) <= not b or a;
    outputs(3520) <= b;
    outputs(3521) <= not (a xor b);
    outputs(3522) <= not (a and b);
    outputs(3523) <= a xor b;
    outputs(3524) <= a xor b;
    outputs(3525) <= a;
    outputs(3526) <= b and not a;
    outputs(3527) <= not a;
    outputs(3528) <= not b or a;
    outputs(3529) <= not b;
    outputs(3530) <= b;
    outputs(3531) <= a;
    outputs(3532) <= not a;
    outputs(3533) <= not (a or b);
    outputs(3534) <= not a;
    outputs(3535) <= not b or a;
    outputs(3536) <= a and b;
    outputs(3537) <= not a;
    outputs(3538) <= not a;
    outputs(3539) <= not b;
    outputs(3540) <= not b;
    outputs(3541) <= not (a xor b);
    outputs(3542) <= b and not a;
    outputs(3543) <= not b or a;
    outputs(3544) <= a xor b;
    outputs(3545) <= a;
    outputs(3546) <= a;
    outputs(3547) <= not (a or b);
    outputs(3548) <= not a or b;
    outputs(3549) <= not (a xor b);
    outputs(3550) <= not b or a;
    outputs(3551) <= a;
    outputs(3552) <= not a;
    outputs(3553) <= not (a xor b);
    outputs(3554) <= a xor b;
    outputs(3555) <= not a;
    outputs(3556) <= not a;
    outputs(3557) <= not (a and b);
    outputs(3558) <= b and not a;
    outputs(3559) <= not a;
    outputs(3560) <= not a or b;
    outputs(3561) <= a or b;
    outputs(3562) <= a xor b;
    outputs(3563) <= not a or b;
    outputs(3564) <= not (a and b);
    outputs(3565) <= not b or a;
    outputs(3566) <= a and b;
    outputs(3567) <= not (a and b);
    outputs(3568) <= not a or b;
    outputs(3569) <= b;
    outputs(3570) <= a and b;
    outputs(3571) <= not (a xor b);
    outputs(3572) <= not a or b;
    outputs(3573) <= not (a and b);
    outputs(3574) <= a or b;
    outputs(3575) <= a;
    outputs(3576) <= a or b;
    outputs(3577) <= not b;
    outputs(3578) <= not b;
    outputs(3579) <= a xor b;
    outputs(3580) <= a and b;
    outputs(3581) <= not b;
    outputs(3582) <= not a;
    outputs(3583) <= not (a or b);
    outputs(3584) <= not (a xor b);
    outputs(3585) <= not a;
    outputs(3586) <= a xor b;
    outputs(3587) <= a;
    outputs(3588) <= b and not a;
    outputs(3589) <= b;
    outputs(3590) <= not (a and b);
    outputs(3591) <= not b or a;
    outputs(3592) <= not (a xor b);
    outputs(3593) <= b;
    outputs(3594) <= not (a xor b);
    outputs(3595) <= a and b;
    outputs(3596) <= not (a or b);
    outputs(3597) <= a and not b;
    outputs(3598) <= not (a xor b);
    outputs(3599) <= not b;
    outputs(3600) <= a;
    outputs(3601) <= a and not b;
    outputs(3602) <= not (a or b);
    outputs(3603) <= a;
    outputs(3604) <= b;
    outputs(3605) <= a;
    outputs(3606) <= a;
    outputs(3607) <= not a;
    outputs(3608) <= a;
    outputs(3609) <= not a or b;
    outputs(3610) <= a xor b;
    outputs(3611) <= not (a and b);
    outputs(3612) <= not a;
    outputs(3613) <= not (a xor b);
    outputs(3614) <= not a or b;
    outputs(3615) <= a;
    outputs(3616) <= not a;
    outputs(3617) <= a or b;
    outputs(3618) <= a;
    outputs(3619) <= not b;
    outputs(3620) <= not (a and b);
    outputs(3621) <= b and not a;
    outputs(3622) <= b;
    outputs(3623) <= b and not a;
    outputs(3624) <= a;
    outputs(3625) <= '1';
    outputs(3626) <= not (a xor b);
    outputs(3627) <= a;
    outputs(3628) <= not a;
    outputs(3629) <= a;
    outputs(3630) <= b;
    outputs(3631) <= a;
    outputs(3632) <= not (a xor b);
    outputs(3633) <= a and b;
    outputs(3634) <= a and not b;
    outputs(3635) <= not b;
    outputs(3636) <= not b;
    outputs(3637) <= a xor b;
    outputs(3638) <= not (a and b);
    outputs(3639) <= b and not a;
    outputs(3640) <= a xor b;
    outputs(3641) <= not (a xor b);
    outputs(3642) <= not (a xor b);
    outputs(3643) <= b and not a;
    outputs(3644) <= a or b;
    outputs(3645) <= b and not a;
    outputs(3646) <= a xor b;
    outputs(3647) <= a and not b;
    outputs(3648) <= not a;
    outputs(3649) <= a xor b;
    outputs(3650) <= a and not b;
    outputs(3651) <= not b or a;
    outputs(3652) <= b;
    outputs(3653) <= a;
    outputs(3654) <= not b;
    outputs(3655) <= not b;
    outputs(3656) <= b;
    outputs(3657) <= not b or a;
    outputs(3658) <= a xor b;
    outputs(3659) <= b;
    outputs(3660) <= not a;
    outputs(3661) <= not (a xor b);
    outputs(3662) <= not (a and b);
    outputs(3663) <= not b or a;
    outputs(3664) <= b;
    outputs(3665) <= not (a xor b);
    outputs(3666) <= a and b;
    outputs(3667) <= not (a xor b);
    outputs(3668) <= not a;
    outputs(3669) <= a;
    outputs(3670) <= b and not a;
    outputs(3671) <= not b;
    outputs(3672) <= b;
    outputs(3673) <= not (a and b);
    outputs(3674) <= not a;
    outputs(3675) <= not b;
    outputs(3676) <= b;
    outputs(3677) <= not b;
    outputs(3678) <= not a;
    outputs(3679) <= not b;
    outputs(3680) <= not (a and b);
    outputs(3681) <= b;
    outputs(3682) <= not (a and b);
    outputs(3683) <= not b;
    outputs(3684) <= not (a and b);
    outputs(3685) <= a xor b;
    outputs(3686) <= b;
    outputs(3687) <= b;
    outputs(3688) <= not (a and b);
    outputs(3689) <= a or b;
    outputs(3690) <= a and b;
    outputs(3691) <= not (a xor b);
    outputs(3692) <= a or b;
    outputs(3693) <= b;
    outputs(3694) <= b;
    outputs(3695) <= a xor b;
    outputs(3696) <= not a;
    outputs(3697) <= not a;
    outputs(3698) <= b and not a;
    outputs(3699) <= not (a xor b);
    outputs(3700) <= not a;
    outputs(3701) <= not (a xor b);
    outputs(3702) <= b;
    outputs(3703) <= not (a and b);
    outputs(3704) <= not (a or b);
    outputs(3705) <= not b;
    outputs(3706) <= not b;
    outputs(3707) <= b;
    outputs(3708) <= a xor b;
    outputs(3709) <= not (a xor b);
    outputs(3710) <= b;
    outputs(3711) <= not b;
    outputs(3712) <= a and b;
    outputs(3713) <= not (a xor b);
    outputs(3714) <= not (a xor b);
    outputs(3715) <= not a;
    outputs(3716) <= a xor b;
    outputs(3717) <= not a or b;
    outputs(3718) <= a xor b;
    outputs(3719) <= a or b;
    outputs(3720) <= a or b;
    outputs(3721) <= not (a xor b);
    outputs(3722) <= a xor b;
    outputs(3723) <= not (a xor b);
    outputs(3724) <= not b;
    outputs(3725) <= not b;
    outputs(3726) <= not (a xor b);
    outputs(3727) <= not b;
    outputs(3728) <= not a or b;
    outputs(3729) <= a;
    outputs(3730) <= b;
    outputs(3731) <= a xor b;
    outputs(3732) <= not b;
    outputs(3733) <= not b or a;
    outputs(3734) <= b and not a;
    outputs(3735) <= not (a xor b);
    outputs(3736) <= a and not b;
    outputs(3737) <= not b or a;
    outputs(3738) <= a or b;
    outputs(3739) <= b and not a;
    outputs(3740) <= a or b;
    outputs(3741) <= b;
    outputs(3742) <= not b;
    outputs(3743) <= a and not b;
    outputs(3744) <= a and b;
    outputs(3745) <= b;
    outputs(3746) <= b and not a;
    outputs(3747) <= not (a and b);
    outputs(3748) <= not a;
    outputs(3749) <= not (a xor b);
    outputs(3750) <= b;
    outputs(3751) <= not b or a;
    outputs(3752) <= not b;
    outputs(3753) <= not (a xor b);
    outputs(3754) <= not (a or b);
    outputs(3755) <= a;
    outputs(3756) <= not a;
    outputs(3757) <= a;
    outputs(3758) <= a;
    outputs(3759) <= not (a xor b);
    outputs(3760) <= a and b;
    outputs(3761) <= not a;
    outputs(3762) <= a xor b;
    outputs(3763) <= not (a xor b);
    outputs(3764) <= not (a xor b);
    outputs(3765) <= not (a and b);
    outputs(3766) <= not (a xor b);
    outputs(3767) <= a;
    outputs(3768) <= a xor b;
    outputs(3769) <= not (a xor b);
    outputs(3770) <= a xor b;
    outputs(3771) <= not b or a;
    outputs(3772) <= not (a xor b);
    outputs(3773) <= b;
    outputs(3774) <= a xor b;
    outputs(3775) <= a;
    outputs(3776) <= not b;
    outputs(3777) <= a and b;
    outputs(3778) <= not (a xor b);
    outputs(3779) <= a and b;
    outputs(3780) <= b;
    outputs(3781) <= b;
    outputs(3782) <= not (a xor b);
    outputs(3783) <= not (a or b);
    outputs(3784) <= not (a and b);
    outputs(3785) <= not (a xor b);
    outputs(3786) <= b and not a;
    outputs(3787) <= a xor b;
    outputs(3788) <= not (a xor b);
    outputs(3789) <= a xor b;
    outputs(3790) <= not (a xor b);
    outputs(3791) <= not a or b;
    outputs(3792) <= a;
    outputs(3793) <= not (a and b);
    outputs(3794) <= a xor b;
    outputs(3795) <= not (a and b);
    outputs(3796) <= not (a xor b);
    outputs(3797) <= not (a xor b);
    outputs(3798) <= a;
    outputs(3799) <= not (a xor b);
    outputs(3800) <= a xor b;
    outputs(3801) <= not a or b;
    outputs(3802) <= not b;
    outputs(3803) <= a and b;
    outputs(3804) <= not b;
    outputs(3805) <= a and b;
    outputs(3806) <= not b;
    outputs(3807) <= not (a xor b);
    outputs(3808) <= not (a xor b);
    outputs(3809) <= a;
    outputs(3810) <= a and not b;
    outputs(3811) <= a;
    outputs(3812) <= a;
    outputs(3813) <= b;
    outputs(3814) <= not b;
    outputs(3815) <= a or b;
    outputs(3816) <= not a or b;
    outputs(3817) <= not (a xor b);
    outputs(3818) <= a xor b;
    outputs(3819) <= a;
    outputs(3820) <= not a;
    outputs(3821) <= b and not a;
    outputs(3822) <= a;
    outputs(3823) <= a;
    outputs(3824) <= a or b;
    outputs(3825) <= not (a and b);
    outputs(3826) <= not a;
    outputs(3827) <= a xor b;
    outputs(3828) <= a or b;
    outputs(3829) <= not (a and b);
    outputs(3830) <= not b;
    outputs(3831) <= not b;
    outputs(3832) <= not (a xor b);
    outputs(3833) <= not (a or b);
    outputs(3834) <= a and b;
    outputs(3835) <= a;
    outputs(3836) <= not (a xor b);
    outputs(3837) <= a;
    outputs(3838) <= a xor b;
    outputs(3839) <= not a or b;
    outputs(3840) <= a xor b;
    outputs(3841) <= not b;
    outputs(3842) <= not a;
    outputs(3843) <= not (a xor b);
    outputs(3844) <= not a;
    outputs(3845) <= not a;
    outputs(3846) <= a and not b;
    outputs(3847) <= not (a or b);
    outputs(3848) <= a and not b;
    outputs(3849) <= not a;
    outputs(3850) <= b;
    outputs(3851) <= not (a or b);
    outputs(3852) <= a or b;
    outputs(3853) <= a and b;
    outputs(3854) <= a and not b;
    outputs(3855) <= not a;
    outputs(3856) <= b;
    outputs(3857) <= a xor b;
    outputs(3858) <= a;
    outputs(3859) <= b;
    outputs(3860) <= not (a and b);
    outputs(3861) <= not (a xor b);
    outputs(3862) <= not (a xor b);
    outputs(3863) <= not a;
    outputs(3864) <= b;
    outputs(3865) <= not (a and b);
    outputs(3866) <= not (a and b);
    outputs(3867) <= a;
    outputs(3868) <= not b;
    outputs(3869) <= not (a xor b);
    outputs(3870) <= b;
    outputs(3871) <= a xor b;
    outputs(3872) <= not a or b;
    outputs(3873) <= a and not b;
    outputs(3874) <= not (a and b);
    outputs(3875) <= not (a xor b);
    outputs(3876) <= not a;
    outputs(3877) <= not a or b;
    outputs(3878) <= not b;
    outputs(3879) <= not a;
    outputs(3880) <= a;
    outputs(3881) <= a or b;
    outputs(3882) <= not (a xor b);
    outputs(3883) <= a;
    outputs(3884) <= a xor b;
    outputs(3885) <= a or b;
    outputs(3886) <= a and not b;
    outputs(3887) <= not (a and b);
    outputs(3888) <= not b;
    outputs(3889) <= not (a and b);
    outputs(3890) <= a xor b;
    outputs(3891) <= not a;
    outputs(3892) <= not a;
    outputs(3893) <= a xor b;
    outputs(3894) <= not b;
    outputs(3895) <= not b;
    outputs(3896) <= not b or a;
    outputs(3897) <= not b;
    outputs(3898) <= a xor b;
    outputs(3899) <= not b;
    outputs(3900) <= a and not b;
    outputs(3901) <= a xor b;
    outputs(3902) <= a or b;
    outputs(3903) <= a and b;
    outputs(3904) <= not a or b;
    outputs(3905) <= a xor b;
    outputs(3906) <= a and b;
    outputs(3907) <= a;
    outputs(3908) <= a and not b;
    outputs(3909) <= not (a xor b);
    outputs(3910) <= b and not a;
    outputs(3911) <= a and b;
    outputs(3912) <= a xor b;
    outputs(3913) <= not b;
    outputs(3914) <= a;
    outputs(3915) <= not (a xor b);
    outputs(3916) <= not a;
    outputs(3917) <= not a;
    outputs(3918) <= a and not b;
    outputs(3919) <= not a;
    outputs(3920) <= not b;
    outputs(3921) <= a xor b;
    outputs(3922) <= a xor b;
    outputs(3923) <= a;
    outputs(3924) <= not (a or b);
    outputs(3925) <= not (a or b);
    outputs(3926) <= not b;
    outputs(3927) <= a or b;
    outputs(3928) <= not b;
    outputs(3929) <= a xor b;
    outputs(3930) <= not a;
    outputs(3931) <= a and b;
    outputs(3932) <= a and b;
    outputs(3933) <= not a or b;
    outputs(3934) <= b;
    outputs(3935) <= a and b;
    outputs(3936) <= a and not b;
    outputs(3937) <= a and not b;
    outputs(3938) <= a;
    outputs(3939) <= a;
    outputs(3940) <= b;
    outputs(3941) <= not (a xor b);
    outputs(3942) <= a;
    outputs(3943) <= b;
    outputs(3944) <= a;
    outputs(3945) <= a or b;
    outputs(3946) <= b;
    outputs(3947) <= a or b;
    outputs(3948) <= not (a xor b);
    outputs(3949) <= b;
    outputs(3950) <= not (a or b);
    outputs(3951) <= not b;
    outputs(3952) <= a and not b;
    outputs(3953) <= not (a or b);
    outputs(3954) <= not (a or b);
    outputs(3955) <= not b;
    outputs(3956) <= a xor b;
    outputs(3957) <= not (a or b);
    outputs(3958) <= not b or a;
    outputs(3959) <= a;
    outputs(3960) <= a or b;
    outputs(3961) <= not a;
    outputs(3962) <= not b;
    outputs(3963) <= a;
    outputs(3964) <= a and b;
    outputs(3965) <= b;
    outputs(3966) <= not b;
    outputs(3967) <= not b;
    outputs(3968) <= a xor b;
    outputs(3969) <= not b or a;
    outputs(3970) <= not b;
    outputs(3971) <= b;
    outputs(3972) <= not b or a;
    outputs(3973) <= not (a and b);
    outputs(3974) <= a;
    outputs(3975) <= not (a or b);
    outputs(3976) <= a;
    outputs(3977) <= a xor b;
    outputs(3978) <= not b or a;
    outputs(3979) <= not b;
    outputs(3980) <= not (a xor b);
    outputs(3981) <= b;
    outputs(3982) <= a or b;
    outputs(3983) <= b;
    outputs(3984) <= a;
    outputs(3985) <= not (a and b);
    outputs(3986) <= b;
    outputs(3987) <= not (a xor b);
    outputs(3988) <= a;
    outputs(3989) <= not b;
    outputs(3990) <= a xor b;
    outputs(3991) <= a;
    outputs(3992) <= not (a xor b);
    outputs(3993) <= a xor b;
    outputs(3994) <= not (a or b);
    outputs(3995) <= not a;
    outputs(3996) <= a or b;
    outputs(3997) <= not (a and b);
    outputs(3998) <= not (a xor b);
    outputs(3999) <= not (a and b);
    outputs(4000) <= a xor b;
    outputs(4001) <= a and b;
    outputs(4002) <= a;
    outputs(4003) <= a xor b;
    outputs(4004) <= a and b;
    outputs(4005) <= not (a xor b);
    outputs(4006) <= not a;
    outputs(4007) <= not b or a;
    outputs(4008) <= not a;
    outputs(4009) <= a;
    outputs(4010) <= a and b;
    outputs(4011) <= a xor b;
    outputs(4012) <= b;
    outputs(4013) <= not (a xor b);
    outputs(4014) <= a and not b;
    outputs(4015) <= not (a xor b);
    outputs(4016) <= b and not a;
    outputs(4017) <= not a;
    outputs(4018) <= not a;
    outputs(4019) <= not b;
    outputs(4020) <= not a or b;
    outputs(4021) <= a xor b;
    outputs(4022) <= a and b;
    outputs(4023) <= a xor b;
    outputs(4024) <= not a or b;
    outputs(4025) <= a or b;
    outputs(4026) <= not a;
    outputs(4027) <= not (a and b);
    outputs(4028) <= not b;
    outputs(4029) <= not (a xor b);
    outputs(4030) <= not (a xor b);
    outputs(4031) <= not a or b;
    outputs(4032) <= a;
    outputs(4033) <= not b;
    outputs(4034) <= not (a or b);
    outputs(4035) <= not (a xor b);
    outputs(4036) <= a and b;
    outputs(4037) <= not (a or b);
    outputs(4038) <= not a;
    outputs(4039) <= not a;
    outputs(4040) <= a xor b;
    outputs(4041) <= not a or b;
    outputs(4042) <= not b;
    outputs(4043) <= not (a or b);
    outputs(4044) <= b;
    outputs(4045) <= not (a xor b);
    outputs(4046) <= b;
    outputs(4047) <= a and not b;
    outputs(4048) <= a and b;
    outputs(4049) <= not (a and b);
    outputs(4050) <= a and not b;
    outputs(4051) <= not (a xor b);
    outputs(4052) <= not (a xor b);
    outputs(4053) <= b;
    outputs(4054) <= a xor b;
    outputs(4055) <= not (a and b);
    outputs(4056) <= not a;
    outputs(4057) <= b and not a;
    outputs(4058) <= a;
    outputs(4059) <= not b;
    outputs(4060) <= not (a xor b);
    outputs(4061) <= a xor b;
    outputs(4062) <= b and not a;
    outputs(4063) <= not (a or b);
    outputs(4064) <= not a;
    outputs(4065) <= a;
    outputs(4066) <= a and not b;
    outputs(4067) <= a xor b;
    outputs(4068) <= a xor b;
    outputs(4069) <= a xor b;
    outputs(4070) <= not b;
    outputs(4071) <= b;
    outputs(4072) <= a and b;
    outputs(4073) <= b;
    outputs(4074) <= not (a and b);
    outputs(4075) <= not b or a;
    outputs(4076) <= a or b;
    outputs(4077) <= a xor b;
    outputs(4078) <= a xor b;
    outputs(4079) <= a and b;
    outputs(4080) <= a;
    outputs(4081) <= not b;
    outputs(4082) <= not a;
    outputs(4083) <= a xor b;
    outputs(4084) <= not a or b;
    outputs(4085) <= not b;
    outputs(4086) <= a xor b;
    outputs(4087) <= a and not b;
    outputs(4088) <= not a or b;
    outputs(4089) <= not (a and b);
    outputs(4090) <= not a;
    outputs(4091) <= not b;
    outputs(4092) <= a xor b;
    outputs(4093) <= a;
    outputs(4094) <= not (a xor b);
    outputs(4095) <= a xor b;
    outputs(4096) <= a and not b;
    outputs(4097) <= not b;
    outputs(4098) <= a and b;
    outputs(4099) <= a and b;
    outputs(4100) <= b and not a;
    outputs(4101) <= not (a or b);
    outputs(4102) <= b;
    outputs(4103) <= b and not a;
    outputs(4104) <= not (a xor b);
    outputs(4105) <= not (a xor b);
    outputs(4106) <= a;
    outputs(4107) <= not a;
    outputs(4108) <= a;
    outputs(4109) <= b;
    outputs(4110) <= not (a xor b);
    outputs(4111) <= a and b;
    outputs(4112) <= a and not b;
    outputs(4113) <= not a or b;
    outputs(4114) <= not b;
    outputs(4115) <= b;
    outputs(4116) <= not b;
    outputs(4117) <= a and not b;
    outputs(4118) <= b;
    outputs(4119) <= a xor b;
    outputs(4120) <= not a;
    outputs(4121) <= a and not b;
    outputs(4122) <= not a;
    outputs(4123) <= a;
    outputs(4124) <= not (a and b);
    outputs(4125) <= a and b;
    outputs(4126) <= not a;
    outputs(4127) <= b;
    outputs(4128) <= not (a xor b);
    outputs(4129) <= b and not a;
    outputs(4130) <= not (a xor b);
    outputs(4131) <= b and not a;
    outputs(4132) <= a xor b;
    outputs(4133) <= a xor b;
    outputs(4134) <= b;
    outputs(4135) <= not (a or b);
    outputs(4136) <= not b;
    outputs(4137) <= a and b;
    outputs(4138) <= not (a xor b);
    outputs(4139) <= a and not b;
    outputs(4140) <= not a;
    outputs(4141) <= a and b;
    outputs(4142) <= not a;
    outputs(4143) <= b;
    outputs(4144) <= a xor b;
    outputs(4145) <= not b;
    outputs(4146) <= a and b;
    outputs(4147) <= a and b;
    outputs(4148) <= not a;
    outputs(4149) <= b;
    outputs(4150) <= a;
    outputs(4151) <= b;
    outputs(4152) <= a or b;
    outputs(4153) <= a and b;
    outputs(4154) <= a xor b;
    outputs(4155) <= not (a and b);
    outputs(4156) <= not (a or b);
    outputs(4157) <= not (a or b);
    outputs(4158) <= a and not b;
    outputs(4159) <= not (a xor b);
    outputs(4160) <= b;
    outputs(4161) <= a xor b;
    outputs(4162) <= not b;
    outputs(4163) <= a;
    outputs(4164) <= not (a xor b);
    outputs(4165) <= b and not a;
    outputs(4166) <= not b;
    outputs(4167) <= not b;
    outputs(4168) <= not (a xor b);
    outputs(4169) <= a xor b;
    outputs(4170) <= a and not b;
    outputs(4171) <= a;
    outputs(4172) <= not b;
    outputs(4173) <= a and b;
    outputs(4174) <= b and not a;
    outputs(4175) <= a;
    outputs(4176) <= not (a and b);
    outputs(4177) <= a or b;
    outputs(4178) <= not a or b;
    outputs(4179) <= not a;
    outputs(4180) <= not (a xor b);
    outputs(4181) <= b and not a;
    outputs(4182) <= b and not a;
    outputs(4183) <= not b;
    outputs(4184) <= not (a or b);
    outputs(4185) <= not (a xor b);
    outputs(4186) <= not (a or b);
    outputs(4187) <= b;
    outputs(4188) <= a and b;
    outputs(4189) <= a;
    outputs(4190) <= not (a xor b);
    outputs(4191) <= not b;
    outputs(4192) <= not (a xor b);
    outputs(4193) <= b;
    outputs(4194) <= a xor b;
    outputs(4195) <= not a;
    outputs(4196) <= b and not a;
    outputs(4197) <= a;
    outputs(4198) <= a xor b;
    outputs(4199) <= not b;
    outputs(4200) <= not (a xor b);
    outputs(4201) <= a and not b;
    outputs(4202) <= b and not a;
    outputs(4203) <= a;
    outputs(4204) <= '0';
    outputs(4205) <= not a;
    outputs(4206) <= not (a or b);
    outputs(4207) <= b;
    outputs(4208) <= a and not b;
    outputs(4209) <= not (a or b);
    outputs(4210) <= b;
    outputs(4211) <= not (a and b);
    outputs(4212) <= not (a or b);
    outputs(4213) <= b and not a;
    outputs(4214) <= not (a and b);
    outputs(4215) <= a xor b;
    outputs(4216) <= b and not a;
    outputs(4217) <= a and not b;
    outputs(4218) <= not a;
    outputs(4219) <= not (a or b);
    outputs(4220) <= not a;
    outputs(4221) <= not (a xor b);
    outputs(4222) <= a and not b;
    outputs(4223) <= a and b;
    outputs(4224) <= not (a xor b);
    outputs(4225) <= not b;
    outputs(4226) <= b and not a;
    outputs(4227) <= not a or b;
    outputs(4228) <= a and b;
    outputs(4229) <= a and b;
    outputs(4230) <= a;
    outputs(4231) <= not b;
    outputs(4232) <= not (a xor b);
    outputs(4233) <= b;
    outputs(4234) <= a and not b;
    outputs(4235) <= a or b;
    outputs(4236) <= a and b;
    outputs(4237) <= b;
    outputs(4238) <= a and not b;
    outputs(4239) <= not b or a;
    outputs(4240) <= not (a xor b);
    outputs(4241) <= a and not b;
    outputs(4242) <= a xor b;
    outputs(4243) <= a xor b;
    outputs(4244) <= b;
    outputs(4245) <= not (a or b);
    outputs(4246) <= a and not b;
    outputs(4247) <= not (a xor b);
    outputs(4248) <= not a;
    outputs(4249) <= not a;
    outputs(4250) <= not (a and b);
    outputs(4251) <= not a;
    outputs(4252) <= not b or a;
    outputs(4253) <= not b;
    outputs(4254) <= a and b;
    outputs(4255) <= not (a xor b);
    outputs(4256) <= a xor b;
    outputs(4257) <= b;
    outputs(4258) <= not (a or b);
    outputs(4259) <= b and not a;
    outputs(4260) <= b and not a;
    outputs(4261) <= not (a or b);
    outputs(4262) <= a xor b;
    outputs(4263) <= a and not b;
    outputs(4264) <= a xor b;
    outputs(4265) <= a and b;
    outputs(4266) <= a;
    outputs(4267) <= a and not b;
    outputs(4268) <= b and not a;
    outputs(4269) <= a;
    outputs(4270) <= b and not a;
    outputs(4271) <= not (a or b);
    outputs(4272) <= b;
    outputs(4273) <= not b;
    outputs(4274) <= not (a or b);
    outputs(4275) <= a and b;
    outputs(4276) <= a and b;
    outputs(4277) <= a;
    outputs(4278) <= not (a xor b);
    outputs(4279) <= not (a or b);
    outputs(4280) <= a and not b;
    outputs(4281) <= b;
    outputs(4282) <= not (a xor b);
    outputs(4283) <= not (a or b);
    outputs(4284) <= b and not a;
    outputs(4285) <= a xor b;
    outputs(4286) <= a and not b;
    outputs(4287) <= not b;
    outputs(4288) <= b;
    outputs(4289) <= not b;
    outputs(4290) <= b;
    outputs(4291) <= a and b;
    outputs(4292) <= not b;
    outputs(4293) <= a;
    outputs(4294) <= a and b;
    outputs(4295) <= not a;
    outputs(4296) <= b;
    outputs(4297) <= not a or b;
    outputs(4298) <= a and not b;
    outputs(4299) <= a and b;
    outputs(4300) <= not (a xor b);
    outputs(4301) <= not (a xor b);
    outputs(4302) <= a and b;
    outputs(4303) <= not (a xor b);
    outputs(4304) <= a and not b;
    outputs(4305) <= a;
    outputs(4306) <= not b;
    outputs(4307) <= not (a xor b);
    outputs(4308) <= a and not b;
    outputs(4309) <= not b;
    outputs(4310) <= a and not b;
    outputs(4311) <= b and not a;
    outputs(4312) <= not (a xor b);
    outputs(4313) <= not (a xor b);
    outputs(4314) <= not (a or b);
    outputs(4315) <= not (a or b);
    outputs(4316) <= not (a xor b);
    outputs(4317) <= '0';
    outputs(4318) <= not b;
    outputs(4319) <= a and b;
    outputs(4320) <= not a;
    outputs(4321) <= not (a xor b);
    outputs(4322) <= b and not a;
    outputs(4323) <= b;
    outputs(4324) <= not b;
    outputs(4325) <= not a;
    outputs(4326) <= not a;
    outputs(4327) <= not (a xor b);
    outputs(4328) <= a and not b;
    outputs(4329) <= not a;
    outputs(4330) <= a xor b;
    outputs(4331) <= b;
    outputs(4332) <= not b;
    outputs(4333) <= a and b;
    outputs(4334) <= not a;
    outputs(4335) <= a;
    outputs(4336) <= a xor b;
    outputs(4337) <= not (a xor b);
    outputs(4338) <= not (a xor b);
    outputs(4339) <= b;
    outputs(4340) <= not b;
    outputs(4341) <= not (a or b);
    outputs(4342) <= a and not b;
    outputs(4343) <= b;
    outputs(4344) <= not (a or b);
    outputs(4345) <= b and not a;
    outputs(4346) <= a and b;
    outputs(4347) <= not b;
    outputs(4348) <= not a;
    outputs(4349) <= a and not b;
    outputs(4350) <= not b or a;
    outputs(4351) <= not (a xor b);
    outputs(4352) <= a and b;
    outputs(4353) <= not b;
    outputs(4354) <= b and not a;
    outputs(4355) <= not a;
    outputs(4356) <= b and not a;
    outputs(4357) <= a and not b;
    outputs(4358) <= b and not a;
    outputs(4359) <= not (a xor b);
    outputs(4360) <= not (a xor b);
    outputs(4361) <= not (a or b);
    outputs(4362) <= a;
    outputs(4363) <= a and b;
    outputs(4364) <= not b;
    outputs(4365) <= not (a xor b);
    outputs(4366) <= a;
    outputs(4367) <= a;
    outputs(4368) <= not a;
    outputs(4369) <= not (a xor b);
    outputs(4370) <= a and b;
    outputs(4371) <= b;
    outputs(4372) <= a;
    outputs(4373) <= b;
    outputs(4374) <= a or b;
    outputs(4375) <= b;
    outputs(4376) <= not b or a;
    outputs(4377) <= b and not a;
    outputs(4378) <= not (a or b);
    outputs(4379) <= a;
    outputs(4380) <= a;
    outputs(4381) <= a xor b;
    outputs(4382) <= not a;
    outputs(4383) <= a and b;
    outputs(4384) <= not a;
    outputs(4385) <= a xor b;
    outputs(4386) <= a and b;
    outputs(4387) <= a xor b;
    outputs(4388) <= a and not b;
    outputs(4389) <= not b;
    outputs(4390) <= a and not b;
    outputs(4391) <= not (a xor b);
    outputs(4392) <= not a;
    outputs(4393) <= not b;
    outputs(4394) <= b and not a;
    outputs(4395) <= not (a xor b);
    outputs(4396) <= not a or b;
    outputs(4397) <= a;
    outputs(4398) <= a xor b;
    outputs(4399) <= not (a or b);
    outputs(4400) <= a and not b;
    outputs(4401) <= not (a or b);
    outputs(4402) <= not (a xor b);
    outputs(4403) <= a and b;
    outputs(4404) <= not a;
    outputs(4405) <= not (a xor b);
    outputs(4406) <= b;
    outputs(4407) <= b and not a;
    outputs(4408) <= b and not a;
    outputs(4409) <= b and not a;
    outputs(4410) <= a xor b;
    outputs(4411) <= not b;
    outputs(4412) <= b;
    outputs(4413) <= a xor b;
    outputs(4414) <= not a;
    outputs(4415) <= not a;
    outputs(4416) <= a;
    outputs(4417) <= not a;
    outputs(4418) <= a and b;
    outputs(4419) <= b and not a;
    outputs(4420) <= not (a xor b);
    outputs(4421) <= not a or b;
    outputs(4422) <= not a;
    outputs(4423) <= a;
    outputs(4424) <= a;
    outputs(4425) <= b;
    outputs(4426) <= a xor b;
    outputs(4427) <= a xor b;
    outputs(4428) <= a xor b;
    outputs(4429) <= not b;
    outputs(4430) <= not b;
    outputs(4431) <= not b;
    outputs(4432) <= not a or b;
    outputs(4433) <= b;
    outputs(4434) <= not (a or b);
    outputs(4435) <= not a;
    outputs(4436) <= not (a xor b);
    outputs(4437) <= b;
    outputs(4438) <= a;
    outputs(4439) <= a or b;
    outputs(4440) <= a and b;
    outputs(4441) <= b;
    outputs(4442) <= not (a xor b);
    outputs(4443) <= not a;
    outputs(4444) <= not b;
    outputs(4445) <= a;
    outputs(4446) <= not (a and b);
    outputs(4447) <= a xor b;
    outputs(4448) <= b and not a;
    outputs(4449) <= not b;
    outputs(4450) <= a;
    outputs(4451) <= b;
    outputs(4452) <= a xor b;
    outputs(4453) <= a and b;
    outputs(4454) <= b and not a;
    outputs(4455) <= b and not a;
    outputs(4456) <= b;
    outputs(4457) <= b and not a;
    outputs(4458) <= not (a xor b);
    outputs(4459) <= a and b;
    outputs(4460) <= not (a xor b);
    outputs(4461) <= not b;
    outputs(4462) <= not (a xor b);
    outputs(4463) <= a xor b;
    outputs(4464) <= not b;
    outputs(4465) <= a;
    outputs(4466) <= a;
    outputs(4467) <= a;
    outputs(4468) <= a and b;
    outputs(4469) <= b and not a;
    outputs(4470) <= a and not b;
    outputs(4471) <= b and not a;
    outputs(4472) <= not (a xor b);
    outputs(4473) <= not b;
    outputs(4474) <= b;
    outputs(4475) <= '0';
    outputs(4476) <= a xor b;
    outputs(4477) <= not (a xor b);
    outputs(4478) <= not b or a;
    outputs(4479) <= not (a or b);
    outputs(4480) <= not b;
    outputs(4481) <= not (a or b);
    outputs(4482) <= b;
    outputs(4483) <= not a;
    outputs(4484) <= b;
    outputs(4485) <= not b;
    outputs(4486) <= b and not a;
    outputs(4487) <= b and not a;
    outputs(4488) <= a and b;
    outputs(4489) <= b and not a;
    outputs(4490) <= a xor b;
    outputs(4491) <= b;
    outputs(4492) <= b and not a;
    outputs(4493) <= not b;
    outputs(4494) <= not (a or b);
    outputs(4495) <= a and not b;
    outputs(4496) <= b;
    outputs(4497) <= b;
    outputs(4498) <= not (a xor b);
    outputs(4499) <= b and not a;
    outputs(4500) <= not b;
    outputs(4501) <= b and not a;
    outputs(4502) <= not a;
    outputs(4503) <= a and b;
    outputs(4504) <= a and b;
    outputs(4505) <= b;
    outputs(4506) <= a and not b;
    outputs(4507) <= not a or b;
    outputs(4508) <= not b;
    outputs(4509) <= a and b;
    outputs(4510) <= a and b;
    outputs(4511) <= a xor b;
    outputs(4512) <= not (a xor b);
    outputs(4513) <= b and not a;
    outputs(4514) <= b;
    outputs(4515) <= b;
    outputs(4516) <= '0';
    outputs(4517) <= a and b;
    outputs(4518) <= not b;
    outputs(4519) <= b and not a;
    outputs(4520) <= a;
    outputs(4521) <= a xor b;
    outputs(4522) <= a and not b;
    outputs(4523) <= b;
    outputs(4524) <= a;
    outputs(4525) <= not b;
    outputs(4526) <= not b;
    outputs(4527) <= a and not b;
    outputs(4528) <= not b;
    outputs(4529) <= a;
    outputs(4530) <= b;
    outputs(4531) <= a xor b;
    outputs(4532) <= not (a xor b);
    outputs(4533) <= a;
    outputs(4534) <= not (a xor b);
    outputs(4535) <= not (a xor b);
    outputs(4536) <= a and not b;
    outputs(4537) <= not b or a;
    outputs(4538) <= not a;
    outputs(4539) <= a and not b;
    outputs(4540) <= b;
    outputs(4541) <= not a;
    outputs(4542) <= b and not a;
    outputs(4543) <= b and not a;
    outputs(4544) <= a and not b;
    outputs(4545) <= not (a xor b);
    outputs(4546) <= a and not b;
    outputs(4547) <= a and not b;
    outputs(4548) <= not (a xor b);
    outputs(4549) <= a;
    outputs(4550) <= a and b;
    outputs(4551) <= b and not a;
    outputs(4552) <= not a;
    outputs(4553) <= not (a or b);
    outputs(4554) <= not (a and b);
    outputs(4555) <= not (a xor b);
    outputs(4556) <= b;
    outputs(4557) <= a and b;
    outputs(4558) <= not a;
    outputs(4559) <= a and b;
    outputs(4560) <= not a;
    outputs(4561) <= not a;
    outputs(4562) <= a;
    outputs(4563) <= a;
    outputs(4564) <= not b;
    outputs(4565) <= a xor b;
    outputs(4566) <= not (a or b);
    outputs(4567) <= not b;
    outputs(4568) <= b;
    outputs(4569) <= not a;
    outputs(4570) <= not b;
    outputs(4571) <= a xor b;
    outputs(4572) <= a xor b;
    outputs(4573) <= a and b;
    outputs(4574) <= not a;
    outputs(4575) <= not (a or b);
    outputs(4576) <= b;
    outputs(4577) <= a;
    outputs(4578) <= a xor b;
    outputs(4579) <= a;
    outputs(4580) <= b and not a;
    outputs(4581) <= not b;
    outputs(4582) <= not a or b;
    outputs(4583) <= b and not a;
    outputs(4584) <= a and not b;
    outputs(4585) <= b and not a;
    outputs(4586) <= b;
    outputs(4587) <= a xor b;
    outputs(4588) <= not b;
    outputs(4589) <= not (a or b);
    outputs(4590) <= not (a xor b);
    outputs(4591) <= not (a and b);
    outputs(4592) <= not (a xor b);
    outputs(4593) <= b and not a;
    outputs(4594) <= not (a xor b);
    outputs(4595) <= not a;
    outputs(4596) <= a and b;
    outputs(4597) <= not (a xor b);
    outputs(4598) <= a;
    outputs(4599) <= '0';
    outputs(4600) <= a;
    outputs(4601) <= not (a or b);
    outputs(4602) <= not a;
    outputs(4603) <= a and not b;
    outputs(4604) <= a xor b;
    outputs(4605) <= a and b;
    outputs(4606) <= not (a or b);
    outputs(4607) <= a;
    outputs(4608) <= not b;
    outputs(4609) <= not (a xor b);
    outputs(4610) <= b and not a;
    outputs(4611) <= a and b;
    outputs(4612) <= not b;
    outputs(4613) <= not b or a;
    outputs(4614) <= not (a or b);
    outputs(4615) <= not (a xor b);
    outputs(4616) <= b and not a;
    outputs(4617) <= b and not a;
    outputs(4618) <= a;
    outputs(4619) <= b and not a;
    outputs(4620) <= a and b;
    outputs(4621) <= b and not a;
    outputs(4622) <= a xor b;
    outputs(4623) <= a xor b;
    outputs(4624) <= not a;
    outputs(4625) <= a and b;
    outputs(4626) <= not (a or b);
    outputs(4627) <= not (a or b);
    outputs(4628) <= b;
    outputs(4629) <= a xor b;
    outputs(4630) <= not b;
    outputs(4631) <= a and not b;
    outputs(4632) <= b;
    outputs(4633) <= not (a xor b);
    outputs(4634) <= a;
    outputs(4635) <= not b or a;
    outputs(4636) <= a or b;
    outputs(4637) <= not (a or b);
    outputs(4638) <= b and not a;
    outputs(4639) <= a and not b;
    outputs(4640) <= a and b;
    outputs(4641) <= not b or a;
    outputs(4642) <= not (a xor b);
    outputs(4643) <= not (a or b);
    outputs(4644) <= a xor b;
    outputs(4645) <= not b or a;
    outputs(4646) <= not a;
    outputs(4647) <= a and not b;
    outputs(4648) <= a and b;
    outputs(4649) <= not a;
    outputs(4650) <= a or b;
    outputs(4651) <= not a;
    outputs(4652) <= not a;
    outputs(4653) <= a and not b;
    outputs(4654) <= a and not b;
    outputs(4655) <= b;
    outputs(4656) <= not b;
    outputs(4657) <= b;
    outputs(4658) <= b and not a;
    outputs(4659) <= a and not b;
    outputs(4660) <= not a;
    outputs(4661) <= a and b;
    outputs(4662) <= b;
    outputs(4663) <= not a;
    outputs(4664) <= a;
    outputs(4665) <= a;
    outputs(4666) <= not (a or b);
    outputs(4667) <= a xor b;
    outputs(4668) <= not (a or b);
    outputs(4669) <= b;
    outputs(4670) <= a and b;
    outputs(4671) <= b;
    outputs(4672) <= a;
    outputs(4673) <= not a or b;
    outputs(4674) <= a xor b;
    outputs(4675) <= not a or b;
    outputs(4676) <= a;
    outputs(4677) <= not b;
    outputs(4678) <= a and not b;
    outputs(4679) <= not (a xor b);
    outputs(4680) <= a xor b;
    outputs(4681) <= not (a xor b);
    outputs(4682) <= b and not a;
    outputs(4683) <= not b;
    outputs(4684) <= a xor b;
    outputs(4685) <= a and b;
    outputs(4686) <= not b or a;
    outputs(4687) <= not (a or b);
    outputs(4688) <= a and b;
    outputs(4689) <= not (a xor b);
    outputs(4690) <= a or b;
    outputs(4691) <= a xor b;
    outputs(4692) <= a;
    outputs(4693) <= not a;
    outputs(4694) <= not (a and b);
    outputs(4695) <= b and not a;
    outputs(4696) <= not b;
    outputs(4697) <= not a;
    outputs(4698) <= not b;
    outputs(4699) <= b and not a;
    outputs(4700) <= b;
    outputs(4701) <= not (a xor b);
    outputs(4702) <= a and not b;
    outputs(4703) <= a and b;
    outputs(4704) <= a xor b;
    outputs(4705) <= not a or b;
    outputs(4706) <= not a;
    outputs(4707) <= a;
    outputs(4708) <= not (a or b);
    outputs(4709) <= a xor b;
    outputs(4710) <= a and not b;
    outputs(4711) <= b;
    outputs(4712) <= a xor b;
    outputs(4713) <= b and not a;
    outputs(4714) <= a;
    outputs(4715) <= not a;
    outputs(4716) <= b;
    outputs(4717) <= b;
    outputs(4718) <= not a or b;
    outputs(4719) <= not (a or b);
    outputs(4720) <= a and b;
    outputs(4721) <= not b;
    outputs(4722) <= a xor b;
    outputs(4723) <= a;
    outputs(4724) <= not (a or b);
    outputs(4725) <= a and not b;
    outputs(4726) <= a and b;
    outputs(4727) <= not (a xor b);
    outputs(4728) <= b;
    outputs(4729) <= not (a xor b);
    outputs(4730) <= b and not a;
    outputs(4731) <= not (a xor b);
    outputs(4732) <= not (a and b);
    outputs(4733) <= not (a or b);
    outputs(4734) <= a;
    outputs(4735) <= a and b;
    outputs(4736) <= a;
    outputs(4737) <= a xor b;
    outputs(4738) <= b and not a;
    outputs(4739) <= not b;
    outputs(4740) <= a and not b;
    outputs(4741) <= not a;
    outputs(4742) <= a and b;
    outputs(4743) <= a;
    outputs(4744) <= a and not b;
    outputs(4745) <= not b;
    outputs(4746) <= not a;
    outputs(4747) <= not (a xor b);
    outputs(4748) <= a xor b;
    outputs(4749) <= a and not b;
    outputs(4750) <= b and not a;
    outputs(4751) <= b;
    outputs(4752) <= not a;
    outputs(4753) <= a and b;
    outputs(4754) <= not b;
    outputs(4755) <= a xor b;
    outputs(4756) <= not b;
    outputs(4757) <= b and not a;
    outputs(4758) <= b;
    outputs(4759) <= b;
    outputs(4760) <= not b;
    outputs(4761) <= not b;
    outputs(4762) <= not (a or b);
    outputs(4763) <= b and not a;
    outputs(4764) <= a xor b;
    outputs(4765) <= '0';
    outputs(4766) <= not b;
    outputs(4767) <= a and not b;
    outputs(4768) <= not b;
    outputs(4769) <= a;
    outputs(4770) <= not (a or b);
    outputs(4771) <= a xor b;
    outputs(4772) <= not (a xor b);
    outputs(4773) <= b;
    outputs(4774) <= a and b;
    outputs(4775) <= a xor b;
    outputs(4776) <= b;
    outputs(4777) <= not (a xor b);
    outputs(4778) <= not a;
    outputs(4779) <= not (a or b);
    outputs(4780) <= a;
    outputs(4781) <= not (a xor b);
    outputs(4782) <= a and b;
    outputs(4783) <= not a;
    outputs(4784) <= b and not a;
    outputs(4785) <= not (a or b);
    outputs(4786) <= a and b;
    outputs(4787) <= a;
    outputs(4788) <= not a;
    outputs(4789) <= a xor b;
    outputs(4790) <= a and b;
    outputs(4791) <= not (a or b);
    outputs(4792) <= b and not a;
    outputs(4793) <= not (a xor b);
    outputs(4794) <= not (a or b);
    outputs(4795) <= not a;
    outputs(4796) <= a xor b;
    outputs(4797) <= not b;
    outputs(4798) <= not (a xor b);
    outputs(4799) <= a and not b;
    outputs(4800) <= a and not b;
    outputs(4801) <= not b;
    outputs(4802) <= not (a or b);
    outputs(4803) <= a xor b;
    outputs(4804) <= b and not a;
    outputs(4805) <= a;
    outputs(4806) <= not a;
    outputs(4807) <= a or b;
    outputs(4808) <= not (a xor b);
    outputs(4809) <= not a or b;
    outputs(4810) <= not (a or b);
    outputs(4811) <= not b;
    outputs(4812) <= b;
    outputs(4813) <= a and b;
    outputs(4814) <= a;
    outputs(4815) <= not (a or b);
    outputs(4816) <= not (a and b);
    outputs(4817) <= a xor b;
    outputs(4818) <= not b;
    outputs(4819) <= not (a or b);
    outputs(4820) <= a xor b;
    outputs(4821) <= not (a or b);
    outputs(4822) <= a and b;
    outputs(4823) <= b;
    outputs(4824) <= b and not a;
    outputs(4825) <= a and not b;
    outputs(4826) <= b and not a;
    outputs(4827) <= a;
    outputs(4828) <= a and not b;
    outputs(4829) <= not b;
    outputs(4830) <= not (a or b);
    outputs(4831) <= not a or b;
    outputs(4832) <= a or b;
    outputs(4833) <= not (a or b);
    outputs(4834) <= not a or b;
    outputs(4835) <= not (a and b);
    outputs(4836) <= not (a or b);
    outputs(4837) <= a;
    outputs(4838) <= not a;
    outputs(4839) <= a xor b;
    outputs(4840) <= not b;
    outputs(4841) <= not (a xor b);
    outputs(4842) <= not b;
    outputs(4843) <= b;
    outputs(4844) <= not b;
    outputs(4845) <= a xor b;
    outputs(4846) <= b and not a;
    outputs(4847) <= a xor b;
    outputs(4848) <= b;
    outputs(4849) <= not b;
    outputs(4850) <= b;
    outputs(4851) <= a and b;
    outputs(4852) <= not a;
    outputs(4853) <= a and b;
    outputs(4854) <= not b;
    outputs(4855) <= not (a xor b);
    outputs(4856) <= a xor b;
    outputs(4857) <= a xor b;
    outputs(4858) <= b and not a;
    outputs(4859) <= a and b;
    outputs(4860) <= a;
    outputs(4861) <= not b;
    outputs(4862) <= not (a or b);
    outputs(4863) <= a and not b;
    outputs(4864) <= a and not b;
    outputs(4865) <= not b;
    outputs(4866) <= b;
    outputs(4867) <= a;
    outputs(4868) <= b;
    outputs(4869) <= not a;
    outputs(4870) <= a and not b;
    outputs(4871) <= not (a or b);
    outputs(4872) <= a and not b;
    outputs(4873) <= a or b;
    outputs(4874) <= a xor b;
    outputs(4875) <= not a;
    outputs(4876) <= a and not b;
    outputs(4877) <= not (a xor b);
    outputs(4878) <= b and not a;
    outputs(4879) <= a;
    outputs(4880) <= a and not b;
    outputs(4881) <= b;
    outputs(4882) <= a;
    outputs(4883) <= b and not a;
    outputs(4884) <= not b;
    outputs(4885) <= a xor b;
    outputs(4886) <= a and b;
    outputs(4887) <= '0';
    outputs(4888) <= not b;
    outputs(4889) <= b;
    outputs(4890) <= a and not b;
    outputs(4891) <= not a;
    outputs(4892) <= not b;
    outputs(4893) <= not (a xor b);
    outputs(4894) <= b and not a;
    outputs(4895) <= not (a xor b);
    outputs(4896) <= not a;
    outputs(4897) <= a and not b;
    outputs(4898) <= a and b;
    outputs(4899) <= b and not a;
    outputs(4900) <= not (a or b);
    outputs(4901) <= b and not a;
    outputs(4902) <= b;
    outputs(4903) <= b;
    outputs(4904) <= b and not a;
    outputs(4905) <= a xor b;
    outputs(4906) <= a xor b;
    outputs(4907) <= not b;
    outputs(4908) <= a and not b;
    outputs(4909) <= not b;
    outputs(4910) <= not (a xor b);
    outputs(4911) <= not b;
    outputs(4912) <= not b or a;
    outputs(4913) <= a and not b;
    outputs(4914) <= not (a xor b);
    outputs(4915) <= a xor b;
    outputs(4916) <= '0';
    outputs(4917) <= not (a or b);
    outputs(4918) <= b;
    outputs(4919) <= not (a xor b);
    outputs(4920) <= not b or a;
    outputs(4921) <= a xor b;
    outputs(4922) <= not b;
    outputs(4923) <= b;
    outputs(4924) <= not (a xor b);
    outputs(4925) <= not b;
    outputs(4926) <= b;
    outputs(4927) <= not a;
    outputs(4928) <= a;
    outputs(4929) <= a;
    outputs(4930) <= b and not a;
    outputs(4931) <= a and b;
    outputs(4932) <= a xor b;
    outputs(4933) <= not a;
    outputs(4934) <= a;
    outputs(4935) <= a;
    outputs(4936) <= b and not a;
    outputs(4937) <= a xor b;
    outputs(4938) <= a and not b;
    outputs(4939) <= b and not a;
    outputs(4940) <= a and not b;
    outputs(4941) <= a;
    outputs(4942) <= not (a or b);
    outputs(4943) <= not b;
    outputs(4944) <= a and not b;
    outputs(4945) <= a and b;
    outputs(4946) <= not b;
    outputs(4947) <= not b;
    outputs(4948) <= a and b;
    outputs(4949) <= a;
    outputs(4950) <= a xor b;
    outputs(4951) <= a xor b;
    outputs(4952) <= a and b;
    outputs(4953) <= not b;
    outputs(4954) <= not a;
    outputs(4955) <= not (a and b);
    outputs(4956) <= not a;
    outputs(4957) <= not b;
    outputs(4958) <= not (a xor b);
    outputs(4959) <= not a;
    outputs(4960) <= a xor b;
    outputs(4961) <= a and not b;
    outputs(4962) <= not (a or b);
    outputs(4963) <= a and b;
    outputs(4964) <= a and not b;
    outputs(4965) <= a;
    outputs(4966) <= b and not a;
    outputs(4967) <= a;
    outputs(4968) <= a xor b;
    outputs(4969) <= a xor b;
    outputs(4970) <= not (a or b);
    outputs(4971) <= a xor b;
    outputs(4972) <= a xor b;
    outputs(4973) <= not (a or b);
    outputs(4974) <= not (a or b);
    outputs(4975) <= a and b;
    outputs(4976) <= a xor b;
    outputs(4977) <= not b;
    outputs(4978) <= a xor b;
    outputs(4979) <= not (a xor b);
    outputs(4980) <= a xor b;
    outputs(4981) <= a and b;
    outputs(4982) <= b and not a;
    outputs(4983) <= not (a xor b);
    outputs(4984) <= b;
    outputs(4985) <= not (a xor b);
    outputs(4986) <= b and not a;
    outputs(4987) <= a and not b;
    outputs(4988) <= not b;
    outputs(4989) <= a and not b;
    outputs(4990) <= not b;
    outputs(4991) <= not b;
    outputs(4992) <= a xor b;
    outputs(4993) <= a and b;
    outputs(4994) <= a xor b;
    outputs(4995) <= not (a xor b);
    outputs(4996) <= a or b;
    outputs(4997) <= a;
    outputs(4998) <= a and not b;
    outputs(4999) <= a and b;
    outputs(5000) <= a;
    outputs(5001) <= a;
    outputs(5002) <= a;
    outputs(5003) <= not a;
    outputs(5004) <= not (a xor b);
    outputs(5005) <= b and not a;
    outputs(5006) <= a and not b;
    outputs(5007) <= a and not b;
    outputs(5008) <= b;
    outputs(5009) <= a and b;
    outputs(5010) <= not (a or b);
    outputs(5011) <= b and not a;
    outputs(5012) <= not (a or b);
    outputs(5013) <= not b;
    outputs(5014) <= b and not a;
    outputs(5015) <= a and b;
    outputs(5016) <= a xor b;
    outputs(5017) <= not a;
    outputs(5018) <= a and not b;
    outputs(5019) <= not a;
    outputs(5020) <= a and b;
    outputs(5021) <= a xor b;
    outputs(5022) <= a xor b;
    outputs(5023) <= not b or a;
    outputs(5024) <= not b;
    outputs(5025) <= a and not b;
    outputs(5026) <= not b or a;
    outputs(5027) <= a and not b;
    outputs(5028) <= not b;
    outputs(5029) <= not a;
    outputs(5030) <= a and not b;
    outputs(5031) <= not (a or b);
    outputs(5032) <= not a;
    outputs(5033) <= a xor b;
    outputs(5034) <= a and not b;
    outputs(5035) <= a and b;
    outputs(5036) <= a and not b;
    outputs(5037) <= b;
    outputs(5038) <= a and b;
    outputs(5039) <= not (a or b);
    outputs(5040) <= not (a xor b);
    outputs(5041) <= not b or a;
    outputs(5042) <= not (a and b);
    outputs(5043) <= a;
    outputs(5044) <= b;
    outputs(5045) <= a and not b;
    outputs(5046) <= a;
    outputs(5047) <= not a;
    outputs(5048) <= not (a or b);
    outputs(5049) <= a xor b;
    outputs(5050) <= not (a or b);
    outputs(5051) <= b and not a;
    outputs(5052) <= not (a xor b);
    outputs(5053) <= b;
    outputs(5054) <= not a;
    outputs(5055) <= a xor b;
    outputs(5056) <= not b;
    outputs(5057) <= not b;
    outputs(5058) <= not (a or b);
    outputs(5059) <= b;
    outputs(5060) <= not a;
    outputs(5061) <= a xor b;
    outputs(5062) <= a and b;
    outputs(5063) <= a xor b;
    outputs(5064) <= a or b;
    outputs(5065) <= b;
    outputs(5066) <= not (a or b);
    outputs(5067) <= a;
    outputs(5068) <= a and b;
    outputs(5069) <= a and b;
    outputs(5070) <= not a;
    outputs(5071) <= not (a xor b);
    outputs(5072) <= not (a xor b);
    outputs(5073) <= not b;
    outputs(5074) <= a xor b;
    outputs(5075) <= a xor b;
    outputs(5076) <= not (a xor b);
    outputs(5077) <= not (a xor b);
    outputs(5078) <= a and not b;
    outputs(5079) <= a and b;
    outputs(5080) <= a xor b;
    outputs(5081) <= not b;
    outputs(5082) <= b;
    outputs(5083) <= not b or a;
    outputs(5084) <= a and not b;
    outputs(5085) <= not a;
    outputs(5086) <= not (a xor b);
    outputs(5087) <= not (a xor b);
    outputs(5088) <= not b;
    outputs(5089) <= not (a xor b);
    outputs(5090) <= not a;
    outputs(5091) <= not b;
    outputs(5092) <= a;
    outputs(5093) <= not b or a;
    outputs(5094) <= not (a xor b);
    outputs(5095) <= not a;
    outputs(5096) <= a and b;
    outputs(5097) <= not a;
    outputs(5098) <= not (a xor b);
    outputs(5099) <= not (a xor b);
    outputs(5100) <= a or b;
    outputs(5101) <= b and not a;
    outputs(5102) <= a and b;
    outputs(5103) <= not b or a;
    outputs(5104) <= a and b;
    outputs(5105) <= b and not a;
    outputs(5106) <= b;
    outputs(5107) <= not (a xor b);
    outputs(5108) <= b and not a;
    outputs(5109) <= not a;
    outputs(5110) <= a xor b;
    outputs(5111) <= a;
    outputs(5112) <= b and not a;
    outputs(5113) <= a and b;
    outputs(5114) <= not b;
    outputs(5115) <= not a;
    outputs(5116) <= a and not b;
    outputs(5117) <= a and b;
    outputs(5118) <= not (a xor b);
    outputs(5119) <= a and not b;
    outputs(5120) <= a or b;
    outputs(5121) <= a;
    outputs(5122) <= a xor b;
    outputs(5123) <= not b or a;
    outputs(5124) <= not b;
    outputs(5125) <= a xor b;
    outputs(5126) <= a;
    outputs(5127) <= not a;
    outputs(5128) <= not (a and b);
    outputs(5129) <= a;
    outputs(5130) <= not a;
    outputs(5131) <= not (a or b);
    outputs(5132) <= not (a xor b);
    outputs(5133) <= not b;
    outputs(5134) <= not (a and b);
    outputs(5135) <= not a or b;
    outputs(5136) <= not b;
    outputs(5137) <= not b;
    outputs(5138) <= not (a xor b);
    outputs(5139) <= b;
    outputs(5140) <= a xor b;
    outputs(5141) <= b;
    outputs(5142) <= a and b;
    outputs(5143) <= b;
    outputs(5144) <= not b or a;
    outputs(5145) <= a and not b;
    outputs(5146) <= b and not a;
    outputs(5147) <= not (a xor b);
    outputs(5148) <= a xor b;
    outputs(5149) <= a or b;
    outputs(5150) <= a xor b;
    outputs(5151) <= not (a xor b);
    outputs(5152) <= a xor b;
    outputs(5153) <= a;
    outputs(5154) <= a xor b;
    outputs(5155) <= a and not b;
    outputs(5156) <= not (a xor b);
    outputs(5157) <= b;
    outputs(5158) <= not (a xor b);
    outputs(5159) <= not (a xor b);
    outputs(5160) <= not a or b;
    outputs(5161) <= a xor b;
    outputs(5162) <= a;
    outputs(5163) <= a;
    outputs(5164) <= a or b;
    outputs(5165) <= not b or a;
    outputs(5166) <= a or b;
    outputs(5167) <= b;
    outputs(5168) <= not (a or b);
    outputs(5169) <= not b or a;
    outputs(5170) <= not a;
    outputs(5171) <= a xor b;
    outputs(5172) <= a xor b;
    outputs(5173) <= a xor b;
    outputs(5174) <= not a;
    outputs(5175) <= not (a xor b);
    outputs(5176) <= a xor b;
    outputs(5177) <= a xor b;
    outputs(5178) <= a;
    outputs(5179) <= not b;
    outputs(5180) <= not (a xor b);
    outputs(5181) <= b and not a;
    outputs(5182) <= a or b;
    outputs(5183) <= b and not a;
    outputs(5184) <= a xor b;
    outputs(5185) <= not (a xor b);
    outputs(5186) <= not b;
    outputs(5187) <= b;
    outputs(5188) <= a xor b;
    outputs(5189) <= not (a or b);
    outputs(5190) <= not (a xor b);
    outputs(5191) <= not a;
    outputs(5192) <= not a;
    outputs(5193) <= a;
    outputs(5194) <= b;
    outputs(5195) <= b;
    outputs(5196) <= not (a xor b);
    outputs(5197) <= not (a xor b);
    outputs(5198) <= not (a xor b);
    outputs(5199) <= a;
    outputs(5200) <= a;
    outputs(5201) <= a and not b;
    outputs(5202) <= a and not b;
    outputs(5203) <= b;
    outputs(5204) <= b;
    outputs(5205) <= not b;
    outputs(5206) <= a;
    outputs(5207) <= not a or b;
    outputs(5208) <= a xor b;
    outputs(5209) <= not a;
    outputs(5210) <= a xor b;
    outputs(5211) <= not (a xor b);
    outputs(5212) <= a xor b;
    outputs(5213) <= not a;
    outputs(5214) <= a xor b;
    outputs(5215) <= a;
    outputs(5216) <= a or b;
    outputs(5217) <= a or b;
    outputs(5218) <= not (a xor b);
    outputs(5219) <= b;
    outputs(5220) <= a;
    outputs(5221) <= not b;
    outputs(5222) <= b;
    outputs(5223) <= not b or a;
    outputs(5224) <= a xor b;
    outputs(5225) <= not (a xor b);
    outputs(5226) <= a;
    outputs(5227) <= a xor b;
    outputs(5228) <= not (a xor b);
    outputs(5229) <= not (a or b);
    outputs(5230) <= a;
    outputs(5231) <= not a;
    outputs(5232) <= not a;
    outputs(5233) <= a xor b;
    outputs(5234) <= a or b;
    outputs(5235) <= not (a xor b);
    outputs(5236) <= a and not b;
    outputs(5237) <= not a or b;
    outputs(5238) <= a;
    outputs(5239) <= a xor b;
    outputs(5240) <= not b;
    outputs(5241) <= not a;
    outputs(5242) <= a;
    outputs(5243) <= a;
    outputs(5244) <= not (a xor b);
    outputs(5245) <= b;
    outputs(5246) <= not (a and b);
    outputs(5247) <= not (a xor b);
    outputs(5248) <= b and not a;
    outputs(5249) <= a xor b;
    outputs(5250) <= b;
    outputs(5251) <= not b or a;
    outputs(5252) <= not a or b;
    outputs(5253) <= a and not b;
    outputs(5254) <= b;
    outputs(5255) <= not (a xor b);
    outputs(5256) <= a xor b;
    outputs(5257) <= a and not b;
    outputs(5258) <= a and b;
    outputs(5259) <= b and not a;
    outputs(5260) <= not (a xor b);
    outputs(5261) <= a xor b;
    outputs(5262) <= a;
    outputs(5263) <= not a;
    outputs(5264) <= b;
    outputs(5265) <= a xor b;
    outputs(5266) <= not b or a;
    outputs(5267) <= not a or b;
    outputs(5268) <= a and b;
    outputs(5269) <= not (a xor b);
    outputs(5270) <= not (a xor b);
    outputs(5271) <= a;
    outputs(5272) <= not (a xor b);
    outputs(5273) <= not a or b;
    outputs(5274) <= a xor b;
    outputs(5275) <= not a or b;
    outputs(5276) <= not (a and b);
    outputs(5277) <= b;
    outputs(5278) <= a xor b;
    outputs(5279) <= not a;
    outputs(5280) <= a and b;
    outputs(5281) <= not a or b;
    outputs(5282) <= b and not a;
    outputs(5283) <= not (a or b);
    outputs(5284) <= b and not a;
    outputs(5285) <= a;
    outputs(5286) <= a;
    outputs(5287) <= b;
    outputs(5288) <= a xor b;
    outputs(5289) <= not a or b;
    outputs(5290) <= not a;
    outputs(5291) <= not a;
    outputs(5292) <= a;
    outputs(5293) <= a xor b;
    outputs(5294) <= a xor b;
    outputs(5295) <= a;
    outputs(5296) <= a and not b;
    outputs(5297) <= not (a or b);
    outputs(5298) <= a xor b;
    outputs(5299) <= a xor b;
    outputs(5300) <= a xor b;
    outputs(5301) <= not b or a;
    outputs(5302) <= a or b;
    outputs(5303) <= not (a xor b);
    outputs(5304) <= b;
    outputs(5305) <= not a;
    outputs(5306) <= a xor b;
    outputs(5307) <= not (a and b);
    outputs(5308) <= a xor b;
    outputs(5309) <= a and not b;
    outputs(5310) <= a xor b;
    outputs(5311) <= not (a xor b);
    outputs(5312) <= b and not a;
    outputs(5313) <= a;
    outputs(5314) <= b;
    outputs(5315) <= not (a and b);
    outputs(5316) <= not (a xor b);
    outputs(5317) <= not (a or b);
    outputs(5318) <= a or b;
    outputs(5319) <= a and not b;
    outputs(5320) <= b and not a;
    outputs(5321) <= not a;
    outputs(5322) <= not (a and b);
    outputs(5323) <= a and b;
    outputs(5324) <= a xor b;
    outputs(5325) <= b;
    outputs(5326) <= not (a and b);
    outputs(5327) <= b;
    outputs(5328) <= a;
    outputs(5329) <= not (a xor b);
    outputs(5330) <= not b;
    outputs(5331) <= not b;
    outputs(5332) <= a;
    outputs(5333) <= a;
    outputs(5334) <= not b;
    outputs(5335) <= not b;
    outputs(5336) <= a xor b;
    outputs(5337) <= a;
    outputs(5338) <= not b;
    outputs(5339) <= a and b;
    outputs(5340) <= not (a and b);
    outputs(5341) <= not b;
    outputs(5342) <= a xor b;
    outputs(5343) <= not a;
    outputs(5344) <= a and not b;
    outputs(5345) <= not b;
    outputs(5346) <= not b or a;
    outputs(5347) <= not (a xor b);
    outputs(5348) <= a xor b;
    outputs(5349) <= a;
    outputs(5350) <= not a;
    outputs(5351) <= a or b;
    outputs(5352) <= a or b;
    outputs(5353) <= a xor b;
    outputs(5354) <= a and b;
    outputs(5355) <= not b;
    outputs(5356) <= b and not a;
    outputs(5357) <= not a;
    outputs(5358) <= b and not a;
    outputs(5359) <= not b;
    outputs(5360) <= not (a or b);
    outputs(5361) <= not b;
    outputs(5362) <= b;
    outputs(5363) <= not (a xor b);
    outputs(5364) <= a;
    outputs(5365) <= not (a xor b);
    outputs(5366) <= a and not b;
    outputs(5367) <= a;
    outputs(5368) <= not (a or b);
    outputs(5369) <= a xor b;
    outputs(5370) <= b and not a;
    outputs(5371) <= b;
    outputs(5372) <= a xor b;
    outputs(5373) <= not (a xor b);
    outputs(5374) <= not (a xor b);
    outputs(5375) <= b and not a;
    outputs(5376) <= not a or b;
    outputs(5377) <= a;
    outputs(5378) <= a xor b;
    outputs(5379) <= a or b;
    outputs(5380) <= a xor b;
    outputs(5381) <= not (a xor b);
    outputs(5382) <= a and not b;
    outputs(5383) <= a;
    outputs(5384) <= not (a and b);
    outputs(5385) <= not a;
    outputs(5386) <= not b;
    outputs(5387) <= b;
    outputs(5388) <= a;
    outputs(5389) <= b;
    outputs(5390) <= a and not b;
    outputs(5391) <= b;
    outputs(5392) <= a and b;
    outputs(5393) <= b;
    outputs(5394) <= not b;
    outputs(5395) <= a or b;
    outputs(5396) <= not a;
    outputs(5397) <= a xor b;
    outputs(5398) <= b and not a;
    outputs(5399) <= a and b;
    outputs(5400) <= a xor b;
    outputs(5401) <= a and b;
    outputs(5402) <= not (a xor b);
    outputs(5403) <= b;
    outputs(5404) <= b;
    outputs(5405) <= b;
    outputs(5406) <= a xor b;
    outputs(5407) <= a and not b;
    outputs(5408) <= b;
    outputs(5409) <= not a;
    outputs(5410) <= a xor b;
    outputs(5411) <= not a;
    outputs(5412) <= b and not a;
    outputs(5413) <= a xor b;
    outputs(5414) <= not (a xor b);
    outputs(5415) <= b and not a;
    outputs(5416) <= not (a or b);
    outputs(5417) <= not b;
    outputs(5418) <= not (a xor b);
    outputs(5419) <= not (a xor b);
    outputs(5420) <= not b;
    outputs(5421) <= not b;
    outputs(5422) <= not b or a;
    outputs(5423) <= not (a or b);
    outputs(5424) <= b and not a;
    outputs(5425) <= not (a xor b);
    outputs(5426) <= a xor b;
    outputs(5427) <= a xor b;
    outputs(5428) <= not (a xor b);
    outputs(5429) <= not b;
    outputs(5430) <= not a;
    outputs(5431) <= not (a and b);
    outputs(5432) <= a xor b;
    outputs(5433) <= not b or a;
    outputs(5434) <= not (a xor b);
    outputs(5435) <= not (a xor b);
    outputs(5436) <= not b;
    outputs(5437) <= not (a xor b);
    outputs(5438) <= not a;
    outputs(5439) <= not b or a;
    outputs(5440) <= not a;
    outputs(5441) <= a or b;
    outputs(5442) <= not b or a;
    outputs(5443) <= a xor b;
    outputs(5444) <= a and not b;
    outputs(5445) <= not a;
    outputs(5446) <= not b;
    outputs(5447) <= not (a xor b);
    outputs(5448) <= b and not a;
    outputs(5449) <= not (a xor b);
    outputs(5450) <= not a;
    outputs(5451) <= not (a and b);
    outputs(5452) <= a;
    outputs(5453) <= not (a xor b);
    outputs(5454) <= a;
    outputs(5455) <= a xor b;
    outputs(5456) <= not a or b;
    outputs(5457) <= a and not b;
    outputs(5458) <= not (a and b);
    outputs(5459) <= b and not a;
    outputs(5460) <= not (a xor b);
    outputs(5461) <= a and b;
    outputs(5462) <= not (a or b);
    outputs(5463) <= not a;
    outputs(5464) <= not (a or b);
    outputs(5465) <= a;
    outputs(5466) <= not (a xor b);
    outputs(5467) <= a or b;
    outputs(5468) <= not b;
    outputs(5469) <= a;
    outputs(5470) <= not (a and b);
    outputs(5471) <= a and not b;
    outputs(5472) <= not b;
    outputs(5473) <= a;
    outputs(5474) <= b and not a;
    outputs(5475) <= not b;
    outputs(5476) <= not a;
    outputs(5477) <= a;
    outputs(5478) <= a and not b;
    outputs(5479) <= not b or a;
    outputs(5480) <= not a;
    outputs(5481) <= a;
    outputs(5482) <= a and not b;
    outputs(5483) <= not a;
    outputs(5484) <= not a;
    outputs(5485) <= a;
    outputs(5486) <= not b;
    outputs(5487) <= not a or b;
    outputs(5488) <= b and not a;
    outputs(5489) <= not (a or b);
    outputs(5490) <= not (a xor b);
    outputs(5491) <= a;
    outputs(5492) <= a xor b;
    outputs(5493) <= b;
    outputs(5494) <= a xor b;
    outputs(5495) <= not a;
    outputs(5496) <= not (a or b);
    outputs(5497) <= a xor b;
    outputs(5498) <= a xor b;
    outputs(5499) <= not a;
    outputs(5500) <= b;
    outputs(5501) <= a xor b;
    outputs(5502) <= not b;
    outputs(5503) <= not (a and b);
    outputs(5504) <= not b;
    outputs(5505) <= not b;
    outputs(5506) <= a;
    outputs(5507) <= a;
    outputs(5508) <= a;
    outputs(5509) <= not (a or b);
    outputs(5510) <= not a;
    outputs(5511) <= not a;
    outputs(5512) <= a xor b;
    outputs(5513) <= a xor b;
    outputs(5514) <= b and not a;
    outputs(5515) <= not b;
    outputs(5516) <= '1';
    outputs(5517) <= a xor b;
    outputs(5518) <= not (a xor b);
    outputs(5519) <= not (a or b);
    outputs(5520) <= b;
    outputs(5521) <= b;
    outputs(5522) <= not a;
    outputs(5523) <= b;
    outputs(5524) <= a;
    outputs(5525) <= a xor b;
    outputs(5526) <= not (a or b);
    outputs(5527) <= not a or b;
    outputs(5528) <= not (a xor b);
    outputs(5529) <= not (a xor b);
    outputs(5530) <= not a;
    outputs(5531) <= a xor b;
    outputs(5532) <= not a or b;
    outputs(5533) <= not (a or b);
    outputs(5534) <= b and not a;
    outputs(5535) <= not (a xor b);
    outputs(5536) <= b;
    outputs(5537) <= a xor b;
    outputs(5538) <= a or b;
    outputs(5539) <= a and not b;
    outputs(5540) <= a;
    outputs(5541) <= a;
    outputs(5542) <= not (a and b);
    outputs(5543) <= not a;
    outputs(5544) <= not a or b;
    outputs(5545) <= not (a xor b);
    outputs(5546) <= not a;
    outputs(5547) <= a xor b;
    outputs(5548) <= not b or a;
    outputs(5549) <= not a or b;
    outputs(5550) <= a and b;
    outputs(5551) <= a;
    outputs(5552) <= a;
    outputs(5553) <= a;
    outputs(5554) <= not a or b;
    outputs(5555) <= a xor b;
    outputs(5556) <= a xor b;
    outputs(5557) <= a;
    outputs(5558) <= b and not a;
    outputs(5559) <= not a;
    outputs(5560) <= a xor b;
    outputs(5561) <= not b;
    outputs(5562) <= not b;
    outputs(5563) <= a or b;
    outputs(5564) <= a and not b;
    outputs(5565) <= not a;
    outputs(5566) <= b;
    outputs(5567) <= not a;
    outputs(5568) <= a and not b;
    outputs(5569) <= a or b;
    outputs(5570) <= b;
    outputs(5571) <= b;
    outputs(5572) <= not a;
    outputs(5573) <= not a;
    outputs(5574) <= not b;
    outputs(5575) <= a xor b;
    outputs(5576) <= a or b;
    outputs(5577) <= not b or a;
    outputs(5578) <= not a;
    outputs(5579) <= not b;
    outputs(5580) <= a and not b;
    outputs(5581) <= not a;
    outputs(5582) <= a;
    outputs(5583) <= b and not a;
    outputs(5584) <= a;
    outputs(5585) <= not b or a;
    outputs(5586) <= b;
    outputs(5587) <= a and b;
    outputs(5588) <= not (a and b);
    outputs(5589) <= a and not b;
    outputs(5590) <= not b or a;
    outputs(5591) <= a and b;
    outputs(5592) <= a;
    outputs(5593) <= b;
    outputs(5594) <= a xor b;
    outputs(5595) <= not (a xor b);
    outputs(5596) <= a or b;
    outputs(5597) <= b;
    outputs(5598) <= not b;
    outputs(5599) <= not (a or b);
    outputs(5600) <= a;
    outputs(5601) <= not a or b;
    outputs(5602) <= not (a xor b);
    outputs(5603) <= a and b;
    outputs(5604) <= a;
    outputs(5605) <= not (a xor b);
    outputs(5606) <= not b or a;
    outputs(5607) <= a and not b;
    outputs(5608) <= b;
    outputs(5609) <= not (a xor b);
    outputs(5610) <= a or b;
    outputs(5611) <= not b;
    outputs(5612) <= not (a and b);
    outputs(5613) <= a or b;
    outputs(5614) <= a and b;
    outputs(5615) <= not a;
    outputs(5616) <= not b or a;
    outputs(5617) <= a and b;
    outputs(5618) <= not (a or b);
    outputs(5619) <= not a;
    outputs(5620) <= b and not a;
    outputs(5621) <= not a or b;
    outputs(5622) <= not a;
    outputs(5623) <= a xor b;
    outputs(5624) <= a xor b;
    outputs(5625) <= a xor b;
    outputs(5626) <= a;
    outputs(5627) <= not b or a;
    outputs(5628) <= a;
    outputs(5629) <= a xor b;
    outputs(5630) <= a and not b;
    outputs(5631) <= a and not b;
    outputs(5632) <= not (a xor b);
    outputs(5633) <= not a;
    outputs(5634) <= b;
    outputs(5635) <= b and not a;
    outputs(5636) <= a and not b;
    outputs(5637) <= b and not a;
    outputs(5638) <= not a;
    outputs(5639) <= a xor b;
    outputs(5640) <= not (a xor b);
    outputs(5641) <= a xor b;
    outputs(5642) <= not a;
    outputs(5643) <= a or b;
    outputs(5644) <= b;
    outputs(5645) <= a and b;
    outputs(5646) <= a xor b;
    outputs(5647) <= not a;
    outputs(5648) <= a xor b;
    outputs(5649) <= a xor b;
    outputs(5650) <= not b;
    outputs(5651) <= b and not a;
    outputs(5652) <= a;
    outputs(5653) <= not b;
    outputs(5654) <= a xor b;
    outputs(5655) <= not (a and b);
    outputs(5656) <= a and not b;
    outputs(5657) <= not a;
    outputs(5658) <= not b;
    outputs(5659) <= not b;
    outputs(5660) <= a xor b;
    outputs(5661) <= b;
    outputs(5662) <= b and not a;
    outputs(5663) <= not b or a;
    outputs(5664) <= not a;
    outputs(5665) <= a xor b;
    outputs(5666) <= a;
    outputs(5667) <= not (a xor b);
    outputs(5668) <= a xor b;
    outputs(5669) <= b and not a;
    outputs(5670) <= a xor b;
    outputs(5671) <= not b;
    outputs(5672) <= not b;
    outputs(5673) <= not b or a;
    outputs(5674) <= not a;
    outputs(5675) <= b and not a;
    outputs(5676) <= not a;
    outputs(5677) <= a and b;
    outputs(5678) <= a xor b;
    outputs(5679) <= a;
    outputs(5680) <= not (a and b);
    outputs(5681) <= a;
    outputs(5682) <= a or b;
    outputs(5683) <= a;
    outputs(5684) <= not (a and b);
    outputs(5685) <= a xor b;
    outputs(5686) <= not b;
    outputs(5687) <= not (a xor b);
    outputs(5688) <= not b;
    outputs(5689) <= not (a xor b);
    outputs(5690) <= a and not b;
    outputs(5691) <= b and not a;
    outputs(5692) <= a xor b;
    outputs(5693) <= not b;
    outputs(5694) <= not (a xor b);
    outputs(5695) <= a xor b;
    outputs(5696) <= not (a xor b);
    outputs(5697) <= not (a or b);
    outputs(5698) <= not a;
    outputs(5699) <= a xor b;
    outputs(5700) <= a;
    outputs(5701) <= a xor b;
    outputs(5702) <= not (a xor b);
    outputs(5703) <= a and not b;
    outputs(5704) <= not a;
    outputs(5705) <= not (a xor b);
    outputs(5706) <= a;
    outputs(5707) <= not (a xor b);
    outputs(5708) <= not b;
    outputs(5709) <= not (a xor b);
    outputs(5710) <= b;
    outputs(5711) <= not b or a;
    outputs(5712) <= not (a or b);
    outputs(5713) <= not b;
    outputs(5714) <= a and not b;
    outputs(5715) <= not (a xor b);
    outputs(5716) <= not a;
    outputs(5717) <= not a or b;
    outputs(5718) <= not (a xor b);
    outputs(5719) <= not (a xor b);
    outputs(5720) <= a;
    outputs(5721) <= not b;
    outputs(5722) <= not (a xor b);
    outputs(5723) <= b;
    outputs(5724) <= a xor b;
    outputs(5725) <= b;
    outputs(5726) <= a and not b;
    outputs(5727) <= not (a xor b);
    outputs(5728) <= not (a and b);
    outputs(5729) <= a xor b;
    outputs(5730) <= a xor b;
    outputs(5731) <= a and not b;
    outputs(5732) <= not (a xor b);
    outputs(5733) <= not (a and b);
    outputs(5734) <= not a;
    outputs(5735) <= not a;
    outputs(5736) <= a;
    outputs(5737) <= not (a or b);
    outputs(5738) <= not b;
    outputs(5739) <= b;
    outputs(5740) <= not (a or b);
    outputs(5741) <= not b;
    outputs(5742) <= a xor b;
    outputs(5743) <= a xor b;
    outputs(5744) <= b;
    outputs(5745) <= a xor b;
    outputs(5746) <= a and not b;
    outputs(5747) <= not a;
    outputs(5748) <= b;
    outputs(5749) <= b;
    outputs(5750) <= not (a xor b);
    outputs(5751) <= not (a xor b);
    outputs(5752) <= not (a xor b);
    outputs(5753) <= not b or a;
    outputs(5754) <= b;
    outputs(5755) <= a;
    outputs(5756) <= not (a and b);
    outputs(5757) <= a xor b;
    outputs(5758) <= not b;
    outputs(5759) <= b;
    outputs(5760) <= a;
    outputs(5761) <= not b;
    outputs(5762) <= a;
    outputs(5763) <= a xor b;
    outputs(5764) <= not b;
    outputs(5765) <= not (a xor b);
    outputs(5766) <= not a;
    outputs(5767) <= not (a xor b);
    outputs(5768) <= not a or b;
    outputs(5769) <= a xor b;
    outputs(5770) <= not a;
    outputs(5771) <= a xor b;
    outputs(5772) <= not (a and b);
    outputs(5773) <= a xor b;
    outputs(5774) <= not b;
    outputs(5775) <= a xor b;
    outputs(5776) <= not (a xor b);
    outputs(5777) <= not (a and b);
    outputs(5778) <= not (a xor b);
    outputs(5779) <= a or b;
    outputs(5780) <= a and not b;
    outputs(5781) <= not a;
    outputs(5782) <= b;
    outputs(5783) <= b and not a;
    outputs(5784) <= not a;
    outputs(5785) <= not (a or b);
    outputs(5786) <= a xor b;
    outputs(5787) <= not b;
    outputs(5788) <= a xor b;
    outputs(5789) <= not (a xor b);
    outputs(5790) <= not a or b;
    outputs(5791) <= a and not b;
    outputs(5792) <= not (a xor b);
    outputs(5793) <= not a;
    outputs(5794) <= a;
    outputs(5795) <= not a or b;
    outputs(5796) <= not a or b;
    outputs(5797) <= b;
    outputs(5798) <= not (a xor b);
    outputs(5799) <= a;
    outputs(5800) <= a xor b;
    outputs(5801) <= not (a xor b);
    outputs(5802) <= a xor b;
    outputs(5803) <= not (a xor b);
    outputs(5804) <= not (a or b);
    outputs(5805) <= a;
    outputs(5806) <= not b or a;
    outputs(5807) <= not b;
    outputs(5808) <= a or b;
    outputs(5809) <= not (a xor b);
    outputs(5810) <= not a;
    outputs(5811) <= not (a and b);
    outputs(5812) <= a xor b;
    outputs(5813) <= not b;
    outputs(5814) <= not (a xor b);
    outputs(5815) <= not (a xor b);
    outputs(5816) <= not a or b;
    outputs(5817) <= b;
    outputs(5818) <= not b;
    outputs(5819) <= a or b;
    outputs(5820) <= a and not b;
    outputs(5821) <= a and b;
    outputs(5822) <= not a;
    outputs(5823) <= a xor b;
    outputs(5824) <= b;
    outputs(5825) <= b and not a;
    outputs(5826) <= a and b;
    outputs(5827) <= a xor b;
    outputs(5828) <= not (a xor b);
    outputs(5829) <= not (a xor b);
    outputs(5830) <= a xor b;
    outputs(5831) <= b and not a;
    outputs(5832) <= a;
    outputs(5833) <= a xor b;
    outputs(5834) <= a and not b;
    outputs(5835) <= not (a xor b);
    outputs(5836) <= b;
    outputs(5837) <= not b or a;
    outputs(5838) <= a;
    outputs(5839) <= not a or b;
    outputs(5840) <= a and b;
    outputs(5841) <= not (a xor b);
    outputs(5842) <= a and b;
    outputs(5843) <= b;
    outputs(5844) <= not (a or b);
    outputs(5845) <= a and not b;
    outputs(5846) <= not (a xor b);
    outputs(5847) <= not a;
    outputs(5848) <= b and not a;
    outputs(5849) <= not (a xor b);
    outputs(5850) <= not b;
    outputs(5851) <= not (a xor b);
    outputs(5852) <= not (a xor b);
    outputs(5853) <= not b or a;
    outputs(5854) <= a;
    outputs(5855) <= not (a xor b);
    outputs(5856) <= not a or b;
    outputs(5857) <= a xor b;
    outputs(5858) <= not (a xor b);
    outputs(5859) <= not (a xor b);
    outputs(5860) <= not a;
    outputs(5861) <= b and not a;
    outputs(5862) <= b;
    outputs(5863) <= not b;
    outputs(5864) <= not a;
    outputs(5865) <= a xor b;
    outputs(5866) <= not a;
    outputs(5867) <= a xor b;
    outputs(5868) <= not b;
    outputs(5869) <= b;
    outputs(5870) <= a;
    outputs(5871) <= not (a xor b);
    outputs(5872) <= a;
    outputs(5873) <= b;
    outputs(5874) <= not b or a;
    outputs(5875) <= not (a or b);
    outputs(5876) <= a;
    outputs(5877) <= '1';
    outputs(5878) <= not a;
    outputs(5879) <= a;
    outputs(5880) <= a and not b;
    outputs(5881) <= not (a xor b);
    outputs(5882) <= a or b;
    outputs(5883) <= not (a xor b);
    outputs(5884) <= not (a xor b);
    outputs(5885) <= a and not b;
    outputs(5886) <= a xor b;
    outputs(5887) <= not b;
    outputs(5888) <= a xor b;
    outputs(5889) <= a;
    outputs(5890) <= not b;
    outputs(5891) <= not (a or b);
    outputs(5892) <= not (a xor b);
    outputs(5893) <= a and not b;
    outputs(5894) <= not a;
    outputs(5895) <= a;
    outputs(5896) <= not a or b;
    outputs(5897) <= not b or a;
    outputs(5898) <= not b;
    outputs(5899) <= not a;
    outputs(5900) <= not a;
    outputs(5901) <= a xor b;
    outputs(5902) <= not (a or b);
    outputs(5903) <= b;
    outputs(5904) <= b;
    outputs(5905) <= a xor b;
    outputs(5906) <= a xor b;
    outputs(5907) <= not (a and b);
    outputs(5908) <= not a;
    outputs(5909) <= not (a or b);
    outputs(5910) <= a xor b;
    outputs(5911) <= a and b;
    outputs(5912) <= a;
    outputs(5913) <= a;
    outputs(5914) <= a;
    outputs(5915) <= not b or a;
    outputs(5916) <= not (a xor b);
    outputs(5917) <= not (a xor b);
    outputs(5918) <= not (a or b);
    outputs(5919) <= a and b;
    outputs(5920) <= not (a xor b);
    outputs(5921) <= not (a xor b);
    outputs(5922) <= a and not b;
    outputs(5923) <= not a;
    outputs(5924) <= b;
    outputs(5925) <= b and not a;
    outputs(5926) <= not a;
    outputs(5927) <= a or b;
    outputs(5928) <= a xor b;
    outputs(5929) <= b;
    outputs(5930) <= a and b;
    outputs(5931) <= a and not b;
    outputs(5932) <= b;
    outputs(5933) <= not (a xor b);
    outputs(5934) <= a and not b;
    outputs(5935) <= a and b;
    outputs(5936) <= not (a xor b);
    outputs(5937) <= a;
    outputs(5938) <= not (a xor b);
    outputs(5939) <= a or b;
    outputs(5940) <= not b or a;
    outputs(5941) <= a xor b;
    outputs(5942) <= not (a xor b);
    outputs(5943) <= b and not a;
    outputs(5944) <= not b;
    outputs(5945) <= not (a xor b);
    outputs(5946) <= a;
    outputs(5947) <= a xor b;
    outputs(5948) <= a xor b;
    outputs(5949) <= a;
    outputs(5950) <= a;
    outputs(5951) <= not b;
    outputs(5952) <= not (a xor b);
    outputs(5953) <= b;
    outputs(5954) <= not (a xor b);
    outputs(5955) <= a;
    outputs(5956) <= a xor b;
    outputs(5957) <= a or b;
    outputs(5958) <= a xor b;
    outputs(5959) <= not a;
    outputs(5960) <= not (a or b);
    outputs(5961) <= not b or a;
    outputs(5962) <= a xor b;
    outputs(5963) <= a and not b;
    outputs(5964) <= a xor b;
    outputs(5965) <= not a;
    outputs(5966) <= a;
    outputs(5967) <= a;
    outputs(5968) <= a or b;
    outputs(5969) <= a and b;
    outputs(5970) <= not b;
    outputs(5971) <= not a;
    outputs(5972) <= not a;
    outputs(5973) <= not a;
    outputs(5974) <= b;
    outputs(5975) <= b;
    outputs(5976) <= a xor b;
    outputs(5977) <= a;
    outputs(5978) <= a xor b;
    outputs(5979) <= not (a xor b);
    outputs(5980) <= a and b;
    outputs(5981) <= not a;
    outputs(5982) <= a;
    outputs(5983) <= a and not b;
    outputs(5984) <= b and not a;
    outputs(5985) <= not (a xor b);
    outputs(5986) <= b;
    outputs(5987) <= a or b;
    outputs(5988) <= not b;
    outputs(5989) <= not (a xor b);
    outputs(5990) <= not (a or b);
    outputs(5991) <= not (a xor b);
    outputs(5992) <= a xor b;
    outputs(5993) <= a xor b;
    outputs(5994) <= a or b;
    outputs(5995) <= not a;
    outputs(5996) <= not (a xor b);
    outputs(5997) <= a xor b;
    outputs(5998) <= a xor b;
    outputs(5999) <= a;
    outputs(6000) <= not (a and b);
    outputs(6001) <= not (a xor b);
    outputs(6002) <= a xor b;
    outputs(6003) <= not (a xor b);
    outputs(6004) <= not a;
    outputs(6005) <= not b or a;
    outputs(6006) <= not (a and b);
    outputs(6007) <= not (a xor b);
    outputs(6008) <= b;
    outputs(6009) <= not (a xor b);
    outputs(6010) <= not (a xor b);
    outputs(6011) <= a xor b;
    outputs(6012) <= a xor b;
    outputs(6013) <= a;
    outputs(6014) <= not a;
    outputs(6015) <= b;
    outputs(6016) <= not b;
    outputs(6017) <= not (a xor b);
    outputs(6018) <= not a or b;
    outputs(6019) <= not a;
    outputs(6020) <= not (a xor b);
    outputs(6021) <= a;
    outputs(6022) <= not (a or b);
    outputs(6023) <= a;
    outputs(6024) <= a and b;
    outputs(6025) <= b;
    outputs(6026) <= a xor b;
    outputs(6027) <= not (a xor b);
    outputs(6028) <= b and not a;
    outputs(6029) <= not (a xor b);
    outputs(6030) <= not a;
    outputs(6031) <= not b;
    outputs(6032) <= a and not b;
    outputs(6033) <= not b;
    outputs(6034) <= not b or a;
    outputs(6035) <= a xor b;
    outputs(6036) <= not a or b;
    outputs(6037) <= b;
    outputs(6038) <= a and b;
    outputs(6039) <= b;
    outputs(6040) <= b;
    outputs(6041) <= a xor b;
    outputs(6042) <= a xor b;
    outputs(6043) <= not (a xor b);
    outputs(6044) <= not (a and b);
    outputs(6045) <= a and not b;
    outputs(6046) <= a and not b;
    outputs(6047) <= a xor b;
    outputs(6048) <= not a;
    outputs(6049) <= not (a xor b);
    outputs(6050) <= a xor b;
    outputs(6051) <= not (a or b);
    outputs(6052) <= not b or a;
    outputs(6053) <= b;
    outputs(6054) <= not (a xor b);
    outputs(6055) <= a or b;
    outputs(6056) <= not (a xor b);
    outputs(6057) <= a xor b;
    outputs(6058) <= a or b;
    outputs(6059) <= b and not a;
    outputs(6060) <= b;
    outputs(6061) <= '0';
    outputs(6062) <= not b or a;
    outputs(6063) <= a xor b;
    outputs(6064) <= not b;
    outputs(6065) <= b;
    outputs(6066) <= a or b;
    outputs(6067) <= not (a xor b);
    outputs(6068) <= a and not b;
    outputs(6069) <= not (a or b);
    outputs(6070) <= b and not a;
    outputs(6071) <= a xor b;
    outputs(6072) <= not b or a;
    outputs(6073) <= not (a xor b);
    outputs(6074) <= b;
    outputs(6075) <= not a;
    outputs(6076) <= not (a xor b);
    outputs(6077) <= b and not a;
    outputs(6078) <= not a or b;
    outputs(6079) <= not a;
    outputs(6080) <= not a;
    outputs(6081) <= not (a xor b);
    outputs(6082) <= not a;
    outputs(6083) <= not (a xor b);
    outputs(6084) <= not (a xor b);
    outputs(6085) <= not a;
    outputs(6086) <= a and not b;
    outputs(6087) <= b;
    outputs(6088) <= not a;
    outputs(6089) <= a;
    outputs(6090) <= not (a xor b);
    outputs(6091) <= b;
    outputs(6092) <= not a or b;
    outputs(6093) <= not a;
    outputs(6094) <= a xor b;
    outputs(6095) <= a or b;
    outputs(6096) <= not a;
    outputs(6097) <= not a;
    outputs(6098) <= a xor b;
    outputs(6099) <= a and b;
    outputs(6100) <= not (a xor b);
    outputs(6101) <= b and not a;
    outputs(6102) <= not a;
    outputs(6103) <= not b or a;
    outputs(6104) <= a xor b;
    outputs(6105) <= not (a xor b);
    outputs(6106) <= not a;
    outputs(6107) <= a xor b;
    outputs(6108) <= b;
    outputs(6109) <= not (a or b);
    outputs(6110) <= not a or b;
    outputs(6111) <= b;
    outputs(6112) <= not (a xor b);
    outputs(6113) <= a and b;
    outputs(6114) <= not b;
    outputs(6115) <= not (a or b);
    outputs(6116) <= not a;
    outputs(6117) <= not b or a;
    outputs(6118) <= not (a xor b);
    outputs(6119) <= not (a xor b);
    outputs(6120) <= a and not b;
    outputs(6121) <= not a or b;
    outputs(6122) <= a xor b;
    outputs(6123) <= b and not a;
    outputs(6124) <= a xor b;
    outputs(6125) <= not b;
    outputs(6126) <= a or b;
    outputs(6127) <= a xor b;
    outputs(6128) <= a or b;
    outputs(6129) <= a xor b;
    outputs(6130) <= not (a or b);
    outputs(6131) <= a and b;
    outputs(6132) <= not a;
    outputs(6133) <= not b;
    outputs(6134) <= not a or b;
    outputs(6135) <= not b or a;
    outputs(6136) <= not (a xor b);
    outputs(6137) <= not (a xor b);
    outputs(6138) <= not b or a;
    outputs(6139) <= not (a xor b);
    outputs(6140) <= not a;
    outputs(6141) <= not a;
    outputs(6142) <= b;
    outputs(6143) <= not b;
    outputs(6144) <= not (a xor b);
    outputs(6145) <= a and b;
    outputs(6146) <= b;
    outputs(6147) <= a or b;
    outputs(6148) <= not (a xor b);
    outputs(6149) <= a xor b;
    outputs(6150) <= a and not b;
    outputs(6151) <= a xor b;
    outputs(6152) <= a and not b;
    outputs(6153) <= not (a or b);
    outputs(6154) <= a xor b;
    outputs(6155) <= b;
    outputs(6156) <= not a or b;
    outputs(6157) <= a;
    outputs(6158) <= b;
    outputs(6159) <= a and b;
    outputs(6160) <= not (a xor b);
    outputs(6161) <= not (a xor b);
    outputs(6162) <= not a;
    outputs(6163) <= not b;
    outputs(6164) <= a;
    outputs(6165) <= not a;
    outputs(6166) <= not b or a;
    outputs(6167) <= not a;
    outputs(6168) <= not b;
    outputs(6169) <= a;
    outputs(6170) <= not b;
    outputs(6171) <= not (a and b);
    outputs(6172) <= not b;
    outputs(6173) <= not a;
    outputs(6174) <= not (a xor b);
    outputs(6175) <= b;
    outputs(6176) <= not a;
    outputs(6177) <= a;
    outputs(6178) <= a xor b;
    outputs(6179) <= a;
    outputs(6180) <= not b;
    outputs(6181) <= not b;
    outputs(6182) <= not b;
    outputs(6183) <= not (a xor b);
    outputs(6184) <= not (a and b);
    outputs(6185) <= not (a xor b);
    outputs(6186) <= b and not a;
    outputs(6187) <= not b;
    outputs(6188) <= not b;
    outputs(6189) <= not (a or b);
    outputs(6190) <= a and not b;
    outputs(6191) <= not a;
    outputs(6192) <= a xor b;
    outputs(6193) <= not (a xor b);
    outputs(6194) <= a or b;
    outputs(6195) <= b and not a;
    outputs(6196) <= b;
    outputs(6197) <= not (a xor b);
    outputs(6198) <= not b;
    outputs(6199) <= not b;
    outputs(6200) <= not a;
    outputs(6201) <= not b;
    outputs(6202) <= not b or a;
    outputs(6203) <= a;
    outputs(6204) <= not b;
    outputs(6205) <= a and not b;
    outputs(6206) <= b;
    outputs(6207) <= a and b;
    outputs(6208) <= not b;
    outputs(6209) <= not a;
    outputs(6210) <= b;
    outputs(6211) <= not (a and b);
    outputs(6212) <= not (a xor b);
    outputs(6213) <= a xor b;
    outputs(6214) <= not b;
    outputs(6215) <= not b;
    outputs(6216) <= a or b;
    outputs(6217) <= not (a xor b);
    outputs(6218) <= a xor b;
    outputs(6219) <= a;
    outputs(6220) <= a or b;
    outputs(6221) <= a or b;
    outputs(6222) <= b;
    outputs(6223) <= not b;
    outputs(6224) <= a and b;
    outputs(6225) <= not (a xor b);
    outputs(6226) <= a and not b;
    outputs(6227) <= not b;
    outputs(6228) <= not (a xor b);
    outputs(6229) <= not (a or b);
    outputs(6230) <= not (a or b);
    outputs(6231) <= not (a xor b);
    outputs(6232) <= a and not b;
    outputs(6233) <= a;
    outputs(6234) <= not a;
    outputs(6235) <= not (a and b);
    outputs(6236) <= not a;
    outputs(6237) <= a and not b;
    outputs(6238) <= a and not b;
    outputs(6239) <= a;
    outputs(6240) <= not (a or b);
    outputs(6241) <= b;
    outputs(6242) <= a and b;
    outputs(6243) <= not (a xor b);
    outputs(6244) <= a or b;
    outputs(6245) <= not (a or b);
    outputs(6246) <= not b;
    outputs(6247) <= a or b;
    outputs(6248) <= not (a or b);
    outputs(6249) <= a;
    outputs(6250) <= a and not b;
    outputs(6251) <= not (a or b);
    outputs(6252) <= a;
    outputs(6253) <= a;
    outputs(6254) <= not a;
    outputs(6255) <= a;
    outputs(6256) <= not a;
    outputs(6257) <= a xor b;
    outputs(6258) <= b and not a;
    outputs(6259) <= b;
    outputs(6260) <= not b;
    outputs(6261) <= a and not b;
    outputs(6262) <= a xor b;
    outputs(6263) <= not a;
    outputs(6264) <= not b or a;
    outputs(6265) <= not (a xor b);
    outputs(6266) <= not (a xor b);
    outputs(6267) <= a and not b;
    outputs(6268) <= not (a or b);
    outputs(6269) <= a and b;
    outputs(6270) <= not a;
    outputs(6271) <= not b;
    outputs(6272) <= a xor b;
    outputs(6273) <= not a or b;
    outputs(6274) <= not (a xor b);
    outputs(6275) <= a and not b;
    outputs(6276) <= not a or b;
    outputs(6277) <= a;
    outputs(6278) <= a xor b;
    outputs(6279) <= not (a xor b);
    outputs(6280) <= not b;
    outputs(6281) <= not (a xor b);
    outputs(6282) <= not a;
    outputs(6283) <= b;
    outputs(6284) <= b;
    outputs(6285) <= not b;
    outputs(6286) <= not (a or b);
    outputs(6287) <= a and b;
    outputs(6288) <= a xor b;
    outputs(6289) <= not (a and b);
    outputs(6290) <= a;
    outputs(6291) <= b;
    outputs(6292) <= not (a xor b);
    outputs(6293) <= not (a or b);
    outputs(6294) <= not a;
    outputs(6295) <= b;
    outputs(6296) <= not (a xor b);
    outputs(6297) <= b;
    outputs(6298) <= a;
    outputs(6299) <= not a;
    outputs(6300) <= not (a or b);
    outputs(6301) <= a;
    outputs(6302) <= b and not a;
    outputs(6303) <= b;
    outputs(6304) <= not b;
    outputs(6305) <= a and not b;
    outputs(6306) <= not (a xor b);
    outputs(6307) <= not (a or b);
    outputs(6308) <= a xor b;
    outputs(6309) <= not b;
    outputs(6310) <= not (a xor b);
    outputs(6311) <= b;
    outputs(6312) <= not b;
    outputs(6313) <= a and b;
    outputs(6314) <= a and b;
    outputs(6315) <= not a;
    outputs(6316) <= b;
    outputs(6317) <= a;
    outputs(6318) <= a and not b;
    outputs(6319) <= b;
    outputs(6320) <= b;
    outputs(6321) <= a;
    outputs(6322) <= not a;
    outputs(6323) <= not a;
    outputs(6324) <= not (a and b);
    outputs(6325) <= not (a xor b);
    outputs(6326) <= a xor b;
    outputs(6327) <= a xor b;
    outputs(6328) <= a xor b;
    outputs(6329) <= a xor b;
    outputs(6330) <= b and not a;
    outputs(6331) <= a xor b;
    outputs(6332) <= a xor b;
    outputs(6333) <= a xor b;
    outputs(6334) <= not (a or b);
    outputs(6335) <= not (a and b);
    outputs(6336) <= not (a and b);
    outputs(6337) <= a xor b;
    outputs(6338) <= not a;
    outputs(6339) <= not (a xor b);
    outputs(6340) <= not a;
    outputs(6341) <= not b;
    outputs(6342) <= b;
    outputs(6343) <= b;
    outputs(6344) <= not b or a;
    outputs(6345) <= not b;
    outputs(6346) <= a xor b;
    outputs(6347) <= not b;
    outputs(6348) <= b and not a;
    outputs(6349) <= a;
    outputs(6350) <= not (a or b);
    outputs(6351) <= not (a or b);
    outputs(6352) <= a xor b;
    outputs(6353) <= not (a or b);
    outputs(6354) <= b and not a;
    outputs(6355) <= a;
    outputs(6356) <= a and b;
    outputs(6357) <= a and not b;
    outputs(6358) <= not b;
    outputs(6359) <= not (a xor b);
    outputs(6360) <= not (a or b);
    outputs(6361) <= a;
    outputs(6362) <= a xor b;
    outputs(6363) <= not a;
    outputs(6364) <= a;
    outputs(6365) <= a;
    outputs(6366) <= not (a xor b);
    outputs(6367) <= b;
    outputs(6368) <= not (a or b);
    outputs(6369) <= b and not a;
    outputs(6370) <= not b;
    outputs(6371) <= not a;
    outputs(6372) <= a xor b;
    outputs(6373) <= a and b;
    outputs(6374) <= a xor b;
    outputs(6375) <= not a or b;
    outputs(6376) <= b and not a;
    outputs(6377) <= a and b;
    outputs(6378) <= not a;
    outputs(6379) <= a and not b;
    outputs(6380) <= not b;
    outputs(6381) <= not b;
    outputs(6382) <= not (a xor b);
    outputs(6383) <= not (a xor b);
    outputs(6384) <= a;
    outputs(6385) <= a xor b;
    outputs(6386) <= not b;
    outputs(6387) <= not a;
    outputs(6388) <= not (a xor b);
    outputs(6389) <= not a;
    outputs(6390) <= b and not a;
    outputs(6391) <= not (a xor b);
    outputs(6392) <= a xor b;
    outputs(6393) <= not b or a;
    outputs(6394) <= not a;
    outputs(6395) <= a and b;
    outputs(6396) <= not a or b;
    outputs(6397) <= not (a xor b);
    outputs(6398) <= b;
    outputs(6399) <= not (a xor b);
    outputs(6400) <= not b or a;
    outputs(6401) <= not (a or b);
    outputs(6402) <= not (a or b);
    outputs(6403) <= a;
    outputs(6404) <= not (a and b);
    outputs(6405) <= not (a xor b);
    outputs(6406) <= b;
    outputs(6407) <= a;
    outputs(6408) <= not a;
    outputs(6409) <= a or b;
    outputs(6410) <= a xor b;
    outputs(6411) <= not (a and b);
    outputs(6412) <= a and b;
    outputs(6413) <= b;
    outputs(6414) <= b and not a;
    outputs(6415) <= not (a xor b);
    outputs(6416) <= a and not b;
    outputs(6417) <= not (a xor b);
    outputs(6418) <= a;
    outputs(6419) <= not (a xor b);
    outputs(6420) <= a and not b;
    outputs(6421) <= a xor b;
    outputs(6422) <= not b or a;
    outputs(6423) <= not (a xor b);
    outputs(6424) <= a xor b;
    outputs(6425) <= not b or a;
    outputs(6426) <= not (a and b);
    outputs(6427) <= a and not b;
    outputs(6428) <= not a;
    outputs(6429) <= a;
    outputs(6430) <= a;
    outputs(6431) <= a xor b;
    outputs(6432) <= not (a xor b);
    outputs(6433) <= a;
    outputs(6434) <= a xor b;
    outputs(6435) <= a xor b;
    outputs(6436) <= not b;
    outputs(6437) <= a;
    outputs(6438) <= a;
    outputs(6439) <= b;
    outputs(6440) <= a and not b;
    outputs(6441) <= a and b;
    outputs(6442) <= a xor b;
    outputs(6443) <= not a or b;
    outputs(6444) <= not b;
    outputs(6445) <= not a;
    outputs(6446) <= not (a xor b);
    outputs(6447) <= not (a xor b);
    outputs(6448) <= a;
    outputs(6449) <= a and not b;
    outputs(6450) <= not a or b;
    outputs(6451) <= a and not b;
    outputs(6452) <= not a or b;
    outputs(6453) <= a and not b;
    outputs(6454) <= not (a xor b);
    outputs(6455) <= not b or a;
    outputs(6456) <= a and not b;
    outputs(6457) <= a xor b;
    outputs(6458) <= not (a xor b);
    outputs(6459) <= a xor b;
    outputs(6460) <= a or b;
    outputs(6461) <= a and b;
    outputs(6462) <= b and not a;
    outputs(6463) <= not (a xor b);
    outputs(6464) <= not (a xor b);
    outputs(6465) <= not (a xor b);
    outputs(6466) <= a and not b;
    outputs(6467) <= b;
    outputs(6468) <= b and not a;
    outputs(6469) <= not (a xor b);
    outputs(6470) <= a xor b;
    outputs(6471) <= a xor b;
    outputs(6472) <= not (a and b);
    outputs(6473) <= not a;
    outputs(6474) <= not (a xor b);
    outputs(6475) <= a and b;
    outputs(6476) <= b;
    outputs(6477) <= a;
    outputs(6478) <= a and not b;
    outputs(6479) <= b;
    outputs(6480) <= a and not b;
    outputs(6481) <= b;
    outputs(6482) <= not (a xor b);
    outputs(6483) <= a and not b;
    outputs(6484) <= a xor b;
    outputs(6485) <= not b;
    outputs(6486) <= not (a xor b);
    outputs(6487) <= not b;
    outputs(6488) <= not (a xor b);
    outputs(6489) <= a;
    outputs(6490) <= a;
    outputs(6491) <= not (a xor b);
    outputs(6492) <= not a;
    outputs(6493) <= not b or a;
    outputs(6494) <= a xor b;
    outputs(6495) <= b and not a;
    outputs(6496) <= not (a xor b);
    outputs(6497) <= a and not b;
    outputs(6498) <= a and not b;
    outputs(6499) <= b;
    outputs(6500) <= not (a or b);
    outputs(6501) <= a xor b;
    outputs(6502) <= not b or a;
    outputs(6503) <= not (a or b);
    outputs(6504) <= not (a or b);
    outputs(6505) <= b and not a;
    outputs(6506) <= not (a or b);
    outputs(6507) <= not a;
    outputs(6508) <= not a;
    outputs(6509) <= a;
    outputs(6510) <= not a;
    outputs(6511) <= a or b;
    outputs(6512) <= a or b;
    outputs(6513) <= a xor b;
    outputs(6514) <= a or b;
    outputs(6515) <= not (a or b);
    outputs(6516) <= a xor b;
    outputs(6517) <= a xor b;
    outputs(6518) <= not (a xor b);
    outputs(6519) <= a xor b;
    outputs(6520) <= a and not b;
    outputs(6521) <= not a or b;
    outputs(6522) <= a or b;
    outputs(6523) <= not a;
    outputs(6524) <= a and b;
    outputs(6525) <= not a;
    outputs(6526) <= b;
    outputs(6527) <= a and b;
    outputs(6528) <= a or b;
    outputs(6529) <= not (a xor b);
    outputs(6530) <= b;
    outputs(6531) <= not a;
    outputs(6532) <= not a;
    outputs(6533) <= not (a or b);
    outputs(6534) <= not b;
    outputs(6535) <= a and b;
    outputs(6536) <= a and not b;
    outputs(6537) <= not (a xor b);
    outputs(6538) <= a;
    outputs(6539) <= not (a or b);
    outputs(6540) <= b;
    outputs(6541) <= not (a xor b);
    outputs(6542) <= b and not a;
    outputs(6543) <= not (a or b);
    outputs(6544) <= a xor b;
    outputs(6545) <= not (a xor b);
    outputs(6546) <= not (a xor b);
    outputs(6547) <= not a;
    outputs(6548) <= a;
    outputs(6549) <= a xor b;
    outputs(6550) <= a and not b;
    outputs(6551) <= a and b;
    outputs(6552) <= not b;
    outputs(6553) <= not (a xor b);
    outputs(6554) <= not b;
    outputs(6555) <= a and not b;
    outputs(6556) <= not (a xor b);
    outputs(6557) <= not b;
    outputs(6558) <= b;
    outputs(6559) <= b and not a;
    outputs(6560) <= a xor b;
    outputs(6561) <= a or b;
    outputs(6562) <= not b;
    outputs(6563) <= not (a and b);
    outputs(6564) <= b and not a;
    outputs(6565) <= not (a and b);
    outputs(6566) <= a;
    outputs(6567) <= not b;
    outputs(6568) <= b;
    outputs(6569) <= not b;
    outputs(6570) <= not (a and b);
    outputs(6571) <= b;
    outputs(6572) <= not b;
    outputs(6573) <= a xor b;
    outputs(6574) <= a;
    outputs(6575) <= a;
    outputs(6576) <= b;
    outputs(6577) <= not b;
    outputs(6578) <= not (a or b);
    outputs(6579) <= not (a or b);
    outputs(6580) <= not a;
    outputs(6581) <= a xor b;
    outputs(6582) <= a xor b;
    outputs(6583) <= a xor b;
    outputs(6584) <= a and not b;
    outputs(6585) <= a or b;
    outputs(6586) <= not a;
    outputs(6587) <= not b;
    outputs(6588) <= a xor b;
    outputs(6589) <= a;
    outputs(6590) <= a xor b;
    outputs(6591) <= a xor b;
    outputs(6592) <= a xor b;
    outputs(6593) <= a and not b;
    outputs(6594) <= not a or b;
    outputs(6595) <= not (a xor b);
    outputs(6596) <= not (a and b);
    outputs(6597) <= a;
    outputs(6598) <= a and b;
    outputs(6599) <= not (a xor b);
    outputs(6600) <= a xor b;
    outputs(6601) <= b;
    outputs(6602) <= not b;
    outputs(6603) <= not (a and b);
    outputs(6604) <= a;
    outputs(6605) <= not b;
    outputs(6606) <= not a;
    outputs(6607) <= not b;
    outputs(6608) <= a xor b;
    outputs(6609) <= a;
    outputs(6610) <= a;
    outputs(6611) <= not b;
    outputs(6612) <= a xor b;
    outputs(6613) <= not b;
    outputs(6614) <= b;
    outputs(6615) <= not b;
    outputs(6616) <= not a;
    outputs(6617) <= a and b;
    outputs(6618) <= a and b;
    outputs(6619) <= not (a xor b);
    outputs(6620) <= b and not a;
    outputs(6621) <= not b;
    outputs(6622) <= a xor b;
    outputs(6623) <= not (a or b);
    outputs(6624) <= b;
    outputs(6625) <= b;
    outputs(6626) <= a and not b;
    outputs(6627) <= a or b;
    outputs(6628) <= a or b;
    outputs(6629) <= b;
    outputs(6630) <= b;
    outputs(6631) <= a;
    outputs(6632) <= a and b;
    outputs(6633) <= b and not a;
    outputs(6634) <= not (a xor b);
    outputs(6635) <= not b;
    outputs(6636) <= not (a xor b);
    outputs(6637) <= not b or a;
    outputs(6638) <= b and not a;
    outputs(6639) <= b;
    outputs(6640) <= not a;
    outputs(6641) <= not a;
    outputs(6642) <= not (a or b);
    outputs(6643) <= not (a xor b);
    outputs(6644) <= not b;
    outputs(6645) <= a;
    outputs(6646) <= not a;
    outputs(6647) <= a xor b;
    outputs(6648) <= a xor b;
    outputs(6649) <= a xor b;
    outputs(6650) <= b;
    outputs(6651) <= not b;
    outputs(6652) <= a xor b;
    outputs(6653) <= a;
    outputs(6654) <= not b or a;
    outputs(6655) <= not (a xor b);
    outputs(6656) <= a;
    outputs(6657) <= a xor b;
    outputs(6658) <= a and not b;
    outputs(6659) <= a xor b;
    outputs(6660) <= not b;
    outputs(6661) <= not (a xor b);
    outputs(6662) <= not b or a;
    outputs(6663) <= a or b;
    outputs(6664) <= a and b;
    outputs(6665) <= a and not b;
    outputs(6666) <= a and b;
    outputs(6667) <= not b or a;
    outputs(6668) <= b and not a;
    outputs(6669) <= not b or a;
    outputs(6670) <= b and not a;
    outputs(6671) <= a and b;
    outputs(6672) <= b and not a;
    outputs(6673) <= not a or b;
    outputs(6674) <= not (a xor b);
    outputs(6675) <= a;
    outputs(6676) <= not b;
    outputs(6677) <= a and b;
    outputs(6678) <= a and not b;
    outputs(6679) <= not (a xor b);
    outputs(6680) <= a;
    outputs(6681) <= not b;
    outputs(6682) <= not b;
    outputs(6683) <= b and not a;
    outputs(6684) <= b;
    outputs(6685) <= b;
    outputs(6686) <= a;
    outputs(6687) <= not a or b;
    outputs(6688) <= not a or b;
    outputs(6689) <= a;
    outputs(6690) <= b;
    outputs(6691) <= b;
    outputs(6692) <= b and not a;
    outputs(6693) <= not a;
    outputs(6694) <= not (a xor b);
    outputs(6695) <= a xor b;
    outputs(6696) <= not (a and b);
    outputs(6697) <= a xor b;
    outputs(6698) <= not (a xor b);
    outputs(6699) <= not (a xor b);
    outputs(6700) <= not a or b;
    outputs(6701) <= not a;
    outputs(6702) <= a;
    outputs(6703) <= a xor b;
    outputs(6704) <= a xor b;
    outputs(6705) <= not (a xor b);
    outputs(6706) <= a and b;
    outputs(6707) <= b;
    outputs(6708) <= not (a xor b);
    outputs(6709) <= b and not a;
    outputs(6710) <= b;
    outputs(6711) <= b;
    outputs(6712) <= not b or a;
    outputs(6713) <= not (a xor b);
    outputs(6714) <= not b or a;
    outputs(6715) <= a or b;
    outputs(6716) <= a;
    outputs(6717) <= a;
    outputs(6718) <= a;
    outputs(6719) <= not (a xor b);
    outputs(6720) <= a or b;
    outputs(6721) <= not a or b;
    outputs(6722) <= b;
    outputs(6723) <= not a;
    outputs(6724) <= a xor b;
    outputs(6725) <= not (a xor b);
    outputs(6726) <= not (a xor b);
    outputs(6727) <= b and not a;
    outputs(6728) <= b and not a;
    outputs(6729) <= not (a xor b);
    outputs(6730) <= a;
    outputs(6731) <= a and not b;
    outputs(6732) <= a xor b;
    outputs(6733) <= not (a xor b);
    outputs(6734) <= b;
    outputs(6735) <= not a;
    outputs(6736) <= not a or b;
    outputs(6737) <= not a;
    outputs(6738) <= not (a xor b);
    outputs(6739) <= a xor b;
    outputs(6740) <= b and not a;
    outputs(6741) <= a and b;
    outputs(6742) <= b and not a;
    outputs(6743) <= not a;
    outputs(6744) <= not b;
    outputs(6745) <= b;
    outputs(6746) <= not b;
    outputs(6747) <= not a;
    outputs(6748) <= '0';
    outputs(6749) <= not (a and b);
    outputs(6750) <= not b;
    outputs(6751) <= not b;
    outputs(6752) <= not (a or b);
    outputs(6753) <= b and not a;
    outputs(6754) <= not (a xor b);
    outputs(6755) <= not (a or b);
    outputs(6756) <= not (a xor b);
    outputs(6757) <= a;
    outputs(6758) <= a xor b;
    outputs(6759) <= a or b;
    outputs(6760) <= a and not b;
    outputs(6761) <= not b or a;
    outputs(6762) <= not b;
    outputs(6763) <= not a;
    outputs(6764) <= not b;
    outputs(6765) <= a;
    outputs(6766) <= not (a xor b);
    outputs(6767) <= a or b;
    outputs(6768) <= not (a and b);
    outputs(6769) <= not (a xor b);
    outputs(6770) <= not (a and b);
    outputs(6771) <= a and not b;
    outputs(6772) <= not a or b;
    outputs(6773) <= b and not a;
    outputs(6774) <= not b;
    outputs(6775) <= a xor b;
    outputs(6776) <= not a or b;
    outputs(6777) <= a and b;
    outputs(6778) <= not b;
    outputs(6779) <= b and not a;
    outputs(6780) <= not (a xor b);
    outputs(6781) <= not b;
    outputs(6782) <= a xor b;
    outputs(6783) <= a xor b;
    outputs(6784) <= b;
    outputs(6785) <= not b;
    outputs(6786) <= a xor b;
    outputs(6787) <= not (a or b);
    outputs(6788) <= a xor b;
    outputs(6789) <= a and b;
    outputs(6790) <= a;
    outputs(6791) <= a xor b;
    outputs(6792) <= not (a or b);
    outputs(6793) <= not a or b;
    outputs(6794) <= b;
    outputs(6795) <= not (a xor b);
    outputs(6796) <= not a;
    outputs(6797) <= not b;
    outputs(6798) <= not (a and b);
    outputs(6799) <= a and not b;
    outputs(6800) <= a;
    outputs(6801) <= a or b;
    outputs(6802) <= not b;
    outputs(6803) <= a or b;
    outputs(6804) <= not b;
    outputs(6805) <= a;
    outputs(6806) <= not (a and b);
    outputs(6807) <= not (a xor b);
    outputs(6808) <= b;
    outputs(6809) <= a;
    outputs(6810) <= b and not a;
    outputs(6811) <= not (a xor b);
    outputs(6812) <= a and not b;
    outputs(6813) <= b;
    outputs(6814) <= not b;
    outputs(6815) <= a xor b;
    outputs(6816) <= not b;
    outputs(6817) <= a xor b;
    outputs(6818) <= not a or b;
    outputs(6819) <= a xor b;
    outputs(6820) <= a and b;
    outputs(6821) <= b and not a;
    outputs(6822) <= a;
    outputs(6823) <= not (a xor b);
    outputs(6824) <= not (a xor b);
    outputs(6825) <= a xor b;
    outputs(6826) <= not b;
    outputs(6827) <= not b;
    outputs(6828) <= a;
    outputs(6829) <= a or b;
    outputs(6830) <= a xor b;
    outputs(6831) <= a xor b;
    outputs(6832) <= not b;
    outputs(6833) <= not a;
    outputs(6834) <= not (a xor b);
    outputs(6835) <= b;
    outputs(6836) <= b and not a;
    outputs(6837) <= not b;
    outputs(6838) <= b;
    outputs(6839) <= not b or a;
    outputs(6840) <= a;
    outputs(6841) <= not b;
    outputs(6842) <= a;
    outputs(6843) <= not b;
    outputs(6844) <= not b;
    outputs(6845) <= b and not a;
    outputs(6846) <= not b;
    outputs(6847) <= not (a or b);
    outputs(6848) <= a;
    outputs(6849) <= b and not a;
    outputs(6850) <= b;
    outputs(6851) <= not (a xor b);
    outputs(6852) <= not b;
    outputs(6853) <= a and not b;
    outputs(6854) <= b;
    outputs(6855) <= not b;
    outputs(6856) <= b and not a;
    outputs(6857) <= a xor b;
    outputs(6858) <= not b;
    outputs(6859) <= a;
    outputs(6860) <= not a;
    outputs(6861) <= a;
    outputs(6862) <= not a or b;
    outputs(6863) <= b;
    outputs(6864) <= not b;
    outputs(6865) <= a;
    outputs(6866) <= a xor b;
    outputs(6867) <= a;
    outputs(6868) <= b;
    outputs(6869) <= a and not b;
    outputs(6870) <= a xor b;
    outputs(6871) <= a;
    outputs(6872) <= a and b;
    outputs(6873) <= not (a and b);
    outputs(6874) <= a;
    outputs(6875) <= not (a or b);
    outputs(6876) <= a and not b;
    outputs(6877) <= a;
    outputs(6878) <= not (a or b);
    outputs(6879) <= not a;
    outputs(6880) <= not (a or b);
    outputs(6881) <= not b;
    outputs(6882) <= not (a or b);
    outputs(6883) <= b;
    outputs(6884) <= not a or b;
    outputs(6885) <= a xor b;
    outputs(6886) <= a and not b;
    outputs(6887) <= not a;
    outputs(6888) <= a;
    outputs(6889) <= not b;
    outputs(6890) <= a or b;
    outputs(6891) <= b;
    outputs(6892) <= b;
    outputs(6893) <= not (a xor b);
    outputs(6894) <= not b;
    outputs(6895) <= not (a and b);
    outputs(6896) <= a;
    outputs(6897) <= a xor b;
    outputs(6898) <= not a or b;
    outputs(6899) <= a and b;
    outputs(6900) <= a xor b;
    outputs(6901) <= b and not a;
    outputs(6902) <= not b;
    outputs(6903) <= not (a or b);
    outputs(6904) <= b and not a;
    outputs(6905) <= a and not b;
    outputs(6906) <= not a;
    outputs(6907) <= not a;
    outputs(6908) <= a xor b;
    outputs(6909) <= not (a or b);
    outputs(6910) <= not b;
    outputs(6911) <= not (a xor b);
    outputs(6912) <= a;
    outputs(6913) <= a;
    outputs(6914) <= a and b;
    outputs(6915) <= a xor b;
    outputs(6916) <= b and not a;
    outputs(6917) <= not (a xor b);
    outputs(6918) <= not (a or b);
    outputs(6919) <= a xor b;
    outputs(6920) <= not a or b;
    outputs(6921) <= a and not b;
    outputs(6922) <= not a;
    outputs(6923) <= not (a xor b);
    outputs(6924) <= not (a xor b);
    outputs(6925) <= not (a xor b);
    outputs(6926) <= a xor b;
    outputs(6927) <= a and b;
    outputs(6928) <= b and not a;
    outputs(6929) <= not a;
    outputs(6930) <= not (a xor b);
    outputs(6931) <= not b;
    outputs(6932) <= not (a and b);
    outputs(6933) <= not b or a;
    outputs(6934) <= not a;
    outputs(6935) <= a and b;
    outputs(6936) <= a;
    outputs(6937) <= a;
    outputs(6938) <= b;
    outputs(6939) <= not b;
    outputs(6940) <= a and b;
    outputs(6941) <= b and not a;
    outputs(6942) <= b and not a;
    outputs(6943) <= a and b;
    outputs(6944) <= a and not b;
    outputs(6945) <= not (a and b);
    outputs(6946) <= a;
    outputs(6947) <= b;
    outputs(6948) <= b;
    outputs(6949) <= not (a xor b);
    outputs(6950) <= a and not b;
    outputs(6951) <= not (a or b);
    outputs(6952) <= not b;
    outputs(6953) <= not b;
    outputs(6954) <= a;
    outputs(6955) <= not (a xor b);
    outputs(6956) <= b;
    outputs(6957) <= b and not a;
    outputs(6958) <= a xor b;
    outputs(6959) <= a;
    outputs(6960) <= b;
    outputs(6961) <= a;
    outputs(6962) <= not (a xor b);
    outputs(6963) <= not (a or b);
    outputs(6964) <= a and b;
    outputs(6965) <= not (a xor b);
    outputs(6966) <= not b;
    outputs(6967) <= not a;
    outputs(6968) <= not b;
    outputs(6969) <= not a;
    outputs(6970) <= not a;
    outputs(6971) <= not b;
    outputs(6972) <= a and b;
    outputs(6973) <= not b or a;
    outputs(6974) <= a;
    outputs(6975) <= a and b;
    outputs(6976) <= b;
    outputs(6977) <= not a;
    outputs(6978) <= not b or a;
    outputs(6979) <= a and not b;
    outputs(6980) <= not a or b;
    outputs(6981) <= not (a and b);
    outputs(6982) <= not b or a;
    outputs(6983) <= not a;
    outputs(6984) <= not b or a;
    outputs(6985) <= b;
    outputs(6986) <= not (a xor b);
    outputs(6987) <= b and not a;
    outputs(6988) <= not (a and b);
    outputs(6989) <= a;
    outputs(6990) <= not (a xor b);
    outputs(6991) <= a or b;
    outputs(6992) <= b;
    outputs(6993) <= a xor b;
    outputs(6994) <= a;
    outputs(6995) <= not b;
    outputs(6996) <= a xor b;
    outputs(6997) <= a;
    outputs(6998) <= a xor b;
    outputs(6999) <= a xor b;
    outputs(7000) <= b and not a;
    outputs(7001) <= not (a xor b);
    outputs(7002) <= a;
    outputs(7003) <= not b;
    outputs(7004) <= not b;
    outputs(7005) <= not a;
    outputs(7006) <= not (a xor b);
    outputs(7007) <= not b;
    outputs(7008) <= not (a xor b);
    outputs(7009) <= a xor b;
    outputs(7010) <= not a;
    outputs(7011) <= not (a xor b);
    outputs(7012) <= not (a and b);
    outputs(7013) <= a xor b;
    outputs(7014) <= b;
    outputs(7015) <= not b;
    outputs(7016) <= not a;
    outputs(7017) <= a and b;
    outputs(7018) <= a;
    outputs(7019) <= not b;
    outputs(7020) <= a xor b;
    outputs(7021) <= not (a or b);
    outputs(7022) <= a;
    outputs(7023) <= a;
    outputs(7024) <= a;
    outputs(7025) <= not a;
    outputs(7026) <= not (a xor b);
    outputs(7027) <= a xor b;
    outputs(7028) <= b;
    outputs(7029) <= not b;
    outputs(7030) <= a xor b;
    outputs(7031) <= not b;
    outputs(7032) <= a xor b;
    outputs(7033) <= not (a xor b);
    outputs(7034) <= b;
    outputs(7035) <= b;
    outputs(7036) <= not (a and b);
    outputs(7037) <= b;
    outputs(7038) <= b and not a;
    outputs(7039) <= not (a xor b);
    outputs(7040) <= not b;
    outputs(7041) <= a and b;
    outputs(7042) <= a xor b;
    outputs(7043) <= not b or a;
    outputs(7044) <= b;
    outputs(7045) <= not b or a;
    outputs(7046) <= not (a xor b);
    outputs(7047) <= a or b;
    outputs(7048) <= a xor b;
    outputs(7049) <= not a;
    outputs(7050) <= a xor b;
    outputs(7051) <= not b or a;
    outputs(7052) <= a;
    outputs(7053) <= not (a and b);
    outputs(7054) <= not (a xor b);
    outputs(7055) <= a and b;
    outputs(7056) <= not b;
    outputs(7057) <= not (a xor b);
    outputs(7058) <= not (a xor b);
    outputs(7059) <= a xor b;
    outputs(7060) <= a xor b;
    outputs(7061) <= b;
    outputs(7062) <= not (a or b);
    outputs(7063) <= not a;
    outputs(7064) <= not a;
    outputs(7065) <= not a or b;
    outputs(7066) <= not b;
    outputs(7067) <= a xor b;
    outputs(7068) <= b;
    outputs(7069) <= a xor b;
    outputs(7070) <= a;
    outputs(7071) <= a xor b;
    outputs(7072) <= a xor b;
    outputs(7073) <= not a;
    outputs(7074) <= not (a xor b);
    outputs(7075) <= a xor b;
    outputs(7076) <= not a;
    outputs(7077) <= a and not b;
    outputs(7078) <= a and b;
    outputs(7079) <= a;
    outputs(7080) <= not (a or b);
    outputs(7081) <= not b;
    outputs(7082) <= a xor b;
    outputs(7083) <= a;
    outputs(7084) <= not b;
    outputs(7085) <= b and not a;
    outputs(7086) <= a or b;
    outputs(7087) <= not b;
    outputs(7088) <= not a;
    outputs(7089) <= not (a xor b);
    outputs(7090) <= not a;
    outputs(7091) <= not (a and b);
    outputs(7092) <= a and b;
    outputs(7093) <= a and not b;
    outputs(7094) <= not b or a;
    outputs(7095) <= not (a xor b);
    outputs(7096) <= not (a or b);
    outputs(7097) <= b and not a;
    outputs(7098) <= not (a xor b);
    outputs(7099) <= b and not a;
    outputs(7100) <= not (a and b);
    outputs(7101) <= b;
    outputs(7102) <= not (a xor b);
    outputs(7103) <= a or b;
    outputs(7104) <= b;
    outputs(7105) <= a and not b;
    outputs(7106) <= not b;
    outputs(7107) <= a and not b;
    outputs(7108) <= not (a or b);
    outputs(7109) <= a;
    outputs(7110) <= not (a xor b);
    outputs(7111) <= b;
    outputs(7112) <= a xor b;
    outputs(7113) <= a;
    outputs(7114) <= a xor b;
    outputs(7115) <= a xor b;
    outputs(7116) <= a and not b;
    outputs(7117) <= a and b;
    outputs(7118) <= not b;
    outputs(7119) <= not a or b;
    outputs(7120) <= a;
    outputs(7121) <= not b;
    outputs(7122) <= a and not b;
    outputs(7123) <= a and b;
    outputs(7124) <= not (a xor b);
    outputs(7125) <= a xor b;
    outputs(7126) <= not (a and b);
    outputs(7127) <= not a;
    outputs(7128) <= not b or a;
    outputs(7129) <= b;
    outputs(7130) <= not a;
    outputs(7131) <= not (a xor b);
    outputs(7132) <= b and not a;
    outputs(7133) <= a or b;
    outputs(7134) <= b;
    outputs(7135) <= not b;
    outputs(7136) <= a and not b;
    outputs(7137) <= not a;
    outputs(7138) <= not b;
    outputs(7139) <= not (a xor b);
    outputs(7140) <= not (a or b);
    outputs(7141) <= a or b;
    outputs(7142) <= b;
    outputs(7143) <= a and b;
    outputs(7144) <= not b or a;
    outputs(7145) <= not a;
    outputs(7146) <= a and not b;
    outputs(7147) <= not a or b;
    outputs(7148) <= not (a and b);
    outputs(7149) <= not (a xor b);
    outputs(7150) <= b;
    outputs(7151) <= b;
    outputs(7152) <= a xor b;
    outputs(7153) <= a;
    outputs(7154) <= not b;
    outputs(7155) <= a;
    outputs(7156) <= not a;
    outputs(7157) <= a xor b;
    outputs(7158) <= not (a xor b);
    outputs(7159) <= a xor b;
    outputs(7160) <= b;
    outputs(7161) <= b;
    outputs(7162) <= b;
    outputs(7163) <= not a;
    outputs(7164) <= not (a xor b);
    outputs(7165) <= a;
    outputs(7166) <= not (a xor b);
    outputs(7167) <= not a;
    outputs(7168) <= a xor b;
    outputs(7169) <= a xor b;
    outputs(7170) <= not b or a;
    outputs(7171) <= not a;
    outputs(7172) <= b and not a;
    outputs(7173) <= not b;
    outputs(7174) <= a and not b;
    outputs(7175) <= not b;
    outputs(7176) <= not (a and b);
    outputs(7177) <= a xor b;
    outputs(7178) <= not a;
    outputs(7179) <= a and not b;
    outputs(7180) <= b;
    outputs(7181) <= b and not a;
    outputs(7182) <= a xor b;
    outputs(7183) <= b and not a;
    outputs(7184) <= b;
    outputs(7185) <= not a;
    outputs(7186) <= not a;
    outputs(7187) <= a;
    outputs(7188) <= b;
    outputs(7189) <= a and b;
    outputs(7190) <= b and not a;
    outputs(7191) <= not a;
    outputs(7192) <= b and not a;
    outputs(7193) <= not a;
    outputs(7194) <= not (a or b);
    outputs(7195) <= not a;
    outputs(7196) <= not (a xor b);
    outputs(7197) <= a and not b;
    outputs(7198) <= not a;
    outputs(7199) <= not (a and b);
    outputs(7200) <= not (a or b);
    outputs(7201) <= a or b;
    outputs(7202) <= not b;
    outputs(7203) <= not a;
    outputs(7204) <= b;
    outputs(7205) <= a and b;
    outputs(7206) <= not a;
    outputs(7207) <= not b;
    outputs(7208) <= a or b;
    outputs(7209) <= not (a xor b);
    outputs(7210) <= a;
    outputs(7211) <= not (a xor b);
    outputs(7212) <= a and b;
    outputs(7213) <= b and not a;
    outputs(7214) <= a or b;
    outputs(7215) <= b;
    outputs(7216) <= b and not a;
    outputs(7217) <= b;
    outputs(7218) <= b;
    outputs(7219) <= not (a xor b);
    outputs(7220) <= not (a or b);
    outputs(7221) <= b;
    outputs(7222) <= a xor b;
    outputs(7223) <= a xor b;
    outputs(7224) <= not b;
    outputs(7225) <= not a;
    outputs(7226) <= not b;
    outputs(7227) <= not a;
    outputs(7228) <= a and not b;
    outputs(7229) <= not (a xor b);
    outputs(7230) <= not (a and b);
    outputs(7231) <= b and not a;
    outputs(7232) <= a and b;
    outputs(7233) <= a and b;
    outputs(7234) <= not (a or b);
    outputs(7235) <= a and b;
    outputs(7236) <= a;
    outputs(7237) <= a xor b;
    outputs(7238) <= not b or a;
    outputs(7239) <= b;
    outputs(7240) <= not (a or b);
    outputs(7241) <= a xor b;
    outputs(7242) <= a xor b;
    outputs(7243) <= a;
    outputs(7244) <= not (a xor b);
    outputs(7245) <= a;
    outputs(7246) <= not (a xor b);
    outputs(7247) <= a and b;
    outputs(7248) <= b;
    outputs(7249) <= not a;
    outputs(7250) <= b and not a;
    outputs(7251) <= not (a xor b);
    outputs(7252) <= b;
    outputs(7253) <= not a;
    outputs(7254) <= a;
    outputs(7255) <= a;
    outputs(7256) <= not b;
    outputs(7257) <= not (a xor b);
    outputs(7258) <= not (a xor b);
    outputs(7259) <= not b;
    outputs(7260) <= not (a xor b);
    outputs(7261) <= a xor b;
    outputs(7262) <= b;
    outputs(7263) <= not a or b;
    outputs(7264) <= a and not b;
    outputs(7265) <= not b;
    outputs(7266) <= not (a or b);
    outputs(7267) <= b;
    outputs(7268) <= not b;
    outputs(7269) <= not (a xor b);
    outputs(7270) <= b;
    outputs(7271) <= not a or b;
    outputs(7272) <= not a;
    outputs(7273) <= a and b;
    outputs(7274) <= not (a xor b);
    outputs(7275) <= not b;
    outputs(7276) <= a;
    outputs(7277) <= a and b;
    outputs(7278) <= not (a xor b);
    outputs(7279) <= a and b;
    outputs(7280) <= not (a xor b);
    outputs(7281) <= not b;
    outputs(7282) <= not (a or b);
    outputs(7283) <= not (a xor b);
    outputs(7284) <= not b;
    outputs(7285) <= not a;
    outputs(7286) <= a;
    outputs(7287) <= a and b;
    outputs(7288) <= not (a xor b);
    outputs(7289) <= not b;
    outputs(7290) <= a;
    outputs(7291) <= not b or a;
    outputs(7292) <= not b or a;
    outputs(7293) <= a xor b;
    outputs(7294) <= a xor b;
    outputs(7295) <= not (a xor b);
    outputs(7296) <= not (a and b);
    outputs(7297) <= a and not b;
    outputs(7298) <= a and b;
    outputs(7299) <= not a;
    outputs(7300) <= not b;
    outputs(7301) <= not a;
    outputs(7302) <= not a;
    outputs(7303) <= b;
    outputs(7304) <= a or b;
    outputs(7305) <= not b;
    outputs(7306) <= not (a xor b);
    outputs(7307) <= a;
    outputs(7308) <= b and not a;
    outputs(7309) <= not a;
    outputs(7310) <= b and not a;
    outputs(7311) <= not (a or b);
    outputs(7312) <= b and not a;
    outputs(7313) <= not a;
    outputs(7314) <= a xor b;
    outputs(7315) <= not b;
    outputs(7316) <= a xor b;
    outputs(7317) <= not b;
    outputs(7318) <= not a;
    outputs(7319) <= not a;
    outputs(7320) <= not (a xor b);
    outputs(7321) <= b;
    outputs(7322) <= b and not a;
    outputs(7323) <= a and not b;
    outputs(7324) <= a xor b;
    outputs(7325) <= a;
    outputs(7326) <= not (a xor b);
    outputs(7327) <= not b;
    outputs(7328) <= a and b;
    outputs(7329) <= a;
    outputs(7330) <= not (a xor b);
    outputs(7331) <= a or b;
    outputs(7332) <= a xor b;
    outputs(7333) <= not (a xor b);
    outputs(7334) <= not a;
    outputs(7335) <= not b;
    outputs(7336) <= a xor b;
    outputs(7337) <= a;
    outputs(7338) <= not b or a;
    outputs(7339) <= not b;
    outputs(7340) <= not a;
    outputs(7341) <= not a;
    outputs(7342) <= not a;
    outputs(7343) <= not (a or b);
    outputs(7344) <= a and not b;
    outputs(7345) <= a and not b;
    outputs(7346) <= a and b;
    outputs(7347) <= b;
    outputs(7348) <= a xor b;
    outputs(7349) <= not b;
    outputs(7350) <= not a;
    outputs(7351) <= a xor b;
    outputs(7352) <= a;
    outputs(7353) <= a xor b;
    outputs(7354) <= a xor b;
    outputs(7355) <= a;
    outputs(7356) <= a and not b;
    outputs(7357) <= not b;
    outputs(7358) <= a;
    outputs(7359) <= not b or a;
    outputs(7360) <= b;
    outputs(7361) <= not a;
    outputs(7362) <= a;
    outputs(7363) <= b and not a;
    outputs(7364) <= not (a xor b);
    outputs(7365) <= not (a and b);
    outputs(7366) <= not b;
    outputs(7367) <= a and b;
    outputs(7368) <= not (a and b);
    outputs(7369) <= a;
    outputs(7370) <= a;
    outputs(7371) <= not a or b;
    outputs(7372) <= a xor b;
    outputs(7373) <= a;
    outputs(7374) <= a and not b;
    outputs(7375) <= not a;
    outputs(7376) <= not (a xor b);
    outputs(7377) <= b and not a;
    outputs(7378) <= not (a or b);
    outputs(7379) <= a and b;
    outputs(7380) <= b;
    outputs(7381) <= not a;
    outputs(7382) <= b and not a;
    outputs(7383) <= a xor b;
    outputs(7384) <= a;
    outputs(7385) <= not a or b;
    outputs(7386) <= b;
    outputs(7387) <= a;
    outputs(7388) <= not (a or b);
    outputs(7389) <= a and not b;
    outputs(7390) <= b;
    outputs(7391) <= b and not a;
    outputs(7392) <= a and not b;
    outputs(7393) <= a;
    outputs(7394) <= a xor b;
    outputs(7395) <= a;
    outputs(7396) <= not b;
    outputs(7397) <= not b;
    outputs(7398) <= a and b;
    outputs(7399) <= not a or b;
    outputs(7400) <= not a;
    outputs(7401) <= not b;
    outputs(7402) <= a;
    outputs(7403) <= not b;
    outputs(7404) <= not a or b;
    outputs(7405) <= a or b;
    outputs(7406) <= not b;
    outputs(7407) <= a and not b;
    outputs(7408) <= not b;
    outputs(7409) <= a xor b;
    outputs(7410) <= b and not a;
    outputs(7411) <= not b;
    outputs(7412) <= a and not b;
    outputs(7413) <= not (a xor b);
    outputs(7414) <= not a;
    outputs(7415) <= not (a and b);
    outputs(7416) <= a xor b;
    outputs(7417) <= not (a and b);
    outputs(7418) <= not (a xor b);
    outputs(7419) <= a and b;
    outputs(7420) <= a;
    outputs(7421) <= b and not a;
    outputs(7422) <= not b;
    outputs(7423) <= not b;
    outputs(7424) <= a xor b;
    outputs(7425) <= a xor b;
    outputs(7426) <= a xor b;
    outputs(7427) <= not (a or b);
    outputs(7428) <= b and not a;
    outputs(7429) <= not a;
    outputs(7430) <= a or b;
    outputs(7431) <= not b;
    outputs(7432) <= b and not a;
    outputs(7433) <= b and not a;
    outputs(7434) <= not b;
    outputs(7435) <= a;
    outputs(7436) <= a;
    outputs(7437) <= a;
    outputs(7438) <= b and not a;
    outputs(7439) <= a xor b;
    outputs(7440) <= a and not b;
    outputs(7441) <= not b;
    outputs(7442) <= b;
    outputs(7443) <= b;
    outputs(7444) <= not (a or b);
    outputs(7445) <= not a;
    outputs(7446) <= not (a xor b);
    outputs(7447) <= not (a and b);
    outputs(7448) <= not (a and b);
    outputs(7449) <= not b;
    outputs(7450) <= a and not b;
    outputs(7451) <= a and b;
    outputs(7452) <= a;
    outputs(7453) <= not (a xor b);
    outputs(7454) <= a and b;
    outputs(7455) <= not (a xor b);
    outputs(7456) <= not b or a;
    outputs(7457) <= a and not b;
    outputs(7458) <= not b;
    outputs(7459) <= b and not a;
    outputs(7460) <= not (a and b);
    outputs(7461) <= not b;
    outputs(7462) <= a xor b;
    outputs(7463) <= a;
    outputs(7464) <= a and not b;
    outputs(7465) <= not b;
    outputs(7466) <= not a;
    outputs(7467) <= b;
    outputs(7468) <= not (a and b);
    outputs(7469) <= not (a xor b);
    outputs(7470) <= not (a and b);
    outputs(7471) <= b and not a;
    outputs(7472) <= b;
    outputs(7473) <= not (a or b);
    outputs(7474) <= not b;
    outputs(7475) <= b and not a;
    outputs(7476) <= not (a xor b);
    outputs(7477) <= a;
    outputs(7478) <= not b;
    outputs(7479) <= not b;
    outputs(7480) <= not (a xor b);
    outputs(7481) <= not (a or b);
    outputs(7482) <= a;
    outputs(7483) <= a xor b;
    outputs(7484) <= not b;
    outputs(7485) <= not a or b;
    outputs(7486) <= not (a xor b);
    outputs(7487) <= a and b;
    outputs(7488) <= a;
    outputs(7489) <= not (a xor b);
    outputs(7490) <= b and not a;
    outputs(7491) <= not (a xor b);
    outputs(7492) <= a;
    outputs(7493) <= not (a xor b);
    outputs(7494) <= b;
    outputs(7495) <= not (a xor b);
    outputs(7496) <= not (a or b);
    outputs(7497) <= not (a xor b);
    outputs(7498) <= not a;
    outputs(7499) <= not b or a;
    outputs(7500) <= not b;
    outputs(7501) <= not (a xor b);
    outputs(7502) <= a xor b;
    outputs(7503) <= a;
    outputs(7504) <= not b;
    outputs(7505) <= not a or b;
    outputs(7506) <= not (a xor b);
    outputs(7507) <= not b or a;
    outputs(7508) <= not b;
    outputs(7509) <= not a;
    outputs(7510) <= not (a or b);
    outputs(7511) <= not (a xor b);
    outputs(7512) <= b;
    outputs(7513) <= not b;
    outputs(7514) <= a xor b;
    outputs(7515) <= b and not a;
    outputs(7516) <= not a or b;
    outputs(7517) <= a xor b;
    outputs(7518) <= a and b;
    outputs(7519) <= a and b;
    outputs(7520) <= a and b;
    outputs(7521) <= a and b;
    outputs(7522) <= not (a or b);
    outputs(7523) <= not a;
    outputs(7524) <= not a;
    outputs(7525) <= not (a xor b);
    outputs(7526) <= not b;
    outputs(7527) <= b;
    outputs(7528) <= a xor b;
    outputs(7529) <= a and not b;
    outputs(7530) <= not (a xor b);
    outputs(7531) <= not (a and b);
    outputs(7532) <= b and not a;
    outputs(7533) <= a and b;
    outputs(7534) <= not b or a;
    outputs(7535) <= a and not b;
    outputs(7536) <= not (a xor b);
    outputs(7537) <= not (a xor b);
    outputs(7538) <= a and not b;
    outputs(7539) <= b and not a;
    outputs(7540) <= not b;
    outputs(7541) <= not (a xor b);
    outputs(7542) <= not a;
    outputs(7543) <= not (a xor b);
    outputs(7544) <= b and not a;
    outputs(7545) <= b;
    outputs(7546) <= b and not a;
    outputs(7547) <= not (a or b);
    outputs(7548) <= not (a and b);
    outputs(7549) <= a and not b;
    outputs(7550) <= a or b;
    outputs(7551) <= b and not a;
    outputs(7552) <= a and not b;
    outputs(7553) <= b;
    outputs(7554) <= a and b;
    outputs(7555) <= not (a or b);
    outputs(7556) <= a and not b;
    outputs(7557) <= a and b;
    outputs(7558) <= a xor b;
    outputs(7559) <= not (a xor b);
    outputs(7560) <= not b;
    outputs(7561) <= not b;
    outputs(7562) <= b;
    outputs(7563) <= not (a or b);
    outputs(7564) <= a and b;
    outputs(7565) <= a;
    outputs(7566) <= b and not a;
    outputs(7567) <= b and not a;
    outputs(7568) <= not a;
    outputs(7569) <= not (a or b);
    outputs(7570) <= b;
    outputs(7571) <= a and b;
    outputs(7572) <= not a;
    outputs(7573) <= a and not b;
    outputs(7574) <= not (a and b);
    outputs(7575) <= a and not b;
    outputs(7576) <= b and not a;
    outputs(7577) <= a and b;
    outputs(7578) <= '0';
    outputs(7579) <= a;
    outputs(7580) <= a;
    outputs(7581) <= a xor b;
    outputs(7582) <= b;
    outputs(7583) <= a and not b;
    outputs(7584) <= a and not b;
    outputs(7585) <= not (a and b);
    outputs(7586) <= b and not a;
    outputs(7587) <= a or b;
    outputs(7588) <= a;
    outputs(7589) <= not (a xor b);
    outputs(7590) <= a xor b;
    outputs(7591) <= not (a xor b);
    outputs(7592) <= not (a or b);
    outputs(7593) <= a xor b;
    outputs(7594) <= b and not a;
    outputs(7595) <= not (a xor b);
    outputs(7596) <= not b or a;
    outputs(7597) <= not a;
    outputs(7598) <= a and b;
    outputs(7599) <= b;
    outputs(7600) <= a and not b;
    outputs(7601) <= not (a or b);
    outputs(7602) <= b and not a;
    outputs(7603) <= b and not a;
    outputs(7604) <= not (a or b);
    outputs(7605) <= not a;
    outputs(7606) <= a and b;
    outputs(7607) <= a xor b;
    outputs(7608) <= not (a xor b);
    outputs(7609) <= a and not b;
    outputs(7610) <= not (a or b);
    outputs(7611) <= a;
    outputs(7612) <= not (a xor b);
    outputs(7613) <= a;
    outputs(7614) <= not a or b;
    outputs(7615) <= a xor b;
    outputs(7616) <= b;
    outputs(7617) <= b;
    outputs(7618) <= not (a xor b);
    outputs(7619) <= not (a xor b);
    outputs(7620) <= not (a or b);
    outputs(7621) <= b;
    outputs(7622) <= a or b;
    outputs(7623) <= a;
    outputs(7624) <= not a;
    outputs(7625) <= b and not a;
    outputs(7626) <= a and b;
    outputs(7627) <= not a or b;
    outputs(7628) <= a and b;
    outputs(7629) <= a and not b;
    outputs(7630) <= a and not b;
    outputs(7631) <= b and not a;
    outputs(7632) <= a xor b;
    outputs(7633) <= not (a or b);
    outputs(7634) <= not a;
    outputs(7635) <= a;
    outputs(7636) <= not a;
    outputs(7637) <= b and not a;
    outputs(7638) <= a;
    outputs(7639) <= a;
    outputs(7640) <= b;
    outputs(7641) <= not b;
    outputs(7642) <= not (a xor b);
    outputs(7643) <= b;
    outputs(7644) <= a;
    outputs(7645) <= not (a or b);
    outputs(7646) <= not a;
    outputs(7647) <= a xor b;
    outputs(7648) <= not (a xor b);
    outputs(7649) <= not a;
    outputs(7650) <= not a;
    outputs(7651) <= a xor b;
    outputs(7652) <= a;
    outputs(7653) <= not (a xor b);
    outputs(7654) <= b;
    outputs(7655) <= b and not a;
    outputs(7656) <= a xor b;
    outputs(7657) <= not (a or b);
    outputs(7658) <= not (a or b);
    outputs(7659) <= not b;
    outputs(7660) <= a xor b;
    outputs(7661) <= not (a and b);
    outputs(7662) <= not a;
    outputs(7663) <= a and b;
    outputs(7664) <= a;
    outputs(7665) <= a and not b;
    outputs(7666) <= not (a xor b);
    outputs(7667) <= a or b;
    outputs(7668) <= not (a or b);
    outputs(7669) <= not (a xor b);
    outputs(7670) <= not a;
    outputs(7671) <= not a or b;
    outputs(7672) <= not b;
    outputs(7673) <= a and b;
    outputs(7674) <= a and not b;
    outputs(7675) <= a xor b;
    outputs(7676) <= a;
    outputs(7677) <= a xor b;
    outputs(7678) <= a;
    outputs(7679) <= b;
    outputs(7680) <= not b or a;
    outputs(7681) <= a or b;
    outputs(7682) <= not a;
    outputs(7683) <= a;
    outputs(7684) <= not a;
    outputs(7685) <= not (a xor b);
    outputs(7686) <= a or b;
    outputs(7687) <= a and b;
    outputs(7688) <= a xor b;
    outputs(7689) <= not (a or b);
    outputs(7690) <= not (a or b);
    outputs(7691) <= not (a or b);
    outputs(7692) <= a xor b;
    outputs(7693) <= not b;
    outputs(7694) <= a xor b;
    outputs(7695) <= not (a xor b);
    outputs(7696) <= b;
    outputs(7697) <= not (a xor b);
    outputs(7698) <= not (a xor b);
    outputs(7699) <= not b;
    outputs(7700) <= a and not b;
    outputs(7701) <= a and not b;
    outputs(7702) <= a;
    outputs(7703) <= a xor b;
    outputs(7704) <= a xor b;
    outputs(7705) <= not b;
    outputs(7706) <= a and b;
    outputs(7707) <= not a;
    outputs(7708) <= b;
    outputs(7709) <= a;
    outputs(7710) <= not (a or b);
    outputs(7711) <= a;
    outputs(7712) <= not (a or b);
    outputs(7713) <= b;
    outputs(7714) <= not (a xor b);
    outputs(7715) <= a and b;
    outputs(7716) <= a;
    outputs(7717) <= a;
    outputs(7718) <= a xor b;
    outputs(7719) <= not a;
    outputs(7720) <= not a;
    outputs(7721) <= not b;
    outputs(7722) <= b;
    outputs(7723) <= a xor b;
    outputs(7724) <= b;
    outputs(7725) <= not a;
    outputs(7726) <= not (a xor b);
    outputs(7727) <= b and not a;
    outputs(7728) <= not a or b;
    outputs(7729) <= a and b;
    outputs(7730) <= not a or b;
    outputs(7731) <= not (a or b);
    outputs(7732) <= a;
    outputs(7733) <= a xor b;
    outputs(7734) <= not b;
    outputs(7735) <= not a;
    outputs(7736) <= a xor b;
    outputs(7737) <= a xor b;
    outputs(7738) <= not (a xor b);
    outputs(7739) <= b and not a;
    outputs(7740) <= a;
    outputs(7741) <= a xor b;
    outputs(7742) <= not b;
    outputs(7743) <= a;
    outputs(7744) <= a and b;
    outputs(7745) <= b;
    outputs(7746) <= b and not a;
    outputs(7747) <= b;
    outputs(7748) <= a and not b;
    outputs(7749) <= b;
    outputs(7750) <= not a;
    outputs(7751) <= a;
    outputs(7752) <= not b;
    outputs(7753) <= a xor b;
    outputs(7754) <= not (a and b);
    outputs(7755) <= a and not b;
    outputs(7756) <= not (a xor b);
    outputs(7757) <= not (a or b);
    outputs(7758) <= b and not a;
    outputs(7759) <= a xor b;
    outputs(7760) <= not b;
    outputs(7761) <= b and not a;
    outputs(7762) <= not (a xor b);
    outputs(7763) <= a and not b;
    outputs(7764) <= not (a xor b);
    outputs(7765) <= not (a xor b);
    outputs(7766) <= not a;
    outputs(7767) <= not b;
    outputs(7768) <= a;
    outputs(7769) <= not b;
    outputs(7770) <= not a;
    outputs(7771) <= b and not a;
    outputs(7772) <= a and not b;
    outputs(7773) <= b;
    outputs(7774) <= b;
    outputs(7775) <= a xor b;
    outputs(7776) <= not a;
    outputs(7777) <= a and b;
    outputs(7778) <= a xor b;
    outputs(7779) <= not b or a;
    outputs(7780) <= not a;
    outputs(7781) <= not (a xor b);
    outputs(7782) <= not (a xor b);
    outputs(7783) <= a xor b;
    outputs(7784) <= b and not a;
    outputs(7785) <= not a or b;
    outputs(7786) <= a xor b;
    outputs(7787) <= not b or a;
    outputs(7788) <= not (a xor b);
    outputs(7789) <= not (a xor b);
    outputs(7790) <= a or b;
    outputs(7791) <= b and not a;
    outputs(7792) <= not b;
    outputs(7793) <= b and not a;
    outputs(7794) <= a xor b;
    outputs(7795) <= not a;
    outputs(7796) <= not (a xor b);
    outputs(7797) <= b;
    outputs(7798) <= a or b;
    outputs(7799) <= not (a or b);
    outputs(7800) <= not a or b;
    outputs(7801) <= a and b;
    outputs(7802) <= a or b;
    outputs(7803) <= not b;
    outputs(7804) <= a and not b;
    outputs(7805) <= b;
    outputs(7806) <= not a;
    outputs(7807) <= not a;
    outputs(7808) <= not (a xor b);
    outputs(7809) <= b and not a;
    outputs(7810) <= a and not b;
    outputs(7811) <= a or b;
    outputs(7812) <= not b;
    outputs(7813) <= a and not b;
    outputs(7814) <= a;
    outputs(7815) <= not (a or b);
    outputs(7816) <= a and b;
    outputs(7817) <= not (a xor b);
    outputs(7818) <= a or b;
    outputs(7819) <= not a or b;
    outputs(7820) <= a xor b;
    outputs(7821) <= a xor b;
    outputs(7822) <= a xor b;
    outputs(7823) <= not (a xor b);
    outputs(7824) <= a or b;
    outputs(7825) <= not b or a;
    outputs(7826) <= not a;
    outputs(7827) <= a and not b;
    outputs(7828) <= not (a or b);
    outputs(7829) <= not a;
    outputs(7830) <= not (a or b);
    outputs(7831) <= not (a xor b);
    outputs(7832) <= a;
    outputs(7833) <= a xor b;
    outputs(7834) <= b and not a;
    outputs(7835) <= a xor b;
    outputs(7836) <= not a;
    outputs(7837) <= b and not a;
    outputs(7838) <= a xor b;
    outputs(7839) <= a and b;
    outputs(7840) <= not (a and b);
    outputs(7841) <= not (a xor b);
    outputs(7842) <= b and not a;
    outputs(7843) <= not (a or b);
    outputs(7844) <= a;
    outputs(7845) <= a xor b;
    outputs(7846) <= b;
    outputs(7847) <= not (a xor b);
    outputs(7848) <= not b;
    outputs(7849) <= not (a xor b);
    outputs(7850) <= b;
    outputs(7851) <= a;
    outputs(7852) <= a and b;
    outputs(7853) <= not b;
    outputs(7854) <= not a;
    outputs(7855) <= b;
    outputs(7856) <= a;
    outputs(7857) <= not (a xor b);
    outputs(7858) <= a and b;
    outputs(7859) <= a and not b;
    outputs(7860) <= not b;
    outputs(7861) <= not a;
    outputs(7862) <= not a or b;
    outputs(7863) <= a;
    outputs(7864) <= not (a or b);
    outputs(7865) <= b and not a;
    outputs(7866) <= not a;
    outputs(7867) <= not a or b;
    outputs(7868) <= not a or b;
    outputs(7869) <= a xor b;
    outputs(7870) <= b and not a;
    outputs(7871) <= not (a xor b);
    outputs(7872) <= b;
    outputs(7873) <= not a;
    outputs(7874) <= a and b;
    outputs(7875) <= not a or b;
    outputs(7876) <= a xor b;
    outputs(7877) <= b;
    outputs(7878) <= b;
    outputs(7879) <= not b;
    outputs(7880) <= a;
    outputs(7881) <= a xor b;
    outputs(7882) <= b and not a;
    outputs(7883) <= a and not b;
    outputs(7884) <= a and b;
    outputs(7885) <= not b or a;
    outputs(7886) <= not b;
    outputs(7887) <= a;
    outputs(7888) <= a xor b;
    outputs(7889) <= not b;
    outputs(7890) <= b;
    outputs(7891) <= not (a xor b);
    outputs(7892) <= a xor b;
    outputs(7893) <= b and not a;
    outputs(7894) <= not (a xor b);
    outputs(7895) <= a and b;
    outputs(7896) <= a and not b;
    outputs(7897) <= a and not b;
    outputs(7898) <= not b;
    outputs(7899) <= a;
    outputs(7900) <= not (a or b);
    outputs(7901) <= not (a or b);
    outputs(7902) <= not b;
    outputs(7903) <= b;
    outputs(7904) <= a xor b;
    outputs(7905) <= not (a or b);
    outputs(7906) <= not (a or b);
    outputs(7907) <= not (a or b);
    outputs(7908) <= a and b;
    outputs(7909) <= not a;
    outputs(7910) <= a and b;
    outputs(7911) <= a;
    outputs(7912) <= not (a xor b);
    outputs(7913) <= a or b;
    outputs(7914) <= b;
    outputs(7915) <= a and not b;
    outputs(7916) <= a and not b;
    outputs(7917) <= not (a or b);
    outputs(7918) <= a;
    outputs(7919) <= not (a xor b);
    outputs(7920) <= b;
    outputs(7921) <= b and not a;
    outputs(7922) <= b and not a;
    outputs(7923) <= not b;
    outputs(7924) <= a and not b;
    outputs(7925) <= not a or b;
    outputs(7926) <= a xor b;
    outputs(7927) <= b;
    outputs(7928) <= b;
    outputs(7929) <= b and not a;
    outputs(7930) <= not b or a;
    outputs(7931) <= a;
    outputs(7932) <= b;
    outputs(7933) <= a;
    outputs(7934) <= a xor b;
    outputs(7935) <= not a;
    outputs(7936) <= b and not a;
    outputs(7937) <= not b;
    outputs(7938) <= a and not b;
    outputs(7939) <= not b;
    outputs(7940) <= not b;
    outputs(7941) <= not b;
    outputs(7942) <= not a;
    outputs(7943) <= not (a or b);
    outputs(7944) <= b;
    outputs(7945) <= not a or b;
    outputs(7946) <= not a;
    outputs(7947) <= not (a or b);
    outputs(7948) <= a and not b;
    outputs(7949) <= a xor b;
    outputs(7950) <= not a;
    outputs(7951) <= not a;
    outputs(7952) <= a xor b;
    outputs(7953) <= b and not a;
    outputs(7954) <= not (a or b);
    outputs(7955) <= b;
    outputs(7956) <= not (a xor b);
    outputs(7957) <= a;
    outputs(7958) <= not b;
    outputs(7959) <= a and not b;
    outputs(7960) <= b and not a;
    outputs(7961) <= a and b;
    outputs(7962) <= not (a xor b);
    outputs(7963) <= not (a or b);
    outputs(7964) <= not b or a;
    outputs(7965) <= not a;
    outputs(7966) <= b and not a;
    outputs(7967) <= b and not a;
    outputs(7968) <= a and b;
    outputs(7969) <= not b;
    outputs(7970) <= not a or b;
    outputs(7971) <= a xor b;
    outputs(7972) <= not (a and b);
    outputs(7973) <= a;
    outputs(7974) <= a xor b;
    outputs(7975) <= b;
    outputs(7976) <= not (a or b);
    outputs(7977) <= a and b;
    outputs(7978) <= a xor b;
    outputs(7979) <= a;
    outputs(7980) <= not (a or b);
    outputs(7981) <= not (a xor b);
    outputs(7982) <= not (a xor b);
    outputs(7983) <= b;
    outputs(7984) <= a xor b;
    outputs(7985) <= a;
    outputs(7986) <= not a;
    outputs(7987) <= not a;
    outputs(7988) <= not (a or b);
    outputs(7989) <= a and not b;
    outputs(7990) <= a;
    outputs(7991) <= not (a or b);
    outputs(7992) <= not b;
    outputs(7993) <= a xor b;
    outputs(7994) <= not (a xor b);
    outputs(7995) <= not (a xor b);
    outputs(7996) <= a and b;
    outputs(7997) <= a;
    outputs(7998) <= b and not a;
    outputs(7999) <= not b;
    outputs(8000) <= a and b;
    outputs(8001) <= a and not b;
    outputs(8002) <= not (a xor b);
    outputs(8003) <= a and not b;
    outputs(8004) <= a or b;
    outputs(8005) <= not (a xor b);
    outputs(8006) <= not (a xor b);
    outputs(8007) <= not (a xor b);
    outputs(8008) <= not b or a;
    outputs(8009) <= not (a or b);
    outputs(8010) <= b;
    outputs(8011) <= not a;
    outputs(8012) <= not (a xor b);
    outputs(8013) <= not b;
    outputs(8014) <= b;
    outputs(8015) <= a and b;
    outputs(8016) <= not (a xor b);
    outputs(8017) <= a;
    outputs(8018) <= b;
    outputs(8019) <= a;
    outputs(8020) <= b;
    outputs(8021) <= not (a or b);
    outputs(8022) <= not b;
    outputs(8023) <= b;
    outputs(8024) <= not (a xor b);
    outputs(8025) <= a;
    outputs(8026) <= b;
    outputs(8027) <= not (a or b);
    outputs(8028) <= b and not a;
    outputs(8029) <= b and not a;
    outputs(8030) <= not b or a;
    outputs(8031) <= not b;
    outputs(8032) <= b and not a;
    outputs(8033) <= a and not b;
    outputs(8034) <= a and b;
    outputs(8035) <= b;
    outputs(8036) <= a and b;
    outputs(8037) <= not a;
    outputs(8038) <= not b;
    outputs(8039) <= a and not b;
    outputs(8040) <= a xor b;
    outputs(8041) <= a and not b;
    outputs(8042) <= a and not b;
    outputs(8043) <= not b or a;
    outputs(8044) <= not b;
    outputs(8045) <= a;
    outputs(8046) <= a and b;
    outputs(8047) <= a xor b;
    outputs(8048) <= a xor b;
    outputs(8049) <= not (a or b);
    outputs(8050) <= b;
    outputs(8051) <= not b;
    outputs(8052) <= not (a xor b);
    outputs(8053) <= not b;
    outputs(8054) <= a;
    outputs(8055) <= a;
    outputs(8056) <= a;
    outputs(8057) <= a;
    outputs(8058) <= not a or b;
    outputs(8059) <= not b or a;
    outputs(8060) <= b;
    outputs(8061) <= b and not a;
    outputs(8062) <= b;
    outputs(8063) <= not a;
    outputs(8064) <= a and b;
    outputs(8065) <= not (a xor b);
    outputs(8066) <= a and not b;
    outputs(8067) <= not b or a;
    outputs(8068) <= not a;
    outputs(8069) <= not (a xor b);
    outputs(8070) <= b;
    outputs(8071) <= a xor b;
    outputs(8072) <= a xor b;
    outputs(8073) <= b;
    outputs(8074) <= not a;
    outputs(8075) <= not a;
    outputs(8076) <= b and not a;
    outputs(8077) <= not b;
    outputs(8078) <= not a;
    outputs(8079) <= not b;
    outputs(8080) <= not (a or b);
    outputs(8081) <= not (a xor b);
    outputs(8082) <= not b;
    outputs(8083) <= a or b;
    outputs(8084) <= not a;
    outputs(8085) <= a and b;
    outputs(8086) <= a or b;
    outputs(8087) <= a xor b;
    outputs(8088) <= a and not b;
    outputs(8089) <= not (a or b);
    outputs(8090) <= not b;
    outputs(8091) <= not b;
    outputs(8092) <= not (a or b);
    outputs(8093) <= a or b;
    outputs(8094) <= not a or b;
    outputs(8095) <= b and not a;
    outputs(8096) <= a xor b;
    outputs(8097) <= not b;
    outputs(8098) <= not b;
    outputs(8099) <= not a;
    outputs(8100) <= b;
    outputs(8101) <= not a;
    outputs(8102) <= a;
    outputs(8103) <= a xor b;
    outputs(8104) <= a and not b;
    outputs(8105) <= b;
    outputs(8106) <= not (a xor b);
    outputs(8107) <= b;
    outputs(8108) <= not a;
    outputs(8109) <= b;
    outputs(8110) <= a xor b;
    outputs(8111) <= not b;
    outputs(8112) <= not a;
    outputs(8113) <= not a or b;
    outputs(8114) <= a xor b;
    outputs(8115) <= not (a or b);
    outputs(8116) <= not a;
    outputs(8117) <= not (a xor b);
    outputs(8118) <= not b;
    outputs(8119) <= a xor b;
    outputs(8120) <= a;
    outputs(8121) <= b;
    outputs(8122) <= b;
    outputs(8123) <= a;
    outputs(8124) <= not a;
    outputs(8125) <= a;
    outputs(8126) <= b;
    outputs(8127) <= not (a xor b);
    outputs(8128) <= not a;
    outputs(8129) <= not (a xor b);
    outputs(8130) <= a and b;
    outputs(8131) <= not (a or b);
    outputs(8132) <= b;
    outputs(8133) <= a and b;
    outputs(8134) <= not a;
    outputs(8135) <= not a;
    outputs(8136) <= not (a xor b);
    outputs(8137) <= not a;
    outputs(8138) <= not a;
    outputs(8139) <= not b;
    outputs(8140) <= b;
    outputs(8141) <= a xor b;
    outputs(8142) <= b;
    outputs(8143) <= a and not b;
    outputs(8144) <= a and not b;
    outputs(8145) <= not b;
    outputs(8146) <= b;
    outputs(8147) <= not (a xor b);
    outputs(8148) <= '0';
    outputs(8149) <= not (a xor b);
    outputs(8150) <= not (a or b);
    outputs(8151) <= b;
    outputs(8152) <= b and not a;
    outputs(8153) <= not (a xor b);
    outputs(8154) <= not a or b;
    outputs(8155) <= a xor b;
    outputs(8156) <= b;
    outputs(8157) <= b;
    outputs(8158) <= a and not b;
    outputs(8159) <= b and not a;
    outputs(8160) <= not (a xor b);
    outputs(8161) <= not (a xor b);
    outputs(8162) <= not a;
    outputs(8163) <= a xor b;
    outputs(8164) <= not (a xor b);
    outputs(8165) <= b;
    outputs(8166) <= not a;
    outputs(8167) <= a and b;
    outputs(8168) <= a xor b;
    outputs(8169) <= not (a or b);
    outputs(8170) <= a and not b;
    outputs(8171) <= b;
    outputs(8172) <= a or b;
    outputs(8173) <= a;
    outputs(8174) <= a and b;
    outputs(8175) <= not a;
    outputs(8176) <= not (a and b);
    outputs(8177) <= b;
    outputs(8178) <= not a;
    outputs(8179) <= b and not a;
    outputs(8180) <= b and not a;
    outputs(8181) <= not (a xor b);
    outputs(8182) <= not b;
    outputs(8183) <= a and not b;
    outputs(8184) <= a and b;
    outputs(8185) <= not a;
    outputs(8186) <= not b;
    outputs(8187) <= a xor b;
    outputs(8188) <= b;
    outputs(8189) <= a xor b;
    outputs(8190) <= a and b;
    outputs(8191) <= a;
    outputs(8192) <= b and not a;
    outputs(8193) <= not (a and b);
    outputs(8194) <= a;
    outputs(8195) <= a xor b;
    outputs(8196) <= a;
    outputs(8197) <= not b;
    outputs(8198) <= b;
    outputs(8199) <= a xor b;
    outputs(8200) <= a;
    outputs(8201) <= a and b;
    outputs(8202) <= not b or a;
    outputs(8203) <= not b;
    outputs(8204) <= b and not a;
    outputs(8205) <= a xor b;
    outputs(8206) <= not (a xor b);
    outputs(8207) <= not (a xor b);
    outputs(8208) <= a xor b;
    outputs(8209) <= b and not a;
    outputs(8210) <= not (a or b);
    outputs(8211) <= b;
    outputs(8212) <= not a;
    outputs(8213) <= not (a xor b);
    outputs(8214) <= a xor b;
    outputs(8215) <= b;
    outputs(8216) <= b;
    outputs(8217) <= not b;
    outputs(8218) <= not (a xor b);
    outputs(8219) <= a xor b;
    outputs(8220) <= b;
    outputs(8221) <= not (a xor b);
    outputs(8222) <= not (a or b);
    outputs(8223) <= not b or a;
    outputs(8224) <= a xor b;
    outputs(8225) <= b;
    outputs(8226) <= b;
    outputs(8227) <= a;
    outputs(8228) <= not a;
    outputs(8229) <= not (a xor b);
    outputs(8230) <= a;
    outputs(8231) <= not (a xor b);
    outputs(8232) <= not a;
    outputs(8233) <= a xor b;
    outputs(8234) <= not b;
    outputs(8235) <= not (a xor b);
    outputs(8236) <= a;
    outputs(8237) <= b;
    outputs(8238) <= a and not b;
    outputs(8239) <= not a;
    outputs(8240) <= not (a xor b);
    outputs(8241) <= b and not a;
    outputs(8242) <= not a or b;
    outputs(8243) <= a xor b;
    outputs(8244) <= a xor b;
    outputs(8245) <= not (a or b);
    outputs(8246) <= not (a or b);
    outputs(8247) <= a;
    outputs(8248) <= not b or a;
    outputs(8249) <= not (a or b);
    outputs(8250) <= not a or b;
    outputs(8251) <= not a or b;
    outputs(8252) <= b;
    outputs(8253) <= a or b;
    outputs(8254) <= a;
    outputs(8255) <= a xor b;
    outputs(8256) <= a;
    outputs(8257) <= a xor b;
    outputs(8258) <= not a;
    outputs(8259) <= a xor b;
    outputs(8260) <= not (a or b);
    outputs(8261) <= b;
    outputs(8262) <= a xor b;
    outputs(8263) <= not (a or b);
    outputs(8264) <= not (a xor b);
    outputs(8265) <= not a or b;
    outputs(8266) <= not (a xor b);
    outputs(8267) <= a and not b;
    outputs(8268) <= not b or a;
    outputs(8269) <= a xor b;
    outputs(8270) <= b;
    outputs(8271) <= not (a xor b);
    outputs(8272) <= a;
    outputs(8273) <= a or b;
    outputs(8274) <= a xor b;
    outputs(8275) <= a;
    outputs(8276) <= a;
    outputs(8277) <= a xor b;
    outputs(8278) <= a xor b;
    outputs(8279) <= a xor b;
    outputs(8280) <= not (a xor b);
    outputs(8281) <= b;
    outputs(8282) <= a xor b;
    outputs(8283) <= not a;
    outputs(8284) <= not b or a;
    outputs(8285) <= a xor b;
    outputs(8286) <= a;
    outputs(8287) <= not (a and b);
    outputs(8288) <= not (a xor b);
    outputs(8289) <= a xor b;
    outputs(8290) <= not (a xor b);
    outputs(8291) <= not a;
    outputs(8292) <= not (a and b);
    outputs(8293) <= not a;
    outputs(8294) <= a xor b;
    outputs(8295) <= not b;
    outputs(8296) <= a xor b;
    outputs(8297) <= not a;
    outputs(8298) <= not (a and b);
    outputs(8299) <= b;
    outputs(8300) <= not (a xor b);
    outputs(8301) <= a;
    outputs(8302) <= a xor b;
    outputs(8303) <= a;
    outputs(8304) <= b;
    outputs(8305) <= a and b;
    outputs(8306) <= b;
    outputs(8307) <= not (a xor b);
    outputs(8308) <= b;
    outputs(8309) <= a xor b;
    outputs(8310) <= not b or a;
    outputs(8311) <= a xor b;
    outputs(8312) <= not (a xor b);
    outputs(8313) <= b;
    outputs(8314) <= a xor b;
    outputs(8315) <= b;
    outputs(8316) <= b;
    outputs(8317) <= a;
    outputs(8318) <= b;
    outputs(8319) <= b and not a;
    outputs(8320) <= not b;
    outputs(8321) <= b;
    outputs(8322) <= a;
    outputs(8323) <= not a;
    outputs(8324) <= not b;
    outputs(8325) <= a or b;
    outputs(8326) <= not (a xor b);
    outputs(8327) <= a;
    outputs(8328) <= b;
    outputs(8329) <= a xor b;
    outputs(8330) <= not (a xor b);
    outputs(8331) <= not a or b;
    outputs(8332) <= not (a xor b);
    outputs(8333) <= not (a xor b);
    outputs(8334) <= not (a and b);
    outputs(8335) <= not a;
    outputs(8336) <= not b or a;
    outputs(8337) <= not b or a;
    outputs(8338) <= not (a xor b);
    outputs(8339) <= a xor b;
    outputs(8340) <= b;
    outputs(8341) <= not (a or b);
    outputs(8342) <= a xor b;
    outputs(8343) <= b;
    outputs(8344) <= a;
    outputs(8345) <= a and b;
    outputs(8346) <= a;
    outputs(8347) <= not b;
    outputs(8348) <= not (a xor b);
    outputs(8349) <= a xor b;
    outputs(8350) <= not b or a;
    outputs(8351) <= not a or b;
    outputs(8352) <= a;
    outputs(8353) <= not a;
    outputs(8354) <= b;
    outputs(8355) <= a and b;
    outputs(8356) <= a;
    outputs(8357) <= not (a or b);
    outputs(8358) <= a xor b;
    outputs(8359) <= not (a xor b);
    outputs(8360) <= not a;
    outputs(8361) <= a xor b;
    outputs(8362) <= not a;
    outputs(8363) <= a xor b;
    outputs(8364) <= a;
    outputs(8365) <= not a or b;
    outputs(8366) <= b;
    outputs(8367) <= not a;
    outputs(8368) <= not (a xor b);
    outputs(8369) <= not (a and b);
    outputs(8370) <= a;
    outputs(8371) <= not b;
    outputs(8372) <= not (a xor b);
    outputs(8373) <= not (a xor b);
    outputs(8374) <= not a;
    outputs(8375) <= not a or b;
    outputs(8376) <= a xor b;
    outputs(8377) <= b;
    outputs(8378) <= not b or a;
    outputs(8379) <= a or b;
    outputs(8380) <= a or b;
    outputs(8381) <= not a;
    outputs(8382) <= not (a xor b);
    outputs(8383) <= a or b;
    outputs(8384) <= a and b;
    outputs(8385) <= b;
    outputs(8386) <= b;
    outputs(8387) <= a and not b;
    outputs(8388) <= not b;
    outputs(8389) <= b;
    outputs(8390) <= b;
    outputs(8391) <= b;
    outputs(8392) <= not (a xor b);
    outputs(8393) <= a and b;
    outputs(8394) <= a xor b;
    outputs(8395) <= b;
    outputs(8396) <= not (a or b);
    outputs(8397) <= a and b;
    outputs(8398) <= not (a and b);
    outputs(8399) <= not (a or b);
    outputs(8400) <= not b;
    outputs(8401) <= not b or a;
    outputs(8402) <= not a;
    outputs(8403) <= a xor b;
    outputs(8404) <= b;
    outputs(8405) <= b;
    outputs(8406) <= not a;
    outputs(8407) <= not b or a;
    outputs(8408) <= a xor b;
    outputs(8409) <= not (a and b);
    outputs(8410) <= not (a and b);
    outputs(8411) <= b and not a;
    outputs(8412) <= not a;
    outputs(8413) <= a xor b;
    outputs(8414) <= not a;
    outputs(8415) <= not (a xor b);
    outputs(8416) <= b;
    outputs(8417) <= a and not b;
    outputs(8418) <= a and b;
    outputs(8419) <= b;
    outputs(8420) <= b;
    outputs(8421) <= a xor b;
    outputs(8422) <= not b;
    outputs(8423) <= not a;
    outputs(8424) <= a or b;
    outputs(8425) <= a xor b;
    outputs(8426) <= not a;
    outputs(8427) <= not a;
    outputs(8428) <= a;
    outputs(8429) <= a xor b;
    outputs(8430) <= not b;
    outputs(8431) <= not a;
    outputs(8432) <= not (a xor b);
    outputs(8433) <= not b;
    outputs(8434) <= not (a and b);
    outputs(8435) <= not b;
    outputs(8436) <= b;
    outputs(8437) <= a and b;
    outputs(8438) <= b and not a;
    outputs(8439) <= b;
    outputs(8440) <= not a;
    outputs(8441) <= not (a xor b);
    outputs(8442) <= not b;
    outputs(8443) <= not (a and b);
    outputs(8444) <= a xor b;
    outputs(8445) <= not a;
    outputs(8446) <= not b;
    outputs(8447) <= not b;
    outputs(8448) <= a xor b;
    outputs(8449) <= not b or a;
    outputs(8450) <= not (a xor b);
    outputs(8451) <= a xor b;
    outputs(8452) <= not (a xor b);
    outputs(8453) <= not (a xor b);
    outputs(8454) <= not a;
    outputs(8455) <= a;
    outputs(8456) <= not (a xor b);
    outputs(8457) <= not (a xor b);
    outputs(8458) <= b;
    outputs(8459) <= '0';
    outputs(8460) <= not b;
    outputs(8461) <= not b;
    outputs(8462) <= not (a xor b);
    outputs(8463) <= a or b;
    outputs(8464) <= not (a and b);
    outputs(8465) <= not a;
    outputs(8466) <= b;
    outputs(8467) <= not a;
    outputs(8468) <= not a or b;
    outputs(8469) <= not b;
    outputs(8470) <= not b;
    outputs(8471) <= a xor b;
    outputs(8472) <= a xor b;
    outputs(8473) <= a xor b;
    outputs(8474) <= not b or a;
    outputs(8475) <= a or b;
    outputs(8476) <= not a;
    outputs(8477) <= a;
    outputs(8478) <= not (a xor b);
    outputs(8479) <= a xor b;
    outputs(8480) <= not b;
    outputs(8481) <= not a or b;
    outputs(8482) <= not a or b;
    outputs(8483) <= not (a xor b);
    outputs(8484) <= a;
    outputs(8485) <= b;
    outputs(8486) <= not b;
    outputs(8487) <= b;
    outputs(8488) <= a;
    outputs(8489) <= a;
    outputs(8490) <= not (a or b);
    outputs(8491) <= not (a xor b);
    outputs(8492) <= a;
    outputs(8493) <= a xor b;
    outputs(8494) <= a and b;
    outputs(8495) <= a xor b;
    outputs(8496) <= not (a xor b);
    outputs(8497) <= a xor b;
    outputs(8498) <= b;
    outputs(8499) <= a and b;
    outputs(8500) <= a;
    outputs(8501) <= not (a xor b);
    outputs(8502) <= not a;
    outputs(8503) <= not b;
    outputs(8504) <= a;
    outputs(8505) <= b;
    outputs(8506) <= not b or a;
    outputs(8507) <= not a;
    outputs(8508) <= b;
    outputs(8509) <= not a;
    outputs(8510) <= not (a or b);
    outputs(8511) <= b;
    outputs(8512) <= a and b;
    outputs(8513) <= not b or a;
    outputs(8514) <= not a or b;
    outputs(8515) <= a xor b;
    outputs(8516) <= not (a xor b);
    outputs(8517) <= not b;
    outputs(8518) <= b;
    outputs(8519) <= a xor b;
    outputs(8520) <= not (a and b);
    outputs(8521) <= a xor b;
    outputs(8522) <= not (a xor b);
    outputs(8523) <= not a or b;
    outputs(8524) <= a;
    outputs(8525) <= a xor b;
    outputs(8526) <= a or b;
    outputs(8527) <= a and b;
    outputs(8528) <= not b;
    outputs(8529) <= not (a xor b);
    outputs(8530) <= a;
    outputs(8531) <= not a or b;
    outputs(8532) <= not (a and b);
    outputs(8533) <= a and not b;
    outputs(8534) <= a;
    outputs(8535) <= b;
    outputs(8536) <= a or b;
    outputs(8537) <= a and b;
    outputs(8538) <= b and not a;
    outputs(8539) <= b;
    outputs(8540) <= a xor b;
    outputs(8541) <= a xor b;
    outputs(8542) <= not b;
    outputs(8543) <= not (a and b);
    outputs(8544) <= b;
    outputs(8545) <= b;
    outputs(8546) <= a and b;
    outputs(8547) <= not a;
    outputs(8548) <= a xor b;
    outputs(8549) <= b and not a;
    outputs(8550) <= b and not a;
    outputs(8551) <= a xor b;
    outputs(8552) <= not b;
    outputs(8553) <= a xor b;
    outputs(8554) <= not b or a;
    outputs(8555) <= a;
    outputs(8556) <= a xor b;
    outputs(8557) <= not a or b;
    outputs(8558) <= a xor b;
    outputs(8559) <= a xor b;
    outputs(8560) <= not a;
    outputs(8561) <= a xor b;
    outputs(8562) <= not a;
    outputs(8563) <= not b;
    outputs(8564) <= a xor b;
    outputs(8565) <= a xor b;
    outputs(8566) <= not a;
    outputs(8567) <= not a;
    outputs(8568) <= not (a and b);
    outputs(8569) <= not (a xor b);
    outputs(8570) <= b;
    outputs(8571) <= b and not a;
    outputs(8572) <= not (a or b);
    outputs(8573) <= not (a xor b);
    outputs(8574) <= a and b;
    outputs(8575) <= a;
    outputs(8576) <= not a;
    outputs(8577) <= not a;
    outputs(8578) <= a xor b;
    outputs(8579) <= a xor b;
    outputs(8580) <= a xor b;
    outputs(8581) <= b;
    outputs(8582) <= not b;
    outputs(8583) <= not b;
    outputs(8584) <= b;
    outputs(8585) <= not a;
    outputs(8586) <= a xor b;
    outputs(8587) <= a xor b;
    outputs(8588) <= a;
    outputs(8589) <= a and b;
    outputs(8590) <= not (a xor b);
    outputs(8591) <= not b;
    outputs(8592) <= not (a and b);
    outputs(8593) <= not a;
    outputs(8594) <= a or b;
    outputs(8595) <= a and not b;
    outputs(8596) <= a xor b;
    outputs(8597) <= not a;
    outputs(8598) <= not (a xor b);
    outputs(8599) <= not (a xor b);
    outputs(8600) <= not b;
    outputs(8601) <= a and not b;
    outputs(8602) <= not a;
    outputs(8603) <= not (a xor b);
    outputs(8604) <= a xor b;
    outputs(8605) <= b;
    outputs(8606) <= not b;
    outputs(8607) <= a;
    outputs(8608) <= not a;
    outputs(8609) <= not b;
    outputs(8610) <= not (a or b);
    outputs(8611) <= a xor b;
    outputs(8612) <= a and not b;
    outputs(8613) <= b;
    outputs(8614) <= not a or b;
    outputs(8615) <= a;
    outputs(8616) <= a or b;
    outputs(8617) <= a xor b;
    outputs(8618) <= a xor b;
    outputs(8619) <= a and not b;
    outputs(8620) <= not a or b;
    outputs(8621) <= a;
    outputs(8622) <= not (a xor b);
    outputs(8623) <= a;
    outputs(8624) <= b and not a;
    outputs(8625) <= not (a xor b);
    outputs(8626) <= not a or b;
    outputs(8627) <= a or b;
    outputs(8628) <= not (a xor b);
    outputs(8629) <= a xor b;
    outputs(8630) <= a and b;
    outputs(8631) <= not (a xor b);
    outputs(8632) <= not (a xor b);
    outputs(8633) <= b;
    outputs(8634) <= not (a xor b);
    outputs(8635) <= a and b;
    outputs(8636) <= not (a xor b);
    outputs(8637) <= a;
    outputs(8638) <= not a;
    outputs(8639) <= not a;
    outputs(8640) <= a;
    outputs(8641) <= a xor b;
    outputs(8642) <= a;
    outputs(8643) <= not b;
    outputs(8644) <= a;
    outputs(8645) <= b;
    outputs(8646) <= b;
    outputs(8647) <= not (a xor b);
    outputs(8648) <= b;
    outputs(8649) <= not (a xor b);
    outputs(8650) <= a and not b;
    outputs(8651) <= not b or a;
    outputs(8652) <= not a;
    outputs(8653) <= b;
    outputs(8654) <= not (a xor b);
    outputs(8655) <= not b;
    outputs(8656) <= not (a and b);
    outputs(8657) <= a xor b;
    outputs(8658) <= not b;
    outputs(8659) <= a xor b;
    outputs(8660) <= a;
    outputs(8661) <= not b;
    outputs(8662) <= b;
    outputs(8663) <= not a;
    outputs(8664) <= not (a xor b);
    outputs(8665) <= not a or b;
    outputs(8666) <= not (a xor b);
    outputs(8667) <= a or b;
    outputs(8668) <= not b;
    outputs(8669) <= not (a xor b);
    outputs(8670) <= b;
    outputs(8671) <= b;
    outputs(8672) <= not b;
    outputs(8673) <= b;
    outputs(8674) <= b and not a;
    outputs(8675) <= not (a xor b);
    outputs(8676) <= b;
    outputs(8677) <= not (a and b);
    outputs(8678) <= not (a and b);
    outputs(8679) <= not b or a;
    outputs(8680) <= not (a or b);
    outputs(8681) <= a xor b;
    outputs(8682) <= a xor b;
    outputs(8683) <= a and not b;
    outputs(8684) <= a;
    outputs(8685) <= not b;
    outputs(8686) <= a xor b;
    outputs(8687) <= not (a or b);
    outputs(8688) <= not a;
    outputs(8689) <= not (a xor b);
    outputs(8690) <= not b;
    outputs(8691) <= not b;
    outputs(8692) <= a;
    outputs(8693) <= not b or a;
    outputs(8694) <= b;
    outputs(8695) <= a and not b;
    outputs(8696) <= not b or a;
    outputs(8697) <= not (a xor b);
    outputs(8698) <= a xor b;
    outputs(8699) <= b and not a;
    outputs(8700) <= not b or a;
    outputs(8701) <= a xor b;
    outputs(8702) <= not a or b;
    outputs(8703) <= not a;
    outputs(8704) <= a;
    outputs(8705) <= a xor b;
    outputs(8706) <= not b;
    outputs(8707) <= not a;
    outputs(8708) <= '1';
    outputs(8709) <= not b;
    outputs(8710) <= not b;
    outputs(8711) <= not (a and b);
    outputs(8712) <= not (a xor b);
    outputs(8713) <= not (a or b);
    outputs(8714) <= not (a or b);
    outputs(8715) <= a xor b;
    outputs(8716) <= a;
    outputs(8717) <= a;
    outputs(8718) <= not b or a;
    outputs(8719) <= b and not a;
    outputs(8720) <= a xor b;
    outputs(8721) <= not (a or b);
    outputs(8722) <= not a or b;
    outputs(8723) <= not a;
    outputs(8724) <= b;
    outputs(8725) <= not a;
    outputs(8726) <= a or b;
    outputs(8727) <= not (a xor b);
    outputs(8728) <= not (a xor b);
    outputs(8729) <= not b;
    outputs(8730) <= a;
    outputs(8731) <= a xor b;
    outputs(8732) <= not a;
    outputs(8733) <= a;
    outputs(8734) <= a xor b;
    outputs(8735) <= a;
    outputs(8736) <= a and b;
    outputs(8737) <= not (a and b);
    outputs(8738) <= a and not b;
    outputs(8739) <= not (a and b);
    outputs(8740) <= a and not b;
    outputs(8741) <= b;
    outputs(8742) <= not (a xor b);
    outputs(8743) <= b;
    outputs(8744) <= not (a or b);
    outputs(8745) <= not b;
    outputs(8746) <= not (a xor b);
    outputs(8747) <= not b or a;
    outputs(8748) <= not b;
    outputs(8749) <= not (a xor b);
    outputs(8750) <= a;
    outputs(8751) <= b;
    outputs(8752) <= a xor b;
    outputs(8753) <= not a;
    outputs(8754) <= a;
    outputs(8755) <= a;
    outputs(8756) <= b;
    outputs(8757) <= a and not b;
    outputs(8758) <= a;
    outputs(8759) <= not b;
    outputs(8760) <= a xor b;
    outputs(8761) <= not b or a;
    outputs(8762) <= a xor b;
    outputs(8763) <= not a or b;
    outputs(8764) <= a;
    outputs(8765) <= not a;
    outputs(8766) <= not b;
    outputs(8767) <= not a or b;
    outputs(8768) <= a or b;
    outputs(8769) <= not b or a;
    outputs(8770) <= not b;
    outputs(8771) <= not b;
    outputs(8772) <= a;
    outputs(8773) <= not a;
    outputs(8774) <= a xor b;
    outputs(8775) <= a and b;
    outputs(8776) <= a xor b;
    outputs(8777) <= not b;
    outputs(8778) <= not (a and b);
    outputs(8779) <= not (a xor b);
    outputs(8780) <= a;
    outputs(8781) <= not (a xor b);
    outputs(8782) <= b and not a;
    outputs(8783) <= not (a xor b);
    outputs(8784) <= not a;
    outputs(8785) <= a xor b;
    outputs(8786) <= a and b;
    outputs(8787) <= a and not b;
    outputs(8788) <= a xor b;
    outputs(8789) <= b and not a;
    outputs(8790) <= not b or a;
    outputs(8791) <= not a or b;
    outputs(8792) <= not b;
    outputs(8793) <= not b or a;
    outputs(8794) <= a xor b;
    outputs(8795) <= b and not a;
    outputs(8796) <= a or b;
    outputs(8797) <= b;
    outputs(8798) <= b;
    outputs(8799) <= a xor b;
    outputs(8800) <= not (a xor b);
    outputs(8801) <= not (a or b);
    outputs(8802) <= b;
    outputs(8803) <= not b;
    outputs(8804) <= not (a xor b);
    outputs(8805) <= a;
    outputs(8806) <= a xor b;
    outputs(8807) <= a and not b;
    outputs(8808) <= b and not a;
    outputs(8809) <= not (a and b);
    outputs(8810) <= not a;
    outputs(8811) <= a xor b;
    outputs(8812) <= b and not a;
    outputs(8813) <= a and not b;
    outputs(8814) <= not b or a;
    outputs(8815) <= a xor b;
    outputs(8816) <= a;
    outputs(8817) <= not b;
    outputs(8818) <= not b;
    outputs(8819) <= a xor b;
    outputs(8820) <= a and not b;
    outputs(8821) <= not a;
    outputs(8822) <= b;
    outputs(8823) <= not (a xor b);
    outputs(8824) <= not a;
    outputs(8825) <= not (a xor b);
    outputs(8826) <= not (a xor b);
    outputs(8827) <= not (a and b);
    outputs(8828) <= a;
    outputs(8829) <= not (a and b);
    outputs(8830) <= a xor b;
    outputs(8831) <= a xor b;
    outputs(8832) <= not (a xor b);
    outputs(8833) <= not (a and b);
    outputs(8834) <= b;
    outputs(8835) <= not (a xor b);
    outputs(8836) <= not (a and b);
    outputs(8837) <= a and b;
    outputs(8838) <= not a or b;
    outputs(8839) <= not b or a;
    outputs(8840) <= not (a xor b);
    outputs(8841) <= not b;
    outputs(8842) <= not (a xor b);
    outputs(8843) <= not (a xor b);
    outputs(8844) <= a xor b;
    outputs(8845) <= b;
    outputs(8846) <= not (a or b);
    outputs(8847) <= a xor b;
    outputs(8848) <= not a;
    outputs(8849) <= a xor b;
    outputs(8850) <= b;
    outputs(8851) <= a and b;
    outputs(8852) <= b;
    outputs(8853) <= b;
    outputs(8854) <= a xor b;
    outputs(8855) <= b;
    outputs(8856) <= not b or a;
    outputs(8857) <= a and not b;
    outputs(8858) <= a;
    outputs(8859) <= b;
    outputs(8860) <= not b;
    outputs(8861) <= not a or b;
    outputs(8862) <= b and not a;
    outputs(8863) <= a or b;
    outputs(8864) <= a and not b;
    outputs(8865) <= b and not a;
    outputs(8866) <= not b;
    outputs(8867) <= a and not b;
    outputs(8868) <= a and b;
    outputs(8869) <= not a;
    outputs(8870) <= not b or a;
    outputs(8871) <= a and not b;
    outputs(8872) <= not (a xor b);
    outputs(8873) <= a xor b;
    outputs(8874) <= not (a xor b);
    outputs(8875) <= not (a xor b);
    outputs(8876) <= a xor b;
    outputs(8877) <= not a;
    outputs(8878) <= not (a or b);
    outputs(8879) <= not (a or b);
    outputs(8880) <= not (a xor b);
    outputs(8881) <= b;
    outputs(8882) <= a xor b;
    outputs(8883) <= not b;
    outputs(8884) <= not (a xor b);
    outputs(8885) <= a xor b;
    outputs(8886) <= a;
    outputs(8887) <= a and b;
    outputs(8888) <= b;
    outputs(8889) <= not b;
    outputs(8890) <= not (a and b);
    outputs(8891) <= a;
    outputs(8892) <= not b;
    outputs(8893) <= a and not b;
    outputs(8894) <= a and b;
    outputs(8895) <= a and b;
    outputs(8896) <= a or b;
    outputs(8897) <= a xor b;
    outputs(8898) <= a and not b;
    outputs(8899) <= a xor b;
    outputs(8900) <= not b or a;
    outputs(8901) <= a;
    outputs(8902) <= not a;
    outputs(8903) <= a and b;
    outputs(8904) <= not (a xor b);
    outputs(8905) <= not (a xor b);
    outputs(8906) <= not a or b;
    outputs(8907) <= not b;
    outputs(8908) <= a xor b;
    outputs(8909) <= a xor b;
    outputs(8910) <= a and b;
    outputs(8911) <= not a;
    outputs(8912) <= a or b;
    outputs(8913) <= not (a or b);
    outputs(8914) <= not a;
    outputs(8915) <= not (a and b);
    outputs(8916) <= a xor b;
    outputs(8917) <= not a;
    outputs(8918) <= a or b;
    outputs(8919) <= a and not b;
    outputs(8920) <= not (a xor b);
    outputs(8921) <= a;
    outputs(8922) <= a xor b;
    outputs(8923) <= a xor b;
    outputs(8924) <= b;
    outputs(8925) <= not (a xor b);
    outputs(8926) <= not (a xor b);
    outputs(8927) <= b;
    outputs(8928) <= a;
    outputs(8929) <= not (a xor b);
    outputs(8930) <= a;
    outputs(8931) <= a xor b;
    outputs(8932) <= not b;
    outputs(8933) <= not b;
    outputs(8934) <= not b;
    outputs(8935) <= a and not b;
    outputs(8936) <= b;
    outputs(8937) <= not a or b;
    outputs(8938) <= b and not a;
    outputs(8939) <= a xor b;
    outputs(8940) <= not (a xor b);
    outputs(8941) <= not b;
    outputs(8942) <= a xor b;
    outputs(8943) <= not (a or b);
    outputs(8944) <= a;
    outputs(8945) <= b and not a;
    outputs(8946) <= b;
    outputs(8947) <= not (a xor b);
    outputs(8948) <= a or b;
    outputs(8949) <= b;
    outputs(8950) <= not (a xor b);
    outputs(8951) <= b and not a;
    outputs(8952) <= not (a and b);
    outputs(8953) <= a;
    outputs(8954) <= not (a xor b);
    outputs(8955) <= not b;
    outputs(8956) <= a xor b;
    outputs(8957) <= a xor b;
    outputs(8958) <= not (a and b);
    outputs(8959) <= b;
    outputs(8960) <= a and b;
    outputs(8961) <= a xor b;
    outputs(8962) <= not b or a;
    outputs(8963) <= b and not a;
    outputs(8964) <= not (a or b);
    outputs(8965) <= not a;
    outputs(8966) <= not (a xor b);
    outputs(8967) <= a and b;
    outputs(8968) <= b;
    outputs(8969) <= a xor b;
    outputs(8970) <= a and not b;
    outputs(8971) <= a and not b;
    outputs(8972) <= not (a xor b);
    outputs(8973) <= a xor b;
    outputs(8974) <= b;
    outputs(8975) <= not (a and b);
    outputs(8976) <= not a;
    outputs(8977) <= b and not a;
    outputs(8978) <= a and b;
    outputs(8979) <= a xor b;
    outputs(8980) <= a or b;
    outputs(8981) <= b and not a;
    outputs(8982) <= not a;
    outputs(8983) <= not a or b;
    outputs(8984) <= not a;
    outputs(8985) <= a xor b;
    outputs(8986) <= not (a xor b);
    outputs(8987) <= not (a xor b);
    outputs(8988) <= not a or b;
    outputs(8989) <= a and not b;
    outputs(8990) <= a;
    outputs(8991) <= not b;
    outputs(8992) <= a;
    outputs(8993) <= b;
    outputs(8994) <= not (a xor b);
    outputs(8995) <= a xor b;
    outputs(8996) <= a;
    outputs(8997) <= b;
    outputs(8998) <= a;
    outputs(8999) <= not (a xor b);
    outputs(9000) <= not b;
    outputs(9001) <= not (a xor b);
    outputs(9002) <= not a;
    outputs(9003) <= not b or a;
    outputs(9004) <= not (a or b);
    outputs(9005) <= b;
    outputs(9006) <= not b;
    outputs(9007) <= a and b;
    outputs(9008) <= not (a and b);
    outputs(9009) <= not (a xor b);
    outputs(9010) <= a xor b;
    outputs(9011) <= a;
    outputs(9012) <= a xor b;
    outputs(9013) <= not b or a;
    outputs(9014) <= not a;
    outputs(9015) <= a xor b;
    outputs(9016) <= not (a xor b);
    outputs(9017) <= not a;
    outputs(9018) <= not a;
    outputs(9019) <= not b;
    outputs(9020) <= not (a and b);
    outputs(9021) <= not (a xor b);
    outputs(9022) <= not b;
    outputs(9023) <= not a;
    outputs(9024) <= not (a xor b);
    outputs(9025) <= not (a and b);
    outputs(9026) <= a;
    outputs(9027) <= not a;
    outputs(9028) <= not (a and b);
    outputs(9029) <= not b;
    outputs(9030) <= a and b;
    outputs(9031) <= not (a xor b);
    outputs(9032) <= not (a and b);
    outputs(9033) <= b and not a;
    outputs(9034) <= b;
    outputs(9035) <= a xor b;
    outputs(9036) <= not b or a;
    outputs(9037) <= a xor b;
    outputs(9038) <= a xor b;
    outputs(9039) <= b and not a;
    outputs(9040) <= not (a and b);
    outputs(9041) <= not b or a;
    outputs(9042) <= not (a xor b);
    outputs(9043) <= b;
    outputs(9044) <= not b;
    outputs(9045) <= not (a and b);
    outputs(9046) <= a xor b;
    outputs(9047) <= not (a xor b);
    outputs(9048) <= not a;
    outputs(9049) <= not (a xor b);
    outputs(9050) <= a;
    outputs(9051) <= not (a xor b);
    outputs(9052) <= not b;
    outputs(9053) <= not (a xor b);
    outputs(9054) <= not (a xor b);
    outputs(9055) <= a xor b;
    outputs(9056) <= not (a or b);
    outputs(9057) <= b;
    outputs(9058) <= not a;
    outputs(9059) <= not (a and b);
    outputs(9060) <= not b;
    outputs(9061) <= a or b;
    outputs(9062) <= not b;
    outputs(9063) <= not (a and b);
    outputs(9064) <= a;
    outputs(9065) <= a;
    outputs(9066) <= '1';
    outputs(9067) <= not b or a;
    outputs(9068) <= not a;
    outputs(9069) <= not a;
    outputs(9070) <= not b;
    outputs(9071) <= not (a or b);
    outputs(9072) <= a and b;
    outputs(9073) <= a xor b;
    outputs(9074) <= a xor b;
    outputs(9075) <= a;
    outputs(9076) <= b;
    outputs(9077) <= b and not a;
    outputs(9078) <= not (a xor b);
    outputs(9079) <= not (a xor b);
    outputs(9080) <= b;
    outputs(9081) <= a and not b;
    outputs(9082) <= a xor b;
    outputs(9083) <= not a;
    outputs(9084) <= a xor b;
    outputs(9085) <= b;
    outputs(9086) <= a xor b;
    outputs(9087) <= a and not b;
    outputs(9088) <= a xor b;
    outputs(9089) <= not (a or b);
    outputs(9090) <= not a;
    outputs(9091) <= a;
    outputs(9092) <= a xor b;
    outputs(9093) <= a;
    outputs(9094) <= not (a or b);
    outputs(9095) <= not b;
    outputs(9096) <= a xor b;
    outputs(9097) <= b;
    outputs(9098) <= a or b;
    outputs(9099) <= b and not a;
    outputs(9100) <= b;
    outputs(9101) <= not a;
    outputs(9102) <= a or b;
    outputs(9103) <= a xor b;
    outputs(9104) <= b and not a;
    outputs(9105) <= not b;
    outputs(9106) <= not (a or b);
    outputs(9107) <= not a;
    outputs(9108) <= a;
    outputs(9109) <= b;
    outputs(9110) <= b;
    outputs(9111) <= not (a xor b);
    outputs(9112) <= not (a xor b);
    outputs(9113) <= not (a xor b);
    outputs(9114) <= not a;
    outputs(9115) <= b;
    outputs(9116) <= not (a xor b);
    outputs(9117) <= b and not a;
    outputs(9118) <= a xor b;
    outputs(9119) <= a xor b;
    outputs(9120) <= a;
    outputs(9121) <= a xor b;
    outputs(9122) <= not (a xor b);
    outputs(9123) <= not b;
    outputs(9124) <= a and not b;
    outputs(9125) <= b and not a;
    outputs(9126) <= b;
    outputs(9127) <= not b or a;
    outputs(9128) <= not (a xor b);
    outputs(9129) <= not (a and b);
    outputs(9130) <= a and b;
    outputs(9131) <= not b;
    outputs(9132) <= not (a and b);
    outputs(9133) <= b;
    outputs(9134) <= not (a xor b);
    outputs(9135) <= not (a or b);
    outputs(9136) <= a xor b;
    outputs(9137) <= not a;
    outputs(9138) <= a xor b;
    outputs(9139) <= not a;
    outputs(9140) <= not b;
    outputs(9141) <= a xor b;
    outputs(9142) <= not a;
    outputs(9143) <= not (a xor b);
    outputs(9144) <= a xor b;
    outputs(9145) <= not (a or b);
    outputs(9146) <= not (a and b);
    outputs(9147) <= a;
    outputs(9148) <= not (a xor b);
    outputs(9149) <= not (a xor b);
    outputs(9150) <= b and not a;
    outputs(9151) <= not b or a;
    outputs(9152) <= a xor b;
    outputs(9153) <= a xor b;
    outputs(9154) <= a xor b;
    outputs(9155) <= a xor b;
    outputs(9156) <= a;
    outputs(9157) <= a or b;
    outputs(9158) <= not (a xor b);
    outputs(9159) <= not (a or b);
    outputs(9160) <= not b;
    outputs(9161) <= b;
    outputs(9162) <= a;
    outputs(9163) <= b;
    outputs(9164) <= not a or b;
    outputs(9165) <= a xor b;
    outputs(9166) <= not a;
    outputs(9167) <= not (a and b);
    outputs(9168) <= not (a xor b);
    outputs(9169) <= not a or b;
    outputs(9170) <= not b;
    outputs(9171) <= not a;
    outputs(9172) <= not (a or b);
    outputs(9173) <= not (a xor b);
    outputs(9174) <= a xor b;
    outputs(9175) <= not b;
    outputs(9176) <= not (a xor b);
    outputs(9177) <= not a or b;
    outputs(9178) <= a xor b;
    outputs(9179) <= a or b;
    outputs(9180) <= not (a xor b);
    outputs(9181) <= not a;
    outputs(9182) <= not (a xor b);
    outputs(9183) <= not a;
    outputs(9184) <= a xor b;
    outputs(9185) <= a xor b;
    outputs(9186) <= b;
    outputs(9187) <= a xor b;
    outputs(9188) <= a xor b;
    outputs(9189) <= not b;
    outputs(9190) <= b;
    outputs(9191) <= not (a xor b);
    outputs(9192) <= b;
    outputs(9193) <= a and b;
    outputs(9194) <= b and not a;
    outputs(9195) <= a and not b;
    outputs(9196) <= a or b;
    outputs(9197) <= not a;
    outputs(9198) <= a;
    outputs(9199) <= a xor b;
    outputs(9200) <= not a;
    outputs(9201) <= a and not b;
    outputs(9202) <= a;
    outputs(9203) <= a or b;
    outputs(9204) <= a and b;
    outputs(9205) <= a or b;
    outputs(9206) <= a;
    outputs(9207) <= not b;
    outputs(9208) <= not b;
    outputs(9209) <= a;
    outputs(9210) <= not b;
    outputs(9211) <= a xor b;
    outputs(9212) <= a xor b;
    outputs(9213) <= not (a or b);
    outputs(9214) <= not a or b;
    outputs(9215) <= a xor b;
    outputs(9216) <= not a;
    outputs(9217) <= a xor b;
    outputs(9218) <= not (a xor b);
    outputs(9219) <= not a;
    outputs(9220) <= b and not a;
    outputs(9221) <= not (a or b);
    outputs(9222) <= a and b;
    outputs(9223) <= a;
    outputs(9224) <= a;
    outputs(9225) <= not (a or b);
    outputs(9226) <= a xor b;
    outputs(9227) <= a and not b;
    outputs(9228) <= a xor b;
    outputs(9229) <= not b or a;
    outputs(9230) <= not (a or b);
    outputs(9231) <= a;
    outputs(9232) <= not b;
    outputs(9233) <= a xor b;
    outputs(9234) <= a xor b;
    outputs(9235) <= not a;
    outputs(9236) <= not (a xor b);
    outputs(9237) <= a and not b;
    outputs(9238) <= not (a xor b);
    outputs(9239) <= not a;
    outputs(9240) <= not b or a;
    outputs(9241) <= not a;
    outputs(9242) <= a xor b;
    outputs(9243) <= not (a xor b);
    outputs(9244) <= b and not a;
    outputs(9245) <= not (a and b);
    outputs(9246) <= a and not b;
    outputs(9247) <= not a;
    outputs(9248) <= b and not a;
    outputs(9249) <= not a or b;
    outputs(9250) <= a xor b;
    outputs(9251) <= not (a xor b);
    outputs(9252) <= a;
    outputs(9253) <= a and not b;
    outputs(9254) <= not (a xor b);
    outputs(9255) <= not (a or b);
    outputs(9256) <= a xor b;
    outputs(9257) <= b;
    outputs(9258) <= not b;
    outputs(9259) <= a;
    outputs(9260) <= not a;
    outputs(9261) <= b and not a;
    outputs(9262) <= not a;
    outputs(9263) <= not (a or b);
    outputs(9264) <= not (a xor b);
    outputs(9265) <= not (a or b);
    outputs(9266) <= not (a or b);
    outputs(9267) <= b;
    outputs(9268) <= not a or b;
    outputs(9269) <= a and not b;
    outputs(9270) <= not b;
    outputs(9271) <= a xor b;
    outputs(9272) <= not (a xor b);
    outputs(9273) <= a;
    outputs(9274) <= a xor b;
    outputs(9275) <= a xor b;
    outputs(9276) <= not b or a;
    outputs(9277) <= b and not a;
    outputs(9278) <= not b or a;
    outputs(9279) <= b and not a;
    outputs(9280) <= not b;
    outputs(9281) <= not a;
    outputs(9282) <= a xor b;
    outputs(9283) <= not (a xor b);
    outputs(9284) <= b;
    outputs(9285) <= a xor b;
    outputs(9286) <= not b;
    outputs(9287) <= a and b;
    outputs(9288) <= a xor b;
    outputs(9289) <= not (a xor b);
    outputs(9290) <= not a;
    outputs(9291) <= a xor b;
    outputs(9292) <= b;
    outputs(9293) <= a xor b;
    outputs(9294) <= not (a xor b);
    outputs(9295) <= not (a or b);
    outputs(9296) <= a;
    outputs(9297) <= not b or a;
    outputs(9298) <= a and not b;
    outputs(9299) <= not b or a;
    outputs(9300) <= a;
    outputs(9301) <= not a;
    outputs(9302) <= a and b;
    outputs(9303) <= not (a or b);
    outputs(9304) <= a and not b;
    outputs(9305) <= a;
    outputs(9306) <= a xor b;
    outputs(9307) <= not b or a;
    outputs(9308) <= a xor b;
    outputs(9309) <= b and not a;
    outputs(9310) <= a xor b;
    outputs(9311) <= not (a and b);
    outputs(9312) <= b and not a;
    outputs(9313) <= not b;
    outputs(9314) <= a and b;
    outputs(9315) <= not (a and b);
    outputs(9316) <= not a;
    outputs(9317) <= not (a xor b);
    outputs(9318) <= not (a or b);
    outputs(9319) <= a and b;
    outputs(9320) <= not (a or b);
    outputs(9321) <= b;
    outputs(9322) <= not (a and b);
    outputs(9323) <= a xor b;
    outputs(9324) <= not b;
    outputs(9325) <= a and not b;
    outputs(9326) <= not (a or b);
    outputs(9327) <= not a or b;
    outputs(9328) <= not (a xor b);
    outputs(9329) <= a and not b;
    outputs(9330) <= not b;
    outputs(9331) <= a xor b;
    outputs(9332) <= not b;
    outputs(9333) <= b;
    outputs(9334) <= not b;
    outputs(9335) <= a and not b;
    outputs(9336) <= not (a and b);
    outputs(9337) <= not (a or b);
    outputs(9338) <= b;
    outputs(9339) <= not (a and b);
    outputs(9340) <= a and b;
    outputs(9341) <= a and b;
    outputs(9342) <= a;
    outputs(9343) <= a;
    outputs(9344) <= b;
    outputs(9345) <= b;
    outputs(9346) <= not (a xor b);
    outputs(9347) <= a xor b;
    outputs(9348) <= a and not b;
    outputs(9349) <= a and not b;
    outputs(9350) <= b;
    outputs(9351) <= not (a xor b);
    outputs(9352) <= not (a and b);
    outputs(9353) <= not (a or b);
    outputs(9354) <= b;
    outputs(9355) <= not (a xor b);
    outputs(9356) <= not (a xor b);
    outputs(9357) <= a and not b;
    outputs(9358) <= a xor b;
    outputs(9359) <= a xor b;
    outputs(9360) <= not (a xor b);
    outputs(9361) <= a;
    outputs(9362) <= not (a and b);
    outputs(9363) <= a xor b;
    outputs(9364) <= a and b;
    outputs(9365) <= a xor b;
    outputs(9366) <= a xor b;
    outputs(9367) <= not b or a;
    outputs(9368) <= a and not b;
    outputs(9369) <= a;
    outputs(9370) <= not (a or b);
    outputs(9371) <= not a;
    outputs(9372) <= b and not a;
    outputs(9373) <= a and b;
    outputs(9374) <= a xor b;
    outputs(9375) <= b;
    outputs(9376) <= b;
    outputs(9377) <= a and b;
    outputs(9378) <= not a;
    outputs(9379) <= b;
    outputs(9380) <= not (a xor b);
    outputs(9381) <= a;
    outputs(9382) <= a and not b;
    outputs(9383) <= not b;
    outputs(9384) <= a xor b;
    outputs(9385) <= a and b;
    outputs(9386) <= not a;
    outputs(9387) <= not (a xor b);
    outputs(9388) <= a;
    outputs(9389) <= not (a or b);
    outputs(9390) <= a and b;
    outputs(9391) <= not (a xor b);
    outputs(9392) <= a or b;
    outputs(9393) <= not (a or b);
    outputs(9394) <= a and b;
    outputs(9395) <= not (a or b);
    outputs(9396) <= not (a xor b);
    outputs(9397) <= a;
    outputs(9398) <= a xor b;
    outputs(9399) <= a;
    outputs(9400) <= b and not a;
    outputs(9401) <= a;
    outputs(9402) <= not a;
    outputs(9403) <= not a;
    outputs(9404) <= b;
    outputs(9405) <= not (a xor b);
    outputs(9406) <= not (a xor b);
    outputs(9407) <= a;
    outputs(9408) <= not (a and b);
    outputs(9409) <= a and b;
    outputs(9410) <= not b;
    outputs(9411) <= not (a xor b);
    outputs(9412) <= b and not a;
    outputs(9413) <= b;
    outputs(9414) <= not (a xor b);
    outputs(9415) <= a and b;
    outputs(9416) <= not b;
    outputs(9417) <= a and not b;
    outputs(9418) <= a;
    outputs(9419) <= b and not a;
    outputs(9420) <= a and b;
    outputs(9421) <= b and not a;
    outputs(9422) <= not a;
    outputs(9423) <= not (a xor b);
    outputs(9424) <= not a;
    outputs(9425) <= not (a xor b);
    outputs(9426) <= a;
    outputs(9427) <= b;
    outputs(9428) <= a xor b;
    outputs(9429) <= not (a xor b);
    outputs(9430) <= a xor b;
    outputs(9431) <= not b or a;
    outputs(9432) <= not (a or b);
    outputs(9433) <= b and not a;
    outputs(9434) <= not (a xor b);
    outputs(9435) <= not (a xor b);
    outputs(9436) <= a xor b;
    outputs(9437) <= b;
    outputs(9438) <= a and b;
    outputs(9439) <= not (a xor b);
    outputs(9440) <= b;
    outputs(9441) <= b and not a;
    outputs(9442) <= not (a xor b);
    outputs(9443) <= not a;
    outputs(9444) <= a and not b;
    outputs(9445) <= a;
    outputs(9446) <= not (a and b);
    outputs(9447) <= a xor b;
    outputs(9448) <= a xor b;
    outputs(9449) <= not (a or b);
    outputs(9450) <= a;
    outputs(9451) <= not a;
    outputs(9452) <= a xor b;
    outputs(9453) <= b and not a;
    outputs(9454) <= b;
    outputs(9455) <= not (a or b);
    outputs(9456) <= a and not b;
    outputs(9457) <= not a;
    outputs(9458) <= a xor b;
    outputs(9459) <= not (a xor b);
    outputs(9460) <= not (a and b);
    outputs(9461) <= not (a and b);
    outputs(9462) <= not (a or b);
    outputs(9463) <= not (a xor b);
    outputs(9464) <= not (a xor b);
    outputs(9465) <= not a or b;
    outputs(9466) <= a or b;
    outputs(9467) <= b;
    outputs(9468) <= a and not b;
    outputs(9469) <= not (a xor b);
    outputs(9470) <= not (a xor b);
    outputs(9471) <= a and b;
    outputs(9472) <= not b;
    outputs(9473) <= a and b;
    outputs(9474) <= not a;
    outputs(9475) <= a;
    outputs(9476) <= a;
    outputs(9477) <= not (a or b);
    outputs(9478) <= not (a or b);
    outputs(9479) <= not (a xor b);
    outputs(9480) <= not b;
    outputs(9481) <= not b;
    outputs(9482) <= not (a xor b);
    outputs(9483) <= a and b;
    outputs(9484) <= a xor b;
    outputs(9485) <= a and not b;
    outputs(9486) <= b;
    outputs(9487) <= not (a xor b);
    outputs(9488) <= a and b;
    outputs(9489) <= not (a or b);
    outputs(9490) <= not (a or b);
    outputs(9491) <= b;
    outputs(9492) <= b;
    outputs(9493) <= a xor b;
    outputs(9494) <= a xor b;
    outputs(9495) <= a and not b;
    outputs(9496) <= a xor b;
    outputs(9497) <= not (a xor b);
    outputs(9498) <= not (a or b);
    outputs(9499) <= b;
    outputs(9500) <= a and not b;
    outputs(9501) <= b and not a;
    outputs(9502) <= not (a and b);
    outputs(9503) <= not (a or b);
    outputs(9504) <= not a;
    outputs(9505) <= not (a and b);
    outputs(9506) <= not (a xor b);
    outputs(9507) <= b and not a;
    outputs(9508) <= not (a xor b);
    outputs(9509) <= a and b;
    outputs(9510) <= b and not a;
    outputs(9511) <= a and not b;
    outputs(9512) <= b;
    outputs(9513) <= a xor b;
    outputs(9514) <= not (a and b);
    outputs(9515) <= not (a xor b);
    outputs(9516) <= a xor b;
    outputs(9517) <= not a;
    outputs(9518) <= a xor b;
    outputs(9519) <= not (a xor b);
    outputs(9520) <= not a or b;
    outputs(9521) <= a and b;
    outputs(9522) <= not (a xor b);
    outputs(9523) <= b and not a;
    outputs(9524) <= a xor b;
    outputs(9525) <= a xor b;
    outputs(9526) <= a xor b;
    outputs(9527) <= not a;
    outputs(9528) <= b;
    outputs(9529) <= b;
    outputs(9530) <= not (a xor b);
    outputs(9531) <= not b;
    outputs(9532) <= b;
    outputs(9533) <= not b or a;
    outputs(9534) <= not (a and b);
    outputs(9535) <= a and not b;
    outputs(9536) <= not a;
    outputs(9537) <= not (a or b);
    outputs(9538) <= a xor b;
    outputs(9539) <= a;
    outputs(9540) <= b and not a;
    outputs(9541) <= not a or b;
    outputs(9542) <= b and not a;
    outputs(9543) <= a and b;
    outputs(9544) <= b;
    outputs(9545) <= not (a or b);
    outputs(9546) <= not b;
    outputs(9547) <= a xor b;
    outputs(9548) <= a and b;
    outputs(9549) <= not a;
    outputs(9550) <= b and not a;
    outputs(9551) <= not (a or b);
    outputs(9552) <= '1';
    outputs(9553) <= not (a xor b);
    outputs(9554) <= not (a or b);
    outputs(9555) <= not b;
    outputs(9556) <= a and not b;
    outputs(9557) <= not (a xor b);
    outputs(9558) <= not b;
    outputs(9559) <= a;
    outputs(9560) <= not a;
    outputs(9561) <= a;
    outputs(9562) <= a and b;
    outputs(9563) <= b and not a;
    outputs(9564) <= a and not b;
    outputs(9565) <= not b;
    outputs(9566) <= b;
    outputs(9567) <= not (a xor b);
    outputs(9568) <= not (a xor b);
    outputs(9569) <= not b or a;
    outputs(9570) <= b and not a;
    outputs(9571) <= not a;
    outputs(9572) <= not (a xor b);
    outputs(9573) <= not b;
    outputs(9574) <= a;
    outputs(9575) <= a xor b;
    outputs(9576) <= not (a xor b);
    outputs(9577) <= not (a or b);
    outputs(9578) <= not b;
    outputs(9579) <= a and b;
    outputs(9580) <= b;
    outputs(9581) <= a;
    outputs(9582) <= not (a or b);
    outputs(9583) <= a xor b;
    outputs(9584) <= b and not a;
    outputs(9585) <= not (a xor b);
    outputs(9586) <= not b;
    outputs(9587) <= a and not b;
    outputs(9588) <= not (a xor b);
    outputs(9589) <= b;
    outputs(9590) <= not b;
    outputs(9591) <= not (a or b);
    outputs(9592) <= b;
    outputs(9593) <= not (a xor b);
    outputs(9594) <= b;
    outputs(9595) <= b and not a;
    outputs(9596) <= b;
    outputs(9597) <= not b or a;
    outputs(9598) <= b;
    outputs(9599) <= b and not a;
    outputs(9600) <= not a;
    outputs(9601) <= not (a and b);
    outputs(9602) <= not a;
    outputs(9603) <= not b or a;
    outputs(9604) <= not (a or b);
    outputs(9605) <= not b;
    outputs(9606) <= not b;
    outputs(9607) <= not (a xor b);
    outputs(9608) <= not b or a;
    outputs(9609) <= b;
    outputs(9610) <= not (a xor b);
    outputs(9611) <= a and b;
    outputs(9612) <= not b;
    outputs(9613) <= b;
    outputs(9614) <= a;
    outputs(9615) <= a xor b;
    outputs(9616) <= not (a xor b);
    outputs(9617) <= b;
    outputs(9618) <= a and not b;
    outputs(9619) <= a and b;
    outputs(9620) <= b;
    outputs(9621) <= not (a xor b);
    outputs(9622) <= a xor b;
    outputs(9623) <= b and not a;
    outputs(9624) <= b and not a;
    outputs(9625) <= a;
    outputs(9626) <= not a;
    outputs(9627) <= not (a or b);
    outputs(9628) <= not a or b;
    outputs(9629) <= not b or a;
    outputs(9630) <= a and b;
    outputs(9631) <= not (a and b);
    outputs(9632) <= a xor b;
    outputs(9633) <= a and b;
    outputs(9634) <= not (a and b);
    outputs(9635) <= not (a and b);
    outputs(9636) <= a and not b;
    outputs(9637) <= not b;
    outputs(9638) <= not a;
    outputs(9639) <= b and not a;
    outputs(9640) <= b and not a;
    outputs(9641) <= a and b;
    outputs(9642) <= not (a xor b);
    outputs(9643) <= a xor b;
    outputs(9644) <= a xor b;
    outputs(9645) <= not b;
    outputs(9646) <= not b;
    outputs(9647) <= not (a xor b);
    outputs(9648) <= not (a xor b);
    outputs(9649) <= a;
    outputs(9650) <= a xor b;
    outputs(9651) <= a and not b;
    outputs(9652) <= b and not a;
    outputs(9653) <= a and not b;
    outputs(9654) <= not b;
    outputs(9655) <= a and b;
    outputs(9656) <= a and b;
    outputs(9657) <= a and not b;
    outputs(9658) <= a and not b;
    outputs(9659) <= a xor b;
    outputs(9660) <= b and not a;
    outputs(9661) <= a or b;
    outputs(9662) <= not (a xor b);
    outputs(9663) <= not a or b;
    outputs(9664) <= a;
    outputs(9665) <= not a;
    outputs(9666) <= a xor b;
    outputs(9667) <= a xor b;
    outputs(9668) <= not a;
    outputs(9669) <= not a;
    outputs(9670) <= not b;
    outputs(9671) <= not (a or b);
    outputs(9672) <= a;
    outputs(9673) <= b;
    outputs(9674) <= not (a xor b);
    outputs(9675) <= a;
    outputs(9676) <= not b or a;
    outputs(9677) <= b and not a;
    outputs(9678) <= not a;
    outputs(9679) <= a;
    outputs(9680) <= a xor b;
    outputs(9681) <= not a;
    outputs(9682) <= not a or b;
    outputs(9683) <= b;
    outputs(9684) <= a or b;
    outputs(9685) <= not a;
    outputs(9686) <= not b;
    outputs(9687) <= a;
    outputs(9688) <= not (a xor b);
    outputs(9689) <= b;
    outputs(9690) <= not a or b;
    outputs(9691) <= not (a xor b);
    outputs(9692) <= not (a and b);
    outputs(9693) <= not (a or b);
    outputs(9694) <= b and not a;
    outputs(9695) <= b;
    outputs(9696) <= b;
    outputs(9697) <= b and not a;
    outputs(9698) <= not b;
    outputs(9699) <= not b;
    outputs(9700) <= a and not b;
    outputs(9701) <= not (a xor b);
    outputs(9702) <= a xor b;
    outputs(9703) <= not (a and b);
    outputs(9704) <= a xor b;
    outputs(9705) <= not a;
    outputs(9706) <= b;
    outputs(9707) <= a and b;
    outputs(9708) <= a;
    outputs(9709) <= a and b;
    outputs(9710) <= not (a xor b);
    outputs(9711) <= b;
    outputs(9712) <= not a;
    outputs(9713) <= not (a xor b);
    outputs(9714) <= a and b;
    outputs(9715) <= a xor b;
    outputs(9716) <= not (a xor b);
    outputs(9717) <= a xor b;
    outputs(9718) <= b;
    outputs(9719) <= b and not a;
    outputs(9720) <= not (a or b);
    outputs(9721) <= not (a and b);
    outputs(9722) <= not b;
    outputs(9723) <= not (a xor b);
    outputs(9724) <= not (a or b);
    outputs(9725) <= a and not b;
    outputs(9726) <= a;
    outputs(9727) <= a xor b;
    outputs(9728) <= b;
    outputs(9729) <= a and b;
    outputs(9730) <= not b;
    outputs(9731) <= a;
    outputs(9732) <= b and not a;
    outputs(9733) <= a;
    outputs(9734) <= a;
    outputs(9735) <= a and b;
    outputs(9736) <= not (a xor b);
    outputs(9737) <= not b;
    outputs(9738) <= a xor b;
    outputs(9739) <= a and b;
    outputs(9740) <= a and b;
    outputs(9741) <= b;
    outputs(9742) <= a;
    outputs(9743) <= a xor b;
    outputs(9744) <= not a;
    outputs(9745) <= a xor b;
    outputs(9746) <= a and b;
    outputs(9747) <= a xor b;
    outputs(9748) <= not b or a;
    outputs(9749) <= not b;
    outputs(9750) <= not (a xor b);
    outputs(9751) <= a;
    outputs(9752) <= not b or a;
    outputs(9753) <= a xor b;
    outputs(9754) <= a xor b;
    outputs(9755) <= not b;
    outputs(9756) <= b;
    outputs(9757) <= a xor b;
    outputs(9758) <= a and not b;
    outputs(9759) <= a and b;
    outputs(9760) <= not (a xor b);
    outputs(9761) <= b;
    outputs(9762) <= a xor b;
    outputs(9763) <= a;
    outputs(9764) <= not b or a;
    outputs(9765) <= a;
    outputs(9766) <= not (a or b);
    outputs(9767) <= a;
    outputs(9768) <= b and not a;
    outputs(9769) <= a and not b;
    outputs(9770) <= not a;
    outputs(9771) <= a and not b;
    outputs(9772) <= a xor b;
    outputs(9773) <= a xor b;
    outputs(9774) <= b;
    outputs(9775) <= a or b;
    outputs(9776) <= not (a or b);
    outputs(9777) <= a and not b;
    outputs(9778) <= not (a xor b);
    outputs(9779) <= not (a xor b);
    outputs(9780) <= b and not a;
    outputs(9781) <= not a;
    outputs(9782) <= a and not b;
    outputs(9783) <= not (a and b);
    outputs(9784) <= not a;
    outputs(9785) <= a or b;
    outputs(9786) <= b;
    outputs(9787) <= a and b;
    outputs(9788) <= not (a or b);
    outputs(9789) <= not b;
    outputs(9790) <= a xor b;
    outputs(9791) <= not (a or b);
    outputs(9792) <= not b;
    outputs(9793) <= a xor b;
    outputs(9794) <= a xor b;
    outputs(9795) <= not b or a;
    outputs(9796) <= b and not a;
    outputs(9797) <= a and b;
    outputs(9798) <= b;
    outputs(9799) <= not b;
    outputs(9800) <= a and b;
    outputs(9801) <= b;
    outputs(9802) <= a and not b;
    outputs(9803) <= not (a xor b);
    outputs(9804) <= a xor b;
    outputs(9805) <= not a;
    outputs(9806) <= not (a xor b);
    outputs(9807) <= not (a or b);
    outputs(9808) <= b and not a;
    outputs(9809) <= b;
    outputs(9810) <= a and b;
    outputs(9811) <= not (a or b);
    outputs(9812) <= a and not b;
    outputs(9813) <= a;
    outputs(9814) <= b;
    outputs(9815) <= not b;
    outputs(9816) <= a and b;
    outputs(9817) <= a and not b;
    outputs(9818) <= b and not a;
    outputs(9819) <= a xor b;
    outputs(9820) <= a and b;
    outputs(9821) <= not b;
    outputs(9822) <= not b;
    outputs(9823) <= not a;
    outputs(9824) <= not (a or b);
    outputs(9825) <= not b or a;
    outputs(9826) <= b and not a;
    outputs(9827) <= a xor b;
    outputs(9828) <= b;
    outputs(9829) <= not (a xor b);
    outputs(9830) <= a;
    outputs(9831) <= not (a xor b);
    outputs(9832) <= not (a xor b);
    outputs(9833) <= not a;
    outputs(9834) <= a;
    outputs(9835) <= b and not a;
    outputs(9836) <= a xor b;
    outputs(9837) <= b and not a;
    outputs(9838) <= a xor b;
    outputs(9839) <= not (a xor b);
    outputs(9840) <= a and not b;
    outputs(9841) <= a or b;
    outputs(9842) <= not (a or b);
    outputs(9843) <= not (a or b);
    outputs(9844) <= b;
    outputs(9845) <= a and not b;
    outputs(9846) <= not b;
    outputs(9847) <= not b or a;
    outputs(9848) <= a and not b;
    outputs(9849) <= not b;
    outputs(9850) <= not (a xor b);
    outputs(9851) <= not (a xor b);
    outputs(9852) <= a and not b;
    outputs(9853) <= a and b;
    outputs(9854) <= b;
    outputs(9855) <= not a;
    outputs(9856) <= a xor b;
    outputs(9857) <= a xor b;
    outputs(9858) <= a and b;
    outputs(9859) <= b;
    outputs(9860) <= a;
    outputs(9861) <= not (a xor b);
    outputs(9862) <= not b;
    outputs(9863) <= not a;
    outputs(9864) <= a and not b;
    outputs(9865) <= a and b;
    outputs(9866) <= a;
    outputs(9867) <= a and not b;
    outputs(9868) <= not a;
    outputs(9869) <= not b;
    outputs(9870) <= not b;
    outputs(9871) <= a xor b;
    outputs(9872) <= a;
    outputs(9873) <= b and not a;
    outputs(9874) <= not b;
    outputs(9875) <= not a;
    outputs(9876) <= not b;
    outputs(9877) <= not (a xor b);
    outputs(9878) <= a and b;
    outputs(9879) <= not a;
    outputs(9880) <= a and not b;
    outputs(9881) <= a;
    outputs(9882) <= a;
    outputs(9883) <= a and b;
    outputs(9884) <= a and b;
    outputs(9885) <= not (a xor b);
    outputs(9886) <= a;
    outputs(9887) <= a;
    outputs(9888) <= a xor b;
    outputs(9889) <= a xor b;
    outputs(9890) <= b and not a;
    outputs(9891) <= not (a xor b);
    outputs(9892) <= b;
    outputs(9893) <= not (a xor b);
    outputs(9894) <= not a or b;
    outputs(9895) <= not (a xor b);
    outputs(9896) <= a xor b;
    outputs(9897) <= not b;
    outputs(9898) <= not a;
    outputs(9899) <= a;
    outputs(9900) <= not (a and b);
    outputs(9901) <= a xor b;
    outputs(9902) <= a;
    outputs(9903) <= b and not a;
    outputs(9904) <= a xor b;
    outputs(9905) <= a and not b;
    outputs(9906) <= a xor b;
    outputs(9907) <= b;
    outputs(9908) <= a and not b;
    outputs(9909) <= not a;
    outputs(9910) <= a;
    outputs(9911) <= not b;
    outputs(9912) <= b;
    outputs(9913) <= a and b;
    outputs(9914) <= not (a or b);
    outputs(9915) <= a;
    outputs(9916) <= a or b;
    outputs(9917) <= not a;
    outputs(9918) <= b and not a;
    outputs(9919) <= not a;
    outputs(9920) <= not (a xor b);
    outputs(9921) <= not b;
    outputs(9922) <= a and not b;
    outputs(9923) <= b;
    outputs(9924) <= not a;
    outputs(9925) <= not (a xor b);
    outputs(9926) <= not a;
    outputs(9927) <= not (a xor b);
    outputs(9928) <= a xor b;
    outputs(9929) <= not (a xor b);
    outputs(9930) <= b and not a;
    outputs(9931) <= a xor b;
    outputs(9932) <= a xor b;
    outputs(9933) <= not a;
    outputs(9934) <= not (a or b);
    outputs(9935) <= a;
    outputs(9936) <= not (a xor b);
    outputs(9937) <= not (a or b);
    outputs(9938) <= not (a xor b);
    outputs(9939) <= not (a xor b);
    outputs(9940) <= a and b;
    outputs(9941) <= a xor b;
    outputs(9942) <= a xor b;
    outputs(9943) <= not (a xor b);
    outputs(9944) <= a;
    outputs(9945) <= b;
    outputs(9946) <= b and not a;
    outputs(9947) <= a and b;
    outputs(9948) <= a xor b;
    outputs(9949) <= not b or a;
    outputs(9950) <= b and not a;
    outputs(9951) <= a and b;
    outputs(9952) <= b;
    outputs(9953) <= a or b;
    outputs(9954) <= not b;
    outputs(9955) <= a xor b;
    outputs(9956) <= a;
    outputs(9957) <= b;
    outputs(9958) <= a or b;
    outputs(9959) <= b and not a;
    outputs(9960) <= not b;
    outputs(9961) <= a xor b;
    outputs(9962) <= not (a or b);
    outputs(9963) <= a or b;
    outputs(9964) <= b;
    outputs(9965) <= a xor b;
    outputs(9966) <= a and b;
    outputs(9967) <= not a;
    outputs(9968) <= not a;
    outputs(9969) <= b and not a;
    outputs(9970) <= a xor b;
    outputs(9971) <= not b;
    outputs(9972) <= a and not b;
    outputs(9973) <= not b or a;
    outputs(9974) <= b;
    outputs(9975) <= not (a or b);
    outputs(9976) <= a and b;
    outputs(9977) <= a and b;
    outputs(9978) <= not b;
    outputs(9979) <= not b or a;
    outputs(9980) <= b and not a;
    outputs(9981) <= a;
    outputs(9982) <= a and b;
    outputs(9983) <= not a;
    outputs(9984) <= not (a xor b);
    outputs(9985) <= not (a or b);
    outputs(9986) <= not a;
    outputs(9987) <= a and not b;
    outputs(9988) <= not b;
    outputs(9989) <= not (a xor b);
    outputs(9990) <= not (a xor b);
    outputs(9991) <= not a;
    outputs(9992) <= not (a xor b);
    outputs(9993) <= not a;
    outputs(9994) <= not (a xor b);
    outputs(9995) <= not b or a;
    outputs(9996) <= not (a xor b);
    outputs(9997) <= not (a xor b);
    outputs(9998) <= a;
    outputs(9999) <= not (a xor b);
    outputs(10000) <= a;
    outputs(10001) <= a and not b;
    outputs(10002) <= not (a xor b);
    outputs(10003) <= a xor b;
    outputs(10004) <= not (a xor b);
    outputs(10005) <= a;
    outputs(10006) <= b and not a;
    outputs(10007) <= b and not a;
    outputs(10008) <= not (a or b);
    outputs(10009) <= not b;
    outputs(10010) <= a xor b;
    outputs(10011) <= a and not b;
    outputs(10012) <= b and not a;
    outputs(10013) <= a;
    outputs(10014) <= a and not b;
    outputs(10015) <= not a;
    outputs(10016) <= not b;
    outputs(10017) <= not (a or b);
    outputs(10018) <= not (a xor b);
    outputs(10019) <= not (a or b);
    outputs(10020) <= a xor b;
    outputs(10021) <= not (a xor b);
    outputs(10022) <= b;
    outputs(10023) <= a and not b;
    outputs(10024) <= b and not a;
    outputs(10025) <= a;
    outputs(10026) <= not a;
    outputs(10027) <= not b or a;
    outputs(10028) <= not a;
    outputs(10029) <= b and not a;
    outputs(10030) <= a and b;
    outputs(10031) <= b;
    outputs(10032) <= a xor b;
    outputs(10033) <= a;
    outputs(10034) <= not b;
    outputs(10035) <= not (a xor b);
    outputs(10036) <= not a;
    outputs(10037) <= not (a xor b);
    outputs(10038) <= not b;
    outputs(10039) <= not b or a;
    outputs(10040) <= not a;
    outputs(10041) <= b and not a;
    outputs(10042) <= not (a or b);
    outputs(10043) <= a and b;
    outputs(10044) <= not (a xor b);
    outputs(10045) <= a and not b;
    outputs(10046) <= a;
    outputs(10047) <= a xor b;
    outputs(10048) <= b;
    outputs(10049) <= not (a xor b);
    outputs(10050) <= a xor b;
    outputs(10051) <= not (a xor b);
    outputs(10052) <= a and b;
    outputs(10053) <= not a;
    outputs(10054) <= a and b;
    outputs(10055) <= not (a xor b);
    outputs(10056) <= not (a xor b);
    outputs(10057) <= b;
    outputs(10058) <= not b;
    outputs(10059) <= not b;
    outputs(10060) <= a or b;
    outputs(10061) <= not a;
    outputs(10062) <= a xor b;
    outputs(10063) <= a xor b;
    outputs(10064) <= a xor b;
    outputs(10065) <= a and not b;
    outputs(10066) <= b;
    outputs(10067) <= b;
    outputs(10068) <= not (a and b);
    outputs(10069) <= a xor b;
    outputs(10070) <= not (a and b);
    outputs(10071) <= b;
    outputs(10072) <= not a;
    outputs(10073) <= a and not b;
    outputs(10074) <= not (a xor b);
    outputs(10075) <= a and not b;
    outputs(10076) <= a xor b;
    outputs(10077) <= not b;
    outputs(10078) <= not b;
    outputs(10079) <= a;
    outputs(10080) <= a xor b;
    outputs(10081) <= a and b;
    outputs(10082) <= not (a or b);
    outputs(10083) <= b and not a;
    outputs(10084) <= not (a or b);
    outputs(10085) <= not (a xor b);
    outputs(10086) <= a xor b;
    outputs(10087) <= not b or a;
    outputs(10088) <= not (a xor b);
    outputs(10089) <= not (a or b);
    outputs(10090) <= b and not a;
    outputs(10091) <= a and not b;
    outputs(10092) <= not b;
    outputs(10093) <= not a;
    outputs(10094) <= a and not b;
    outputs(10095) <= b and not a;
    outputs(10096) <= not b;
    outputs(10097) <= not b;
    outputs(10098) <= not a;
    outputs(10099) <= a xor b;
    outputs(10100) <= a xor b;
    outputs(10101) <= a xor b;
    outputs(10102) <= b;
    outputs(10103) <= b;
    outputs(10104) <= b;
    outputs(10105) <= b;
    outputs(10106) <= b and not a;
    outputs(10107) <= a or b;
    outputs(10108) <= a and b;
    outputs(10109) <= b and not a;
    outputs(10110) <= a xor b;
    outputs(10111) <= not (a or b);
    outputs(10112) <= not b;
    outputs(10113) <= not (a xor b);
    outputs(10114) <= a and not b;
    outputs(10115) <= a or b;
    outputs(10116) <= a;
    outputs(10117) <= a or b;
    outputs(10118) <= b;
    outputs(10119) <= a xor b;
    outputs(10120) <= not (a xor b);
    outputs(10121) <= a and b;
    outputs(10122) <= a xor b;
    outputs(10123) <= a and b;
    outputs(10124) <= a xor b;
    outputs(10125) <= not (a xor b);
    outputs(10126) <= not b;
    outputs(10127) <= a xor b;
    outputs(10128) <= not (a or b);
    outputs(10129) <= a and not b;
    outputs(10130) <= not b;
    outputs(10131) <= not (a xor b);
    outputs(10132) <= a xor b;
    outputs(10133) <= a and b;
    outputs(10134) <= a xor b;
    outputs(10135) <= not (a xor b);
    outputs(10136) <= a xor b;
    outputs(10137) <= b;
    outputs(10138) <= not a;
    outputs(10139) <= a xor b;
    outputs(10140) <= a and b;
    outputs(10141) <= not (a and b);
    outputs(10142) <= a and b;
    outputs(10143) <= b;
    outputs(10144) <= a;
    outputs(10145) <= a xor b;
    outputs(10146) <= b;
    outputs(10147) <= a;
    outputs(10148) <= not a;
    outputs(10149) <= not a or b;
    outputs(10150) <= not b;
    outputs(10151) <= not (a xor b);
    outputs(10152) <= a and not b;
    outputs(10153) <= b;
    outputs(10154) <= a;
    outputs(10155) <= a xor b;
    outputs(10156) <= b;
    outputs(10157) <= not b;
    outputs(10158) <= b and not a;
    outputs(10159) <= a and b;
    outputs(10160) <= not (a or b);
    outputs(10161) <= not b;
    outputs(10162) <= not (a or b);
    outputs(10163) <= not (a xor b);
    outputs(10164) <= a;
    outputs(10165) <= not (a xor b);
    outputs(10166) <= a xor b;
    outputs(10167) <= a xor b;
    outputs(10168) <= a and b;
    outputs(10169) <= b;
    outputs(10170) <= b;
    outputs(10171) <= a and not b;
    outputs(10172) <= not (a xor b);
    outputs(10173) <= not b or a;
    outputs(10174) <= not (a xor b);
    outputs(10175) <= a;
    outputs(10176) <= a xor b;
    outputs(10177) <= a xor b;
    outputs(10178) <= not b;
    outputs(10179) <= a;
    outputs(10180) <= a xor b;
    outputs(10181) <= not (a or b);
    outputs(10182) <= a;
    outputs(10183) <= a;
    outputs(10184) <= not (a xor b);
    outputs(10185) <= not a;
    outputs(10186) <= b;
    outputs(10187) <= b;
    outputs(10188) <= not (a or b);
    outputs(10189) <= not a;
    outputs(10190) <= not a;
    outputs(10191) <= a and b;
    outputs(10192) <= not (a or b);
    outputs(10193) <= not b;
    outputs(10194) <= not b;
    outputs(10195) <= b and not a;
    outputs(10196) <= a and b;
    outputs(10197) <= a xor b;
    outputs(10198) <= not (a xor b);
    outputs(10199) <= not (a xor b);
    outputs(10200) <= b;
    outputs(10201) <= not b;
    outputs(10202) <= not (a xor b);
    outputs(10203) <= a and b;
    outputs(10204) <= '0';
    outputs(10205) <= a;
    outputs(10206) <= not a;
    outputs(10207) <= not a;
    outputs(10208) <= not a;
    outputs(10209) <= a and b;
    outputs(10210) <= a and b;
    outputs(10211) <= not (a xor b);
    outputs(10212) <= not a;
    outputs(10213) <= not (a and b);
    outputs(10214) <= not (a or b);
    outputs(10215) <= not b;
    outputs(10216) <= not (a xor b);
    outputs(10217) <= a and b;
    outputs(10218) <= a and not b;
    outputs(10219) <= b and not a;
    outputs(10220) <= not b;
    outputs(10221) <= a;
    outputs(10222) <= not (a and b);
    outputs(10223) <= a xor b;
    outputs(10224) <= a and not b;
    outputs(10225) <= a and not b;
    outputs(10226) <= a and b;
    outputs(10227) <= a xor b;
    outputs(10228) <= a xor b;
    outputs(10229) <= not (a or b);
    outputs(10230) <= b;
    outputs(10231) <= a and b;
    outputs(10232) <= a and not b;
    outputs(10233) <= a xor b;
    outputs(10234) <= a;
    outputs(10235) <= not b;
    outputs(10236) <= b and not a;
    outputs(10237) <= not (a or b);
    outputs(10238) <= b;
    outputs(10239) <= b and not a;
end Behavioral;
