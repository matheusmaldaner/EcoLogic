library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(2559 downto 0);

begin

    layer0_outputs(0) <= not((inputs(127)) or (inputs(35)));
    layer0_outputs(1) <= (inputs(47)) xor (inputs(21));
    layer0_outputs(2) <= not(inputs(35));
    layer0_outputs(3) <= inputs(141);
    layer0_outputs(4) <= not(inputs(92)) or (inputs(254));
    layer0_outputs(5) <= not((inputs(156)) or (inputs(33)));
    layer0_outputs(6) <= (inputs(242)) or (inputs(140));
    layer0_outputs(7) <= inputs(213);
    layer0_outputs(8) <= (inputs(217)) xor (inputs(249));
    layer0_outputs(9) <= (inputs(241)) and not (inputs(93));
    layer0_outputs(10) <= (inputs(65)) or (inputs(93));
    layer0_outputs(11) <= not((inputs(17)) or (inputs(204)));
    layer0_outputs(12) <= not((inputs(85)) or (inputs(133)));
    layer0_outputs(13) <= not(inputs(26));
    layer0_outputs(14) <= not(inputs(92));
    layer0_outputs(15) <= not(inputs(172)) or (inputs(0));
    layer0_outputs(16) <= not(inputs(183)) or (inputs(102));
    layer0_outputs(17) <= (inputs(53)) or (inputs(225));
    layer0_outputs(18) <= inputs(115);
    layer0_outputs(19) <= not(inputs(176)) or (inputs(100));
    layer0_outputs(20) <= '1';
    layer0_outputs(21) <= not((inputs(95)) xor (inputs(38)));
    layer0_outputs(22) <= not(inputs(119));
    layer0_outputs(23) <= not(inputs(219)) or (inputs(97));
    layer0_outputs(24) <= not(inputs(98));
    layer0_outputs(25) <= not((inputs(68)) or (inputs(12)));
    layer0_outputs(26) <= not(inputs(244)) or (inputs(39));
    layer0_outputs(27) <= not(inputs(56)) or (inputs(0));
    layer0_outputs(28) <= '0';
    layer0_outputs(29) <= inputs(229);
    layer0_outputs(30) <= not(inputs(96));
    layer0_outputs(31) <= '0';
    layer0_outputs(32) <= not(inputs(69));
    layer0_outputs(33) <= not(inputs(172));
    layer0_outputs(34) <= not((inputs(118)) or (inputs(174)));
    layer0_outputs(35) <= not(inputs(114)) or (inputs(65));
    layer0_outputs(36) <= '1';
    layer0_outputs(37) <= (inputs(139)) or (inputs(205));
    layer0_outputs(38) <= not(inputs(69));
    layer0_outputs(39) <= (inputs(183)) and not (inputs(174));
    layer0_outputs(40) <= (inputs(49)) or (inputs(34));
    layer0_outputs(41) <= inputs(52);
    layer0_outputs(42) <= not(inputs(70));
    layer0_outputs(43) <= not(inputs(163));
    layer0_outputs(44) <= not(inputs(146)) or (inputs(93));
    layer0_outputs(45) <= not((inputs(91)) or (inputs(65)));
    layer0_outputs(46) <= not(inputs(244));
    layer0_outputs(47) <= not(inputs(107));
    layer0_outputs(48) <= not(inputs(51));
    layer0_outputs(49) <= (inputs(21)) or (inputs(86));
    layer0_outputs(50) <= inputs(183);
    layer0_outputs(51) <= not((inputs(87)) or (inputs(85)));
    layer0_outputs(52) <= '0';
    layer0_outputs(53) <= (inputs(211)) or (inputs(16));
    layer0_outputs(54) <= (inputs(226)) or (inputs(225));
    layer0_outputs(55) <= not(inputs(138));
    layer0_outputs(56) <= (inputs(195)) or (inputs(20));
    layer0_outputs(57) <= inputs(173);
    layer0_outputs(58) <= inputs(162);
    layer0_outputs(59) <= inputs(149);
    layer0_outputs(60) <= (inputs(43)) and not (inputs(246));
    layer0_outputs(61) <= not(inputs(166)) or (inputs(172));
    layer0_outputs(62) <= not(inputs(140)) or (inputs(147));
    layer0_outputs(63) <= not((inputs(13)) or (inputs(21)));
    layer0_outputs(64) <= '0';
    layer0_outputs(65) <= not((inputs(82)) or (inputs(86)));
    layer0_outputs(66) <= (inputs(26)) and not (inputs(175));
    layer0_outputs(67) <= (inputs(117)) or (inputs(248));
    layer0_outputs(68) <= (inputs(250)) or (inputs(229));
    layer0_outputs(69) <= not(inputs(120));
    layer0_outputs(70) <= (inputs(42)) and not (inputs(252));
    layer0_outputs(71) <= not((inputs(138)) or (inputs(7)));
    layer0_outputs(72) <= (inputs(108)) or (inputs(121));
    layer0_outputs(73) <= not((inputs(82)) or (inputs(194)));
    layer0_outputs(74) <= (inputs(57)) and not (inputs(58));
    layer0_outputs(75) <= (inputs(201)) or (inputs(116));
    layer0_outputs(76) <= not((inputs(107)) or (inputs(12)));
    layer0_outputs(77) <= '0';
    layer0_outputs(78) <= not((inputs(17)) or (inputs(90)));
    layer0_outputs(79) <= (inputs(220)) and not (inputs(249));
    layer0_outputs(80) <= inputs(25);
    layer0_outputs(81) <= inputs(181);
    layer0_outputs(82) <= not(inputs(131)) or (inputs(48));
    layer0_outputs(83) <= (inputs(213)) or (inputs(173));
    layer0_outputs(84) <= (inputs(18)) and not (inputs(185));
    layer0_outputs(85) <= not(inputs(105));
    layer0_outputs(86) <= not(inputs(167));
    layer0_outputs(87) <= not(inputs(232));
    layer0_outputs(88) <= not(inputs(99));
    layer0_outputs(89) <= (inputs(177)) or (inputs(176));
    layer0_outputs(90) <= (inputs(86)) or (inputs(129));
    layer0_outputs(91) <= inputs(179);
    layer0_outputs(92) <= not(inputs(136)) or (inputs(79));
    layer0_outputs(93) <= (inputs(2)) and not (inputs(13));
    layer0_outputs(94) <= not((inputs(242)) or (inputs(89)));
    layer0_outputs(95) <= not((inputs(207)) or (inputs(37)));
    layer0_outputs(96) <= (inputs(157)) or (inputs(227));
    layer0_outputs(97) <= not((inputs(142)) and (inputs(174)));
    layer0_outputs(98) <= inputs(215);
    layer0_outputs(99) <= (inputs(40)) and not (inputs(127));
    layer0_outputs(100) <= not(inputs(70));
    layer0_outputs(101) <= not(inputs(230));
    layer0_outputs(102) <= (inputs(171)) xor (inputs(0));
    layer0_outputs(103) <= (inputs(172)) and not (inputs(253));
    layer0_outputs(104) <= inputs(90);
    layer0_outputs(105) <= inputs(221);
    layer0_outputs(106) <= (inputs(193)) or (inputs(248));
    layer0_outputs(107) <= not(inputs(176)) or (inputs(42));
    layer0_outputs(108) <= (inputs(110)) xor (inputs(135));
    layer0_outputs(109) <= '0';
    layer0_outputs(110) <= (inputs(101)) or (inputs(146));
    layer0_outputs(111) <= (inputs(84)) and not (inputs(110));
    layer0_outputs(112) <= not((inputs(244)) or (inputs(32)));
    layer0_outputs(113) <= not((inputs(188)) xor (inputs(137)));
    layer0_outputs(114) <= inputs(248);
    layer0_outputs(115) <= (inputs(139)) or (inputs(123));
    layer0_outputs(116) <= not(inputs(122));
    layer0_outputs(117) <= inputs(84);
    layer0_outputs(118) <= (inputs(210)) or (inputs(9));
    layer0_outputs(119) <= not(inputs(165));
    layer0_outputs(120) <= (inputs(127)) and not (inputs(57));
    layer0_outputs(121) <= inputs(133);
    layer0_outputs(122) <= inputs(74);
    layer0_outputs(123) <= '1';
    layer0_outputs(124) <= inputs(220);
    layer0_outputs(125) <= (inputs(174)) or (inputs(20));
    layer0_outputs(126) <= '0';
    layer0_outputs(127) <= not((inputs(218)) or (inputs(165)));
    layer0_outputs(128) <= (inputs(154)) or (inputs(110));
    layer0_outputs(129) <= (inputs(174)) or (inputs(180));
    layer0_outputs(130) <= not((inputs(158)) or (inputs(240)));
    layer0_outputs(131) <= not(inputs(240));
    layer0_outputs(132) <= '1';
    layer0_outputs(133) <= inputs(149);
    layer0_outputs(134) <= not(inputs(116));
    layer0_outputs(135) <= not(inputs(224));
    layer0_outputs(136) <= (inputs(195)) or (inputs(69));
    layer0_outputs(137) <= (inputs(39)) or (inputs(45));
    layer0_outputs(138) <= not((inputs(244)) xor (inputs(197)));
    layer0_outputs(139) <= not(inputs(152)) or (inputs(56));
    layer0_outputs(140) <= (inputs(225)) or (inputs(23));
    layer0_outputs(141) <= (inputs(24)) and (inputs(199));
    layer0_outputs(142) <= not(inputs(245)) or (inputs(94));
    layer0_outputs(143) <= (inputs(37)) or (inputs(210));
    layer0_outputs(144) <= not(inputs(99));
    layer0_outputs(145) <= not((inputs(168)) or (inputs(254)));
    layer0_outputs(146) <= inputs(179);
    layer0_outputs(147) <= not((inputs(234)) or (inputs(140)));
    layer0_outputs(148) <= not(inputs(82)) or (inputs(60));
    layer0_outputs(149) <= not(inputs(103)) or (inputs(111));
    layer0_outputs(150) <= inputs(26);
    layer0_outputs(151) <= (inputs(198)) and not (inputs(146));
    layer0_outputs(152) <= not((inputs(239)) or (inputs(20)));
    layer0_outputs(153) <= not((inputs(45)) or (inputs(43)));
    layer0_outputs(154) <= (inputs(73)) or (inputs(72));
    layer0_outputs(155) <= not(inputs(10));
    layer0_outputs(156) <= (inputs(150)) or (inputs(88));
    layer0_outputs(157) <= not(inputs(248));
    layer0_outputs(158) <= inputs(195);
    layer0_outputs(159) <= (inputs(165)) or (inputs(197));
    layer0_outputs(160) <= inputs(231);
    layer0_outputs(161) <= (inputs(62)) or (inputs(87));
    layer0_outputs(162) <= not(inputs(174));
    layer0_outputs(163) <= not(inputs(247));
    layer0_outputs(164) <= (inputs(118)) or (inputs(175));
    layer0_outputs(165) <= not((inputs(112)) or (inputs(185)));
    layer0_outputs(166) <= not(inputs(25)) or (inputs(157));
    layer0_outputs(167) <= not(inputs(84));
    layer0_outputs(168) <= not((inputs(46)) or (inputs(90)));
    layer0_outputs(169) <= inputs(143);
    layer0_outputs(170) <= (inputs(26)) and (inputs(199));
    layer0_outputs(171) <= (inputs(84)) or (inputs(10));
    layer0_outputs(172) <= inputs(133);
    layer0_outputs(173) <= (inputs(207)) and not (inputs(160));
    layer0_outputs(174) <= (inputs(159)) and not (inputs(71));
    layer0_outputs(175) <= inputs(93);
    layer0_outputs(176) <= not((inputs(85)) xor (inputs(54)));
    layer0_outputs(177) <= not(inputs(152));
    layer0_outputs(178) <= not(inputs(98));
    layer0_outputs(179) <= (inputs(60)) and not (inputs(176));
    layer0_outputs(180) <= (inputs(196)) or (inputs(209));
    layer0_outputs(181) <= '0';
    layer0_outputs(182) <= not((inputs(200)) or (inputs(95)));
    layer0_outputs(183) <= (inputs(2)) and not (inputs(107));
    layer0_outputs(184) <= not(inputs(126));
    layer0_outputs(185) <= (inputs(224)) or (inputs(207));
    layer0_outputs(186) <= not((inputs(163)) or (inputs(254)));
    layer0_outputs(187) <= (inputs(245)) and not (inputs(2));
    layer0_outputs(188) <= not((inputs(219)) or (inputs(143)));
    layer0_outputs(189) <= inputs(79);
    layer0_outputs(190) <= (inputs(139)) or (inputs(239));
    layer0_outputs(191) <= (inputs(3)) and not (inputs(239));
    layer0_outputs(192) <= not((inputs(31)) xor (inputs(12)));
    layer0_outputs(193) <= not(inputs(113));
    layer0_outputs(194) <= not((inputs(172)) or (inputs(159)));
    layer0_outputs(195) <= not(inputs(167)) or (inputs(118));
    layer0_outputs(196) <= (inputs(73)) and (inputs(231));
    layer0_outputs(197) <= not((inputs(218)) or (inputs(155)));
    layer0_outputs(198) <= inputs(90);
    layer0_outputs(199) <= inputs(217);
    layer0_outputs(200) <= not(inputs(126));
    layer0_outputs(201) <= not(inputs(141));
    layer0_outputs(202) <= inputs(62);
    layer0_outputs(203) <= not(inputs(182));
    layer0_outputs(204) <= inputs(245);
    layer0_outputs(205) <= (inputs(116)) and (inputs(152));
    layer0_outputs(206) <= inputs(198);
    layer0_outputs(207) <= inputs(74);
    layer0_outputs(208) <= (inputs(50)) and not (inputs(30));
    layer0_outputs(209) <= inputs(27);
    layer0_outputs(210) <= inputs(78);
    layer0_outputs(211) <= not(inputs(231));
    layer0_outputs(212) <= not(inputs(178));
    layer0_outputs(213) <= not(inputs(25));
    layer0_outputs(214) <= not(inputs(229));
    layer0_outputs(215) <= not(inputs(143));
    layer0_outputs(216) <= inputs(75);
    layer0_outputs(217) <= not(inputs(60)) or (inputs(105));
    layer0_outputs(218) <= not((inputs(192)) or (inputs(236)));
    layer0_outputs(219) <= not(inputs(221));
    layer0_outputs(220) <= not(inputs(89)) or (inputs(130));
    layer0_outputs(221) <= (inputs(56)) and not (inputs(49));
    layer0_outputs(222) <= not(inputs(185));
    layer0_outputs(223) <= (inputs(181)) or (inputs(210));
    layer0_outputs(224) <= inputs(121);
    layer0_outputs(225) <= not(inputs(104)) or (inputs(224));
    layer0_outputs(226) <= inputs(31);
    layer0_outputs(227) <= inputs(118);
    layer0_outputs(228) <= not((inputs(17)) and (inputs(156)));
    layer0_outputs(229) <= not((inputs(106)) or (inputs(3)));
    layer0_outputs(230) <= (inputs(223)) and not (inputs(14));
    layer0_outputs(231) <= not(inputs(206));
    layer0_outputs(232) <= inputs(114);
    layer0_outputs(233) <= not(inputs(221)) or (inputs(11));
    layer0_outputs(234) <= inputs(126);
    layer0_outputs(235) <= inputs(129);
    layer0_outputs(236) <= inputs(137);
    layer0_outputs(237) <= (inputs(234)) or (inputs(84));
    layer0_outputs(238) <= not(inputs(184));
    layer0_outputs(239) <= (inputs(39)) and not (inputs(172));
    layer0_outputs(240) <= not((inputs(144)) or (inputs(159)));
    layer0_outputs(241) <= not(inputs(51)) or (inputs(253));
    layer0_outputs(242) <= not(inputs(152)) or (inputs(220));
    layer0_outputs(243) <= inputs(226);
    layer0_outputs(244) <= inputs(69);
    layer0_outputs(245) <= inputs(18);
    layer0_outputs(246) <= (inputs(152)) xor (inputs(153));
    layer0_outputs(247) <= not(inputs(91)) or (inputs(123));
    layer0_outputs(248) <= not(inputs(28));
    layer0_outputs(249) <= not(inputs(247));
    layer0_outputs(250) <= not((inputs(234)) xor (inputs(185)));
    layer0_outputs(251) <= inputs(182);
    layer0_outputs(252) <= inputs(106);
    layer0_outputs(253) <= inputs(191);
    layer0_outputs(254) <= not((inputs(68)) or (inputs(166)));
    layer0_outputs(255) <= not(inputs(118));
    layer0_outputs(256) <= not((inputs(152)) or (inputs(244)));
    layer0_outputs(257) <= not((inputs(248)) or (inputs(101)));
    layer0_outputs(258) <= (inputs(252)) and not (inputs(145));
    layer0_outputs(259) <= (inputs(17)) or (inputs(164));
    layer0_outputs(260) <= (inputs(177)) and not (inputs(199));
    layer0_outputs(261) <= inputs(243);
    layer0_outputs(262) <= inputs(219);
    layer0_outputs(263) <= not(inputs(52));
    layer0_outputs(264) <= (inputs(240)) xor (inputs(34));
    layer0_outputs(265) <= not((inputs(178)) or (inputs(7)));
    layer0_outputs(266) <= '0';
    layer0_outputs(267) <= (inputs(232)) and not (inputs(127));
    layer0_outputs(268) <= inputs(38);
    layer0_outputs(269) <= (inputs(54)) and (inputs(136));
    layer0_outputs(270) <= not(inputs(83));
    layer0_outputs(271) <= (inputs(62)) or (inputs(7));
    layer0_outputs(272) <= not((inputs(153)) and (inputs(224)));
    layer0_outputs(273) <= (inputs(58)) and not (inputs(63));
    layer0_outputs(274) <= not((inputs(129)) or (inputs(189)));
    layer0_outputs(275) <= inputs(206);
    layer0_outputs(276) <= (inputs(28)) or (inputs(198));
    layer0_outputs(277) <= inputs(166);
    layer0_outputs(278) <= not(inputs(194));
    layer0_outputs(279) <= inputs(23);
    layer0_outputs(280) <= (inputs(182)) or (inputs(14));
    layer0_outputs(281) <= not(inputs(122));
    layer0_outputs(282) <= not(inputs(231));
    layer0_outputs(283) <= not((inputs(52)) or (inputs(219)));
    layer0_outputs(284) <= inputs(170);
    layer0_outputs(285) <= inputs(34);
    layer0_outputs(286) <= (inputs(72)) and (inputs(72));
    layer0_outputs(287) <= not(inputs(44)) or (inputs(131));
    layer0_outputs(288) <= '1';
    layer0_outputs(289) <= inputs(131);
    layer0_outputs(290) <= (inputs(196)) and not (inputs(34));
    layer0_outputs(291) <= not((inputs(214)) or (inputs(148)));
    layer0_outputs(292) <= inputs(182);
    layer0_outputs(293) <= not((inputs(39)) or (inputs(254)));
    layer0_outputs(294) <= not(inputs(188));
    layer0_outputs(295) <= (inputs(32)) and (inputs(17));
    layer0_outputs(296) <= not(inputs(157));
    layer0_outputs(297) <= not((inputs(208)) or (inputs(55)));
    layer0_outputs(298) <= (inputs(228)) or (inputs(42));
    layer0_outputs(299) <= not(inputs(146));
    layer0_outputs(300) <= inputs(154);
    layer0_outputs(301) <= not(inputs(101));
    layer0_outputs(302) <= not((inputs(99)) or (inputs(101)));
    layer0_outputs(303) <= not((inputs(122)) xor (inputs(177)));
    layer0_outputs(304) <= not(inputs(183));
    layer0_outputs(305) <= not(inputs(188)) or (inputs(95));
    layer0_outputs(306) <= not((inputs(55)) or (inputs(17)));
    layer0_outputs(307) <= (inputs(105)) or (inputs(19));
    layer0_outputs(308) <= inputs(135);
    layer0_outputs(309) <= inputs(140);
    layer0_outputs(310) <= not(inputs(36)) or (inputs(126));
    layer0_outputs(311) <= inputs(77);
    layer0_outputs(312) <= not(inputs(183)) or (inputs(209));
    layer0_outputs(313) <= inputs(213);
    layer0_outputs(314) <= not(inputs(100));
    layer0_outputs(315) <= not((inputs(219)) and (inputs(147)));
    layer0_outputs(316) <= (inputs(88)) and not (inputs(114));
    layer0_outputs(317) <= not(inputs(138));
    layer0_outputs(318) <= (inputs(235)) and not (inputs(175));
    layer0_outputs(319) <= (inputs(56)) and not (inputs(180));
    layer0_outputs(320) <= (inputs(124)) or (inputs(74));
    layer0_outputs(321) <= inputs(194);
    layer0_outputs(322) <= (inputs(248)) and not (inputs(5));
    layer0_outputs(323) <= (inputs(203)) xor (inputs(230));
    layer0_outputs(324) <= inputs(98);
    layer0_outputs(325) <= inputs(212);
    layer0_outputs(326) <= (inputs(113)) or (inputs(133));
    layer0_outputs(327) <= not(inputs(246)) or (inputs(215));
    layer0_outputs(328) <= not(inputs(203));
    layer0_outputs(329) <= (inputs(69)) or (inputs(35));
    layer0_outputs(330) <= not(inputs(71)) or (inputs(2));
    layer0_outputs(331) <= (inputs(244)) or (inputs(148));
    layer0_outputs(332) <= not(inputs(2));
    layer0_outputs(333) <= not(inputs(58)) or (inputs(52));
    layer0_outputs(334) <= inputs(38);
    layer0_outputs(335) <= (inputs(162)) or (inputs(234));
    layer0_outputs(336) <= not(inputs(85)) or (inputs(16));
    layer0_outputs(337) <= not((inputs(128)) or (inputs(188)));
    layer0_outputs(338) <= not(inputs(111)) or (inputs(239));
    layer0_outputs(339) <= (inputs(18)) or (inputs(131));
    layer0_outputs(340) <= not((inputs(117)) and (inputs(29)));
    layer0_outputs(341) <= not(inputs(169));
    layer0_outputs(342) <= not((inputs(20)) or (inputs(19)));
    layer0_outputs(343) <= not(inputs(215)) or (inputs(156));
    layer0_outputs(344) <= not(inputs(161));
    layer0_outputs(345) <= (inputs(117)) and not (inputs(221));
    layer0_outputs(346) <= (inputs(120)) and not (inputs(2));
    layer0_outputs(347) <= not(inputs(156)) or (inputs(53));
    layer0_outputs(348) <= not(inputs(132)) or (inputs(1));
    layer0_outputs(349) <= inputs(165);
    layer0_outputs(350) <= inputs(53);
    layer0_outputs(351) <= (inputs(171)) and not (inputs(46));
    layer0_outputs(352) <= not(inputs(40)) or (inputs(155));
    layer0_outputs(353) <= not((inputs(238)) or (inputs(179)));
    layer0_outputs(354) <= not(inputs(105));
    layer0_outputs(355) <= not(inputs(204)) or (inputs(61));
    layer0_outputs(356) <= inputs(55);
    layer0_outputs(357) <= not((inputs(56)) or (inputs(30)));
    layer0_outputs(358) <= (inputs(252)) or (inputs(8));
    layer0_outputs(359) <= not((inputs(27)) xor (inputs(64)));
    layer0_outputs(360) <= not(inputs(23)) or (inputs(28));
    layer0_outputs(361) <= not(inputs(166));
    layer0_outputs(362) <= inputs(203);
    layer0_outputs(363) <= not(inputs(154));
    layer0_outputs(364) <= (inputs(44)) or (inputs(217));
    layer0_outputs(365) <= (inputs(92)) and not (inputs(225));
    layer0_outputs(366) <= '1';
    layer0_outputs(367) <= not(inputs(92));
    layer0_outputs(368) <= inputs(114);
    layer0_outputs(369) <= inputs(196);
    layer0_outputs(370) <= not(inputs(193));
    layer0_outputs(371) <= '0';
    layer0_outputs(372) <= (inputs(252)) or (inputs(36));
    layer0_outputs(373) <= not((inputs(218)) or (inputs(94)));
    layer0_outputs(374) <= inputs(196);
    layer0_outputs(375) <= '0';
    layer0_outputs(376) <= not(inputs(93));
    layer0_outputs(377) <= not((inputs(171)) or (inputs(222)));
    layer0_outputs(378) <= not(inputs(68)) or (inputs(32));
    layer0_outputs(379) <= not((inputs(5)) or (inputs(237)));
    layer0_outputs(380) <= not(inputs(133));
    layer0_outputs(381) <= not(inputs(77));
    layer0_outputs(382) <= not(inputs(157));
    layer0_outputs(383) <= inputs(48);
    layer0_outputs(384) <= (inputs(10)) and not (inputs(225));
    layer0_outputs(385) <= (inputs(143)) or (inputs(204));
    layer0_outputs(386) <= not(inputs(115));
    layer0_outputs(387) <= (inputs(169)) or (inputs(82));
    layer0_outputs(388) <= '1';
    layer0_outputs(389) <= (inputs(189)) or (inputs(37));
    layer0_outputs(390) <= inputs(229);
    layer0_outputs(391) <= not(inputs(247));
    layer0_outputs(392) <= not(inputs(152)) or (inputs(102));
    layer0_outputs(393) <= inputs(250);
    layer0_outputs(394) <= inputs(164);
    layer0_outputs(395) <= not(inputs(209));
    layer0_outputs(396) <= (inputs(225)) xor (inputs(0));
    layer0_outputs(397) <= not(inputs(154));
    layer0_outputs(398) <= inputs(62);
    layer0_outputs(399) <= not(inputs(146));
    layer0_outputs(400) <= '1';
    layer0_outputs(401) <= (inputs(28)) xor (inputs(59));
    layer0_outputs(402) <= (inputs(153)) and not (inputs(46));
    layer0_outputs(403) <= (inputs(67)) or (inputs(109));
    layer0_outputs(404) <= not(inputs(5)) or (inputs(129));
    layer0_outputs(405) <= (inputs(157)) and not (inputs(186));
    layer0_outputs(406) <= inputs(8);
    layer0_outputs(407) <= not(inputs(133));
    layer0_outputs(408) <= (inputs(57)) or (inputs(40));
    layer0_outputs(409) <= not(inputs(135)) or (inputs(50));
    layer0_outputs(410) <= not(inputs(53)) or (inputs(2));
    layer0_outputs(411) <= (inputs(238)) or (inputs(213));
    layer0_outputs(412) <= inputs(8);
    layer0_outputs(413) <= not(inputs(106));
    layer0_outputs(414) <= not(inputs(221));
    layer0_outputs(415) <= not(inputs(237)) or (inputs(171));
    layer0_outputs(416) <= not(inputs(89)) or (inputs(66));
    layer0_outputs(417) <= inputs(206);
    layer0_outputs(418) <= inputs(21);
    layer0_outputs(419) <= (inputs(126)) or (inputs(162));
    layer0_outputs(420) <= not((inputs(13)) or (inputs(137)));
    layer0_outputs(421) <= (inputs(239)) or (inputs(120));
    layer0_outputs(422) <= (inputs(142)) and not (inputs(255));
    layer0_outputs(423) <= not(inputs(151));
    layer0_outputs(424) <= inputs(133);
    layer0_outputs(425) <= inputs(41);
    layer0_outputs(426) <= not(inputs(228)) or (inputs(156));
    layer0_outputs(427) <= not(inputs(220)) or (inputs(58));
    layer0_outputs(428) <= inputs(77);
    layer0_outputs(429) <= not(inputs(148));
    layer0_outputs(430) <= not((inputs(48)) or (inputs(192)));
    layer0_outputs(431) <= (inputs(66)) or (inputs(55));
    layer0_outputs(432) <= inputs(162);
    layer0_outputs(433) <= not((inputs(114)) or (inputs(194)));
    layer0_outputs(434) <= (inputs(235)) or (inputs(186));
    layer0_outputs(435) <= not(inputs(100));
    layer0_outputs(436) <= not((inputs(98)) or (inputs(158)));
    layer0_outputs(437) <= (inputs(30)) or (inputs(205));
    layer0_outputs(438) <= inputs(115);
    layer0_outputs(439) <= not((inputs(50)) xor (inputs(111)));
    layer0_outputs(440) <= not(inputs(22));
    layer0_outputs(441) <= (inputs(59)) or (inputs(194));
    layer0_outputs(442) <= not(inputs(96)) or (inputs(188));
    layer0_outputs(443) <= inputs(212);
    layer0_outputs(444) <= not(inputs(217)) or (inputs(19));
    layer0_outputs(445) <= (inputs(148)) and not (inputs(118));
    layer0_outputs(446) <= not(inputs(98));
    layer0_outputs(447) <= (inputs(21)) and not (inputs(55));
    layer0_outputs(448) <= not((inputs(130)) or (inputs(63)));
    layer0_outputs(449) <= (inputs(25)) and not (inputs(222));
    layer0_outputs(450) <= not(inputs(178));
    layer0_outputs(451) <= not(inputs(227));
    layer0_outputs(452) <= (inputs(148)) and not (inputs(142));
    layer0_outputs(453) <= '1';
    layer0_outputs(454) <= (inputs(181)) and not (inputs(241));
    layer0_outputs(455) <= not(inputs(88));
    layer0_outputs(456) <= not(inputs(60)) or (inputs(222));
    layer0_outputs(457) <= not((inputs(69)) or (inputs(159)));
    layer0_outputs(458) <= (inputs(36)) and (inputs(41));
    layer0_outputs(459) <= not((inputs(193)) or (inputs(174)));
    layer0_outputs(460) <= inputs(21);
    layer0_outputs(461) <= not(inputs(169)) or (inputs(92));
    layer0_outputs(462) <= not(inputs(37));
    layer0_outputs(463) <= inputs(30);
    layer0_outputs(464) <= not(inputs(131));
    layer0_outputs(465) <= (inputs(80)) and not (inputs(158));
    layer0_outputs(466) <= not((inputs(79)) or (inputs(138)));
    layer0_outputs(467) <= inputs(168);
    layer0_outputs(468) <= not((inputs(176)) or (inputs(90)));
    layer0_outputs(469) <= inputs(93);
    layer0_outputs(470) <= inputs(47);
    layer0_outputs(471) <= (inputs(115)) or (inputs(160));
    layer0_outputs(472) <= (inputs(19)) or (inputs(79));
    layer0_outputs(473) <= not(inputs(57)) or (inputs(14));
    layer0_outputs(474) <= not(inputs(43));
    layer0_outputs(475) <= not(inputs(61));
    layer0_outputs(476) <= not(inputs(28));
    layer0_outputs(477) <= not(inputs(83)) or (inputs(175));
    layer0_outputs(478) <= not(inputs(110));
    layer0_outputs(479) <= (inputs(32)) or (inputs(221));
    layer0_outputs(480) <= inputs(208);
    layer0_outputs(481) <= not(inputs(144)) or (inputs(255));
    layer0_outputs(482) <= inputs(127);
    layer0_outputs(483) <= inputs(17);
    layer0_outputs(484) <= not((inputs(112)) or (inputs(178)));
    layer0_outputs(485) <= inputs(176);
    layer0_outputs(486) <= not(inputs(240));
    layer0_outputs(487) <= inputs(175);
    layer0_outputs(488) <= inputs(94);
    layer0_outputs(489) <= (inputs(25)) and not (inputs(97));
    layer0_outputs(490) <= inputs(20);
    layer0_outputs(491) <= (inputs(61)) or (inputs(91));
    layer0_outputs(492) <= '1';
    layer0_outputs(493) <= not((inputs(30)) or (inputs(113)));
    layer0_outputs(494) <= inputs(25);
    layer0_outputs(495) <= not((inputs(99)) or (inputs(98)));
    layer0_outputs(496) <= not((inputs(215)) or (inputs(191)));
    layer0_outputs(497) <= not((inputs(120)) xor (inputs(124)));
    layer0_outputs(498) <= not((inputs(189)) and (inputs(54)));
    layer0_outputs(499) <= inputs(15);
    layer0_outputs(500) <= not(inputs(5)) or (inputs(112));
    layer0_outputs(501) <= inputs(203);
    layer0_outputs(502) <= not(inputs(125)) or (inputs(109));
    layer0_outputs(503) <= not(inputs(86)) or (inputs(254));
    layer0_outputs(504) <= not(inputs(90));
    layer0_outputs(505) <= (inputs(210)) or (inputs(238));
    layer0_outputs(506) <= inputs(43);
    layer0_outputs(507) <= not(inputs(22));
    layer0_outputs(508) <= not((inputs(83)) and (inputs(236)));
    layer0_outputs(509) <= not(inputs(68));
    layer0_outputs(510) <= (inputs(71)) or (inputs(4));
    layer0_outputs(511) <= not(inputs(117));
    layer0_outputs(512) <= not((inputs(175)) or (inputs(59)));
    layer0_outputs(513) <= not(inputs(116));
    layer0_outputs(514) <= not((inputs(176)) or (inputs(216)));
    layer0_outputs(515) <= (inputs(191)) or (inputs(171));
    layer0_outputs(516) <= (inputs(172)) or (inputs(161));
    layer0_outputs(517) <= not((inputs(128)) and (inputs(81)));
    layer0_outputs(518) <= inputs(167);
    layer0_outputs(519) <= not(inputs(59));
    layer0_outputs(520) <= not(inputs(60));
    layer0_outputs(521) <= not(inputs(14)) or (inputs(63));
    layer0_outputs(522) <= not(inputs(22));
    layer0_outputs(523) <= (inputs(55)) or (inputs(30));
    layer0_outputs(524) <= not(inputs(39));
    layer0_outputs(525) <= inputs(210);
    layer0_outputs(526) <= (inputs(200)) or (inputs(131));
    layer0_outputs(527) <= not(inputs(14));
    layer0_outputs(528) <= not((inputs(79)) or (inputs(222)));
    layer0_outputs(529) <= inputs(78);
    layer0_outputs(530) <= not(inputs(132)) or (inputs(33));
    layer0_outputs(531) <= not(inputs(103));
    layer0_outputs(532) <= not(inputs(230));
    layer0_outputs(533) <= (inputs(184)) and not (inputs(79));
    layer0_outputs(534) <= inputs(255);
    layer0_outputs(535) <= not(inputs(235));
    layer0_outputs(536) <= not(inputs(91)) or (inputs(161));
    layer0_outputs(537) <= not((inputs(193)) or (inputs(51)));
    layer0_outputs(538) <= not((inputs(77)) or (inputs(3)));
    layer0_outputs(539) <= (inputs(158)) xor (inputs(134));
    layer0_outputs(540) <= inputs(160);
    layer0_outputs(541) <= not((inputs(183)) or (inputs(241)));
    layer0_outputs(542) <= inputs(123);
    layer0_outputs(543) <= '1';
    layer0_outputs(544) <= inputs(8);
    layer0_outputs(545) <= (inputs(6)) xor (inputs(51));
    layer0_outputs(546) <= not(inputs(209));
    layer0_outputs(547) <= (inputs(103)) and not (inputs(51));
    layer0_outputs(548) <= inputs(99);
    layer0_outputs(549) <= not((inputs(251)) or (inputs(133)));
    layer0_outputs(550) <= not(inputs(136)) or (inputs(205));
    layer0_outputs(551) <= not(inputs(136)) or (inputs(23));
    layer0_outputs(552) <= inputs(183);
    layer0_outputs(553) <= (inputs(184)) and (inputs(155));
    layer0_outputs(554) <= not((inputs(66)) or (inputs(25)));
    layer0_outputs(555) <= not((inputs(180)) or (inputs(46)));
    layer0_outputs(556) <= (inputs(78)) or (inputs(45));
    layer0_outputs(557) <= not(inputs(26));
    layer0_outputs(558) <= not(inputs(27));
    layer0_outputs(559) <= not((inputs(205)) or (inputs(18)));
    layer0_outputs(560) <= not(inputs(250));
    layer0_outputs(561) <= not(inputs(132)) or (inputs(192));
    layer0_outputs(562) <= (inputs(223)) and not (inputs(33));
    layer0_outputs(563) <= (inputs(137)) and not (inputs(246));
    layer0_outputs(564) <= not(inputs(150));
    layer0_outputs(565) <= inputs(167);
    layer0_outputs(566) <= '1';
    layer0_outputs(567) <= (inputs(139)) or (inputs(253));
    layer0_outputs(568) <= not(inputs(209)) or (inputs(237));
    layer0_outputs(569) <= not(inputs(233));
    layer0_outputs(570) <= not((inputs(204)) or (inputs(187)));
    layer0_outputs(571) <= (inputs(172)) and not (inputs(162));
    layer0_outputs(572) <= not((inputs(226)) or (inputs(206)));
    layer0_outputs(573) <= inputs(246);
    layer0_outputs(574) <= (inputs(137)) and not (inputs(172));
    layer0_outputs(575) <= (inputs(151)) xor (inputs(166));
    layer0_outputs(576) <= not(inputs(105));
    layer0_outputs(577) <= inputs(157);
    layer0_outputs(578) <= not((inputs(45)) and (inputs(152)));
    layer0_outputs(579) <= (inputs(109)) or (inputs(190));
    layer0_outputs(580) <= not((inputs(16)) and (inputs(234)));
    layer0_outputs(581) <= not(inputs(158));
    layer0_outputs(582) <= not(inputs(75));
    layer0_outputs(583) <= inputs(212);
    layer0_outputs(584) <= inputs(163);
    layer0_outputs(585) <= not(inputs(232));
    layer0_outputs(586) <= (inputs(239)) and not (inputs(16));
    layer0_outputs(587) <= not(inputs(29)) or (inputs(216));
    layer0_outputs(588) <= not(inputs(91));
    layer0_outputs(589) <= (inputs(204)) or (inputs(192));
    layer0_outputs(590) <= not((inputs(176)) or (inputs(202)));
    layer0_outputs(591) <= (inputs(16)) and (inputs(5));
    layer0_outputs(592) <= (inputs(254)) or (inputs(126));
    layer0_outputs(593) <= not((inputs(51)) and (inputs(51)));
    layer0_outputs(594) <= not((inputs(46)) or (inputs(241)));
    layer0_outputs(595) <= not(inputs(97));
    layer0_outputs(596) <= not((inputs(170)) or (inputs(223)));
    layer0_outputs(597) <= inputs(129);
    layer0_outputs(598) <= (inputs(205)) or (inputs(176));
    layer0_outputs(599) <= inputs(120);
    layer0_outputs(600) <= (inputs(85)) or (inputs(131));
    layer0_outputs(601) <= inputs(23);
    layer0_outputs(602) <= not(inputs(127));
    layer0_outputs(603) <= (inputs(55)) and not (inputs(62));
    layer0_outputs(604) <= not(inputs(101));
    layer0_outputs(605) <= not(inputs(40));
    layer0_outputs(606) <= (inputs(102)) and not (inputs(32));
    layer0_outputs(607) <= (inputs(156)) and not (inputs(1));
    layer0_outputs(608) <= (inputs(137)) and not (inputs(231));
    layer0_outputs(609) <= not(inputs(212));
    layer0_outputs(610) <= not(inputs(179));
    layer0_outputs(611) <= (inputs(241)) or (inputs(247));
    layer0_outputs(612) <= not((inputs(140)) or (inputs(123)));
    layer0_outputs(613) <= (inputs(72)) and not (inputs(32));
    layer0_outputs(614) <= (inputs(198)) and not (inputs(82));
    layer0_outputs(615) <= (inputs(254)) or (inputs(147));
    layer0_outputs(616) <= not(inputs(220));
    layer0_outputs(617) <= not((inputs(177)) or (inputs(141)));
    layer0_outputs(618) <= not(inputs(46));
    layer0_outputs(619) <= inputs(232);
    layer0_outputs(620) <= not(inputs(21)) or (inputs(118));
    layer0_outputs(621) <= inputs(95);
    layer0_outputs(622) <= (inputs(221)) and not (inputs(59));
    layer0_outputs(623) <= not(inputs(18));
    layer0_outputs(624) <= not(inputs(133)) or (inputs(64));
    layer0_outputs(625) <= inputs(79);
    layer0_outputs(626) <= (inputs(155)) and not (inputs(101));
    layer0_outputs(627) <= not(inputs(22)) or (inputs(97));
    layer0_outputs(628) <= not(inputs(90));
    layer0_outputs(629) <= inputs(163);
    layer0_outputs(630) <= not(inputs(90)) or (inputs(255));
    layer0_outputs(631) <= not((inputs(176)) or (inputs(68)));
    layer0_outputs(632) <= not(inputs(164)) or (inputs(95));
    layer0_outputs(633) <= not((inputs(83)) xor (inputs(22)));
    layer0_outputs(634) <= (inputs(181)) and not (inputs(15));
    layer0_outputs(635) <= not((inputs(128)) or (inputs(239)));
    layer0_outputs(636) <= not((inputs(96)) or (inputs(121)));
    layer0_outputs(637) <= not((inputs(242)) or (inputs(200)));
    layer0_outputs(638) <= inputs(216);
    layer0_outputs(639) <= not(inputs(137));
    layer0_outputs(640) <= not(inputs(152)) or (inputs(160));
    layer0_outputs(641) <= (inputs(71)) and not (inputs(255));
    layer0_outputs(642) <= not(inputs(225));
    layer0_outputs(643) <= inputs(208);
    layer0_outputs(644) <= not(inputs(39)) or (inputs(149));
    layer0_outputs(645) <= not((inputs(233)) xor (inputs(188)));
    layer0_outputs(646) <= not((inputs(193)) or (inputs(131)));
    layer0_outputs(647) <= not((inputs(168)) and (inputs(121)));
    layer0_outputs(648) <= not(inputs(72)) or (inputs(248));
    layer0_outputs(649) <= not((inputs(212)) or (inputs(214)));
    layer0_outputs(650) <= (inputs(112)) and not (inputs(140));
    layer0_outputs(651) <= not(inputs(188));
    layer0_outputs(652) <= not((inputs(177)) or (inputs(31)));
    layer0_outputs(653) <= (inputs(206)) or (inputs(54));
    layer0_outputs(654) <= (inputs(108)) or (inputs(139));
    layer0_outputs(655) <= not((inputs(112)) or (inputs(209)));
    layer0_outputs(656) <= not(inputs(138)) or (inputs(34));
    layer0_outputs(657) <= not(inputs(157));
    layer0_outputs(658) <= inputs(152);
    layer0_outputs(659) <= not(inputs(98));
    layer0_outputs(660) <= (inputs(170)) and not (inputs(231));
    layer0_outputs(661) <= (inputs(89)) and not (inputs(86));
    layer0_outputs(662) <= (inputs(19)) and not (inputs(235));
    layer0_outputs(663) <= not(inputs(142));
    layer0_outputs(664) <= (inputs(250)) or (inputs(63));
    layer0_outputs(665) <= not(inputs(213));
    layer0_outputs(666) <= (inputs(68)) and not (inputs(63));
    layer0_outputs(667) <= (inputs(222)) or (inputs(175));
    layer0_outputs(668) <= (inputs(251)) or (inputs(146));
    layer0_outputs(669) <= not(inputs(203)) or (inputs(18));
    layer0_outputs(670) <= not(inputs(229)) or (inputs(2));
    layer0_outputs(671) <= inputs(146);
    layer0_outputs(672) <= (inputs(86)) and not (inputs(127));
    layer0_outputs(673) <= not(inputs(151));
    layer0_outputs(674) <= (inputs(97)) and not (inputs(249));
    layer0_outputs(675) <= not(inputs(105));
    layer0_outputs(676) <= (inputs(226)) or (inputs(39));
    layer0_outputs(677) <= (inputs(142)) and not (inputs(94));
    layer0_outputs(678) <= (inputs(218)) and not (inputs(124));
    layer0_outputs(679) <= (inputs(89)) and not (inputs(54));
    layer0_outputs(680) <= not(inputs(203));
    layer0_outputs(681) <= inputs(236);
    layer0_outputs(682) <= '0';
    layer0_outputs(683) <= not((inputs(125)) or (inputs(110)));
    layer0_outputs(684) <= inputs(206);
    layer0_outputs(685) <= not(inputs(231));
    layer0_outputs(686) <= (inputs(49)) and not (inputs(86));
    layer0_outputs(687) <= (inputs(217)) and not (inputs(4));
    layer0_outputs(688) <= not((inputs(229)) or (inputs(7)));
    layer0_outputs(689) <= '1';
    layer0_outputs(690) <= (inputs(145)) or (inputs(206));
    layer0_outputs(691) <= (inputs(148)) xor (inputs(80));
    layer0_outputs(692) <= inputs(179);
    layer0_outputs(693) <= not(inputs(169)) or (inputs(111));
    layer0_outputs(694) <= (inputs(237)) or (inputs(20));
    layer0_outputs(695) <= not((inputs(170)) or (inputs(64)));
    layer0_outputs(696) <= not(inputs(192));
    layer0_outputs(697) <= (inputs(189)) or (inputs(95));
    layer0_outputs(698) <= (inputs(6)) or (inputs(12));
    layer0_outputs(699) <= (inputs(146)) and not (inputs(150));
    layer0_outputs(700) <= not(inputs(178)) or (inputs(176));
    layer0_outputs(701) <= inputs(181);
    layer0_outputs(702) <= (inputs(86)) and not (inputs(46));
    layer0_outputs(703) <= not(inputs(242)) or (inputs(236));
    layer0_outputs(704) <= (inputs(97)) and not (inputs(7));
    layer0_outputs(705) <= (inputs(248)) and not (inputs(186));
    layer0_outputs(706) <= inputs(219);
    layer0_outputs(707) <= not((inputs(110)) or (inputs(162)));
    layer0_outputs(708) <= not(inputs(22));
    layer0_outputs(709) <= not(inputs(247));
    layer0_outputs(710) <= not(inputs(108));
    layer0_outputs(711) <= (inputs(185)) and (inputs(95));
    layer0_outputs(712) <= not(inputs(73)) or (inputs(21));
    layer0_outputs(713) <= not(inputs(106));
    layer0_outputs(714) <= '1';
    layer0_outputs(715) <= (inputs(39)) and not (inputs(118));
    layer0_outputs(716) <= not(inputs(85)) or (inputs(48));
    layer0_outputs(717) <= not(inputs(188)) or (inputs(51));
    layer0_outputs(718) <= not(inputs(100));
    layer0_outputs(719) <= not((inputs(205)) or (inputs(161)));
    layer0_outputs(720) <= not((inputs(233)) and (inputs(57)));
    layer0_outputs(721) <= inputs(132);
    layer0_outputs(722) <= not(inputs(52)) or (inputs(137));
    layer0_outputs(723) <= (inputs(126)) or (inputs(239));
    layer0_outputs(724) <= not((inputs(223)) xor (inputs(204)));
    layer0_outputs(725) <= inputs(169);
    layer0_outputs(726) <= inputs(148);
    layer0_outputs(727) <= (inputs(176)) or (inputs(107));
    layer0_outputs(728) <= not(inputs(252)) or (inputs(234));
    layer0_outputs(729) <= not(inputs(182)) or (inputs(58));
    layer0_outputs(730) <= not(inputs(83));
    layer0_outputs(731) <= inputs(63);
    layer0_outputs(732) <= not(inputs(171));
    layer0_outputs(733) <= inputs(182);
    layer0_outputs(734) <= not((inputs(6)) or (inputs(81)));
    layer0_outputs(735) <= not(inputs(230));
    layer0_outputs(736) <= (inputs(168)) or (inputs(59));
    layer0_outputs(737) <= not(inputs(34));
    layer0_outputs(738) <= inputs(29);
    layer0_outputs(739) <= not((inputs(32)) or (inputs(59)));
    layer0_outputs(740) <= inputs(115);
    layer0_outputs(741) <= (inputs(42)) and not (inputs(116));
    layer0_outputs(742) <= not((inputs(107)) or (inputs(4)));
    layer0_outputs(743) <= not(inputs(163));
    layer0_outputs(744) <= not(inputs(228));
    layer0_outputs(745) <= not(inputs(21));
    layer0_outputs(746) <= not((inputs(29)) or (inputs(161)));
    layer0_outputs(747) <= not(inputs(88));
    layer0_outputs(748) <= not(inputs(179));
    layer0_outputs(749) <= not((inputs(179)) or (inputs(100)));
    layer0_outputs(750) <= not((inputs(134)) or (inputs(143)));
    layer0_outputs(751) <= (inputs(36)) and not (inputs(191));
    layer0_outputs(752) <= (inputs(122)) and not (inputs(31));
    layer0_outputs(753) <= not(inputs(27)) or (inputs(185));
    layer0_outputs(754) <= inputs(99);
    layer0_outputs(755) <= (inputs(38)) and not (inputs(19));
    layer0_outputs(756) <= inputs(141);
    layer0_outputs(757) <= not(inputs(104));
    layer0_outputs(758) <= not(inputs(187));
    layer0_outputs(759) <= not(inputs(132)) or (inputs(167));
    layer0_outputs(760) <= not(inputs(2));
    layer0_outputs(761) <= not((inputs(24)) and (inputs(25)));
    layer0_outputs(762) <= (inputs(1)) or (inputs(21));
    layer0_outputs(763) <= not(inputs(38)) or (inputs(158));
    layer0_outputs(764) <= not(inputs(170)) or (inputs(141));
    layer0_outputs(765) <= (inputs(96)) or (inputs(181));
    layer0_outputs(766) <= not((inputs(61)) and (inputs(92)));
    layer0_outputs(767) <= not(inputs(144)) or (inputs(48));
    layer0_outputs(768) <= inputs(235);
    layer0_outputs(769) <= inputs(123);
    layer0_outputs(770) <= (inputs(16)) or (inputs(200));
    layer0_outputs(771) <= (inputs(240)) or (inputs(145));
    layer0_outputs(772) <= (inputs(88)) and not (inputs(0));
    layer0_outputs(773) <= (inputs(86)) and not (inputs(50));
    layer0_outputs(774) <= (inputs(173)) xor (inputs(238));
    layer0_outputs(775) <= (inputs(102)) or (inputs(71));
    layer0_outputs(776) <= inputs(91);
    layer0_outputs(777) <= (inputs(210)) and not (inputs(14));
    layer0_outputs(778) <= (inputs(82)) or (inputs(116));
    layer0_outputs(779) <= not(inputs(69));
    layer0_outputs(780) <= not((inputs(35)) or (inputs(228)));
    layer0_outputs(781) <= (inputs(87)) and not (inputs(254));
    layer0_outputs(782) <= not(inputs(93));
    layer0_outputs(783) <= '1';
    layer0_outputs(784) <= (inputs(247)) and not (inputs(74));
    layer0_outputs(785) <= not(inputs(180));
    layer0_outputs(786) <= '1';
    layer0_outputs(787) <= (inputs(52)) and not (inputs(199));
    layer0_outputs(788) <= not(inputs(146));
    layer0_outputs(789) <= not((inputs(94)) or (inputs(21)));
    layer0_outputs(790) <= (inputs(220)) or (inputs(28));
    layer0_outputs(791) <= inputs(85);
    layer0_outputs(792) <= (inputs(151)) and (inputs(136));
    layer0_outputs(793) <= inputs(172);
    layer0_outputs(794) <= not(inputs(136));
    layer0_outputs(795) <= not(inputs(133)) or (inputs(158));
    layer0_outputs(796) <= not((inputs(160)) xor (inputs(123)));
    layer0_outputs(797) <= inputs(234);
    layer0_outputs(798) <= (inputs(102)) or (inputs(85));
    layer0_outputs(799) <= not((inputs(24)) or (inputs(46)));
    layer0_outputs(800) <= (inputs(38)) and not (inputs(114));
    layer0_outputs(801) <= (inputs(121)) and not (inputs(241));
    layer0_outputs(802) <= (inputs(142)) or (inputs(211));
    layer0_outputs(803) <= not(inputs(252));
    layer0_outputs(804) <= (inputs(148)) or (inputs(239));
    layer0_outputs(805) <= inputs(60);
    layer0_outputs(806) <= not(inputs(195));
    layer0_outputs(807) <= not((inputs(40)) or (inputs(22)));
    layer0_outputs(808) <= inputs(244);
    layer0_outputs(809) <= (inputs(253)) and not (inputs(80));
    layer0_outputs(810) <= (inputs(221)) and not (inputs(186));
    layer0_outputs(811) <= not(inputs(223)) or (inputs(221));
    layer0_outputs(812) <= not((inputs(161)) or (inputs(139)));
    layer0_outputs(813) <= (inputs(38)) and not (inputs(192));
    layer0_outputs(814) <= not(inputs(99));
    layer0_outputs(815) <= inputs(168);
    layer0_outputs(816) <= (inputs(197)) and not (inputs(167));
    layer0_outputs(817) <= not(inputs(163));
    layer0_outputs(818) <= (inputs(211)) or (inputs(114));
    layer0_outputs(819) <= inputs(24);
    layer0_outputs(820) <= not(inputs(209));
    layer0_outputs(821) <= not((inputs(214)) xor (inputs(83)));
    layer0_outputs(822) <= (inputs(68)) and not (inputs(217));
    layer0_outputs(823) <= inputs(104);
    layer0_outputs(824) <= not((inputs(50)) or (inputs(91)));
    layer0_outputs(825) <= not((inputs(7)) or (inputs(28)));
    layer0_outputs(826) <= (inputs(123)) and not (inputs(224));
    layer0_outputs(827) <= not(inputs(238));
    layer0_outputs(828) <= (inputs(136)) and not (inputs(157));
    layer0_outputs(829) <= (inputs(247)) and not (inputs(29));
    layer0_outputs(830) <= (inputs(232)) and not (inputs(164));
    layer0_outputs(831) <= (inputs(76)) xor (inputs(95));
    layer0_outputs(832) <= not((inputs(129)) xor (inputs(6)));
    layer0_outputs(833) <= (inputs(237)) and not (inputs(5));
    layer0_outputs(834) <= (inputs(240)) or (inputs(220));
    layer0_outputs(835) <= (inputs(240)) or (inputs(185));
    layer0_outputs(836) <= inputs(9);
    layer0_outputs(837) <= inputs(185);
    layer0_outputs(838) <= not(inputs(26)) or (inputs(162));
    layer0_outputs(839) <= not(inputs(74)) or (inputs(2));
    layer0_outputs(840) <= not(inputs(167));
    layer0_outputs(841) <= not(inputs(145));
    layer0_outputs(842) <= inputs(118);
    layer0_outputs(843) <= '1';
    layer0_outputs(844) <= not(inputs(210));
    layer0_outputs(845) <= '1';
    layer0_outputs(846) <= not(inputs(68)) or (inputs(51));
    layer0_outputs(847) <= not((inputs(238)) or (inputs(119)));
    layer0_outputs(848) <= (inputs(47)) and not (inputs(241));
    layer0_outputs(849) <= '0';
    layer0_outputs(850) <= inputs(182);
    layer0_outputs(851) <= (inputs(78)) and not (inputs(128));
    layer0_outputs(852) <= not((inputs(219)) or (inputs(177)));
    layer0_outputs(853) <= (inputs(195)) and not (inputs(237));
    layer0_outputs(854) <= not(inputs(120));
    layer0_outputs(855) <= not((inputs(235)) or (inputs(251)));
    layer0_outputs(856) <= (inputs(120)) and not (inputs(199));
    layer0_outputs(857) <= (inputs(161)) or (inputs(157));
    layer0_outputs(858) <= inputs(167);
    layer0_outputs(859) <= (inputs(135)) or (inputs(253));
    layer0_outputs(860) <= not(inputs(163));
    layer0_outputs(861) <= not(inputs(166));
    layer0_outputs(862) <= not(inputs(143));
    layer0_outputs(863) <= not(inputs(174));
    layer0_outputs(864) <= not(inputs(184));
    layer0_outputs(865) <= inputs(198);
    layer0_outputs(866) <= not(inputs(3));
    layer0_outputs(867) <= inputs(119);
    layer0_outputs(868) <= (inputs(246)) or (inputs(240));
    layer0_outputs(869) <= (inputs(121)) or (inputs(135));
    layer0_outputs(870) <= (inputs(178)) or (inputs(194));
    layer0_outputs(871) <= not(inputs(109));
    layer0_outputs(872) <= (inputs(103)) and not (inputs(123));
    layer0_outputs(873) <= inputs(1);
    layer0_outputs(874) <= not(inputs(204)) or (inputs(29));
    layer0_outputs(875) <= not(inputs(190));
    layer0_outputs(876) <= inputs(126);
    layer0_outputs(877) <= (inputs(175)) or (inputs(56));
    layer0_outputs(878) <= not((inputs(112)) or (inputs(237)));
    layer0_outputs(879) <= inputs(67);
    layer0_outputs(880) <= inputs(132);
    layer0_outputs(881) <= inputs(67);
    layer0_outputs(882) <= not((inputs(162)) or (inputs(181)));
    layer0_outputs(883) <= not(inputs(167));
    layer0_outputs(884) <= not(inputs(245));
    layer0_outputs(885) <= not(inputs(121));
    layer0_outputs(886) <= inputs(13);
    layer0_outputs(887) <= inputs(154);
    layer0_outputs(888) <= not(inputs(206));
    layer0_outputs(889) <= not((inputs(126)) xor (inputs(136)));
    layer0_outputs(890) <= inputs(218);
    layer0_outputs(891) <= not(inputs(60)) or (inputs(249));
    layer0_outputs(892) <= not(inputs(9)) or (inputs(194));
    layer0_outputs(893) <= (inputs(238)) or (inputs(109));
    layer0_outputs(894) <= not(inputs(223));
    layer0_outputs(895) <= not(inputs(68));
    layer0_outputs(896) <= not((inputs(240)) or (inputs(55)));
    layer0_outputs(897) <= not((inputs(197)) or (inputs(113)));
    layer0_outputs(898) <= not(inputs(177));
    layer0_outputs(899) <= inputs(237);
    layer0_outputs(900) <= not(inputs(26)) or (inputs(115));
    layer0_outputs(901) <= not((inputs(72)) and (inputs(44)));
    layer0_outputs(902) <= inputs(23);
    layer0_outputs(903) <= not(inputs(54)) or (inputs(207));
    layer0_outputs(904) <= inputs(75);
    layer0_outputs(905) <= (inputs(87)) xor (inputs(114));
    layer0_outputs(906) <= not(inputs(134));
    layer0_outputs(907) <= (inputs(211)) and not (inputs(48));
    layer0_outputs(908) <= inputs(106);
    layer0_outputs(909) <= (inputs(221)) or (inputs(27));
    layer0_outputs(910) <= (inputs(181)) xor (inputs(185));
    layer0_outputs(911) <= not(inputs(225));
    layer0_outputs(912) <= inputs(168);
    layer0_outputs(913) <= inputs(153);
    layer0_outputs(914) <= not(inputs(10));
    layer0_outputs(915) <= not(inputs(82));
    layer0_outputs(916) <= inputs(131);
    layer0_outputs(917) <= (inputs(163)) and (inputs(74));
    layer0_outputs(918) <= not(inputs(28));
    layer0_outputs(919) <= '0';
    layer0_outputs(920) <= not((inputs(49)) or (inputs(47)));
    layer0_outputs(921) <= not((inputs(96)) or (inputs(70)));
    layer0_outputs(922) <= not((inputs(89)) or (inputs(88)));
    layer0_outputs(923) <= inputs(98);
    layer0_outputs(924) <= not((inputs(76)) or (inputs(236)));
    layer0_outputs(925) <= (inputs(70)) or (inputs(232));
    layer0_outputs(926) <= inputs(226);
    layer0_outputs(927) <= (inputs(229)) and (inputs(109));
    layer0_outputs(928) <= inputs(20);
    layer0_outputs(929) <= not(inputs(184)) or (inputs(80));
    layer0_outputs(930) <= (inputs(69)) and not (inputs(106));
    layer0_outputs(931) <= not(inputs(92)) or (inputs(46));
    layer0_outputs(932) <= not(inputs(93));
    layer0_outputs(933) <= not(inputs(151));
    layer0_outputs(934) <= not((inputs(113)) xor (inputs(68)));
    layer0_outputs(935) <= (inputs(106)) xor (inputs(204));
    layer0_outputs(936) <= not(inputs(243));
    layer0_outputs(937) <= (inputs(233)) and not (inputs(165));
    layer0_outputs(938) <= inputs(72);
    layer0_outputs(939) <= (inputs(200)) or (inputs(32));
    layer0_outputs(940) <= not((inputs(113)) or (inputs(67)));
    layer0_outputs(941) <= not((inputs(75)) or (inputs(73)));
    layer0_outputs(942) <= not(inputs(145));
    layer0_outputs(943) <= (inputs(178)) or (inputs(110));
    layer0_outputs(944) <= (inputs(165)) or (inputs(192));
    layer0_outputs(945) <= inputs(145);
    layer0_outputs(946) <= inputs(104);
    layer0_outputs(947) <= inputs(132);
    layer0_outputs(948) <= (inputs(10)) or (inputs(24));
    layer0_outputs(949) <= (inputs(117)) and not (inputs(3));
    layer0_outputs(950) <= not(inputs(195)) or (inputs(10));
    layer0_outputs(951) <= not((inputs(130)) or (inputs(243)));
    layer0_outputs(952) <= not((inputs(3)) xor (inputs(48)));
    layer0_outputs(953) <= (inputs(230)) and not (inputs(110));
    layer0_outputs(954) <= (inputs(187)) or (inputs(253));
    layer0_outputs(955) <= not((inputs(144)) or (inputs(205)));
    layer0_outputs(956) <= not((inputs(71)) or (inputs(243)));
    layer0_outputs(957) <= not(inputs(122));
    layer0_outputs(958) <= inputs(232);
    layer0_outputs(959) <= not(inputs(98));
    layer0_outputs(960) <= not((inputs(173)) or (inputs(179)));
    layer0_outputs(961) <= (inputs(113)) and not (inputs(7));
    layer0_outputs(962) <= not((inputs(138)) or (inputs(115)));
    layer0_outputs(963) <= not(inputs(163));
    layer0_outputs(964) <= inputs(196);
    layer0_outputs(965) <= (inputs(55)) and not (inputs(226));
    layer0_outputs(966) <= inputs(9);
    layer0_outputs(967) <= '1';
    layer0_outputs(968) <= (inputs(185)) and (inputs(146));
    layer0_outputs(969) <= inputs(109);
    layer0_outputs(970) <= not(inputs(203));
    layer0_outputs(971) <= inputs(56);
    layer0_outputs(972) <= not(inputs(3)) or (inputs(239));
    layer0_outputs(973) <= not((inputs(47)) or (inputs(11)));
    layer0_outputs(974) <= (inputs(180)) and not (inputs(240));
    layer0_outputs(975) <= (inputs(122)) or (inputs(36));
    layer0_outputs(976) <= (inputs(2)) or (inputs(150));
    layer0_outputs(977) <= inputs(59);
    layer0_outputs(978) <= (inputs(25)) and not (inputs(142));
    layer0_outputs(979) <= not(inputs(247)) or (inputs(5));
    layer0_outputs(980) <= not(inputs(167));
    layer0_outputs(981) <= not(inputs(134));
    layer0_outputs(982) <= inputs(153);
    layer0_outputs(983) <= inputs(160);
    layer0_outputs(984) <= not(inputs(42)) or (inputs(239));
    layer0_outputs(985) <= (inputs(205)) or (inputs(102));
    layer0_outputs(986) <= inputs(169);
    layer0_outputs(987) <= (inputs(186)) and not (inputs(133));
    layer0_outputs(988) <= (inputs(165)) and (inputs(232));
    layer0_outputs(989) <= (inputs(107)) and not (inputs(207));
    layer0_outputs(990) <= not((inputs(143)) or (inputs(121)));
    layer0_outputs(991) <= (inputs(73)) or (inputs(0));
    layer0_outputs(992) <= (inputs(212)) and not (inputs(22));
    layer0_outputs(993) <= not((inputs(146)) xor (inputs(120)));
    layer0_outputs(994) <= not(inputs(181));
    layer0_outputs(995) <= not((inputs(177)) or (inputs(64)));
    layer0_outputs(996) <= '1';
    layer0_outputs(997) <= not((inputs(57)) xor (inputs(22)));
    layer0_outputs(998) <= (inputs(108)) and (inputs(35));
    layer0_outputs(999) <= not((inputs(79)) or (inputs(52)));
    layer0_outputs(1000) <= (inputs(71)) and not (inputs(220));
    layer0_outputs(1001) <= (inputs(50)) and not (inputs(83));
    layer0_outputs(1002) <= (inputs(208)) or (inputs(114));
    layer0_outputs(1003) <= not(inputs(245));
    layer0_outputs(1004) <= (inputs(175)) xor (inputs(234));
    layer0_outputs(1005) <= inputs(197);
    layer0_outputs(1006) <= not(inputs(8)) or (inputs(241));
    layer0_outputs(1007) <= inputs(107);
    layer0_outputs(1008) <= inputs(100);
    layer0_outputs(1009) <= (inputs(22)) and not (inputs(131));
    layer0_outputs(1010) <= not(inputs(118));
    layer0_outputs(1011) <= inputs(253);
    layer0_outputs(1012) <= inputs(126);
    layer0_outputs(1013) <= not((inputs(107)) or (inputs(1)));
    layer0_outputs(1014) <= (inputs(28)) xor (inputs(94));
    layer0_outputs(1015) <= (inputs(23)) or (inputs(208));
    layer0_outputs(1016) <= '1';
    layer0_outputs(1017) <= not((inputs(80)) or (inputs(195)));
    layer0_outputs(1018) <= '0';
    layer0_outputs(1019) <= (inputs(234)) and not (inputs(40));
    layer0_outputs(1020) <= not(inputs(103));
    layer0_outputs(1021) <= inputs(212);
    layer0_outputs(1022) <= (inputs(236)) and not (inputs(112));
    layer0_outputs(1023) <= inputs(229);
    layer0_outputs(1024) <= not((inputs(255)) xor (inputs(188)));
    layer0_outputs(1025) <= inputs(104);
    layer0_outputs(1026) <= (inputs(178)) or (inputs(189));
    layer0_outputs(1027) <= not((inputs(217)) or (inputs(50)));
    layer0_outputs(1028) <= not(inputs(232));
    layer0_outputs(1029) <= (inputs(236)) or (inputs(77));
    layer0_outputs(1030) <= (inputs(70)) or (inputs(25));
    layer0_outputs(1031) <= (inputs(228)) and not (inputs(58));
    layer0_outputs(1032) <= not(inputs(86)) or (inputs(3));
    layer0_outputs(1033) <= inputs(127);
    layer0_outputs(1034) <= (inputs(40)) or (inputs(243));
    layer0_outputs(1035) <= not(inputs(215)) or (inputs(236));
    layer0_outputs(1036) <= (inputs(229)) and not (inputs(165));
    layer0_outputs(1037) <= not(inputs(150));
    layer0_outputs(1038) <= not(inputs(66)) or (inputs(143));
    layer0_outputs(1039) <= inputs(211);
    layer0_outputs(1040) <= not(inputs(63));
    layer0_outputs(1041) <= (inputs(191)) or (inputs(249));
    layer0_outputs(1042) <= inputs(75);
    layer0_outputs(1043) <= (inputs(249)) or (inputs(66));
    layer0_outputs(1044) <= not((inputs(113)) or (inputs(219)));
    layer0_outputs(1045) <= (inputs(37)) and not (inputs(244));
    layer0_outputs(1046) <= not(inputs(117));
    layer0_outputs(1047) <= not(inputs(131));
    layer0_outputs(1048) <= not(inputs(136)) or (inputs(236));
    layer0_outputs(1049) <= '0';
    layer0_outputs(1050) <= (inputs(2)) and not (inputs(67));
    layer0_outputs(1051) <= not(inputs(112)) or (inputs(14));
    layer0_outputs(1052) <= not(inputs(233));
    layer0_outputs(1053) <= (inputs(216)) and not (inputs(32));
    layer0_outputs(1054) <= inputs(42);
    layer0_outputs(1055) <= inputs(212);
    layer0_outputs(1056) <= (inputs(207)) and not (inputs(208));
    layer0_outputs(1057) <= (inputs(226)) or (inputs(248));
    layer0_outputs(1058) <= not(inputs(96));
    layer0_outputs(1059) <= not(inputs(42));
    layer0_outputs(1060) <= (inputs(240)) or (inputs(71));
    layer0_outputs(1061) <= (inputs(198)) and not (inputs(106));
    layer0_outputs(1062) <= (inputs(194)) and not (inputs(249));
    layer0_outputs(1063) <= (inputs(93)) or (inputs(19));
    layer0_outputs(1064) <= not(inputs(228));
    layer0_outputs(1065) <= (inputs(49)) and (inputs(144));
    layer0_outputs(1066) <= not((inputs(169)) or (inputs(81)));
    layer0_outputs(1067) <= (inputs(171)) or (inputs(220));
    layer0_outputs(1068) <= (inputs(119)) or (inputs(36));
    layer0_outputs(1069) <= '0';
    layer0_outputs(1070) <= not(inputs(111)) or (inputs(3));
    layer0_outputs(1071) <= (inputs(118)) and not (inputs(0));
    layer0_outputs(1072) <= inputs(168);
    layer0_outputs(1073) <= not(inputs(81));
    layer0_outputs(1074) <= (inputs(32)) or (inputs(171));
    layer0_outputs(1075) <= inputs(151);
    layer0_outputs(1076) <= (inputs(193)) or (inputs(158));
    layer0_outputs(1077) <= not((inputs(31)) xor (inputs(197)));
    layer0_outputs(1078) <= inputs(99);
    layer0_outputs(1079) <= inputs(85);
    layer0_outputs(1080) <= inputs(178);
    layer0_outputs(1081) <= not((inputs(132)) and (inputs(72)));
    layer0_outputs(1082) <= not(inputs(83));
    layer0_outputs(1083) <= not(inputs(11));
    layer0_outputs(1084) <= inputs(38);
    layer0_outputs(1085) <= (inputs(106)) and not (inputs(143));
    layer0_outputs(1086) <= inputs(13);
    layer0_outputs(1087) <= not((inputs(220)) or (inputs(164)));
    layer0_outputs(1088) <= inputs(124);
    layer0_outputs(1089) <= inputs(217);
    layer0_outputs(1090) <= inputs(211);
    layer0_outputs(1091) <= inputs(113);
    layer0_outputs(1092) <= inputs(23);
    layer0_outputs(1093) <= not(inputs(112)) or (inputs(17));
    layer0_outputs(1094) <= not(inputs(74)) or (inputs(4));
    layer0_outputs(1095) <= not(inputs(20));
    layer0_outputs(1096) <= not(inputs(151)) or (inputs(237));
    layer0_outputs(1097) <= not(inputs(60));
    layer0_outputs(1098) <= not(inputs(119));
    layer0_outputs(1099) <= not(inputs(149)) or (inputs(77));
    layer0_outputs(1100) <= (inputs(152)) and not (inputs(132));
    layer0_outputs(1101) <= not((inputs(72)) or (inputs(9)));
    layer0_outputs(1102) <= not(inputs(145));
    layer0_outputs(1103) <= not(inputs(189));
    layer0_outputs(1104) <= not(inputs(109));
    layer0_outputs(1105) <= inputs(63);
    layer0_outputs(1106) <= not(inputs(108));
    layer0_outputs(1107) <= inputs(191);
    layer0_outputs(1108) <= (inputs(153)) and (inputs(217));
    layer0_outputs(1109) <= inputs(249);
    layer0_outputs(1110) <= not(inputs(43));
    layer0_outputs(1111) <= (inputs(55)) and not (inputs(158));
    layer0_outputs(1112) <= not((inputs(170)) xor (inputs(139)));
    layer0_outputs(1113) <= not(inputs(37));
    layer0_outputs(1114) <= not(inputs(58)) or (inputs(79));
    layer0_outputs(1115) <= not(inputs(147)) or (inputs(58));
    layer0_outputs(1116) <= not(inputs(129));
    layer0_outputs(1117) <= not(inputs(247)) or (inputs(254));
    layer0_outputs(1118) <= (inputs(104)) and not (inputs(210));
    layer0_outputs(1119) <= (inputs(159)) or (inputs(121));
    layer0_outputs(1120) <= not((inputs(147)) or (inputs(173)));
    layer0_outputs(1121) <= not(inputs(120));
    layer0_outputs(1122) <= not(inputs(147));
    layer0_outputs(1123) <= not((inputs(225)) or (inputs(173)));
    layer0_outputs(1124) <= '0';
    layer0_outputs(1125) <= not((inputs(4)) or (inputs(205)));
    layer0_outputs(1126) <= not((inputs(218)) or (inputs(248)));
    layer0_outputs(1127) <= not(inputs(162));
    layer0_outputs(1128) <= (inputs(160)) and not (inputs(56));
    layer0_outputs(1129) <= not(inputs(229));
    layer0_outputs(1130) <= inputs(180);
    layer0_outputs(1131) <= (inputs(43)) and not (inputs(105));
    layer0_outputs(1132) <= not((inputs(240)) or (inputs(182)));
    layer0_outputs(1133) <= inputs(167);
    layer0_outputs(1134) <= not(inputs(179));
    layer0_outputs(1135) <= inputs(200);
    layer0_outputs(1136) <= (inputs(71)) or (inputs(180));
    layer0_outputs(1137) <= not(inputs(152));
    layer0_outputs(1138) <= inputs(218);
    layer0_outputs(1139) <= not(inputs(87));
    layer0_outputs(1140) <= not((inputs(110)) or (inputs(74)));
    layer0_outputs(1141) <= not((inputs(154)) xor (inputs(102)));
    layer0_outputs(1142) <= (inputs(70)) and not (inputs(1));
    layer0_outputs(1143) <= inputs(14);
    layer0_outputs(1144) <= not((inputs(80)) xor (inputs(222)));
    layer0_outputs(1145) <= inputs(10);
    layer0_outputs(1146) <= not(inputs(36));
    layer0_outputs(1147) <= '1';
    layer0_outputs(1148) <= not((inputs(4)) or (inputs(189)));
    layer0_outputs(1149) <= inputs(197);
    layer0_outputs(1150) <= not(inputs(75));
    layer0_outputs(1151) <= not(inputs(217));
    layer0_outputs(1152) <= inputs(12);
    layer0_outputs(1153) <= (inputs(209)) and not (inputs(15));
    layer0_outputs(1154) <= (inputs(88)) and not (inputs(205));
    layer0_outputs(1155) <= inputs(86);
    layer0_outputs(1156) <= (inputs(252)) or (inputs(150));
    layer0_outputs(1157) <= not(inputs(88)) or (inputs(148));
    layer0_outputs(1158) <= inputs(26);
    layer0_outputs(1159) <= (inputs(214)) and (inputs(202));
    layer0_outputs(1160) <= not(inputs(222));
    layer0_outputs(1161) <= not(inputs(101));
    layer0_outputs(1162) <= (inputs(109)) or (inputs(44));
    layer0_outputs(1163) <= not(inputs(100));
    layer0_outputs(1164) <= not(inputs(136));
    layer0_outputs(1165) <= inputs(207);
    layer0_outputs(1166) <= '1';
    layer0_outputs(1167) <= (inputs(255)) or (inputs(150));
    layer0_outputs(1168) <= not(inputs(29)) or (inputs(207));
    layer0_outputs(1169) <= (inputs(136)) and not (inputs(195));
    layer0_outputs(1170) <= inputs(42);
    layer0_outputs(1171) <= not(inputs(96));
    layer0_outputs(1172) <= not(inputs(247)) or (inputs(31));
    layer0_outputs(1173) <= not(inputs(88)) or (inputs(39));
    layer0_outputs(1174) <= inputs(165);
    layer0_outputs(1175) <= inputs(19);
    layer0_outputs(1176) <= not(inputs(36));
    layer0_outputs(1177) <= not(inputs(78)) or (inputs(115));
    layer0_outputs(1178) <= not(inputs(72)) or (inputs(238));
    layer0_outputs(1179) <= inputs(41);
    layer0_outputs(1180) <= (inputs(126)) xor (inputs(104));
    layer0_outputs(1181) <= not(inputs(211));
    layer0_outputs(1182) <= not((inputs(194)) or (inputs(115)));
    layer0_outputs(1183) <= (inputs(179)) or (inputs(158));
    layer0_outputs(1184) <= not((inputs(178)) or (inputs(92)));
    layer0_outputs(1185) <= (inputs(7)) and not (inputs(87));
    layer0_outputs(1186) <= not(inputs(212));
    layer0_outputs(1187) <= not((inputs(122)) and (inputs(116)));
    layer0_outputs(1188) <= inputs(40);
    layer0_outputs(1189) <= not((inputs(147)) xor (inputs(116)));
    layer0_outputs(1190) <= not(inputs(106));
    layer0_outputs(1191) <= not(inputs(110)) or (inputs(168));
    layer0_outputs(1192) <= not(inputs(124)) or (inputs(181));
    layer0_outputs(1193) <= not(inputs(42));
    layer0_outputs(1194) <= (inputs(134)) and not (inputs(128));
    layer0_outputs(1195) <= not((inputs(107)) or (inputs(252)));
    layer0_outputs(1196) <= not(inputs(195));
    layer0_outputs(1197) <= inputs(212);
    layer0_outputs(1198) <= not(inputs(62));
    layer0_outputs(1199) <= not((inputs(164)) or (inputs(16)));
    layer0_outputs(1200) <= (inputs(80)) xor (inputs(110));
    layer0_outputs(1201) <= not((inputs(85)) and (inputs(114)));
    layer0_outputs(1202) <= not((inputs(218)) xor (inputs(62)));
    layer0_outputs(1203) <= not((inputs(224)) or (inputs(230)));
    layer0_outputs(1204) <= not((inputs(198)) or (inputs(195)));
    layer0_outputs(1205) <= not(inputs(151));
    layer0_outputs(1206) <= not(inputs(4));
    layer0_outputs(1207) <= not((inputs(76)) or (inputs(92)));
    layer0_outputs(1208) <= not((inputs(34)) or (inputs(113)));
    layer0_outputs(1209) <= (inputs(247)) and not (inputs(70));
    layer0_outputs(1210) <= not((inputs(58)) or (inputs(170)));
    layer0_outputs(1211) <= not((inputs(206)) or (inputs(185)));
    layer0_outputs(1212) <= (inputs(224)) or (inputs(161));
    layer0_outputs(1213) <= not((inputs(108)) or (inputs(7)));
    layer0_outputs(1214) <= not(inputs(182));
    layer0_outputs(1215) <= not((inputs(116)) or (inputs(255)));
    layer0_outputs(1216) <= not((inputs(80)) and (inputs(54)));
    layer0_outputs(1217) <= (inputs(24)) and (inputs(29));
    layer0_outputs(1218) <= not((inputs(254)) or (inputs(253)));
    layer0_outputs(1219) <= not((inputs(238)) or (inputs(91)));
    layer0_outputs(1220) <= inputs(88);
    layer0_outputs(1221) <= not(inputs(81));
    layer0_outputs(1222) <= not((inputs(20)) or (inputs(190)));
    layer0_outputs(1223) <= not((inputs(186)) and (inputs(214)));
    layer0_outputs(1224) <= not(inputs(21));
    layer0_outputs(1225) <= (inputs(213)) and not (inputs(74));
    layer0_outputs(1226) <= not((inputs(218)) or (inputs(202)));
    layer0_outputs(1227) <= not(inputs(164));
    layer0_outputs(1228) <= (inputs(63)) or (inputs(9));
    layer0_outputs(1229) <= (inputs(144)) or (inputs(232));
    layer0_outputs(1230) <= not(inputs(226));
    layer0_outputs(1231) <= not((inputs(105)) or (inputs(30)));
    layer0_outputs(1232) <= '1';
    layer0_outputs(1233) <= '0';
    layer0_outputs(1234) <= inputs(215);
    layer0_outputs(1235) <= inputs(156);
    layer0_outputs(1236) <= inputs(244);
    layer0_outputs(1237) <= (inputs(192)) or (inputs(239));
    layer0_outputs(1238) <= (inputs(68)) and not (inputs(51));
    layer0_outputs(1239) <= inputs(46);
    layer0_outputs(1240) <= not((inputs(76)) xor (inputs(77)));
    layer0_outputs(1241) <= not((inputs(127)) or (inputs(43)));
    layer0_outputs(1242) <= (inputs(81)) and not (inputs(178));
    layer0_outputs(1243) <= not(inputs(230));
    layer0_outputs(1244) <= inputs(176);
    layer0_outputs(1245) <= not((inputs(57)) and (inputs(139)));
    layer0_outputs(1246) <= inputs(107);
    layer0_outputs(1247) <= (inputs(195)) or (inputs(178));
    layer0_outputs(1248) <= (inputs(140)) xor (inputs(174));
    layer0_outputs(1249) <= inputs(128);
    layer0_outputs(1250) <= not(inputs(203)) or (inputs(18));
    layer0_outputs(1251) <= not(inputs(142));
    layer0_outputs(1252) <= inputs(104);
    layer0_outputs(1253) <= (inputs(121)) xor (inputs(93));
    layer0_outputs(1254) <= not(inputs(99));
    layer0_outputs(1255) <= not(inputs(60));
    layer0_outputs(1256) <= not((inputs(242)) or (inputs(104)));
    layer0_outputs(1257) <= not(inputs(126));
    layer0_outputs(1258) <= not((inputs(18)) or (inputs(244)));
    layer0_outputs(1259) <= not(inputs(184));
    layer0_outputs(1260) <= not((inputs(119)) or (inputs(236)));
    layer0_outputs(1261) <= inputs(149);
    layer0_outputs(1262) <= (inputs(213)) or (inputs(94));
    layer0_outputs(1263) <= not((inputs(139)) or (inputs(70)));
    layer0_outputs(1264) <= (inputs(244)) and (inputs(210));
    layer0_outputs(1265) <= inputs(98);
    layer0_outputs(1266) <= (inputs(33)) or (inputs(217));
    layer0_outputs(1267) <= inputs(17);
    layer0_outputs(1268) <= not((inputs(239)) or (inputs(55)));
    layer0_outputs(1269) <= not(inputs(158)) or (inputs(163));
    layer0_outputs(1270) <= not((inputs(2)) or (inputs(239)));
    layer0_outputs(1271) <= not((inputs(69)) and (inputs(137)));
    layer0_outputs(1272) <= not(inputs(145));
    layer0_outputs(1273) <= (inputs(47)) or (inputs(60));
    layer0_outputs(1274) <= (inputs(215)) and not (inputs(15));
    layer0_outputs(1275) <= (inputs(78)) or (inputs(36));
    layer0_outputs(1276) <= (inputs(194)) or (inputs(54));
    layer0_outputs(1277) <= not((inputs(218)) xor (inputs(121)));
    layer0_outputs(1278) <= not(inputs(86)) or (inputs(16));
    layer0_outputs(1279) <= (inputs(119)) and (inputs(40));
    layer0_outputs(1280) <= not((inputs(145)) or (inputs(254)));
    layer0_outputs(1281) <= inputs(76);
    layer0_outputs(1282) <= inputs(60);
    layer0_outputs(1283) <= not((inputs(120)) and (inputs(108)));
    layer0_outputs(1284) <= '1';
    layer0_outputs(1285) <= not(inputs(196)) or (inputs(175));
    layer0_outputs(1286) <= inputs(120);
    layer0_outputs(1287) <= (inputs(229)) and not (inputs(3));
    layer0_outputs(1288) <= not((inputs(219)) or (inputs(235)));
    layer0_outputs(1289) <= not(inputs(133)) or (inputs(95));
    layer0_outputs(1290) <= (inputs(36)) or (inputs(254));
    layer0_outputs(1291) <= not(inputs(133));
    layer0_outputs(1292) <= (inputs(234)) and not (inputs(126));
    layer0_outputs(1293) <= (inputs(217)) and (inputs(231));
    layer0_outputs(1294) <= inputs(37);
    layer0_outputs(1295) <= not(inputs(151));
    layer0_outputs(1296) <= inputs(166);
    layer0_outputs(1297) <= not(inputs(164));
    layer0_outputs(1298) <= inputs(185);
    layer0_outputs(1299) <= (inputs(75)) and not (inputs(79));
    layer0_outputs(1300) <= '1';
    layer0_outputs(1301) <= '0';
    layer0_outputs(1302) <= not((inputs(81)) or (inputs(29)));
    layer0_outputs(1303) <= inputs(218);
    layer0_outputs(1304) <= (inputs(34)) and not (inputs(236));
    layer0_outputs(1305) <= inputs(92);
    layer0_outputs(1306) <= inputs(47);
    layer0_outputs(1307) <= inputs(192);
    layer0_outputs(1308) <= inputs(100);
    layer0_outputs(1309) <= not(inputs(76));
    layer0_outputs(1310) <= not(inputs(255));
    layer0_outputs(1311) <= (inputs(154)) and not (inputs(230));
    layer0_outputs(1312) <= (inputs(252)) xor (inputs(187));
    layer0_outputs(1313) <= (inputs(58)) and not (inputs(32));
    layer0_outputs(1314) <= not(inputs(227));
    layer0_outputs(1315) <= not(inputs(108)) or (inputs(18));
    layer0_outputs(1316) <= inputs(121);
    layer0_outputs(1317) <= not(inputs(103)) or (inputs(162));
    layer0_outputs(1318) <= not(inputs(182));
    layer0_outputs(1319) <= inputs(159);
    layer0_outputs(1320) <= (inputs(128)) or (inputs(154));
    layer0_outputs(1321) <= not((inputs(6)) or (inputs(204)));
    layer0_outputs(1322) <= '0';
    layer0_outputs(1323) <= not(inputs(146));
    layer0_outputs(1324) <= (inputs(90)) and not (inputs(110));
    layer0_outputs(1325) <= inputs(30);
    layer0_outputs(1326) <= not((inputs(239)) or (inputs(147)));
    layer0_outputs(1327) <= not(inputs(89)) or (inputs(35));
    layer0_outputs(1328) <= inputs(179);
    layer0_outputs(1329) <= inputs(237);
    layer0_outputs(1330) <= not(inputs(55));
    layer0_outputs(1331) <= (inputs(185)) or (inputs(124));
    layer0_outputs(1332) <= (inputs(38)) or (inputs(8));
    layer0_outputs(1333) <= inputs(219);
    layer0_outputs(1334) <= not(inputs(246));
    layer0_outputs(1335) <= (inputs(7)) or (inputs(80));
    layer0_outputs(1336) <= not((inputs(19)) or (inputs(241)));
    layer0_outputs(1337) <= (inputs(24)) and (inputs(12));
    layer0_outputs(1338) <= '1';
    layer0_outputs(1339) <= not(inputs(137)) or (inputs(6));
    layer0_outputs(1340) <= (inputs(18)) xor (inputs(191));
    layer0_outputs(1341) <= not((inputs(139)) or (inputs(14)));
    layer0_outputs(1342) <= (inputs(151)) and not (inputs(189));
    layer0_outputs(1343) <= not(inputs(48)) or (inputs(250));
    layer0_outputs(1344) <= (inputs(212)) and not (inputs(4));
    layer0_outputs(1345) <= '0';
    layer0_outputs(1346) <= (inputs(247)) and not (inputs(145));
    layer0_outputs(1347) <= not((inputs(105)) or (inputs(103)));
    layer0_outputs(1348) <= inputs(173);
    layer0_outputs(1349) <= not(inputs(117));
    layer0_outputs(1350) <= inputs(97);
    layer0_outputs(1351) <= (inputs(181)) xor (inputs(227));
    layer0_outputs(1352) <= not((inputs(78)) or (inputs(219)));
    layer0_outputs(1353) <= (inputs(171)) and (inputs(41));
    layer0_outputs(1354) <= inputs(247);
    layer0_outputs(1355) <= not(inputs(118));
    layer0_outputs(1356) <= not(inputs(38));
    layer0_outputs(1357) <= inputs(228);
    layer0_outputs(1358) <= (inputs(233)) or (inputs(112));
    layer0_outputs(1359) <= not((inputs(209)) or (inputs(181)));
    layer0_outputs(1360) <= not((inputs(89)) or (inputs(16)));
    layer0_outputs(1361) <= (inputs(96)) or (inputs(130));
    layer0_outputs(1362) <= '0';
    layer0_outputs(1363) <= (inputs(92)) and not (inputs(98));
    layer0_outputs(1364) <= not((inputs(89)) or (inputs(236)));
    layer0_outputs(1365) <= not(inputs(117));
    layer0_outputs(1366) <= inputs(131);
    layer0_outputs(1367) <= inputs(47);
    layer0_outputs(1368) <= (inputs(151)) and not (inputs(29));
    layer0_outputs(1369) <= inputs(223);
    layer0_outputs(1370) <= not(inputs(40)) or (inputs(150));
    layer0_outputs(1371) <= not((inputs(114)) or (inputs(197)));
    layer0_outputs(1372) <= (inputs(72)) xor (inputs(244));
    layer0_outputs(1373) <= inputs(104);
    layer0_outputs(1374) <= not((inputs(110)) or (inputs(88)));
    layer0_outputs(1375) <= not((inputs(230)) or (inputs(194)));
    layer0_outputs(1376) <= (inputs(75)) and not (inputs(161));
    layer0_outputs(1377) <= (inputs(88)) and not (inputs(56));
    layer0_outputs(1378) <= not(inputs(74)) or (inputs(57));
    layer0_outputs(1379) <= inputs(132);
    layer0_outputs(1380) <= not(inputs(233));
    layer0_outputs(1381) <= not((inputs(132)) or (inputs(143)));
    layer0_outputs(1382) <= (inputs(96)) and not (inputs(171));
    layer0_outputs(1383) <= (inputs(117)) and not (inputs(224));
    layer0_outputs(1384) <= inputs(246);
    layer0_outputs(1385) <= inputs(234);
    layer0_outputs(1386) <= not(inputs(24));
    layer0_outputs(1387) <= (inputs(23)) and not (inputs(181));
    layer0_outputs(1388) <= not(inputs(230));
    layer0_outputs(1389) <= (inputs(252)) or (inputs(69));
    layer0_outputs(1390) <= (inputs(213)) and (inputs(61));
    layer0_outputs(1391) <= not((inputs(182)) or (inputs(254)));
    layer0_outputs(1392) <= (inputs(180)) and not (inputs(113));
    layer0_outputs(1393) <= inputs(148);
    layer0_outputs(1394) <= (inputs(107)) and not (inputs(245));
    layer0_outputs(1395) <= (inputs(11)) and not (inputs(222));
    layer0_outputs(1396) <= inputs(216);
    layer0_outputs(1397) <= not((inputs(52)) xor (inputs(144)));
    layer0_outputs(1398) <= not((inputs(159)) or (inputs(187)));
    layer0_outputs(1399) <= not(inputs(31));
    layer0_outputs(1400) <= not((inputs(208)) or (inputs(200)));
    layer0_outputs(1401) <= inputs(211);
    layer0_outputs(1402) <= (inputs(243)) and (inputs(240));
    layer0_outputs(1403) <= not((inputs(207)) or (inputs(150)));
    layer0_outputs(1404) <= (inputs(251)) or (inputs(131));
    layer0_outputs(1405) <= not(inputs(175)) or (inputs(41));
    layer0_outputs(1406) <= not(inputs(201)) or (inputs(201));
    layer0_outputs(1407) <= inputs(167);
    layer0_outputs(1408) <= not(inputs(246)) or (inputs(16));
    layer0_outputs(1409) <= not(inputs(237));
    layer0_outputs(1410) <= not(inputs(215));
    layer0_outputs(1411) <= not(inputs(225)) or (inputs(190));
    layer0_outputs(1412) <= inputs(152);
    layer0_outputs(1413) <= inputs(156);
    layer0_outputs(1414) <= inputs(255);
    layer0_outputs(1415) <= inputs(205);
    layer0_outputs(1416) <= not((inputs(138)) or (inputs(85)));
    layer0_outputs(1417) <= not((inputs(95)) or (inputs(81)));
    layer0_outputs(1418) <= (inputs(6)) and (inputs(58));
    layer0_outputs(1419) <= not(inputs(231));
    layer0_outputs(1420) <= not(inputs(254)) or (inputs(245));
    layer0_outputs(1421) <= not(inputs(173)) or (inputs(254));
    layer0_outputs(1422) <= (inputs(57)) and not (inputs(33));
    layer0_outputs(1423) <= not(inputs(138)) or (inputs(243));
    layer0_outputs(1424) <= not(inputs(130)) or (inputs(40));
    layer0_outputs(1425) <= inputs(246);
    layer0_outputs(1426) <= not((inputs(178)) or (inputs(230)));
    layer0_outputs(1427) <= not(inputs(120));
    layer0_outputs(1428) <= (inputs(198)) and not (inputs(59));
    layer0_outputs(1429) <= (inputs(130)) or (inputs(132));
    layer0_outputs(1430) <= (inputs(125)) and not (inputs(65));
    layer0_outputs(1431) <= inputs(75);
    layer0_outputs(1432) <= not(inputs(204)) or (inputs(79));
    layer0_outputs(1433) <= inputs(116);
    layer0_outputs(1434) <= '0';
    layer0_outputs(1435) <= not(inputs(98));
    layer0_outputs(1436) <= (inputs(203)) and not (inputs(137));
    layer0_outputs(1437) <= (inputs(15)) or (inputs(237));
    layer0_outputs(1438) <= '1';
    layer0_outputs(1439) <= not((inputs(1)) or (inputs(65)));
    layer0_outputs(1440) <= (inputs(108)) or (inputs(241));
    layer0_outputs(1441) <= '0';
    layer0_outputs(1442) <= not((inputs(232)) or (inputs(116)));
    layer0_outputs(1443) <= not((inputs(85)) or (inputs(193)));
    layer0_outputs(1444) <= (inputs(156)) or (inputs(4));
    layer0_outputs(1445) <= not((inputs(148)) and (inputs(220)));
    layer0_outputs(1446) <= inputs(168);
    layer0_outputs(1447) <= not((inputs(202)) or (inputs(3)));
    layer0_outputs(1448) <= (inputs(33)) or (inputs(145));
    layer0_outputs(1449) <= not(inputs(243));
    layer0_outputs(1450) <= (inputs(103)) and not (inputs(180));
    layer0_outputs(1451) <= not(inputs(152));
    layer0_outputs(1452) <= not((inputs(162)) or (inputs(194)));
    layer0_outputs(1453) <= not(inputs(140));
    layer0_outputs(1454) <= not(inputs(40));
    layer0_outputs(1455) <= not(inputs(228));
    layer0_outputs(1456) <= (inputs(43)) and not (inputs(240));
    layer0_outputs(1457) <= (inputs(162)) or (inputs(136));
    layer0_outputs(1458) <= not(inputs(95)) or (inputs(155));
    layer0_outputs(1459) <= not(inputs(216));
    layer0_outputs(1460) <= not(inputs(228)) or (inputs(30));
    layer0_outputs(1461) <= (inputs(219)) or (inputs(222));
    layer0_outputs(1462) <= inputs(153);
    layer0_outputs(1463) <= '1';
    layer0_outputs(1464) <= inputs(214);
    layer0_outputs(1465) <= not(inputs(55));
    layer0_outputs(1466) <= not(inputs(123));
    layer0_outputs(1467) <= '0';
    layer0_outputs(1468) <= not(inputs(107)) or (inputs(83));
    layer0_outputs(1469) <= inputs(51);
    layer0_outputs(1470) <= (inputs(219)) or (inputs(47));
    layer0_outputs(1471) <= (inputs(120)) and not (inputs(6));
    layer0_outputs(1472) <= inputs(4);
    layer0_outputs(1473) <= not(inputs(13));
    layer0_outputs(1474) <= not(inputs(136));
    layer0_outputs(1475) <= not((inputs(164)) or (inputs(162)));
    layer0_outputs(1476) <= (inputs(252)) or (inputs(150));
    layer0_outputs(1477) <= inputs(86);
    layer0_outputs(1478) <= not(inputs(94));
    layer0_outputs(1479) <= (inputs(125)) or (inputs(166));
    layer0_outputs(1480) <= inputs(76);
    layer0_outputs(1481) <= not(inputs(191)) or (inputs(249));
    layer0_outputs(1482) <= not((inputs(17)) or (inputs(154)));
    layer0_outputs(1483) <= not((inputs(127)) xor (inputs(151)));
    layer0_outputs(1484) <= inputs(223);
    layer0_outputs(1485) <= not((inputs(161)) or (inputs(19)));
    layer0_outputs(1486) <= not(inputs(68)) or (inputs(172));
    layer0_outputs(1487) <= not((inputs(174)) or (inputs(147)));
    layer0_outputs(1488) <= inputs(53);
    layer0_outputs(1489) <= not((inputs(97)) or (inputs(102)));
    layer0_outputs(1490) <= not(inputs(18));
    layer0_outputs(1491) <= not((inputs(246)) or (inputs(80)));
    layer0_outputs(1492) <= (inputs(239)) or (inputs(187));
    layer0_outputs(1493) <= (inputs(167)) or (inputs(169));
    layer0_outputs(1494) <= (inputs(127)) or (inputs(210));
    layer0_outputs(1495) <= (inputs(166)) and not (inputs(96));
    layer0_outputs(1496) <= not(inputs(83));
    layer0_outputs(1497) <= (inputs(138)) or (inputs(48));
    layer0_outputs(1498) <= not(inputs(153));
    layer0_outputs(1499) <= (inputs(159)) or (inputs(225));
    layer0_outputs(1500) <= (inputs(174)) or (inputs(245));
    layer0_outputs(1501) <= not(inputs(149));
    layer0_outputs(1502) <= (inputs(226)) or (inputs(177));
    layer0_outputs(1503) <= (inputs(108)) and not (inputs(237));
    layer0_outputs(1504) <= not((inputs(241)) or (inputs(168)));
    layer0_outputs(1505) <= not(inputs(230)) or (inputs(190));
    layer0_outputs(1506) <= not(inputs(31));
    layer0_outputs(1507) <= not(inputs(26)) or (inputs(102));
    layer0_outputs(1508) <= inputs(173);
    layer0_outputs(1509) <= (inputs(189)) and not (inputs(73));
    layer0_outputs(1510) <= not(inputs(228));
    layer0_outputs(1511) <= '1';
    layer0_outputs(1512) <= (inputs(67)) or (inputs(252));
    layer0_outputs(1513) <= not((inputs(225)) or (inputs(161)));
    layer0_outputs(1514) <= not(inputs(84));
    layer0_outputs(1515) <= not(inputs(127));
    layer0_outputs(1516) <= not((inputs(20)) or (inputs(148)));
    layer0_outputs(1517) <= not((inputs(2)) and (inputs(159)));
    layer0_outputs(1518) <= inputs(84);
    layer0_outputs(1519) <= inputs(156);
    layer0_outputs(1520) <= not((inputs(146)) or (inputs(171)));
    layer0_outputs(1521) <= not((inputs(103)) or (inputs(103)));
    layer0_outputs(1522) <= not((inputs(70)) or (inputs(179)));
    layer0_outputs(1523) <= (inputs(170)) and not (inputs(124));
    layer0_outputs(1524) <= not(inputs(3));
    layer0_outputs(1525) <= not(inputs(253)) or (inputs(234));
    layer0_outputs(1526) <= not((inputs(141)) and (inputs(138)));
    layer0_outputs(1527) <= (inputs(76)) or (inputs(239));
    layer0_outputs(1528) <= (inputs(165)) and not (inputs(29));
    layer0_outputs(1529) <= not((inputs(92)) or (inputs(48)));
    layer0_outputs(1530) <= not(inputs(112));
    layer0_outputs(1531) <= not((inputs(211)) or (inputs(204)));
    layer0_outputs(1532) <= not(inputs(184));
    layer0_outputs(1533) <= not((inputs(227)) or (inputs(136)));
    layer0_outputs(1534) <= (inputs(35)) and not (inputs(24));
    layer0_outputs(1535) <= not(inputs(121));
    layer0_outputs(1536) <= not(inputs(12)) or (inputs(144));
    layer0_outputs(1537) <= not((inputs(188)) or (inputs(5)));
    layer0_outputs(1538) <= not(inputs(69));
    layer0_outputs(1539) <= inputs(151);
    layer0_outputs(1540) <= inputs(52);
    layer0_outputs(1541) <= not(inputs(180));
    layer0_outputs(1542) <= not(inputs(212));
    layer0_outputs(1543) <= (inputs(244)) and not (inputs(189));
    layer0_outputs(1544) <= (inputs(194)) or (inputs(208));
    layer0_outputs(1545) <= '1';
    layer0_outputs(1546) <= not((inputs(186)) or (inputs(26)));
    layer0_outputs(1547) <= inputs(82);
    layer0_outputs(1548) <= '0';
    layer0_outputs(1549) <= (inputs(206)) xor (inputs(140));
    layer0_outputs(1550) <= (inputs(89)) and not (inputs(55));
    layer0_outputs(1551) <= inputs(179);
    layer0_outputs(1552) <= not((inputs(241)) xor (inputs(13)));
    layer0_outputs(1553) <= not(inputs(26));
    layer0_outputs(1554) <= not(inputs(179)) or (inputs(153));
    layer0_outputs(1555) <= (inputs(88)) and not (inputs(157));
    layer0_outputs(1556) <= not((inputs(80)) or (inputs(238)));
    layer0_outputs(1557) <= (inputs(158)) or (inputs(191));
    layer0_outputs(1558) <= inputs(76);
    layer0_outputs(1559) <= '0';
    layer0_outputs(1560) <= not(inputs(180));
    layer0_outputs(1561) <= not(inputs(22));
    layer0_outputs(1562) <= inputs(15);
    layer0_outputs(1563) <= inputs(244);
    layer0_outputs(1564) <= not(inputs(170));
    layer0_outputs(1565) <= not(inputs(84)) or (inputs(123));
    layer0_outputs(1566) <= inputs(82);
    layer0_outputs(1567) <= not(inputs(200));
    layer0_outputs(1568) <= (inputs(135)) and not (inputs(120));
    layer0_outputs(1569) <= (inputs(197)) or (inputs(176));
    layer0_outputs(1570) <= not(inputs(67));
    layer0_outputs(1571) <= inputs(43);
    layer0_outputs(1572) <= not(inputs(246)) or (inputs(174));
    layer0_outputs(1573) <= (inputs(67)) and not (inputs(189));
    layer0_outputs(1574) <= inputs(208);
    layer0_outputs(1575) <= '1';
    layer0_outputs(1576) <= inputs(39);
    layer0_outputs(1577) <= not((inputs(20)) xor (inputs(52)));
    layer0_outputs(1578) <= (inputs(0)) or (inputs(222));
    layer0_outputs(1579) <= not((inputs(164)) or (inputs(147)));
    layer0_outputs(1580) <= not((inputs(102)) or (inputs(98)));
    layer0_outputs(1581) <= not(inputs(13));
    layer0_outputs(1582) <= inputs(58);
    layer0_outputs(1583) <= (inputs(44)) and not (inputs(245));
    layer0_outputs(1584) <= not(inputs(146));
    layer0_outputs(1585) <= '0';
    layer0_outputs(1586) <= (inputs(154)) or (inputs(237));
    layer0_outputs(1587) <= not(inputs(98));
    layer0_outputs(1588) <= inputs(209);
    layer0_outputs(1589) <= inputs(117);
    layer0_outputs(1590) <= not((inputs(118)) or (inputs(69)));
    layer0_outputs(1591) <= not(inputs(230)) or (inputs(47));
    layer0_outputs(1592) <= not((inputs(90)) or (inputs(180)));
    layer0_outputs(1593) <= not(inputs(108));
    layer0_outputs(1594) <= (inputs(94)) or (inputs(206));
    layer0_outputs(1595) <= not((inputs(163)) or (inputs(64)));
    layer0_outputs(1596) <= not((inputs(182)) or (inputs(5)));
    layer0_outputs(1597) <= (inputs(24)) xor (inputs(110));
    layer0_outputs(1598) <= not(inputs(138)) or (inputs(142));
    layer0_outputs(1599) <= inputs(100);
    layer0_outputs(1600) <= inputs(106);
    layer0_outputs(1601) <= not((inputs(34)) or (inputs(135)));
    layer0_outputs(1602) <= inputs(229);
    layer0_outputs(1603) <= (inputs(138)) and not (inputs(194));
    layer0_outputs(1604) <= inputs(168);
    layer0_outputs(1605) <= not(inputs(24));
    layer0_outputs(1606) <= not(inputs(207)) or (inputs(224));
    layer0_outputs(1607) <= inputs(164);
    layer0_outputs(1608) <= not(inputs(183));
    layer0_outputs(1609) <= inputs(8);
    layer0_outputs(1610) <= not(inputs(45));
    layer0_outputs(1611) <= inputs(242);
    layer0_outputs(1612) <= not((inputs(205)) or (inputs(86)));
    layer0_outputs(1613) <= (inputs(0)) or (inputs(16));
    layer0_outputs(1614) <= not(inputs(221)) or (inputs(81));
    layer0_outputs(1615) <= (inputs(255)) or (inputs(237));
    layer0_outputs(1616) <= inputs(68);
    layer0_outputs(1617) <= not(inputs(164));
    layer0_outputs(1618) <= (inputs(112)) and (inputs(144));
    layer0_outputs(1619) <= not((inputs(218)) or (inputs(191)));
    layer0_outputs(1620) <= inputs(228);
    layer0_outputs(1621) <= inputs(134);
    layer0_outputs(1622) <= not((inputs(149)) or (inputs(166)));
    layer0_outputs(1623) <= inputs(183);
    layer0_outputs(1624) <= not((inputs(99)) or (inputs(218)));
    layer0_outputs(1625) <= (inputs(39)) xor (inputs(7));
    layer0_outputs(1626) <= inputs(127);
    layer0_outputs(1627) <= inputs(137);
    layer0_outputs(1628) <= '0';
    layer0_outputs(1629) <= not(inputs(8));
    layer0_outputs(1630) <= not(inputs(21)) or (inputs(238));
    layer0_outputs(1631) <= inputs(202);
    layer0_outputs(1632) <= (inputs(37)) and not (inputs(107));
    layer0_outputs(1633) <= not((inputs(63)) or (inputs(101)));
    layer0_outputs(1634) <= '1';
    layer0_outputs(1635) <= (inputs(100)) or (inputs(102));
    layer0_outputs(1636) <= not(inputs(166));
    layer0_outputs(1637) <= (inputs(23)) and not (inputs(220));
    layer0_outputs(1638) <= not(inputs(210));
    layer0_outputs(1639) <= not(inputs(109)) or (inputs(130));
    layer0_outputs(1640) <= not(inputs(106));
    layer0_outputs(1641) <= not((inputs(215)) or (inputs(231)));
    layer0_outputs(1642) <= inputs(213);
    layer0_outputs(1643) <= inputs(227);
    layer0_outputs(1644) <= not(inputs(84));
    layer0_outputs(1645) <= not((inputs(76)) or (inputs(48)));
    layer0_outputs(1646) <= not(inputs(129));
    layer0_outputs(1647) <= not((inputs(131)) or (inputs(67)));
    layer0_outputs(1648) <= (inputs(38)) and (inputs(80));
    layer0_outputs(1649) <= not(inputs(251));
    layer0_outputs(1650) <= inputs(153);
    layer0_outputs(1651) <= '0';
    layer0_outputs(1652) <= not(inputs(38));
    layer0_outputs(1653) <= not((inputs(37)) or (inputs(70)));
    layer0_outputs(1654) <= not((inputs(15)) or (inputs(238)));
    layer0_outputs(1655) <= '0';
    layer0_outputs(1656) <= not(inputs(24));
    layer0_outputs(1657) <= '0';
    layer0_outputs(1658) <= (inputs(213)) xor (inputs(196));
    layer0_outputs(1659) <= not((inputs(75)) or (inputs(142)));
    layer0_outputs(1660) <= not(inputs(136)) or (inputs(223));
    layer0_outputs(1661) <= inputs(36);
    layer0_outputs(1662) <= not(inputs(247)) or (inputs(29));
    layer0_outputs(1663) <= not(inputs(230));
    layer0_outputs(1664) <= '1';
    layer0_outputs(1665) <= not(inputs(121)) or (inputs(64));
    layer0_outputs(1666) <= not((inputs(169)) or (inputs(24)));
    layer0_outputs(1667) <= not((inputs(201)) or (inputs(177)));
    layer0_outputs(1668) <= not((inputs(175)) or (inputs(213)));
    layer0_outputs(1669) <= (inputs(119)) and not (inputs(149));
    layer0_outputs(1670) <= (inputs(140)) or (inputs(156));
    layer0_outputs(1671) <= inputs(145);
    layer0_outputs(1672) <= not(inputs(99)) or (inputs(66));
    layer0_outputs(1673) <= inputs(226);
    layer0_outputs(1674) <= not(inputs(142));
    layer0_outputs(1675) <= not(inputs(106));
    layer0_outputs(1676) <= not(inputs(37)) or (inputs(46));
    layer0_outputs(1677) <= inputs(207);
    layer0_outputs(1678) <= (inputs(95)) or (inputs(177));
    layer0_outputs(1679) <= not(inputs(163));
    layer0_outputs(1680) <= not(inputs(137)) or (inputs(190));
    layer0_outputs(1681) <= '1';
    layer0_outputs(1682) <= not((inputs(192)) or (inputs(241)));
    layer0_outputs(1683) <= (inputs(25)) xor (inputs(251));
    layer0_outputs(1684) <= inputs(134);
    layer0_outputs(1685) <= (inputs(25)) and not (inputs(14));
    layer0_outputs(1686) <= not(inputs(187)) or (inputs(169));
    layer0_outputs(1687) <= not(inputs(178));
    layer0_outputs(1688) <= not(inputs(233)) or (inputs(130));
    layer0_outputs(1689) <= not((inputs(81)) xor (inputs(71)));
    layer0_outputs(1690) <= inputs(98);
    layer0_outputs(1691) <= not(inputs(231));
    layer0_outputs(1692) <= (inputs(95)) xor (inputs(59));
    layer0_outputs(1693) <= inputs(84);
    layer0_outputs(1694) <= not((inputs(91)) or (inputs(240)));
    layer0_outputs(1695) <= not(inputs(182));
    layer0_outputs(1696) <= (inputs(248)) or (inputs(115));
    layer0_outputs(1697) <= inputs(122);
    layer0_outputs(1698) <= not(inputs(114));
    layer0_outputs(1699) <= inputs(119);
    layer0_outputs(1700) <= (inputs(53)) and not (inputs(173));
    layer0_outputs(1701) <= not(inputs(23)) or (inputs(195));
    layer0_outputs(1702) <= (inputs(115)) and not (inputs(223));
    layer0_outputs(1703) <= (inputs(192)) or (inputs(1));
    layer0_outputs(1704) <= inputs(79);
    layer0_outputs(1705) <= (inputs(130)) or (inputs(169));
    layer0_outputs(1706) <= inputs(155);
    layer0_outputs(1707) <= not(inputs(80));
    layer0_outputs(1708) <= (inputs(107)) and not (inputs(153));
    layer0_outputs(1709) <= not(inputs(141));
    layer0_outputs(1710) <= not(inputs(134));
    layer0_outputs(1711) <= not((inputs(151)) xor (inputs(139)));
    layer0_outputs(1712) <= not(inputs(192));
    layer0_outputs(1713) <= (inputs(70)) and not (inputs(32));
    layer0_outputs(1714) <= not(inputs(45));
    layer0_outputs(1715) <= not((inputs(147)) or (inputs(62)));
    layer0_outputs(1716) <= (inputs(242)) or (inputs(46));
    layer0_outputs(1717) <= '0';
    layer0_outputs(1718) <= not(inputs(193));
    layer0_outputs(1719) <= inputs(90);
    layer0_outputs(1720) <= not(inputs(202));
    layer0_outputs(1721) <= not(inputs(199));
    layer0_outputs(1722) <= (inputs(246)) and not (inputs(16));
    layer0_outputs(1723) <= inputs(181);
    layer0_outputs(1724) <= inputs(105);
    layer0_outputs(1725) <= not(inputs(216));
    layer0_outputs(1726) <= inputs(140);
    layer0_outputs(1727) <= not(inputs(179));
    layer0_outputs(1728) <= (inputs(221)) and not (inputs(13));
    layer0_outputs(1729) <= not(inputs(36));
    layer0_outputs(1730) <= not(inputs(60));
    layer0_outputs(1731) <= inputs(186);
    layer0_outputs(1732) <= (inputs(18)) or (inputs(202));
    layer0_outputs(1733) <= not(inputs(2));
    layer0_outputs(1734) <= (inputs(119)) and (inputs(21));
    layer0_outputs(1735) <= not(inputs(163));
    layer0_outputs(1736) <= not((inputs(49)) or (inputs(47)));
    layer0_outputs(1737) <= not((inputs(99)) or (inputs(179)));
    layer0_outputs(1738) <= inputs(103);
    layer0_outputs(1739) <= not((inputs(190)) xor (inputs(34)));
    layer0_outputs(1740) <= not((inputs(131)) or (inputs(143)));
    layer0_outputs(1741) <= inputs(75);
    layer0_outputs(1742) <= (inputs(111)) or (inputs(183));
    layer0_outputs(1743) <= not((inputs(217)) or (inputs(240)));
    layer0_outputs(1744) <= (inputs(9)) and not (inputs(141));
    layer0_outputs(1745) <= (inputs(160)) or (inputs(44));
    layer0_outputs(1746) <= (inputs(129)) xor (inputs(148));
    layer0_outputs(1747) <= not(inputs(100)) or (inputs(212));
    layer0_outputs(1748) <= inputs(68);
    layer0_outputs(1749) <= not(inputs(45));
    layer0_outputs(1750) <= not(inputs(101));
    layer0_outputs(1751) <= not(inputs(165));
    layer0_outputs(1752) <= not(inputs(204));
    layer0_outputs(1753) <= not((inputs(180)) or (inputs(188)));
    layer0_outputs(1754) <= not(inputs(106)) or (inputs(233));
    layer0_outputs(1755) <= (inputs(249)) and not (inputs(173));
    layer0_outputs(1756) <= (inputs(113)) or (inputs(70));
    layer0_outputs(1757) <= inputs(69);
    layer0_outputs(1758) <= not(inputs(124));
    layer0_outputs(1759) <= (inputs(190)) or (inputs(231));
    layer0_outputs(1760) <= inputs(155);
    layer0_outputs(1761) <= (inputs(8)) and not (inputs(214));
    layer0_outputs(1762) <= not(inputs(39));
    layer0_outputs(1763) <= '0';
    layer0_outputs(1764) <= not((inputs(151)) and (inputs(231)));
    layer0_outputs(1765) <= not((inputs(84)) or (inputs(130)));
    layer0_outputs(1766) <= inputs(99);
    layer0_outputs(1767) <= (inputs(136)) and not (inputs(224));
    layer0_outputs(1768) <= not((inputs(14)) or (inputs(222)));
    layer0_outputs(1769) <= not(inputs(93));
    layer0_outputs(1770) <= (inputs(253)) xor (inputs(68));
    layer0_outputs(1771) <= (inputs(141)) and not (inputs(14));
    layer0_outputs(1772) <= not((inputs(4)) or (inputs(50)));
    layer0_outputs(1773) <= inputs(164);
    layer0_outputs(1774) <= not(inputs(139)) or (inputs(227));
    layer0_outputs(1775) <= not(inputs(125));
    layer0_outputs(1776) <= inputs(213);
    layer0_outputs(1777) <= inputs(60);
    layer0_outputs(1778) <= not((inputs(211)) or (inputs(66)));
    layer0_outputs(1779) <= (inputs(119)) or (inputs(251));
    layer0_outputs(1780) <= not(inputs(173)) or (inputs(65));
    layer0_outputs(1781) <= (inputs(26)) or (inputs(254));
    layer0_outputs(1782) <= inputs(131);
    layer0_outputs(1783) <= not(inputs(101));
    layer0_outputs(1784) <= inputs(117);
    layer0_outputs(1785) <= (inputs(73)) or (inputs(79));
    layer0_outputs(1786) <= not(inputs(179));
    layer0_outputs(1787) <= inputs(164);
    layer0_outputs(1788) <= inputs(88);
    layer0_outputs(1789) <= not(inputs(122)) or (inputs(114));
    layer0_outputs(1790) <= inputs(135);
    layer0_outputs(1791) <= (inputs(131)) or (inputs(138));
    layer0_outputs(1792) <= not(inputs(83)) or (inputs(175));
    layer0_outputs(1793) <= not(inputs(112)) or (inputs(204));
    layer0_outputs(1794) <= not(inputs(229)) or (inputs(128));
    layer0_outputs(1795) <= not(inputs(13)) or (inputs(226));
    layer0_outputs(1796) <= inputs(101);
    layer0_outputs(1797) <= not((inputs(187)) or (inputs(160)));
    layer0_outputs(1798) <= not(inputs(232)) or (inputs(224));
    layer0_outputs(1799) <= inputs(61);
    layer0_outputs(1800) <= (inputs(70)) and not (inputs(253));
    layer0_outputs(1801) <= (inputs(130)) and not (inputs(103));
    layer0_outputs(1802) <= not((inputs(192)) or (inputs(208)));
    layer0_outputs(1803) <= inputs(193);
    layer0_outputs(1804) <= not(inputs(106));
    layer0_outputs(1805) <= (inputs(160)) and not (inputs(48));
    layer0_outputs(1806) <= not(inputs(159));
    layer0_outputs(1807) <= (inputs(11)) xor (inputs(20));
    layer0_outputs(1808) <= not((inputs(122)) or (inputs(205)));
    layer0_outputs(1809) <= not((inputs(255)) xor (inputs(34)));
    layer0_outputs(1810) <= '1';
    layer0_outputs(1811) <= inputs(56);
    layer0_outputs(1812) <= (inputs(172)) or (inputs(97));
    layer0_outputs(1813) <= not(inputs(199)) or (inputs(99));
    layer0_outputs(1814) <= not(inputs(109));
    layer0_outputs(1815) <= (inputs(1)) or (inputs(183));
    layer0_outputs(1816) <= inputs(207);
    layer0_outputs(1817) <= '1';
    layer0_outputs(1818) <= not((inputs(64)) or (inputs(186)));
    layer0_outputs(1819) <= not(inputs(15)) or (inputs(78));
    layer0_outputs(1820) <= not(inputs(40)) or (inputs(31));
    layer0_outputs(1821) <= inputs(87);
    layer0_outputs(1822) <= not(inputs(53));
    layer0_outputs(1823) <= not(inputs(130)) or (inputs(19));
    layer0_outputs(1824) <= not((inputs(11)) or (inputs(128)));
    layer0_outputs(1825) <= '1';
    layer0_outputs(1826) <= (inputs(105)) and not (inputs(94));
    layer0_outputs(1827) <= not(inputs(101));
    layer0_outputs(1828) <= inputs(115);
    layer0_outputs(1829) <= not((inputs(65)) xor (inputs(52)));
    layer0_outputs(1830) <= (inputs(83)) or (inputs(95));
    layer0_outputs(1831) <= not((inputs(172)) xor (inputs(236)));
    layer0_outputs(1832) <= not(inputs(22)) or (inputs(27));
    layer0_outputs(1833) <= (inputs(227)) or (inputs(101));
    layer0_outputs(1834) <= not(inputs(93));
    layer0_outputs(1835) <= inputs(116);
    layer0_outputs(1836) <= not(inputs(151));
    layer0_outputs(1837) <= (inputs(45)) or (inputs(122));
    layer0_outputs(1838) <= not(inputs(200));
    layer0_outputs(1839) <= not(inputs(115)) or (inputs(146));
    layer0_outputs(1840) <= (inputs(92)) or (inputs(77));
    layer0_outputs(1841) <= not((inputs(165)) xor (inputs(211)));
    layer0_outputs(1842) <= inputs(123);
    layer0_outputs(1843) <= not(inputs(121)) or (inputs(33));
    layer0_outputs(1844) <= inputs(165);
    layer0_outputs(1845) <= not(inputs(91)) or (inputs(212));
    layer0_outputs(1846) <= not(inputs(22));
    layer0_outputs(1847) <= not(inputs(85)) or (inputs(111));
    layer0_outputs(1848) <= not((inputs(32)) or (inputs(3)));
    layer0_outputs(1849) <= inputs(193);
    layer0_outputs(1850) <= (inputs(1)) or (inputs(73));
    layer0_outputs(1851) <= not(inputs(23));
    layer0_outputs(1852) <= not(inputs(84));
    layer0_outputs(1853) <= (inputs(223)) or (inputs(22));
    layer0_outputs(1854) <= not(inputs(134)) or (inputs(33));
    layer0_outputs(1855) <= (inputs(245)) xor (inputs(198));
    layer0_outputs(1856) <= not(inputs(12)) or (inputs(34));
    layer0_outputs(1857) <= not(inputs(51)) or (inputs(141));
    layer0_outputs(1858) <= not(inputs(183));
    layer0_outputs(1859) <= not((inputs(53)) or (inputs(176)));
    layer0_outputs(1860) <= (inputs(229)) or (inputs(3));
    layer0_outputs(1861) <= not(inputs(169));
    layer0_outputs(1862) <= not(inputs(216)) or (inputs(33));
    layer0_outputs(1863) <= (inputs(191)) or (inputs(226));
    layer0_outputs(1864) <= not(inputs(27));
    layer0_outputs(1865) <= not((inputs(112)) or (inputs(211)));
    layer0_outputs(1866) <= not((inputs(157)) or (inputs(179)));
    layer0_outputs(1867) <= not((inputs(82)) or (inputs(232)));
    layer0_outputs(1868) <= not(inputs(69)) or (inputs(238));
    layer0_outputs(1869) <= (inputs(23)) and not (inputs(113));
    layer0_outputs(1870) <= '0';
    layer0_outputs(1871) <= not((inputs(127)) or (inputs(194)));
    layer0_outputs(1872) <= (inputs(106)) or (inputs(135));
    layer0_outputs(1873) <= (inputs(84)) xor (inputs(96));
    layer0_outputs(1874) <= (inputs(155)) and not (inputs(196));
    layer0_outputs(1875) <= not((inputs(226)) or (inputs(180)));
    layer0_outputs(1876) <= not((inputs(183)) or (inputs(122)));
    layer0_outputs(1877) <= (inputs(157)) and (inputs(154));
    layer0_outputs(1878) <= inputs(105);
    layer0_outputs(1879) <= not(inputs(23));
    layer0_outputs(1880) <= (inputs(160)) or (inputs(248));
    layer0_outputs(1881) <= not(inputs(219));
    layer0_outputs(1882) <= not(inputs(227));
    layer0_outputs(1883) <= inputs(100);
    layer0_outputs(1884) <= not(inputs(114));
    layer0_outputs(1885) <= not((inputs(107)) or (inputs(182)));
    layer0_outputs(1886) <= (inputs(119)) or (inputs(63));
    layer0_outputs(1887) <= not(inputs(20)) or (inputs(127));
    layer0_outputs(1888) <= not(inputs(212)) or (inputs(130));
    layer0_outputs(1889) <= not(inputs(165));
    layer0_outputs(1890) <= '0';
    layer0_outputs(1891) <= not(inputs(53)) or (inputs(221));
    layer0_outputs(1892) <= (inputs(46)) or (inputs(74));
    layer0_outputs(1893) <= (inputs(242)) and not (inputs(159));
    layer0_outputs(1894) <= not((inputs(204)) or (inputs(65)));
    layer0_outputs(1895) <= not(inputs(87)) or (inputs(89));
    layer0_outputs(1896) <= (inputs(76)) or (inputs(209));
    layer0_outputs(1897) <= not(inputs(246)) or (inputs(253));
    layer0_outputs(1898) <= not(inputs(104));
    layer0_outputs(1899) <= (inputs(97)) or (inputs(208));
    layer0_outputs(1900) <= not((inputs(222)) or (inputs(204)));
    layer0_outputs(1901) <= (inputs(161)) or (inputs(204));
    layer0_outputs(1902) <= not(inputs(113));
    layer0_outputs(1903) <= not(inputs(93));
    layer0_outputs(1904) <= inputs(247);
    layer0_outputs(1905) <= (inputs(57)) or (inputs(189));
    layer0_outputs(1906) <= (inputs(128)) or (inputs(172));
    layer0_outputs(1907) <= (inputs(24)) or (inputs(95));
    layer0_outputs(1908) <= not(inputs(117)) or (inputs(70));
    layer0_outputs(1909) <= inputs(99);
    layer0_outputs(1910) <= inputs(211);
    layer0_outputs(1911) <= not(inputs(150));
    layer0_outputs(1912) <= not((inputs(3)) xor (inputs(49)));
    layer0_outputs(1913) <= (inputs(32)) xor (inputs(92));
    layer0_outputs(1914) <= (inputs(105)) and not (inputs(126));
    layer0_outputs(1915) <= '0';
    layer0_outputs(1916) <= not(inputs(178));
    layer0_outputs(1917) <= not(inputs(168)) or (inputs(232));
    layer0_outputs(1918) <= (inputs(253)) and not (inputs(207));
    layer0_outputs(1919) <= not(inputs(141));
    layer0_outputs(1920) <= (inputs(22)) or (inputs(142));
    layer0_outputs(1921) <= inputs(27);
    layer0_outputs(1922) <= (inputs(156)) or (inputs(220));
    layer0_outputs(1923) <= not(inputs(130));
    layer0_outputs(1924) <= not((inputs(224)) or (inputs(118)));
    layer0_outputs(1925) <= (inputs(134)) or (inputs(63));
    layer0_outputs(1926) <= inputs(181);
    layer0_outputs(1927) <= (inputs(0)) and (inputs(168));
    layer0_outputs(1928) <= inputs(38);
    layer0_outputs(1929) <= not((inputs(111)) or (inputs(197)));
    layer0_outputs(1930) <= (inputs(13)) and not (inputs(61));
    layer0_outputs(1931) <= not(inputs(215)) or (inputs(10));
    layer0_outputs(1932) <= not((inputs(69)) or (inputs(77)));
    layer0_outputs(1933) <= inputs(162);
    layer0_outputs(1934) <= (inputs(74)) and not (inputs(144));
    layer0_outputs(1935) <= (inputs(145)) or (inputs(71));
    layer0_outputs(1936) <= not((inputs(197)) or (inputs(174)));
    layer0_outputs(1937) <= not((inputs(243)) or (inputs(48)));
    layer0_outputs(1938) <= not(inputs(119));
    layer0_outputs(1939) <= not((inputs(145)) or (inputs(163)));
    layer0_outputs(1940) <= not(inputs(118)) or (inputs(156));
    layer0_outputs(1941) <= (inputs(180)) and (inputs(180));
    layer0_outputs(1942) <= inputs(89);
    layer0_outputs(1943) <= not((inputs(156)) or (inputs(115)));
    layer0_outputs(1944) <= not(inputs(125));
    layer0_outputs(1945) <= not(inputs(165));
    layer0_outputs(1946) <= (inputs(54)) and (inputs(214));
    layer0_outputs(1947) <= not((inputs(94)) or (inputs(60)));
    layer0_outputs(1948) <= (inputs(125)) or (inputs(219));
    layer0_outputs(1949) <= not(inputs(100));
    layer0_outputs(1950) <= not(inputs(205));
    layer0_outputs(1951) <= not((inputs(124)) or (inputs(26)));
    layer0_outputs(1952) <= not(inputs(166)) or (inputs(102));
    layer0_outputs(1953) <= inputs(237);
    layer0_outputs(1954) <= not(inputs(231));
    layer0_outputs(1955) <= (inputs(29)) or (inputs(209));
    layer0_outputs(1956) <= not(inputs(60)) or (inputs(192));
    layer0_outputs(1957) <= inputs(195);
    layer0_outputs(1958) <= not((inputs(10)) or (inputs(223)));
    layer0_outputs(1959) <= not(inputs(117));
    layer0_outputs(1960) <= not(inputs(135)) or (inputs(187));
    layer0_outputs(1961) <= not(inputs(247));
    layer0_outputs(1962) <= (inputs(116)) or (inputs(158));
    layer0_outputs(1963) <= not(inputs(55));
    layer0_outputs(1964) <= (inputs(186)) and not (inputs(50));
    layer0_outputs(1965) <= not((inputs(218)) and (inputs(215)));
    layer0_outputs(1966) <= inputs(106);
    layer0_outputs(1967) <= inputs(39);
    layer0_outputs(1968) <= not((inputs(223)) or (inputs(124)));
    layer0_outputs(1969) <= (inputs(253)) or (inputs(218));
    layer0_outputs(1970) <= not(inputs(50)) or (inputs(31));
    layer0_outputs(1971) <= not(inputs(249));
    layer0_outputs(1972) <= not(inputs(128)) or (inputs(223));
    layer0_outputs(1973) <= (inputs(250)) and not (inputs(21));
    layer0_outputs(1974) <= not(inputs(119)) or (inputs(161));
    layer0_outputs(1975) <= not((inputs(93)) or (inputs(95)));
    layer0_outputs(1976) <= inputs(109);
    layer0_outputs(1977) <= not(inputs(115));
    layer0_outputs(1978) <= inputs(40);
    layer0_outputs(1979) <= not(inputs(67)) or (inputs(18));
    layer0_outputs(1980) <= (inputs(209)) or (inputs(126));
    layer0_outputs(1981) <= not((inputs(249)) and (inputs(58)));
    layer0_outputs(1982) <= '1';
    layer0_outputs(1983) <= (inputs(132)) or (inputs(114));
    layer0_outputs(1984) <= (inputs(85)) and not (inputs(19));
    layer0_outputs(1985) <= inputs(78);
    layer0_outputs(1986) <= not(inputs(187)) or (inputs(111));
    layer0_outputs(1987) <= not(inputs(209));
    layer0_outputs(1988) <= (inputs(2)) and not (inputs(222));
    layer0_outputs(1989) <= inputs(43);
    layer0_outputs(1990) <= (inputs(190)) or (inputs(144));
    layer0_outputs(1991) <= (inputs(214)) and not (inputs(156));
    layer0_outputs(1992) <= (inputs(134)) and not (inputs(17));
    layer0_outputs(1993) <= not(inputs(28)) or (inputs(208));
    layer0_outputs(1994) <= (inputs(210)) and not (inputs(215));
    layer0_outputs(1995) <= inputs(39);
    layer0_outputs(1996) <= (inputs(6)) and not (inputs(151));
    layer0_outputs(1997) <= not((inputs(180)) or (inputs(195)));
    layer0_outputs(1998) <= (inputs(200)) or (inputs(132));
    layer0_outputs(1999) <= inputs(104);
    layer0_outputs(2000) <= inputs(56);
    layer0_outputs(2001) <= not(inputs(25));
    layer0_outputs(2002) <= not(inputs(182));
    layer0_outputs(2003) <= not(inputs(72));
    layer0_outputs(2004) <= not(inputs(189)) or (inputs(16));
    layer0_outputs(2005) <= not(inputs(210)) or (inputs(152));
    layer0_outputs(2006) <= not(inputs(84)) or (inputs(30));
    layer0_outputs(2007) <= not(inputs(193)) or (inputs(45));
    layer0_outputs(2008) <= (inputs(36)) or (inputs(191));
    layer0_outputs(2009) <= inputs(133);
    layer0_outputs(2010) <= (inputs(163)) or (inputs(19));
    layer0_outputs(2011) <= not(inputs(181));
    layer0_outputs(2012) <= (inputs(42)) and not (inputs(96));
    layer0_outputs(2013) <= (inputs(9)) and not (inputs(5));
    layer0_outputs(2014) <= not(inputs(58)) or (inputs(185));
    layer0_outputs(2015) <= not(inputs(163));
    layer0_outputs(2016) <= (inputs(191)) or (inputs(195));
    layer0_outputs(2017) <= not((inputs(54)) or (inputs(27)));
    layer0_outputs(2018) <= not(inputs(180));
    layer0_outputs(2019) <= inputs(163);
    layer0_outputs(2020) <= (inputs(150)) and not (inputs(90));
    layer0_outputs(2021) <= '0';
    layer0_outputs(2022) <= (inputs(156)) and not (inputs(223));
    layer0_outputs(2023) <= (inputs(121)) and not (inputs(234));
    layer0_outputs(2024) <= (inputs(15)) and not (inputs(64));
    layer0_outputs(2025) <= inputs(255);
    layer0_outputs(2026) <= not((inputs(19)) or (inputs(188)));
    layer0_outputs(2027) <= not(inputs(35));
    layer0_outputs(2028) <= (inputs(24)) and (inputs(90));
    layer0_outputs(2029) <= inputs(156);
    layer0_outputs(2030) <= not(inputs(117));
    layer0_outputs(2031) <= (inputs(21)) and not (inputs(211));
    layer0_outputs(2032) <= not(inputs(159)) or (inputs(140));
    layer0_outputs(2033) <= (inputs(50)) or (inputs(93));
    layer0_outputs(2034) <= not(inputs(62));
    layer0_outputs(2035) <= not((inputs(87)) or (inputs(50)));
    layer0_outputs(2036) <= not(inputs(148)) or (inputs(66));
    layer0_outputs(2037) <= not(inputs(136)) or (inputs(42));
    layer0_outputs(2038) <= not(inputs(254));
    layer0_outputs(2039) <= inputs(233);
    layer0_outputs(2040) <= (inputs(27)) and not (inputs(1));
    layer0_outputs(2041) <= (inputs(17)) or (inputs(150));
    layer0_outputs(2042) <= (inputs(155)) and not (inputs(113));
    layer0_outputs(2043) <= (inputs(147)) xor (inputs(175));
    layer0_outputs(2044) <= not(inputs(104)) or (inputs(18));
    layer0_outputs(2045) <= not(inputs(196));
    layer0_outputs(2046) <= inputs(69);
    layer0_outputs(2047) <= (inputs(193)) and not (inputs(15));
    layer0_outputs(2048) <= not(inputs(24));
    layer0_outputs(2049) <= not((inputs(9)) or (inputs(210)));
    layer0_outputs(2050) <= inputs(25);
    layer0_outputs(2051) <= not((inputs(146)) or (inputs(212)));
    layer0_outputs(2052) <= inputs(35);
    layer0_outputs(2053) <= (inputs(222)) and not (inputs(250));
    layer0_outputs(2054) <= inputs(63);
    layer0_outputs(2055) <= inputs(154);
    layer0_outputs(2056) <= (inputs(24)) or (inputs(41));
    layer0_outputs(2057) <= not(inputs(230)) or (inputs(3));
    layer0_outputs(2058) <= inputs(115);
    layer0_outputs(2059) <= not(inputs(53));
    layer0_outputs(2060) <= not((inputs(85)) or (inputs(69)));
    layer0_outputs(2061) <= (inputs(142)) or (inputs(47));
    layer0_outputs(2062) <= not((inputs(167)) xor (inputs(78)));
    layer0_outputs(2063) <= inputs(129);
    layer0_outputs(2064) <= inputs(223);
    layer0_outputs(2065) <= not(inputs(244)) or (inputs(65));
    layer0_outputs(2066) <= (inputs(97)) or (inputs(197));
    layer0_outputs(2067) <= '1';
    layer0_outputs(2068) <= inputs(247);
    layer0_outputs(2069) <= not(inputs(83));
    layer0_outputs(2070) <= not((inputs(42)) and (inputs(111)));
    layer0_outputs(2071) <= not((inputs(147)) or (inputs(14)));
    layer0_outputs(2072) <= not(inputs(8));
    layer0_outputs(2073) <= inputs(115);
    layer0_outputs(2074) <= (inputs(155)) and not (inputs(64));
    layer0_outputs(2075) <= (inputs(45)) xor (inputs(92));
    layer0_outputs(2076) <= (inputs(191)) or (inputs(157));
    layer0_outputs(2077) <= not(inputs(25));
    layer0_outputs(2078) <= (inputs(149)) and not (inputs(35));
    layer0_outputs(2079) <= not(inputs(231)) or (inputs(148));
    layer0_outputs(2080) <= (inputs(170)) or (inputs(112));
    layer0_outputs(2081) <= not(inputs(67)) or (inputs(142));
    layer0_outputs(2082) <= not(inputs(87));
    layer0_outputs(2083) <= (inputs(224)) xor (inputs(63));
    layer0_outputs(2084) <= not(inputs(253));
    layer0_outputs(2085) <= (inputs(247)) and (inputs(9));
    layer0_outputs(2086) <= inputs(97);
    layer0_outputs(2087) <= (inputs(132)) or (inputs(169));
    layer0_outputs(2088) <= (inputs(113)) and (inputs(122));
    layer0_outputs(2089) <= (inputs(87)) or (inputs(122));
    layer0_outputs(2090) <= (inputs(164)) or (inputs(68));
    layer0_outputs(2091) <= not(inputs(121));
    layer0_outputs(2092) <= not((inputs(218)) or (inputs(202)));
    layer0_outputs(2093) <= not((inputs(25)) and (inputs(124)));
    layer0_outputs(2094) <= not((inputs(174)) or (inputs(191)));
    layer0_outputs(2095) <= not((inputs(79)) or (inputs(76)));
    layer0_outputs(2096) <= not(inputs(61)) or (inputs(16));
    layer0_outputs(2097) <= (inputs(38)) or (inputs(157));
    layer0_outputs(2098) <= not((inputs(171)) or (inputs(67)));
    layer0_outputs(2099) <= (inputs(160)) or (inputs(63));
    layer0_outputs(2100) <= inputs(235);
    layer0_outputs(2101) <= not(inputs(122));
    layer0_outputs(2102) <= (inputs(33)) or (inputs(77));
    layer0_outputs(2103) <= not((inputs(183)) xor (inputs(183)));
    layer0_outputs(2104) <= (inputs(187)) and not (inputs(54));
    layer0_outputs(2105) <= '1';
    layer0_outputs(2106) <= '0';
    layer0_outputs(2107) <= not(inputs(153));
    layer0_outputs(2108) <= inputs(146);
    layer0_outputs(2109) <= (inputs(56)) and not (inputs(110));
    layer0_outputs(2110) <= (inputs(184)) and (inputs(212));
    layer0_outputs(2111) <= not(inputs(141)) or (inputs(223));
    layer0_outputs(2112) <= (inputs(99)) xor (inputs(57));
    layer0_outputs(2113) <= not(inputs(87));
    layer0_outputs(2114) <= (inputs(165)) or (inputs(77));
    layer0_outputs(2115) <= not(inputs(162));
    layer0_outputs(2116) <= not((inputs(44)) or (inputs(60)));
    layer0_outputs(2117) <= not(inputs(183)) or (inputs(101));
    layer0_outputs(2118) <= not(inputs(130));
    layer0_outputs(2119) <= not(inputs(75));
    layer0_outputs(2120) <= (inputs(8)) or (inputs(96));
    layer0_outputs(2121) <= (inputs(124)) or (inputs(7));
    layer0_outputs(2122) <= not(inputs(120));
    layer0_outputs(2123) <= (inputs(200)) or (inputs(169));
    layer0_outputs(2124) <= inputs(67);
    layer0_outputs(2125) <= (inputs(251)) and not (inputs(5));
    layer0_outputs(2126) <= not(inputs(27)) or (inputs(142));
    layer0_outputs(2127) <= (inputs(194)) and not (inputs(171));
    layer0_outputs(2128) <= (inputs(170)) or (inputs(100));
    layer0_outputs(2129) <= inputs(153);
    layer0_outputs(2130) <= not((inputs(84)) xor (inputs(0)));
    layer0_outputs(2131) <= (inputs(198)) or (inputs(30));
    layer0_outputs(2132) <= not(inputs(46));
    layer0_outputs(2133) <= inputs(169);
    layer0_outputs(2134) <= not(inputs(87));
    layer0_outputs(2135) <= (inputs(221)) or (inputs(154));
    layer0_outputs(2136) <= (inputs(13)) or (inputs(165));
    layer0_outputs(2137) <= inputs(193);
    layer0_outputs(2138) <= not(inputs(207));
    layer0_outputs(2139) <= (inputs(52)) or (inputs(123));
    layer0_outputs(2140) <= (inputs(213)) and not (inputs(27));
    layer0_outputs(2141) <= not(inputs(192));
    layer0_outputs(2142) <= not(inputs(50));
    layer0_outputs(2143) <= inputs(108);
    layer0_outputs(2144) <= inputs(99);
    layer0_outputs(2145) <= not(inputs(116)) or (inputs(4));
    layer0_outputs(2146) <= not((inputs(21)) or (inputs(82)));
    layer0_outputs(2147) <= not(inputs(164));
    layer0_outputs(2148) <= (inputs(116)) and not (inputs(230));
    layer0_outputs(2149) <= '1';
    layer0_outputs(2150) <= (inputs(162)) or (inputs(206));
    layer0_outputs(2151) <= not(inputs(73)) or (inputs(82));
    layer0_outputs(2152) <= not(inputs(198));
    layer0_outputs(2153) <= not(inputs(201));
    layer0_outputs(2154) <= not(inputs(253)) or (inputs(222));
    layer0_outputs(2155) <= not((inputs(31)) or (inputs(213)));
    layer0_outputs(2156) <= (inputs(68)) and (inputs(9));
    layer0_outputs(2157) <= not(inputs(45));
    layer0_outputs(2158) <= (inputs(217)) and (inputs(203));
    layer0_outputs(2159) <= (inputs(92)) or (inputs(218));
    layer0_outputs(2160) <= not((inputs(48)) or (inputs(11)));
    layer0_outputs(2161) <= not((inputs(84)) or (inputs(49)));
    layer0_outputs(2162) <= '1';
    layer0_outputs(2163) <= not(inputs(128));
    layer0_outputs(2164) <= inputs(231);
    layer0_outputs(2165) <= not(inputs(134));
    layer0_outputs(2166) <= (inputs(118)) or (inputs(37));
    layer0_outputs(2167) <= inputs(13);
    layer0_outputs(2168) <= not(inputs(77)) or (inputs(1));
    layer0_outputs(2169) <= not((inputs(98)) or (inputs(117)));
    layer0_outputs(2170) <= (inputs(103)) or (inputs(45));
    layer0_outputs(2171) <= not(inputs(145));
    layer0_outputs(2172) <= not((inputs(26)) or (inputs(56)));
    layer0_outputs(2173) <= inputs(168);
    layer0_outputs(2174) <= (inputs(22)) or (inputs(35));
    layer0_outputs(2175) <= inputs(27);
    layer0_outputs(2176) <= inputs(103);
    layer0_outputs(2177) <= (inputs(0)) and not (inputs(82));
    layer0_outputs(2178) <= (inputs(97)) and not (inputs(92));
    layer0_outputs(2179) <= inputs(43);
    layer0_outputs(2180) <= not((inputs(170)) xor (inputs(137)));
    layer0_outputs(2181) <= not((inputs(239)) or (inputs(149)));
    layer0_outputs(2182) <= not(inputs(207));
    layer0_outputs(2183) <= not(inputs(248)) or (inputs(161));
    layer0_outputs(2184) <= (inputs(201)) and (inputs(132));
    layer0_outputs(2185) <= not((inputs(111)) or (inputs(187)));
    layer0_outputs(2186) <= not(inputs(198)) or (inputs(101));
    layer0_outputs(2187) <= inputs(28);
    layer0_outputs(2188) <= not((inputs(152)) or (inputs(135)));
    layer0_outputs(2189) <= (inputs(188)) or (inputs(63));
    layer0_outputs(2190) <= (inputs(224)) xor (inputs(24));
    layer0_outputs(2191) <= (inputs(226)) or (inputs(56));
    layer0_outputs(2192) <= not(inputs(76));
    layer0_outputs(2193) <= not((inputs(220)) or (inputs(212)));
    layer0_outputs(2194) <= (inputs(171)) and not (inputs(248));
    layer0_outputs(2195) <= not(inputs(248));
    layer0_outputs(2196) <= not(inputs(167));
    layer0_outputs(2197) <= '1';
    layer0_outputs(2198) <= inputs(109);
    layer0_outputs(2199) <= not(inputs(8));
    layer0_outputs(2200) <= inputs(2);
    layer0_outputs(2201) <= not(inputs(115));
    layer0_outputs(2202) <= '0';
    layer0_outputs(2203) <= not(inputs(252));
    layer0_outputs(2204) <= '0';
    layer0_outputs(2205) <= (inputs(20)) xor (inputs(53));
    layer0_outputs(2206) <= '0';
    layer0_outputs(2207) <= (inputs(116)) or (inputs(222));
    layer0_outputs(2208) <= (inputs(140)) and not (inputs(252));
    layer0_outputs(2209) <= (inputs(227)) and not (inputs(158));
    layer0_outputs(2210) <= not(inputs(52));
    layer0_outputs(2211) <= not((inputs(34)) or (inputs(51)));
    layer0_outputs(2212) <= not((inputs(0)) xor (inputs(95)));
    layer0_outputs(2213) <= not((inputs(4)) or (inputs(188)));
    layer0_outputs(2214) <= not((inputs(118)) or (inputs(177)));
    layer0_outputs(2215) <= not(inputs(75)) or (inputs(13));
    layer0_outputs(2216) <= not((inputs(61)) or (inputs(133)));
    layer0_outputs(2217) <= inputs(153);
    layer0_outputs(2218) <= (inputs(251)) and not (inputs(246));
    layer0_outputs(2219) <= not(inputs(184));
    layer0_outputs(2220) <= (inputs(169)) or (inputs(113));
    layer0_outputs(2221) <= not((inputs(112)) or (inputs(102)));
    layer0_outputs(2222) <= (inputs(68)) and not (inputs(219));
    layer0_outputs(2223) <= inputs(154);
    layer0_outputs(2224) <= not((inputs(67)) or (inputs(61)));
    layer0_outputs(2225) <= (inputs(193)) or (inputs(67));
    layer0_outputs(2226) <= not(inputs(229));
    layer0_outputs(2227) <= not(inputs(169)) or (inputs(84));
    layer0_outputs(2228) <= (inputs(92)) or (inputs(97));
    layer0_outputs(2229) <= not((inputs(234)) xor (inputs(147)));
    layer0_outputs(2230) <= not((inputs(77)) or (inputs(179)));
    layer0_outputs(2231) <= (inputs(90)) and not (inputs(128));
    layer0_outputs(2232) <= inputs(145);
    layer0_outputs(2233) <= inputs(124);
    layer0_outputs(2234) <= (inputs(96)) or (inputs(34));
    layer0_outputs(2235) <= not((inputs(45)) or (inputs(65)));
    layer0_outputs(2236) <= inputs(75);
    layer0_outputs(2237) <= (inputs(104)) and not (inputs(129));
    layer0_outputs(2238) <= inputs(119);
    layer0_outputs(2239) <= inputs(202);
    layer0_outputs(2240) <= not(inputs(105));
    layer0_outputs(2241) <= (inputs(146)) or (inputs(11));
    layer0_outputs(2242) <= (inputs(23)) and not (inputs(71));
    layer0_outputs(2243) <= not(inputs(120));
    layer0_outputs(2244) <= (inputs(126)) or (inputs(216));
    layer0_outputs(2245) <= inputs(120);
    layer0_outputs(2246) <= inputs(164);
    layer0_outputs(2247) <= not(inputs(72));
    layer0_outputs(2248) <= not((inputs(211)) or (inputs(230)));
    layer0_outputs(2249) <= not(inputs(148));
    layer0_outputs(2250) <= not(inputs(217)) or (inputs(1));
    layer0_outputs(2251) <= '1';
    layer0_outputs(2252) <= not((inputs(237)) or (inputs(111)));
    layer0_outputs(2253) <= not((inputs(128)) or (inputs(245)));
    layer0_outputs(2254) <= inputs(100);
    layer0_outputs(2255) <= inputs(129);
    layer0_outputs(2256) <= inputs(231);
    layer0_outputs(2257) <= (inputs(76)) and not (inputs(160));
    layer0_outputs(2258) <= not((inputs(162)) or (inputs(203)));
    layer0_outputs(2259) <= inputs(116);
    layer0_outputs(2260) <= not((inputs(50)) or (inputs(20)));
    layer0_outputs(2261) <= inputs(225);
    layer0_outputs(2262) <= (inputs(44)) or (inputs(228));
    layer0_outputs(2263) <= not(inputs(135));
    layer0_outputs(2264) <= inputs(202);
    layer0_outputs(2265) <= inputs(80);
    layer0_outputs(2266) <= not(inputs(59));
    layer0_outputs(2267) <= (inputs(145)) or (inputs(94));
    layer0_outputs(2268) <= inputs(194);
    layer0_outputs(2269) <= not((inputs(246)) xor (inputs(104)));
    layer0_outputs(2270) <= not(inputs(83)) or (inputs(208));
    layer0_outputs(2271) <= inputs(197);
    layer0_outputs(2272) <= '1';
    layer0_outputs(2273) <= (inputs(104)) and (inputs(216));
    layer0_outputs(2274) <= (inputs(111)) or (inputs(224));
    layer0_outputs(2275) <= not((inputs(169)) or (inputs(143)));
    layer0_outputs(2276) <= (inputs(124)) and not (inputs(245));
    layer0_outputs(2277) <= not(inputs(210));
    layer0_outputs(2278) <= not(inputs(194));
    layer0_outputs(2279) <= '0';
    layer0_outputs(2280) <= (inputs(252)) and not (inputs(104));
    layer0_outputs(2281) <= not(inputs(164));
    layer0_outputs(2282) <= (inputs(209)) and not (inputs(130));
    layer0_outputs(2283) <= not(inputs(26)) or (inputs(166));
    layer0_outputs(2284) <= inputs(227);
    layer0_outputs(2285) <= not(inputs(249)) or (inputs(74));
    layer0_outputs(2286) <= not((inputs(155)) or (inputs(190)));
    layer0_outputs(2287) <= not((inputs(81)) or (inputs(195)));
    layer0_outputs(2288) <= not(inputs(141));
    layer0_outputs(2289) <= inputs(146);
    layer0_outputs(2290) <= not((inputs(234)) xor (inputs(186)));
    layer0_outputs(2291) <= (inputs(66)) xor (inputs(149));
    layer0_outputs(2292) <= not(inputs(25)) or (inputs(171));
    layer0_outputs(2293) <= not(inputs(74)) or (inputs(33));
    layer0_outputs(2294) <= not(inputs(111));
    layer0_outputs(2295) <= not((inputs(234)) xor (inputs(101)));
    layer0_outputs(2296) <= inputs(61);
    layer0_outputs(2297) <= not(inputs(149)) or (inputs(193));
    layer0_outputs(2298) <= (inputs(214)) or (inputs(71));
    layer0_outputs(2299) <= inputs(68);
    layer0_outputs(2300) <= (inputs(32)) or (inputs(30));
    layer0_outputs(2301) <= not(inputs(228)) or (inputs(9));
    layer0_outputs(2302) <= not(inputs(130)) or (inputs(211));
    layer0_outputs(2303) <= (inputs(141)) or (inputs(196));
    layer0_outputs(2304) <= not((inputs(231)) or (inputs(161)));
    layer0_outputs(2305) <= '1';
    layer0_outputs(2306) <= inputs(117);
    layer0_outputs(2307) <= not((inputs(108)) xor (inputs(3)));
    layer0_outputs(2308) <= inputs(74);
    layer0_outputs(2309) <= not(inputs(86));
    layer0_outputs(2310) <= not((inputs(145)) or (inputs(60)));
    layer0_outputs(2311) <= not(inputs(173)) or (inputs(65));
    layer0_outputs(2312) <= (inputs(247)) or (inputs(201));
    layer0_outputs(2313) <= '0';
    layer0_outputs(2314) <= inputs(228);
    layer0_outputs(2315) <= not(inputs(178)) or (inputs(95));
    layer0_outputs(2316) <= (inputs(8)) and (inputs(0));
    layer0_outputs(2317) <= not(inputs(74)) or (inputs(146));
    layer0_outputs(2318) <= not(inputs(170));
    layer0_outputs(2319) <= not(inputs(59));
    layer0_outputs(2320) <= (inputs(134)) and not (inputs(86));
    layer0_outputs(2321) <= not((inputs(200)) and (inputs(249)));
    layer0_outputs(2322) <= not((inputs(81)) or (inputs(147)));
    layer0_outputs(2323) <= not((inputs(158)) or (inputs(59)));
    layer0_outputs(2324) <= (inputs(206)) and not (inputs(175));
    layer0_outputs(2325) <= not((inputs(75)) or (inputs(48)));
    layer0_outputs(2326) <= (inputs(249)) and not (inputs(255));
    layer0_outputs(2327) <= inputs(136);
    layer0_outputs(2328) <= not((inputs(177)) xor (inputs(23)));
    layer0_outputs(2329) <= (inputs(149)) and not (inputs(49));
    layer0_outputs(2330) <= not(inputs(229));
    layer0_outputs(2331) <= not(inputs(173)) or (inputs(154));
    layer0_outputs(2332) <= not(inputs(105)) or (inputs(144));
    layer0_outputs(2333) <= not(inputs(73));
    layer0_outputs(2334) <= (inputs(247)) and not (inputs(49));
    layer0_outputs(2335) <= not(inputs(23)) or (inputs(71));
    layer0_outputs(2336) <= (inputs(254)) or (inputs(155));
    layer0_outputs(2337) <= (inputs(118)) and not (inputs(52));
    layer0_outputs(2338) <= not(inputs(100));
    layer0_outputs(2339) <= not(inputs(196));
    layer0_outputs(2340) <= (inputs(56)) and not (inputs(127));
    layer0_outputs(2341) <= inputs(248);
    layer0_outputs(2342) <= not((inputs(18)) or (inputs(64)));
    layer0_outputs(2343) <= not(inputs(150));
    layer0_outputs(2344) <= (inputs(107)) and (inputs(79));
    layer0_outputs(2345) <= inputs(168);
    layer0_outputs(2346) <= not(inputs(35));
    layer0_outputs(2347) <= not(inputs(192));
    layer0_outputs(2348) <= not((inputs(36)) or (inputs(14)));
    layer0_outputs(2349) <= not(inputs(246)) or (inputs(4));
    layer0_outputs(2350) <= (inputs(73)) or (inputs(214));
    layer0_outputs(2351) <= (inputs(165)) and (inputs(248));
    layer0_outputs(2352) <= (inputs(137)) and not (inputs(31));
    layer0_outputs(2353) <= not(inputs(229));
    layer0_outputs(2354) <= inputs(184);
    layer0_outputs(2355) <= not((inputs(83)) or (inputs(103)));
    layer0_outputs(2356) <= '0';
    layer0_outputs(2357) <= not(inputs(89));
    layer0_outputs(2358) <= (inputs(235)) or (inputs(104));
    layer0_outputs(2359) <= not((inputs(217)) or (inputs(34)));
    layer0_outputs(2360) <= not(inputs(88));
    layer0_outputs(2361) <= (inputs(75)) or (inputs(144));
    layer0_outputs(2362) <= not(inputs(172)) or (inputs(166));
    layer0_outputs(2363) <= not(inputs(119)) or (inputs(143));
    layer0_outputs(2364) <= not((inputs(123)) xor (inputs(142)));
    layer0_outputs(2365) <= (inputs(51)) and not (inputs(114));
    layer0_outputs(2366) <= (inputs(66)) xor (inputs(68));
    layer0_outputs(2367) <= (inputs(21)) or (inputs(77));
    layer0_outputs(2368) <= (inputs(32)) or (inputs(39));
    layer0_outputs(2369) <= not(inputs(90));
    layer0_outputs(2370) <= not((inputs(172)) xor (inputs(125)));
    layer0_outputs(2371) <= not(inputs(91));
    layer0_outputs(2372) <= inputs(108);
    layer0_outputs(2373) <= (inputs(193)) or (inputs(106));
    layer0_outputs(2374) <= (inputs(39)) and (inputs(134));
    layer0_outputs(2375) <= not(inputs(83)) or (inputs(138));
    layer0_outputs(2376) <= not(inputs(63)) or (inputs(33));
    layer0_outputs(2377) <= inputs(57);
    layer0_outputs(2378) <= not(inputs(14));
    layer0_outputs(2379) <= not(inputs(177));
    layer0_outputs(2380) <= not(inputs(177));
    layer0_outputs(2381) <= (inputs(58)) and not (inputs(215));
    layer0_outputs(2382) <= (inputs(199)) or (inputs(144));
    layer0_outputs(2383) <= inputs(156);
    layer0_outputs(2384) <= inputs(102);
    layer0_outputs(2385) <= (inputs(158)) or (inputs(141));
    layer0_outputs(2386) <= inputs(109);
    layer0_outputs(2387) <= not((inputs(208)) or (inputs(172)));
    layer0_outputs(2388) <= not((inputs(193)) or (inputs(178)));
    layer0_outputs(2389) <= not(inputs(242)) or (inputs(173));
    layer0_outputs(2390) <= inputs(214);
    layer0_outputs(2391) <= not(inputs(91));
    layer0_outputs(2392) <= inputs(24);
    layer0_outputs(2393) <= not(inputs(23));
    layer0_outputs(2394) <= not(inputs(33)) or (inputs(81));
    layer0_outputs(2395) <= inputs(211);
    layer0_outputs(2396) <= not((inputs(251)) and (inputs(206)));
    layer0_outputs(2397) <= (inputs(207)) or (inputs(47));
    layer0_outputs(2398) <= not(inputs(60));
    layer0_outputs(2399) <= (inputs(207)) or (inputs(194));
    layer0_outputs(2400) <= inputs(53);
    layer0_outputs(2401) <= not(inputs(147));
    layer0_outputs(2402) <= not(inputs(81)) or (inputs(250));
    layer0_outputs(2403) <= not((inputs(35)) or (inputs(38)));
    layer0_outputs(2404) <= not(inputs(251));
    layer0_outputs(2405) <= (inputs(238)) or (inputs(182));
    layer0_outputs(2406) <= (inputs(137)) and not (inputs(72));
    layer0_outputs(2407) <= not(inputs(103));
    layer0_outputs(2408) <= inputs(199);
    layer0_outputs(2409) <= not(inputs(28));
    layer0_outputs(2410) <= inputs(61);
    layer0_outputs(2411) <= '0';
    layer0_outputs(2412) <= inputs(245);
    layer0_outputs(2413) <= (inputs(28)) and not (inputs(191));
    layer0_outputs(2414) <= (inputs(18)) and (inputs(96));
    layer0_outputs(2415) <= (inputs(14)) or (inputs(242));
    layer0_outputs(2416) <= (inputs(44)) and not (inputs(238));
    layer0_outputs(2417) <= not(inputs(147));
    layer0_outputs(2418) <= inputs(137);
    layer0_outputs(2419) <= not((inputs(37)) or (inputs(135)));
    layer0_outputs(2420) <= (inputs(181)) or (inputs(208));
    layer0_outputs(2421) <= inputs(167);
    layer0_outputs(2422) <= (inputs(143)) and not (inputs(229));
    layer0_outputs(2423) <= (inputs(89)) and not (inputs(17));
    layer0_outputs(2424) <= not((inputs(27)) or (inputs(50)));
    layer0_outputs(2425) <= not(inputs(41)) or (inputs(200));
    layer0_outputs(2426) <= inputs(198);
    layer0_outputs(2427) <= (inputs(185)) xor (inputs(236));
    layer0_outputs(2428) <= not(inputs(149));
    layer0_outputs(2429) <= not(inputs(232));
    layer0_outputs(2430) <= (inputs(164)) or (inputs(236));
    layer0_outputs(2431) <= (inputs(38)) or (inputs(106));
    layer0_outputs(2432) <= not(inputs(193));
    layer0_outputs(2433) <= not(inputs(72));
    layer0_outputs(2434) <= not((inputs(9)) or (inputs(137)));
    layer0_outputs(2435) <= (inputs(139)) or (inputs(191));
    layer0_outputs(2436) <= not(inputs(40));
    layer0_outputs(2437) <= (inputs(226)) or (inputs(64));
    layer0_outputs(2438) <= not((inputs(169)) or (inputs(94)));
    layer0_outputs(2439) <= not(inputs(126));
    layer0_outputs(2440) <= not((inputs(48)) or (inputs(197)));
    layer0_outputs(2441) <= not((inputs(116)) or (inputs(255)));
    layer0_outputs(2442) <= (inputs(224)) or (inputs(3));
    layer0_outputs(2443) <= not(inputs(167));
    layer0_outputs(2444) <= (inputs(67)) or (inputs(66));
    layer0_outputs(2445) <= (inputs(170)) or (inputs(81));
    layer0_outputs(2446) <= not((inputs(93)) or (inputs(163)));
    layer0_outputs(2447) <= (inputs(60)) and (inputs(233));
    layer0_outputs(2448) <= inputs(120);
    layer0_outputs(2449) <= (inputs(221)) or (inputs(120));
    layer0_outputs(2450) <= not((inputs(188)) or (inputs(94)));
    layer0_outputs(2451) <= (inputs(6)) and not (inputs(238));
    layer0_outputs(2452) <= not((inputs(15)) or (inputs(119)));
    layer0_outputs(2453) <= not(inputs(214));
    layer0_outputs(2454) <= not((inputs(233)) or (inputs(202)));
    layer0_outputs(2455) <= (inputs(131)) and not (inputs(232));
    layer0_outputs(2456) <= not((inputs(153)) and (inputs(155)));
    layer0_outputs(2457) <= not((inputs(176)) or (inputs(181)));
    layer0_outputs(2458) <= (inputs(110)) and not (inputs(45));
    layer0_outputs(2459) <= not(inputs(104));
    layer0_outputs(2460) <= (inputs(239)) xor (inputs(210));
    layer0_outputs(2461) <= (inputs(0)) xor (inputs(227));
    layer0_outputs(2462) <= (inputs(30)) or (inputs(5));
    layer0_outputs(2463) <= not(inputs(44)) or (inputs(206));
    layer0_outputs(2464) <= inputs(189);
    layer0_outputs(2465) <= (inputs(64)) and (inputs(2));
    layer0_outputs(2466) <= (inputs(124)) or (inputs(53));
    layer0_outputs(2467) <= inputs(113);
    layer0_outputs(2468) <= not(inputs(186));
    layer0_outputs(2469) <= not((inputs(160)) or (inputs(140)));
    layer0_outputs(2470) <= not(inputs(135));
    layer0_outputs(2471) <= not((inputs(22)) or (inputs(123)));
    layer0_outputs(2472) <= not((inputs(153)) and (inputs(213)));
    layer0_outputs(2473) <= not((inputs(57)) and (inputs(101)));
    layer0_outputs(2474) <= not((inputs(78)) or (inputs(66)));
    layer0_outputs(2475) <= (inputs(44)) xor (inputs(57));
    layer0_outputs(2476) <= not(inputs(195));
    layer0_outputs(2477) <= not(inputs(170));
    layer0_outputs(2478) <= (inputs(249)) and not (inputs(11));
    layer0_outputs(2479) <= not(inputs(122));
    layer0_outputs(2480) <= not(inputs(108));
    layer0_outputs(2481) <= inputs(31);
    layer0_outputs(2482) <= not(inputs(37)) or (inputs(206));
    layer0_outputs(2483) <= not(inputs(100));
    layer0_outputs(2484) <= inputs(230);
    layer0_outputs(2485) <= (inputs(225)) or (inputs(239));
    layer0_outputs(2486) <= not(inputs(219));
    layer0_outputs(2487) <= inputs(231);
    layer0_outputs(2488) <= not((inputs(182)) and (inputs(186)));
    layer0_outputs(2489) <= '0';
    layer0_outputs(2490) <= (inputs(85)) or (inputs(233));
    layer0_outputs(2491) <= (inputs(117)) and not (inputs(238));
    layer0_outputs(2492) <= (inputs(65)) xor (inputs(17));
    layer0_outputs(2493) <= not(inputs(105));
    layer0_outputs(2494) <= not(inputs(205));
    layer0_outputs(2495) <= not(inputs(216));
    layer0_outputs(2496) <= not((inputs(67)) or (inputs(204)));
    layer0_outputs(2497) <= not(inputs(147)) or (inputs(129));
    layer0_outputs(2498) <= not(inputs(91));
    layer0_outputs(2499) <= not((inputs(255)) or (inputs(242)));
    layer0_outputs(2500) <= not((inputs(102)) or (inputs(144)));
    layer0_outputs(2501) <= '1';
    layer0_outputs(2502) <= inputs(152);
    layer0_outputs(2503) <= '1';
    layer0_outputs(2504) <= not((inputs(165)) or (inputs(81)));
    layer0_outputs(2505) <= not((inputs(66)) or (inputs(149)));
    layer0_outputs(2506) <= not(inputs(208));
    layer0_outputs(2507) <= not((inputs(254)) xor (inputs(85)));
    layer0_outputs(2508) <= inputs(135);
    layer0_outputs(2509) <= (inputs(91)) or (inputs(108));
    layer0_outputs(2510) <= (inputs(254)) or (inputs(84));
    layer0_outputs(2511) <= not((inputs(166)) or (inputs(73)));
    layer0_outputs(2512) <= inputs(144);
    layer0_outputs(2513) <= inputs(214);
    layer0_outputs(2514) <= not((inputs(253)) xor (inputs(251)));
    layer0_outputs(2515) <= inputs(211);
    layer0_outputs(2516) <= (inputs(90)) and not (inputs(233));
    layer0_outputs(2517) <= not((inputs(85)) or (inputs(79)));
    layer0_outputs(2518) <= not(inputs(237));
    layer0_outputs(2519) <= (inputs(227)) and not (inputs(82));
    layer0_outputs(2520) <= not(inputs(160)) or (inputs(1));
    layer0_outputs(2521) <= not(inputs(173));
    layer0_outputs(2522) <= not((inputs(224)) or (inputs(64)));
    layer0_outputs(2523) <= (inputs(33)) or (inputs(61));
    layer0_outputs(2524) <= inputs(243);
    layer0_outputs(2525) <= not((inputs(113)) xor (inputs(148)));
    layer0_outputs(2526) <= not((inputs(115)) or (inputs(158)));
    layer0_outputs(2527) <= (inputs(3)) or (inputs(12));
    layer0_outputs(2528) <= not(inputs(21));
    layer0_outputs(2529) <= not(inputs(227));
    layer0_outputs(2530) <= inputs(148);
    layer0_outputs(2531) <= inputs(186);
    layer0_outputs(2532) <= inputs(42);
    layer0_outputs(2533) <= not(inputs(177));
    layer0_outputs(2534) <= not(inputs(54)) or (inputs(1));
    layer0_outputs(2535) <= not(inputs(16));
    layer0_outputs(2536) <= (inputs(133)) and not (inputs(129));
    layer0_outputs(2537) <= '0';
    layer0_outputs(2538) <= not(inputs(241));
    layer0_outputs(2539) <= not(inputs(97));
    layer0_outputs(2540) <= (inputs(71)) or (inputs(242));
    layer0_outputs(2541) <= not(inputs(228)) or (inputs(112));
    layer0_outputs(2542) <= inputs(196);
    layer0_outputs(2543) <= inputs(255);
    layer0_outputs(2544) <= (inputs(26)) and not (inputs(226));
    layer0_outputs(2545) <= not(inputs(92));
    layer0_outputs(2546) <= (inputs(227)) or (inputs(139));
    layer0_outputs(2547) <= not(inputs(85));
    layer0_outputs(2548) <= not((inputs(33)) and (inputs(35)));
    layer0_outputs(2549) <= not(inputs(100));
    layer0_outputs(2550) <= not(inputs(188)) or (inputs(46));
    layer0_outputs(2551) <= inputs(209);
    layer0_outputs(2552) <= not(inputs(83)) or (inputs(140));
    layer0_outputs(2553) <= inputs(150);
    layer0_outputs(2554) <= not(inputs(76));
    layer0_outputs(2555) <= (inputs(56)) or (inputs(83));
    layer0_outputs(2556) <= (inputs(164)) and not (inputs(15));
    layer0_outputs(2557) <= '1';
    layer0_outputs(2558) <= inputs(210);
    layer0_outputs(2559) <= (inputs(109)) or (inputs(126));
    outputs(0) <= not(layer0_outputs(2173)) or (layer0_outputs(917));
    outputs(1) <= not(layer0_outputs(1865));
    outputs(2) <= layer0_outputs(354);
    outputs(3) <= layer0_outputs(1494);
    outputs(4) <= not(layer0_outputs(595)) or (layer0_outputs(1430));
    outputs(5) <= (layer0_outputs(229)) and not (layer0_outputs(373));
    outputs(6) <= layer0_outputs(794);
    outputs(7) <= (layer0_outputs(441)) or (layer0_outputs(2356));
    outputs(8) <= (layer0_outputs(1764)) and not (layer0_outputs(2516));
    outputs(9) <= (layer0_outputs(1632)) and (layer0_outputs(764));
    outputs(10) <= not(layer0_outputs(1522));
    outputs(11) <= not((layer0_outputs(1842)) and (layer0_outputs(1381)));
    outputs(12) <= layer0_outputs(583);
    outputs(13) <= layer0_outputs(854);
    outputs(14) <= (layer0_outputs(1805)) and (layer0_outputs(1420));
    outputs(15) <= layer0_outputs(1799);
    outputs(16) <= not((layer0_outputs(756)) xor (layer0_outputs(400)));
    outputs(17) <= not(layer0_outputs(215)) or (layer0_outputs(83));
    outputs(18) <= layer0_outputs(83);
    outputs(19) <= not(layer0_outputs(941));
    outputs(20) <= (layer0_outputs(501)) and not (layer0_outputs(2344));
    outputs(21) <= layer0_outputs(1136);
    outputs(22) <= not((layer0_outputs(1613)) xor (layer0_outputs(2429)));
    outputs(23) <= not(layer0_outputs(1257)) or (layer0_outputs(1964));
    outputs(24) <= (layer0_outputs(1033)) and not (layer0_outputs(542));
    outputs(25) <= not(layer0_outputs(2129));
    outputs(26) <= layer0_outputs(1270);
    outputs(27) <= layer0_outputs(145);
    outputs(28) <= layer0_outputs(2263);
    outputs(29) <= not(layer0_outputs(257));
    outputs(30) <= layer0_outputs(1425);
    outputs(31) <= not(layer0_outputs(1491));
    outputs(32) <= not(layer0_outputs(1698));
    outputs(33) <= not(layer0_outputs(581));
    outputs(34) <= (layer0_outputs(1898)) and (layer0_outputs(1456));
    outputs(35) <= (layer0_outputs(907)) and not (layer0_outputs(1324));
    outputs(36) <= (layer0_outputs(2188)) and (layer0_outputs(587));
    outputs(37) <= not(layer0_outputs(2245));
    outputs(38) <= (layer0_outputs(1885)) and not (layer0_outputs(2125));
    outputs(39) <= not(layer0_outputs(402));
    outputs(40) <= not(layer0_outputs(1478));
    outputs(41) <= not(layer0_outputs(1609)) or (layer0_outputs(2334));
    outputs(42) <= not((layer0_outputs(1866)) or (layer0_outputs(984)));
    outputs(43) <= layer0_outputs(1451);
    outputs(44) <= layer0_outputs(1643);
    outputs(45) <= not(layer0_outputs(2258));
    outputs(46) <= not(layer0_outputs(2323));
    outputs(47) <= not(layer0_outputs(206));
    outputs(48) <= not(layer0_outputs(1207));
    outputs(49) <= layer0_outputs(981);
    outputs(50) <= not((layer0_outputs(2473)) and (layer0_outputs(410)));
    outputs(51) <= (layer0_outputs(1750)) xor (layer0_outputs(1846));
    outputs(52) <= not((layer0_outputs(1085)) or (layer0_outputs(1554)));
    outputs(53) <= not(layer0_outputs(2288));
    outputs(54) <= not(layer0_outputs(2171));
    outputs(55) <= not(layer0_outputs(1769)) or (layer0_outputs(2296));
    outputs(56) <= layer0_outputs(600);
    outputs(57) <= not(layer0_outputs(1584));
    outputs(58) <= not(layer0_outputs(277));
    outputs(59) <= layer0_outputs(977);
    outputs(60) <= layer0_outputs(175);
    outputs(61) <= (layer0_outputs(1409)) and not (layer0_outputs(1662));
    outputs(62) <= not(layer0_outputs(1261));
    outputs(63) <= not(layer0_outputs(450));
    outputs(64) <= (layer0_outputs(1887)) and not (layer0_outputs(982));
    outputs(65) <= layer0_outputs(2386);
    outputs(66) <= not((layer0_outputs(2483)) or (layer0_outputs(1101)));
    outputs(67) <= not(layer0_outputs(1972)) or (layer0_outputs(930));
    outputs(68) <= layer0_outputs(983);
    outputs(69) <= layer0_outputs(793);
    outputs(70) <= not(layer0_outputs(50)) or (layer0_outputs(2208));
    outputs(71) <= not(layer0_outputs(1634)) or (layer0_outputs(980));
    outputs(72) <= layer0_outputs(1756);
    outputs(73) <= (layer0_outputs(1000)) or (layer0_outputs(260));
    outputs(74) <= not(layer0_outputs(2462));
    outputs(75) <= (layer0_outputs(2037)) and not (layer0_outputs(1407));
    outputs(76) <= not((layer0_outputs(648)) and (layer0_outputs(1496)));
    outputs(77) <= (layer0_outputs(1889)) and not (layer0_outputs(1999));
    outputs(78) <= layer0_outputs(2479);
    outputs(79) <= layer0_outputs(1488);
    outputs(80) <= not(layer0_outputs(850));
    outputs(81) <= not(layer0_outputs(2330)) or (layer0_outputs(1236));
    outputs(82) <= not(layer0_outputs(2418));
    outputs(83) <= not(layer0_outputs(1081)) or (layer0_outputs(146));
    outputs(84) <= (layer0_outputs(119)) and (layer0_outputs(29));
    outputs(85) <= (layer0_outputs(1614)) and (layer0_outputs(1425));
    outputs(86) <= (layer0_outputs(1353)) or (layer0_outputs(1390));
    outputs(87) <= not(layer0_outputs(532));
    outputs(88) <= not((layer0_outputs(1350)) xor (layer0_outputs(348)));
    outputs(89) <= (layer0_outputs(2555)) and not (layer0_outputs(236));
    outputs(90) <= layer0_outputs(2047);
    outputs(91) <= (layer0_outputs(1037)) and not (layer0_outputs(278));
    outputs(92) <= layer0_outputs(1189);
    outputs(93) <= not((layer0_outputs(1568)) or (layer0_outputs(1779)));
    outputs(94) <= not(layer0_outputs(1831));
    outputs(95) <= not(layer0_outputs(1070)) or (layer0_outputs(1801));
    outputs(96) <= not(layer0_outputs(456));
    outputs(97) <= (layer0_outputs(549)) and not (layer0_outputs(841));
    outputs(98) <= (layer0_outputs(1910)) and not (layer0_outputs(318));
    outputs(99) <= layer0_outputs(1403);
    outputs(100) <= not(layer0_outputs(381));
    outputs(101) <= not(layer0_outputs(867));
    outputs(102) <= not((layer0_outputs(1251)) and (layer0_outputs(2005)));
    outputs(103) <= (layer0_outputs(957)) and not (layer0_outputs(2421));
    outputs(104) <= layer0_outputs(1436);
    outputs(105) <= (layer0_outputs(2443)) and (layer0_outputs(1940));
    outputs(106) <= (layer0_outputs(363)) and not (layer0_outputs(1522));
    outputs(107) <= not(layer0_outputs(982));
    outputs(108) <= (layer0_outputs(1305)) or (layer0_outputs(577));
    outputs(109) <= layer0_outputs(1036);
    outputs(110) <= not((layer0_outputs(681)) or (layer0_outputs(716)));
    outputs(111) <= not(layer0_outputs(748)) or (layer0_outputs(1502));
    outputs(112) <= layer0_outputs(1248);
    outputs(113) <= (layer0_outputs(2107)) and (layer0_outputs(885));
    outputs(114) <= layer0_outputs(847);
    outputs(115) <= (layer0_outputs(2419)) or (layer0_outputs(927));
    outputs(116) <= not(layer0_outputs(986));
    outputs(117) <= (layer0_outputs(639)) and not (layer0_outputs(2133));
    outputs(118) <= not(layer0_outputs(683));
    outputs(119) <= not(layer0_outputs(2095));
    outputs(120) <= not(layer0_outputs(2322)) or (layer0_outputs(1933));
    outputs(121) <= layer0_outputs(2264);
    outputs(122) <= not(layer0_outputs(1977));
    outputs(123) <= layer0_outputs(488);
    outputs(124) <= not(layer0_outputs(1814));
    outputs(125) <= layer0_outputs(1876);
    outputs(126) <= not(layer0_outputs(1315));
    outputs(127) <= layer0_outputs(2289);
    outputs(128) <= not(layer0_outputs(1872));
    outputs(129) <= layer0_outputs(1291);
    outputs(130) <= not(layer0_outputs(1370));
    outputs(131) <= not(layer0_outputs(1117)) or (layer0_outputs(110));
    outputs(132) <= not(layer0_outputs(105));
    outputs(133) <= (layer0_outputs(1264)) or (layer0_outputs(1265));
    outputs(134) <= not(layer0_outputs(2131));
    outputs(135) <= not(layer0_outputs(2295));
    outputs(136) <= not((layer0_outputs(467)) or (layer0_outputs(1252)));
    outputs(137) <= not(layer0_outputs(658));
    outputs(138) <= not((layer0_outputs(651)) and (layer0_outputs(979)));
    outputs(139) <= (layer0_outputs(2165)) and not (layer0_outputs(386));
    outputs(140) <= (layer0_outputs(94)) and not (layer0_outputs(2215));
    outputs(141) <= (layer0_outputs(1364)) and not (layer0_outputs(899));
    outputs(142) <= (layer0_outputs(1394)) xor (layer0_outputs(407));
    outputs(143) <= layer0_outputs(1938);
    outputs(144) <= layer0_outputs(221);
    outputs(145) <= (layer0_outputs(2044)) and not (layer0_outputs(2405));
    outputs(146) <= (layer0_outputs(1905)) or (layer0_outputs(2400));
    outputs(147) <= layer0_outputs(423);
    outputs(148) <= layer0_outputs(160);
    outputs(149) <= (layer0_outputs(894)) and not (layer0_outputs(1779));
    outputs(150) <= (layer0_outputs(12)) or (layer0_outputs(691));
    outputs(151) <= not(layer0_outputs(1286));
    outputs(152) <= layer0_outputs(1626);
    outputs(153) <= layer0_outputs(2372);
    outputs(154) <= (layer0_outputs(55)) and not (layer0_outputs(1604));
    outputs(155) <= not(layer0_outputs(631));
    outputs(156) <= not(layer0_outputs(733));
    outputs(157) <= (layer0_outputs(317)) and (layer0_outputs(2164));
    outputs(158) <= layer0_outputs(1702);
    outputs(159) <= not(layer0_outputs(1421));
    outputs(160) <= (layer0_outputs(1270)) and not (layer0_outputs(1674));
    outputs(161) <= not(layer0_outputs(2533));
    outputs(162) <= (layer0_outputs(1552)) and not (layer0_outputs(2098));
    outputs(163) <= not((layer0_outputs(2294)) or (layer0_outputs(2435)));
    outputs(164) <= not((layer0_outputs(1963)) or (layer0_outputs(2324)));
    outputs(165) <= (layer0_outputs(343)) and not (layer0_outputs(2057));
    outputs(166) <= layer0_outputs(1503);
    outputs(167) <= not((layer0_outputs(270)) and (layer0_outputs(1003)));
    outputs(168) <= not(layer0_outputs(1465));
    outputs(169) <= layer0_outputs(1782);
    outputs(170) <= layer0_outputs(1601);
    outputs(171) <= not(layer0_outputs(2337)) or (layer0_outputs(2026));
    outputs(172) <= layer0_outputs(1800);
    outputs(173) <= not((layer0_outputs(1130)) xor (layer0_outputs(1376)));
    outputs(174) <= (layer0_outputs(1713)) and (layer0_outputs(1989));
    outputs(175) <= layer0_outputs(892);
    outputs(176) <= not((layer0_outputs(93)) or (layer0_outputs(2331)));
    outputs(177) <= not((layer0_outputs(2287)) and (layer0_outputs(1715)));
    outputs(178) <= layer0_outputs(1746);
    outputs(179) <= not((layer0_outputs(1201)) and (layer0_outputs(874)));
    outputs(180) <= not(layer0_outputs(1316));
    outputs(181) <= (layer0_outputs(1924)) and not (layer0_outputs(2217));
    outputs(182) <= layer0_outputs(1037);
    outputs(183) <= (layer0_outputs(1423)) and not (layer0_outputs(1669));
    outputs(184) <= not(layer0_outputs(2401));
    outputs(185) <= not(layer0_outputs(599));
    outputs(186) <= layer0_outputs(742);
    outputs(187) <= not(layer0_outputs(1438)) or (layer0_outputs(1142));
    outputs(188) <= not((layer0_outputs(1797)) or (layer0_outputs(848)));
    outputs(189) <= not(layer0_outputs(581));
    outputs(190) <= not((layer0_outputs(590)) or (layer0_outputs(797)));
    outputs(191) <= not((layer0_outputs(245)) or (layer0_outputs(473)));
    outputs(192) <= (layer0_outputs(693)) or (layer0_outputs(529));
    outputs(193) <= not(layer0_outputs(2503)) or (layer0_outputs(1913));
    outputs(194) <= not(layer0_outputs(1449)) or (layer0_outputs(290));
    outputs(195) <= not(layer0_outputs(1820));
    outputs(196) <= (layer0_outputs(1760)) xor (layer0_outputs(1358));
    outputs(197) <= (layer0_outputs(2522)) and (layer0_outputs(85));
    outputs(198) <= layer0_outputs(1039);
    outputs(199) <= layer0_outputs(118);
    outputs(200) <= not(layer0_outputs(1182));
    outputs(201) <= not((layer0_outputs(992)) xor (layer0_outputs(1979)));
    outputs(202) <= not(layer0_outputs(1232)) or (layer0_outputs(17));
    outputs(203) <= not((layer0_outputs(2017)) or (layer0_outputs(2320)));
    outputs(204) <= layer0_outputs(420);
    outputs(205) <= not(layer0_outputs(1823)) or (layer0_outputs(2086));
    outputs(206) <= not(layer0_outputs(815));
    outputs(207) <= not(layer0_outputs(707));
    outputs(208) <= not(layer0_outputs(147));
    outputs(209) <= not(layer0_outputs(960));
    outputs(210) <= (layer0_outputs(426)) and (layer0_outputs(2184));
    outputs(211) <= not(layer0_outputs(391));
    outputs(212) <= layer0_outputs(754);
    outputs(213) <= layer0_outputs(2395);
    outputs(214) <= not(layer0_outputs(1584));
    outputs(215) <= layer0_outputs(1012);
    outputs(216) <= not((layer0_outputs(815)) or (layer0_outputs(2100)));
    outputs(217) <= not((layer0_outputs(382)) and (layer0_outputs(193)));
    outputs(218) <= not(layer0_outputs(1826));
    outputs(219) <= not(layer0_outputs(1600));
    outputs(220) <= not(layer0_outputs(1052)) or (layer0_outputs(1464));
    outputs(221) <= not(layer0_outputs(2495));
    outputs(222) <= not((layer0_outputs(946)) or (layer0_outputs(1815)));
    outputs(223) <= (layer0_outputs(1813)) and not (layer0_outputs(2290));
    outputs(224) <= not(layer0_outputs(4));
    outputs(225) <= not(layer0_outputs(453)) or (layer0_outputs(1164));
    outputs(226) <= (layer0_outputs(425)) and not (layer0_outputs(82));
    outputs(227) <= not(layer0_outputs(338));
    outputs(228) <= not(layer0_outputs(1891)) or (layer0_outputs(506));
    outputs(229) <= layer0_outputs(86);
    outputs(230) <= (layer0_outputs(1768)) and (layer0_outputs(916));
    outputs(231) <= (layer0_outputs(1481)) and not (layer0_outputs(1816));
    outputs(232) <= layer0_outputs(2377);
    outputs(233) <= layer0_outputs(413);
    outputs(234) <= layer0_outputs(1188);
    outputs(235) <= not(layer0_outputs(558)) or (layer0_outputs(41));
    outputs(236) <= not(layer0_outputs(1735));
    outputs(237) <= not(layer0_outputs(138));
    outputs(238) <= (layer0_outputs(2179)) and not (layer0_outputs(373));
    outputs(239) <= not(layer0_outputs(450));
    outputs(240) <= layer0_outputs(2410);
    outputs(241) <= not(layer0_outputs(2253)) or (layer0_outputs(641));
    outputs(242) <= layer0_outputs(321);
    outputs(243) <= layer0_outputs(1836);
    outputs(244) <= not(layer0_outputs(2278));
    outputs(245) <= not(layer0_outputs(670));
    outputs(246) <= (layer0_outputs(948)) and not (layer0_outputs(252));
    outputs(247) <= not((layer0_outputs(2448)) or (layer0_outputs(1717)));
    outputs(248) <= (layer0_outputs(80)) and not (layer0_outputs(1369));
    outputs(249) <= not(layer0_outputs(1497));
    outputs(250) <= not(layer0_outputs(835)) or (layer0_outputs(895));
    outputs(251) <= not(layer0_outputs(1687)) or (layer0_outputs(1642));
    outputs(252) <= (layer0_outputs(1382)) or (layer0_outputs(676));
    outputs(253) <= not(layer0_outputs(2238));
    outputs(254) <= (layer0_outputs(584)) or (layer0_outputs(2137));
    outputs(255) <= not((layer0_outputs(59)) or (layer0_outputs(1381)));
    outputs(256) <= (layer0_outputs(5)) and not (layer0_outputs(1261));
    outputs(257) <= (layer0_outputs(2213)) and not (layer0_outputs(1895));
    outputs(258) <= (layer0_outputs(559)) and not (layer0_outputs(350));
    outputs(259) <= layer0_outputs(2338);
    outputs(260) <= not((layer0_outputs(2064)) or (layer0_outputs(190)));
    outputs(261) <= not((layer0_outputs(243)) or (layer0_outputs(1913)));
    outputs(262) <= (layer0_outputs(570)) and not (layer0_outputs(351));
    outputs(263) <= (layer0_outputs(1102)) and (layer0_outputs(1215));
    outputs(264) <= not(layer0_outputs(1660));
    outputs(265) <= (layer0_outputs(1516)) and (layer0_outputs(1169));
    outputs(266) <= (layer0_outputs(655)) and not (layer0_outputs(2134));
    outputs(267) <= not(layer0_outputs(647));
    outputs(268) <= (layer0_outputs(366)) and not (layer0_outputs(857));
    outputs(269) <= (layer0_outputs(872)) and (layer0_outputs(1644));
    outputs(270) <= (layer0_outputs(1587)) and (layer0_outputs(1373));
    outputs(271) <= (layer0_outputs(251)) and not (layer0_outputs(1096));
    outputs(272) <= not((layer0_outputs(1043)) or (layer0_outputs(92)));
    outputs(273) <= not(layer0_outputs(1960));
    outputs(274) <= layer0_outputs(283);
    outputs(275) <= not((layer0_outputs(542)) or (layer0_outputs(1695)));
    outputs(276) <= layer0_outputs(2048);
    outputs(277) <= (layer0_outputs(1546)) and (layer0_outputs(47));
    outputs(278) <= (layer0_outputs(99)) and not (layer0_outputs(1357));
    outputs(279) <= (layer0_outputs(780)) and (layer0_outputs(2498));
    outputs(280) <= (layer0_outputs(1940)) and (layer0_outputs(1434));
    outputs(281) <= (layer0_outputs(1285)) and (layer0_outputs(2502));
    outputs(282) <= (layer0_outputs(730)) and (layer0_outputs(1715));
    outputs(283) <= (layer0_outputs(2401)) and not (layer0_outputs(1096));
    outputs(284) <= (layer0_outputs(514)) and not (layer0_outputs(237));
    outputs(285) <= (layer0_outputs(746)) and (layer0_outputs(1359));
    outputs(286) <= not((layer0_outputs(2128)) or (layer0_outputs(1293)));
    outputs(287) <= not((layer0_outputs(124)) or (layer0_outputs(2336)));
    outputs(288) <= not(layer0_outputs(922));
    outputs(289) <= (layer0_outputs(1166)) and not (layer0_outputs(118));
    outputs(290) <= not((layer0_outputs(1304)) or (layer0_outputs(1015)));
    outputs(291) <= (layer0_outputs(1219)) and (layer0_outputs(1199));
    outputs(292) <= not((layer0_outputs(993)) or (layer0_outputs(592)));
    outputs(293) <= (layer0_outputs(1968)) and (layer0_outputs(1072));
    outputs(294) <= not(layer0_outputs(75));
    outputs(295) <= not(layer0_outputs(2241));
    outputs(296) <= (layer0_outputs(194)) and not (layer0_outputs(551));
    outputs(297) <= (layer0_outputs(1943)) and not (layer0_outputs(1434));
    outputs(298) <= (layer0_outputs(971)) and not (layer0_outputs(2460));
    outputs(299) <= (layer0_outputs(2260)) and (layer0_outputs(2176));
    outputs(300) <= layer0_outputs(1932);
    outputs(301) <= (layer0_outputs(12)) and (layer0_outputs(327));
    outputs(302) <= (layer0_outputs(468)) and (layer0_outputs(1095));
    outputs(303) <= (layer0_outputs(554)) and not (layer0_outputs(1351));
    outputs(304) <= (layer0_outputs(1610)) and (layer0_outputs(2185));
    outputs(305) <= layer0_outputs(1808);
    outputs(306) <= (layer0_outputs(1654)) and (layer0_outputs(1841));
    outputs(307) <= layer0_outputs(168);
    outputs(308) <= (layer0_outputs(197)) and not (layer0_outputs(1080));
    outputs(309) <= (layer0_outputs(2324)) and not (layer0_outputs(1232));
    outputs(310) <= (layer0_outputs(1280)) and (layer0_outputs(1666));
    outputs(311) <= '0';
    outputs(312) <= (layer0_outputs(43)) and (layer0_outputs(1202));
    outputs(313) <= not((layer0_outputs(1131)) or (layer0_outputs(2225)));
    outputs(314) <= (layer0_outputs(1617)) and (layer0_outputs(1758));
    outputs(315) <= (layer0_outputs(940)) and not (layer0_outputs(383));
    outputs(316) <= (layer0_outputs(1624)) and not (layer0_outputs(1312));
    outputs(317) <= '0';
    outputs(318) <= '0';
    outputs(319) <= (layer0_outputs(1189)) and not (layer0_outputs(121));
    outputs(320) <= (layer0_outputs(734)) and (layer0_outputs(555));
    outputs(321) <= (layer0_outputs(602)) and not (layer0_outputs(1451));
    outputs(322) <= not((layer0_outputs(804)) or (layer0_outputs(227)));
    outputs(323) <= (layer0_outputs(2438)) and (layer0_outputs(155));
    outputs(324) <= not((layer0_outputs(1683)) or (layer0_outputs(2159)));
    outputs(325) <= not((layer0_outputs(2242)) or (layer0_outputs(1589)));
    outputs(326) <= (layer0_outputs(1629)) and (layer0_outputs(1894));
    outputs(327) <= (layer0_outputs(1755)) and not (layer0_outputs(1236));
    outputs(328) <= (layer0_outputs(1592)) and not (layer0_outputs(2267));
    outputs(329) <= (layer0_outputs(603)) and not (layer0_outputs(441));
    outputs(330) <= not((layer0_outputs(339)) or (layer0_outputs(615)));
    outputs(331) <= not((layer0_outputs(1063)) or (layer0_outputs(2440)));
    outputs(332) <= not((layer0_outputs(358)) or (layer0_outputs(2268)));
    outputs(333) <= (layer0_outputs(1822)) and not (layer0_outputs(1625));
    outputs(334) <= not(layer0_outputs(1026));
    outputs(335) <= (layer0_outputs(898)) and not (layer0_outputs(1019));
    outputs(336) <= not((layer0_outputs(1927)) or (layer0_outputs(364)));
    outputs(337) <= not((layer0_outputs(129)) xor (layer0_outputs(904)));
    outputs(338) <= not((layer0_outputs(1281)) or (layer0_outputs(2128)));
    outputs(339) <= not(layer0_outputs(762));
    outputs(340) <= (layer0_outputs(448)) and not (layer0_outputs(1379));
    outputs(341) <= (layer0_outputs(2214)) and (layer0_outputs(2472));
    outputs(342) <= (layer0_outputs(1416)) and not (layer0_outputs(1518));
    outputs(343) <= (layer0_outputs(55)) and (layer0_outputs(1640));
    outputs(344) <= (layer0_outputs(45)) and (layer0_outputs(2252));
    outputs(345) <= not((layer0_outputs(1317)) or (layer0_outputs(232)));
    outputs(346) <= not((layer0_outputs(2063)) or (layer0_outputs(653)));
    outputs(347) <= (layer0_outputs(2542)) and (layer0_outputs(2023));
    outputs(348) <= (layer0_outputs(457)) and not (layer0_outputs(1329));
    outputs(349) <= (layer0_outputs(812)) and (layer0_outputs(749));
    outputs(350) <= not((layer0_outputs(694)) or (layer0_outputs(1178)));
    outputs(351) <= (layer0_outputs(250)) and (layer0_outputs(655));
    outputs(352) <= (layer0_outputs(1154)) and not (layer0_outputs(1157));
    outputs(353) <= (layer0_outputs(229)) and not (layer0_outputs(2102));
    outputs(354) <= (layer0_outputs(1956)) and not (layer0_outputs(2256));
    outputs(355) <= not((layer0_outputs(2546)) or (layer0_outputs(1721)));
    outputs(356) <= not((layer0_outputs(2200)) or (layer0_outputs(529)));
    outputs(357) <= (layer0_outputs(1729)) and (layer0_outputs(241));
    outputs(358) <= (layer0_outputs(1730)) and not (layer0_outputs(72));
    outputs(359) <= (layer0_outputs(512)) and not (layer0_outputs(2240));
    outputs(360) <= not((layer0_outputs(1456)) or (layer0_outputs(2445)));
    outputs(361) <= (layer0_outputs(1785)) and (layer0_outputs(1263));
    outputs(362) <= not(layer0_outputs(389));
    outputs(363) <= not((layer0_outputs(260)) or (layer0_outputs(2285)));
    outputs(364) <= (layer0_outputs(1762)) and not (layer0_outputs(1751));
    outputs(365) <= (layer0_outputs(1682)) and not (layer0_outputs(668));
    outputs(366) <= layer0_outputs(1633);
    outputs(367) <= (layer0_outputs(1652)) and (layer0_outputs(1579));
    outputs(368) <= (layer0_outputs(1520)) and (layer0_outputs(219));
    outputs(369) <= not((layer0_outputs(562)) or (layer0_outputs(61)));
    outputs(370) <= not((layer0_outputs(2259)) or (layer0_outputs(2257)));
    outputs(371) <= (layer0_outputs(1439)) and not (layer0_outputs(2466));
    outputs(372) <= (layer0_outputs(1432)) and not (layer0_outputs(2462));
    outputs(373) <= (layer0_outputs(788)) and not (layer0_outputs(1597));
    outputs(374) <= not((layer0_outputs(2114)) or (layer0_outputs(2174)));
    outputs(375) <= (layer0_outputs(1709)) and (layer0_outputs(2539));
    outputs(376) <= (layer0_outputs(750)) and not (layer0_outputs(2016));
    outputs(377) <= (layer0_outputs(1501)) and not (layer0_outputs(2285));
    outputs(378) <= not((layer0_outputs(1835)) or (layer0_outputs(2075)));
    outputs(379) <= not((layer0_outputs(654)) or (layer0_outputs(2220)));
    outputs(380) <= (layer0_outputs(317)) and (layer0_outputs(1847));
    outputs(381) <= (layer0_outputs(2229)) and not (layer0_outputs(1702));
    outputs(382) <= (layer0_outputs(1644)) and not (layer0_outputs(27));
    outputs(383) <= not((layer0_outputs(434)) or (layer0_outputs(1899)));
    outputs(384) <= not((layer0_outputs(1179)) or (layer0_outputs(150)));
    outputs(385) <= (layer0_outputs(990)) and (layer0_outputs(2353));
    outputs(386) <= layer0_outputs(151);
    outputs(387) <= (layer0_outputs(1570)) and not (layer0_outputs(2220));
    outputs(388) <= (layer0_outputs(1169)) and not (layer0_outputs(1031));
    outputs(389) <= not(layer0_outputs(2159));
    outputs(390) <= (layer0_outputs(0)) and (layer0_outputs(153));
    outputs(391) <= '0';
    outputs(392) <= (layer0_outputs(302)) and not (layer0_outputs(1185));
    outputs(393) <= (layer0_outputs(1163)) and not (layer0_outputs(463));
    outputs(394) <= (layer0_outputs(1595)) and not (layer0_outputs(1980));
    outputs(395) <= (layer0_outputs(112)) and (layer0_outputs(2169));
    outputs(396) <= (layer0_outputs(1288)) and not (layer0_outputs(586));
    outputs(397) <= (layer0_outputs(1221)) and not (layer0_outputs(1440));
    outputs(398) <= (layer0_outputs(2138)) and not (layer0_outputs(2523));
    outputs(399) <= (layer0_outputs(679)) and not (layer0_outputs(1404));
    outputs(400) <= (layer0_outputs(1959)) and (layer0_outputs(617));
    outputs(401) <= (layer0_outputs(1570)) and not (layer0_outputs(2373));
    outputs(402) <= (layer0_outputs(1144)) and not (layer0_outputs(1836));
    outputs(403) <= (layer0_outputs(680)) and (layer0_outputs(25));
    outputs(404) <= (layer0_outputs(875)) and not (layer0_outputs(1470));
    outputs(405) <= not(layer0_outputs(26));
    outputs(406) <= not((layer0_outputs(885)) or (layer0_outputs(2120)));
    outputs(407) <= (layer0_outputs(1580)) and not (layer0_outputs(2300));
    outputs(408) <= (layer0_outputs(1884)) and not (layer0_outputs(2255));
    outputs(409) <= (layer0_outputs(2315)) and not (layer0_outputs(980));
    outputs(410) <= not((layer0_outputs(1837)) or (layer0_outputs(790)));
    outputs(411) <= not(layer0_outputs(909));
    outputs(412) <= not((layer0_outputs(836)) or (layer0_outputs(1969)));
    outputs(413) <= (layer0_outputs(2525)) and (layer0_outputs(1513));
    outputs(414) <= (layer0_outputs(1458)) and not (layer0_outputs(1812));
    outputs(415) <= layer0_outputs(2471);
    outputs(416) <= not((layer0_outputs(1574)) or (layer0_outputs(1625)));
    outputs(417) <= (layer0_outputs(193)) and (layer0_outputs(1146));
    outputs(418) <= (layer0_outputs(1044)) and (layer0_outputs(781));
    outputs(419) <= (layer0_outputs(733)) and (layer0_outputs(1040));
    outputs(420) <= (layer0_outputs(76)) and not (layer0_outputs(1021));
    outputs(421) <= not((layer0_outputs(1331)) or (layer0_outputs(149)));
    outputs(422) <= not((layer0_outputs(1791)) or (layer0_outputs(961)));
    outputs(423) <= not((layer0_outputs(471)) or (layer0_outputs(927)));
    outputs(424) <= not(layer0_outputs(2470));
    outputs(425) <= (layer0_outputs(814)) and (layer0_outputs(2353));
    outputs(426) <= (layer0_outputs(265)) and not (layer0_outputs(1909));
    outputs(427) <= (layer0_outputs(1687)) and not (layer0_outputs(544));
    outputs(428) <= (layer0_outputs(1148)) and not (layer0_outputs(674));
    outputs(429) <= (layer0_outputs(414)) and (layer0_outputs(2359));
    outputs(430) <= (layer0_outputs(959)) and (layer0_outputs(39));
    outputs(431) <= not((layer0_outputs(1293)) or (layer0_outputs(2087)));
    outputs(432) <= not((layer0_outputs(1922)) or (layer0_outputs(1627)));
    outputs(433) <= (layer0_outputs(633)) and not (layer0_outputs(747));
    outputs(434) <= (layer0_outputs(521)) xor (layer0_outputs(802));
    outputs(435) <= (layer0_outputs(652)) and not (layer0_outputs(501));
    outputs(436) <= (layer0_outputs(547)) and not (layer0_outputs(2076));
    outputs(437) <= layer0_outputs(2146);
    outputs(438) <= (layer0_outputs(642)) and not (layer0_outputs(136));
    outputs(439) <= not((layer0_outputs(1567)) or (layer0_outputs(1544)));
    outputs(440) <= layer0_outputs(1095);
    outputs(441) <= (layer0_outputs(1268)) and not (layer0_outputs(1132));
    outputs(442) <= not((layer0_outputs(1849)) or (layer0_outputs(517)));
    outputs(443) <= (layer0_outputs(1951)) and not (layer0_outputs(177));
    outputs(444) <= not((layer0_outputs(127)) xor (layer0_outputs(1231)));
    outputs(445) <= (layer0_outputs(1149)) and not (layer0_outputs(2256));
    outputs(446) <= layer0_outputs(1176);
    outputs(447) <= (layer0_outputs(960)) and (layer0_outputs(194));
    outputs(448) <= not(layer0_outputs(1347));
    outputs(449) <= layer0_outputs(999);
    outputs(450) <= (layer0_outputs(530)) and (layer0_outputs(1561));
    outputs(451) <= not((layer0_outputs(2110)) or (layer0_outputs(2166)));
    outputs(452) <= '0';
    outputs(453) <= (layer0_outputs(1852)) and not (layer0_outputs(37));
    outputs(454) <= layer0_outputs(1555);
    outputs(455) <= (layer0_outputs(1875)) and (layer0_outputs(65));
    outputs(456) <= (layer0_outputs(732)) and not (layer0_outputs(117));
    outputs(457) <= (layer0_outputs(316)) and not (layer0_outputs(1379));
    outputs(458) <= not(layer0_outputs(2299));
    outputs(459) <= not((layer0_outputs(2433)) or (layer0_outputs(411)));
    outputs(460) <= layer0_outputs(1263);
    outputs(461) <= not((layer0_outputs(2028)) or (layer0_outputs(933)));
    outputs(462) <= not((layer0_outputs(606)) or (layer0_outputs(1267)));
    outputs(463) <= (layer0_outputs(1737)) and (layer0_outputs(2506));
    outputs(464) <= (layer0_outputs(1778)) and not (layer0_outputs(1745));
    outputs(465) <= (layer0_outputs(1220)) and not (layer0_outputs(1242));
    outputs(466) <= layer0_outputs(1061);
    outputs(467) <= (layer0_outputs(73)) and (layer0_outputs(1530));
    outputs(468) <= (layer0_outputs(1118)) and (layer0_outputs(1768));
    outputs(469) <= (layer0_outputs(1283)) and (layer0_outputs(792));
    outputs(470) <= (layer0_outputs(2514)) and not (layer0_outputs(1770));
    outputs(471) <= (layer0_outputs(852)) and not (layer0_outputs(880));
    outputs(472) <= (layer0_outputs(724)) and not (layer0_outputs(49));
    outputs(473) <= (layer0_outputs(1447)) and (layer0_outputs(1749));
    outputs(474) <= (layer0_outputs(1841)) and not (layer0_outputs(1335));
    outputs(475) <= (layer0_outputs(2404)) and not (layer0_outputs(2435));
    outputs(476) <= (layer0_outputs(2340)) and (layer0_outputs(2287));
    outputs(477) <= not((layer0_outputs(566)) xor (layer0_outputs(1336)));
    outputs(478) <= (layer0_outputs(1790)) and not (layer0_outputs(22));
    outputs(479) <= (layer0_outputs(1341)) and not (layer0_outputs(727));
    outputs(480) <= not((layer0_outputs(447)) or (layer0_outputs(2470)));
    outputs(481) <= (layer0_outputs(2488)) and (layer0_outputs(955));
    outputs(482) <= (layer0_outputs(2216)) and not (layer0_outputs(2073));
    outputs(483) <= (layer0_outputs(536)) and not (layer0_outputs(1023));
    outputs(484) <= not((layer0_outputs(66)) or (layer0_outputs(403)));
    outputs(485) <= (layer0_outputs(1590)) and not (layer0_outputs(2262));
    outputs(486) <= (layer0_outputs(761)) and not (layer0_outputs(1651));
    outputs(487) <= not((layer0_outputs(2076)) or (layer0_outputs(2139)));
    outputs(488) <= layer0_outputs(1113);
    outputs(489) <= not(layer0_outputs(691));
    outputs(490) <= (layer0_outputs(1868)) and (layer0_outputs(1859));
    outputs(491) <= not((layer0_outputs(1512)) or (layer0_outputs(339)));
    outputs(492) <= (layer0_outputs(4)) and (layer0_outputs(2051));
    outputs(493) <= (layer0_outputs(165)) and (layer0_outputs(1208));
    outputs(494) <= (layer0_outputs(1718)) and not (layer0_outputs(409));
    outputs(495) <= not((layer0_outputs(225)) or (layer0_outputs(2117)));
    outputs(496) <= not((layer0_outputs(1063)) or (layer0_outputs(933)));
    outputs(497) <= (layer0_outputs(1646)) and (layer0_outputs(1342));
    outputs(498) <= (layer0_outputs(286)) and not (layer0_outputs(1601));
    outputs(499) <= (layer0_outputs(378)) and not (layer0_outputs(2218));
    outputs(500) <= (layer0_outputs(1439)) and not (layer0_outputs(329));
    outputs(501) <= not((layer0_outputs(2135)) or (layer0_outputs(1367)));
    outputs(502) <= (layer0_outputs(1859)) and (layer0_outputs(2258));
    outputs(503) <= not((layer0_outputs(2052)) or (layer0_outputs(1925)));
    outputs(504) <= layer0_outputs(812);
    outputs(505) <= (layer0_outputs(1211)) and not (layer0_outputs(67));
    outputs(506) <= (layer0_outputs(1241)) and not (layer0_outputs(2267));
    outputs(507) <= not((layer0_outputs(2427)) or (layer0_outputs(437)));
    outputs(508) <= (layer0_outputs(477)) and (layer0_outputs(1866));
    outputs(509) <= (layer0_outputs(2095)) and not (layer0_outputs(2097));
    outputs(510) <= (layer0_outputs(2155)) and not (layer0_outputs(1361));
    outputs(511) <= (layer0_outputs(2370)) and (layer0_outputs(1279));
    outputs(512) <= not(layer0_outputs(1917));
    outputs(513) <= layer0_outputs(1075);
    outputs(514) <= (layer0_outputs(2136)) or (layer0_outputs(180));
    outputs(515) <= not(layer0_outputs(1983));
    outputs(516) <= layer0_outputs(25);
    outputs(517) <= layer0_outputs(2271);
    outputs(518) <= (layer0_outputs(314)) and not (layer0_outputs(541));
    outputs(519) <= layer0_outputs(604);
    outputs(520) <= layer0_outputs(98);
    outputs(521) <= not(layer0_outputs(1667));
    outputs(522) <= (layer0_outputs(561)) and (layer0_outputs(834));
    outputs(523) <= layer0_outputs(505);
    outputs(524) <= not(layer0_outputs(341));
    outputs(525) <= not(layer0_outputs(742));
    outputs(526) <= (layer0_outputs(390)) xor (layer0_outputs(1561));
    outputs(527) <= (layer0_outputs(366)) and (layer0_outputs(1698));
    outputs(528) <= layer0_outputs(1298);
    outputs(529) <= not(layer0_outputs(49)) or (layer0_outputs(97));
    outputs(530) <= not(layer0_outputs(357)) or (layer0_outputs(768));
    outputs(531) <= not(layer0_outputs(699));
    outputs(532) <= (layer0_outputs(2531)) or (layer0_outputs(284));
    outputs(533) <= layer0_outputs(1333);
    outputs(534) <= (layer0_outputs(1783)) and (layer0_outputs(1378));
    outputs(535) <= layer0_outputs(2201);
    outputs(536) <= not(layer0_outputs(1838));
    outputs(537) <= not(layer0_outputs(440)) or (layer0_outputs(1484));
    outputs(538) <= layer0_outputs(865);
    outputs(539) <= not(layer0_outputs(377));
    outputs(540) <= not(layer0_outputs(1821));
    outputs(541) <= not((layer0_outputs(2144)) or (layer0_outputs(368)));
    outputs(542) <= not(layer0_outputs(342)) or (layer0_outputs(472));
    outputs(543) <= (layer0_outputs(912)) and not (layer0_outputs(1562));
    outputs(544) <= not((layer0_outputs(2020)) xor (layer0_outputs(1114)));
    outputs(545) <= (layer0_outputs(1385)) xor (layer0_outputs(1812));
    outputs(546) <= not(layer0_outputs(2342)) or (layer0_outputs(208));
    outputs(547) <= not(layer0_outputs(1937));
    outputs(548) <= not(layer0_outputs(2318));
    outputs(549) <= layer0_outputs(2221);
    outputs(550) <= layer0_outputs(2355);
    outputs(551) <= layer0_outputs(2270);
    outputs(552) <= not(layer0_outputs(1786));
    outputs(553) <= not((layer0_outputs(956)) and (layer0_outputs(177)));
    outputs(554) <= layer0_outputs(779);
    outputs(555) <= not(layer0_outputs(610));
    outputs(556) <= not(layer0_outputs(1426));
    outputs(557) <= not(layer0_outputs(864));
    outputs(558) <= not(layer0_outputs(111));
    outputs(559) <= layer0_outputs(1615);
    outputs(560) <= (layer0_outputs(1798)) or (layer0_outputs(2064));
    outputs(561) <= not(layer0_outputs(1213)) or (layer0_outputs(2157));
    outputs(562) <= not(layer0_outputs(1125));
    outputs(563) <= not(layer0_outputs(451)) or (layer0_outputs(53));
    outputs(564) <= (layer0_outputs(2370)) and (layer0_outputs(105));
    outputs(565) <= not(layer0_outputs(2468));
    outputs(566) <= (layer0_outputs(2362)) and not (layer0_outputs(2544));
    outputs(567) <= not(layer0_outputs(1321));
    outputs(568) <= layer0_outputs(701);
    outputs(569) <= layer0_outputs(2282);
    outputs(570) <= (layer0_outputs(1098)) and (layer0_outputs(380));
    outputs(571) <= (layer0_outputs(1424)) and not (layer0_outputs(637));
    outputs(572) <= not(layer0_outputs(1155)) or (layer0_outputs(1539));
    outputs(573) <= not(layer0_outputs(405));
    outputs(574) <= layer0_outputs(1538);
    outputs(575) <= (layer0_outputs(1816)) or (layer0_outputs(2096));
    outputs(576) <= layer0_outputs(2399);
    outputs(577) <= layer0_outputs(659);
    outputs(578) <= layer0_outputs(1247);
    outputs(579) <= (layer0_outputs(1004)) or (layer0_outputs(1212));
    outputs(580) <= not(layer0_outputs(2491));
    outputs(581) <= layer0_outputs(1167);
    outputs(582) <= (layer0_outputs(2056)) and not (layer0_outputs(744));
    outputs(583) <= (layer0_outputs(1153)) and not (layer0_outputs(2279));
    outputs(584) <= (layer0_outputs(1296)) or (layer0_outputs(185));
    outputs(585) <= (layer0_outputs(521)) and (layer0_outputs(1302));
    outputs(586) <= not(layer0_outputs(195));
    outputs(587) <= (layer0_outputs(630)) and (layer0_outputs(862));
    outputs(588) <= layer0_outputs(943);
    outputs(589) <= not(layer0_outputs(1636));
    outputs(590) <= (layer0_outputs(1115)) or (layer0_outputs(957));
    outputs(591) <= not(layer0_outputs(791));
    outputs(592) <= not(layer0_outputs(1726));
    outputs(593) <= layer0_outputs(1703);
    outputs(594) <= layer0_outputs(1174);
    outputs(595) <= (layer0_outputs(1399)) and (layer0_outputs(1843));
    outputs(596) <= not(layer0_outputs(161));
    outputs(597) <= layer0_outputs(1416);
    outputs(598) <= layer0_outputs(976);
    outputs(599) <= not(layer0_outputs(2254));
    outputs(600) <= (layer0_outputs(378)) and not (layer0_outputs(1708));
    outputs(601) <= not(layer0_outputs(2227));
    outputs(602) <= not(layer0_outputs(379));
    outputs(603) <= layer0_outputs(2268);
    outputs(604) <= not(layer0_outputs(1925));
    outputs(605) <= layer0_outputs(2209);
    outputs(606) <= (layer0_outputs(2469)) xor (layer0_outputs(1848));
    outputs(607) <= (layer0_outputs(85)) or (layer0_outputs(432));
    outputs(608) <= layer0_outputs(2216);
    outputs(609) <= layer0_outputs(146);
    outputs(610) <= not((layer0_outputs(1252)) or (layer0_outputs(1078)));
    outputs(611) <= (layer0_outputs(228)) and not (layer0_outputs(1119));
    outputs(612) <= not(layer0_outputs(1186));
    outputs(613) <= not(layer0_outputs(1222));
    outputs(614) <= layer0_outputs(79);
    outputs(615) <= layer0_outputs(258);
    outputs(616) <= (layer0_outputs(1819)) and not (layer0_outputs(304));
    outputs(617) <= not((layer0_outputs(1676)) and (layer0_outputs(801)));
    outputs(618) <= (layer0_outputs(1486)) and not (layer0_outputs(1079));
    outputs(619) <= (layer0_outputs(330)) or (layer0_outputs(1677));
    outputs(620) <= layer0_outputs(1647);
    outputs(621) <= not(layer0_outputs(95)) or (layer0_outputs(52));
    outputs(622) <= (layer0_outputs(1168)) and not (layer0_outputs(1361));
    outputs(623) <= not(layer0_outputs(2348)) or (layer0_outputs(2223));
    outputs(624) <= layer0_outputs(725);
    outputs(625) <= layer0_outputs(134);
    outputs(626) <= not(layer0_outputs(1152));
    outputs(627) <= layer0_outputs(493);
    outputs(628) <= not(layer0_outputs(1992));
    outputs(629) <= not((layer0_outputs(108)) xor (layer0_outputs(639)));
    outputs(630) <= (layer0_outputs(1032)) and not (layer0_outputs(368));
    outputs(631) <= not(layer0_outputs(1828));
    outputs(632) <= layer0_outputs(1161);
    outputs(633) <= not((layer0_outputs(1970)) and (layer0_outputs(840)));
    outputs(634) <= not(layer0_outputs(535));
    outputs(635) <= layer0_outputs(50);
    outputs(636) <= not((layer0_outputs(1071)) or (layer0_outputs(471)));
    outputs(637) <= not((layer0_outputs(995)) and (layer0_outputs(869)));
    outputs(638) <= layer0_outputs(1993);
    outputs(639) <= layer0_outputs(1773);
    outputs(640) <= layer0_outputs(1062);
    outputs(641) <= layer0_outputs(349);
    outputs(642) <= not(layer0_outputs(1043));
    outputs(643) <= (layer0_outputs(492)) and not (layer0_outputs(2457));
    outputs(644) <= not(layer0_outputs(293)) or (layer0_outputs(2365));
    outputs(645) <= layer0_outputs(2354);
    outputs(646) <= not(layer0_outputs(1873));
    outputs(647) <= not(layer0_outputs(2073));
    outputs(648) <= (layer0_outputs(1296)) or (layer0_outputs(2553));
    outputs(649) <= (layer0_outputs(2157)) or (layer0_outputs(2025));
    outputs(650) <= layer0_outputs(1159);
    outputs(651) <= layer0_outputs(604);
    outputs(652) <= (layer0_outputs(264)) or (layer0_outputs(1893));
    outputs(653) <= not(layer0_outputs(1537));
    outputs(654) <= not((layer0_outputs(1377)) or (layer0_outputs(1012)));
    outputs(655) <= not(layer0_outputs(360));
    outputs(656) <= (layer0_outputs(942)) and (layer0_outputs(531));
    outputs(657) <= layer0_outputs(979);
    outputs(658) <= layer0_outputs(1502);
    outputs(659) <= (layer0_outputs(595)) and (layer0_outputs(2014));
    outputs(660) <= layer0_outputs(1884);
    outputs(661) <= not(layer0_outputs(1308));
    outputs(662) <= layer0_outputs(614);
    outputs(663) <= (layer0_outputs(551)) and (layer0_outputs(1173));
    outputs(664) <= (layer0_outputs(1300)) and (layer0_outputs(1022));
    outputs(665) <= not(layer0_outputs(1883));
    outputs(666) <= not(layer0_outputs(326));
    outputs(667) <= layer0_outputs(1897);
    outputs(668) <= (layer0_outputs(1168)) and not (layer0_outputs(1888));
    outputs(669) <= layer0_outputs(87);
    outputs(670) <= not((layer0_outputs(353)) and (layer0_outputs(1950)));
    outputs(671) <= not((layer0_outputs(708)) and (layer0_outputs(2084)));
    outputs(672) <= not(layer0_outputs(2117));
    outputs(673) <= (layer0_outputs(33)) xor (layer0_outputs(147));
    outputs(674) <= not(layer0_outputs(596));
    outputs(675) <= not(layer0_outputs(1541));
    outputs(676) <= layer0_outputs(257);
    outputs(677) <= not((layer0_outputs(23)) or (layer0_outputs(2092)));
    outputs(678) <= (layer0_outputs(2483)) and not (layer0_outputs(2440));
    outputs(679) <= not((layer0_outputs(699)) or (layer0_outputs(127)));
    outputs(680) <= not((layer0_outputs(2541)) or (layer0_outputs(346)));
    outputs(681) <= not(layer0_outputs(379));
    outputs(682) <= layer0_outputs(65);
    outputs(683) <= not(layer0_outputs(392));
    outputs(684) <= not((layer0_outputs(539)) and (layer0_outputs(498)));
    outputs(685) <= not((layer0_outputs(535)) or (layer0_outputs(924)));
    outputs(686) <= (layer0_outputs(1854)) and (layer0_outputs(1569));
    outputs(687) <= (layer0_outputs(1448)) or (layer0_outputs(839));
    outputs(688) <= not(layer0_outputs(2412)) or (layer0_outputs(1074));
    outputs(689) <= layer0_outputs(509);
    outputs(690) <= layer0_outputs(417);
    outputs(691) <= (layer0_outputs(1837)) xor (layer0_outputs(156));
    outputs(692) <= (layer0_outputs(2174)) and not (layer0_outputs(2086));
    outputs(693) <= not(layer0_outputs(2229));
    outputs(694) <= (layer0_outputs(1092)) and (layer0_outputs(1269));
    outputs(695) <= not((layer0_outputs(361)) or (layer0_outputs(1875)));
    outputs(696) <= layer0_outputs(525);
    outputs(697) <= not(layer0_outputs(1619));
    outputs(698) <= layer0_outputs(1149);
    outputs(699) <= (layer0_outputs(634)) and not (layer0_outputs(1930));
    outputs(700) <= not((layer0_outputs(1813)) and (layer0_outputs(415)));
    outputs(701) <= not(layer0_outputs(422));
    outputs(702) <= (layer0_outputs(1586)) or (layer0_outputs(1328));
    outputs(703) <= not(layer0_outputs(187));
    outputs(704) <= layer0_outputs(1686);
    outputs(705) <= not((layer0_outputs(2497)) and (layer0_outputs(451)));
    outputs(706) <= layer0_outputs(1901);
    outputs(707) <= layer0_outputs(2284);
    outputs(708) <= layer0_outputs(1067);
    outputs(709) <= layer0_outputs(2515);
    outputs(710) <= not(layer0_outputs(1400));
    outputs(711) <= not(layer0_outputs(1297)) or (layer0_outputs(2083));
    outputs(712) <= layer0_outputs(467);
    outputs(713) <= not(layer0_outputs(1778));
    outputs(714) <= not(layer0_outputs(1818));
    outputs(715) <= layer0_outputs(520);
    outputs(716) <= layer0_outputs(259);
    outputs(717) <= not((layer0_outputs(1962)) or (layer0_outputs(823)));
    outputs(718) <= not((layer0_outputs(619)) or (layer0_outputs(222)));
    outputs(719) <= not(layer0_outputs(1398)) or (layer0_outputs(2398));
    outputs(720) <= not(layer0_outputs(361));
    outputs(721) <= (layer0_outputs(2263)) or (layer0_outputs(2010));
    outputs(722) <= (layer0_outputs(1672)) and (layer0_outputs(1896));
    outputs(723) <= not(layer0_outputs(2281));
    outputs(724) <= layer0_outputs(34);
    outputs(725) <= not((layer0_outputs(152)) and (layer0_outputs(875)));
    outputs(726) <= not(layer0_outputs(2007));
    outputs(727) <= not((layer0_outputs(2315)) and (layer0_outputs(1683)));
    outputs(728) <= not(layer0_outputs(1132));
    outputs(729) <= (layer0_outputs(1949)) and (layer0_outputs(215));
    outputs(730) <= (layer0_outputs(109)) xor (layer0_outputs(140));
    outputs(731) <= not(layer0_outputs(2277));
    outputs(732) <= not((layer0_outputs(2499)) and (layer0_outputs(439)));
    outputs(733) <= not(layer0_outputs(1504));
    outputs(734) <= layer0_outputs(321);
    outputs(735) <= layer0_outputs(926);
    outputs(736) <= not(layer0_outputs(1204));
    outputs(737) <= not((layer0_outputs(1510)) or (layer0_outputs(1832)));
    outputs(738) <= not(layer0_outputs(1649)) or (layer0_outputs(550));
    outputs(739) <= (layer0_outputs(2542)) and not (layer0_outputs(289));
    outputs(740) <= layer0_outputs(2114);
    outputs(741) <= not(layer0_outputs(2388)) or (layer0_outputs(1974));
    outputs(742) <= layer0_outputs(1156);
    outputs(743) <= layer0_outputs(987);
    outputs(744) <= (layer0_outputs(1961)) and not (layer0_outputs(2219));
    outputs(745) <= layer0_outputs(1803);
    outputs(746) <= not(layer0_outputs(1480)) or (layer0_outputs(2235));
    outputs(747) <= not(layer0_outputs(1354));
    outputs(748) <= not((layer0_outputs(459)) and (layer0_outputs(2307)));
    outputs(749) <= layer0_outputs(158);
    outputs(750) <= not(layer0_outputs(1556));
    outputs(751) <= not(layer0_outputs(426)) or (layer0_outputs(1990));
    outputs(752) <= (layer0_outputs(1289)) and (layer0_outputs(1731));
    outputs(753) <= not(layer0_outputs(721));
    outputs(754) <= (layer0_outputs(1202)) xor (layer0_outputs(828));
    outputs(755) <= layer0_outputs(81);
    outputs(756) <= not(layer0_outputs(1444)) or (layer0_outputs(1453));
    outputs(757) <= layer0_outputs(1824);
    outputs(758) <= layer0_outputs(2110);
    outputs(759) <= layer0_outputs(634);
    outputs(760) <= not(layer0_outputs(438));
    outputs(761) <= layer0_outputs(448);
    outputs(762) <= not(layer0_outputs(947));
    outputs(763) <= not(layer0_outputs(438));
    outputs(764) <= not(layer0_outputs(370)) or (layer0_outputs(777));
    outputs(765) <= layer0_outputs(1659);
    outputs(766) <= not(layer0_outputs(1014));
    outputs(767) <= (layer0_outputs(348)) and (layer0_outputs(1365));
    outputs(768) <= (layer0_outputs(2068)) and not (layer0_outputs(2291));
    outputs(769) <= layer0_outputs(959);
    outputs(770) <= not(layer0_outputs(2362)) or (layer0_outputs(2189));
    outputs(771) <= (layer0_outputs(330)) and not (layer0_outputs(2452));
    outputs(772) <= not(layer0_outputs(2096));
    outputs(773) <= not(layer0_outputs(2494)) or (layer0_outputs(470));
    outputs(774) <= layer0_outputs(2505);
    outputs(775) <= not(layer0_outputs(249)) or (layer0_outputs(487));
    outputs(776) <= not(layer0_outputs(233));
    outputs(777) <= (layer0_outputs(2460)) and not (layer0_outputs(1547));
    outputs(778) <= (layer0_outputs(2061)) and not (layer0_outputs(597));
    outputs(779) <= (layer0_outputs(2312)) and not (layer0_outputs(1156));
    outputs(780) <= layer0_outputs(2350);
    outputs(781) <= not(layer0_outputs(616));
    outputs(782) <= layer0_outputs(1508);
    outputs(783) <= layer0_outputs(1292);
    outputs(784) <= layer0_outputs(1557);
    outputs(785) <= layer0_outputs(216);
    outputs(786) <= not(layer0_outputs(1540));
    outputs(787) <= (layer0_outputs(136)) xor (layer0_outputs(786));
    outputs(788) <= not((layer0_outputs(2330)) or (layer0_outputs(280)));
    outputs(789) <= not(layer0_outputs(455));
    outputs(790) <= (layer0_outputs(515)) and (layer0_outputs(652));
    outputs(791) <= not(layer0_outputs(2091));
    outputs(792) <= (layer0_outputs(1902)) and not (layer0_outputs(1918));
    outputs(793) <= (layer0_outputs(1994)) or (layer0_outputs(418));
    outputs(794) <= not(layer0_outputs(81));
    outputs(795) <= (layer0_outputs(2309)) and (layer0_outputs(1067));
    outputs(796) <= (layer0_outputs(2045)) and (layer0_outputs(2238));
    outputs(797) <= not((layer0_outputs(1310)) xor (layer0_outputs(435)));
    outputs(798) <= (layer0_outputs(2312)) and not (layer0_outputs(1190));
    outputs(799) <= (layer0_outputs(251)) xor (layer0_outputs(1681));
    outputs(800) <= not(layer0_outputs(1640));
    outputs(801) <= (layer0_outputs(254)) and (layer0_outputs(1679));
    outputs(802) <= layer0_outputs(1099);
    outputs(803) <= (layer0_outputs(1124)) or (layer0_outputs(706));
    outputs(804) <= layer0_outputs(537);
    outputs(805) <= not(layer0_outputs(1455));
    outputs(806) <= not(layer0_outputs(1521));
    outputs(807) <= layer0_outputs(929);
    outputs(808) <= not(layer0_outputs(168));
    outputs(809) <= (layer0_outputs(1323)) and (layer0_outputs(2412));
    outputs(810) <= (layer0_outputs(611)) and not (layer0_outputs(2140));
    outputs(811) <= layer0_outputs(953);
    outputs(812) <= not(layer0_outputs(627));
    outputs(813) <= not(layer0_outputs(1674)) or (layer0_outputs(587));
    outputs(814) <= not((layer0_outputs(46)) or (layer0_outputs(2422)));
    outputs(815) <= (layer0_outputs(270)) and (layer0_outputs(673));
    outputs(816) <= not(layer0_outputs(69));
    outputs(817) <= not(layer0_outputs(2195));
    outputs(818) <= not((layer0_outputs(1167)) or (layer0_outputs(1830)));
    outputs(819) <= not(layer0_outputs(90));
    outputs(820) <= layer0_outputs(1303);
    outputs(821) <= layer0_outputs(167);
    outputs(822) <= (layer0_outputs(1030)) and not (layer0_outputs(1881));
    outputs(823) <= (layer0_outputs(1786)) and (layer0_outputs(392));
    outputs(824) <= not(layer0_outputs(1569));
    outputs(825) <= layer0_outputs(1732);
    outputs(826) <= layer0_outputs(830);
    outputs(827) <= not((layer0_outputs(1685)) xor (layer0_outputs(1147)));
    outputs(828) <= (layer0_outputs(1443)) and not (layer0_outputs(740));
    outputs(829) <= layer0_outputs(38);
    outputs(830) <= (layer0_outputs(2135)) and not (layer0_outputs(919));
    outputs(831) <= not(layer0_outputs(1466));
    outputs(832) <= not((layer0_outputs(724)) xor (layer0_outputs(1124)));
    outputs(833) <= (layer0_outputs(107)) and not (layer0_outputs(87));
    outputs(834) <= not((layer0_outputs(1103)) and (layer0_outputs(568)));
    outputs(835) <= not((layer0_outputs(34)) or (layer0_outputs(944)));
    outputs(836) <= (layer0_outputs(1259)) and not (layer0_outputs(1265));
    outputs(837) <= not((layer0_outputs(1083)) or (layer0_outputs(683)));
    outputs(838) <= (layer0_outputs(861)) and (layer0_outputs(795));
    outputs(839) <= not((layer0_outputs(916)) or (layer0_outputs(943)));
    outputs(840) <= (layer0_outputs(2012)) and not (layer0_outputs(837));
    outputs(841) <= not((layer0_outputs(1535)) or (layer0_outputs(452)));
    outputs(842) <= (layer0_outputs(2154)) and (layer0_outputs(115));
    outputs(843) <= (layer0_outputs(777)) and not (layer0_outputs(128));
    outputs(844) <= layer0_outputs(1066);
    outputs(845) <= not(layer0_outputs(888)) or (layer0_outputs(1053));
    outputs(846) <= (layer0_outputs(156)) and (layer0_outputs(1385));
    outputs(847) <= (layer0_outputs(433)) and not (layer0_outputs(1276));
    outputs(848) <= not(layer0_outputs(282));
    outputs(849) <= layer0_outputs(915);
    outputs(850) <= (layer0_outputs(571)) and not (layer0_outputs(2046));
    outputs(851) <= not(layer0_outputs(1213));
    outputs(852) <= layer0_outputs(2438);
    outputs(853) <= (layer0_outputs(1461)) or (layer0_outputs(1996));
    outputs(854) <= (layer0_outputs(1783)) and not (layer0_outputs(2434));
    outputs(855) <= not((layer0_outputs(2467)) or (layer0_outputs(1713)));
    outputs(856) <= layer0_outputs(1716);
    outputs(857) <= layer0_outputs(8);
    outputs(858) <= not(layer0_outputs(1998));
    outputs(859) <= (layer0_outputs(1878)) and (layer0_outputs(2358));
    outputs(860) <= layer0_outputs(1560);
    outputs(861) <= not((layer0_outputs(1283)) and (layer0_outputs(832)));
    outputs(862) <= (layer0_outputs(2089)) and not (layer0_outputs(552));
    outputs(863) <= layer0_outputs(966);
    outputs(864) <= not(layer0_outputs(884)) or (layer0_outputs(183));
    outputs(865) <= layer0_outputs(1904);
    outputs(866) <= not(layer0_outputs(2463)) or (layer0_outputs(1728));
    outputs(867) <= not((layer0_outputs(625)) xor (layer0_outputs(2317)));
    outputs(868) <= (layer0_outputs(236)) and not (layer0_outputs(1797));
    outputs(869) <= layer0_outputs(302);
    outputs(870) <= not(layer0_outputs(2079));
    outputs(871) <= not(layer0_outputs(287));
    outputs(872) <= not(layer0_outputs(2243));
    outputs(873) <= layer0_outputs(1740);
    outputs(874) <= layer0_outputs(840);
    outputs(875) <= (layer0_outputs(2392)) and not (layer0_outputs(11));
    outputs(876) <= (layer0_outputs(2121)) and not (layer0_outputs(1599));
    outputs(877) <= not(layer0_outputs(1938));
    outputs(878) <= not(layer0_outputs(1123)) or (layer0_outputs(2279));
    outputs(879) <= (layer0_outputs(817)) and (layer0_outputs(1254));
    outputs(880) <= not(layer0_outputs(197));
    outputs(881) <= (layer0_outputs(1209)) and not (layer0_outputs(2001));
    outputs(882) <= not((layer0_outputs(2478)) xor (layer0_outputs(475)));
    outputs(883) <= (layer0_outputs(2161)) or (layer0_outputs(1105));
    outputs(884) <= layer0_outputs(1719);
    outputs(885) <= not(layer0_outputs(2124));
    outputs(886) <= not(layer0_outputs(289));
    outputs(887) <= not(layer0_outputs(2151));
    outputs(888) <= not(layer0_outputs(2444));
    outputs(889) <= not(layer0_outputs(387));
    outputs(890) <= layer0_outputs(1878);
    outputs(891) <= layer0_outputs(860);
    outputs(892) <= (layer0_outputs(2404)) xor (layer0_outputs(1352));
    outputs(893) <= not((layer0_outputs(1562)) or (layer0_outputs(159)));
    outputs(894) <= not(layer0_outputs(1111));
    outputs(895) <= layer0_outputs(262);
    outputs(896) <= not((layer0_outputs(220)) or (layer0_outputs(305)));
    outputs(897) <= layer0_outputs(2337);
    outputs(898) <= (layer0_outputs(338)) and (layer0_outputs(293));
    outputs(899) <= layer0_outputs(30);
    outputs(900) <= (layer0_outputs(1609)) and not (layer0_outputs(1429));
    outputs(901) <= not(layer0_outputs(1991)) or (layer0_outputs(1088));
    outputs(902) <= not(layer0_outputs(1830));
    outputs(903) <= not(layer0_outputs(277));
    outputs(904) <= (layer0_outputs(940)) and not (layer0_outputs(592));
    outputs(905) <= (layer0_outputs(1735)) and not (layer0_outputs(1843));
    outputs(906) <= not(layer0_outputs(986));
    outputs(907) <= layer0_outputs(1109);
    outputs(908) <= layer0_outputs(1788);
    outputs(909) <= layer0_outputs(1673);
    outputs(910) <= not(layer0_outputs(416));
    outputs(911) <= (layer0_outputs(508)) and not (layer0_outputs(1446));
    outputs(912) <= not(layer0_outputs(1691));
    outputs(913) <= (layer0_outputs(398)) or (layer0_outputs(417));
    outputs(914) <= layer0_outputs(1268);
    outputs(915) <= not((layer0_outputs(949)) or (layer0_outputs(369)));
    outputs(916) <= (layer0_outputs(1346)) and (layer0_outputs(1857));
    outputs(917) <= layer0_outputs(2383);
    outputs(918) <= layer0_outputs(2230);
    outputs(919) <= (layer0_outputs(2050)) and not (layer0_outputs(1469));
    outputs(920) <= not(layer0_outputs(2101));
    outputs(921) <= layer0_outputs(2176);
    outputs(922) <= not(layer0_outputs(2311)) or (layer0_outputs(1217));
    outputs(923) <= not(layer0_outputs(1412));
    outputs(924) <= not(layer0_outputs(630));
    outputs(925) <= layer0_outputs(1235);
    outputs(926) <= layer0_outputs(1538);
    outputs(927) <= not(layer0_outputs(213)) or (layer0_outputs(1472));
    outputs(928) <= (layer0_outputs(1492)) or (layer0_outputs(2419));
    outputs(929) <= layer0_outputs(262);
    outputs(930) <= layer0_outputs(1685);
    outputs(931) <= layer0_outputs(1734);
    outputs(932) <= not(layer0_outputs(2066));
    outputs(933) <= not((layer0_outputs(1251)) xor (layer0_outputs(626)));
    outputs(934) <= not(layer0_outputs(1742));
    outputs(935) <= (layer0_outputs(2168)) xor (layer0_outputs(519));
    outputs(936) <= layer0_outputs(2504);
    outputs(937) <= layer0_outputs(937);
    outputs(938) <= (layer0_outputs(1920)) and (layer0_outputs(1182));
    outputs(939) <= layer0_outputs(1670);
    outputs(940) <= not(layer0_outputs(1386));
    outputs(941) <= layer0_outputs(950);
    outputs(942) <= (layer0_outputs(102)) and not (layer0_outputs(2178));
    outputs(943) <= not(layer0_outputs(1757));
    outputs(944) <= (layer0_outputs(1316)) and (layer0_outputs(481));
    outputs(945) <= layer0_outputs(1082);
    outputs(946) <= not((layer0_outputs(250)) or (layer0_outputs(1616)));
    outputs(947) <= not((layer0_outputs(360)) or (layer0_outputs(234)));
    outputs(948) <= (layer0_outputs(306)) or (layer0_outputs(191));
    outputs(949) <= not((layer0_outputs(91)) or (layer0_outputs(1705)));
    outputs(950) <= not((layer0_outputs(802)) xor (layer0_outputs(1139)));
    outputs(951) <= not(layer0_outputs(2521));
    outputs(952) <= not((layer0_outputs(1606)) and (layer0_outputs(2077)));
    outputs(953) <= (layer0_outputs(410)) and not (layer0_outputs(431));
    outputs(954) <= (layer0_outputs(698)) and not (layer0_outputs(208));
    outputs(955) <= (layer0_outputs(547)) and not (layer0_outputs(1604));
    outputs(956) <= not(layer0_outputs(1623)) or (layer0_outputs(371));
    outputs(957) <= layer0_outputs(2147);
    outputs(958) <= not(layer0_outputs(1427)) or (layer0_outputs(705));
    outputs(959) <= layer0_outputs(1622);
    outputs(960) <= (layer0_outputs(810)) or (layer0_outputs(1771));
    outputs(961) <= (layer0_outputs(856)) and not (layer0_outputs(778));
    outputs(962) <= not(layer0_outputs(838));
    outputs(963) <= not((layer0_outputs(1375)) or (layer0_outputs(1133)));
    outputs(964) <= layer0_outputs(1266);
    outputs(965) <= not(layer0_outputs(62));
    outputs(966) <= (layer0_outputs(1163)) and (layer0_outputs(1858));
    outputs(967) <= layer0_outputs(963);
    outputs(968) <= not(layer0_outputs(372));
    outputs(969) <= (layer0_outputs(1295)) and not (layer0_outputs(913));
    outputs(970) <= (layer0_outputs(88)) and (layer0_outputs(752));
    outputs(971) <= layer0_outputs(2170);
    outputs(972) <= not(layer0_outputs(58));
    outputs(973) <= not(layer0_outputs(1539));
    outputs(974) <= not(layer0_outputs(1789));
    outputs(975) <= not(layer0_outputs(1675));
    outputs(976) <= not(layer0_outputs(2132)) or (layer0_outputs(2042));
    outputs(977) <= not(layer0_outputs(1782));
    outputs(978) <= not(layer0_outputs(2408));
    outputs(979) <= layer0_outputs(312);
    outputs(980) <= layer0_outputs(857);
    outputs(981) <= (layer0_outputs(2071)) and (layer0_outputs(1617));
    outputs(982) <= (layer0_outputs(890)) and not (layer0_outputs(799));
    outputs(983) <= (layer0_outputs(494)) and not (layer0_outputs(2459));
    outputs(984) <= not(layer0_outputs(2434));
    outputs(985) <= not(layer0_outputs(1641));
    outputs(986) <= layer0_outputs(1699);
    outputs(987) <= (layer0_outputs(1767)) or (layer0_outputs(1367));
    outputs(988) <= not((layer0_outputs(41)) or (layer0_outputs(2232)));
    outputs(989) <= not(layer0_outputs(1468));
    outputs(990) <= not(layer0_outputs(791));
    outputs(991) <= not(layer0_outputs(1075));
    outputs(992) <= layer0_outputs(145);
    outputs(993) <= not((layer0_outputs(2226)) and (layer0_outputs(1269)));
    outputs(994) <= not(layer0_outputs(1926));
    outputs(995) <= layer0_outputs(659);
    outputs(996) <= not((layer0_outputs(2387)) and (layer0_outputs(580)));
    outputs(997) <= not(layer0_outputs(1476));
    outputs(998) <= (layer0_outputs(1869)) and not (layer0_outputs(532));
    outputs(999) <= not((layer0_outputs(586)) or (layer0_outputs(1164)));
    outputs(1000) <= not(layer0_outputs(1984));
    outputs(1001) <= not(layer0_outputs(2333)) or (layer0_outputs(505));
    outputs(1002) <= not(layer0_outputs(292));
    outputs(1003) <= layer0_outputs(1550);
    outputs(1004) <= (layer0_outputs(868)) and (layer0_outputs(2007));
    outputs(1005) <= not(layer0_outputs(1986));
    outputs(1006) <= not(layer0_outputs(2390));
    outputs(1007) <= (layer0_outputs(1371)) and (layer0_outputs(103));
    outputs(1008) <= layer0_outputs(2504);
    outputs(1009) <= (layer0_outputs(267)) and not (layer0_outputs(660));
    outputs(1010) <= (layer0_outputs(2321)) and not (layer0_outputs(1974));
    outputs(1011) <= (layer0_outputs(42)) and not (layer0_outputs(1010));
    outputs(1012) <= layer0_outputs(1631);
    outputs(1013) <= (layer0_outputs(1721)) and not (layer0_outputs(2357));
    outputs(1014) <= (layer0_outputs(1218)) and not (layer0_outputs(675));
    outputs(1015) <= not(layer0_outputs(2364)) or (layer0_outputs(125));
    outputs(1016) <= layer0_outputs(1220);
    outputs(1017) <= (layer0_outputs(1234)) xor (layer0_outputs(821));
    outputs(1018) <= layer0_outputs(2104);
    outputs(1019) <= not((layer0_outputs(2458)) or (layer0_outputs(671)));
    outputs(1020) <= not(layer0_outputs(1780));
    outputs(1021) <= not(layer0_outputs(1148));
    outputs(1022) <= not(layer0_outputs(1688));
    outputs(1023) <= (layer0_outputs(593)) and not (layer0_outputs(1831));
    outputs(1024) <= not(layer0_outputs(638)) or (layer0_outputs(2512));
    outputs(1025) <= not(layer0_outputs(1034));
    outputs(1026) <= (layer0_outputs(1629)) and (layer0_outputs(2432));
    outputs(1027) <= not(layer0_outputs(508)) or (layer0_outputs(1671));
    outputs(1028) <= (layer0_outputs(2360)) and not (layer0_outputs(1055));
    outputs(1029) <= not(layer0_outputs(2350));
    outputs(1030) <= not(layer0_outputs(2441));
    outputs(1031) <= not(layer0_outputs(1576));
    outputs(1032) <= not(layer0_outputs(477));
    outputs(1033) <= (layer0_outputs(2055)) and (layer0_outputs(1144));
    outputs(1034) <= not(layer0_outputs(1678));
    outputs(1035) <= not(layer0_outputs(1291));
    outputs(1036) <= layer0_outputs(95);
    outputs(1037) <= not(layer0_outputs(1514));
    outputs(1038) <= (layer0_outputs(2457)) and not (layer0_outputs(622));
    outputs(1039) <= not(layer0_outputs(624));
    outputs(1040) <= (layer0_outputs(2328)) and not (layer0_outputs(2524));
    outputs(1041) <= (layer0_outputs(453)) and (layer0_outputs(1421));
    outputs(1042) <= (layer0_outputs(1828)) or (layer0_outputs(2088));
    outputs(1043) <= not(layer0_outputs(698));
    outputs(1044) <= (layer0_outputs(1752)) and not (layer0_outputs(69));
    outputs(1045) <= not(layer0_outputs(412));
    outputs(1046) <= not(layer0_outputs(1849));
    outputs(1047) <= not((layer0_outputs(640)) or (layer0_outputs(2261)));
    outputs(1048) <= (layer0_outputs(1196)) and not (layer0_outputs(2392));
    outputs(1049) <= layer0_outputs(214);
    outputs(1050) <= (layer0_outputs(1345)) or (layer0_outputs(2304));
    outputs(1051) <= (layer0_outputs(1997)) and not (layer0_outputs(2540));
    outputs(1052) <= layer0_outputs(887);
    outputs(1053) <= not((layer0_outputs(2085)) or (layer0_outputs(140)));
    outputs(1054) <= (layer0_outputs(2041)) and (layer0_outputs(1634));
    outputs(1055) <= not(layer0_outputs(1));
    outputs(1056) <= layer0_outputs(1460);
    outputs(1057) <= layer0_outputs(1790);
    outputs(1058) <= not((layer0_outputs(851)) or (layer0_outputs(1464)));
    outputs(1059) <= (layer0_outputs(620)) and (layer0_outputs(1230));
    outputs(1060) <= (layer0_outputs(651)) and (layer0_outputs(666));
    outputs(1061) <= not((layer0_outputs(2485)) or (layer0_outputs(1470)));
    outputs(1062) <= not(layer0_outputs(2544));
    outputs(1063) <= (layer0_outputs(498)) and not (layer0_outputs(429));
    outputs(1064) <= layer0_outputs(2172);
    outputs(1065) <= (layer0_outputs(1577)) and not (layer0_outputs(2054));
    outputs(1066) <= not(layer0_outputs(298));
    outputs(1067) <= (layer0_outputs(786)) and not (layer0_outputs(1486));
    outputs(1068) <= not(layer0_outputs(390));
    outputs(1069) <= not(layer0_outputs(635)) or (layer0_outputs(531));
    outputs(1070) <= not(layer0_outputs(1673));
    outputs(1071) <= not(layer0_outputs(1498));
    outputs(1072) <= layer0_outputs(2455);
    outputs(1073) <= not((layer0_outputs(713)) or (layer0_outputs(1094)));
    outputs(1074) <= layer0_outputs(1126);
    outputs(1075) <= layer0_outputs(2029);
    outputs(1076) <= not(layer0_outputs(2302));
    outputs(1077) <= layer0_outputs(2049);
    outputs(1078) <= not(layer0_outputs(143));
    outputs(1079) <= layer0_outputs(2339);
    outputs(1080) <= layer0_outputs(880);
    outputs(1081) <= not(layer0_outputs(1424));
    outputs(1082) <= not((layer0_outputs(1978)) or (layer0_outputs(1643)));
    outputs(1083) <= layer0_outputs(1311);
    outputs(1084) <= layer0_outputs(2327);
    outputs(1085) <= layer0_outputs(2450);
    outputs(1086) <= not((layer0_outputs(1484)) or (layer0_outputs(70)));
    outputs(1087) <= not(layer0_outputs(1967));
    outputs(1088) <= (layer0_outputs(1028)) and not (layer0_outputs(1001));
    outputs(1089) <= not((layer0_outputs(697)) or (layer0_outputs(938)));
    outputs(1090) <= layer0_outputs(1879);
    outputs(1091) <= layer0_outputs(605);
    outputs(1092) <= layer0_outputs(1077);
    outputs(1093) <= not(layer0_outputs(1131));
    outputs(1094) <= layer0_outputs(300);
    outputs(1095) <= not((layer0_outputs(24)) and (layer0_outputs(1047)));
    outputs(1096) <= not(layer0_outputs(619));
    outputs(1097) <= (layer0_outputs(1596)) and not (layer0_outputs(1563));
    outputs(1098) <= not(layer0_outputs(2190));
    outputs(1099) <= layer0_outputs(2407);
    outputs(1100) <= not((layer0_outputs(1338)) xor (layer0_outputs(1027)));
    outputs(1101) <= not(layer0_outputs(902));
    outputs(1102) <= layer0_outputs(110);
    outputs(1103) <= (layer0_outputs(702)) or (layer0_outputs(117));
    outputs(1104) <= layer0_outputs(1078);
    outputs(1105) <= layer0_outputs(112);
    outputs(1106) <= (layer0_outputs(1736)) and (layer0_outputs(863));
    outputs(1107) <= layer0_outputs(852);
    outputs(1108) <= (layer0_outputs(1791)) and not (layer0_outputs(1031));
    outputs(1109) <= layer0_outputs(1342);
    outputs(1110) <= (layer0_outputs(440)) and not (layer0_outputs(784));
    outputs(1111) <= (layer0_outputs(1638)) and not (layer0_outputs(1876));
    outputs(1112) <= not(layer0_outputs(116)) or (layer0_outputs(2276));
    outputs(1113) <= not(layer0_outputs(861)) or (layer0_outputs(1452));
    outputs(1114) <= not(layer0_outputs(2390));
    outputs(1115) <= layer0_outputs(572);
    outputs(1116) <= layer0_outputs(297);
    outputs(1117) <= layer0_outputs(2090);
    outputs(1118) <= (layer0_outputs(1756)) or (layer0_outputs(1407));
    outputs(1119) <= not((layer0_outputs(1272)) and (layer0_outputs(1005)));
    outputs(1120) <= layer0_outputs(1380);
    outputs(1121) <= (layer0_outputs(1059)) and (layer0_outputs(1064));
    outputs(1122) <= not(layer0_outputs(1332));
    outputs(1123) <= layer0_outputs(365);
    outputs(1124) <= layer0_outputs(1682);
    outputs(1125) <= layer0_outputs(761);
    outputs(1126) <= layer0_outputs(2148);
    outputs(1127) <= layer0_outputs(1874);
    outputs(1128) <= layer0_outputs(1462);
    outputs(1129) <= not((layer0_outputs(2297)) or (layer0_outputs(731)));
    outputs(1130) <= (layer0_outputs(989)) and (layer0_outputs(2009));
    outputs(1131) <= (layer0_outputs(1809)) and (layer0_outputs(278));
    outputs(1132) <= layer0_outputs(2372);
    outputs(1133) <= layer0_outputs(703);
    outputs(1134) <= not((layer0_outputs(2183)) xor (layer0_outputs(2141)));
    outputs(1135) <= (layer0_outputs(1559)) or (layer0_outputs(1743));
    outputs(1136) <= (layer0_outputs(1091)) or (layer0_outputs(309));
    outputs(1137) <= not((layer0_outputs(705)) or (layer0_outputs(814)));
    outputs(1138) <= not(layer0_outputs(1869));
    outputs(1139) <= not(layer0_outputs(76));
    outputs(1140) <= layer0_outputs(831);
    outputs(1141) <= layer0_outputs(218);
    outputs(1142) <= not(layer0_outputs(656));
    outputs(1143) <= layer0_outputs(2450);
    outputs(1144) <= layer0_outputs(1394);
    outputs(1145) <= not(layer0_outputs(206));
    outputs(1146) <= not(layer0_outputs(611));
    outputs(1147) <= not((layer0_outputs(1190)) or (layer0_outputs(966)));
    outputs(1148) <= (layer0_outputs(1324)) and not (layer0_outputs(1279));
    outputs(1149) <= layer0_outputs(1510);
    outputs(1150) <= (layer0_outputs(1650)) and (layer0_outputs(2329));
    outputs(1151) <= not(layer0_outputs(1581)) or (layer0_outputs(1413));
    outputs(1152) <= layer0_outputs(2529);
    outputs(1153) <= not((layer0_outputs(1295)) xor (layer0_outputs(181)));
    outputs(1154) <= not(layer0_outputs(159)) or (layer0_outputs(1143));
    outputs(1155) <= (layer0_outputs(497)) or (layer0_outputs(1467));
    outputs(1156) <= not((layer0_outputs(124)) xor (layer0_outputs(1231)));
    outputs(1157) <= (layer0_outputs(1325)) or (layer0_outputs(1011));
    outputs(1158) <= not(layer0_outputs(1240)) or (layer0_outputs(1773));
    outputs(1159) <= not(layer0_outputs(1116));
    outputs(1160) <= not(layer0_outputs(1795)) or (layer0_outputs(1748));
    outputs(1161) <= not(layer0_outputs(819));
    outputs(1162) <= not(layer0_outputs(1228));
    outputs(1163) <= not(layer0_outputs(1335));
    outputs(1164) <= (layer0_outputs(2346)) and not (layer0_outputs(1474));
    outputs(1165) <= (layer0_outputs(805)) and not (layer0_outputs(1571));
    outputs(1166) <= layer0_outputs(2144);
    outputs(1167) <= (layer0_outputs(1621)) and not (layer0_outputs(2158));
    outputs(1168) <= not(layer0_outputs(1121)) or (layer0_outputs(462));
    outputs(1169) <= not(layer0_outputs(204));
    outputs(1170) <= not((layer0_outputs(870)) or (layer0_outputs(253)));
    outputs(1171) <= layer0_outputs(214);
    outputs(1172) <= not(layer0_outputs(68));
    outputs(1173) <= not(layer0_outputs(160));
    outputs(1174) <= not(layer0_outputs(443));
    outputs(1175) <= not(layer0_outputs(624)) or (layer0_outputs(2063));
    outputs(1176) <= not(layer0_outputs(369));
    outputs(1177) <= not(layer0_outputs(1774));
    outputs(1178) <= not((layer0_outputs(9)) or (layer0_outputs(2071)));
    outputs(1179) <= layer0_outputs(2491);
    outputs(1180) <= (layer0_outputs(387)) and (layer0_outputs(2506));
    outputs(1181) <= (layer0_outputs(1479)) or (layer0_outputs(346));
    outputs(1182) <= not(layer0_outputs(578)) or (layer0_outputs(1870));
    outputs(1183) <= layer0_outputs(2467);
    outputs(1184) <= not(layer0_outputs(824));
    outputs(1185) <= layer0_outputs(1374);
    outputs(1186) <= (layer0_outputs(2393)) and (layer0_outputs(1554));
    outputs(1187) <= not(layer0_outputs(601));
    outputs(1188) <= (layer0_outputs(231)) and not (layer0_outputs(1907));
    outputs(1189) <= (layer0_outputs(1668)) and not (layer0_outputs(2428));
    outputs(1190) <= (layer0_outputs(2494)) and not (layer0_outputs(261));
    outputs(1191) <= (layer0_outputs(213)) and (layer0_outputs(2003));
    outputs(1192) <= (layer0_outputs(2223)) and not (layer0_outputs(480));
    outputs(1193) <= not(layer0_outputs(242));
    outputs(1194) <= not(layer0_outputs(1038)) or (layer0_outputs(822));
    outputs(1195) <= not(layer0_outputs(44));
    outputs(1196) <= not(layer0_outputs(1659)) or (layer0_outputs(2280));
    outputs(1197) <= (layer0_outputs(736)) and (layer0_outputs(975));
    outputs(1198) <= (layer0_outputs(820)) and not (layer0_outputs(407));
    outputs(1199) <= layer0_outputs(2388);
    outputs(1200) <= not(layer0_outputs(139));
    outputs(1201) <= layer0_outputs(237);
    outputs(1202) <= not(layer0_outputs(92));
    outputs(1203) <= not((layer0_outputs(2205)) and (layer0_outputs(2163)));
    outputs(1204) <= (layer0_outputs(1446)) and not (layer0_outputs(86));
    outputs(1205) <= (layer0_outputs(1216)) and not (layer0_outputs(2428));
    outputs(1206) <= not(layer0_outputs(134));
    outputs(1207) <= not(layer0_outputs(598));
    outputs(1208) <= not(layer0_outputs(2343));
    outputs(1209) <= not(layer0_outputs(2181));
    outputs(1210) <= not(layer0_outputs(1187));
    outputs(1211) <= not(layer0_outputs(2249));
    outputs(1212) <= layer0_outputs(2143);
    outputs(1213) <= not(layer0_outputs(1765));
    outputs(1214) <= not(layer0_outputs(54));
    outputs(1215) <= layer0_outputs(2023);
    outputs(1216) <= not(layer0_outputs(1854));
    outputs(1217) <= not(layer0_outputs(313)) or (layer0_outputs(674));
    outputs(1218) <= not((layer0_outputs(1517)) and (layer0_outputs(846)));
    outputs(1219) <= (layer0_outputs(75)) and (layer0_outputs(1388));
    outputs(1220) <= not(layer0_outputs(1171)) or (layer0_outputs(1079));
    outputs(1221) <= not(layer0_outputs(167));
    outputs(1222) <= not(layer0_outputs(1504));
    outputs(1223) <= not(layer0_outputs(1747));
    outputs(1224) <= not(layer0_outputs(1636));
    outputs(1225) <= not((layer0_outputs(161)) or (layer0_outputs(598)));
    outputs(1226) <= (layer0_outputs(1697)) or (layer0_outputs(1467));
    outputs(1227) <= not(layer0_outputs(1346));
    outputs(1228) <= not((layer0_outputs(1399)) and (layer0_outputs(2318)));
    outputs(1229) <= not(layer0_outputs(939));
    outputs(1230) <= (layer0_outputs(2329)) or (layer0_outputs(1091));
    outputs(1231) <= (layer0_outputs(2212)) and (layer0_outputs(152));
    outputs(1232) <= not(layer0_outputs(1041));
    outputs(1233) <= not((layer0_outputs(1089)) or (layer0_outputs(1349)));
    outputs(1234) <= layer0_outputs(59);
    outputs(1235) <= layer0_outputs(736);
    outputs(1236) <= not(layer0_outputs(1280)) or (layer0_outputs(164));
    outputs(1237) <= layer0_outputs(1454);
    outputs(1238) <= (layer0_outputs(2379)) and (layer0_outputs(881));
    outputs(1239) <= layer0_outputs(879);
    outputs(1240) <= (layer0_outputs(149)) and not (layer0_outputs(1594));
    outputs(1241) <= not((layer0_outputs(1349)) xor (layer0_outputs(2246)));
    outputs(1242) <= not(layer0_outputs(1137));
    outputs(1243) <= (layer0_outputs(2453)) and not (layer0_outputs(397));
    outputs(1244) <= layer0_outputs(1366);
    outputs(1245) <= not(layer0_outputs(356));
    outputs(1246) <= (layer0_outputs(726)) or (layer0_outputs(2009));
    outputs(1247) <= not(layer0_outputs(1811));
    outputs(1248) <= layer0_outputs(2347);
    outputs(1249) <= (layer0_outputs(2538)) and (layer0_outputs(1691));
    outputs(1250) <= not((layer0_outputs(578)) and (layer0_outputs(2271)));
    outputs(1251) <= layer0_outputs(1603);
    outputs(1252) <= layer0_outputs(585);
    outputs(1253) <= (layer0_outputs(1352)) and not (layer0_outputs(341));
    outputs(1254) <= layer0_outputs(896);
    outputs(1255) <= not(layer0_outputs(1054));
    outputs(1256) <= layer0_outputs(1518);
    outputs(1257) <= not(layer0_outputs(1473)) or (layer0_outputs(597));
    outputs(1258) <= (layer0_outputs(1273)) or (layer0_outputs(1024));
    outputs(1259) <= not(layer0_outputs(718));
    outputs(1260) <= layer0_outputs(1203);
    outputs(1261) <= (layer0_outputs(212)) and (layer0_outputs(1308));
    outputs(1262) <= not(layer0_outputs(981));
    outputs(1263) <= (layer0_outputs(413)) xor (layer0_outputs(2272));
    outputs(1264) <= layer0_outputs(1605);
    outputs(1265) <= layer0_outputs(917);
    outputs(1266) <= not(layer0_outputs(1262));
    outputs(1267) <= not(layer0_outputs(1494));
    outputs(1268) <= (layer0_outputs(844)) and not (layer0_outputs(418));
    outputs(1269) <= (layer0_outputs(842)) or (layer0_outputs(2424));
    outputs(1270) <= not((layer0_outputs(2038)) and (layer0_outputs(1680)));
    outputs(1271) <= layer0_outputs(563);
    outputs(1272) <= (layer0_outputs(1794)) and (layer0_outputs(507));
    outputs(1273) <= not(layer0_outputs(2551));
    outputs(1274) <= layer0_outputs(2228);
    outputs(1275) <= not((layer0_outputs(1466)) or (layer0_outputs(2558)));
    outputs(1276) <= (layer0_outputs(2436)) and not (layer0_outputs(715));
    outputs(1277) <= layer0_outputs(908);
    outputs(1278) <= (layer0_outputs(1882)) and (layer0_outputs(1963));
    outputs(1279) <= layer0_outputs(445);
    outputs(1280) <= not((layer0_outputs(1888)) and (layer0_outputs(826)));
    outputs(1281) <= not(layer0_outputs(1161));
    outputs(1282) <= (layer0_outputs(1477)) and (layer0_outputs(640));
    outputs(1283) <= (layer0_outputs(1030)) and not (layer0_outputs(997));
    outputs(1284) <= not(layer0_outputs(2010));
    outputs(1285) <= layer0_outputs(925);
    outputs(1286) <= not(layer0_outputs(1741));
    outputs(1287) <= (layer0_outputs(743)) and (layer0_outputs(798));
    outputs(1288) <= (layer0_outputs(2230)) and not (layer0_outputs(2017));
    outputs(1289) <= layer0_outputs(1272);
    outputs(1290) <= (layer0_outputs(2310)) and (layer0_outputs(1608));
    outputs(1291) <= (layer0_outputs(556)) xor (layer0_outputs(2527));
    outputs(1292) <= not(layer0_outputs(320));
    outputs(1293) <= not(layer0_outputs(2079));
    outputs(1294) <= not(layer0_outputs(142)) or (layer0_outputs(1958));
    outputs(1295) <= (layer0_outputs(942)) xor (layer0_outputs(2345));
    outputs(1296) <= not(layer0_outputs(1100));
    outputs(1297) <= not((layer0_outputs(2078)) xor (layer0_outputs(482)));
    outputs(1298) <= not((layer0_outputs(2452)) or (layer0_outputs(1065)));
    outputs(1299) <= (layer0_outputs(2103)) and (layer0_outputs(1776));
    outputs(1300) <= not(layer0_outputs(2059));
    outputs(1301) <= not(layer0_outputs(679));
    outputs(1302) <= not((layer0_outputs(2108)) or (layer0_outputs(101)));
    outputs(1303) <= not((layer0_outputs(1536)) and (layer0_outputs(2534)));
    outputs(1304) <= (layer0_outputs(2480)) xor (layer0_outputs(1942));
    outputs(1305) <= not((layer0_outputs(570)) xor (layer0_outputs(2382)));
    outputs(1306) <= layer0_outputs(1955);
    outputs(1307) <= layer0_outputs(2282);
    outputs(1308) <= not(layer0_outputs(2363));
    outputs(1309) <= layer0_outputs(1939);
    outputs(1310) <= (layer0_outputs(2469)) xor (layer0_outputs(464));
    outputs(1311) <= not(layer0_outputs(1411)) or (layer0_outputs(1354));
    outputs(1312) <= layer0_outputs(1097);
    outputs(1313) <= layer0_outputs(1690);
    outputs(1314) <= layer0_outputs(645);
    outputs(1315) <= layer0_outputs(1002);
    outputs(1316) <= not(layer0_outputs(1491)) or (layer0_outputs(1821));
    outputs(1317) <= (layer0_outputs(993)) and not (layer0_outputs(1842));
    outputs(1318) <= (layer0_outputs(1408)) xor (layer0_outputs(654));
    outputs(1319) <= layer0_outputs(582);
    outputs(1320) <= layer0_outputs(18);
    outputs(1321) <= not(layer0_outputs(780));
    outputs(1322) <= (layer0_outputs(355)) xor (layer0_outputs(442));
    outputs(1323) <= not((layer0_outputs(2421)) or (layer0_outputs(207)));
    outputs(1324) <= layer0_outputs(1372);
    outputs(1325) <= not(layer0_outputs(178));
    outputs(1326) <= (layer0_outputs(287)) and not (layer0_outputs(859));
    outputs(1327) <= not(layer0_outputs(2308));
    outputs(1328) <= not(layer0_outputs(141));
    outputs(1329) <= (layer0_outputs(1483)) and (layer0_outputs(1227));
    outputs(1330) <= layer0_outputs(2167);
    outputs(1331) <= not((layer0_outputs(1418)) or (layer0_outputs(394)));
    outputs(1332) <= (layer0_outputs(99)) and not (layer0_outputs(2496));
    outputs(1333) <= layer0_outputs(1140);
    outputs(1334) <= (layer0_outputs(1158)) and (layer0_outputs(787));
    outputs(1335) <= (layer0_outputs(1739)) and not (layer0_outputs(1159));
    outputs(1336) <= (layer0_outputs(1620)) and not (layer0_outputs(833));
    outputs(1337) <= not((layer0_outputs(1969)) or (layer0_outputs(31)));
    outputs(1338) <= not((layer0_outputs(1755)) or (layer0_outputs(1742)));
    outputs(1339) <= layer0_outputs(2062);
    outputs(1340) <= (layer0_outputs(18)) and not (layer0_outputs(1746));
    outputs(1341) <= layer0_outputs(2127);
    outputs(1342) <= not(layer0_outputs(386));
    outputs(1343) <= not((layer0_outputs(1461)) xor (layer0_outputs(856)));
    outputs(1344) <= not(layer0_outputs(1314));
    outputs(1345) <= (layer0_outputs(238)) and (layer0_outputs(788));
    outputs(1346) <= (layer0_outputs(1662)) xor (layer0_outputs(2031));
    outputs(1347) <= not((layer0_outputs(621)) or (layer0_outputs(2035)));
    outputs(1348) <= layer0_outputs(1086);
    outputs(1349) <= not(layer0_outputs(395));
    outputs(1350) <= not(layer0_outputs(1393));
    outputs(1351) <= not(layer0_outputs(934));
    outputs(1352) <= not(layer0_outputs(58));
    outputs(1353) <= layer0_outputs(1929);
    outputs(1354) <= (layer0_outputs(1256)) and (layer0_outputs(803));
    outputs(1355) <= not((layer0_outputs(831)) or (layer0_outputs(469)));
    outputs(1356) <= (layer0_outputs(1160)) xor (layer0_outputs(129));
    outputs(1357) <= not(layer0_outputs(1302));
    outputs(1358) <= not((layer0_outputs(2331)) xor (layer0_outputs(455)));
    outputs(1359) <= (layer0_outputs(669)) and not (layer0_outputs(1618));
    outputs(1360) <= not((layer0_outputs(297)) and (layer0_outputs(1762)));
    outputs(1361) <= (layer0_outputs(2288)) and (layer0_outputs(2480));
    outputs(1362) <= layer0_outputs(548);
    outputs(1363) <= not((layer0_outputs(2376)) and (layer0_outputs(2423)));
    outputs(1364) <= not((layer0_outputs(1590)) and (layer0_outputs(1612)));
    outputs(1365) <= not(layer0_outputs(1549));
    outputs(1366) <= (layer0_outputs(2212)) and not (layer0_outputs(1594));
    outputs(1367) <= not((layer0_outputs(2224)) and (layer0_outputs(2552)));
    outputs(1368) <= not((layer0_outputs(1856)) xor (layer0_outputs(855)));
    outputs(1369) <= (layer0_outputs(2233)) xor (layer0_outputs(757));
    outputs(1370) <= not((layer0_outputs(876)) or (layer0_outputs(968)));
    outputs(1371) <= not(layer0_outputs(2348)) or (layer0_outputs(2455));
    outputs(1372) <= (layer0_outputs(929)) and not (layer0_outputs(1392));
    outputs(1373) <= not((layer0_outputs(1480)) or (layer0_outputs(1771)));
    outputs(1374) <= (layer0_outputs(312)) and not (layer0_outputs(1534));
    outputs(1375) <= not((layer0_outputs(1029)) or (layer0_outputs(644)));
    outputs(1376) <= layer0_outputs(775);
    outputs(1377) <= (layer0_outputs(186)) and (layer0_outputs(1287));
    outputs(1378) <= layer0_outputs(1195);
    outputs(1379) <= not(layer0_outputs(858));
    outputs(1380) <= not(layer0_outputs(1941));
    outputs(1381) <= (layer0_outputs(953)) and (layer0_outputs(209));
    outputs(1382) <= layer0_outputs(1244);
    outputs(1383) <= not(layer0_outputs(1552));
    outputs(1384) <= (layer0_outputs(821)) or (layer0_outputs(465));
    outputs(1385) <= layer0_outputs(1008);
    outputs(1386) <= layer0_outputs(2490);
    outputs(1387) <= not(layer0_outputs(1492));
    outputs(1388) <= not(layer0_outputs(2361));
    outputs(1389) <= layer0_outputs(90);
    outputs(1390) <= (layer0_outputs(1158)) and (layer0_outputs(1823));
    outputs(1391) <= not((layer0_outputs(660)) or (layer0_outputs(2512)));
    outputs(1392) <= (layer0_outputs(2192)) and not (layer0_outputs(1496));
    outputs(1393) <= layer0_outputs(2446);
    outputs(1394) <= (layer0_outputs(1097)) and not (layer0_outputs(311));
    outputs(1395) <= (layer0_outputs(1310)) and not (layer0_outputs(1454));
    outputs(1396) <= (layer0_outputs(299)) and (layer0_outputs(1693));
    outputs(1397) <= (layer0_outputs(1260)) xor (layer0_outputs(2427));
    outputs(1398) <= not(layer0_outputs(495));
    outputs(1399) <= not((layer0_outputs(259)) or (layer0_outputs(1704)));
    outputs(1400) <= layer0_outputs(2551);
    outputs(1401) <= (layer0_outputs(871)) and not (layer0_outputs(776));
    outputs(1402) <= (layer0_outputs(1191)) and not (layer0_outputs(725));
    outputs(1403) <= (layer0_outputs(1406)) and not (layer0_outputs(2248));
    outputs(1404) <= (layer0_outputs(1277)) and not (layer0_outputs(273));
    outputs(1405) <= not(layer0_outputs(2028)) or (layer0_outputs(1870));
    outputs(1406) <= not(layer0_outputs(614)) or (layer0_outputs(1306));
    outputs(1407) <= not(layer0_outputs(661));
    outputs(1408) <= not((layer0_outputs(2286)) xor (layer0_outputs(2183)));
    outputs(1409) <= not(layer0_outputs(1281));
    outputs(1410) <= not(layer0_outputs(107)) or (layer0_outputs(628));
    outputs(1411) <= not(layer0_outputs(513));
    outputs(1412) <= layer0_outputs(548);
    outputs(1413) <= not(layer0_outputs(419));
    outputs(1414) <= (layer0_outputs(1104)) and not (layer0_outputs(2221));
    outputs(1415) <= (layer0_outputs(700)) and (layer0_outputs(738));
    outputs(1416) <= not(layer0_outputs(950)) or (layer0_outputs(499));
    outputs(1417) <= not(layer0_outputs(2358)) or (layer0_outputs(1648));
    outputs(1418) <= (layer0_outputs(165)) xor (layer0_outputs(1991));
    outputs(1419) <= not(layer0_outputs(1977));
    outputs(1420) <= layer0_outputs(319);
    outputs(1421) <= not(layer0_outputs(1340));
    outputs(1422) <= (layer0_outputs(2486)) xor (layer0_outputs(2449));
    outputs(1423) <= layer0_outputs(2275);
    outputs(1424) <= not((layer0_outputs(2409)) and (layer0_outputs(2121)));
    outputs(1425) <= not((layer0_outputs(1360)) xor (layer0_outputs(657)));
    outputs(1426) <= not(layer0_outputs(216));
    outputs(1427) <= not(layer0_outputs(336));
    outputs(1428) <= (layer0_outputs(2247)) and (layer0_outputs(2437));
    outputs(1429) <= layer0_outputs(781);
    outputs(1430) <= not(layer0_outputs(1505)) or (layer0_outputs(2465));
    outputs(1431) <= (layer0_outputs(827)) and (layer0_outputs(817));
    outputs(1432) <= not(layer0_outputs(1607));
    outputs(1433) <= not(layer0_outputs(1489));
    outputs(1434) <= layer0_outputs(2026);
    outputs(1435) <= not(layer0_outputs(2509));
    outputs(1436) <= layer0_outputs(710);
    outputs(1437) <= not(layer0_outputs(73));
    outputs(1438) <= not((layer0_outputs(2305)) and (layer0_outputs(1003)));
    outputs(1439) <= layer0_outputs(111);
    outputs(1440) <= layer0_outputs(1351);
    outputs(1441) <= (layer0_outputs(2479)) and not (layer0_outputs(91));
    outputs(1442) <= not((layer0_outputs(591)) or (layer0_outputs(1966)));
    outputs(1443) <= layer0_outputs(1535);
    outputs(1444) <= (layer0_outputs(2391)) and (layer0_outputs(1391));
    outputs(1445) <= (layer0_outputs(841)) and not (layer0_outputs(1495));
    outputs(1446) <= not((layer0_outputs(2198)) or (layer0_outputs(196)));
    outputs(1447) <= layer0_outputs(941);
    outputs(1448) <= not(layer0_outputs(2030));
    outputs(1449) <= not((layer0_outputs(752)) or (layer0_outputs(1393)));
    outputs(1450) <= not(layer0_outputs(511));
    outputs(1451) <= (layer0_outputs(1127)) and (layer0_outputs(663));
    outputs(1452) <= not(layer0_outputs(2378));
    outputs(1453) <= (layer0_outputs(1239)) and not (layer0_outputs(449));
    outputs(1454) <= not((layer0_outputs(1193)) and (layer0_outputs(1040)));
    outputs(1455) <= not(layer0_outputs(608));
    outputs(1456) <= not(layer0_outputs(1587));
    outputs(1457) <= layer0_outputs(1184);
    outputs(1458) <= not(layer0_outputs(122));
    outputs(1459) <= not(layer0_outputs(1877));
    outputs(1460) <= (layer0_outputs(1968)) and (layer0_outputs(1475));
    outputs(1461) <= layer0_outputs(757);
    outputs(1462) <= layer0_outputs(2109);
    outputs(1463) <= not(layer0_outputs(567)) or (layer0_outputs(849));
    outputs(1464) <= (layer0_outputs(247)) and (layer0_outputs(1589));
    outputs(1465) <= not((layer0_outputs(646)) or (layer0_outputs(629)));
    outputs(1466) <= (layer0_outputs(1429)) and (layer0_outputs(466));
    outputs(1467) <= not((layer0_outputs(1436)) xor (layer0_outputs(1025)));
    outputs(1468) <= (layer0_outputs(2394)) and (layer0_outputs(1541));
    outputs(1469) <= layer0_outputs(1769);
    outputs(1470) <= not(layer0_outputs(2142));
    outputs(1471) <= (layer0_outputs(2187)) and (layer0_outputs(2461));
    outputs(1472) <= not((layer0_outputs(2217)) xor (layer0_outputs(1886)));
    outputs(1473) <= layer0_outputs(71);
    outputs(1474) <= (layer0_outputs(1621)) and not (layer0_outputs(2053));
    outputs(1475) <= not((layer0_outputs(921)) and (layer0_outputs(524)));
    outputs(1476) <= layer0_outputs(1155);
    outputs(1477) <= (layer0_outputs(748)) xor (layer0_outputs(1118));
    outputs(1478) <= (layer0_outputs(1474)) and not (layer0_outputs(2143));
    outputs(1479) <= (layer0_outputs(1323)) and (layer0_outputs(350));
    outputs(1480) <= not(layer0_outputs(2507)) or (layer0_outputs(1585));
    outputs(1481) <= not(layer0_outputs(1025)) or (layer0_outputs(447));
    outputs(1482) <= not(layer0_outputs(1058));
    outputs(1483) <= not(layer0_outputs(1072));
    outputs(1484) <= not(layer0_outputs(446));
    outputs(1485) <= layer0_outputs(1899);
    outputs(1486) <= not(layer0_outputs(2098)) or (layer0_outputs(2298));
    outputs(1487) <= not(layer0_outputs(1868));
    outputs(1488) <= layer0_outputs(1592);
    outputs(1489) <= (layer0_outputs(2261)) and (layer0_outputs(1919));
    outputs(1490) <= not((layer0_outputs(566)) and (layer0_outputs(1847)));
    outputs(1491) <= not((layer0_outputs(434)) xor (layer0_outputs(2245)));
    outputs(1492) <= not(layer0_outputs(1558));
    outputs(1493) <= (layer0_outputs(1120)) and (layer0_outputs(1405));
    outputs(1494) <= layer0_outputs(2171);
    outputs(1495) <= layer0_outputs(43);
    outputs(1496) <= not(layer0_outputs(2447));
    outputs(1497) <= not(layer0_outputs(2475));
    outputs(1498) <= (layer0_outputs(879)) and not (layer0_outputs(1080));
    outputs(1499) <= not(layer0_outputs(273));
    outputs(1500) <= not(layer0_outputs(935));
    outputs(1501) <= (layer0_outputs(1401)) and not (layer0_outputs(1430));
    outputs(1502) <= (layer0_outputs(1532)) and not (layer0_outputs(2328));
    outputs(1503) <= not((layer0_outputs(807)) xor (layer0_outputs(89)));
    outputs(1504) <= (layer0_outputs(2199)) and (layer0_outputs(143));
    outputs(1505) <= not((layer0_outputs(2484)) xor (layer0_outputs(891)));
    outputs(1506) <= (layer0_outputs(1036)) and (layer0_outputs(883));
    outputs(1507) <= layer0_outputs(1122);
    outputs(1508) <= not(layer0_outputs(518));
    outputs(1509) <= layer0_outputs(2083);
    outputs(1510) <= not(layer0_outputs(1934));
    outputs(1511) <= layer0_outputs(14);
    outputs(1512) <= layer0_outputs(1111);
    outputs(1513) <= not(layer0_outputs(42));
    outputs(1514) <= not(layer0_outputs(615));
    outputs(1515) <= not(layer0_outputs(1767));
    outputs(1516) <= not(layer0_outputs(1827));
    outputs(1517) <= not(layer0_outputs(1368));
    outputs(1518) <= not(layer0_outputs(1647));
    outputs(1519) <= not(layer0_outputs(1435));
    outputs(1520) <= not(layer0_outputs(2352));
    outputs(1521) <= layer0_outputs(2254);
    outputs(1522) <= (layer0_outputs(790)) and (layer0_outputs(334));
    outputs(1523) <= layer0_outputs(1758);
    outputs(1524) <= not(layer0_outputs(402));
    outputs(1525) <= (layer0_outputs(1106)) and (layer0_outputs(315));
    outputs(1526) <= layer0_outputs(504);
    outputs(1527) <= (layer0_outputs(2514)) and (layer0_outputs(1886));
    outputs(1528) <= (layer0_outputs(2101)) and not (layer0_outputs(969));
    outputs(1529) <= layer0_outputs(1903);
    outputs(1530) <= not((layer0_outputs(1793)) and (layer0_outputs(1418)));
    outputs(1531) <= not(layer0_outputs(1010));
    outputs(1532) <= not((layer0_outputs(189)) or (layer0_outputs(2538)));
    outputs(1533) <= not((layer0_outputs(400)) and (layer0_outputs(530)));
    outputs(1534) <= not(layer0_outputs(1479));
    outputs(1535) <= (layer0_outputs(2262)) and not (layer0_outputs(876));
    outputs(1536) <= (layer0_outputs(2375)) and (layer0_outputs(176));
    outputs(1537) <= not(layer0_outputs(1945));
    outputs(1538) <= not(layer0_outputs(2417));
    outputs(1539) <= (layer0_outputs(727)) xor (layer0_outputs(2439));
    outputs(1540) <= layer0_outputs(504);
    outputs(1541) <= (layer0_outputs(2060)) xor (layer0_outputs(2082));
    outputs(1542) <= not((layer0_outputs(1180)) or (layer0_outputs(869)));
    outputs(1543) <= not((layer0_outputs(491)) or (layer0_outputs(685)));
    outputs(1544) <= layer0_outputs(2369);
    outputs(1545) <= layer0_outputs(1610);
    outputs(1546) <= layer0_outputs(1500);
    outputs(1547) <= (layer0_outputs(1106)) and not (layer0_outputs(1214));
    outputs(1548) <= layer0_outputs(533);
    outputs(1549) <= not((layer0_outputs(1068)) or (layer0_outputs(511)));
    outputs(1550) <= (layer0_outputs(176)) and (layer0_outputs(1219));
    outputs(1551) <= layer0_outputs(158);
    outputs(1552) <= not(layer0_outputs(1689)) or (layer0_outputs(1142));
    outputs(1553) <= layer0_outputs(2371);
    outputs(1554) <= not((layer0_outputs(427)) and (layer0_outputs(1460)));
    outputs(1555) <= not((layer0_outputs(1998)) xor (layer0_outputs(1284)));
    outputs(1556) <= not(layer0_outputs(1432));
    outputs(1557) <= (layer0_outputs(593)) and not (layer0_outputs(1459));
    outputs(1558) <= (layer0_outputs(322)) and not (layer0_outputs(1011));
    outputs(1559) <= not(layer0_outputs(239));
    outputs(1560) <= (layer0_outputs(2192)) and not (layer0_outputs(463));
    outputs(1561) <= (layer0_outputs(1910)) and not (layer0_outputs(202));
    outputs(1562) <= not(layer0_outputs(1226));
    outputs(1563) <= layer0_outputs(701);
    outputs(1564) <= (layer0_outputs(22)) and (layer0_outputs(1336));
    outputs(1565) <= layer0_outputs(2039);
    outputs(1566) <= not(layer0_outputs(403));
    outputs(1567) <= (layer0_outputs(1417)) and not (layer0_outputs(2274));
    outputs(1568) <= layer0_outputs(1274);
    outputs(1569) <= (layer0_outputs(94)) and not (layer0_outputs(2175));
    outputs(1570) <= layer0_outputs(404);
    outputs(1571) <= not(layer0_outputs(963));
    outputs(1572) <= not(layer0_outputs(1246));
    outputs(1573) <= not(layer0_outputs(1278));
    outputs(1574) <= not(layer0_outputs(1896));
    outputs(1575) <= not((layer0_outputs(787)) or (layer0_outputs(249)));
    outputs(1576) <= layer0_outputs(1108);
    outputs(1577) <= not(layer0_outputs(2523));
    outputs(1578) <= not(layer0_outputs(291));
    outputs(1579) <= not(layer0_outputs(2477));
    outputs(1580) <= layer0_outputs(205);
    outputs(1581) <= not(layer0_outputs(1892));
    outputs(1582) <= not(layer0_outputs(1799));
    outputs(1583) <= (layer0_outputs(1817)) xor (layer0_outputs(800));
    outputs(1584) <= (layer0_outputs(2528)) and not (layer0_outputs(1936));
    outputs(1585) <= layer0_outputs(497);
    outputs(1586) <= layer0_outputs(1061);
    outputs(1587) <= not((layer0_outputs(272)) and (layer0_outputs(1603)));
    outputs(1588) <= layer0_outputs(2016);
    outputs(1589) <= not(layer0_outputs(2431));
    outputs(1590) <= not(layer0_outputs(1015));
    outputs(1591) <= layer0_outputs(1255);
    outputs(1592) <= (layer0_outputs(870)) and (layer0_outputs(430));
    outputs(1593) <= not((layer0_outputs(1311)) or (layer0_outputs(2550)));
    outputs(1594) <= not(layer0_outputs(1437));
    outputs(1595) <= layer0_outputs(1960);
    outputs(1596) <= (layer0_outputs(1814)) and not (layer0_outputs(2327));
    outputs(1597) <= (layer0_outputs(1529)) and (layer0_outputs(765));
    outputs(1598) <= not(layer0_outputs(1638)) or (layer0_outputs(1383));
    outputs(1599) <= (layer0_outputs(1877)) or (layer0_outputs(1787));
    outputs(1600) <= not(layer0_outputs(271));
    outputs(1601) <= (layer0_outputs(557)) and not (layer0_outputs(1179));
    outputs(1602) <= not(layer0_outputs(1679));
    outputs(1603) <= layer0_outputs(67);
    outputs(1604) <= not(layer0_outputs(2248));
    outputs(1605) <= not(layer0_outputs(2368));
    outputs(1606) <= not(layer0_outputs(1369));
    outputs(1607) <= (layer0_outputs(1864)) and (layer0_outputs(2266));
    outputs(1608) <= not(layer0_outputs(157));
    outputs(1609) <= (layer0_outputs(1225)) and not (layer0_outputs(189));
    outputs(1610) <= layer0_outputs(57);
    outputs(1611) <= not(layer0_outputs(1989));
    outputs(1612) <= not((layer0_outputs(2454)) or (layer0_outputs(632)));
    outputs(1613) <= not((layer0_outputs(1068)) and (layer0_outputs(2286)));
    outputs(1614) <= (layer0_outputs(1309)) and not (layer0_outputs(1388));
    outputs(1615) <= not(layer0_outputs(2065)) or (layer0_outputs(2204));
    outputs(1616) <= not(layer0_outputs(2400));
    outputs(1617) <= not(layer0_outputs(2045)) or (layer0_outputs(174));
    outputs(1618) <= not(layer0_outputs(560)) or (layer0_outputs(1038));
    outputs(1619) <= not(layer0_outputs(2367));
    outputs(1620) <= not(layer0_outputs(1916));
    outputs(1621) <= not(layer0_outputs(461));
    outputs(1622) <= layer0_outputs(303);
    outputs(1623) <= (layer0_outputs(753)) and (layer0_outputs(825));
    outputs(1624) <= layer0_outputs(454);
    outputs(1625) <= not((layer0_outputs(1997)) or (layer0_outputs(2344)));
    outputs(1626) <= not(layer0_outputs(355));
    outputs(1627) <= (layer0_outputs(1183)) or (layer0_outputs(349));
    outputs(1628) <= (layer0_outputs(2408)) and not (layer0_outputs(2200));
    outputs(1629) <= layer0_outputs(1256);
    outputs(1630) <= not(layer0_outputs(391));
    outputs(1631) <= layer0_outputs(1650);
    outputs(1632) <= (layer0_outputs(866)) and not (layer0_outputs(717));
    outputs(1633) <= not(layer0_outputs(1564));
    outputs(1634) <= not(layer0_outputs(421)) or (layer0_outputs(1933));
    outputs(1635) <= (layer0_outputs(1711)) xor (layer0_outputs(169));
    outputs(1636) <= (layer0_outputs(1138)) and not (layer0_outputs(661));
    outputs(1637) <= not(layer0_outputs(1042));
    outputs(1638) <= not((layer0_outputs(2381)) or (layer0_outputs(2180)));
    outputs(1639) <= layer0_outputs(2409);
    outputs(1640) <= not((layer0_outputs(2416)) or (layer0_outputs(610)));
    outputs(1641) <= (layer0_outputs(2030)) xor (layer0_outputs(1221));
    outputs(1642) <= not(layer0_outputs(1600));
    outputs(1643) <= (layer0_outputs(2545)) and not (layer0_outputs(1578));
    outputs(1644) <= (layer0_outputs(2459)) and (layer0_outputs(2154));
    outputs(1645) <= not((layer0_outputs(1045)) or (layer0_outputs(2180)));
    outputs(1646) <= not(layer0_outputs(207));
    outputs(1647) <= (layer0_outputs(2369)) and not (layer0_outputs(1934));
    outputs(1648) <= not(layer0_outputs(1753));
    outputs(1649) <= (layer0_outputs(2246)) or (layer0_outputs(1019));
    outputs(1650) <= not((layer0_outputs(1371)) or (layer0_outputs(1282)));
    outputs(1651) <= not((layer0_outputs(1397)) xor (layer0_outputs(878)));
    outputs(1652) <= not(layer0_outputs(1117));
    outputs(1653) <= not(layer0_outputs(1961)) or (layer0_outputs(120));
    outputs(1654) <= not(layer0_outputs(17));
    outputs(1655) <= layer0_outputs(2341);
    outputs(1656) <= not(layer0_outputs(656));
    outputs(1657) <= not(layer0_outputs(1243));
    outputs(1658) <= (layer0_outputs(922)) and not (layer0_outputs(1976));
    outputs(1659) <= not(layer0_outputs(2002));
    outputs(1660) <= not(layer0_outputs(1858));
    outputs(1661) <= layer0_outputs(692);
    outputs(1662) <= layer0_outputs(1834);
    outputs(1663) <= layer0_outputs(988);
    outputs(1664) <= not((layer0_outputs(279)) or (layer0_outputs(175)));
    outputs(1665) <= (layer0_outputs(1187)) and not (layer0_outputs(2299));
    outputs(1666) <= (layer0_outputs(2490)) and not (layer0_outputs(198));
    outputs(1667) <= (layer0_outputs(2333)) and (layer0_outputs(1905));
    outputs(1668) <= (layer0_outputs(2014)) and not (layer0_outputs(1200));
    outputs(1669) <= layer0_outputs(628);
    outputs(1670) <= (layer0_outputs(2078)) and not (layer0_outputs(1863));
    outputs(1671) <= not(layer0_outputs(1738));
    outputs(1672) <= (layer0_outputs(1195)) and not (layer0_outputs(1890));
    outputs(1673) <= not(layer0_outputs(616)) or (layer0_outputs(988));
    outputs(1674) <= (layer0_outputs(2415)) xor (layer0_outputs(36));
    outputs(1675) <= not(layer0_outputs(44)) or (layer0_outputs(2133));
    outputs(1676) <= (layer0_outputs(1427)) and not (layer0_outputs(1112));
    outputs(1677) <= (layer0_outputs(2080)) and not (layer0_outputs(1419));
    outputs(1678) <= (layer0_outputs(1328)) and not (layer0_outputs(2559));
    outputs(1679) <= layer0_outputs(773);
    outputs(1680) <= layer0_outputs(1224);
    outputs(1681) <= layer0_outputs(796);
    outputs(1682) <= not(layer0_outputs(1120));
    outputs(1683) <= (layer0_outputs(1861)) xor (layer0_outputs(116));
    outputs(1684) <= (layer0_outputs(1465)) and (layer0_outputs(1370));
    outputs(1685) <= layer0_outputs(629);
    outputs(1686) <= not(layer0_outputs(860));
    outputs(1687) <= not((layer0_outputs(2057)) or (layer0_outputs(1953)));
    outputs(1688) <= (layer0_outputs(340)) and (layer0_outputs(2364));
    outputs(1689) <= layer0_outputs(133);
    outputs(1690) <= layer0_outputs(1509);
    outputs(1691) <= layer0_outputs(1110);
    outputs(1692) <= not((layer0_outputs(2406)) xor (layer0_outputs(1210)));
    outputs(1693) <= (layer0_outputs(376)) and not (layer0_outputs(975));
    outputs(1694) <= (layer0_outputs(1857)) and not (layer0_outputs(1862));
    outputs(1695) <= (layer0_outputs(78)) and not (layer0_outputs(1275));
    outputs(1696) <= not(layer0_outputs(461));
    outputs(1697) <= (layer0_outputs(538)) and not (layer0_outputs(2492));
    outputs(1698) <= not((layer0_outputs(1986)) and (layer0_outputs(337)));
    outputs(1699) <= (layer0_outputs(432)) or (layer0_outputs(793));
    outputs(1700) <= (layer0_outputs(2084)) or (layer0_outputs(668));
    outputs(1701) <= not((layer0_outputs(1126)) or (layer0_outputs(1050)));
    outputs(1702) <= not(layer0_outputs(104));
    outputs(1703) <= not((layer0_outputs(718)) xor (layer0_outputs(1086)));
    outputs(1704) <= layer0_outputs(367);
    outputs(1705) <= not(layer0_outputs(1582));
    outputs(1706) <= not(layer0_outputs(82)) or (layer0_outputs(889));
    outputs(1707) <= (layer0_outputs(905)) or (layer0_outputs(2043));
    outputs(1708) <= not(layer0_outputs(2456));
    outputs(1709) <= (layer0_outputs(45)) and (layer0_outputs(1005));
    outputs(1710) <= not((layer0_outputs(171)) and (layer0_outputs(1738)));
    outputs(1711) <= not(layer0_outputs(1445)) or (layer0_outputs(1128));
    outputs(1712) <= not(layer0_outputs(1853));
    outputs(1713) <= not((layer0_outputs(2373)) and (layer0_outputs(2004)));
    outputs(1714) <= not((layer0_outputs(2242)) or (layer0_outputs(1591)));
    outputs(1715) <= not(layer0_outputs(700));
    outputs(1716) <= layer0_outputs(829);
    outputs(1717) <= layer0_outputs(200);
    outputs(1718) <= (layer0_outputs(267)) and not (layer0_outputs(2236));
    outputs(1719) <= not(layer0_outputs(2296));
    outputs(1720) <= not(layer0_outputs(2532)) or (layer0_outputs(1932));
    outputs(1721) <= not(layer0_outputs(2290)) or (layer0_outputs(2326));
    outputs(1722) <= not((layer0_outputs(962)) xor (layer0_outputs(435)));
    outputs(1723) <= layer0_outputs(958);
    outputs(1724) <= layer0_outputs(1586);
    outputs(1725) <= (layer0_outputs(1809)) and not (layer0_outputs(307));
    outputs(1726) <= (layer0_outputs(2160)) and not (layer0_outputs(1781));
    outputs(1727) <= (layer0_outputs(528)) and not (layer0_outputs(173));
    outputs(1728) <= not(layer0_outputs(1737));
    outputs(1729) <= layer0_outputs(2382);
    outputs(1730) <= (layer0_outputs(1374)) and not (layer0_outputs(859));
    outputs(1731) <= not(layer0_outputs(296)) or (layer0_outputs(606));
    outputs(1732) <= layer0_outputs(789);
    outputs(1733) <= (layer0_outputs(1292)) and not (layer0_outputs(383));
    outputs(1734) <= (layer0_outputs(2132)) and not (layer0_outputs(2374));
    outputs(1735) <= layer0_outputs(519);
    outputs(1736) <= layer0_outputs(1729);
    outputs(1737) <= (layer0_outputs(782)) and not (layer0_outputs(1531));
    outputs(1738) <= not(layer0_outputs(1785));
    outputs(1739) <= not(layer0_outputs(1716));
    outputs(1740) <= layer0_outputs(2224);
    outputs(1741) <= (layer0_outputs(1903)) and not (layer0_outputs(601));
    outputs(1742) <= not(layer0_outputs(2349));
    outputs(1743) <= not(layer0_outputs(1450)) or (layer0_outputs(52));
    outputs(1744) <= not(layer0_outputs(806));
    outputs(1745) <= layer0_outputs(1344);
    outputs(1746) <= (layer0_outputs(932)) and (layer0_outputs(573));
    outputs(1747) <= layer0_outputs(1183);
    outputs(1748) <= not((layer0_outputs(893)) or (layer0_outputs(732)));
    outputs(1749) <= not(layer0_outputs(1376));
    outputs(1750) <= not(layer0_outputs(569));
    outputs(1751) <= not(layer0_outputs(211));
    outputs(1752) <= not(layer0_outputs(122));
    outputs(1753) <= not(layer0_outputs(1440));
    outputs(1754) <= not((layer0_outputs(1781)) or (layer0_outputs(1487)));
    outputs(1755) <= layer0_outputs(300);
    outputs(1756) <= not(layer0_outputs(1709)) or (layer0_outputs(1413));
    outputs(1757) <= (layer0_outputs(2522)) and not (layer0_outputs(805));
    outputs(1758) <= not(layer0_outputs(1380));
    outputs(1759) <= (layer0_outputs(563)) xor (layer0_outputs(1825));
    outputs(1760) <= not(layer0_outputs(649));
    outputs(1761) <= not(layer0_outputs(646)) or (layer0_outputs(2403));
    outputs(1762) <= not(layer0_outputs(2396)) or (layer0_outputs(1128));
    outputs(1763) <= layer0_outputs(1197);
    outputs(1764) <= (layer0_outputs(1722)) and not (layer0_outputs(1099));
    outputs(1765) <= (layer0_outputs(799)) and not (layer0_outputs(2301));
    outputs(1766) <= not(layer0_outputs(1253));
    outputs(1767) <= (layer0_outputs(1975)) and not (layer0_outputs(1999));
    outputs(1768) <= not(layer0_outputs(150));
    outputs(1769) <= layer0_outputs(850);
    outputs(1770) <= not(layer0_outputs(1954));
    outputs(1771) <= not(layer0_outputs(1115));
    outputs(1772) <= not((layer0_outputs(1028)) or (layer0_outputs(928)));
    outputs(1773) <= layer0_outputs(1360);
    outputs(1774) <= (layer0_outputs(478)) and not (layer0_outputs(758));
    outputs(1775) <= layer0_outputs(2291);
    outputs(1776) <= layer0_outputs(2116);
    outputs(1777) <= (layer0_outputs(1694)) and not (layer0_outputs(10));
    outputs(1778) <= (layer0_outputs(520)) and (layer0_outputs(1880));
    outputs(1779) <= layer0_outputs(351);
    outputs(1780) <= not((layer0_outputs(1290)) or (layer0_outputs(1699)));
    outputs(1781) <= (layer0_outputs(2351)) or (layer0_outputs(232));
    outputs(1782) <= layer0_outputs(2074);
    outputs(1783) <= (layer0_outputs(424)) or (layer0_outputs(1973));
    outputs(1784) <= (layer0_outputs(374)) and not (layer0_outputs(1669));
    outputs(1785) <= not((layer0_outputs(1337)) or (layer0_outputs(1503)));
    outputs(1786) <= (layer0_outputs(722)) and (layer0_outputs(2426));
    outputs(1787) <= not(layer0_outputs(2196));
    outputs(1788) <= not(layer0_outputs(1527));
    outputs(1789) <= not(layer0_outputs(1475));
    outputs(1790) <= (layer0_outputs(2042)) and (layer0_outputs(1722));
    outputs(1791) <= (layer0_outputs(1730)) and not (layer0_outputs(908));
    outputs(1792) <= layer0_outputs(60);
    outputs(1793) <= not((layer0_outputs(54)) or (layer0_outputs(1990)));
    outputs(1794) <= layer0_outputs(1780);
    outputs(1795) <= not(layer0_outputs(2530)) or (layer0_outputs(1304));
    outputs(1796) <= (layer0_outputs(2360)) and (layer0_outputs(1314));
    outputs(1797) <= not(layer0_outputs(1490));
    outputs(1798) <= not((layer0_outputs(1935)) or (layer0_outputs(1835)));
    outputs(1799) <= layer0_outputs(1622);
    outputs(1800) <= (layer0_outputs(1689)) and not (layer0_outputs(1237));
    outputs(1801) <= layer0_outputs(1442);
    outputs(1802) <= (layer0_outputs(2153)) and not (layer0_outputs(352));
    outputs(1803) <= not(layer0_outputs(1473)) or (layer0_outputs(246));
    outputs(1804) <= not(layer0_outputs(71)) or (layer0_outputs(731));
    outputs(1805) <= (layer0_outputs(1426)) and (layer0_outputs(60));
    outputs(1806) <= (layer0_outputs(1487)) and (layer0_outputs(1802));
    outputs(1807) <= layer0_outputs(514);
    outputs(1808) <= (layer0_outputs(305)) and not (layer0_outputs(2));
    outputs(1809) <= layer0_outputs(2033);
    outputs(1810) <= (layer0_outputs(1151)) and not (layer0_outputs(613));
    outputs(1811) <= (layer0_outputs(1900)) and not (layer0_outputs(575));
    outputs(1812) <= (layer0_outputs(1326)) and not (layer0_outputs(2399));
    outputs(1813) <= (layer0_outputs(888)) and not (layer0_outputs(2225));
    outputs(1814) <= layer0_outputs(1359);
    outputs(1815) <= not((layer0_outputs(1245)) and (layer0_outputs(2235)));
    outputs(1816) <= layer0_outputs(1881);
    outputs(1817) <= layer0_outputs(1288);
    outputs(1818) <= (layer0_outputs(2379)) and not (layer0_outputs(923));
    outputs(1819) <= (layer0_outputs(1560)) and not (layer0_outputs(588));
    outputs(1820) <= (layer0_outputs(1533)) or (layer0_outputs(886));
    outputs(1821) <= layer0_outputs(910);
    outputs(1822) <= (layer0_outputs(1882)) and (layer0_outputs(1134));
    outputs(1823) <= (layer0_outputs(142)) and not (layer0_outputs(540));
    outputs(1824) <= (layer0_outputs(2355)) and (layer0_outputs(1009));
    outputs(1825) <= (layer0_outputs(1612)) and not (layer0_outputs(2411));
    outputs(1826) <= not(layer0_outputs(1880));
    outputs(1827) <= layer0_outputs(800);
    outputs(1828) <= (layer0_outputs(1923)) and (layer0_outputs(457));
    outputs(1829) <= (layer0_outputs(436)) and (layer0_outputs(2433));
    outputs(1830) <= not(layer0_outputs(1193));
    outputs(1831) <= not((layer0_outputs(1450)) or (layer0_outputs(1368)));
    outputs(1832) <= (layer0_outputs(490)) and not (layer0_outputs(1366));
    outputs(1833) <= not((layer0_outputs(667)) or (layer0_outputs(737)));
    outputs(1834) <= not(layer0_outputs(763));
    outputs(1835) <= not(layer0_outputs(1772));
    outputs(1836) <= not(layer0_outputs(745));
    outputs(1837) <= (layer0_outputs(39)) and not (layer0_outputs(944));
    outputs(1838) <= not(layer0_outputs(2346));
    outputs(1839) <= (layer0_outputs(2181)) and not (layer0_outputs(324));
    outputs(1840) <= not((layer0_outputs(228)) and (layer0_outputs(1060)));
    outputs(1841) <= not((layer0_outputs(1914)) or (layer0_outputs(932)));
    outputs(1842) <= not((layer0_outputs(918)) or (layer0_outputs(1348)));
    outputs(1843) <= not((layer0_outputs(2556)) or (layer0_outputs(1401)));
    outputs(1844) <= not(layer0_outputs(2149)) or (layer0_outputs(2509));
    outputs(1845) <= not(layer0_outputs(1956));
    outputs(1846) <= layer0_outputs(556);
    outputs(1847) <= layer0_outputs(1777);
    outputs(1848) <= (layer0_outputs(314)) and (layer0_outputs(2368));
    outputs(1849) <= layer0_outputs(1246);
    outputs(1850) <= layer0_outputs(741);
    outputs(1851) <= not(layer0_outputs(2487));
    outputs(1852) <= (layer0_outputs(1889)) and (layer0_outputs(2386));
    outputs(1853) <= not(layer0_outputs(972));
    outputs(1854) <= layer0_outputs(2413);
    outputs(1855) <= layer0_outputs(211);
    outputs(1856) <= layer0_outputs(40);
    outputs(1857) <= (layer0_outputs(658)) xor (layer0_outputs(468));
    outputs(1858) <= not((layer0_outputs(485)) or (layer0_outputs(1706)));
    outputs(1859) <= layer0_outputs(291);
    outputs(1860) <= not((layer0_outputs(154)) or (layer0_outputs(534)));
    outputs(1861) <= not(layer0_outputs(248));
    outputs(1862) <= not((layer0_outputs(2126)) or (layer0_outputs(2273)));
    outputs(1863) <= not(layer0_outputs(1696));
    outputs(1864) <= (layer0_outputs(1987)) and (layer0_outputs(2269));
    outputs(1865) <= (layer0_outputs(844)) and (layer0_outputs(635));
    outputs(1866) <= not((layer0_outputs(332)) and (layer0_outputs(687)));
    outputs(1867) <= (layer0_outputs(1181)) and not (layer0_outputs(667));
    outputs(1868) <= layer0_outputs(1995);
    outputs(1869) <= not(layer0_outputs(2423));
    outputs(1870) <= layer0_outputs(785);
    outputs(1871) <= layer0_outputs(2549);
    outputs(1872) <= (layer0_outputs(898)) and (layer0_outputs(662));
    outputs(1873) <= not(layer0_outputs(2449));
    outputs(1874) <= layer0_outputs(2018);
    outputs(1875) <= (layer0_outputs(2488)) and not (layer0_outputs(763));
    outputs(1876) <= (layer0_outputs(2243)) and not (layer0_outputs(525));
    outputs(1877) <= layer0_outputs(1170);
    outputs(1878) <= (layer0_outputs(1579)) and not (layer0_outputs(331));
    outputs(1879) <= not((layer0_outputs(1247)) or (layer0_outputs(1645)));
    outputs(1880) <= not(layer0_outputs(1008));
    outputs(1881) <= (layer0_outputs(1852)) and not (layer0_outputs(106));
    outputs(1882) <= not((layer0_outputs(2239)) and (layer0_outputs(594)));
    outputs(1883) <= not(layer0_outputs(1457));
    outputs(1884) <= not(layer0_outputs(1749));
    outputs(1885) <= not(layer0_outputs(306)) or (layer0_outputs(191));
    outputs(1886) <= (layer0_outputs(148)) and (layer0_outputs(433));
    outputs(1887) <= layer0_outputs(545);
    outputs(1888) <= not(layer0_outputs(132)) or (layer0_outputs(1103));
    outputs(1889) <= (layer0_outputs(2037)) and not (layer0_outputs(2430));
    outputs(1890) <= (layer0_outputs(1853)) and not (layer0_outputs(2100));
    outputs(1891) <= not(layer0_outputs(243));
    outputs(1892) <= not(layer0_outputs(1822)) or (layer0_outputs(2451));
    outputs(1893) <= not(layer0_outputs(476));
    outputs(1894) <= layer0_outputs(1134);
    outputs(1895) <= not((layer0_outputs(737)) and (layer0_outputs(2317)));
    outputs(1896) <= (layer0_outputs(2526)) and not (layer0_outputs(2510));
    outputs(1897) <= layer0_outputs(1410);
    outputs(1898) <= (layer0_outputs(680)) and not (layer0_outputs(926));
    outputs(1899) <= (layer0_outputs(751)) and (layer0_outputs(1978));
    outputs(1900) <= (layer0_outputs(1260)) and not (layer0_outputs(235));
    outputs(1901) <= (layer0_outputs(1497)) and not (layer0_outputs(358));
    outputs(1902) <= layer0_outputs(1365);
    outputs(1903) <= layer0_outputs(66);
    outputs(1904) <= not(layer0_outputs(1942));
    outputs(1905) <= not((layer0_outputs(1277)) or (layer0_outputs(804)));
    outputs(1906) <= (layer0_outputs(715)) and (layer0_outputs(1112));
    outputs(1907) <= not(layer0_outputs(1536));
    outputs(1908) <= (layer0_outputs(1214)) xor (layer0_outputs(182));
    outputs(1909) <= (layer0_outputs(182)) and (layer0_outputs(2429));
    outputs(1910) <= layer0_outputs(1375);
    outputs(1911) <= (layer0_outputs(399)) and not (layer0_outputs(2164));
    outputs(1912) <= (layer0_outputs(2113)) and not (layer0_outputs(2510));
    outputs(1913) <= not(layer0_outputs(618));
    outputs(1914) <= not(layer0_outputs(745));
    outputs(1915) <= layer0_outputs(2193);
    outputs(1916) <= not(layer0_outputs(2150));
    outputs(1917) <= not(layer0_outputs(842));
    outputs(1918) <= not(layer0_outputs(13));
    outputs(1919) <= layer0_outputs(1840);
    outputs(1920) <= (layer0_outputs(1928)) and not (layer0_outputs(1588));
    outputs(1921) <= (layer0_outputs(347)) and not (layer0_outputs(1796));
    outputs(1922) <= not((layer0_outputs(411)) or (layer0_outputs(1244)));
    outputs(1923) <= (layer0_outputs(2338)) and not (layer0_outputs(600));
    outputs(1924) <= not((layer0_outputs(2172)) or (layer0_outputs(768)));
    outputs(1925) <= layer0_outputs(1976);
    outputs(1926) <= (layer0_outputs(51)) and not (layer0_outputs(1909));
    outputs(1927) <= not(layer0_outputs(726));
    outputs(1928) <= not(layer0_outputs(1373));
    outputs(1929) <= layer0_outputs(1334);
    outputs(1930) <= (layer0_outputs(546)) and not (layer0_outputs(1789));
    outputs(1931) <= not(layer0_outputs(1630));
    outputs(1932) <= (layer0_outputs(489)) and (layer0_outputs(1243));
    outputs(1933) <= not(layer0_outputs(325));
    outputs(1934) <= layer0_outputs(513);
    outputs(1935) <= not(layer0_outputs(1701));
    outputs(1936) <= layer0_outputs(56);
    outputs(1937) <= (layer0_outputs(608)) xor (layer0_outputs(1353));
    outputs(1938) <= not(layer0_outputs(1176)) or (layer0_outputs(1988));
    outputs(1939) <= not((layer0_outputs(474)) or (layer0_outputs(1805)));
    outputs(1940) <= not(layer0_outputs(1235));
    outputs(1941) <= layer0_outputs(2533);
    outputs(1942) <= (layer0_outputs(764)) xor (layer0_outputs(1048));
    outputs(1943) <= (layer0_outputs(1420)) and (layer0_outputs(749));
    outputs(1944) <= (layer0_outputs(1250)) and not (layer0_outputs(1384));
    outputs(1945) <= (layer0_outputs(2177)) or (layer0_outputs(1014));
    outputs(1946) <= layer0_outputs(709);
    outputs(1947) <= (layer0_outputs(218)) and not (layer0_outputs(1241));
    outputs(1948) <= (layer0_outputs(444)) and (layer0_outputs(2281));
    outputs(1949) <= (layer0_outputs(2122)) and not (layer0_outputs(2463));
    outputs(1950) <= (layer0_outputs(2322)) and not (layer0_outputs(227));
    outputs(1951) <= not(layer0_outputs(1238));
    outputs(1952) <= (layer0_outputs(472)) or (layer0_outputs(1322));
    outputs(1953) <= not(layer0_outputs(217));
    outputs(1954) <= layer0_outputs(741);
    outputs(1955) <= (layer0_outputs(1911)) and not (layer0_outputs(1523));
    outputs(1956) <= (layer0_outputs(1637)) and (layer0_outputs(767));
    outputs(1957) <= not(layer0_outputs(627));
    outputs(1958) <= not((layer0_outputs(79)) or (layer0_outputs(864)));
    outputs(1959) <= (layer0_outputs(1686)) and not (layer0_outputs(1731));
    outputs(1960) <= (layer0_outputs(2056)) and (layer0_outputs(484));
    outputs(1961) <= layer0_outputs(2527);
    outputs(1962) <= layer0_outputs(1129);
    outputs(1963) <= not(layer0_outputs(2335));
    outputs(1964) <= (layer0_outputs(1253)) and not (layer0_outputs(1728));
    outputs(1965) <= (layer0_outputs(2094)) and not (layer0_outputs(1471));
    outputs(1966) <= (layer0_outputs(758)) and not (layer0_outputs(1165));
    outputs(1967) <= (layer0_outputs(1806)) and not (layer0_outputs(2019));
    outputs(1968) <= not(layer0_outputs(335));
    outputs(1969) <= layer0_outputs(2441);
    outputs(1970) <= layer0_outputs(162);
    outputs(1971) <= (layer0_outputs(1223)) and not (layer0_outputs(1671));
    outputs(1972) <= not((layer0_outputs(2025)) or (layer0_outputs(1855)));
    outputs(1973) <= not(layer0_outputs(359));
    outputs(1974) <= (layer0_outputs(1162)) and (layer0_outputs(1712));
    outputs(1975) <= not(layer0_outputs(2013));
    outputs(1976) <= not(layer0_outputs(1993));
    outputs(1977) <= layer0_outputs(255);
    outputs(1978) <= (layer0_outputs(669)) and not (layer0_outputs(692));
    outputs(1979) <= (layer0_outputs(826)) and not (layer0_outputs(607));
    outputs(1980) <= (layer0_outputs(484)) and not (layer0_outputs(2027));
    outputs(1981) <= (layer0_outputs(1254)) and not (layer0_outputs(1249));
    outputs(1982) <= not(layer0_outputs(1224));
    outputs(1983) <= not((layer0_outputs(540)) or (layer0_outputs(1499)));
    outputs(1984) <= (layer0_outputs(458)) and not (layer0_outputs(2411));
    outputs(1985) <= (layer0_outputs(882)) and (layer0_outputs(135));
    outputs(1986) <= not(layer0_outputs(393));
    outputs(1987) <= layer0_outputs(15);
    outputs(1988) <= not(layer0_outputs(871)) or (layer0_outputs(873));
    outputs(1989) <= (layer0_outputs(712)) and (layer0_outputs(549));
    outputs(1990) <= not(layer0_outputs(589));
    outputs(1991) <= not(layer0_outputs(2259));
    outputs(1992) <= layer0_outputs(1741);
    outputs(1993) <= (layer0_outputs(460)) and not (layer0_outputs(672));
    outputs(1994) <= not((layer0_outputs(708)) or (layer0_outputs(2485)));
    outputs(1995) <= layer0_outputs(2052);
    outputs(1996) <= (layer0_outputs(1818)) xor (layer0_outputs(1018));
    outputs(1997) <= not(layer0_outputs(1599));
    outputs(1998) <= not(layer0_outputs(1696));
    outputs(1999) <= not(layer0_outputs(973));
    outputs(2000) <= not((layer0_outputs(2335)) or (layer0_outputs(633)));
    outputs(2001) <= (layer0_outputs(135)) and not (layer0_outputs(2482));
    outputs(2002) <= (layer0_outputs(162)) and not (layer0_outputs(420));
    outputs(2003) <= (layer0_outputs(2012)) and (layer0_outputs(1139));
    outputs(2004) <= not((layer0_outputs(1384)) and (layer0_outputs(845)));
    outputs(2005) <= not(layer0_outputs(644));
    outputs(2006) <= not(layer0_outputs(443));
    outputs(2007) <= (layer0_outputs(1215)) and not (layer0_outputs(2325));
    outputs(2008) <= not(layer0_outputs(1146));
    outputs(2009) <= layer0_outputs(1949);
    outputs(2010) <= layer0_outputs(1203);
    outputs(2011) <= layer0_outputs(144);
    outputs(2012) <= layer0_outputs(751);
    outputs(2013) <= (layer0_outputs(1943)) and (layer0_outputs(179));
    outputs(2014) <= (layer0_outputs(2182)) and not (layer0_outputs(774));
    outputs(2015) <= layer0_outputs(1867);
    outputs(2016) <= layer0_outputs(1954);
    outputs(2017) <= not(layer0_outputs(342));
    outputs(2018) <= not(layer0_outputs(1833));
    outputs(2019) <= not((layer0_outputs(1051)) xor (layer0_outputs(2234)));
    outputs(2020) <= not((layer0_outputs(170)) xor (layer0_outputs(2406)));
    outputs(2021) <= not((layer0_outputs(2319)) or (layer0_outputs(275)));
    outputs(2022) <= not((layer0_outputs(2292)) or (layer0_outputs(2207)));
    outputs(2023) <= not(layer0_outputs(1620));
    outputs(2024) <= (layer0_outputs(2416)) and (layer0_outputs(382));
    outputs(2025) <= (layer0_outputs(813)) and (layer0_outputs(2500));
    outputs(2026) <= (layer0_outputs(1583)) and (layer0_outputs(819));
    outputs(2027) <= (layer0_outputs(2497)) and not (layer0_outputs(1605));
    outputs(2028) <= (layer0_outputs(2431)) and (layer0_outputs(436));
    outputs(2029) <= not((layer0_outputs(2156)) or (layer0_outputs(187)));
    outputs(2030) <= (layer0_outputs(1196)) and not (layer0_outputs(2292));
    outputs(2031) <= (layer0_outputs(1827)) and (layer0_outputs(1044));
    outputs(2032) <= not(layer0_outputs(1733)) or (layer0_outputs(897));
    outputs(2033) <= (layer0_outputs(1959)) and (layer0_outputs(1410));
    outputs(2034) <= not(layer0_outputs(421)) or (layer0_outputs(1301));
    outputs(2035) <= (layer0_outputs(657)) and not (layer0_outputs(500));
    outputs(2036) <= not(layer0_outputs(166));
    outputs(2037) <= layer0_outputs(1939);
    outputs(2038) <= not((layer0_outputs(823)) or (layer0_outputs(2077)));
    outputs(2039) <= (layer0_outputs(1921)) and not (layer0_outputs(2194));
    outputs(2040) <= (layer0_outputs(1920)) and (layer0_outputs(1965));
    outputs(2041) <= (layer0_outputs(1661)) and (layer0_outputs(1024));
    outputs(2042) <= layer0_outputs(1988);
    outputs(2043) <= layer0_outputs(1443);
    outputs(2044) <= (layer0_outputs(1481)) and not (layer0_outputs(1507));
    outputs(2045) <= layer0_outputs(750);
    outputs(2046) <= not((layer0_outputs(2306)) or (layer0_outputs(1766)));
    outputs(2047) <= layer0_outputs(1337);
    outputs(2048) <= (layer0_outputs(2448)) and not (layer0_outputs(166));
    outputs(2049) <= not(layer0_outputs(1205));
    outputs(2050) <= not(layer0_outputs(241));
    outputs(2051) <= not(layer0_outputs(163));
    outputs(2052) <= (layer0_outputs(2054)) or (layer0_outputs(974));
    outputs(2053) <= (layer0_outputs(829)) and not (layer0_outputs(2029));
    outputs(2054) <= (layer0_outputs(32)) xor (layer0_outputs(2520));
    outputs(2055) <= (layer0_outputs(2265)) or (layer0_outputs(2124));
    outputs(2056) <= (layer0_outputs(184)) or (layer0_outputs(396));
    outputs(2057) <= not((layer0_outputs(2493)) or (layer0_outputs(809)));
    outputs(2058) <= (layer0_outputs(1864)) xor (layer0_outputs(1073));
    outputs(2059) <= layer0_outputs(2508);
    outputs(2060) <= (layer0_outputs(874)) and not (layer0_outputs(2112));
    outputs(2061) <= not((layer0_outputs(1970)) and (layer0_outputs(2018)));
    outputs(2062) <= layer0_outputs(121);
    outputs(2063) <= not(layer0_outputs(1411)) or (layer0_outputs(1273));
    outputs(2064) <= not(layer0_outputs(740));
    outputs(2065) <= (layer0_outputs(2127)) or (layer0_outputs(2366));
    outputs(2066) <= not((layer0_outputs(1455)) or (layer0_outputs(1017)));
    outputs(2067) <= not(layer0_outputs(1751));
    outputs(2068) <= layer0_outputs(473);
    outputs(2069) <= not((layer0_outputs(557)) and (layer0_outputs(720)));
    outputs(2070) <= not(layer0_outputs(735));
    outputs(2071) <= layer0_outputs(1084);
    outputs(2072) <= (layer0_outputs(1930)) xor (layer0_outputs(2138));
    outputs(2073) <= not(layer0_outputs(1408));
    outputs(2074) <= (layer0_outputs(1602)) and (layer0_outputs(2301));
    outputs(2075) <= not(layer0_outputs(1945));
    outputs(2076) <= layer0_outputs(2447);
    outputs(2077) <= layer0_outputs(478);
    outputs(2078) <= not(layer0_outputs(999));
    outputs(2079) <= (layer0_outputs(1839)) and (layer0_outputs(946));
    outputs(2080) <= layer0_outputs(2384);
    outputs(2081) <= (layer0_outputs(130)) and not (layer0_outputs(2443));
    outputs(2082) <= layer0_outputs(827);
    outputs(2083) <= layer0_outputs(1392);
    outputs(2084) <= layer0_outputs(1684);
    outputs(2085) <= not(layer0_outputs(1851));
    outputs(2086) <= not(layer0_outputs(1829)) or (layer0_outputs(428));
    outputs(2087) <= not(layer0_outputs(235));
    outputs(2088) <= not(layer0_outputs(1680));
    outputs(2089) <= not(layer0_outputs(1565));
    outputs(2090) <= (layer0_outputs(144)) xor (layer0_outputs(2442));
    outputs(2091) <= not(layer0_outputs(340)) or (layer0_outputs(905));
    outputs(2092) <= not(layer0_outputs(362)) or (layer0_outputs(678));
    outputs(2093) <= layer0_outputs(244);
    outputs(2094) <= layer0_outputs(204);
    outputs(2095) <= not(layer0_outputs(1879)) or (layer0_outputs(1985));
    outputs(2096) <= layer0_outputs(1525);
    outputs(2097) <= (layer0_outputs(1391)) xor (layer0_outputs(1320));
    outputs(2098) <= not((layer0_outputs(2303)) xor (layer0_outputs(1705)));
    outputs(2099) <= layer0_outputs(599);
    outputs(2100) <= not(layer0_outputs(1850));
    outputs(2101) <= layer0_outputs(760);
    outputs(2102) <= not(layer0_outputs(1630));
    outputs(2103) <= not(layer0_outputs(1356));
    outputs(2104) <= (layer0_outputs(663)) and not (layer0_outputs(32));
    outputs(2105) <= (layer0_outputs(303)) and (layer0_outputs(1777));
    outputs(2106) <= not((layer0_outputs(1055)) xor (layer0_outputs(721)));
    outputs(2107) <= not(layer0_outputs(743));
    outputs(2108) <= not(layer0_outputs(1631));
    outputs(2109) <= (layer0_outputs(1218)) and not (layer0_outputs(589));
    outputs(2110) <= (layer0_outputs(491)) and not (layer0_outputs(499));
    outputs(2111) <= not(layer0_outputs(1020));
    outputs(2112) <= not(layer0_outputs(157));
    outputs(2113) <= (layer0_outputs(1571)) or (layer0_outputs(2405));
    outputs(2114) <= layer0_outputs(2163);
    outputs(2115) <= layer0_outputs(2508);
    outputs(2116) <= layer0_outputs(853);
    outputs(2117) <= not(layer0_outputs(2371));
    outputs(2118) <= (layer0_outputs(1635)) and (layer0_outputs(1515));
    outputs(2119) <= layer0_outputs(1744);
    outputs(2120) <= layer0_outputs(326);
    outputs(2121) <= not((layer0_outputs(2389)) and (layer0_outputs(2471)));
    outputs(2122) <= layer0_outputs(490);
    outputs(2123) <= not(layer0_outputs(2103)) or (layer0_outputs(796));
    outputs(2124) <= (layer0_outputs(1912)) and not (layer0_outputs(965));
    outputs(2125) <= not(layer0_outputs(1764));
    outputs(2126) <= layer0_outputs(612);
    outputs(2127) <= layer0_outputs(867);
    outputs(2128) <= not((layer0_outputs(1326)) xor (layer0_outputs(1396)));
    outputs(2129) <= layer0_outputs(2410);
    outputs(2130) <= layer0_outputs(2420);
    outputs(2131) <= layer0_outputs(1941);
    outputs(2132) <= (layer0_outputs(2093)) and (layer0_outputs(1744));
    outputs(2133) <= layer0_outputs(1658);
    outputs(2134) <= not((layer0_outputs(2474)) or (layer0_outputs(1249)));
    outputs(2135) <= layer0_outputs(1476);
    outputs(2136) <= not(layer0_outputs(2278)) or (layer0_outputs(40));
    outputs(2137) <= (layer0_outputs(1333)) xor (layer0_outputs(2107));
    outputs(2138) <= (layer0_outputs(308)) and not (layer0_outputs(1386));
    outputs(2139) <= not(layer0_outputs(1971)) or (layer0_outputs(454));
    outputs(2140) <= not((layer0_outputs(992)) or (layer0_outputs(2146)));
    outputs(2141) <= not((layer0_outputs(263)) or (layer0_outputs(1655)));
    outputs(2142) <= not(layer0_outputs(1501));
    outputs(2143) <= not(layer0_outputs(558));
    outputs(2144) <= not((layer0_outputs(906)) or (layer0_outputs(445)));
    outputs(2145) <= layer0_outputs(1543);
    outputs(2146) <= (layer0_outputs(2050)) or (layer0_outputs(686));
    outputs(2147) <= not(layer0_outputs(2417));
    outputs(2148) <= (layer0_outputs(2033)) or (layer0_outputs(1409));
    outputs(2149) <= (layer0_outputs(2518)) and (layer0_outputs(1658));
    outputs(2150) <= not(layer0_outputs(1483));
    outputs(2151) <= (layer0_outputs(332)) and not (layer0_outputs(1727));
    outputs(2152) <= (layer0_outputs(2302)) and not (layer0_outputs(1653));
    outputs(2153) <= layer0_outputs(184);
    outputs(2154) <= layer0_outputs(2367);
    outputs(2155) <= (layer0_outputs(80)) and not (layer0_outputs(893));
    outputs(2156) <= layer0_outputs(2231);
    outputs(2157) <= not(layer0_outputs(1347));
    outputs(2158) <= (layer0_outputs(974)) and (layer0_outputs(760));
    outputs(2159) <= not(layer0_outputs(1981)) or (layer0_outputs(1632));
    outputs(2160) <= layer0_outputs(2213);
    outputs(2161) <= (layer0_outputs(1085)) and not (layer0_outputs(100));
    outputs(2162) <= not((layer0_outputs(359)) and (layer0_outputs(2027)));
    outputs(2163) <= not(layer0_outputs(550));
    outputs(2164) <= layer0_outputs(171);
    outputs(2165) <= (layer0_outputs(1807)) and (layer0_outputs(274));
    outputs(2166) <= not(layer0_outputs(2069)) or (layer0_outputs(1108));
    outputs(2167) <= not(layer0_outputs(865)) or (layer0_outputs(419));
    outputs(2168) <= (layer0_outputs(1723)) and (layer0_outputs(1602));
    outputs(2169) <= not((layer0_outputs(1795)) xor (layer0_outputs(2518)));
    outputs(2170) <= not((layer0_outputs(38)) or (layer0_outputs(516)));
    outputs(2171) <= (layer0_outputs(331)) and not (layer0_outputs(675));
    outputs(2172) <= layer0_outputs(978);
    outputs(2173) <= not((layer0_outputs(2145)) xor (layer0_outputs(1477)));
    outputs(2174) <= not((layer0_outputs(2521)) xor (layer0_outputs(131)));
    outputs(2175) <= not(layer0_outputs(934));
    outputs(2176) <= not(layer0_outputs(313));
    outputs(2177) <= (layer0_outputs(2019)) and (layer0_outputs(201));
    outputs(2178) <= not(layer0_outputs(564));
    outputs(2179) <= not(layer0_outputs(1006));
    outputs(2180) <= layer0_outputs(1757);
    outputs(2181) <= not(layer0_outputs(1750));
    outputs(2182) <= layer0_outputs(1257);
    outputs(2183) <= (layer0_outputs(68)) and not (layer0_outputs(1345));
    outputs(2184) <= not(layer0_outputs(2169)) or (layer0_outputs(1802));
    outputs(2185) <= (layer0_outputs(1447)) and not (layer0_outputs(186));
    outputs(2186) <= layer0_outputs(797);
    outputs(2187) <= not(layer0_outputs(2517));
    outputs(2188) <= not((layer0_outputs(2385)) or (layer0_outputs(1422)));
    outputs(2189) <= layer0_outputs(188);
    outputs(2190) <= not(layer0_outputs(128));
    outputs(2191) <= (layer0_outputs(2070)) and not (layer0_outputs(770));
    outputs(2192) <= not(layer0_outputs(2108));
    outputs(2193) <= not(layer0_outputs(1048));
    outputs(2194) <= layer0_outputs(114);
    outputs(2195) <= layer0_outputs(133);
    outputs(2196) <= layer0_outputs(35);
    outputs(2197) <= layer0_outputs(1784);
    outputs(2198) <= not(layer0_outputs(1732)) or (layer0_outputs(1493));
    outputs(2199) <= not(layer0_outputs(2072));
    outputs(2200) <= layer0_outputs(298);
    outputs(2201) <= layer0_outputs(424);
    outputs(2202) <= (layer0_outputs(612)) and not (layer0_outputs(2091));
    outputs(2203) <= not(layer0_outputs(734));
    outputs(2204) <= not(layer0_outputs(729));
    outputs(2205) <= not(layer0_outputs(2309));
    outputs(2206) <= not(layer0_outputs(310));
    outputs(2207) <= not(layer0_outputs(247));
    outputs(2208) <= not((layer0_outputs(2481)) xor (layer0_outputs(2140)));
    outputs(2209) <= not(layer0_outputs(1129));
    outputs(2210) <= (layer0_outputs(970)) and not (layer0_outputs(1285));
    outputs(2211) <= not((layer0_outputs(723)) or (layer0_outputs(824)));
    outputs(2212) <= (layer0_outputs(2125)) xor (layer0_outputs(2251));
    outputs(2213) <= not(layer0_outputs(2088));
    outputs(2214) <= layer0_outputs(717);
    outputs(2215) <= not(layer0_outputs(1760));
    outputs(2216) <= not(layer0_outputs(1971)) or (layer0_outputs(1305));
    outputs(2217) <= not(layer0_outputs(2534));
    outputs(2218) <= not((layer0_outputs(1449)) xor (layer0_outputs(2341)));
    outputs(2219) <= layer0_outputs(1614);
    outputs(2220) <= (layer0_outputs(767)) and not (layer0_outputs(1088));
    outputs(2221) <= not(layer0_outputs(1633));
    outputs(2222) <= not(layer0_outputs(2006));
    outputs(2223) <= not(layer0_outputs(730));
    outputs(2224) <= layer0_outputs(2237);
    outputs(2225) <= layer0_outputs(1923);
    outputs(2226) <= (layer0_outputs(1902)) and (layer0_outputs(1944));
    outputs(2227) <= not(layer0_outputs(1198)) or (layer0_outputs(1090));
    outputs(2228) <= not(layer0_outputs(583)) or (layer0_outputs(188));
    outputs(2229) <= not(layer0_outputs(1240));
    outputs(2230) <= (layer0_outputs(178)) and (layer0_outputs(2526));
    outputs(2231) <= not((layer0_outputs(855)) xor (layer0_outputs(281)));
    outputs(2232) <= not(layer0_outputs(577));
    outputs(2233) <= not((layer0_outputs(2043)) xor (layer0_outputs(883)));
    outputs(2234) <= (layer0_outputs(449)) or (layer0_outputs(1145));
    outputs(2235) <= not(layer0_outputs(576));
    outputs(2236) <= layer0_outputs(1462);
    outputs(2237) <= (layer0_outputs(1597)) and (layer0_outputs(2093));
    outputs(2238) <= layer0_outputs(2234);
    outputs(2239) <= not(layer0_outputs(2554));
    outputs(2240) <= not(layer0_outputs(503));
    outputs(2241) <= not((layer0_outputs(1720)) xor (layer0_outputs(2530)));
    outputs(2242) <= '1';
    outputs(2243) <= not(layer0_outputs(1397));
    outputs(2244) <= not(layer0_outputs(2049));
    outputs(2245) <= layer0_outputs(323);
    outputs(2246) <= not(layer0_outputs(1121));
    outputs(2247) <= not(layer0_outputs(2240));
    outputs(2248) <= not(layer0_outputs(607));
    outputs(2249) <= (layer0_outputs(602)) and not (layer0_outputs(1565));
    outputs(2250) <= not(layer0_outputs(3));
    outputs(2251) <= (layer0_outputs(2247)) and not (layer0_outputs(818));
    outputs(2252) <= (layer0_outputs(279)) and not (layer0_outputs(2255));
    outputs(2253) <= (layer0_outputs(1445)) and not (layer0_outputs(579));
    outputs(2254) <= (layer0_outputs(1628)) xor (layer0_outputs(1914));
    outputs(2255) <= (layer0_outputs(23)) and not (layer0_outputs(1572));
    outputs(2256) <= not(layer0_outputs(900));
    outputs(2257) <= not(layer0_outputs(2034)) or (layer0_outputs(292));
    outputs(2258) <= layer0_outputs(1341);
    outputs(2259) <= not((layer0_outputs(591)) xor (layer0_outputs(1572)));
    outputs(2260) <= not(layer0_outputs(901)) or (layer0_outputs(113));
    outputs(2261) <= layer0_outputs(452);
    outputs(2262) <= layer0_outputs(565);
    outputs(2263) <= not(layer0_outputs(1557));
    outputs(2264) <= layer0_outputs(872);
    outputs(2265) <= not(layer0_outputs(1595));
    outputs(2266) <= not(layer0_outputs(1297));
    outputs(2267) <= not(layer0_outputs(703));
    outputs(2268) <= (layer0_outputs(665)) and (layer0_outputs(1564));
    outputs(2269) <= not(layer0_outputs(1364));
    outputs(2270) <= layer0_outputs(1672);
    outputs(2271) <= not(layer0_outputs(1505));
    outputs(2272) <= layer0_outputs(1287);
    outputs(2273) <= layer0_outputs(2535);
    outputs(2274) <= not(layer0_outputs(685));
    outputs(2275) <= not((layer0_outputs(838)) and (layer0_outputs(1046)));
    outputs(2276) <= layer0_outputs(406);
    outputs(2277) <= not((layer0_outputs(2250)) xor (layer0_outputs(907)));
    outputs(2278) <= not(layer0_outputs(2015));
    outputs(2279) <= not(layer0_outputs(688));
    outputs(2280) <= not(layer0_outputs(2074));
    outputs(2281) <= (layer0_outputs(200)) and not (layer0_outputs(2));
    outputs(2282) <= not(layer0_outputs(1765)) or (layer0_outputs(590));
    outputs(2283) <= not((layer0_outputs(256)) or (layer0_outputs(1706)));
    outputs(2284) <= not((layer0_outputs(1994)) xor (layer0_outputs(1962)));
    outputs(2285) <= (layer0_outputs(1171)) and not (layer0_outputs(806));
    outputs(2286) <= not((layer0_outputs(2211)) and (layer0_outputs(21)));
    outputs(2287) <= layer0_outputs(828);
    outputs(2288) <= not((layer0_outputs(275)) xor (layer0_outputs(1726)));
    outputs(2289) <= (layer0_outputs(1775)) and not (layer0_outputs(230));
    outputs(2290) <= not(layer0_outputs(1227)) or (layer0_outputs(2068));
    outputs(2291) <= not(layer0_outputs(138));
    outputs(2292) <= not(layer0_outputs(2547));
    outputs(2293) <= (layer0_outputs(7)) xor (layer0_outputs(1039));
    outputs(2294) <= layer0_outputs(1174);
    outputs(2295) <= not(layer0_outputs(1615));
    outputs(2296) <= not((layer0_outputs(2343)) and (layer0_outputs(2142)));
    outputs(2297) <= layer0_outputs(1724);
    outputs(2298) <= not((layer0_outputs(1172)) xor (layer0_outputs(2519)));
    outputs(2299) <= (layer0_outputs(948)) and (layer0_outputs(1723));
    outputs(2300) <= (layer0_outputs(1800)) or (layer0_outputs(1363));
    outputs(2301) <= not((layer0_outputs(1069)) xor (layer0_outputs(1710)));
    outputs(2302) <= not(layer0_outputs(301));
    outputs(2303) <= layer0_outputs(1194);
    outputs(2304) <= not(layer0_outputs(1057));
    outputs(2305) <= layer0_outputs(2190);
    outputs(2306) <= (layer0_outputs(2257)) and not (layer0_outputs(928));
    outputs(2307) <= (layer0_outputs(778)) and (layer0_outputs(994));
    outputs(2308) <= (layer0_outputs(1591)) and (layer0_outputs(2432));
    outputs(2309) <= layer0_outputs(459);
    outputs(2310) <= (layer0_outputs(1398)) and (layer0_outputs(404));
    outputs(2311) <= not(layer0_outputs(830));
    outputs(2312) <= (layer0_outputs(132)) xor (layer0_outputs(759));
    outputs(2313) <= (layer0_outputs(1047)) and (layer0_outputs(2002));
    outputs(2314) <= not(layer0_outputs(223));
    outputs(2315) <= layer0_outputs(1452);
    outputs(2316) <= not(layer0_outputs(1804));
    outputs(2317) <= layer0_outputs(894);
    outputs(2318) <= (layer0_outputs(212)) and not (layer0_outputs(2303));
    outputs(2319) <= (layer0_outputs(2120)) and (layer0_outputs(1258));
    outputs(2320) <= layer0_outputs(881);
    outputs(2321) <= not(layer0_outputs(6));
    outputs(2322) <= layer0_outputs(2207);
    outputs(2323) <= not((layer0_outputs(931)) and (layer0_outputs(2272)));
    outputs(2324) <= (layer0_outputs(1937)) and not (layer0_outputs(1948));
    outputs(2325) <= layer0_outputs(5);
    outputs(2326) <= layer0_outputs(357);
    outputs(2327) <= (layer0_outputs(1897)) and not (layer0_outputs(1135));
    outputs(2328) <= not(layer0_outputs(2507));
    outputs(2329) <= not(layer0_outputs(1860));
    outputs(2330) <= (layer0_outputs(481)) and (layer0_outputs(744));
    outputs(2331) <= not(layer0_outputs(495));
    outputs(2332) <= not(layer0_outputs(1787));
    outputs(2333) <= (layer0_outputs(1186)) and (layer0_outputs(1007));
    outputs(2334) <= not(layer0_outputs(2123));
    outputs(2335) <= not((layer0_outputs(1109)) or (layer0_outputs(1498)));
    outputs(2336) <= (layer0_outputs(1743)) and not (layer0_outputs(895));
    outputs(2337) <= (layer0_outputs(546)) and (layer0_outputs(203));
    outputs(2338) <= (layer0_outputs(246)) and not (layer0_outputs(962));
    outputs(2339) <= not((layer0_outputs(1883)) xor (layer0_outputs(2118)));
    outputs(2340) <= layer0_outputs(1389);
    outputs(2341) <= (layer0_outputs(555)) and not (layer0_outputs(945));
    outputs(2342) <= (layer0_outputs(2525)) and not (layer0_outputs(74));
    outputs(2343) <= (layer0_outputs(1403)) and not (layer0_outputs(868));
    outputs(2344) <= not(layer0_outputs(2099));
    outputs(2345) <= not(layer0_outputs(2391));
    outputs(2346) <= (layer0_outputs(1693)) and not (layer0_outputs(1955));
    outputs(2347) <= not((layer0_outputs(28)) xor (layer0_outputs(2393)));
    outputs(2348) <= (layer0_outputs(444)) and (layer0_outputs(1180));
    outputs(2349) <= not(layer0_outputs(2044));
    outputs(2350) <= (layer0_outputs(1145)) and not (layer0_outputs(245));
    outputs(2351) <= (layer0_outputs(1242)) or (layer0_outputs(2486));
    outputs(2352) <= (layer0_outputs(890)) xor (layer0_outputs(696));
    outputs(2353) <= (layer0_outputs(190)) and not (layer0_outputs(1135));
    outputs(2354) <= (layer0_outputs(2222)) and not (layer0_outputs(694));
    outputs(2355) <= (layer0_outputs(2476)) and not (layer0_outputs(1089));
    outputs(2356) <= not(layer0_outputs(1656));
    outputs(2357) <= not(layer0_outputs(1855));
    outputs(2358) <= layer0_outputs(649);
    outputs(2359) <= layer0_outputs(2495);
    outputs(2360) <= (layer0_outputs(617)) and not (layer0_outputs(223));
    outputs(2361) <= not((layer0_outputs(515)) or (layer0_outputs(1339)));
    outputs(2362) <= not(layer0_outputs(2059));
    outputs(2363) <= (layer0_outputs(282)) and not (layer0_outputs(939));
    outputs(2364) <= not(layer0_outputs(892));
    outputs(2365) <= (layer0_outputs(476)) xor (layer0_outputs(1985));
    outputs(2366) <= not(layer0_outputs(774));
    outputs(2367) <= (layer0_outputs(231)) and (layer0_outputs(2550));
    outputs(2368) <= (layer0_outputs(307)) and not (layer0_outputs(937));
    outputs(2369) <= (layer0_outputs(1299)) and not (layer0_outputs(480));
    outputs(2370) <= (layer0_outputs(269)) and not (layer0_outputs(1100));
    outputs(2371) <= not((layer0_outputs(848)) or (layer0_outputs(576)));
    outputs(2372) <= (layer0_outputs(911)) and not (layer0_outputs(374));
    outputs(2373) <= layer0_outputs(956);
    outputs(2374) <= not(layer0_outputs(396));
    outputs(2375) <= (layer0_outputs(72)) and (layer0_outputs(430));
    outputs(2376) <= (layer0_outputs(1581)) and (layer0_outputs(2222));
    outputs(2377) <= not(layer0_outputs(1357));
    outputs(2378) <= not(layer0_outputs(1553));
    outputs(2379) <= layer0_outputs(2139);
    outputs(2380) <= (layer0_outputs(2446)) and not (layer0_outputs(2244));
    outputs(2381) <= layer0_outputs(252);
    outputs(2382) <= not(layer0_outputs(1947));
    outputs(2383) <= (layer0_outputs(2179)) and (layer0_outputs(2062));
    outputs(2384) <= not(layer0_outputs(2119));
    outputs(2385) <= not((layer0_outputs(301)) or (layer0_outputs(1776)));
    outputs(2386) <= not((layer0_outputs(839)) or (layer0_outputs(1611)));
    outputs(2387) <= (layer0_outputs(1929)) and not (layer0_outputs(1811));
    outputs(2388) <= not(layer0_outputs(510));
    outputs(2389) <= not((layer0_outputs(524)) or (layer0_outputs(264)));
    outputs(2390) <= (layer0_outputs(274)) and (layer0_outputs(1826));
    outputs(2391) <= (layer0_outputs(502)) and not (layer0_outputs(225));
    outputs(2392) <= not((layer0_outputs(2487)) or (layer0_outputs(573)));
    outputs(2393) <= not(layer0_outputs(523));
    outputs(2394) <= not(layer0_outputs(98));
    outputs(2395) <= (layer0_outputs(2004)) and not (layer0_outputs(1829));
    outputs(2396) <= (layer0_outputs(1596)) and not (layer0_outputs(2420));
    outputs(2397) <= not(layer0_outputs(1747)) or (layer0_outputs(1641));
    outputs(2398) <= (layer0_outputs(2231)) and not (layer0_outputs(437));
    outputs(2399) <= layer0_outputs(2011);
    outputs(2400) <= (layer0_outputs(401)) and not (layer0_outputs(1423));
    outputs(2401) <= layer0_outputs(1720);
    outputs(2402) <= layer0_outputs(1488);
    outputs(2403) <= layer0_outputs(2226);
    outputs(2404) <= layer0_outputs(572);
    outputs(2405) <= not(layer0_outputs(1670));
    outputs(2406) <= (layer0_outputs(747)) xor (layer0_outputs(1639));
    outputs(2407) <= (layer0_outputs(755)) and not (layer0_outputs(643));
    outputs(2408) <= not(layer0_outputs(2385));
    outputs(2409) <= (layer0_outputs(496)) and (layer0_outputs(1177));
    outputs(2410) <= not(layer0_outputs(1598));
    outputs(2411) <= not(layer0_outputs(153));
    outputs(2412) <= not(layer0_outputs(1598));
    outputs(2413) <= not(layer0_outputs(877));
    outputs(2414) <= (layer0_outputs(1526)) xor (layer0_outputs(2493));
    outputs(2415) <= layer0_outputs(923);
    outputs(2416) <= (layer0_outputs(1387)) and not (layer0_outputs(2006));
    outputs(2417) <= not(layer0_outputs(2293));
    outputs(2418) <= not((layer0_outputs(1307)) or (layer0_outputs(1356)));
    outputs(2419) <= not(layer0_outputs(1839)) or (layer0_outputs(1383));
    outputs(2420) <= (layer0_outputs(642)) and (layer0_outputs(2013));
    outputs(2421) <= not((layer0_outputs(1406)) and (layer0_outputs(47)));
    outputs(2422) <= (layer0_outputs(1123)) and (layer0_outputs(1984));
    outputs(2423) <= (layer0_outputs(1806)) and not (layer0_outputs(2298));
    outputs(2424) <= layer0_outputs(707);
    outputs(2425) <= (layer0_outputs(2396)) and (layer0_outputs(1092));
    outputs(2426) <= layer0_outputs(2536);
    outputs(2427) <= (layer0_outputs(1023)) xor (layer0_outputs(1300));
    outputs(2428) <= (layer0_outputs(623)) and not (layer0_outputs(2266));
    outputs(2429) <= layer0_outputs(130);
    outputs(2430) <= not((layer0_outputs(1437)) or (layer0_outputs(2397)));
    outputs(2431) <= (layer0_outputs(1524)) and (layer0_outputs(772));
    outputs(2432) <= layer0_outputs(1334);
    outputs(2433) <= not((layer0_outputs(199)) or (layer0_outputs(1076)));
    outputs(2434) <= layer0_outputs(1313);
    outputs(2435) <= not(layer0_outputs(1141));
    outputs(2436) <= not((layer0_outputs(2484)) or (layer0_outputs(522)));
    outputs(2437) <= (layer0_outputs(1911)) and not (layer0_outputs(1138));
    outputs(2438) <= not((layer0_outputs(2158)) or (layer0_outputs(971)));
    outputs(2439) <= (layer0_outputs(755)) and (layer0_outputs(1725));
    outputs(2440) <= (layer0_outputs(1748)) and (layer0_outputs(1793));
    outputs(2441) <= not((layer0_outputs(2136)) or (layer0_outputs(784)));
    outputs(2442) <= not(layer0_outputs(2038));
    outputs(2443) <= (layer0_outputs(1087)) and not (layer0_outputs(1885));
    outputs(2444) <= layer0_outputs(384);
    outputs(2445) <= not(layer0_outputs(924));
    outputs(2446) <= layer0_outputs(1045);
    outputs(2447) <= (layer0_outputs(1739)) and (layer0_outputs(365));
    outputs(2448) <= not((layer0_outputs(811)) and (layer0_outputs(2191)));
    outputs(2449) <= layer0_outputs(2366);
    outputs(2450) <= layer0_outputs(1724);
    outputs(2451) <= (layer0_outputs(1387)) and not (layer0_outputs(103));
    outputs(2452) <= not(layer0_outputs(1551));
    outputs(2453) <= (layer0_outputs(205)) and not (layer0_outputs(1237));
    outputs(2454) <= not(layer0_outputs(710));
    outputs(2455) <= (layer0_outputs(244)) xor (layer0_outputs(1953));
    outputs(2456) <= not(layer0_outputs(2134));
    outputs(2457) <= layer0_outputs(1734);
    outputs(2458) <= (layer0_outputs(328)) and not (layer0_outputs(753));
    outputs(2459) <= not(layer0_outputs(2314));
    outputs(2460) <= not((layer0_outputs(2430)) or (layer0_outputs(1613)));
    outputs(2461) <= not(layer0_outputs(914));
    outputs(2462) <= (layer0_outputs(952)) and not (layer0_outputs(1325));
    outputs(2463) <= layer0_outputs(104);
    outputs(2464) <= layer0_outputs(1485);
    outputs(2465) <= layer0_outputs(1871);
    outputs(2466) <= layer0_outputs(1077);
    outputs(2467) <= not(layer0_outputs(408));
    outputs(2468) <= (layer0_outputs(936)) and not (layer0_outputs(2383));
    outputs(2469) <= not((layer0_outputs(1808)) or (layer0_outputs(53)));
    outputs(2470) <= layer0_outputs(866);
    outputs(2471) <= layer0_outputs(801);
    outputs(2472) <= (layer0_outputs(1245)) and not (layer0_outputs(2354));
    outputs(2473) <= (layer0_outputs(1052)) and (layer0_outputs(395));
    outputs(2474) <= layer0_outputs(1516);
    outputs(2475) <= not(layer0_outputs(2126));
    outputs(2476) <= (layer0_outputs(1916)) and not (layer0_outputs(945));
    outputs(2477) <= not((layer0_outputs(1389)) xor (layer0_outputs(1160)));
    outputs(2478) <= layer0_outputs(813);
    outputs(2479) <= (layer0_outputs(2080)) xor (layer0_outputs(1412));
    outputs(2480) <= layer0_outputs(494);
    outputs(2481) <= not(layer0_outputs(1553));
    outputs(2482) <= layer0_outputs(2011);
    outputs(2483) <= not((layer0_outputs(1000)) or (layer0_outputs(808)));
    outputs(2484) <= (layer0_outputs(884)) and not (layer0_outputs(487));
    outputs(2485) <= layer0_outputs(2193);
    outputs(2486) <= layer0_outputs(1700);
    outputs(2487) <= not(layer0_outputs(1665)) or (layer0_outputs(409));
    outputs(2488) <= not(layer0_outputs(263));
    outputs(2489) <= layer0_outputs(195);
    outputs(2490) <= (layer0_outputs(952)) and not (layer0_outputs(1107));
    outputs(2491) <= not((layer0_outputs(1500)) or (layer0_outputs(1495)));
    outputs(2492) <= layer0_outputs(496);
    outputs(2493) <= not(layer0_outputs(526)) or (layer0_outputs(574));
    outputs(2494) <= layer0_outputs(2040);
    outputs(2495) <= layer0_outputs(2276);
    outputs(2496) <= (layer0_outputs(681)) and (layer0_outputs(921));
    outputs(2497) <= not(layer0_outputs(1255));
    outputs(2498) <= layer0_outputs(544);
    outputs(2499) <= (layer0_outputs(1718)) and not (layer0_outputs(853));
    outputs(2500) <= (layer0_outputs(559)) and not (layer0_outputs(181));
    outputs(2501) <= layer0_outputs(2304);
    outputs(2502) <= not(layer0_outputs(1551));
    outputs(2503) <= not((layer0_outputs(1209)) or (layer0_outputs(816)));
    outputs(2504) <= not((layer0_outputs(690)) or (layer0_outputs(1964)));
    outputs(2505) <= not(layer0_outputs(2402));
    outputs(2506) <= layer0_outputs(1766);
    outputs(2507) <= not(layer0_outputs(584));
    outputs(2508) <= layer0_outputs(101);
    outputs(2509) <= not(layer0_outputs(914)) or (layer0_outputs(902));
    outputs(2510) <= not((layer0_outputs(2001)) or (layer0_outputs(509)));
    outputs(2511) <= not(layer0_outputs(155));
    outputs(2512) <= (layer0_outputs(1719)) and (layer0_outputs(1201));
    outputs(2513) <= (layer0_outputs(789)) and not (layer0_outputs(319));
    outputs(2514) <= not((layer0_outputs(2152)) xor (layer0_outputs(1794)));
    outputs(2515) <= not(layer0_outputs(1448));
    outputs(2516) <= (layer0_outputs(1668)) and not (layer0_outputs(1957));
    outputs(2517) <= not((layer0_outputs(816)) or (layer0_outputs(1090)));
    outputs(2518) <= (layer0_outputs(2332)) xor (layer0_outputs(1606));
    outputs(2519) <= layer0_outputs(978);
    outputs(2520) <= (layer0_outputs(1952)) and not (layer0_outputs(1056));
    outputs(2521) <= (layer0_outputs(1871)) and (layer0_outputs(1663));
    outputs(2522) <= not((layer0_outputs(1402)) xor (layer0_outputs(56)));
    outputs(2523) <= not((layer0_outputs(2461)) or (layer0_outputs(1844)));
    outputs(2524) <= (layer0_outputs(1965)) and not (layer0_outputs(2547));
    outputs(2525) <= layer0_outputs(754);
    outputs(2526) <= layer0_outputs(1294);
    outputs(2527) <= layer0_outputs(1542);
    outputs(2528) <= (layer0_outputs(769)) and not (layer0_outputs(2173));
    outputs(2529) <= (layer0_outputs(353)) and (layer0_outputs(61));
    outputs(2530) <= not(layer0_outputs(48));
    outputs(2531) <= (layer0_outputs(2474)) xor (layer0_outputs(2517));
    outputs(2532) <= not(layer0_outputs(915));
    outputs(2533) <= (layer0_outputs(1317)) xor (layer0_outputs(1710));
    outputs(2534) <= (layer0_outputs(1299)) and not (layer0_outputs(516));
    outputs(2535) <= (layer0_outputs(2249)) and (layer0_outputs(772));
    outputs(2536) <= (layer0_outputs(1873)) and not (layer0_outputs(964));
    outputs(2537) <= layer0_outputs(666);
    outputs(2538) <= not(layer0_outputs(2289));
    outputs(2539) <= (layer0_outputs(719)) and (layer0_outputs(1912));
    outputs(2540) <= (layer0_outputs(2236)) and not (layer0_outputs(255));
    outputs(2541) <= layer0_outputs(609);
    outputs(2542) <= (layer0_outputs(1753)) and not (layer0_outputs(220));
    outputs(2543) <= layer0_outputs(2529);
    outputs(2544) <= (layer0_outputs(1661)) and not (layer0_outputs(276));
    outputs(2545) <= not((layer0_outputs(1754)) or (layer0_outputs(2515)));
    outputs(2546) <= not((layer0_outputs(1508)) or (layer0_outputs(2000)));
    outputs(2547) <= (layer0_outputs(345)) and not (layer0_outputs(938));
    outputs(2548) <= (layer0_outputs(822)) and (layer0_outputs(2439));
    outputs(2549) <= not(layer0_outputs(280));
    outputs(2550) <= layer0_outputs(2277);
    outputs(2551) <= not(layer0_outputs(114));
    outputs(2552) <= not(layer0_outputs(1652));
    outputs(2553) <= not(layer0_outputs(2326));
    outputs(2554) <= (layer0_outputs(1084)) and (layer0_outputs(735));
    outputs(2555) <= not(layer0_outputs(1271));
    outputs(2556) <= layer0_outputs(1708);
    outputs(2557) <= layer0_outputs(1154);
    outputs(2558) <= not((layer0_outputs(1607)) or (layer0_outputs(180)));
    outputs(2559) <= not((layer0_outputs(376)) and (layer0_outputs(803)));

end Behavioral;
