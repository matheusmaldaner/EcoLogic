module logic_network(
    input wire [255:0] inputs,
    output wire [9:0] outputs
);

    wire [5119:0] layer0_outputs;
    wire [5119:0] layer1_outputs;
    wire [5119:0] layer2_outputs;
    wire [5119:0] layer3_outputs;
    wire [5119:0] layer4_outputs;
    wire [5119:0] layer5_outputs;
    wire [5119:0] layer6_outputs;

    assign layer0_outputs[0] = ~(inputs[3]) | (inputs[95]);
    assign layer0_outputs[1] = 1'b0;
    assign layer0_outputs[2] = (inputs[246]) & ~(inputs[173]);
    assign layer0_outputs[3] = inputs[56];
    assign layer0_outputs[4] = (inputs[44]) & ~(inputs[231]);
    assign layer0_outputs[5] = ~((inputs[191]) | (inputs[115]));
    assign layer0_outputs[6] = inputs[94];
    assign layer0_outputs[7] = inputs[112];
    assign layer0_outputs[8] = ~(inputs[215]) | (inputs[26]);
    assign layer0_outputs[9] = ~((inputs[20]) | (inputs[102]));
    assign layer0_outputs[10] = (inputs[178]) | (inputs[153]);
    assign layer0_outputs[11] = ~(inputs[46]) | (inputs[155]);
    assign layer0_outputs[12] = 1'b0;
    assign layer0_outputs[13] = inputs[78];
    assign layer0_outputs[14] = (inputs[47]) & ~(inputs[81]);
    assign layer0_outputs[15] = ~(inputs[108]);
    assign layer0_outputs[16] = (inputs[42]) & ~(inputs[235]);
    assign layer0_outputs[17] = (inputs[32]) & (inputs[171]);
    assign layer0_outputs[18] = (inputs[190]) & ~(inputs[170]);
    assign layer0_outputs[19] = (inputs[13]) & ~(inputs[146]);
    assign layer0_outputs[20] = ~((inputs[127]) | (inputs[95]));
    assign layer0_outputs[21] = ~(inputs[110]) | (inputs[84]);
    assign layer0_outputs[22] = inputs[138];
    assign layer0_outputs[23] = (inputs[236]) & ~(inputs[180]);
    assign layer0_outputs[24] = (inputs[18]) & ~(inputs[60]);
    assign layer0_outputs[25] = inputs[216];
    assign layer0_outputs[26] = 1'b1;
    assign layer0_outputs[27] = ~(inputs[136]) | (inputs[154]);
    assign layer0_outputs[28] = (inputs[77]) & ~(inputs[19]);
    assign layer0_outputs[29] = inputs[76];
    assign layer0_outputs[30] = (inputs[231]) ^ (inputs[15]);
    assign layer0_outputs[31] = ~((inputs[41]) ^ (inputs[8]));
    assign layer0_outputs[32] = 1'b1;
    assign layer0_outputs[33] = (inputs[6]) & ~(inputs[50]);
    assign layer0_outputs[34] = ~((inputs[173]) & (inputs[58]));
    assign layer0_outputs[35] = inputs[47];
    assign layer0_outputs[36] = (inputs[126]) & (inputs[186]);
    assign layer0_outputs[37] = ~((inputs[204]) & (inputs[107]));
    assign layer0_outputs[38] = (inputs[235]) & (inputs[66]);
    assign layer0_outputs[39] = inputs[156];
    assign layer0_outputs[40] = ~((inputs[43]) | (inputs[102]));
    assign layer0_outputs[41] = (inputs[162]) & ~(inputs[66]);
    assign layer0_outputs[42] = (inputs[198]) & (inputs[200]);
    assign layer0_outputs[43] = (inputs[89]) & ~(inputs[254]);
    assign layer0_outputs[44] = 1'b0;
    assign layer0_outputs[45] = ~((inputs[206]) & (inputs[193]));
    assign layer0_outputs[46] = (inputs[128]) & ~(inputs[42]);
    assign layer0_outputs[47] = ~((inputs[239]) | (inputs[187]));
    assign layer0_outputs[48] = ~(inputs[248]);
    assign layer0_outputs[49] = (inputs[170]) | (inputs[42]);
    assign layer0_outputs[50] = ~(inputs[71]);
    assign layer0_outputs[51] = ~(inputs[153]) | (inputs[199]);
    assign layer0_outputs[52] = inputs[57];
    assign layer0_outputs[53] = (inputs[184]) | (inputs[24]);
    assign layer0_outputs[54] = ~(inputs[207]) | (inputs[34]);
    assign layer0_outputs[55] = (inputs[10]) ^ (inputs[12]);
    assign layer0_outputs[56] = (inputs[169]) & ~(inputs[178]);
    assign layer0_outputs[57] = ~(inputs[162]);
    assign layer0_outputs[58] = inputs[7];
    assign layer0_outputs[59] = ~((inputs[111]) ^ (inputs[178]));
    assign layer0_outputs[60] = inputs[153];
    assign layer0_outputs[61] = (inputs[44]) & ~(inputs[95]);
    assign layer0_outputs[62] = (inputs[161]) & (inputs[243]);
    assign layer0_outputs[63] = inputs[8];
    assign layer0_outputs[64] = ~(inputs[177]);
    assign layer0_outputs[65] = (inputs[192]) & (inputs[80]);
    assign layer0_outputs[66] = (inputs[54]) ^ (inputs[207]);
    assign layer0_outputs[67] = ~((inputs[39]) ^ (inputs[144]));
    assign layer0_outputs[68] = ~((inputs[75]) | (inputs[16]));
    assign layer0_outputs[69] = (inputs[111]) | (inputs[116]);
    assign layer0_outputs[70] = ~(inputs[113]);
    assign layer0_outputs[71] = 1'b1;
    assign layer0_outputs[72] = ~((inputs[98]) ^ (inputs[65]));
    assign layer0_outputs[73] = ~((inputs[148]) & (inputs[152]));
    assign layer0_outputs[74] = inputs[222];
    assign layer0_outputs[75] = ~(inputs[96]);
    assign layer0_outputs[76] = inputs[124];
    assign layer0_outputs[77] = (inputs[51]) & ~(inputs[247]);
    assign layer0_outputs[78] = (inputs[16]) & ~(inputs[196]);
    assign layer0_outputs[79] = ~(inputs[167]);
    assign layer0_outputs[80] = inputs[186];
    assign layer0_outputs[81] = inputs[57];
    assign layer0_outputs[82] = ~((inputs[190]) ^ (inputs[30]));
    assign layer0_outputs[83] = ~(inputs[60]) | (inputs[28]);
    assign layer0_outputs[84] = ~(inputs[149]);
    assign layer0_outputs[85] = ~((inputs[11]) ^ (inputs[3]));
    assign layer0_outputs[86] = ~(inputs[156]);
    assign layer0_outputs[87] = ~(inputs[106]);
    assign layer0_outputs[88] = (inputs[120]) & (inputs[56]);
    assign layer0_outputs[89] = 1'b0;
    assign layer0_outputs[90] = inputs[51];
    assign layer0_outputs[91] = 1'b1;
    assign layer0_outputs[92] = 1'b1;
    assign layer0_outputs[93] = 1'b1;
    assign layer0_outputs[94] = ~(inputs[188]) | (inputs[254]);
    assign layer0_outputs[95] = ~(inputs[160]);
    assign layer0_outputs[96] = (inputs[178]) ^ (inputs[133]);
    assign layer0_outputs[97] = inputs[219];
    assign layer0_outputs[98] = (inputs[149]) & ~(inputs[29]);
    assign layer0_outputs[99] = ~((inputs[101]) | (inputs[47]));
    assign layer0_outputs[100] = (inputs[200]) | (inputs[233]);
    assign layer0_outputs[101] = ~(inputs[168]) | (inputs[121]);
    assign layer0_outputs[102] = inputs[6];
    assign layer0_outputs[103] = ~(inputs[8]) | (inputs[43]);
    assign layer0_outputs[104] = ~((inputs[163]) & (inputs[54]));
    assign layer0_outputs[105] = inputs[197];
    assign layer0_outputs[106] = 1'b0;
    assign layer0_outputs[107] = ~((inputs[176]) ^ (inputs[239]));
    assign layer0_outputs[108] = inputs[13];
    assign layer0_outputs[109] = (inputs[68]) & ~(inputs[42]);
    assign layer0_outputs[110] = (inputs[245]) & ~(inputs[255]);
    assign layer0_outputs[111] = ~((inputs[115]) & (inputs[140]));
    assign layer0_outputs[112] = (inputs[175]) & ~(inputs[83]);
    assign layer0_outputs[113] = (inputs[97]) | (inputs[130]);
    assign layer0_outputs[114] = (inputs[24]) & (inputs[60]);
    assign layer0_outputs[115] = ~(inputs[164]);
    assign layer0_outputs[116] = (inputs[214]) | (inputs[198]);
    assign layer0_outputs[117] = (inputs[4]) & ~(inputs[42]);
    assign layer0_outputs[118] = inputs[214];
    assign layer0_outputs[119] = (inputs[171]) | (inputs[56]);
    assign layer0_outputs[120] = (inputs[157]) & ~(inputs[96]);
    assign layer0_outputs[121] = ~(inputs[173]);
    assign layer0_outputs[122] = 1'b0;
    assign layer0_outputs[123] = ~(inputs[176]) | (inputs[124]);
    assign layer0_outputs[124] = ~(inputs[129]) | (inputs[230]);
    assign layer0_outputs[125] = ~(inputs[156]) | (inputs[23]);
    assign layer0_outputs[126] = (inputs[55]) & (inputs[49]);
    assign layer0_outputs[127] = (inputs[200]) | (inputs[241]);
    assign layer0_outputs[128] = (inputs[178]) & ~(inputs[106]);
    assign layer0_outputs[129] = inputs[74];
    assign layer0_outputs[130] = ~(inputs[90]);
    assign layer0_outputs[131] = ~((inputs[25]) | (inputs[123]));
    assign layer0_outputs[132] = ~(inputs[157]);
    assign layer0_outputs[133] = ~((inputs[253]) ^ (inputs[162]));
    assign layer0_outputs[134] = ~(inputs[169]) | (inputs[17]);
    assign layer0_outputs[135] = 1'b0;
    assign layer0_outputs[136] = inputs[174];
    assign layer0_outputs[137] = 1'b1;
    assign layer0_outputs[138] = (inputs[178]) & ~(inputs[166]);
    assign layer0_outputs[139] = ~(inputs[64]) | (inputs[252]);
    assign layer0_outputs[140] = ~((inputs[214]) | (inputs[103]));
    assign layer0_outputs[141] = (inputs[189]) | (inputs[134]);
    assign layer0_outputs[142] = (inputs[110]) | (inputs[253]);
    assign layer0_outputs[143] = inputs[160];
    assign layer0_outputs[144] = ~((inputs[156]) & (inputs[29]));
    assign layer0_outputs[145] = ~(inputs[191]);
    assign layer0_outputs[146] = inputs[187];
    assign layer0_outputs[147] = ~(inputs[78]);
    assign layer0_outputs[148] = inputs[111];
    assign layer0_outputs[149] = (inputs[194]) | (inputs[164]);
    assign layer0_outputs[150] = ~((inputs[47]) ^ (inputs[55]));
    assign layer0_outputs[151] = inputs[76];
    assign layer0_outputs[152] = inputs[203];
    assign layer0_outputs[153] = ~(inputs[68]);
    assign layer0_outputs[154] = ~((inputs[93]) | (inputs[149]));
    assign layer0_outputs[155] = (inputs[180]) | (inputs[55]);
    assign layer0_outputs[156] = 1'b1;
    assign layer0_outputs[157] = ~((inputs[233]) | (inputs[250]));
    assign layer0_outputs[158] = ~(inputs[249]);
    assign layer0_outputs[159] = (inputs[188]) | (inputs[40]);
    assign layer0_outputs[160] = (inputs[33]) & (inputs[174]);
    assign layer0_outputs[161] = 1'b0;
    assign layer0_outputs[162] = 1'b0;
    assign layer0_outputs[163] = (inputs[99]) & ~(inputs[135]);
    assign layer0_outputs[164] = inputs[74];
    assign layer0_outputs[165] = 1'b0;
    assign layer0_outputs[166] = ~(inputs[29]) | (inputs[84]);
    assign layer0_outputs[167] = (inputs[37]) & ~(inputs[148]);
    assign layer0_outputs[168] = (inputs[192]) | (inputs[254]);
    assign layer0_outputs[169] = (inputs[28]) & ~(inputs[28]);
    assign layer0_outputs[170] = ~(inputs[93]) | (inputs[31]);
    assign layer0_outputs[171] = 1'b1;
    assign layer0_outputs[172] = inputs[156];
    assign layer0_outputs[173] = (inputs[125]) ^ (inputs[6]);
    assign layer0_outputs[174] = ~((inputs[106]) ^ (inputs[2]));
    assign layer0_outputs[175] = ~((inputs[243]) & (inputs[47]));
    assign layer0_outputs[176] = 1'b0;
    assign layer0_outputs[177] = 1'b0;
    assign layer0_outputs[178] = ~(inputs[110]);
    assign layer0_outputs[179] = (inputs[20]) | (inputs[56]);
    assign layer0_outputs[180] = 1'b0;
    assign layer0_outputs[181] = (inputs[40]) & ~(inputs[119]);
    assign layer0_outputs[182] = ~(inputs[197]);
    assign layer0_outputs[183] = 1'b0;
    assign layer0_outputs[184] = ~((inputs[161]) | (inputs[30]));
    assign layer0_outputs[185] = ~((inputs[70]) ^ (inputs[16]));
    assign layer0_outputs[186] = ~(inputs[63]) | (inputs[203]);
    assign layer0_outputs[187] = inputs[41];
    assign layer0_outputs[188] = ~(inputs[0]);
    assign layer0_outputs[189] = ~((inputs[175]) ^ (inputs[251]));
    assign layer0_outputs[190] = ~(inputs[111]);
    assign layer0_outputs[191] = ~((inputs[121]) | (inputs[16]));
    assign layer0_outputs[192] = ~((inputs[109]) & (inputs[35]));
    assign layer0_outputs[193] = (inputs[76]) & ~(inputs[195]);
    assign layer0_outputs[194] = ~(inputs[199]);
    assign layer0_outputs[195] = (inputs[236]) & (inputs[38]);
    assign layer0_outputs[196] = inputs[247];
    assign layer0_outputs[197] = ~(inputs[118]);
    assign layer0_outputs[198] = ~((inputs[59]) | (inputs[182]));
    assign layer0_outputs[199] = (inputs[139]) | (inputs[129]);
    assign layer0_outputs[200] = inputs[66];
    assign layer0_outputs[201] = ~(inputs[126]);
    assign layer0_outputs[202] = (inputs[226]) & ~(inputs[136]);
    assign layer0_outputs[203] = (inputs[129]) & ~(inputs[189]);
    assign layer0_outputs[204] = (inputs[192]) & ~(inputs[53]);
    assign layer0_outputs[205] = inputs[89];
    assign layer0_outputs[206] = ~((inputs[141]) ^ (inputs[231]));
    assign layer0_outputs[207] = ~((inputs[218]) ^ (inputs[94]));
    assign layer0_outputs[208] = (inputs[188]) & ~(inputs[219]);
    assign layer0_outputs[209] = (inputs[53]) | (inputs[236]);
    assign layer0_outputs[210] = ~(inputs[230]);
    assign layer0_outputs[211] = (inputs[197]) & ~(inputs[252]);
    assign layer0_outputs[212] = inputs[52];
    assign layer0_outputs[213] = (inputs[25]) | (inputs[142]);
    assign layer0_outputs[214] = (inputs[107]) & ~(inputs[170]);
    assign layer0_outputs[215] = ~((inputs[13]) | (inputs[87]));
    assign layer0_outputs[216] = inputs[67];
    assign layer0_outputs[217] = ~(inputs[137]);
    assign layer0_outputs[218] = (inputs[93]) | (inputs[42]);
    assign layer0_outputs[219] = ~(inputs[180]) | (inputs[186]);
    assign layer0_outputs[220] = ~((inputs[75]) & (inputs[19]));
    assign layer0_outputs[221] = (inputs[135]) & ~(inputs[54]);
    assign layer0_outputs[222] = (inputs[22]) & (inputs[254]);
    assign layer0_outputs[223] = inputs[31];
    assign layer0_outputs[224] = inputs[113];
    assign layer0_outputs[225] = ~((inputs[219]) | (inputs[51]));
    assign layer0_outputs[226] = (inputs[63]) | (inputs[17]);
    assign layer0_outputs[227] = ~(inputs[0]);
    assign layer0_outputs[228] = ~((inputs[240]) & (inputs[44]));
    assign layer0_outputs[229] = (inputs[235]) ^ (inputs[45]);
    assign layer0_outputs[230] = (inputs[238]) & ~(inputs[202]);
    assign layer0_outputs[231] = ~((inputs[81]) & (inputs[226]));
    assign layer0_outputs[232] = ~((inputs[175]) ^ (inputs[64]));
    assign layer0_outputs[233] = ~(inputs[28]);
    assign layer0_outputs[234] = ~(inputs[73]);
    assign layer0_outputs[235] = 1'b1;
    assign layer0_outputs[236] = inputs[117];
    assign layer0_outputs[237] = (inputs[144]) | (inputs[63]);
    assign layer0_outputs[238] = inputs[240];
    assign layer0_outputs[239] = ~(inputs[89]);
    assign layer0_outputs[240] = ~(inputs[191]) | (inputs[130]);
    assign layer0_outputs[241] = 1'b0;
    assign layer0_outputs[242] = inputs[178];
    assign layer0_outputs[243] = (inputs[242]) & ~(inputs[233]);
    assign layer0_outputs[244] = ~(inputs[59]) | (inputs[28]);
    assign layer0_outputs[245] = ~((inputs[250]) ^ (inputs[68]));
    assign layer0_outputs[246] = (inputs[167]) & ~(inputs[112]);
    assign layer0_outputs[247] = ~(inputs[87]) | (inputs[148]);
    assign layer0_outputs[248] = inputs[45];
    assign layer0_outputs[249] = (inputs[187]) | (inputs[104]);
    assign layer0_outputs[250] = ~(inputs[68]) | (inputs[177]);
    assign layer0_outputs[251] = (inputs[143]) & ~(inputs[13]);
    assign layer0_outputs[252] = (inputs[162]) & ~(inputs[162]);
    assign layer0_outputs[253] = ~(inputs[86]);
    assign layer0_outputs[254] = ~((inputs[148]) & (inputs[62]));
    assign layer0_outputs[255] = (inputs[74]) & ~(inputs[36]);
    assign layer0_outputs[256] = (inputs[84]) | (inputs[9]);
    assign layer0_outputs[257] = (inputs[97]) & ~(inputs[174]);
    assign layer0_outputs[258] = inputs[132];
    assign layer0_outputs[259] = (inputs[51]) | (inputs[154]);
    assign layer0_outputs[260] = inputs[69];
    assign layer0_outputs[261] = ~((inputs[88]) | (inputs[115]));
    assign layer0_outputs[262] = (inputs[219]) & ~(inputs[5]);
    assign layer0_outputs[263] = ~(inputs[39]);
    assign layer0_outputs[264] = ~(inputs[27]);
    assign layer0_outputs[265] = (inputs[142]) & ~(inputs[207]);
    assign layer0_outputs[266] = ~(inputs[101]);
    assign layer0_outputs[267] = ~((inputs[248]) & (inputs[161]));
    assign layer0_outputs[268] = (inputs[204]) & (inputs[119]);
    assign layer0_outputs[269] = (inputs[23]) ^ (inputs[78]);
    assign layer0_outputs[270] = (inputs[155]) & (inputs[109]);
    assign layer0_outputs[271] = 1'b1;
    assign layer0_outputs[272] = (inputs[193]) | (inputs[251]);
    assign layer0_outputs[273] = (inputs[112]) | (inputs[149]);
    assign layer0_outputs[274] = 1'b1;
    assign layer0_outputs[275] = ~(inputs[123]) | (inputs[244]);
    assign layer0_outputs[276] = (inputs[231]) | (inputs[170]);
    assign layer0_outputs[277] = (inputs[34]) & (inputs[251]);
    assign layer0_outputs[278] = ~(inputs[35]) | (inputs[95]);
    assign layer0_outputs[279] = inputs[109];
    assign layer0_outputs[280] = ~(inputs[61]);
    assign layer0_outputs[281] = (inputs[86]) | (inputs[149]);
    assign layer0_outputs[282] = (inputs[220]) & ~(inputs[64]);
    assign layer0_outputs[283] = (inputs[53]) & ~(inputs[165]);
    assign layer0_outputs[284] = ~((inputs[5]) | (inputs[9]));
    assign layer0_outputs[285] = (inputs[188]) ^ (inputs[117]);
    assign layer0_outputs[286] = (inputs[142]) & ~(inputs[55]);
    assign layer0_outputs[287] = (inputs[103]) & ~(inputs[54]);
    assign layer0_outputs[288] = ~((inputs[88]) | (inputs[62]));
    assign layer0_outputs[289] = (inputs[224]) & ~(inputs[82]);
    assign layer0_outputs[290] = ~(inputs[126]) | (inputs[111]);
    assign layer0_outputs[291] = ~((inputs[71]) & (inputs[241]));
    assign layer0_outputs[292] = 1'b1;
    assign layer0_outputs[293] = inputs[175];
    assign layer0_outputs[294] = ~(inputs[145]) | (inputs[57]);
    assign layer0_outputs[295] = ~(inputs[246]);
    assign layer0_outputs[296] = ~(inputs[154]) | (inputs[187]);
    assign layer0_outputs[297] = ~(inputs[46]);
    assign layer0_outputs[298] = ~(inputs[129]) | (inputs[120]);
    assign layer0_outputs[299] = ~((inputs[198]) ^ (inputs[213]));
    assign layer0_outputs[300] = ~((inputs[182]) | (inputs[229]));
    assign layer0_outputs[301] = (inputs[38]) | (inputs[53]);
    assign layer0_outputs[302] = 1'b0;
    assign layer0_outputs[303] = (inputs[227]) & ~(inputs[8]);
    assign layer0_outputs[304] = inputs[92];
    assign layer0_outputs[305] = ~(inputs[187]) | (inputs[5]);
    assign layer0_outputs[306] = ~((inputs[234]) & (inputs[142]));
    assign layer0_outputs[307] = ~(inputs[111]) | (inputs[7]);
    assign layer0_outputs[308] = 1'b1;
    assign layer0_outputs[309] = ~(inputs[19]) | (inputs[123]);
    assign layer0_outputs[310] = (inputs[24]) & ~(inputs[172]);
    assign layer0_outputs[311] = 1'b0;
    assign layer0_outputs[312] = (inputs[221]) & ~(inputs[158]);
    assign layer0_outputs[313] = ~((inputs[49]) & (inputs[19]));
    assign layer0_outputs[314] = 1'b0;
    assign layer0_outputs[315] = ~(inputs[177]) | (inputs[173]);
    assign layer0_outputs[316] = ~((inputs[73]) & (inputs[186]));
    assign layer0_outputs[317] = ~(inputs[225]);
    assign layer0_outputs[318] = ~(inputs[61]);
    assign layer0_outputs[319] = (inputs[144]) | (inputs[112]);
    assign layer0_outputs[320] = (inputs[142]) ^ (inputs[191]);
    assign layer0_outputs[321] = ~((inputs[240]) ^ (inputs[184]));
    assign layer0_outputs[322] = (inputs[151]) | (inputs[6]);
    assign layer0_outputs[323] = ~(inputs[37]) | (inputs[150]);
    assign layer0_outputs[324] = 1'b0;
    assign layer0_outputs[325] = ~((inputs[39]) ^ (inputs[70]));
    assign layer0_outputs[326] = ~((inputs[109]) & (inputs[55]));
    assign layer0_outputs[327] = (inputs[183]) & ~(inputs[131]);
    assign layer0_outputs[328] = inputs[139];
    assign layer0_outputs[329] = inputs[2];
    assign layer0_outputs[330] = ~(inputs[161]);
    assign layer0_outputs[331] = 1'b1;
    assign layer0_outputs[332] = ~((inputs[118]) & (inputs[87]));
    assign layer0_outputs[333] = inputs[109];
    assign layer0_outputs[334] = ~((inputs[184]) ^ (inputs[189]));
    assign layer0_outputs[335] = ~((inputs[79]) | (inputs[159]));
    assign layer0_outputs[336] = ~(inputs[136]);
    assign layer0_outputs[337] = (inputs[134]) ^ (inputs[226]);
    assign layer0_outputs[338] = ~(inputs[163]) | (inputs[102]);
    assign layer0_outputs[339] = inputs[134];
    assign layer0_outputs[340] = (inputs[176]) | (inputs[110]);
    assign layer0_outputs[341] = 1'b1;
    assign layer0_outputs[342] = (inputs[147]) | (inputs[99]);
    assign layer0_outputs[343] = inputs[91];
    assign layer0_outputs[344] = inputs[96];
    assign layer0_outputs[345] = ~(inputs[126]) | (inputs[119]);
    assign layer0_outputs[346] = ~(inputs[106]) | (inputs[139]);
    assign layer0_outputs[347] = 1'b1;
    assign layer0_outputs[348] = (inputs[214]) | (inputs[239]);
    assign layer0_outputs[349] = ~(inputs[213]);
    assign layer0_outputs[350] = 1'b0;
    assign layer0_outputs[351] = ~((inputs[123]) | (inputs[193]));
    assign layer0_outputs[352] = (inputs[143]) & ~(inputs[17]);
    assign layer0_outputs[353] = 1'b0;
    assign layer0_outputs[354] = (inputs[84]) & (inputs[145]);
    assign layer0_outputs[355] = (inputs[217]) ^ (inputs[196]);
    assign layer0_outputs[356] = (inputs[11]) ^ (inputs[137]);
    assign layer0_outputs[357] = ~((inputs[164]) | (inputs[156]));
    assign layer0_outputs[358] = 1'b0;
    assign layer0_outputs[359] = inputs[89];
    assign layer0_outputs[360] = inputs[246];
    assign layer0_outputs[361] = 1'b0;
    assign layer0_outputs[362] = inputs[3];
    assign layer0_outputs[363] = ~(inputs[251]) | (inputs[157]);
    assign layer0_outputs[364] = ~(inputs[250]);
    assign layer0_outputs[365] = (inputs[186]) & (inputs[199]);
    assign layer0_outputs[366] = (inputs[228]) | (inputs[98]);
    assign layer0_outputs[367] = ~(inputs[131]);
    assign layer0_outputs[368] = ~(inputs[46]);
    assign layer0_outputs[369] = (inputs[237]) & (inputs[120]);
    assign layer0_outputs[370] = (inputs[50]) & (inputs[215]);
    assign layer0_outputs[371] = inputs[192];
    assign layer0_outputs[372] = (inputs[197]) & (inputs[146]);
    assign layer0_outputs[373] = ~(inputs[250]) | (inputs[142]);
    assign layer0_outputs[374] = ~((inputs[173]) | (inputs[72]));
    assign layer0_outputs[375] = ~(inputs[112]);
    assign layer0_outputs[376] = inputs[233];
    assign layer0_outputs[377] = ~(inputs[222]) | (inputs[249]);
    assign layer0_outputs[378] = ~((inputs[139]) ^ (inputs[3]));
    assign layer0_outputs[379] = inputs[44];
    assign layer0_outputs[380] = ~((inputs[195]) & (inputs[10]));
    assign layer0_outputs[381] = (inputs[86]) | (inputs[92]);
    assign layer0_outputs[382] = (inputs[53]) ^ (inputs[115]);
    assign layer0_outputs[383] = 1'b1;
    assign layer0_outputs[384] = ~(inputs[124]) | (inputs[250]);
    assign layer0_outputs[385] = ~((inputs[58]) | (inputs[223]));
    assign layer0_outputs[386] = inputs[231];
    assign layer0_outputs[387] = ~(inputs[137]);
    assign layer0_outputs[388] = ~((inputs[46]) & (inputs[173]));
    assign layer0_outputs[389] = (inputs[231]) | (inputs[144]);
    assign layer0_outputs[390] = 1'b1;
    assign layer0_outputs[391] = inputs[131];
    assign layer0_outputs[392] = ~((inputs[196]) ^ (inputs[80]));
    assign layer0_outputs[393] = inputs[68];
    assign layer0_outputs[394] = ~(inputs[191]);
    assign layer0_outputs[395] = ~((inputs[166]) | (inputs[126]));
    assign layer0_outputs[396] = inputs[137];
    assign layer0_outputs[397] = ~(inputs[96]);
    assign layer0_outputs[398] = ~(inputs[212]);
    assign layer0_outputs[399] = ~(inputs[21]);
    assign layer0_outputs[400] = ~((inputs[108]) | (inputs[254]));
    assign layer0_outputs[401] = inputs[190];
    assign layer0_outputs[402] = inputs[249];
    assign layer0_outputs[403] = ~((inputs[115]) & (inputs[253]));
    assign layer0_outputs[404] = inputs[192];
    assign layer0_outputs[405] = ~(inputs[170]) | (inputs[212]);
    assign layer0_outputs[406] = (inputs[46]) | (inputs[241]);
    assign layer0_outputs[407] = ~((inputs[113]) ^ (inputs[95]));
    assign layer0_outputs[408] = ~(inputs[192]) | (inputs[193]);
    assign layer0_outputs[409] = ~(inputs[148]);
    assign layer0_outputs[410] = (inputs[127]) & ~(inputs[65]);
    assign layer0_outputs[411] = inputs[105];
    assign layer0_outputs[412] = 1'b0;
    assign layer0_outputs[413] = (inputs[133]) ^ (inputs[147]);
    assign layer0_outputs[414] = (inputs[38]) | (inputs[172]);
    assign layer0_outputs[415] = inputs[136];
    assign layer0_outputs[416] = (inputs[126]) & ~(inputs[1]);
    assign layer0_outputs[417] = ~(inputs[66]) | (inputs[2]);
    assign layer0_outputs[418] = (inputs[175]) & ~(inputs[244]);
    assign layer0_outputs[419] = (inputs[33]) | (inputs[222]);
    assign layer0_outputs[420] = ~((inputs[163]) & (inputs[115]));
    assign layer0_outputs[421] = (inputs[153]) | (inputs[114]);
    assign layer0_outputs[422] = ~((inputs[32]) | (inputs[195]));
    assign layer0_outputs[423] = ~(inputs[55]);
    assign layer0_outputs[424] = ~(inputs[219]);
    assign layer0_outputs[425] = (inputs[40]) & (inputs[217]);
    assign layer0_outputs[426] = (inputs[59]) & ~(inputs[169]);
    assign layer0_outputs[427] = ~(inputs[40]);
    assign layer0_outputs[428] = (inputs[7]) & ~(inputs[64]);
    assign layer0_outputs[429] = inputs[22];
    assign layer0_outputs[430] = (inputs[83]) & ~(inputs[88]);
    assign layer0_outputs[431] = inputs[45];
    assign layer0_outputs[432] = (inputs[24]) | (inputs[120]);
    assign layer0_outputs[433] = ~(inputs[191]) | (inputs[241]);
    assign layer0_outputs[434] = (inputs[32]) & ~(inputs[208]);
    assign layer0_outputs[435] = ~(inputs[188]) | (inputs[108]);
    assign layer0_outputs[436] = ~(inputs[191]);
    assign layer0_outputs[437] = inputs[46];
    assign layer0_outputs[438] = (inputs[80]) | (inputs[204]);
    assign layer0_outputs[439] = ~(inputs[54]);
    assign layer0_outputs[440] = ~((inputs[164]) | (inputs[170]));
    assign layer0_outputs[441] = (inputs[213]) ^ (inputs[13]);
    assign layer0_outputs[442] = (inputs[61]) & ~(inputs[180]);
    assign layer0_outputs[443] = 1'b0;
    assign layer0_outputs[444] = ~((inputs[64]) | (inputs[211]));
    assign layer0_outputs[445] = inputs[156];
    assign layer0_outputs[446] = ~(inputs[209]) | (inputs[180]);
    assign layer0_outputs[447] = ~((inputs[59]) & (inputs[21]));
    assign layer0_outputs[448] = ~((inputs[206]) | (inputs[173]));
    assign layer0_outputs[449] = ~((inputs[79]) & (inputs[136]));
    assign layer0_outputs[450] = ~(inputs[53]) | (inputs[248]);
    assign layer0_outputs[451] = (inputs[204]) | (inputs[141]);
    assign layer0_outputs[452] = ~(inputs[134]) | (inputs[112]);
    assign layer0_outputs[453] = (inputs[19]) & ~(inputs[163]);
    assign layer0_outputs[454] = (inputs[2]) & (inputs[156]);
    assign layer0_outputs[455] = 1'b1;
    assign layer0_outputs[456] = ~((inputs[125]) & (inputs[139]));
    assign layer0_outputs[457] = (inputs[241]) & ~(inputs[68]);
    assign layer0_outputs[458] = (inputs[219]) | (inputs[63]);
    assign layer0_outputs[459] = ~(inputs[221]) | (inputs[3]);
    assign layer0_outputs[460] = ~(inputs[188]);
    assign layer0_outputs[461] = (inputs[179]) | (inputs[71]);
    assign layer0_outputs[462] = ~(inputs[168]) | (inputs[179]);
    assign layer0_outputs[463] = (inputs[123]) | (inputs[49]);
    assign layer0_outputs[464] = ~((inputs[179]) ^ (inputs[235]));
    assign layer0_outputs[465] = ~(inputs[55]);
    assign layer0_outputs[466] = 1'b1;
    assign layer0_outputs[467] = ~(inputs[216]) | (inputs[252]);
    assign layer0_outputs[468] = (inputs[185]) & ~(inputs[67]);
    assign layer0_outputs[469] = 1'b1;
    assign layer0_outputs[470] = 1'b0;
    assign layer0_outputs[471] = 1'b0;
    assign layer0_outputs[472] = 1'b0;
    assign layer0_outputs[473] = (inputs[164]) & ~(inputs[26]);
    assign layer0_outputs[474] = ~((inputs[9]) ^ (inputs[0]));
    assign layer0_outputs[475] = (inputs[181]) & ~(inputs[50]);
    assign layer0_outputs[476] = ~(inputs[162]) | (inputs[239]);
    assign layer0_outputs[477] = (inputs[72]) | (inputs[138]);
    assign layer0_outputs[478] = ~((inputs[64]) | (inputs[239]));
    assign layer0_outputs[479] = (inputs[79]) & (inputs[14]);
    assign layer0_outputs[480] = inputs[13];
    assign layer0_outputs[481] = ~(inputs[240]) | (inputs[123]);
    assign layer0_outputs[482] = ~(inputs[162]) | (inputs[102]);
    assign layer0_outputs[483] = ~((inputs[78]) | (inputs[207]));
    assign layer0_outputs[484] = ~(inputs[194]) | (inputs[188]);
    assign layer0_outputs[485] = ~(inputs[116]);
    assign layer0_outputs[486] = inputs[143];
    assign layer0_outputs[487] = (inputs[150]) ^ (inputs[237]);
    assign layer0_outputs[488] = (inputs[79]) | (inputs[147]);
    assign layer0_outputs[489] = 1'b1;
    assign layer0_outputs[490] = 1'b1;
    assign layer0_outputs[491] = (inputs[171]) & (inputs[191]);
    assign layer0_outputs[492] = (inputs[148]) | (inputs[5]);
    assign layer0_outputs[493] = 1'b0;
    assign layer0_outputs[494] = 1'b1;
    assign layer0_outputs[495] = (inputs[78]) | (inputs[227]);
    assign layer0_outputs[496] = (inputs[177]) & (inputs[210]);
    assign layer0_outputs[497] = ~((inputs[71]) & (inputs[163]));
    assign layer0_outputs[498] = ~(inputs[13]);
    assign layer0_outputs[499] = ~(inputs[208]);
    assign layer0_outputs[500] = ~(inputs[151]);
    assign layer0_outputs[501] = 1'b0;
    assign layer0_outputs[502] = ~(inputs[34]) | (inputs[11]);
    assign layer0_outputs[503] = ~((inputs[110]) ^ (inputs[91]));
    assign layer0_outputs[504] = ~(inputs[149]) | (inputs[82]);
    assign layer0_outputs[505] = 1'b0;
    assign layer0_outputs[506] = ~(inputs[171]) | (inputs[241]);
    assign layer0_outputs[507] = (inputs[86]) & ~(inputs[211]);
    assign layer0_outputs[508] = 1'b1;
    assign layer0_outputs[509] = ~((inputs[141]) | (inputs[70]));
    assign layer0_outputs[510] = (inputs[134]) & ~(inputs[248]);
    assign layer0_outputs[511] = ~(inputs[182]);
    assign layer0_outputs[512] = inputs[187];
    assign layer0_outputs[513] = ~((inputs[215]) | (inputs[213]));
    assign layer0_outputs[514] = ~((inputs[205]) & (inputs[79]));
    assign layer0_outputs[515] = (inputs[225]) & ~(inputs[162]);
    assign layer0_outputs[516] = ~((inputs[83]) & (inputs[142]));
    assign layer0_outputs[517] = (inputs[100]) & ~(inputs[209]);
    assign layer0_outputs[518] = ~((inputs[4]) ^ (inputs[158]));
    assign layer0_outputs[519] = ~(inputs[204]);
    assign layer0_outputs[520] = ~((inputs[174]) & (inputs[216]));
    assign layer0_outputs[521] = (inputs[27]) & ~(inputs[93]);
    assign layer0_outputs[522] = inputs[177];
    assign layer0_outputs[523] = 1'b1;
    assign layer0_outputs[524] = inputs[71];
    assign layer0_outputs[525] = inputs[51];
    assign layer0_outputs[526] = (inputs[14]) & (inputs[29]);
    assign layer0_outputs[527] = ~(inputs[128]) | (inputs[226]);
    assign layer0_outputs[528] = inputs[58];
    assign layer0_outputs[529] = ~((inputs[36]) & (inputs[121]));
    assign layer0_outputs[530] = ~((inputs[116]) ^ (inputs[243]));
    assign layer0_outputs[531] = inputs[101];
    assign layer0_outputs[532] = (inputs[33]) & (inputs[88]);
    assign layer0_outputs[533] = ~((inputs[33]) ^ (inputs[98]));
    assign layer0_outputs[534] = ~((inputs[75]) | (inputs[31]));
    assign layer0_outputs[535] = ~(inputs[180]) | (inputs[212]);
    assign layer0_outputs[536] = ~((inputs[31]) & (inputs[135]));
    assign layer0_outputs[537] = (inputs[48]) ^ (inputs[57]);
    assign layer0_outputs[538] = ~((inputs[101]) & (inputs[40]));
    assign layer0_outputs[539] = ~((inputs[41]) | (inputs[171]));
    assign layer0_outputs[540] = inputs[238];
    assign layer0_outputs[541] = ~((inputs[246]) & (inputs[76]));
    assign layer0_outputs[542] = (inputs[227]) | (inputs[125]);
    assign layer0_outputs[543] = inputs[215];
    assign layer0_outputs[544] = inputs[13];
    assign layer0_outputs[545] = 1'b1;
    assign layer0_outputs[546] = (inputs[231]) & (inputs[39]);
    assign layer0_outputs[547] = (inputs[89]) | (inputs[95]);
    assign layer0_outputs[548] = (inputs[182]) | (inputs[81]);
    assign layer0_outputs[549] = inputs[116];
    assign layer0_outputs[550] = ~((inputs[213]) | (inputs[254]));
    assign layer0_outputs[551] = 1'b0;
    assign layer0_outputs[552] = 1'b0;
    assign layer0_outputs[553] = 1'b0;
    assign layer0_outputs[554] = (inputs[88]) & ~(inputs[230]);
    assign layer0_outputs[555] = (inputs[83]) & ~(inputs[237]);
    assign layer0_outputs[556] = (inputs[98]) & ~(inputs[212]);
    assign layer0_outputs[557] = ~((inputs[165]) & (inputs[223]));
    assign layer0_outputs[558] = (inputs[7]) & ~(inputs[110]);
    assign layer0_outputs[559] = ~(inputs[220]);
    assign layer0_outputs[560] = (inputs[254]) & ~(inputs[72]);
    assign layer0_outputs[561] = (inputs[79]) & ~(inputs[110]);
    assign layer0_outputs[562] = ~(inputs[243]) | (inputs[99]);
    assign layer0_outputs[563] = ~((inputs[157]) | (inputs[255]));
    assign layer0_outputs[564] = (inputs[165]) ^ (inputs[15]);
    assign layer0_outputs[565] = ~((inputs[28]) & (inputs[88]));
    assign layer0_outputs[566] = (inputs[20]) ^ (inputs[135]);
    assign layer0_outputs[567] = ~((inputs[139]) | (inputs[64]));
    assign layer0_outputs[568] = (inputs[81]) | (inputs[216]);
    assign layer0_outputs[569] = inputs[9];
    assign layer0_outputs[570] = (inputs[82]) | (inputs[245]);
    assign layer0_outputs[571] = ~(inputs[106]);
    assign layer0_outputs[572] = (inputs[20]) ^ (inputs[243]);
    assign layer0_outputs[573] = inputs[232];
    assign layer0_outputs[574] = ~(inputs[209]);
    assign layer0_outputs[575] = ~(inputs[99]) | (inputs[99]);
    assign layer0_outputs[576] = 1'b1;
    assign layer0_outputs[577] = ~((inputs[65]) & (inputs[129]));
    assign layer0_outputs[578] = ~((inputs[51]) | (inputs[206]));
    assign layer0_outputs[579] = ~(inputs[191]);
    assign layer0_outputs[580] = ~(inputs[52]) | (inputs[98]);
    assign layer0_outputs[581] = ~(inputs[171]);
    assign layer0_outputs[582] = 1'b0;
    assign layer0_outputs[583] = ~((inputs[122]) | (inputs[150]));
    assign layer0_outputs[584] = ~(inputs[242]);
    assign layer0_outputs[585] = 1'b0;
    assign layer0_outputs[586] = ~(inputs[197]) | (inputs[125]);
    assign layer0_outputs[587] = (inputs[127]) & ~(inputs[242]);
    assign layer0_outputs[588] = (inputs[247]) & ~(inputs[133]);
    assign layer0_outputs[589] = ~(inputs[50]);
    assign layer0_outputs[590] = ~(inputs[228]);
    assign layer0_outputs[591] = 1'b0;
    assign layer0_outputs[592] = ~(inputs[108]);
    assign layer0_outputs[593] = ~(inputs[170]) | (inputs[133]);
    assign layer0_outputs[594] = ~(inputs[196]);
    assign layer0_outputs[595] = ~(inputs[105]);
    assign layer0_outputs[596] = (inputs[80]) & ~(inputs[101]);
    assign layer0_outputs[597] = ~(inputs[1]) | (inputs[108]);
    assign layer0_outputs[598] = 1'b0;
    assign layer0_outputs[599] = ~((inputs[219]) ^ (inputs[130]));
    assign layer0_outputs[600] = 1'b1;
    assign layer0_outputs[601] = ~(inputs[39]);
    assign layer0_outputs[602] = ~(inputs[207]) | (inputs[81]);
    assign layer0_outputs[603] = inputs[145];
    assign layer0_outputs[604] = ~(inputs[210]);
    assign layer0_outputs[605] = ~(inputs[120]) | (inputs[169]);
    assign layer0_outputs[606] = ~(inputs[125]);
    assign layer0_outputs[607] = (inputs[134]) & ~(inputs[181]);
    assign layer0_outputs[608] = 1'b1;
    assign layer0_outputs[609] = ~((inputs[181]) ^ (inputs[31]));
    assign layer0_outputs[610] = (inputs[126]) ^ (inputs[125]);
    assign layer0_outputs[611] = (inputs[199]) & ~(inputs[221]);
    assign layer0_outputs[612] = ~((inputs[172]) & (inputs[229]));
    assign layer0_outputs[613] = (inputs[13]) | (inputs[118]);
    assign layer0_outputs[614] = ~((inputs[203]) | (inputs[56]));
    assign layer0_outputs[615] = ~((inputs[241]) & (inputs[139]));
    assign layer0_outputs[616] = ~((inputs[108]) & (inputs[16]));
    assign layer0_outputs[617] = ~((inputs[51]) ^ (inputs[229]));
    assign layer0_outputs[618] = (inputs[89]) & ~(inputs[78]);
    assign layer0_outputs[619] = (inputs[151]) & ~(inputs[172]);
    assign layer0_outputs[620] = ~(inputs[55]) | (inputs[207]);
    assign layer0_outputs[621] = inputs[97];
    assign layer0_outputs[622] = (inputs[196]) & ~(inputs[87]);
    assign layer0_outputs[623] = (inputs[62]) & ~(inputs[135]);
    assign layer0_outputs[624] = ~(inputs[221]) | (inputs[216]);
    assign layer0_outputs[625] = 1'b1;
    assign layer0_outputs[626] = ~(inputs[38]) | (inputs[20]);
    assign layer0_outputs[627] = ~(inputs[63]);
    assign layer0_outputs[628] = ~(inputs[162]);
    assign layer0_outputs[629] = ~((inputs[203]) & (inputs[41]));
    assign layer0_outputs[630] = (inputs[104]) & ~(inputs[225]);
    assign layer0_outputs[631] = ~(inputs[158]) | (inputs[16]);
    assign layer0_outputs[632] = ~((inputs[101]) | (inputs[93]));
    assign layer0_outputs[633] = ~(inputs[104]);
    assign layer0_outputs[634] = ~((inputs[144]) & (inputs[68]));
    assign layer0_outputs[635] = (inputs[107]) & (inputs[83]);
    assign layer0_outputs[636] = ~((inputs[46]) ^ (inputs[152]));
    assign layer0_outputs[637] = (inputs[178]) | (inputs[210]);
    assign layer0_outputs[638] = (inputs[230]) & ~(inputs[184]);
    assign layer0_outputs[639] = ~(inputs[182]);
    assign layer0_outputs[640] = ~(inputs[121]);
    assign layer0_outputs[641] = ~(inputs[243]) | (inputs[148]);
    assign layer0_outputs[642] = inputs[155];
    assign layer0_outputs[643] = ~((inputs[47]) | (inputs[174]));
    assign layer0_outputs[644] = 1'b1;
    assign layer0_outputs[645] = (inputs[13]) ^ (inputs[247]);
    assign layer0_outputs[646] = ~(inputs[156]);
    assign layer0_outputs[647] = ~(inputs[4]) | (inputs[121]);
    assign layer0_outputs[648] = (inputs[107]) | (inputs[89]);
    assign layer0_outputs[649] = (inputs[119]) & ~(inputs[164]);
    assign layer0_outputs[650] = ~(inputs[14]);
    assign layer0_outputs[651] = ~(inputs[197]);
    assign layer0_outputs[652] = ~(inputs[106]) | (inputs[132]);
    assign layer0_outputs[653] = ~(inputs[227]) | (inputs[48]);
    assign layer0_outputs[654] = inputs[206];
    assign layer0_outputs[655] = (inputs[120]) | (inputs[47]);
    assign layer0_outputs[656] = ~((inputs[103]) ^ (inputs[97]));
    assign layer0_outputs[657] = ~(inputs[194]);
    assign layer0_outputs[658] = ~(inputs[137]) | (inputs[225]);
    assign layer0_outputs[659] = (inputs[81]) | (inputs[125]);
    assign layer0_outputs[660] = (inputs[113]) & (inputs[74]);
    assign layer0_outputs[661] = inputs[222];
    assign layer0_outputs[662] = ~(inputs[136]) | (inputs[156]);
    assign layer0_outputs[663] = (inputs[60]) ^ (inputs[26]);
    assign layer0_outputs[664] = ~((inputs[11]) | (inputs[127]));
    assign layer0_outputs[665] = ~(inputs[107]);
    assign layer0_outputs[666] = (inputs[154]) & ~(inputs[143]);
    assign layer0_outputs[667] = inputs[72];
    assign layer0_outputs[668] = ~(inputs[255]) | (inputs[79]);
    assign layer0_outputs[669] = (inputs[88]) & ~(inputs[14]);
    assign layer0_outputs[670] = (inputs[133]) & ~(inputs[42]);
    assign layer0_outputs[671] = (inputs[137]) ^ (inputs[221]);
    assign layer0_outputs[672] = ~(inputs[30]) | (inputs[58]);
    assign layer0_outputs[673] = (inputs[2]) & (inputs[78]);
    assign layer0_outputs[674] = (inputs[14]) & (inputs[190]);
    assign layer0_outputs[675] = inputs[218];
    assign layer0_outputs[676] = (inputs[166]) & ~(inputs[223]);
    assign layer0_outputs[677] = (inputs[92]) & ~(inputs[250]);
    assign layer0_outputs[678] = ~(inputs[171]);
    assign layer0_outputs[679] = ~((inputs[204]) | (inputs[25]));
    assign layer0_outputs[680] = ~(inputs[192]) | (inputs[33]);
    assign layer0_outputs[681] = (inputs[60]) | (inputs[223]);
    assign layer0_outputs[682] = ~(inputs[252]) | (inputs[126]);
    assign layer0_outputs[683] = (inputs[171]) & ~(inputs[172]);
    assign layer0_outputs[684] = inputs[108];
    assign layer0_outputs[685] = 1'b0;
    assign layer0_outputs[686] = (inputs[233]) & ~(inputs[167]);
    assign layer0_outputs[687] = ~(inputs[37]) | (inputs[90]);
    assign layer0_outputs[688] = (inputs[93]) | (inputs[252]);
    assign layer0_outputs[689] = ~(inputs[94]) | (inputs[35]);
    assign layer0_outputs[690] = ~(inputs[57]) | (inputs[25]);
    assign layer0_outputs[691] = ~(inputs[62]);
    assign layer0_outputs[692] = ~((inputs[70]) | (inputs[198]));
    assign layer0_outputs[693] = (inputs[171]) | (inputs[202]);
    assign layer0_outputs[694] = (inputs[206]) & (inputs[160]);
    assign layer0_outputs[695] = ~((inputs[250]) | (inputs[193]));
    assign layer0_outputs[696] = (inputs[60]) & ~(inputs[207]);
    assign layer0_outputs[697] = ~(inputs[250]);
    assign layer0_outputs[698] = ~(inputs[81]);
    assign layer0_outputs[699] = inputs[72];
    assign layer0_outputs[700] = 1'b1;
    assign layer0_outputs[701] = 1'b1;
    assign layer0_outputs[702] = inputs[45];
    assign layer0_outputs[703] = ~((inputs[51]) & (inputs[83]));
    assign layer0_outputs[704] = (inputs[142]) & ~(inputs[3]);
    assign layer0_outputs[705] = ~(inputs[24]);
    assign layer0_outputs[706] = (inputs[126]) | (inputs[186]);
    assign layer0_outputs[707] = (inputs[102]) | (inputs[114]);
    assign layer0_outputs[708] = (inputs[235]) ^ (inputs[61]);
    assign layer0_outputs[709] = ~((inputs[228]) | (inputs[100]));
    assign layer0_outputs[710] = inputs[113];
    assign layer0_outputs[711] = (inputs[51]) ^ (inputs[81]);
    assign layer0_outputs[712] = ~(inputs[57]);
    assign layer0_outputs[713] = ~(inputs[151]) | (inputs[121]);
    assign layer0_outputs[714] = ~((inputs[157]) | (inputs[100]));
    assign layer0_outputs[715] = ~(inputs[141]) | (inputs[255]);
    assign layer0_outputs[716] = 1'b0;
    assign layer0_outputs[717] = (inputs[95]) | (inputs[50]);
    assign layer0_outputs[718] = 1'b1;
    assign layer0_outputs[719] = 1'b1;
    assign layer0_outputs[720] = 1'b1;
    assign layer0_outputs[721] = ~(inputs[216]) | (inputs[194]);
    assign layer0_outputs[722] = ~(inputs[147]);
    assign layer0_outputs[723] = 1'b1;
    assign layer0_outputs[724] = inputs[237];
    assign layer0_outputs[725] = (inputs[65]) | (inputs[118]);
    assign layer0_outputs[726] = 1'b0;
    assign layer0_outputs[727] = ~((inputs[146]) & (inputs[157]));
    assign layer0_outputs[728] = ~((inputs[99]) | (inputs[228]));
    assign layer0_outputs[729] = ~(inputs[234]);
    assign layer0_outputs[730] = ~(inputs[61]) | (inputs[96]);
    assign layer0_outputs[731] = ~((inputs[255]) | (inputs[36]));
    assign layer0_outputs[732] = 1'b1;
    assign layer0_outputs[733] = (inputs[24]) ^ (inputs[148]);
    assign layer0_outputs[734] = (inputs[195]) & ~(inputs[229]);
    assign layer0_outputs[735] = (inputs[12]) & ~(inputs[49]);
    assign layer0_outputs[736] = 1'b0;
    assign layer0_outputs[737] = 1'b0;
    assign layer0_outputs[738] = ~((inputs[252]) | (inputs[44]));
    assign layer0_outputs[739] = ~((inputs[212]) | (inputs[188]));
    assign layer0_outputs[740] = (inputs[27]) | (inputs[45]);
    assign layer0_outputs[741] = ~((inputs[28]) | (inputs[122]));
    assign layer0_outputs[742] = inputs[251];
    assign layer0_outputs[743] = (inputs[245]) & (inputs[219]);
    assign layer0_outputs[744] = (inputs[118]) & ~(inputs[233]);
    assign layer0_outputs[745] = 1'b1;
    assign layer0_outputs[746] = ~(inputs[99]);
    assign layer0_outputs[747] = ~(inputs[236]);
    assign layer0_outputs[748] = ~(inputs[6]) | (inputs[22]);
    assign layer0_outputs[749] = 1'b1;
    assign layer0_outputs[750] = ~((inputs[220]) | (inputs[161]));
    assign layer0_outputs[751] = ~(inputs[31]) | (inputs[175]);
    assign layer0_outputs[752] = ~(inputs[86]);
    assign layer0_outputs[753] = inputs[6];
    assign layer0_outputs[754] = ~(inputs[32]);
    assign layer0_outputs[755] = (inputs[32]) & ~(inputs[224]);
    assign layer0_outputs[756] = (inputs[19]) & ~(inputs[190]);
    assign layer0_outputs[757] = 1'b1;
    assign layer0_outputs[758] = ~(inputs[13]) | (inputs[232]);
    assign layer0_outputs[759] = ~(inputs[240]) | (inputs[9]);
    assign layer0_outputs[760] = ~(inputs[153]);
    assign layer0_outputs[761] = ~(inputs[248]) | (inputs[115]);
    assign layer0_outputs[762] = (inputs[84]) & ~(inputs[87]);
    assign layer0_outputs[763] = (inputs[154]) & ~(inputs[199]);
    assign layer0_outputs[764] = ~(inputs[185]);
    assign layer0_outputs[765] = ~((inputs[32]) ^ (inputs[14]));
    assign layer0_outputs[766] = (inputs[83]) & (inputs[254]);
    assign layer0_outputs[767] = ~(inputs[1]) | (inputs[93]);
    assign layer0_outputs[768] = (inputs[137]) & ~(inputs[53]);
    assign layer0_outputs[769] = (inputs[183]) ^ (inputs[17]);
    assign layer0_outputs[770] = 1'b1;
    assign layer0_outputs[771] = ~(inputs[140]);
    assign layer0_outputs[772] = 1'b1;
    assign layer0_outputs[773] = 1'b0;
    assign layer0_outputs[774] = (inputs[128]) ^ (inputs[82]);
    assign layer0_outputs[775] = (inputs[49]) ^ (inputs[113]);
    assign layer0_outputs[776] = ~((inputs[195]) | (inputs[210]));
    assign layer0_outputs[777] = (inputs[157]) | (inputs[124]);
    assign layer0_outputs[778] = ~((inputs[122]) ^ (inputs[177]));
    assign layer0_outputs[779] = 1'b1;
    assign layer0_outputs[780] = ~((inputs[86]) ^ (inputs[111]));
    assign layer0_outputs[781] = 1'b1;
    assign layer0_outputs[782] = inputs[202];
    assign layer0_outputs[783] = ~(inputs[46]) | (inputs[201]);
    assign layer0_outputs[784] = (inputs[143]) | (inputs[42]);
    assign layer0_outputs[785] = inputs[64];
    assign layer0_outputs[786] = inputs[231];
    assign layer0_outputs[787] = ~(inputs[80]);
    assign layer0_outputs[788] = ~(inputs[163]);
    assign layer0_outputs[789] = inputs[246];
    assign layer0_outputs[790] = ~((inputs[235]) | (inputs[193]));
    assign layer0_outputs[791] = ~((inputs[143]) ^ (inputs[35]));
    assign layer0_outputs[792] = inputs[247];
    assign layer0_outputs[793] = ~(inputs[105]);
    assign layer0_outputs[794] = ~(inputs[85]) | (inputs[177]);
    assign layer0_outputs[795] = ~((inputs[147]) | (inputs[164]));
    assign layer0_outputs[796] = (inputs[32]) | (inputs[45]);
    assign layer0_outputs[797] = inputs[49];
    assign layer0_outputs[798] = (inputs[210]) & ~(inputs[194]);
    assign layer0_outputs[799] = (inputs[83]) & (inputs[144]);
    assign layer0_outputs[800] = (inputs[149]) & ~(inputs[161]);
    assign layer0_outputs[801] = 1'b1;
    assign layer0_outputs[802] = ~(inputs[252]) | (inputs[121]);
    assign layer0_outputs[803] = inputs[28];
    assign layer0_outputs[804] = ~(inputs[181]) | (inputs[50]);
    assign layer0_outputs[805] = 1'b1;
    assign layer0_outputs[806] = ~((inputs[36]) & (inputs[239]));
    assign layer0_outputs[807] = inputs[41];
    assign layer0_outputs[808] = ~(inputs[203]);
    assign layer0_outputs[809] = inputs[78];
    assign layer0_outputs[810] = ~(inputs[110]) | (inputs[103]);
    assign layer0_outputs[811] = 1'b1;
    assign layer0_outputs[812] = inputs[155];
    assign layer0_outputs[813] = ~((inputs[103]) | (inputs[85]));
    assign layer0_outputs[814] = ~(inputs[37]);
    assign layer0_outputs[815] = ~(inputs[88]) | (inputs[101]);
    assign layer0_outputs[816] = 1'b0;
    assign layer0_outputs[817] = ~((inputs[17]) ^ (inputs[251]));
    assign layer0_outputs[818] = ~(inputs[234]);
    assign layer0_outputs[819] = ~(inputs[15]);
    assign layer0_outputs[820] = inputs[12];
    assign layer0_outputs[821] = 1'b0;
    assign layer0_outputs[822] = ~(inputs[161]);
    assign layer0_outputs[823] = (inputs[25]) ^ (inputs[93]);
    assign layer0_outputs[824] = ~(inputs[76]) | (inputs[237]);
    assign layer0_outputs[825] = ~(inputs[175]);
    assign layer0_outputs[826] = (inputs[14]) ^ (inputs[128]);
    assign layer0_outputs[827] = ~(inputs[158]) | (inputs[247]);
    assign layer0_outputs[828] = (inputs[91]) & (inputs[14]);
    assign layer0_outputs[829] = ~(inputs[44]) | (inputs[103]);
    assign layer0_outputs[830] = ~(inputs[136]) | (inputs[27]);
    assign layer0_outputs[831] = ~(inputs[234]);
    assign layer0_outputs[832] = ~((inputs[18]) ^ (inputs[115]));
    assign layer0_outputs[833] = (inputs[167]) | (inputs[28]);
    assign layer0_outputs[834] = (inputs[116]) ^ (inputs[189]);
    assign layer0_outputs[835] = (inputs[147]) & ~(inputs[92]);
    assign layer0_outputs[836] = 1'b1;
    assign layer0_outputs[837] = ~((inputs[17]) & (inputs[129]));
    assign layer0_outputs[838] = (inputs[91]) & ~(inputs[244]);
    assign layer0_outputs[839] = 1'b1;
    assign layer0_outputs[840] = (inputs[52]) | (inputs[154]);
    assign layer0_outputs[841] = ~(inputs[5]) | (inputs[70]);
    assign layer0_outputs[842] = ~(inputs[223]) | (inputs[131]);
    assign layer0_outputs[843] = ~((inputs[181]) & (inputs[10]));
    assign layer0_outputs[844] = ~(inputs[205]);
    assign layer0_outputs[845] = ~(inputs[49]) | (inputs[90]);
    assign layer0_outputs[846] = ~(inputs[166]) | (inputs[98]);
    assign layer0_outputs[847] = inputs[173];
    assign layer0_outputs[848] = (inputs[116]) & ~(inputs[94]);
    assign layer0_outputs[849] = (inputs[239]) & ~(inputs[153]);
    assign layer0_outputs[850] = ~(inputs[2]);
    assign layer0_outputs[851] = ~((inputs[189]) ^ (inputs[3]));
    assign layer0_outputs[852] = ~(inputs[160]) | (inputs[162]);
    assign layer0_outputs[853] = ~(inputs[211]) | (inputs[4]);
    assign layer0_outputs[854] = ~(inputs[42]) | (inputs[228]);
    assign layer0_outputs[855] = ~(inputs[137]);
    assign layer0_outputs[856] = ~(inputs[85]);
    assign layer0_outputs[857] = 1'b0;
    assign layer0_outputs[858] = (inputs[103]) | (inputs[104]);
    assign layer0_outputs[859] = (inputs[175]) & (inputs[54]);
    assign layer0_outputs[860] = ~((inputs[113]) & (inputs[118]));
    assign layer0_outputs[861] = 1'b0;
    assign layer0_outputs[862] = ~(inputs[54]);
    assign layer0_outputs[863] = ~(inputs[118]);
    assign layer0_outputs[864] = inputs[72];
    assign layer0_outputs[865] = ~((inputs[255]) | (inputs[46]));
    assign layer0_outputs[866] = (inputs[191]) & ~(inputs[206]);
    assign layer0_outputs[867] = (inputs[232]) & ~(inputs[206]);
    assign layer0_outputs[868] = (inputs[149]) ^ (inputs[5]);
    assign layer0_outputs[869] = ~(inputs[217]) | (inputs[227]);
    assign layer0_outputs[870] = ~(inputs[238]);
    assign layer0_outputs[871] = inputs[218];
    assign layer0_outputs[872] = ~((inputs[250]) & (inputs[239]));
    assign layer0_outputs[873] = ~(inputs[177]) | (inputs[178]);
    assign layer0_outputs[874] = ~(inputs[35]) | (inputs[217]);
    assign layer0_outputs[875] = ~(inputs[236]) | (inputs[2]);
    assign layer0_outputs[876] = 1'b0;
    assign layer0_outputs[877] = ~((inputs[187]) | (inputs[123]));
    assign layer0_outputs[878] = ~((inputs[102]) | (inputs[238]));
    assign layer0_outputs[879] = ~(inputs[224]);
    assign layer0_outputs[880] = inputs[212];
    assign layer0_outputs[881] = ~((inputs[210]) & (inputs[233]));
    assign layer0_outputs[882] = ~(inputs[217]) | (inputs[125]);
    assign layer0_outputs[883] = 1'b1;
    assign layer0_outputs[884] = (inputs[197]) ^ (inputs[24]);
    assign layer0_outputs[885] = inputs[22];
    assign layer0_outputs[886] = ~(inputs[63]);
    assign layer0_outputs[887] = (inputs[76]) & (inputs[67]);
    assign layer0_outputs[888] = ~(inputs[196]);
    assign layer0_outputs[889] = 1'b1;
    assign layer0_outputs[890] = ~((inputs[86]) | (inputs[131]));
    assign layer0_outputs[891] = inputs[115];
    assign layer0_outputs[892] = ~(inputs[227]) | (inputs[244]);
    assign layer0_outputs[893] = ~((inputs[81]) ^ (inputs[17]));
    assign layer0_outputs[894] = inputs[1];
    assign layer0_outputs[895] = inputs[8];
    assign layer0_outputs[896] = inputs[174];
    assign layer0_outputs[897] = (inputs[179]) & ~(inputs[93]);
    assign layer0_outputs[898] = ~(inputs[66]) | (inputs[32]);
    assign layer0_outputs[899] = ~(inputs[183]) | (inputs[169]);
    assign layer0_outputs[900] = 1'b1;
    assign layer0_outputs[901] = (inputs[48]) ^ (inputs[237]);
    assign layer0_outputs[902] = (inputs[105]) & ~(inputs[184]);
    assign layer0_outputs[903] = inputs[24];
    assign layer0_outputs[904] = (inputs[109]) & ~(inputs[26]);
    assign layer0_outputs[905] = 1'b0;
    assign layer0_outputs[906] = (inputs[155]) & ~(inputs[82]);
    assign layer0_outputs[907] = ~(inputs[233]);
    assign layer0_outputs[908] = 1'b1;
    assign layer0_outputs[909] = (inputs[119]) & ~(inputs[229]);
    assign layer0_outputs[910] = inputs[3];
    assign layer0_outputs[911] = inputs[38];
    assign layer0_outputs[912] = (inputs[148]) & ~(inputs[217]);
    assign layer0_outputs[913] = (inputs[165]) & (inputs[20]);
    assign layer0_outputs[914] = (inputs[24]) & ~(inputs[32]);
    assign layer0_outputs[915] = ~((inputs[53]) | (inputs[196]));
    assign layer0_outputs[916] = inputs[181];
    assign layer0_outputs[917] = (inputs[31]) & ~(inputs[36]);
    assign layer0_outputs[918] = (inputs[163]) ^ (inputs[91]);
    assign layer0_outputs[919] = 1'b0;
    assign layer0_outputs[920] = (inputs[117]) & ~(inputs[185]);
    assign layer0_outputs[921] = ~((inputs[29]) & (inputs[50]));
    assign layer0_outputs[922] = 1'b1;
    assign layer0_outputs[923] = ~(inputs[68]);
    assign layer0_outputs[924] = ~((inputs[66]) & (inputs[0]));
    assign layer0_outputs[925] = ~((inputs[213]) & (inputs[79]));
    assign layer0_outputs[926] = inputs[139];
    assign layer0_outputs[927] = (inputs[71]) & ~(inputs[168]);
    assign layer0_outputs[928] = (inputs[46]) & ~(inputs[227]);
    assign layer0_outputs[929] = (inputs[193]) & ~(inputs[18]);
    assign layer0_outputs[930] = inputs[3];
    assign layer0_outputs[931] = ~(inputs[147]) | (inputs[232]);
    assign layer0_outputs[932] = ~(inputs[33]);
    assign layer0_outputs[933] = ~(inputs[19]);
    assign layer0_outputs[934] = (inputs[133]) & ~(inputs[190]);
    assign layer0_outputs[935] = (inputs[122]) | (inputs[8]);
    assign layer0_outputs[936] = 1'b0;
    assign layer0_outputs[937] = inputs[119];
    assign layer0_outputs[938] = ~(inputs[167]) | (inputs[78]);
    assign layer0_outputs[939] = inputs[89];
    assign layer0_outputs[940] = 1'b1;
    assign layer0_outputs[941] = ~(inputs[24]) | (inputs[226]);
    assign layer0_outputs[942] = ~(inputs[97]) | (inputs[8]);
    assign layer0_outputs[943] = ~((inputs[116]) | (inputs[9]));
    assign layer0_outputs[944] = (inputs[77]) & (inputs[9]);
    assign layer0_outputs[945] = (inputs[136]) & ~(inputs[226]);
    assign layer0_outputs[946] = (inputs[247]) & (inputs[199]);
    assign layer0_outputs[947] = ~((inputs[115]) ^ (inputs[251]));
    assign layer0_outputs[948] = (inputs[27]) & ~(inputs[55]);
    assign layer0_outputs[949] = ~(inputs[167]);
    assign layer0_outputs[950] = inputs[193];
    assign layer0_outputs[951] = inputs[158];
    assign layer0_outputs[952] = inputs[216];
    assign layer0_outputs[953] = 1'b0;
    assign layer0_outputs[954] = 1'b1;
    assign layer0_outputs[955] = ~((inputs[178]) ^ (inputs[103]));
    assign layer0_outputs[956] = inputs[137];
    assign layer0_outputs[957] = ~(inputs[186]) | (inputs[69]);
    assign layer0_outputs[958] = (inputs[186]) & (inputs[213]);
    assign layer0_outputs[959] = ~(inputs[33]);
    assign layer0_outputs[960] = 1'b0;
    assign layer0_outputs[961] = ~(inputs[108]) | (inputs[192]);
    assign layer0_outputs[962] = ~(inputs[164]);
    assign layer0_outputs[963] = inputs[65];
    assign layer0_outputs[964] = ~(inputs[118]) | (inputs[146]);
    assign layer0_outputs[965] = inputs[12];
    assign layer0_outputs[966] = 1'b1;
    assign layer0_outputs[967] = 1'b1;
    assign layer0_outputs[968] = ~(inputs[6]) | (inputs[149]);
    assign layer0_outputs[969] = (inputs[107]) | (inputs[227]);
    assign layer0_outputs[970] = 1'b1;
    assign layer0_outputs[971] = ~(inputs[7]);
    assign layer0_outputs[972] = (inputs[102]) | (inputs[109]);
    assign layer0_outputs[973] = 1'b1;
    assign layer0_outputs[974] = 1'b1;
    assign layer0_outputs[975] = (inputs[52]) & ~(inputs[227]);
    assign layer0_outputs[976] = (inputs[55]) & ~(inputs[69]);
    assign layer0_outputs[977] = (inputs[196]) ^ (inputs[11]);
    assign layer0_outputs[978] = ~((inputs[107]) ^ (inputs[180]));
    assign layer0_outputs[979] = (inputs[43]) & ~(inputs[19]);
    assign layer0_outputs[980] = 1'b0;
    assign layer0_outputs[981] = inputs[198];
    assign layer0_outputs[982] = 1'b0;
    assign layer0_outputs[983] = (inputs[111]) ^ (inputs[214]);
    assign layer0_outputs[984] = (inputs[137]) ^ (inputs[14]);
    assign layer0_outputs[985] = ~((inputs[45]) & (inputs[37]));
    assign layer0_outputs[986] = ~(inputs[238]) | (inputs[88]);
    assign layer0_outputs[987] = ~((inputs[88]) | (inputs[10]));
    assign layer0_outputs[988] = (inputs[79]) & ~(inputs[184]);
    assign layer0_outputs[989] = ~(inputs[185]) | (inputs[5]);
    assign layer0_outputs[990] = ~((inputs[227]) ^ (inputs[17]));
    assign layer0_outputs[991] = (inputs[207]) & ~(inputs[174]);
    assign layer0_outputs[992] = (inputs[5]) | (inputs[123]);
    assign layer0_outputs[993] = ~(inputs[53]);
    assign layer0_outputs[994] = inputs[9];
    assign layer0_outputs[995] = (inputs[1]) | (inputs[17]);
    assign layer0_outputs[996] = (inputs[24]) ^ (inputs[79]);
    assign layer0_outputs[997] = inputs[230];
    assign layer0_outputs[998] = ~((inputs[222]) ^ (inputs[100]));
    assign layer0_outputs[999] = ~(inputs[6]);
    assign layer0_outputs[1000] = ~(inputs[228]) | (inputs[164]);
    assign layer0_outputs[1001] = (inputs[52]) | (inputs[1]);
    assign layer0_outputs[1002] = ~(inputs[214]) | (inputs[92]);
    assign layer0_outputs[1003] = ~(inputs[194]);
    assign layer0_outputs[1004] = (inputs[36]) | (inputs[137]);
    assign layer0_outputs[1005] = inputs[119];
    assign layer0_outputs[1006] = ~(inputs[170]) | (inputs[25]);
    assign layer0_outputs[1007] = (inputs[74]) & ~(inputs[219]);
    assign layer0_outputs[1008] = ~((inputs[129]) & (inputs[166]));
    assign layer0_outputs[1009] = ~(inputs[63]) | (inputs[46]);
    assign layer0_outputs[1010] = ~(inputs[10]) | (inputs[172]);
    assign layer0_outputs[1011] = ~((inputs[57]) | (inputs[171]));
    assign layer0_outputs[1012] = (inputs[42]) & ~(inputs[46]);
    assign layer0_outputs[1013] = (inputs[224]) ^ (inputs[60]);
    assign layer0_outputs[1014] = (inputs[213]) & ~(inputs[22]);
    assign layer0_outputs[1015] = 1'b1;
    assign layer0_outputs[1016] = (inputs[151]) | (inputs[219]);
    assign layer0_outputs[1017] = ~((inputs[53]) ^ (inputs[94]));
    assign layer0_outputs[1018] = (inputs[81]) & ~(inputs[55]);
    assign layer0_outputs[1019] = ~((inputs[63]) ^ (inputs[172]));
    assign layer0_outputs[1020] = (inputs[205]) & (inputs[172]);
    assign layer0_outputs[1021] = (inputs[172]) & ~(inputs[15]);
    assign layer0_outputs[1022] = (inputs[246]) & ~(inputs[24]);
    assign layer0_outputs[1023] = inputs[33];
    assign layer0_outputs[1024] = 1'b0;
    assign layer0_outputs[1025] = ~(inputs[219]);
    assign layer0_outputs[1026] = ~(inputs[128]);
    assign layer0_outputs[1027] = ~(inputs[81]);
    assign layer0_outputs[1028] = inputs[88];
    assign layer0_outputs[1029] = (inputs[193]) ^ (inputs[106]);
    assign layer0_outputs[1030] = 1'b0;
    assign layer0_outputs[1031] = (inputs[37]) & ~(inputs[60]);
    assign layer0_outputs[1032] = 1'b1;
    assign layer0_outputs[1033] = inputs[144];
    assign layer0_outputs[1034] = (inputs[32]) ^ (inputs[133]);
    assign layer0_outputs[1035] = ~(inputs[192]) | (inputs[38]);
    assign layer0_outputs[1036] = inputs[56];
    assign layer0_outputs[1037] = inputs[70];
    assign layer0_outputs[1038] = (inputs[207]) & ~(inputs[121]);
    assign layer0_outputs[1039] = (inputs[161]) | (inputs[162]);
    assign layer0_outputs[1040] = ~(inputs[220]);
    assign layer0_outputs[1041] = (inputs[32]) | (inputs[105]);
    assign layer0_outputs[1042] = inputs[25];
    assign layer0_outputs[1043] = (inputs[70]) & ~(inputs[240]);
    assign layer0_outputs[1044] = ~(inputs[18]) | (inputs[201]);
    assign layer0_outputs[1045] = (inputs[95]) & ~(inputs[251]);
    assign layer0_outputs[1046] = (inputs[229]) & ~(inputs[34]);
    assign layer0_outputs[1047] = inputs[205];
    assign layer0_outputs[1048] = 1'b1;
    assign layer0_outputs[1049] = 1'b0;
    assign layer0_outputs[1050] = 1'b1;
    assign layer0_outputs[1051] = inputs[242];
    assign layer0_outputs[1052] = (inputs[77]) | (inputs[102]);
    assign layer0_outputs[1053] = 1'b0;
    assign layer0_outputs[1054] = 1'b0;
    assign layer0_outputs[1055] = ~((inputs[40]) ^ (inputs[199]));
    assign layer0_outputs[1056] = ~(inputs[145]);
    assign layer0_outputs[1057] = (inputs[166]) & (inputs[171]);
    assign layer0_outputs[1058] = 1'b0;
    assign layer0_outputs[1059] = ~(inputs[234]) | (inputs[29]);
    assign layer0_outputs[1060] = ~(inputs[168]);
    assign layer0_outputs[1061] = ~(inputs[36]);
    assign layer0_outputs[1062] = (inputs[69]) ^ (inputs[9]);
    assign layer0_outputs[1063] = 1'b0;
    assign layer0_outputs[1064] = 1'b0;
    assign layer0_outputs[1065] = ~((inputs[201]) ^ (inputs[138]));
    assign layer0_outputs[1066] = inputs[136];
    assign layer0_outputs[1067] = inputs[151];
    assign layer0_outputs[1068] = ~(inputs[151]) | (inputs[206]);
    assign layer0_outputs[1069] = (inputs[86]) ^ (inputs[208]);
    assign layer0_outputs[1070] = ~(inputs[216]) | (inputs[45]);
    assign layer0_outputs[1071] = ~(inputs[99]);
    assign layer0_outputs[1072] = ~(inputs[72]) | (inputs[136]);
    assign layer0_outputs[1073] = inputs[65];
    assign layer0_outputs[1074] = (inputs[89]) & (inputs[48]);
    assign layer0_outputs[1075] = ~(inputs[13]) | (inputs[203]);
    assign layer0_outputs[1076] = (inputs[160]) & (inputs[230]);
    assign layer0_outputs[1077] = ~((inputs[43]) ^ (inputs[35]));
    assign layer0_outputs[1078] = ~(inputs[97]) | (inputs[182]);
    assign layer0_outputs[1079] = ~((inputs[55]) & (inputs[74]));
    assign layer0_outputs[1080] = (inputs[121]) & ~(inputs[182]);
    assign layer0_outputs[1081] = (inputs[7]) & ~(inputs[223]);
    assign layer0_outputs[1082] = ~((inputs[64]) | (inputs[128]));
    assign layer0_outputs[1083] = inputs[101];
    assign layer0_outputs[1084] = (inputs[255]) & (inputs[93]);
    assign layer0_outputs[1085] = (inputs[122]) & (inputs[18]);
    assign layer0_outputs[1086] = ~((inputs[251]) | (inputs[163]));
    assign layer0_outputs[1087] = (inputs[17]) & ~(inputs[76]);
    assign layer0_outputs[1088] = (inputs[200]) & (inputs[183]);
    assign layer0_outputs[1089] = inputs[211];
    assign layer0_outputs[1090] = ~(inputs[25]) | (inputs[144]);
    assign layer0_outputs[1091] = (inputs[133]) ^ (inputs[251]);
    assign layer0_outputs[1092] = inputs[169];
    assign layer0_outputs[1093] = ~((inputs[109]) ^ (inputs[241]));
    assign layer0_outputs[1094] = 1'b1;
    assign layer0_outputs[1095] = (inputs[21]) & (inputs[90]);
    assign layer0_outputs[1096] = (inputs[252]) & ~(inputs[6]);
    assign layer0_outputs[1097] = inputs[29];
    assign layer0_outputs[1098] = (inputs[47]) & ~(inputs[33]);
    assign layer0_outputs[1099] = inputs[252];
    assign layer0_outputs[1100] = (inputs[166]) & ~(inputs[163]);
    assign layer0_outputs[1101] = (inputs[206]) | (inputs[188]);
    assign layer0_outputs[1102] = (inputs[56]) | (inputs[148]);
    assign layer0_outputs[1103] = ~((inputs[255]) & (inputs[210]));
    assign layer0_outputs[1104] = ~(inputs[129]);
    assign layer0_outputs[1105] = ~((inputs[167]) | (inputs[6]));
    assign layer0_outputs[1106] = (inputs[25]) & (inputs[58]);
    assign layer0_outputs[1107] = ~(inputs[41]) | (inputs[85]);
    assign layer0_outputs[1108] = ~(inputs[114]) | (inputs[243]);
    assign layer0_outputs[1109] = ~((inputs[80]) ^ (inputs[85]));
    assign layer0_outputs[1110] = ~(inputs[157]);
    assign layer0_outputs[1111] = 1'b1;
    assign layer0_outputs[1112] = (inputs[44]) & (inputs[234]);
    assign layer0_outputs[1113] = ~((inputs[220]) | (inputs[80]));
    assign layer0_outputs[1114] = ~(inputs[176]);
    assign layer0_outputs[1115] = inputs[143];
    assign layer0_outputs[1116] = (inputs[134]) ^ (inputs[207]);
    assign layer0_outputs[1117] = ~(inputs[247]);
    assign layer0_outputs[1118] = (inputs[208]) & ~(inputs[228]);
    assign layer0_outputs[1119] = ~((inputs[207]) | (inputs[28]));
    assign layer0_outputs[1120] = (inputs[92]) & ~(inputs[229]);
    assign layer0_outputs[1121] = inputs[23];
    assign layer0_outputs[1122] = (inputs[177]) ^ (inputs[105]);
    assign layer0_outputs[1123] = ~(inputs[157]) | (inputs[73]);
    assign layer0_outputs[1124] = ~(inputs[102]) | (inputs[152]);
    assign layer0_outputs[1125] = ~(inputs[132]) | (inputs[236]);
    assign layer0_outputs[1126] = ~(inputs[27]);
    assign layer0_outputs[1127] = inputs[27];
    assign layer0_outputs[1128] = 1'b0;
    assign layer0_outputs[1129] = ~((inputs[171]) | (inputs[202]));
    assign layer0_outputs[1130] = inputs[181];
    assign layer0_outputs[1131] = ~(inputs[127]);
    assign layer0_outputs[1132] = 1'b0;
    assign layer0_outputs[1133] = inputs[164];
    assign layer0_outputs[1134] = (inputs[149]) | (inputs[174]);
    assign layer0_outputs[1135] = ~((inputs[55]) & (inputs[55]));
    assign layer0_outputs[1136] = (inputs[134]) & ~(inputs[36]);
    assign layer0_outputs[1137] = (inputs[67]) & ~(inputs[196]);
    assign layer0_outputs[1138] = ~((inputs[178]) & (inputs[150]));
    assign layer0_outputs[1139] = 1'b0;
    assign layer0_outputs[1140] = ~(inputs[151]) | (inputs[144]);
    assign layer0_outputs[1141] = 1'b0;
    assign layer0_outputs[1142] = (inputs[35]) ^ (inputs[68]);
    assign layer0_outputs[1143] = (inputs[48]) & (inputs[41]);
    assign layer0_outputs[1144] = (inputs[117]) & ~(inputs[114]);
    assign layer0_outputs[1145] = ~(inputs[44]) | (inputs[90]);
    assign layer0_outputs[1146] = 1'b0;
    assign layer0_outputs[1147] = (inputs[143]) | (inputs[150]);
    assign layer0_outputs[1148] = 1'b1;
    assign layer0_outputs[1149] = ~(inputs[217]) | (inputs[29]);
    assign layer0_outputs[1150] = (inputs[121]) & ~(inputs[180]);
    assign layer0_outputs[1151] = 1'b0;
    assign layer0_outputs[1152] = ~((inputs[49]) ^ (inputs[172]));
    assign layer0_outputs[1153] = (inputs[151]) & ~(inputs[82]);
    assign layer0_outputs[1154] = (inputs[128]) & (inputs[4]);
    assign layer0_outputs[1155] = ~(inputs[189]);
    assign layer0_outputs[1156] = (inputs[57]) | (inputs[93]);
    assign layer0_outputs[1157] = inputs[43];
    assign layer0_outputs[1158] = 1'b0;
    assign layer0_outputs[1159] = ~((inputs[152]) & (inputs[137]));
    assign layer0_outputs[1160] = ~(inputs[223]);
    assign layer0_outputs[1161] = ~((inputs[62]) ^ (inputs[244]));
    assign layer0_outputs[1162] = ~(inputs[29]);
    assign layer0_outputs[1163] = inputs[149];
    assign layer0_outputs[1164] = ~(inputs[202]) | (inputs[99]);
    assign layer0_outputs[1165] = ~((inputs[41]) | (inputs[51]));
    assign layer0_outputs[1166] = ~(inputs[250]) | (inputs[5]);
    assign layer0_outputs[1167] = inputs[74];
    assign layer0_outputs[1168] = (inputs[12]) | (inputs[215]);
    assign layer0_outputs[1169] = inputs[169];
    assign layer0_outputs[1170] = (inputs[137]) & ~(inputs[38]);
    assign layer0_outputs[1171] = ~(inputs[188]) | (inputs[81]);
    assign layer0_outputs[1172] = (inputs[242]) & ~(inputs[187]);
    assign layer0_outputs[1173] = ~((inputs[80]) & (inputs[114]));
    assign layer0_outputs[1174] = ~(inputs[161]) | (inputs[253]);
    assign layer0_outputs[1175] = ~(inputs[45]) | (inputs[122]);
    assign layer0_outputs[1176] = ~((inputs[3]) & (inputs[23]));
    assign layer0_outputs[1177] = ~((inputs[192]) ^ (inputs[51]));
    assign layer0_outputs[1178] = ~(inputs[88]);
    assign layer0_outputs[1179] = ~((inputs[205]) & (inputs[157]));
    assign layer0_outputs[1180] = 1'b1;
    assign layer0_outputs[1181] = (inputs[173]) | (inputs[43]);
    assign layer0_outputs[1182] = ~(inputs[185]) | (inputs[35]);
    assign layer0_outputs[1183] = (inputs[66]) | (inputs[181]);
    assign layer0_outputs[1184] = 1'b0;
    assign layer0_outputs[1185] = 1'b1;
    assign layer0_outputs[1186] = ~(inputs[207]);
    assign layer0_outputs[1187] = (inputs[114]) & ~(inputs[70]);
    assign layer0_outputs[1188] = 1'b0;
    assign layer0_outputs[1189] = (inputs[96]) | (inputs[30]);
    assign layer0_outputs[1190] = inputs[145];
    assign layer0_outputs[1191] = (inputs[104]) & ~(inputs[81]);
    assign layer0_outputs[1192] = 1'b0;
    assign layer0_outputs[1193] = ~(inputs[224]) | (inputs[2]);
    assign layer0_outputs[1194] = inputs[53];
    assign layer0_outputs[1195] = ~((inputs[253]) ^ (inputs[145]));
    assign layer0_outputs[1196] = ~(inputs[222]);
    assign layer0_outputs[1197] = (inputs[159]) ^ (inputs[199]);
    assign layer0_outputs[1198] = (inputs[115]) & ~(inputs[20]);
    assign layer0_outputs[1199] = (inputs[105]) | (inputs[97]);
    assign layer0_outputs[1200] = ~(inputs[150]);
    assign layer0_outputs[1201] = ~(inputs[51]);
    assign layer0_outputs[1202] = (inputs[37]) & ~(inputs[92]);
    assign layer0_outputs[1203] = (inputs[215]) | (inputs[101]);
    assign layer0_outputs[1204] = ~(inputs[69]);
    assign layer0_outputs[1205] = 1'b1;
    assign layer0_outputs[1206] = ~((inputs[232]) ^ (inputs[9]));
    assign layer0_outputs[1207] = inputs[102];
    assign layer0_outputs[1208] = ~((inputs[20]) ^ (inputs[38]));
    assign layer0_outputs[1209] = ~((inputs[39]) | (inputs[165]));
    assign layer0_outputs[1210] = ~(inputs[194]);
    assign layer0_outputs[1211] = (inputs[148]) | (inputs[25]);
    assign layer0_outputs[1212] = 1'b1;
    assign layer0_outputs[1213] = ~(inputs[102]);
    assign layer0_outputs[1214] = inputs[172];
    assign layer0_outputs[1215] = inputs[157];
    assign layer0_outputs[1216] = ~((inputs[242]) ^ (inputs[33]));
    assign layer0_outputs[1217] = (inputs[200]) ^ (inputs[249]);
    assign layer0_outputs[1218] = (inputs[169]) | (inputs[92]);
    assign layer0_outputs[1219] = ~(inputs[205]);
    assign layer0_outputs[1220] = ~(inputs[193]);
    assign layer0_outputs[1221] = (inputs[166]) & ~(inputs[44]);
    assign layer0_outputs[1222] = (inputs[130]) & ~(inputs[156]);
    assign layer0_outputs[1223] = (inputs[127]) ^ (inputs[210]);
    assign layer0_outputs[1224] = ~((inputs[213]) & (inputs[175]));
    assign layer0_outputs[1225] = (inputs[59]) & ~(inputs[233]);
    assign layer0_outputs[1226] = (inputs[188]) & ~(inputs[24]);
    assign layer0_outputs[1227] = ~((inputs[132]) | (inputs[118]));
    assign layer0_outputs[1228] = 1'b1;
    assign layer0_outputs[1229] = ~((inputs[151]) | (inputs[253]));
    assign layer0_outputs[1230] = (inputs[210]) | (inputs[63]);
    assign layer0_outputs[1231] = inputs[108];
    assign layer0_outputs[1232] = ~((inputs[253]) | (inputs[5]));
    assign layer0_outputs[1233] = ~(inputs[102]);
    assign layer0_outputs[1234] = (inputs[228]) & ~(inputs[251]);
    assign layer0_outputs[1235] = inputs[131];
    assign layer0_outputs[1236] = (inputs[249]) & (inputs[35]);
    assign layer0_outputs[1237] = (inputs[207]) & (inputs[224]);
    assign layer0_outputs[1238] = inputs[21];
    assign layer0_outputs[1239] = (inputs[100]) | (inputs[19]);
    assign layer0_outputs[1240] = ~((inputs[57]) & (inputs[203]));
    assign layer0_outputs[1241] = ~(inputs[79]) | (inputs[97]);
    assign layer0_outputs[1242] = (inputs[53]) & ~(inputs[146]);
    assign layer0_outputs[1243] = inputs[63];
    assign layer0_outputs[1244] = inputs[229];
    assign layer0_outputs[1245] = ~((inputs[167]) | (inputs[223]));
    assign layer0_outputs[1246] = (inputs[142]) | (inputs[21]);
    assign layer0_outputs[1247] = inputs[170];
    assign layer0_outputs[1248] = ~((inputs[82]) ^ (inputs[184]));
    assign layer0_outputs[1249] = 1'b1;
    assign layer0_outputs[1250] = ~(inputs[121]) | (inputs[166]);
    assign layer0_outputs[1251] = ~(inputs[128]);
    assign layer0_outputs[1252] = ~((inputs[93]) | (inputs[159]));
    assign layer0_outputs[1253] = ~((inputs[130]) ^ (inputs[116]));
    assign layer0_outputs[1254] = (inputs[74]) | (inputs[162]);
    assign layer0_outputs[1255] = inputs[240];
    assign layer0_outputs[1256] = (inputs[129]) & (inputs[170]);
    assign layer0_outputs[1257] = ~((inputs[177]) ^ (inputs[122]));
    assign layer0_outputs[1258] = 1'b0;
    assign layer0_outputs[1259] = ~(inputs[26]);
    assign layer0_outputs[1260] = ~(inputs[63]);
    assign layer0_outputs[1261] = inputs[68];
    assign layer0_outputs[1262] = (inputs[138]) & ~(inputs[225]);
    assign layer0_outputs[1263] = ~(inputs[232]) | (inputs[43]);
    assign layer0_outputs[1264] = (inputs[242]) & ~(inputs[235]);
    assign layer0_outputs[1265] = ~((inputs[169]) & (inputs[108]));
    assign layer0_outputs[1266] = inputs[44];
    assign layer0_outputs[1267] = (inputs[254]) & (inputs[36]);
    assign layer0_outputs[1268] = (inputs[130]) & ~(inputs[173]);
    assign layer0_outputs[1269] = (inputs[245]) & ~(inputs[183]);
    assign layer0_outputs[1270] = (inputs[192]) & ~(inputs[176]);
    assign layer0_outputs[1271] = ~(inputs[56]) | (inputs[114]);
    assign layer0_outputs[1272] = ~(inputs[190]);
    assign layer0_outputs[1273] = (inputs[205]) & (inputs[143]);
    assign layer0_outputs[1274] = ~((inputs[101]) | (inputs[117]));
    assign layer0_outputs[1275] = 1'b1;
    assign layer0_outputs[1276] = ~((inputs[89]) ^ (inputs[251]));
    assign layer0_outputs[1277] = ~(inputs[5]);
    assign layer0_outputs[1278] = 1'b1;
    assign layer0_outputs[1279] = (inputs[219]) | (inputs[122]);
    assign layer0_outputs[1280] = (inputs[2]) & (inputs[228]);
    assign layer0_outputs[1281] = (inputs[118]) & ~(inputs[225]);
    assign layer0_outputs[1282] = ~(inputs[208]);
    assign layer0_outputs[1283] = ~((inputs[127]) & (inputs[81]));
    assign layer0_outputs[1284] = (inputs[27]) & ~(inputs[196]);
    assign layer0_outputs[1285] = ~((inputs[208]) & (inputs[184]));
    assign layer0_outputs[1286] = (inputs[182]) ^ (inputs[80]);
    assign layer0_outputs[1287] = (inputs[81]) & ~(inputs[39]);
    assign layer0_outputs[1288] = ~(inputs[12]) | (inputs[85]);
    assign layer0_outputs[1289] = 1'b0;
    assign layer0_outputs[1290] = 1'b0;
    assign layer0_outputs[1291] = inputs[88];
    assign layer0_outputs[1292] = inputs[146];
    assign layer0_outputs[1293] = (inputs[39]) & ~(inputs[245]);
    assign layer0_outputs[1294] = ~((inputs[207]) ^ (inputs[29]));
    assign layer0_outputs[1295] = 1'b1;
    assign layer0_outputs[1296] = inputs[85];
    assign layer0_outputs[1297] = (inputs[22]) | (inputs[201]);
    assign layer0_outputs[1298] = ~(inputs[117]) | (inputs[159]);
    assign layer0_outputs[1299] = (inputs[33]) | (inputs[104]);
    assign layer0_outputs[1300] = ~(inputs[40]);
    assign layer0_outputs[1301] = ~(inputs[51]);
    assign layer0_outputs[1302] = (inputs[70]) | (inputs[215]);
    assign layer0_outputs[1303] = 1'b0;
    assign layer0_outputs[1304] = inputs[21];
    assign layer0_outputs[1305] = ~(inputs[148]) | (inputs[86]);
    assign layer0_outputs[1306] = ~(inputs[149]) | (inputs[37]);
    assign layer0_outputs[1307] = (inputs[102]) ^ (inputs[235]);
    assign layer0_outputs[1308] = ~((inputs[251]) & (inputs[141]));
    assign layer0_outputs[1309] = ~(inputs[29]);
    assign layer0_outputs[1310] = inputs[61];
    assign layer0_outputs[1311] = (inputs[204]) | (inputs[101]);
    assign layer0_outputs[1312] = 1'b0;
    assign layer0_outputs[1313] = ~((inputs[210]) ^ (inputs[175]));
    assign layer0_outputs[1314] = inputs[151];
    assign layer0_outputs[1315] = ~((inputs[113]) & (inputs[58]));
    assign layer0_outputs[1316] = (inputs[233]) ^ (inputs[208]);
    assign layer0_outputs[1317] = ~(inputs[124]) | (inputs[160]);
    assign layer0_outputs[1318] = ~((inputs[215]) & (inputs[193]));
    assign layer0_outputs[1319] = ~((inputs[201]) ^ (inputs[247]));
    assign layer0_outputs[1320] = ~((inputs[177]) | (inputs[118]));
    assign layer0_outputs[1321] = (inputs[252]) | (inputs[73]);
    assign layer0_outputs[1322] = 1'b0;
    assign layer0_outputs[1323] = inputs[58];
    assign layer0_outputs[1324] = (inputs[225]) & ~(inputs[171]);
    assign layer0_outputs[1325] = ~((inputs[91]) | (inputs[30]));
    assign layer0_outputs[1326] = inputs[136];
    assign layer0_outputs[1327] = ~(inputs[94]);
    assign layer0_outputs[1328] = ~(inputs[72]) | (inputs[143]);
    assign layer0_outputs[1329] = 1'b1;
    assign layer0_outputs[1330] = (inputs[208]) & ~(inputs[175]);
    assign layer0_outputs[1331] = inputs[138];
    assign layer0_outputs[1332] = (inputs[183]) & (inputs[10]);
    assign layer0_outputs[1333] = (inputs[118]) & (inputs[34]);
    assign layer0_outputs[1334] = ~(inputs[161]) | (inputs[67]);
    assign layer0_outputs[1335] = (inputs[6]) & (inputs[180]);
    assign layer0_outputs[1336] = 1'b0;
    assign layer0_outputs[1337] = ~((inputs[176]) ^ (inputs[119]));
    assign layer0_outputs[1338] = ~(inputs[98]);
    assign layer0_outputs[1339] = ~(inputs[239]) | (inputs[176]);
    assign layer0_outputs[1340] = ~((inputs[158]) & (inputs[255]));
    assign layer0_outputs[1341] = ~((inputs[143]) ^ (inputs[2]));
    assign layer0_outputs[1342] = ~(inputs[156]);
    assign layer0_outputs[1343] = (inputs[158]) & ~(inputs[127]);
    assign layer0_outputs[1344] = ~((inputs[174]) & (inputs[21]));
    assign layer0_outputs[1345] = inputs[252];
    assign layer0_outputs[1346] = (inputs[58]) & (inputs[32]);
    assign layer0_outputs[1347] = (inputs[143]) | (inputs[54]);
    assign layer0_outputs[1348] = (inputs[188]) & ~(inputs[28]);
    assign layer0_outputs[1349] = (inputs[172]) & (inputs[196]);
    assign layer0_outputs[1350] = ~(inputs[94]) | (inputs[246]);
    assign layer0_outputs[1351] = 1'b1;
    assign layer0_outputs[1352] = ~((inputs[137]) | (inputs[21]));
    assign layer0_outputs[1353] = inputs[34];
    assign layer0_outputs[1354] = (inputs[198]) & ~(inputs[220]);
    assign layer0_outputs[1355] = 1'b1;
    assign layer0_outputs[1356] = ~(inputs[206]);
    assign layer0_outputs[1357] = ~(inputs[71]);
    assign layer0_outputs[1358] = ~((inputs[23]) ^ (inputs[236]));
    assign layer0_outputs[1359] = 1'b1;
    assign layer0_outputs[1360] = ~((inputs[204]) ^ (inputs[135]));
    assign layer0_outputs[1361] = 1'b1;
    assign layer0_outputs[1362] = (inputs[200]) | (inputs[176]);
    assign layer0_outputs[1363] = inputs[126];
    assign layer0_outputs[1364] = 1'b1;
    assign layer0_outputs[1365] = 1'b0;
    assign layer0_outputs[1366] = (inputs[226]) & ~(inputs[30]);
    assign layer0_outputs[1367] = ~(inputs[153]);
    assign layer0_outputs[1368] = inputs[105];
    assign layer0_outputs[1369] = inputs[238];
    assign layer0_outputs[1370] = ~((inputs[74]) | (inputs[181]));
    assign layer0_outputs[1371] = inputs[184];
    assign layer0_outputs[1372] = ~((inputs[178]) | (inputs[180]));
    assign layer0_outputs[1373] = (inputs[120]) & ~(inputs[18]);
    assign layer0_outputs[1374] = (inputs[208]) & ~(inputs[144]);
    assign layer0_outputs[1375] = ~((inputs[21]) ^ (inputs[58]));
    assign layer0_outputs[1376] = inputs[5];
    assign layer0_outputs[1377] = ~((inputs[128]) & (inputs[166]));
    assign layer0_outputs[1378] = ~((inputs[137]) | (inputs[137]));
    assign layer0_outputs[1379] = (inputs[108]) & (inputs[108]);
    assign layer0_outputs[1380] = (inputs[62]) & ~(inputs[101]);
    assign layer0_outputs[1381] = (inputs[3]) & ~(inputs[150]);
    assign layer0_outputs[1382] = ~(inputs[116]);
    assign layer0_outputs[1383] = ~(inputs[237]);
    assign layer0_outputs[1384] = 1'b1;
    assign layer0_outputs[1385] = 1'b1;
    assign layer0_outputs[1386] = ~((inputs[45]) | (inputs[211]));
    assign layer0_outputs[1387] = 1'b1;
    assign layer0_outputs[1388] = ~((inputs[160]) | (inputs[161]));
    assign layer0_outputs[1389] = 1'b1;
    assign layer0_outputs[1390] = ~(inputs[246]);
    assign layer0_outputs[1391] = ~(inputs[158]);
    assign layer0_outputs[1392] = (inputs[40]) & ~(inputs[97]);
    assign layer0_outputs[1393] = ~((inputs[152]) | (inputs[222]));
    assign layer0_outputs[1394] = ~(inputs[235]) | (inputs[51]);
    assign layer0_outputs[1395] = ~(inputs[159]);
    assign layer0_outputs[1396] = 1'b0;
    assign layer0_outputs[1397] = ~(inputs[14]) | (inputs[10]);
    assign layer0_outputs[1398] = inputs[136];
    assign layer0_outputs[1399] = inputs[60];
    assign layer0_outputs[1400] = ~((inputs[232]) & (inputs[244]));
    assign layer0_outputs[1401] = (inputs[56]) & (inputs[236]);
    assign layer0_outputs[1402] = ~(inputs[221]) | (inputs[151]);
    assign layer0_outputs[1403] = ~((inputs[236]) | (inputs[242]));
    assign layer0_outputs[1404] = 1'b1;
    assign layer0_outputs[1405] = ~((inputs[192]) | (inputs[250]));
    assign layer0_outputs[1406] = (inputs[215]) & (inputs[25]);
    assign layer0_outputs[1407] = inputs[142];
    assign layer0_outputs[1408] = ~(inputs[198]) | (inputs[139]);
    assign layer0_outputs[1409] = ~((inputs[182]) | (inputs[197]));
    assign layer0_outputs[1410] = 1'b0;
    assign layer0_outputs[1411] = 1'b1;
    assign layer0_outputs[1412] = ~((inputs[210]) ^ (inputs[61]));
    assign layer0_outputs[1413] = (inputs[113]) | (inputs[13]);
    assign layer0_outputs[1414] = ~((inputs[52]) | (inputs[138]));
    assign layer0_outputs[1415] = ~((inputs[160]) & (inputs[218]));
    assign layer0_outputs[1416] = 1'b0;
    assign layer0_outputs[1417] = (inputs[168]) & ~(inputs[252]);
    assign layer0_outputs[1418] = inputs[245];
    assign layer0_outputs[1419] = ~(inputs[132]);
    assign layer0_outputs[1420] = (inputs[147]) ^ (inputs[94]);
    assign layer0_outputs[1421] = inputs[64];
    assign layer0_outputs[1422] = (inputs[149]) & ~(inputs[43]);
    assign layer0_outputs[1423] = ~(inputs[49]);
    assign layer0_outputs[1424] = ~((inputs[203]) ^ (inputs[29]));
    assign layer0_outputs[1425] = (inputs[125]) | (inputs[87]);
    assign layer0_outputs[1426] = (inputs[193]) & ~(inputs[72]);
    assign layer0_outputs[1427] = (inputs[101]) | (inputs[106]);
    assign layer0_outputs[1428] = ~(inputs[31]) | (inputs[138]);
    assign layer0_outputs[1429] = 1'b1;
    assign layer0_outputs[1430] = ~((inputs[12]) ^ (inputs[86]));
    assign layer0_outputs[1431] = 1'b1;
    assign layer0_outputs[1432] = ~((inputs[21]) | (inputs[170]));
    assign layer0_outputs[1433] = inputs[66];
    assign layer0_outputs[1434] = (inputs[252]) | (inputs[208]);
    assign layer0_outputs[1435] = (inputs[172]) | (inputs[202]);
    assign layer0_outputs[1436] = (inputs[16]) & ~(inputs[21]);
    assign layer0_outputs[1437] = (inputs[105]) & ~(inputs[8]);
    assign layer0_outputs[1438] = (inputs[205]) & ~(inputs[140]);
    assign layer0_outputs[1439] = (inputs[92]) ^ (inputs[61]);
    assign layer0_outputs[1440] = 1'b1;
    assign layer0_outputs[1441] = (inputs[46]) ^ (inputs[188]);
    assign layer0_outputs[1442] = inputs[75];
    assign layer0_outputs[1443] = ~((inputs[30]) & (inputs[70]));
    assign layer0_outputs[1444] = inputs[120];
    assign layer0_outputs[1445] = 1'b0;
    assign layer0_outputs[1446] = (inputs[45]) & ~(inputs[13]);
    assign layer0_outputs[1447] = ~((inputs[40]) | (inputs[210]));
    assign layer0_outputs[1448] = 1'b1;
    assign layer0_outputs[1449] = (inputs[176]) ^ (inputs[52]);
    assign layer0_outputs[1450] = ~((inputs[150]) ^ (inputs[223]));
    assign layer0_outputs[1451] = 1'b1;
    assign layer0_outputs[1452] = ~(inputs[248]);
    assign layer0_outputs[1453] = (inputs[92]) | (inputs[11]);
    assign layer0_outputs[1454] = (inputs[48]) & (inputs[107]);
    assign layer0_outputs[1455] = (inputs[87]) | (inputs[93]);
    assign layer0_outputs[1456] = (inputs[39]) & ~(inputs[134]);
    assign layer0_outputs[1457] = inputs[68];
    assign layer0_outputs[1458] = inputs[105];
    assign layer0_outputs[1459] = (inputs[117]) & (inputs[105]);
    assign layer0_outputs[1460] = (inputs[186]) & ~(inputs[243]);
    assign layer0_outputs[1461] = ~(inputs[69]);
    assign layer0_outputs[1462] = ~(inputs[14]);
    assign layer0_outputs[1463] = inputs[39];
    assign layer0_outputs[1464] = 1'b0;
    assign layer0_outputs[1465] = ~((inputs[247]) & (inputs[78]));
    assign layer0_outputs[1466] = ~((inputs[154]) | (inputs[195]));
    assign layer0_outputs[1467] = inputs[158];
    assign layer0_outputs[1468] = ~((inputs[161]) ^ (inputs[15]));
    assign layer0_outputs[1469] = ~((inputs[26]) | (inputs[140]));
    assign layer0_outputs[1470] = (inputs[102]) ^ (inputs[65]);
    assign layer0_outputs[1471] = ~(inputs[120]) | (inputs[23]);
    assign layer0_outputs[1472] = ~((inputs[191]) | (inputs[27]));
    assign layer0_outputs[1473] = (inputs[47]) ^ (inputs[187]);
    assign layer0_outputs[1474] = ~(inputs[124]);
    assign layer0_outputs[1475] = 1'b0;
    assign layer0_outputs[1476] = ~(inputs[79]) | (inputs[174]);
    assign layer0_outputs[1477] = (inputs[127]) & ~(inputs[163]);
    assign layer0_outputs[1478] = 1'b0;
    assign layer0_outputs[1479] = (inputs[55]) & (inputs[246]);
    assign layer0_outputs[1480] = inputs[148];
    assign layer0_outputs[1481] = (inputs[202]) ^ (inputs[130]);
    assign layer0_outputs[1482] = ~(inputs[27]);
    assign layer0_outputs[1483] = inputs[4];
    assign layer0_outputs[1484] = ~(inputs[78]) | (inputs[47]);
    assign layer0_outputs[1485] = ~(inputs[141]);
    assign layer0_outputs[1486] = (inputs[211]) | (inputs[134]);
    assign layer0_outputs[1487] = ~(inputs[177]);
    assign layer0_outputs[1488] = (inputs[129]) & ~(inputs[77]);
    assign layer0_outputs[1489] = ~(inputs[138]) | (inputs[178]);
    assign layer0_outputs[1490] = (inputs[1]) & (inputs[154]);
    assign layer0_outputs[1491] = ~((inputs[85]) | (inputs[229]));
    assign layer0_outputs[1492] = inputs[52];
    assign layer0_outputs[1493] = inputs[185];
    assign layer0_outputs[1494] = ~((inputs[126]) & (inputs[34]));
    assign layer0_outputs[1495] = 1'b1;
    assign layer0_outputs[1496] = 1'b0;
    assign layer0_outputs[1497] = 1'b0;
    assign layer0_outputs[1498] = inputs[61];
    assign layer0_outputs[1499] = (inputs[24]) & ~(inputs[243]);
    assign layer0_outputs[1500] = ~((inputs[107]) | (inputs[91]));
    assign layer0_outputs[1501] = 1'b1;
    assign layer0_outputs[1502] = ~(inputs[240]);
    assign layer0_outputs[1503] = (inputs[212]) & ~(inputs[176]);
    assign layer0_outputs[1504] = 1'b0;
    assign layer0_outputs[1505] = (inputs[122]) & ~(inputs[78]);
    assign layer0_outputs[1506] = 1'b1;
    assign layer0_outputs[1507] = ~((inputs[22]) | (inputs[209]));
    assign layer0_outputs[1508] = ~((inputs[17]) & (inputs[185]));
    assign layer0_outputs[1509] = (inputs[255]) & ~(inputs[4]);
    assign layer0_outputs[1510] = ~((inputs[159]) ^ (inputs[80]));
    assign layer0_outputs[1511] = ~((inputs[191]) & (inputs[113]));
    assign layer0_outputs[1512] = ~(inputs[99]) | (inputs[66]);
    assign layer0_outputs[1513] = inputs[68];
    assign layer0_outputs[1514] = inputs[116];
    assign layer0_outputs[1515] = ~(inputs[53]);
    assign layer0_outputs[1516] = (inputs[84]) & (inputs[79]);
    assign layer0_outputs[1517] = ~((inputs[19]) | (inputs[117]));
    assign layer0_outputs[1518] = ~((inputs[1]) ^ (inputs[177]));
    assign layer0_outputs[1519] = inputs[9];
    assign layer0_outputs[1520] = inputs[136];
    assign layer0_outputs[1521] = ~((inputs[29]) | (inputs[253]));
    assign layer0_outputs[1522] = ~(inputs[50]) | (inputs[30]);
    assign layer0_outputs[1523] = 1'b1;
    assign layer0_outputs[1524] = ~(inputs[7]);
    assign layer0_outputs[1525] = 1'b0;
    assign layer0_outputs[1526] = (inputs[186]) & ~(inputs[58]);
    assign layer0_outputs[1527] = ~(inputs[54]) | (inputs[110]);
    assign layer0_outputs[1528] = ~((inputs[220]) | (inputs[132]));
    assign layer0_outputs[1529] = 1'b1;
    assign layer0_outputs[1530] = (inputs[57]) | (inputs[244]);
    assign layer0_outputs[1531] = (inputs[49]) & (inputs[196]);
    assign layer0_outputs[1532] = inputs[48];
    assign layer0_outputs[1533] = (inputs[143]) & ~(inputs[36]);
    assign layer0_outputs[1534] = ~((inputs[222]) | (inputs[24]));
    assign layer0_outputs[1535] = ~((inputs[133]) & (inputs[167]));
    assign layer0_outputs[1536] = ~(inputs[132]);
    assign layer0_outputs[1537] = 1'b0;
    assign layer0_outputs[1538] = (inputs[254]) & (inputs[228]);
    assign layer0_outputs[1539] = (inputs[74]) ^ (inputs[73]);
    assign layer0_outputs[1540] = inputs[56];
    assign layer0_outputs[1541] = (inputs[117]) | (inputs[109]);
    assign layer0_outputs[1542] = (inputs[89]) & (inputs[64]);
    assign layer0_outputs[1543] = ~(inputs[144]);
    assign layer0_outputs[1544] = (inputs[234]) & (inputs[39]);
    assign layer0_outputs[1545] = (inputs[97]) & ~(inputs[2]);
    assign layer0_outputs[1546] = (inputs[255]) & (inputs[168]);
    assign layer0_outputs[1547] = (inputs[230]) | (inputs[224]);
    assign layer0_outputs[1548] = ~((inputs[116]) | (inputs[216]));
    assign layer0_outputs[1549] = inputs[109];
    assign layer0_outputs[1550] = ~(inputs[231]) | (inputs[177]);
    assign layer0_outputs[1551] = (inputs[185]) & ~(inputs[206]);
    assign layer0_outputs[1552] = ~((inputs[238]) | (inputs[105]));
    assign layer0_outputs[1553] = ~(inputs[6]);
    assign layer0_outputs[1554] = ~(inputs[90]);
    assign layer0_outputs[1555] = 1'b1;
    assign layer0_outputs[1556] = ~(inputs[10]);
    assign layer0_outputs[1557] = ~(inputs[41]) | (inputs[7]);
    assign layer0_outputs[1558] = 1'b1;
    assign layer0_outputs[1559] = 1'b1;
    assign layer0_outputs[1560] = ~((inputs[59]) ^ (inputs[72]));
    assign layer0_outputs[1561] = (inputs[245]) ^ (inputs[34]);
    assign layer0_outputs[1562] = 1'b1;
    assign layer0_outputs[1563] = (inputs[10]) & ~(inputs[26]);
    assign layer0_outputs[1564] = (inputs[120]) | (inputs[68]);
    assign layer0_outputs[1565] = ~(inputs[134]) | (inputs[59]);
    assign layer0_outputs[1566] = inputs[207];
    assign layer0_outputs[1567] = ~(inputs[169]);
    assign layer0_outputs[1568] = ~(inputs[52]);
    assign layer0_outputs[1569] = 1'b0;
    assign layer0_outputs[1570] = (inputs[189]) ^ (inputs[23]);
    assign layer0_outputs[1571] = ~((inputs[72]) | (inputs[35]));
    assign layer0_outputs[1572] = ~(inputs[179]) | (inputs[173]);
    assign layer0_outputs[1573] = ~(inputs[82]) | (inputs[11]);
    assign layer0_outputs[1574] = (inputs[63]) | (inputs[47]);
    assign layer0_outputs[1575] = ~((inputs[240]) & (inputs[249]));
    assign layer0_outputs[1576] = (inputs[112]) & (inputs[5]);
    assign layer0_outputs[1577] = ~(inputs[52]);
    assign layer0_outputs[1578] = (inputs[9]) & ~(inputs[80]);
    assign layer0_outputs[1579] = ~(inputs[15]) | (inputs[44]);
    assign layer0_outputs[1580] = inputs[189];
    assign layer0_outputs[1581] = (inputs[30]) & ~(inputs[112]);
    assign layer0_outputs[1582] = inputs[15];
    assign layer0_outputs[1583] = (inputs[167]) & ~(inputs[99]);
    assign layer0_outputs[1584] = 1'b1;
    assign layer0_outputs[1585] = 1'b0;
    assign layer0_outputs[1586] = ~(inputs[36]) | (inputs[65]);
    assign layer0_outputs[1587] = (inputs[195]) & ~(inputs[15]);
    assign layer0_outputs[1588] = (inputs[231]) & (inputs[95]);
    assign layer0_outputs[1589] = (inputs[63]) & ~(inputs[80]);
    assign layer0_outputs[1590] = ~(inputs[151]);
    assign layer0_outputs[1591] = inputs[214];
    assign layer0_outputs[1592] = 1'b0;
    assign layer0_outputs[1593] = inputs[214];
    assign layer0_outputs[1594] = (inputs[255]) & ~(inputs[144]);
    assign layer0_outputs[1595] = inputs[67];
    assign layer0_outputs[1596] = ~(inputs[148]) | (inputs[255]);
    assign layer0_outputs[1597] = ~((inputs[45]) | (inputs[192]));
    assign layer0_outputs[1598] = inputs[242];
    assign layer0_outputs[1599] = (inputs[167]) & ~(inputs[3]);
    assign layer0_outputs[1600] = ~(inputs[222]);
    assign layer0_outputs[1601] = ~((inputs[115]) & (inputs[203]));
    assign layer0_outputs[1602] = ~(inputs[139]) | (inputs[94]);
    assign layer0_outputs[1603] = 1'b0;
    assign layer0_outputs[1604] = ~((inputs[251]) ^ (inputs[171]));
    assign layer0_outputs[1605] = 1'b0;
    assign layer0_outputs[1606] = ~((inputs[123]) ^ (inputs[222]));
    assign layer0_outputs[1607] = 1'b0;
    assign layer0_outputs[1608] = ~((inputs[239]) & (inputs[96]));
    assign layer0_outputs[1609] = ~((inputs[33]) ^ (inputs[159]));
    assign layer0_outputs[1610] = 1'b1;
    assign layer0_outputs[1611] = 1'b1;
    assign layer0_outputs[1612] = ~((inputs[94]) ^ (inputs[166]));
    assign layer0_outputs[1613] = ~((inputs[150]) | (inputs[100]));
    assign layer0_outputs[1614] = (inputs[153]) | (inputs[35]);
    assign layer0_outputs[1615] = ~(inputs[152]);
    assign layer0_outputs[1616] = (inputs[216]) | (inputs[12]);
    assign layer0_outputs[1617] = ~(inputs[224]) | (inputs[104]);
    assign layer0_outputs[1618] = ~(inputs[211]);
    assign layer0_outputs[1619] = (inputs[152]) ^ (inputs[243]);
    assign layer0_outputs[1620] = 1'b1;
    assign layer0_outputs[1621] = (inputs[30]) ^ (inputs[7]);
    assign layer0_outputs[1622] = ~(inputs[236]);
    assign layer0_outputs[1623] = inputs[222];
    assign layer0_outputs[1624] = ~(inputs[40]) | (inputs[231]);
    assign layer0_outputs[1625] = ~((inputs[98]) | (inputs[137]));
    assign layer0_outputs[1626] = (inputs[94]) & ~(inputs[130]);
    assign layer0_outputs[1627] = (inputs[216]) & ~(inputs[12]);
    assign layer0_outputs[1628] = (inputs[172]) & ~(inputs[121]);
    assign layer0_outputs[1629] = 1'b1;
    assign layer0_outputs[1630] = inputs[74];
    assign layer0_outputs[1631] = ~(inputs[135]);
    assign layer0_outputs[1632] = (inputs[116]) ^ (inputs[130]);
    assign layer0_outputs[1633] = inputs[91];
    assign layer0_outputs[1634] = ~(inputs[158]) | (inputs[216]);
    assign layer0_outputs[1635] = ~((inputs[66]) ^ (inputs[106]));
    assign layer0_outputs[1636] = (inputs[83]) & (inputs[55]);
    assign layer0_outputs[1637] = ~(inputs[31]);
    assign layer0_outputs[1638] = 1'b0;
    assign layer0_outputs[1639] = 1'b0;
    assign layer0_outputs[1640] = 1'b0;
    assign layer0_outputs[1641] = (inputs[23]) & (inputs[238]);
    assign layer0_outputs[1642] = (inputs[118]) & ~(inputs[98]);
    assign layer0_outputs[1643] = ~(inputs[136]);
    assign layer0_outputs[1644] = (inputs[125]) & (inputs[20]);
    assign layer0_outputs[1645] = 1'b1;
    assign layer0_outputs[1646] = (inputs[123]) & ~(inputs[157]);
    assign layer0_outputs[1647] = inputs[159];
    assign layer0_outputs[1648] = (inputs[79]) & (inputs[51]);
    assign layer0_outputs[1649] = (inputs[14]) & (inputs[214]);
    assign layer0_outputs[1650] = ~(inputs[45]);
    assign layer0_outputs[1651] = (inputs[246]) & (inputs[26]);
    assign layer0_outputs[1652] = (inputs[186]) | (inputs[45]);
    assign layer0_outputs[1653] = inputs[183];
    assign layer0_outputs[1654] = (inputs[3]) | (inputs[166]);
    assign layer0_outputs[1655] = ~(inputs[238]) | (inputs[86]);
    assign layer0_outputs[1656] = (inputs[166]) & ~(inputs[237]);
    assign layer0_outputs[1657] = inputs[24];
    assign layer0_outputs[1658] = ~((inputs[89]) | (inputs[97]));
    assign layer0_outputs[1659] = ~((inputs[225]) | (inputs[81]));
    assign layer0_outputs[1660] = ~((inputs[68]) ^ (inputs[140]));
    assign layer0_outputs[1661] = ~(inputs[183]);
    assign layer0_outputs[1662] = ~(inputs[75]);
    assign layer0_outputs[1663] = ~(inputs[10]);
    assign layer0_outputs[1664] = inputs[10];
    assign layer0_outputs[1665] = ~(inputs[5]) | (inputs[169]);
    assign layer0_outputs[1666] = (inputs[194]) & ~(inputs[86]);
    assign layer0_outputs[1667] = ~(inputs[116]) | (inputs[171]);
    assign layer0_outputs[1668] = (inputs[192]) & ~(inputs[133]);
    assign layer0_outputs[1669] = (inputs[79]) ^ (inputs[93]);
    assign layer0_outputs[1670] = (inputs[168]) | (inputs[82]);
    assign layer0_outputs[1671] = 1'b0;
    assign layer0_outputs[1672] = inputs[164];
    assign layer0_outputs[1673] = (inputs[170]) & (inputs[89]);
    assign layer0_outputs[1674] = ~(inputs[184]) | (inputs[15]);
    assign layer0_outputs[1675] = ~(inputs[242]);
    assign layer0_outputs[1676] = ~((inputs[56]) | (inputs[172]));
    assign layer0_outputs[1677] = ~(inputs[146]);
    assign layer0_outputs[1678] = inputs[16];
    assign layer0_outputs[1679] = ~(inputs[131]);
    assign layer0_outputs[1680] = ~((inputs[190]) | (inputs[85]));
    assign layer0_outputs[1681] = ~((inputs[113]) ^ (inputs[130]));
    assign layer0_outputs[1682] = (inputs[158]) & ~(inputs[203]);
    assign layer0_outputs[1683] = ~(inputs[150]);
    assign layer0_outputs[1684] = (inputs[111]) & (inputs[12]);
    assign layer0_outputs[1685] = ~(inputs[34]);
    assign layer0_outputs[1686] = ~(inputs[3]) | (inputs[238]);
    assign layer0_outputs[1687] = ~((inputs[137]) ^ (inputs[13]));
    assign layer0_outputs[1688] = 1'b1;
    assign layer0_outputs[1689] = 1'b0;
    assign layer0_outputs[1690] = (inputs[131]) & ~(inputs[101]);
    assign layer0_outputs[1691] = 1'b1;
    assign layer0_outputs[1692] = ~((inputs[198]) ^ (inputs[35]));
    assign layer0_outputs[1693] = 1'b0;
    assign layer0_outputs[1694] = ~(inputs[233]) | (inputs[59]);
    assign layer0_outputs[1695] = (inputs[81]) & ~(inputs[19]);
    assign layer0_outputs[1696] = (inputs[108]) & ~(inputs[237]);
    assign layer0_outputs[1697] = 1'b1;
    assign layer0_outputs[1698] = inputs[58];
    assign layer0_outputs[1699] = (inputs[112]) & (inputs[141]);
    assign layer0_outputs[1700] = (inputs[184]) & ~(inputs[224]);
    assign layer0_outputs[1701] = (inputs[187]) | (inputs[189]);
    assign layer0_outputs[1702] = ~((inputs[211]) | (inputs[253]));
    assign layer0_outputs[1703] = 1'b1;
    assign layer0_outputs[1704] = (inputs[79]) & (inputs[72]);
    assign layer0_outputs[1705] = ~(inputs[125]);
    assign layer0_outputs[1706] = (inputs[112]) & (inputs[121]);
    assign layer0_outputs[1707] = (inputs[154]) & ~(inputs[212]);
    assign layer0_outputs[1708] = (inputs[190]) & ~(inputs[4]);
    assign layer0_outputs[1709] = (inputs[93]) ^ (inputs[47]);
    assign layer0_outputs[1710] = ~(inputs[144]) | (inputs[234]);
    assign layer0_outputs[1711] = ~((inputs[252]) ^ (inputs[18]));
    assign layer0_outputs[1712] = (inputs[50]) ^ (inputs[33]);
    assign layer0_outputs[1713] = ~(inputs[63]) | (inputs[185]);
    assign layer0_outputs[1714] = inputs[235];
    assign layer0_outputs[1715] = 1'b1;
    assign layer0_outputs[1716] = inputs[203];
    assign layer0_outputs[1717] = ~(inputs[250]);
    assign layer0_outputs[1718] = (inputs[35]) & ~(inputs[43]);
    assign layer0_outputs[1719] = 1'b0;
    assign layer0_outputs[1720] = ~((inputs[49]) | (inputs[105]));
    assign layer0_outputs[1721] = ~(inputs[117]) | (inputs[68]);
    assign layer0_outputs[1722] = inputs[32];
    assign layer0_outputs[1723] = 1'b0;
    assign layer0_outputs[1724] = ~((inputs[24]) & (inputs[19]));
    assign layer0_outputs[1725] = (inputs[200]) & (inputs[244]);
    assign layer0_outputs[1726] = inputs[122];
    assign layer0_outputs[1727] = (inputs[21]) | (inputs[83]);
    assign layer0_outputs[1728] = 1'b1;
    assign layer0_outputs[1729] = 1'b1;
    assign layer0_outputs[1730] = ~(inputs[150]) | (inputs[71]);
    assign layer0_outputs[1731] = ~(inputs[127]) | (inputs[125]);
    assign layer0_outputs[1732] = ~((inputs[176]) & (inputs[47]));
    assign layer0_outputs[1733] = 1'b0;
    assign layer0_outputs[1734] = (inputs[157]) | (inputs[215]);
    assign layer0_outputs[1735] = ~(inputs[155]) | (inputs[79]);
    assign layer0_outputs[1736] = ~(inputs[106]) | (inputs[179]);
    assign layer0_outputs[1737] = ~(inputs[20]);
    assign layer0_outputs[1738] = (inputs[198]) ^ (inputs[207]);
    assign layer0_outputs[1739] = ~((inputs[146]) ^ (inputs[149]));
    assign layer0_outputs[1740] = (inputs[194]) ^ (inputs[233]);
    assign layer0_outputs[1741] = ~(inputs[117]) | (inputs[172]);
    assign layer0_outputs[1742] = (inputs[237]) & ~(inputs[223]);
    assign layer0_outputs[1743] = (inputs[196]) | (inputs[211]);
    assign layer0_outputs[1744] = (inputs[133]) & ~(inputs[222]);
    assign layer0_outputs[1745] = (inputs[239]) & (inputs[27]);
    assign layer0_outputs[1746] = (inputs[82]) ^ (inputs[36]);
    assign layer0_outputs[1747] = (inputs[11]) & (inputs[138]);
    assign layer0_outputs[1748] = ~(inputs[53]) | (inputs[94]);
    assign layer0_outputs[1749] = ~(inputs[152]) | (inputs[154]);
    assign layer0_outputs[1750] = ~((inputs[78]) | (inputs[111]));
    assign layer0_outputs[1751] = (inputs[104]) & ~(inputs[204]);
    assign layer0_outputs[1752] = (inputs[56]) & ~(inputs[64]);
    assign layer0_outputs[1753] = ~(inputs[174]);
    assign layer0_outputs[1754] = 1'b1;
    assign layer0_outputs[1755] = ~((inputs[223]) | (inputs[164]));
    assign layer0_outputs[1756] = (inputs[36]) & (inputs[130]);
    assign layer0_outputs[1757] = 1'b1;
    assign layer0_outputs[1758] = ~((inputs[21]) | (inputs[229]));
    assign layer0_outputs[1759] = 1'b0;
    assign layer0_outputs[1760] = ~((inputs[108]) | (inputs[55]));
    assign layer0_outputs[1761] = ~(inputs[237]) | (inputs[69]);
    assign layer0_outputs[1762] = 1'b1;
    assign layer0_outputs[1763] = ~((inputs[130]) | (inputs[60]));
    assign layer0_outputs[1764] = inputs[124];
    assign layer0_outputs[1765] = inputs[77];
    assign layer0_outputs[1766] = ~((inputs[237]) | (inputs[148]));
    assign layer0_outputs[1767] = ~(inputs[6]);
    assign layer0_outputs[1768] = ~(inputs[196]) | (inputs[239]);
    assign layer0_outputs[1769] = ~((inputs[205]) ^ (inputs[166]));
    assign layer0_outputs[1770] = ~((inputs[242]) ^ (inputs[188]));
    assign layer0_outputs[1771] = (inputs[196]) & ~(inputs[26]);
    assign layer0_outputs[1772] = ~(inputs[182]) | (inputs[217]);
    assign layer0_outputs[1773] = ~(inputs[145]);
    assign layer0_outputs[1774] = ~(inputs[163]) | (inputs[115]);
    assign layer0_outputs[1775] = inputs[137];
    assign layer0_outputs[1776] = (inputs[4]) & (inputs[34]);
    assign layer0_outputs[1777] = inputs[31];
    assign layer0_outputs[1778] = ~(inputs[232]) | (inputs[126]);
    assign layer0_outputs[1779] = inputs[223];
    assign layer0_outputs[1780] = ~(inputs[236]) | (inputs[232]);
    assign layer0_outputs[1781] = ~(inputs[237]);
    assign layer0_outputs[1782] = ~((inputs[112]) & (inputs[27]));
    assign layer0_outputs[1783] = inputs[1];
    assign layer0_outputs[1784] = (inputs[87]) & ~(inputs[209]);
    assign layer0_outputs[1785] = 1'b1;
    assign layer0_outputs[1786] = 1'b0;
    assign layer0_outputs[1787] = (inputs[110]) | (inputs[46]);
    assign layer0_outputs[1788] = (inputs[161]) ^ (inputs[206]);
    assign layer0_outputs[1789] = ~((inputs[196]) & (inputs[139]));
    assign layer0_outputs[1790] = (inputs[2]) & ~(inputs[26]);
    assign layer0_outputs[1791] = ~(inputs[231]);
    assign layer0_outputs[1792] = (inputs[48]) ^ (inputs[129]);
    assign layer0_outputs[1793] = (inputs[163]) & ~(inputs[127]);
    assign layer0_outputs[1794] = ~(inputs[216]) | (inputs[90]);
    assign layer0_outputs[1795] = 1'b0;
    assign layer0_outputs[1796] = (inputs[119]) | (inputs[135]);
    assign layer0_outputs[1797] = (inputs[136]) ^ (inputs[224]);
    assign layer0_outputs[1798] = ~(inputs[181]) | (inputs[97]);
    assign layer0_outputs[1799] = ~(inputs[117]);
    assign layer0_outputs[1800] = ~(inputs[225]);
    assign layer0_outputs[1801] = ~((inputs[89]) & (inputs[42]));
    assign layer0_outputs[1802] = ~((inputs[25]) ^ (inputs[203]));
    assign layer0_outputs[1803] = 1'b0;
    assign layer0_outputs[1804] = inputs[149];
    assign layer0_outputs[1805] = (inputs[174]) & (inputs[169]);
    assign layer0_outputs[1806] = 1'b1;
    assign layer0_outputs[1807] = ~(inputs[254]);
    assign layer0_outputs[1808] = inputs[221];
    assign layer0_outputs[1809] = ~((inputs[86]) | (inputs[129]));
    assign layer0_outputs[1810] = (inputs[130]) & ~(inputs[179]);
    assign layer0_outputs[1811] = ~((inputs[12]) & (inputs[228]));
    assign layer0_outputs[1812] = ~(inputs[85]) | (inputs[222]);
    assign layer0_outputs[1813] = (inputs[220]) & ~(inputs[134]);
    assign layer0_outputs[1814] = ~((inputs[147]) | (inputs[43]));
    assign layer0_outputs[1815] = ~((inputs[13]) & (inputs[88]));
    assign layer0_outputs[1816] = (inputs[10]) ^ (inputs[4]);
    assign layer0_outputs[1817] = (inputs[204]) & ~(inputs[101]);
    assign layer0_outputs[1818] = (inputs[84]) & (inputs[206]);
    assign layer0_outputs[1819] = ~((inputs[228]) | (inputs[172]));
    assign layer0_outputs[1820] = 1'b1;
    assign layer0_outputs[1821] = (inputs[119]) ^ (inputs[40]);
    assign layer0_outputs[1822] = ~(inputs[8]);
    assign layer0_outputs[1823] = 1'b1;
    assign layer0_outputs[1824] = ~(inputs[243]) | (inputs[111]);
    assign layer0_outputs[1825] = (inputs[169]) | (inputs[229]);
    assign layer0_outputs[1826] = inputs[16];
    assign layer0_outputs[1827] = (inputs[1]) & ~(inputs[137]);
    assign layer0_outputs[1828] = ~(inputs[196]);
    assign layer0_outputs[1829] = ~(inputs[109]) | (inputs[23]);
    assign layer0_outputs[1830] = ~(inputs[175]) | (inputs[70]);
    assign layer0_outputs[1831] = inputs[109];
    assign layer0_outputs[1832] = 1'b0;
    assign layer0_outputs[1833] = ~((inputs[184]) & (inputs[188]));
    assign layer0_outputs[1834] = (inputs[234]) & ~(inputs[125]);
    assign layer0_outputs[1835] = 1'b1;
    assign layer0_outputs[1836] = (inputs[207]) ^ (inputs[219]);
    assign layer0_outputs[1837] = ~(inputs[113]) | (inputs[62]);
    assign layer0_outputs[1838] = ~(inputs[46]) | (inputs[230]);
    assign layer0_outputs[1839] = (inputs[189]) & (inputs[91]);
    assign layer0_outputs[1840] = inputs[69];
    assign layer0_outputs[1841] = (inputs[103]) & (inputs[42]);
    assign layer0_outputs[1842] = (inputs[46]) & ~(inputs[21]);
    assign layer0_outputs[1843] = ~(inputs[94]);
    assign layer0_outputs[1844] = ~(inputs[48]) | (inputs[88]);
    assign layer0_outputs[1845] = ~((inputs[253]) & (inputs[75]));
    assign layer0_outputs[1846] = inputs[91];
    assign layer0_outputs[1847] = ~((inputs[184]) | (inputs[142]));
    assign layer0_outputs[1848] = (inputs[200]) & ~(inputs[244]);
    assign layer0_outputs[1849] = inputs[33];
    assign layer0_outputs[1850] = ~((inputs[149]) & (inputs[118]));
    assign layer0_outputs[1851] = ~(inputs[61]);
    assign layer0_outputs[1852] = (inputs[118]) | (inputs[60]);
    assign layer0_outputs[1853] = 1'b1;
    assign layer0_outputs[1854] = (inputs[40]) & ~(inputs[104]);
    assign layer0_outputs[1855] = ~((inputs[124]) ^ (inputs[45]));
    assign layer0_outputs[1856] = ~((inputs[11]) | (inputs[126]));
    assign layer0_outputs[1857] = ~(inputs[218]) | (inputs[202]);
    assign layer0_outputs[1858] = inputs[34];
    assign layer0_outputs[1859] = inputs[5];
    assign layer0_outputs[1860] = (inputs[180]) & ~(inputs[244]);
    assign layer0_outputs[1861] = (inputs[39]) & ~(inputs[60]);
    assign layer0_outputs[1862] = inputs[56];
    assign layer0_outputs[1863] = (inputs[191]) & ~(inputs[163]);
    assign layer0_outputs[1864] = ~((inputs[183]) ^ (inputs[19]));
    assign layer0_outputs[1865] = ~(inputs[159]) | (inputs[185]);
    assign layer0_outputs[1866] = (inputs[94]) & ~(inputs[248]);
    assign layer0_outputs[1867] = 1'b1;
    assign layer0_outputs[1868] = ~(inputs[81]) | (inputs[92]);
    assign layer0_outputs[1869] = ~((inputs[152]) | (inputs[46]));
    assign layer0_outputs[1870] = ~(inputs[132]) | (inputs[61]);
    assign layer0_outputs[1871] = 1'b0;
    assign layer0_outputs[1872] = ~((inputs[87]) | (inputs[71]));
    assign layer0_outputs[1873] = inputs[181];
    assign layer0_outputs[1874] = ~((inputs[80]) | (inputs[86]));
    assign layer0_outputs[1875] = (inputs[85]) & ~(inputs[140]);
    assign layer0_outputs[1876] = (inputs[180]) & ~(inputs[67]);
    assign layer0_outputs[1877] = ~((inputs[141]) | (inputs[91]));
    assign layer0_outputs[1878] = (inputs[18]) | (inputs[44]);
    assign layer0_outputs[1879] = inputs[194];
    assign layer0_outputs[1880] = ~((inputs[111]) ^ (inputs[47]));
    assign layer0_outputs[1881] = (inputs[236]) & ~(inputs[147]);
    assign layer0_outputs[1882] = ~((inputs[0]) | (inputs[202]));
    assign layer0_outputs[1883] = ~(inputs[14]);
    assign layer0_outputs[1884] = 1'b1;
    assign layer0_outputs[1885] = (inputs[96]) & ~(inputs[218]);
    assign layer0_outputs[1886] = inputs[22];
    assign layer0_outputs[1887] = 1'b0;
    assign layer0_outputs[1888] = (inputs[224]) ^ (inputs[198]);
    assign layer0_outputs[1889] = (inputs[61]) & ~(inputs[205]);
    assign layer0_outputs[1890] = inputs[162];
    assign layer0_outputs[1891] = ~((inputs[130]) | (inputs[196]));
    assign layer0_outputs[1892] = ~((inputs[9]) | (inputs[19]));
    assign layer0_outputs[1893] = ~(inputs[68]);
    assign layer0_outputs[1894] = (inputs[203]) & (inputs[3]);
    assign layer0_outputs[1895] = inputs[154];
    assign layer0_outputs[1896] = ~((inputs[236]) | (inputs[126]));
    assign layer0_outputs[1897] = ~(inputs[192]);
    assign layer0_outputs[1898] = ~(inputs[79]) | (inputs[39]);
    assign layer0_outputs[1899] = (inputs[155]) & ~(inputs[201]);
    assign layer0_outputs[1900] = inputs[180];
    assign layer0_outputs[1901] = 1'b1;
    assign layer0_outputs[1902] = (inputs[59]) | (inputs[162]);
    assign layer0_outputs[1903] = ~(inputs[189]);
    assign layer0_outputs[1904] = (inputs[230]) ^ (inputs[67]);
    assign layer0_outputs[1905] = ~((inputs[171]) ^ (inputs[136]));
    assign layer0_outputs[1906] = inputs[4];
    assign layer0_outputs[1907] = (inputs[85]) & ~(inputs[95]);
    assign layer0_outputs[1908] = (inputs[72]) & ~(inputs[179]);
    assign layer0_outputs[1909] = inputs[26];
    assign layer0_outputs[1910] = ~((inputs[24]) | (inputs[9]));
    assign layer0_outputs[1911] = (inputs[15]) ^ (inputs[240]);
    assign layer0_outputs[1912] = (inputs[36]) | (inputs[173]);
    assign layer0_outputs[1913] = (inputs[242]) & ~(inputs[161]);
    assign layer0_outputs[1914] = ~(inputs[67]);
    assign layer0_outputs[1915] = (inputs[100]) ^ (inputs[193]);
    assign layer0_outputs[1916] = ~((inputs[31]) ^ (inputs[121]));
    assign layer0_outputs[1917] = (inputs[53]) & ~(inputs[155]);
    assign layer0_outputs[1918] = ~((inputs[135]) | (inputs[9]));
    assign layer0_outputs[1919] = ~(inputs[1]);
    assign layer0_outputs[1920] = inputs[201];
    assign layer0_outputs[1921] = ~(inputs[231]);
    assign layer0_outputs[1922] = (inputs[70]) ^ (inputs[220]);
    assign layer0_outputs[1923] = (inputs[183]) | (inputs[180]);
    assign layer0_outputs[1924] = ~(inputs[179]);
    assign layer0_outputs[1925] = 1'b0;
    assign layer0_outputs[1926] = ~(inputs[200]) | (inputs[184]);
    assign layer0_outputs[1927] = ~((inputs[132]) ^ (inputs[120]));
    assign layer0_outputs[1928] = (inputs[28]) | (inputs[249]);
    assign layer0_outputs[1929] = ~(inputs[91]);
    assign layer0_outputs[1930] = (inputs[199]) & ~(inputs[43]);
    assign layer0_outputs[1931] = ~((inputs[241]) | (inputs[120]));
    assign layer0_outputs[1932] = ~((inputs[150]) | (inputs[28]));
    assign layer0_outputs[1933] = 1'b1;
    assign layer0_outputs[1934] = (inputs[221]) | (inputs[150]);
    assign layer0_outputs[1935] = ~(inputs[147]) | (inputs[190]);
    assign layer0_outputs[1936] = (inputs[140]) ^ (inputs[20]);
    assign layer0_outputs[1937] = ~(inputs[47]);
    assign layer0_outputs[1938] = 1'b1;
    assign layer0_outputs[1939] = 1'b1;
    assign layer0_outputs[1940] = (inputs[145]) & ~(inputs[125]);
    assign layer0_outputs[1941] = ~(inputs[142]) | (inputs[139]);
    assign layer0_outputs[1942] = ~(inputs[116]) | (inputs[129]);
    assign layer0_outputs[1943] = ~((inputs[51]) & (inputs[163]));
    assign layer0_outputs[1944] = (inputs[2]) & ~(inputs[97]);
    assign layer0_outputs[1945] = inputs[170];
    assign layer0_outputs[1946] = ~((inputs[12]) & (inputs[15]));
    assign layer0_outputs[1947] = ~(inputs[225]) | (inputs[245]);
    assign layer0_outputs[1948] = 1'b0;
    assign layer0_outputs[1949] = ~((inputs[247]) | (inputs[107]));
    assign layer0_outputs[1950] = inputs[62];
    assign layer0_outputs[1951] = ~(inputs[192]);
    assign layer0_outputs[1952] = inputs[23];
    assign layer0_outputs[1953] = (inputs[216]) ^ (inputs[252]);
    assign layer0_outputs[1954] = 1'b1;
    assign layer0_outputs[1955] = inputs[92];
    assign layer0_outputs[1956] = 1'b0;
    assign layer0_outputs[1957] = 1'b1;
    assign layer0_outputs[1958] = ~((inputs[10]) & (inputs[176]));
    assign layer0_outputs[1959] = ~((inputs[8]) ^ (inputs[160]));
    assign layer0_outputs[1960] = ~(inputs[234]);
    assign layer0_outputs[1961] = inputs[41];
    assign layer0_outputs[1962] = 1'b0;
    assign layer0_outputs[1963] = ~(inputs[198]);
    assign layer0_outputs[1964] = (inputs[15]) ^ (inputs[61]);
    assign layer0_outputs[1965] = ~((inputs[205]) ^ (inputs[79]));
    assign layer0_outputs[1966] = 1'b1;
    assign layer0_outputs[1967] = (inputs[145]) | (inputs[38]);
    assign layer0_outputs[1968] = ~(inputs[211]);
    assign layer0_outputs[1969] = ~(inputs[185]);
    assign layer0_outputs[1970] = (inputs[112]) & ~(inputs[33]);
    assign layer0_outputs[1971] = ~((inputs[36]) ^ (inputs[92]));
    assign layer0_outputs[1972] = ~(inputs[184]);
    assign layer0_outputs[1973] = (inputs[219]) | (inputs[133]);
    assign layer0_outputs[1974] = (inputs[66]) & ~(inputs[96]);
    assign layer0_outputs[1975] = (inputs[228]) ^ (inputs[207]);
    assign layer0_outputs[1976] = ~((inputs[97]) & (inputs[148]));
    assign layer0_outputs[1977] = ~(inputs[197]) | (inputs[61]);
    assign layer0_outputs[1978] = (inputs[90]) ^ (inputs[166]);
    assign layer0_outputs[1979] = ~((inputs[83]) | (inputs[165]));
    assign layer0_outputs[1980] = ~((inputs[200]) & (inputs[75]));
    assign layer0_outputs[1981] = (inputs[165]) | (inputs[157]);
    assign layer0_outputs[1982] = ~(inputs[225]);
    assign layer0_outputs[1983] = ~(inputs[51]) | (inputs[245]);
    assign layer0_outputs[1984] = ~(inputs[133]);
    assign layer0_outputs[1985] = 1'b1;
    assign layer0_outputs[1986] = inputs[8];
    assign layer0_outputs[1987] = ~(inputs[214]);
    assign layer0_outputs[1988] = (inputs[140]) & ~(inputs[204]);
    assign layer0_outputs[1989] = ~((inputs[239]) & (inputs[99]));
    assign layer0_outputs[1990] = (inputs[128]) & ~(inputs[0]);
    assign layer0_outputs[1991] = ~(inputs[6]);
    assign layer0_outputs[1992] = (inputs[50]) & ~(inputs[220]);
    assign layer0_outputs[1993] = ~(inputs[120]);
    assign layer0_outputs[1994] = (inputs[129]) ^ (inputs[124]);
    assign layer0_outputs[1995] = (inputs[135]) & ~(inputs[176]);
    assign layer0_outputs[1996] = 1'b0;
    assign layer0_outputs[1997] = (inputs[140]) & ~(inputs[222]);
    assign layer0_outputs[1998] = 1'b1;
    assign layer0_outputs[1999] = 1'b1;
    assign layer0_outputs[2000] = 1'b1;
    assign layer0_outputs[2001] = ~((inputs[28]) ^ (inputs[125]));
    assign layer0_outputs[2002] = ~(inputs[82]);
    assign layer0_outputs[2003] = ~(inputs[164]) | (inputs[5]);
    assign layer0_outputs[2004] = ~(inputs[10]);
    assign layer0_outputs[2005] = (inputs[154]) | (inputs[234]);
    assign layer0_outputs[2006] = inputs[71];
    assign layer0_outputs[2007] = ~(inputs[178]);
    assign layer0_outputs[2008] = (inputs[12]) ^ (inputs[145]);
    assign layer0_outputs[2009] = 1'b0;
    assign layer0_outputs[2010] = ~(inputs[86]) | (inputs[237]);
    assign layer0_outputs[2011] = ~(inputs[186]) | (inputs[46]);
    assign layer0_outputs[2012] = ~(inputs[243]) | (inputs[45]);
    assign layer0_outputs[2013] = 1'b1;
    assign layer0_outputs[2014] = ~(inputs[206]) | (inputs[245]);
    assign layer0_outputs[2015] = ~((inputs[253]) ^ (inputs[64]));
    assign layer0_outputs[2016] = (inputs[186]) | (inputs[22]);
    assign layer0_outputs[2017] = (inputs[194]) & ~(inputs[90]);
    assign layer0_outputs[2018] = (inputs[163]) ^ (inputs[200]);
    assign layer0_outputs[2019] = inputs[218];
    assign layer0_outputs[2020] = ~(inputs[161]);
    assign layer0_outputs[2021] = ~((inputs[249]) | (inputs[89]));
    assign layer0_outputs[2022] = ~((inputs[9]) ^ (inputs[60]));
    assign layer0_outputs[2023] = (inputs[221]) ^ (inputs[63]);
    assign layer0_outputs[2024] = inputs[27];
    assign layer0_outputs[2025] = ~((inputs[148]) | (inputs[24]));
    assign layer0_outputs[2026] = (inputs[185]) | (inputs[153]);
    assign layer0_outputs[2027] = ~((inputs[215]) | (inputs[104]));
    assign layer0_outputs[2028] = ~(inputs[132]) | (inputs[206]);
    assign layer0_outputs[2029] = ~(inputs[131]);
    assign layer0_outputs[2030] = ~(inputs[34]);
    assign layer0_outputs[2031] = (inputs[208]) & ~(inputs[172]);
    assign layer0_outputs[2032] = 1'b0;
    assign layer0_outputs[2033] = ~((inputs[179]) | (inputs[119]));
    assign layer0_outputs[2034] = ~(inputs[86]);
    assign layer0_outputs[2035] = (inputs[88]) & ~(inputs[156]);
    assign layer0_outputs[2036] = ~((inputs[124]) | (inputs[36]));
    assign layer0_outputs[2037] = ~((inputs[118]) ^ (inputs[49]));
    assign layer0_outputs[2038] = (inputs[23]) | (inputs[182]);
    assign layer0_outputs[2039] = ~((inputs[143]) ^ (inputs[248]));
    assign layer0_outputs[2040] = (inputs[39]) & ~(inputs[213]);
    assign layer0_outputs[2041] = ~((inputs[38]) ^ (inputs[17]));
    assign layer0_outputs[2042] = ~((inputs[53]) | (inputs[154]));
    assign layer0_outputs[2043] = 1'b0;
    assign layer0_outputs[2044] = (inputs[197]) & ~(inputs[159]);
    assign layer0_outputs[2045] = (inputs[46]) & ~(inputs[66]);
    assign layer0_outputs[2046] = 1'b0;
    assign layer0_outputs[2047] = ~((inputs[158]) | (inputs[186]));
    assign layer0_outputs[2048] = ~(inputs[42]);
    assign layer0_outputs[2049] = ~((inputs[185]) & (inputs[182]));
    assign layer0_outputs[2050] = (inputs[103]) & ~(inputs[234]);
    assign layer0_outputs[2051] = ~(inputs[48]);
    assign layer0_outputs[2052] = ~((inputs[49]) ^ (inputs[231]));
    assign layer0_outputs[2053] = (inputs[179]) | (inputs[252]);
    assign layer0_outputs[2054] = 1'b1;
    assign layer0_outputs[2055] = ~(inputs[110]) | (inputs[18]);
    assign layer0_outputs[2056] = ~(inputs[152]);
    assign layer0_outputs[2057] = inputs[181];
    assign layer0_outputs[2058] = ~(inputs[78]);
    assign layer0_outputs[2059] = ~(inputs[91]) | (inputs[4]);
    assign layer0_outputs[2060] = (inputs[190]) & ~(inputs[252]);
    assign layer0_outputs[2061] = ~((inputs[39]) | (inputs[12]));
    assign layer0_outputs[2062] = 1'b1;
    assign layer0_outputs[2063] = ~(inputs[92]);
    assign layer0_outputs[2064] = (inputs[252]) & (inputs[64]);
    assign layer0_outputs[2065] = (inputs[188]) | (inputs[57]);
    assign layer0_outputs[2066] = (inputs[186]) | (inputs[4]);
    assign layer0_outputs[2067] = ~(inputs[250]);
    assign layer0_outputs[2068] = (inputs[147]) | (inputs[231]);
    assign layer0_outputs[2069] = 1'b1;
    assign layer0_outputs[2070] = (inputs[180]) | (inputs[158]);
    assign layer0_outputs[2071] = ~(inputs[165]) | (inputs[202]);
    assign layer0_outputs[2072] = ~((inputs[4]) | (inputs[249]));
    assign layer0_outputs[2073] = ~((inputs[240]) ^ (inputs[159]));
    assign layer0_outputs[2074] = (inputs[174]) | (inputs[21]);
    assign layer0_outputs[2075] = ~((inputs[94]) ^ (inputs[3]));
    assign layer0_outputs[2076] = ~((inputs[75]) & (inputs[23]));
    assign layer0_outputs[2077] = ~(inputs[206]);
    assign layer0_outputs[2078] = 1'b1;
    assign layer0_outputs[2079] = ~((inputs[131]) | (inputs[87]));
    assign layer0_outputs[2080] = 1'b1;
    assign layer0_outputs[2081] = 1'b0;
    assign layer0_outputs[2082] = ~(inputs[36]) | (inputs[1]);
    assign layer0_outputs[2083] = ~((inputs[117]) | (inputs[39]));
    assign layer0_outputs[2084] = ~((inputs[74]) & (inputs[241]));
    assign layer0_outputs[2085] = ~(inputs[87]) | (inputs[161]);
    assign layer0_outputs[2086] = 1'b0;
    assign layer0_outputs[2087] = ~(inputs[238]);
    assign layer0_outputs[2088] = ~((inputs[205]) | (inputs[244]));
    assign layer0_outputs[2089] = 1'b0;
    assign layer0_outputs[2090] = (inputs[6]) & ~(inputs[241]);
    assign layer0_outputs[2091] = ~((inputs[102]) | (inputs[44]));
    assign layer0_outputs[2092] = (inputs[151]) | (inputs[97]);
    assign layer0_outputs[2093] = (inputs[114]) ^ (inputs[198]);
    assign layer0_outputs[2094] = ~(inputs[228]);
    assign layer0_outputs[2095] = (inputs[88]) ^ (inputs[20]);
    assign layer0_outputs[2096] = 1'b0;
    assign layer0_outputs[2097] = 1'b1;
    assign layer0_outputs[2098] = (inputs[176]) & ~(inputs[158]);
    assign layer0_outputs[2099] = inputs[124];
    assign layer0_outputs[2100] = ~((inputs[106]) | (inputs[50]));
    assign layer0_outputs[2101] = ~((inputs[178]) & (inputs[219]));
    assign layer0_outputs[2102] = ~(inputs[208]) | (inputs[182]);
    assign layer0_outputs[2103] = (inputs[110]) ^ (inputs[54]);
    assign layer0_outputs[2104] = (inputs[84]) | (inputs[76]);
    assign layer0_outputs[2105] = ~(inputs[13]);
    assign layer0_outputs[2106] = ~(inputs[52]);
    assign layer0_outputs[2107] = (inputs[73]) & ~(inputs[130]);
    assign layer0_outputs[2108] = (inputs[115]) | (inputs[183]);
    assign layer0_outputs[2109] = ~((inputs[90]) | (inputs[217]));
    assign layer0_outputs[2110] = ~(inputs[91]) | (inputs[29]);
    assign layer0_outputs[2111] = (inputs[249]) ^ (inputs[27]);
    assign layer0_outputs[2112] = ~(inputs[66]);
    assign layer0_outputs[2113] = 1'b0;
    assign layer0_outputs[2114] = ~((inputs[147]) | (inputs[123]));
    assign layer0_outputs[2115] = (inputs[164]) ^ (inputs[238]);
    assign layer0_outputs[2116] = (inputs[66]) ^ (inputs[7]);
    assign layer0_outputs[2117] = ~(inputs[98]);
    assign layer0_outputs[2118] = (inputs[145]) | (inputs[128]);
    assign layer0_outputs[2119] = ~(inputs[230]);
    assign layer0_outputs[2120] = ~(inputs[34]);
    assign layer0_outputs[2121] = ~(inputs[164]);
    assign layer0_outputs[2122] = (inputs[22]) ^ (inputs[35]);
    assign layer0_outputs[2123] = ~(inputs[15]);
    assign layer0_outputs[2124] = ~((inputs[233]) | (inputs[204]));
    assign layer0_outputs[2125] = ~((inputs[31]) ^ (inputs[185]));
    assign layer0_outputs[2126] = 1'b1;
    assign layer0_outputs[2127] = (inputs[6]) & ~(inputs[65]);
    assign layer0_outputs[2128] = ~(inputs[232]) | (inputs[101]);
    assign layer0_outputs[2129] = ~((inputs[192]) | (inputs[17]));
    assign layer0_outputs[2130] = ~(inputs[12]) | (inputs[121]);
    assign layer0_outputs[2131] = ~((inputs[66]) | (inputs[22]));
    assign layer0_outputs[2132] = ~((inputs[166]) | (inputs[205]));
    assign layer0_outputs[2133] = 1'b1;
    assign layer0_outputs[2134] = (inputs[232]) & (inputs[16]);
    assign layer0_outputs[2135] = ~(inputs[14]);
    assign layer0_outputs[2136] = inputs[211];
    assign layer0_outputs[2137] = ~((inputs[110]) | (inputs[12]));
    assign layer0_outputs[2138] = ~((inputs[203]) | (inputs[234]));
    assign layer0_outputs[2139] = ~(inputs[59]) | (inputs[38]);
    assign layer0_outputs[2140] = (inputs[75]) & ~(inputs[219]);
    assign layer0_outputs[2141] = ~(inputs[54]);
    assign layer0_outputs[2142] = ~(inputs[128]);
    assign layer0_outputs[2143] = ~(inputs[8]) | (inputs[88]);
    assign layer0_outputs[2144] = 1'b0;
    assign layer0_outputs[2145] = ~(inputs[65]) | (inputs[238]);
    assign layer0_outputs[2146] = inputs[57];
    assign layer0_outputs[2147] = 1'b0;
    assign layer0_outputs[2148] = ~((inputs[180]) & (inputs[39]));
    assign layer0_outputs[2149] = ~(inputs[87]);
    assign layer0_outputs[2150] = (inputs[243]) & ~(inputs[232]);
    assign layer0_outputs[2151] = inputs[13];
    assign layer0_outputs[2152] = ~((inputs[220]) | (inputs[37]));
    assign layer0_outputs[2153] = inputs[106];
    assign layer0_outputs[2154] = (inputs[157]) & (inputs[123]);
    assign layer0_outputs[2155] = (inputs[159]) & ~(inputs[52]);
    assign layer0_outputs[2156] = (inputs[124]) & ~(inputs[20]);
    assign layer0_outputs[2157] = (inputs[50]) & (inputs[49]);
    assign layer0_outputs[2158] = ~(inputs[29]);
    assign layer0_outputs[2159] = inputs[222];
    assign layer0_outputs[2160] = ~((inputs[23]) | (inputs[104]));
    assign layer0_outputs[2161] = ~((inputs[140]) | (inputs[160]));
    assign layer0_outputs[2162] = inputs[61];
    assign layer0_outputs[2163] = (inputs[221]) & (inputs[69]);
    assign layer0_outputs[2164] = 1'b0;
    assign layer0_outputs[2165] = ~((inputs[89]) | (inputs[73]));
    assign layer0_outputs[2166] = ~(inputs[137]);
    assign layer0_outputs[2167] = ~(inputs[62]) | (inputs[46]);
    assign layer0_outputs[2168] = inputs[220];
    assign layer0_outputs[2169] = 1'b0;
    assign layer0_outputs[2170] = (inputs[63]) & ~(inputs[92]);
    assign layer0_outputs[2171] = ~(inputs[38]) | (inputs[114]);
    assign layer0_outputs[2172] = 1'b0;
    assign layer0_outputs[2173] = (inputs[37]) ^ (inputs[59]);
    assign layer0_outputs[2174] = inputs[76];
    assign layer0_outputs[2175] = ~((inputs[233]) ^ (inputs[156]));
    assign layer0_outputs[2176] = ~(inputs[45]) | (inputs[221]);
    assign layer0_outputs[2177] = inputs[150];
    assign layer0_outputs[2178] = ~(inputs[56]) | (inputs[49]);
    assign layer0_outputs[2179] = ~(inputs[37]);
    assign layer0_outputs[2180] = ~((inputs[224]) ^ (inputs[206]));
    assign layer0_outputs[2181] = inputs[143];
    assign layer0_outputs[2182] = ~((inputs[160]) & (inputs[110]));
    assign layer0_outputs[2183] = 1'b1;
    assign layer0_outputs[2184] = ~(inputs[7]) | (inputs[182]);
    assign layer0_outputs[2185] = 1'b1;
    assign layer0_outputs[2186] = 1'b1;
    assign layer0_outputs[2187] = 1'b0;
    assign layer0_outputs[2188] = inputs[100];
    assign layer0_outputs[2189] = ~(inputs[191]);
    assign layer0_outputs[2190] = (inputs[156]) & ~(inputs[200]);
    assign layer0_outputs[2191] = ~(inputs[44]) | (inputs[200]);
    assign layer0_outputs[2192] = inputs[127];
    assign layer0_outputs[2193] = ~(inputs[225]) | (inputs[43]);
    assign layer0_outputs[2194] = ~((inputs[99]) | (inputs[190]));
    assign layer0_outputs[2195] = ~(inputs[63]);
    assign layer0_outputs[2196] = ~(inputs[29]);
    assign layer0_outputs[2197] = 1'b0;
    assign layer0_outputs[2198] = ~(inputs[243]) | (inputs[64]);
    assign layer0_outputs[2199] = inputs[122];
    assign layer0_outputs[2200] = (inputs[42]) & ~(inputs[147]);
    assign layer0_outputs[2201] = ~((inputs[210]) ^ (inputs[241]));
    assign layer0_outputs[2202] = ~((inputs[64]) ^ (inputs[213]));
    assign layer0_outputs[2203] = 1'b0;
    assign layer0_outputs[2204] = (inputs[209]) & (inputs[52]);
    assign layer0_outputs[2205] = ~((inputs[180]) & (inputs[96]));
    assign layer0_outputs[2206] = (inputs[246]) & (inputs[65]);
    assign layer0_outputs[2207] = inputs[246];
    assign layer0_outputs[2208] = ~(inputs[38]);
    assign layer0_outputs[2209] = (inputs[122]) & ~(inputs[64]);
    assign layer0_outputs[2210] = inputs[55];
    assign layer0_outputs[2211] = ~(inputs[181]) | (inputs[229]);
    assign layer0_outputs[2212] = (inputs[227]) & (inputs[179]);
    assign layer0_outputs[2213] = 1'b1;
    assign layer0_outputs[2214] = inputs[127];
    assign layer0_outputs[2215] = (inputs[40]) & ~(inputs[190]);
    assign layer0_outputs[2216] = ~(inputs[184]);
    assign layer0_outputs[2217] = 1'b1;
    assign layer0_outputs[2218] = (inputs[68]) | (inputs[179]);
    assign layer0_outputs[2219] = ~(inputs[189]) | (inputs[10]);
    assign layer0_outputs[2220] = (inputs[168]) & ~(inputs[41]);
    assign layer0_outputs[2221] = ~(inputs[237]) | (inputs[202]);
    assign layer0_outputs[2222] = ~(inputs[214]);
    assign layer0_outputs[2223] = ~(inputs[230]) | (inputs[239]);
    assign layer0_outputs[2224] = 1'b1;
    assign layer0_outputs[2225] = ~((inputs[75]) & (inputs[42]));
    assign layer0_outputs[2226] = ~(inputs[254]);
    assign layer0_outputs[2227] = (inputs[219]) & ~(inputs[108]);
    assign layer0_outputs[2228] = ~(inputs[81]);
    assign layer0_outputs[2229] = (inputs[97]) ^ (inputs[215]);
    assign layer0_outputs[2230] = ~((inputs[250]) ^ (inputs[205]));
    assign layer0_outputs[2231] = (inputs[2]) | (inputs[227]);
    assign layer0_outputs[2232] = (inputs[14]) & (inputs[178]);
    assign layer0_outputs[2233] = 1'b0;
    assign layer0_outputs[2234] = (inputs[78]) | (inputs[117]);
    assign layer0_outputs[2235] = ~((inputs[58]) | (inputs[56]));
    assign layer0_outputs[2236] = ~(inputs[157]) | (inputs[113]);
    assign layer0_outputs[2237] = 1'b0;
    assign layer0_outputs[2238] = (inputs[19]) & (inputs[43]);
    assign layer0_outputs[2239] = ~(inputs[62]);
    assign layer0_outputs[2240] = (inputs[229]) & (inputs[94]);
    assign layer0_outputs[2241] = (inputs[145]) & ~(inputs[208]);
    assign layer0_outputs[2242] = (inputs[213]) | (inputs[193]);
    assign layer0_outputs[2243] = (inputs[151]) & ~(inputs[88]);
    assign layer0_outputs[2244] = (inputs[92]) & ~(inputs[101]);
    assign layer0_outputs[2245] = 1'b0;
    assign layer0_outputs[2246] = ~((inputs[226]) & (inputs[237]));
    assign layer0_outputs[2247] = 1'b0;
    assign layer0_outputs[2248] = (inputs[250]) | (inputs[105]);
    assign layer0_outputs[2249] = ~(inputs[92]);
    assign layer0_outputs[2250] = ~(inputs[80]);
    assign layer0_outputs[2251] = ~(inputs[194]) | (inputs[119]);
    assign layer0_outputs[2252] = 1'b0;
    assign layer0_outputs[2253] = (inputs[66]) & ~(inputs[95]);
    assign layer0_outputs[2254] = (inputs[233]) | (inputs[120]);
    assign layer0_outputs[2255] = ~((inputs[5]) ^ (inputs[65]));
    assign layer0_outputs[2256] = 1'b0;
    assign layer0_outputs[2257] = ~(inputs[209]) | (inputs[56]);
    assign layer0_outputs[2258] = 1'b1;
    assign layer0_outputs[2259] = 1'b0;
    assign layer0_outputs[2260] = 1'b0;
    assign layer0_outputs[2261] = (inputs[75]) & ~(inputs[67]);
    assign layer0_outputs[2262] = inputs[173];
    assign layer0_outputs[2263] = 1'b1;
    assign layer0_outputs[2264] = ~(inputs[135]);
    assign layer0_outputs[2265] = (inputs[4]) | (inputs[83]);
    assign layer0_outputs[2266] = inputs[199];
    assign layer0_outputs[2267] = 1'b1;
    assign layer0_outputs[2268] = inputs[65];
    assign layer0_outputs[2269] = (inputs[135]) & ~(inputs[28]);
    assign layer0_outputs[2270] = ~(inputs[135]);
    assign layer0_outputs[2271] = (inputs[41]) | (inputs[37]);
    assign layer0_outputs[2272] = (inputs[199]) & (inputs[175]);
    assign layer0_outputs[2273] = (inputs[127]) & ~(inputs[4]);
    assign layer0_outputs[2274] = ~(inputs[141]) | (inputs[66]);
    assign layer0_outputs[2275] = ~(inputs[204]);
    assign layer0_outputs[2276] = (inputs[191]) & (inputs[154]);
    assign layer0_outputs[2277] = (inputs[145]) ^ (inputs[204]);
    assign layer0_outputs[2278] = inputs[69];
    assign layer0_outputs[2279] = inputs[130];
    assign layer0_outputs[2280] = (inputs[14]) & ~(inputs[19]);
    assign layer0_outputs[2281] = ~((inputs[202]) | (inputs[229]));
    assign layer0_outputs[2282] = (inputs[183]) ^ (inputs[28]);
    assign layer0_outputs[2283] = ~(inputs[98]);
    assign layer0_outputs[2284] = (inputs[27]) ^ (inputs[120]);
    assign layer0_outputs[2285] = ~((inputs[128]) | (inputs[227]));
    assign layer0_outputs[2286] = (inputs[17]) | (inputs[109]);
    assign layer0_outputs[2287] = 1'b1;
    assign layer0_outputs[2288] = (inputs[167]) & ~(inputs[195]);
    assign layer0_outputs[2289] = ~((inputs[122]) & (inputs[150]));
    assign layer0_outputs[2290] = 1'b1;
    assign layer0_outputs[2291] = ~(inputs[42]);
    assign layer0_outputs[2292] = (inputs[253]) & (inputs[87]);
    assign layer0_outputs[2293] = ~(inputs[101]);
    assign layer0_outputs[2294] = 1'b1;
    assign layer0_outputs[2295] = (inputs[160]) ^ (inputs[31]);
    assign layer0_outputs[2296] = ~(inputs[195]) | (inputs[33]);
    assign layer0_outputs[2297] = inputs[136];
    assign layer0_outputs[2298] = ~((inputs[178]) ^ (inputs[119]));
    assign layer0_outputs[2299] = ~((inputs[166]) | (inputs[125]));
    assign layer0_outputs[2300] = ~((inputs[213]) | (inputs[90]));
    assign layer0_outputs[2301] = ~(inputs[173]) | (inputs[241]);
    assign layer0_outputs[2302] = ~(inputs[204]) | (inputs[252]);
    assign layer0_outputs[2303] = ~(inputs[132]) | (inputs[157]);
    assign layer0_outputs[2304] = inputs[97];
    assign layer0_outputs[2305] = ~((inputs[185]) & (inputs[28]));
    assign layer0_outputs[2306] = ~(inputs[16]) | (inputs[132]);
    assign layer0_outputs[2307] = (inputs[218]) & (inputs[180]);
    assign layer0_outputs[2308] = ~((inputs[177]) | (inputs[80]));
    assign layer0_outputs[2309] = ~(inputs[163]) | (inputs[242]);
    assign layer0_outputs[2310] = inputs[75];
    assign layer0_outputs[2311] = ~(inputs[96]);
    assign layer0_outputs[2312] = (inputs[69]) | (inputs[67]);
    assign layer0_outputs[2313] = ~(inputs[180]) | (inputs[235]);
    assign layer0_outputs[2314] = ~((inputs[123]) | (inputs[17]));
    assign layer0_outputs[2315] = 1'b1;
    assign layer0_outputs[2316] = 1'b1;
    assign layer0_outputs[2317] = 1'b1;
    assign layer0_outputs[2318] = ~(inputs[198]) | (inputs[198]);
    assign layer0_outputs[2319] = ~((inputs[14]) | (inputs[101]));
    assign layer0_outputs[2320] = ~(inputs[203]) | (inputs[15]);
    assign layer0_outputs[2321] = (inputs[94]) & ~(inputs[0]);
    assign layer0_outputs[2322] = (inputs[81]) ^ (inputs[23]);
    assign layer0_outputs[2323] = ~((inputs[75]) & (inputs[110]));
    assign layer0_outputs[2324] = ~(inputs[9]) | (inputs[173]);
    assign layer0_outputs[2325] = ~((inputs[99]) | (inputs[142]));
    assign layer0_outputs[2326] = (inputs[183]) & ~(inputs[96]);
    assign layer0_outputs[2327] = ~((inputs[238]) & (inputs[119]));
    assign layer0_outputs[2328] = inputs[249];
    assign layer0_outputs[2329] = ~(inputs[187]) | (inputs[155]);
    assign layer0_outputs[2330] = (inputs[68]) | (inputs[22]);
    assign layer0_outputs[2331] = 1'b1;
    assign layer0_outputs[2332] = (inputs[64]) & (inputs[79]);
    assign layer0_outputs[2333] = ~((inputs[155]) | (inputs[32]));
    assign layer0_outputs[2334] = 1'b0;
    assign layer0_outputs[2335] = ~((inputs[54]) | (inputs[54]));
    assign layer0_outputs[2336] = ~(inputs[135]);
    assign layer0_outputs[2337] = 1'b1;
    assign layer0_outputs[2338] = ~(inputs[19]);
    assign layer0_outputs[2339] = ~((inputs[181]) | (inputs[25]));
    assign layer0_outputs[2340] = ~(inputs[2]);
    assign layer0_outputs[2341] = (inputs[139]) & ~(inputs[177]);
    assign layer0_outputs[2342] = ~((inputs[4]) | (inputs[6]));
    assign layer0_outputs[2343] = (inputs[84]) & ~(inputs[160]);
    assign layer0_outputs[2344] = ~(inputs[179]);
    assign layer0_outputs[2345] = (inputs[208]) & (inputs[180]);
    assign layer0_outputs[2346] = ~(inputs[226]);
    assign layer0_outputs[2347] = (inputs[249]) ^ (inputs[13]);
    assign layer0_outputs[2348] = ~(inputs[39]) | (inputs[247]);
    assign layer0_outputs[2349] = ~((inputs[218]) | (inputs[82]));
    assign layer0_outputs[2350] = (inputs[21]) ^ (inputs[95]);
    assign layer0_outputs[2351] = (inputs[25]) | (inputs[26]);
    assign layer0_outputs[2352] = ~(inputs[149]) | (inputs[224]);
    assign layer0_outputs[2353] = (inputs[154]) & (inputs[166]);
    assign layer0_outputs[2354] = (inputs[64]) & ~(inputs[94]);
    assign layer0_outputs[2355] = (inputs[82]) ^ (inputs[158]);
    assign layer0_outputs[2356] = 1'b1;
    assign layer0_outputs[2357] = ~(inputs[190]);
    assign layer0_outputs[2358] = (inputs[244]) & (inputs[216]);
    assign layer0_outputs[2359] = inputs[13];
    assign layer0_outputs[2360] = ~(inputs[148]);
    assign layer0_outputs[2361] = ~(inputs[234]) | (inputs[150]);
    assign layer0_outputs[2362] = ~((inputs[64]) ^ (inputs[7]));
    assign layer0_outputs[2363] = (inputs[116]) & ~(inputs[142]);
    assign layer0_outputs[2364] = ~((inputs[31]) & (inputs[161]));
    assign layer0_outputs[2365] = ~(inputs[135]);
    assign layer0_outputs[2366] = (inputs[165]) | (inputs[173]);
    assign layer0_outputs[2367] = ~(inputs[145]) | (inputs[125]);
    assign layer0_outputs[2368] = inputs[50];
    assign layer0_outputs[2369] = ~((inputs[74]) & (inputs[117]));
    assign layer0_outputs[2370] = ~((inputs[201]) ^ (inputs[25]));
    assign layer0_outputs[2371] = (inputs[237]) & (inputs[4]);
    assign layer0_outputs[2372] = (inputs[189]) | (inputs[136]);
    assign layer0_outputs[2373] = ~(inputs[219]) | (inputs[72]);
    assign layer0_outputs[2374] = (inputs[110]) & ~(inputs[189]);
    assign layer0_outputs[2375] = (inputs[138]) | (inputs[137]);
    assign layer0_outputs[2376] = ~(inputs[4]) | (inputs[54]);
    assign layer0_outputs[2377] = ~(inputs[141]) | (inputs[6]);
    assign layer0_outputs[2378] = ~(inputs[116]);
    assign layer0_outputs[2379] = (inputs[68]) | (inputs[81]);
    assign layer0_outputs[2380] = 1'b1;
    assign layer0_outputs[2381] = 1'b1;
    assign layer0_outputs[2382] = 1'b1;
    assign layer0_outputs[2383] = ~((inputs[34]) ^ (inputs[226]));
    assign layer0_outputs[2384] = inputs[102];
    assign layer0_outputs[2385] = ~(inputs[225]) | (inputs[170]);
    assign layer0_outputs[2386] = ~((inputs[41]) & (inputs[122]));
    assign layer0_outputs[2387] = ~(inputs[97]) | (inputs[160]);
    assign layer0_outputs[2388] = 1'b1;
    assign layer0_outputs[2389] = (inputs[131]) & (inputs[38]);
    assign layer0_outputs[2390] = (inputs[181]) | (inputs[101]);
    assign layer0_outputs[2391] = (inputs[5]) & ~(inputs[32]);
    assign layer0_outputs[2392] = ~((inputs[43]) | (inputs[160]));
    assign layer0_outputs[2393] = ~(inputs[195]) | (inputs[31]);
    assign layer0_outputs[2394] = ~(inputs[217]);
    assign layer0_outputs[2395] = 1'b1;
    assign layer0_outputs[2396] = (inputs[74]) & ~(inputs[170]);
    assign layer0_outputs[2397] = 1'b1;
    assign layer0_outputs[2398] = ~((inputs[191]) | (inputs[165]));
    assign layer0_outputs[2399] = ~((inputs[162]) & (inputs[50]));
    assign layer0_outputs[2400] = ~(inputs[23]) | (inputs[164]);
    assign layer0_outputs[2401] = ~((inputs[209]) ^ (inputs[58]));
    assign layer0_outputs[2402] = (inputs[60]) & ~(inputs[200]);
    assign layer0_outputs[2403] = inputs[4];
    assign layer0_outputs[2404] = (inputs[247]) & ~(inputs[182]);
    assign layer0_outputs[2405] = 1'b1;
    assign layer0_outputs[2406] = ~(inputs[21]);
    assign layer0_outputs[2407] = ~(inputs[51]) | (inputs[7]);
    assign layer0_outputs[2408] = ~((inputs[186]) | (inputs[58]));
    assign layer0_outputs[2409] = ~(inputs[4]) | (inputs[107]);
    assign layer0_outputs[2410] = ~((inputs[91]) | (inputs[162]));
    assign layer0_outputs[2411] = (inputs[156]) & ~(inputs[180]);
    assign layer0_outputs[2412] = ~(inputs[248]) | (inputs[221]);
    assign layer0_outputs[2413] = 1'b1;
    assign layer0_outputs[2414] = ~(inputs[99]) | (inputs[192]);
    assign layer0_outputs[2415] = 1'b1;
    assign layer0_outputs[2416] = (inputs[209]) | (inputs[145]);
    assign layer0_outputs[2417] = (inputs[243]) & ~(inputs[49]);
    assign layer0_outputs[2418] = (inputs[227]) & (inputs[66]);
    assign layer0_outputs[2419] = (inputs[205]) & (inputs[154]);
    assign layer0_outputs[2420] = inputs[46];
    assign layer0_outputs[2421] = ~((inputs[34]) & (inputs[219]));
    assign layer0_outputs[2422] = ~((inputs[186]) ^ (inputs[33]));
    assign layer0_outputs[2423] = 1'b0;
    assign layer0_outputs[2424] = inputs[19];
    assign layer0_outputs[2425] = (inputs[238]) | (inputs[236]);
    assign layer0_outputs[2426] = ~((inputs[220]) | (inputs[195]));
    assign layer0_outputs[2427] = ~((inputs[21]) & (inputs[83]));
    assign layer0_outputs[2428] = ~((inputs[37]) ^ (inputs[74]));
    assign layer0_outputs[2429] = ~(inputs[107]) | (inputs[173]);
    assign layer0_outputs[2430] = 1'b1;
    assign layer0_outputs[2431] = 1'b0;
    assign layer0_outputs[2432] = (inputs[52]) & ~(inputs[71]);
    assign layer0_outputs[2433] = 1'b1;
    assign layer0_outputs[2434] = ~((inputs[210]) | (inputs[48]));
    assign layer0_outputs[2435] = (inputs[178]) & (inputs[80]);
    assign layer0_outputs[2436] = inputs[71];
    assign layer0_outputs[2437] = inputs[188];
    assign layer0_outputs[2438] = ~(inputs[242]);
    assign layer0_outputs[2439] = ~(inputs[138]) | (inputs[204]);
    assign layer0_outputs[2440] = (inputs[159]) & ~(inputs[176]);
    assign layer0_outputs[2441] = (inputs[25]) & (inputs[109]);
    assign layer0_outputs[2442] = ~((inputs[68]) ^ (inputs[255]));
    assign layer0_outputs[2443] = (inputs[125]) | (inputs[95]);
    assign layer0_outputs[2444] = ~(inputs[177]);
    assign layer0_outputs[2445] = (inputs[136]) & ~(inputs[55]);
    assign layer0_outputs[2446] = (inputs[142]) & ~(inputs[11]);
    assign layer0_outputs[2447] = 1'b1;
    assign layer0_outputs[2448] = ~(inputs[104]);
    assign layer0_outputs[2449] = (inputs[98]) & (inputs[116]);
    assign layer0_outputs[2450] = ~(inputs[209]) | (inputs[48]);
    assign layer0_outputs[2451] = 1'b1;
    assign layer0_outputs[2452] = (inputs[135]) & ~(inputs[162]);
    assign layer0_outputs[2453] = 1'b0;
    assign layer0_outputs[2454] = (inputs[179]) | (inputs[158]);
    assign layer0_outputs[2455] = ~(inputs[83]);
    assign layer0_outputs[2456] = ~(inputs[95]) | (inputs[253]);
    assign layer0_outputs[2457] = ~((inputs[3]) | (inputs[53]));
    assign layer0_outputs[2458] = inputs[195];
    assign layer0_outputs[2459] = (inputs[101]) ^ (inputs[0]);
    assign layer0_outputs[2460] = ~(inputs[62]) | (inputs[248]);
    assign layer0_outputs[2461] = ~((inputs[170]) | (inputs[69]));
    assign layer0_outputs[2462] = 1'b0;
    assign layer0_outputs[2463] = ~((inputs[169]) & (inputs[140]));
    assign layer0_outputs[2464] = ~((inputs[144]) & (inputs[102]));
    assign layer0_outputs[2465] = (inputs[48]) | (inputs[241]);
    assign layer0_outputs[2466] = (inputs[228]) & (inputs[251]);
    assign layer0_outputs[2467] = ~((inputs[188]) | (inputs[96]));
    assign layer0_outputs[2468] = (inputs[244]) & ~(inputs[102]);
    assign layer0_outputs[2469] = ~(inputs[4]) | (inputs[211]);
    assign layer0_outputs[2470] = ~(inputs[187]);
    assign layer0_outputs[2471] = (inputs[25]) ^ (inputs[220]);
    assign layer0_outputs[2472] = (inputs[197]) | (inputs[178]);
    assign layer0_outputs[2473] = (inputs[23]) ^ (inputs[101]);
    assign layer0_outputs[2474] = ~((inputs[172]) | (inputs[146]));
    assign layer0_outputs[2475] = ~(inputs[225]) | (inputs[173]);
    assign layer0_outputs[2476] = inputs[141];
    assign layer0_outputs[2477] = ~((inputs[250]) & (inputs[31]));
    assign layer0_outputs[2478] = (inputs[21]) & ~(inputs[53]);
    assign layer0_outputs[2479] = (inputs[208]) ^ (inputs[87]);
    assign layer0_outputs[2480] = inputs[186];
    assign layer0_outputs[2481] = inputs[186];
    assign layer0_outputs[2482] = inputs[61];
    assign layer0_outputs[2483] = (inputs[252]) | (inputs[65]);
    assign layer0_outputs[2484] = ~(inputs[239]);
    assign layer0_outputs[2485] = 1'b0;
    assign layer0_outputs[2486] = 1'b1;
    assign layer0_outputs[2487] = ~(inputs[222]) | (inputs[125]);
    assign layer0_outputs[2488] = ~(inputs[183]);
    assign layer0_outputs[2489] = (inputs[129]) & (inputs[39]);
    assign layer0_outputs[2490] = (inputs[147]) & ~(inputs[122]);
    assign layer0_outputs[2491] = 1'b0;
    assign layer0_outputs[2492] = ~((inputs[196]) & (inputs[20]));
    assign layer0_outputs[2493] = (inputs[244]) & ~(inputs[207]);
    assign layer0_outputs[2494] = inputs[101];
    assign layer0_outputs[2495] = ~(inputs[84]) | (inputs[19]);
    assign layer0_outputs[2496] = (inputs[219]) & ~(inputs[138]);
    assign layer0_outputs[2497] = (inputs[155]) & ~(inputs[1]);
    assign layer0_outputs[2498] = 1'b0;
    assign layer0_outputs[2499] = inputs[71];
    assign layer0_outputs[2500] = (inputs[140]) | (inputs[172]);
    assign layer0_outputs[2501] = inputs[7];
    assign layer0_outputs[2502] = ~(inputs[164]) | (inputs[95]);
    assign layer0_outputs[2503] = ~(inputs[150]);
    assign layer0_outputs[2504] = inputs[132];
    assign layer0_outputs[2505] = inputs[234];
    assign layer0_outputs[2506] = (inputs[200]) & ~(inputs[48]);
    assign layer0_outputs[2507] = 1'b1;
    assign layer0_outputs[2508] = (inputs[159]) & ~(inputs[6]);
    assign layer0_outputs[2509] = ~(inputs[244]);
    assign layer0_outputs[2510] = 1'b1;
    assign layer0_outputs[2511] = (inputs[66]) & (inputs[67]);
    assign layer0_outputs[2512] = ~((inputs[80]) | (inputs[251]));
    assign layer0_outputs[2513] = ~(inputs[72]);
    assign layer0_outputs[2514] = inputs[119];
    assign layer0_outputs[2515] = (inputs[109]) ^ (inputs[90]);
    assign layer0_outputs[2516] = 1'b1;
    assign layer0_outputs[2517] = ~(inputs[25]) | (inputs[234]);
    assign layer0_outputs[2518] = ~(inputs[223]) | (inputs[38]);
    assign layer0_outputs[2519] = ~(inputs[18]) | (inputs[203]);
    assign layer0_outputs[2520] = ~(inputs[203]) | (inputs[180]);
    assign layer0_outputs[2521] = ~(inputs[191]) | (inputs[72]);
    assign layer0_outputs[2522] = ~(inputs[14]);
    assign layer0_outputs[2523] = (inputs[164]) & (inputs[246]);
    assign layer0_outputs[2524] = ~(inputs[107]);
    assign layer0_outputs[2525] = (inputs[169]) | (inputs[82]);
    assign layer0_outputs[2526] = ~((inputs[120]) | (inputs[128]));
    assign layer0_outputs[2527] = inputs[155];
    assign layer0_outputs[2528] = 1'b0;
    assign layer0_outputs[2529] = (inputs[40]) | (inputs[126]);
    assign layer0_outputs[2530] = ~(inputs[104]) | (inputs[49]);
    assign layer0_outputs[2531] = ~(inputs[146]) | (inputs[249]);
    assign layer0_outputs[2532] = ~((inputs[10]) | (inputs[157]));
    assign layer0_outputs[2533] = (inputs[253]) & ~(inputs[125]);
    assign layer0_outputs[2534] = ~((inputs[27]) | (inputs[136]));
    assign layer0_outputs[2535] = 1'b0;
    assign layer0_outputs[2536] = (inputs[11]) & ~(inputs[166]);
    assign layer0_outputs[2537] = 1'b0;
    assign layer0_outputs[2538] = (inputs[223]) ^ (inputs[75]);
    assign layer0_outputs[2539] = ~(inputs[210]);
    assign layer0_outputs[2540] = ~(inputs[138]);
    assign layer0_outputs[2541] = inputs[49];
    assign layer0_outputs[2542] = ~((inputs[197]) | (inputs[189]));
    assign layer0_outputs[2543] = (inputs[186]) & ~(inputs[223]);
    assign layer0_outputs[2544] = ~(inputs[153]) | (inputs[24]);
    assign layer0_outputs[2545] = ~(inputs[173]);
    assign layer0_outputs[2546] = inputs[120];
    assign layer0_outputs[2547] = (inputs[29]) | (inputs[222]);
    assign layer0_outputs[2548] = ~(inputs[113]);
    assign layer0_outputs[2549] = ~(inputs[213]);
    assign layer0_outputs[2550] = (inputs[35]) & ~(inputs[51]);
    assign layer0_outputs[2551] = ~((inputs[196]) | (inputs[229]));
    assign layer0_outputs[2552] = 1'b0;
    assign layer0_outputs[2553] = (inputs[156]) | (inputs[133]);
    assign layer0_outputs[2554] = (inputs[129]) | (inputs[149]);
    assign layer0_outputs[2555] = ~((inputs[14]) & (inputs[81]));
    assign layer0_outputs[2556] = 1'b1;
    assign layer0_outputs[2557] = 1'b1;
    assign layer0_outputs[2558] = 1'b1;
    assign layer0_outputs[2559] = ~(inputs[113]) | (inputs[49]);
    assign layer0_outputs[2560] = ~(inputs[188]) | (inputs[220]);
    assign layer0_outputs[2561] = 1'b1;
    assign layer0_outputs[2562] = ~(inputs[167]) | (inputs[98]);
    assign layer0_outputs[2563] = inputs[61];
    assign layer0_outputs[2564] = inputs[229];
    assign layer0_outputs[2565] = (inputs[145]) & ~(inputs[161]);
    assign layer0_outputs[2566] = ~(inputs[39]);
    assign layer0_outputs[2567] = ~((inputs[111]) ^ (inputs[182]));
    assign layer0_outputs[2568] = ~((inputs[167]) ^ (inputs[113]));
    assign layer0_outputs[2569] = (inputs[156]) | (inputs[174]);
    assign layer0_outputs[2570] = ~((inputs[169]) & (inputs[8]));
    assign layer0_outputs[2571] = (inputs[107]) & (inputs[12]);
    assign layer0_outputs[2572] = ~((inputs[147]) | (inputs[87]));
    assign layer0_outputs[2573] = ~(inputs[119]);
    assign layer0_outputs[2574] = 1'b1;
    assign layer0_outputs[2575] = inputs[242];
    assign layer0_outputs[2576] = ~(inputs[113]);
    assign layer0_outputs[2577] = (inputs[96]) & (inputs[239]);
    assign layer0_outputs[2578] = (inputs[138]) & ~(inputs[158]);
    assign layer0_outputs[2579] = ~(inputs[147]);
    assign layer0_outputs[2580] = 1'b1;
    assign layer0_outputs[2581] = inputs[128];
    assign layer0_outputs[2582] = inputs[148];
    assign layer0_outputs[2583] = (inputs[152]) & ~(inputs[73]);
    assign layer0_outputs[2584] = ~((inputs[109]) | (inputs[214]));
    assign layer0_outputs[2585] = ~(inputs[127]);
    assign layer0_outputs[2586] = ~(inputs[60]);
    assign layer0_outputs[2587] = 1'b1;
    assign layer0_outputs[2588] = inputs[45];
    assign layer0_outputs[2589] = ~(inputs[253]);
    assign layer0_outputs[2590] = ~(inputs[87]) | (inputs[1]);
    assign layer0_outputs[2591] = (inputs[63]) ^ (inputs[95]);
    assign layer0_outputs[2592] = (inputs[189]) & ~(inputs[22]);
    assign layer0_outputs[2593] = ~((inputs[83]) | (inputs[195]));
    assign layer0_outputs[2594] = ~(inputs[174]);
    assign layer0_outputs[2595] = (inputs[103]) & (inputs[157]);
    assign layer0_outputs[2596] = (inputs[60]) ^ (inputs[215]);
    assign layer0_outputs[2597] = inputs[197];
    assign layer0_outputs[2598] = ~(inputs[185]);
    assign layer0_outputs[2599] = (inputs[211]) & (inputs[61]);
    assign layer0_outputs[2600] = (inputs[71]) ^ (inputs[71]);
    assign layer0_outputs[2601] = inputs[190];
    assign layer0_outputs[2602] = (inputs[248]) | (inputs[131]);
    assign layer0_outputs[2603] = inputs[24];
    assign layer0_outputs[2604] = inputs[235];
    assign layer0_outputs[2605] = ~((inputs[218]) | (inputs[70]));
    assign layer0_outputs[2606] = 1'b1;
    assign layer0_outputs[2607] = inputs[171];
    assign layer0_outputs[2608] = (inputs[64]) & (inputs[55]);
    assign layer0_outputs[2609] = (inputs[123]) ^ (inputs[50]);
    assign layer0_outputs[2610] = 1'b0;
    assign layer0_outputs[2611] = ~((inputs[213]) | (inputs[163]));
    assign layer0_outputs[2612] = (inputs[171]) & ~(inputs[249]);
    assign layer0_outputs[2613] = ~((inputs[20]) | (inputs[205]));
    assign layer0_outputs[2614] = (inputs[145]) & ~(inputs[11]);
    assign layer0_outputs[2615] = 1'b1;
    assign layer0_outputs[2616] = (inputs[244]) ^ (inputs[136]);
    assign layer0_outputs[2617] = ~(inputs[7]);
    assign layer0_outputs[2618] = (inputs[177]) ^ (inputs[220]);
    assign layer0_outputs[2619] = (inputs[160]) & (inputs[15]);
    assign layer0_outputs[2620] = ~((inputs[43]) ^ (inputs[133]));
    assign layer0_outputs[2621] = ~(inputs[93]) | (inputs[32]);
    assign layer0_outputs[2622] = (inputs[107]) & ~(inputs[210]);
    assign layer0_outputs[2623] = inputs[165];
    assign layer0_outputs[2624] = 1'b0;
    assign layer0_outputs[2625] = inputs[59];
    assign layer0_outputs[2626] = 1'b1;
    assign layer0_outputs[2627] = ~((inputs[236]) | (inputs[47]));
    assign layer0_outputs[2628] = 1'b1;
    assign layer0_outputs[2629] = ~(inputs[82]) | (inputs[128]);
    assign layer0_outputs[2630] = ~(inputs[69]) | (inputs[219]);
    assign layer0_outputs[2631] = (inputs[158]) ^ (inputs[64]);
    assign layer0_outputs[2632] = (inputs[102]) & ~(inputs[184]);
    assign layer0_outputs[2633] = ~((inputs[109]) ^ (inputs[215]));
    assign layer0_outputs[2634] = (inputs[24]) & ~(inputs[178]);
    assign layer0_outputs[2635] = ~(inputs[57]);
    assign layer0_outputs[2636] = (inputs[152]) | (inputs[67]);
    assign layer0_outputs[2637] = inputs[2];
    assign layer0_outputs[2638] = (inputs[81]) & ~(inputs[140]);
    assign layer0_outputs[2639] = (inputs[157]) | (inputs[42]);
    assign layer0_outputs[2640] = 1'b0;
    assign layer0_outputs[2641] = ~(inputs[244]) | (inputs[158]);
    assign layer0_outputs[2642] = 1'b1;
    assign layer0_outputs[2643] = ~((inputs[89]) ^ (inputs[252]));
    assign layer0_outputs[2644] = inputs[165];
    assign layer0_outputs[2645] = (inputs[86]) | (inputs[61]);
    assign layer0_outputs[2646] = ~(inputs[41]);
    assign layer0_outputs[2647] = ~(inputs[22]) | (inputs[108]);
    assign layer0_outputs[2648] = ~(inputs[120]);
    assign layer0_outputs[2649] = ~((inputs[122]) & (inputs[224]));
    assign layer0_outputs[2650] = inputs[2];
    assign layer0_outputs[2651] = 1'b0;
    assign layer0_outputs[2652] = ~((inputs[98]) & (inputs[168]));
    assign layer0_outputs[2653] = ~((inputs[69]) & (inputs[33]));
    assign layer0_outputs[2654] = ~((inputs[254]) & (inputs[225]));
    assign layer0_outputs[2655] = (inputs[145]) ^ (inputs[1]);
    assign layer0_outputs[2656] = ~((inputs[212]) & (inputs[6]));
    assign layer0_outputs[2657] = (inputs[35]) & ~(inputs[76]);
    assign layer0_outputs[2658] = ~((inputs[36]) & (inputs[10]));
    assign layer0_outputs[2659] = ~(inputs[195]) | (inputs[98]);
    assign layer0_outputs[2660] = (inputs[189]) ^ (inputs[49]);
    assign layer0_outputs[2661] = (inputs[77]) ^ (inputs[9]);
    assign layer0_outputs[2662] = inputs[72];
    assign layer0_outputs[2663] = inputs[202];
    assign layer0_outputs[2664] = (inputs[95]) ^ (inputs[110]);
    assign layer0_outputs[2665] = inputs[187];
    assign layer0_outputs[2666] = 1'b0;
    assign layer0_outputs[2667] = ~(inputs[38]);
    assign layer0_outputs[2668] = (inputs[146]) ^ (inputs[218]);
    assign layer0_outputs[2669] = inputs[66];
    assign layer0_outputs[2670] = ~((inputs[175]) | (inputs[218]));
    assign layer0_outputs[2671] = ~((inputs[61]) & (inputs[199]));
    assign layer0_outputs[2672] = 1'b0;
    assign layer0_outputs[2673] = inputs[188];
    assign layer0_outputs[2674] = inputs[8];
    assign layer0_outputs[2675] = ~(inputs[93]) | (inputs[102]);
    assign layer0_outputs[2676] = (inputs[239]) & ~(inputs[68]);
    assign layer0_outputs[2677] = ~((inputs[245]) & (inputs[125]));
    assign layer0_outputs[2678] = (inputs[226]) ^ (inputs[136]);
    assign layer0_outputs[2679] = (inputs[121]) & ~(inputs[126]);
    assign layer0_outputs[2680] = inputs[170];
    assign layer0_outputs[2681] = 1'b1;
    assign layer0_outputs[2682] = inputs[220];
    assign layer0_outputs[2683] = ~((inputs[168]) | (inputs[182]));
    assign layer0_outputs[2684] = 1'b1;
    assign layer0_outputs[2685] = (inputs[28]) ^ (inputs[62]);
    assign layer0_outputs[2686] = ~((inputs[150]) ^ (inputs[204]));
    assign layer0_outputs[2687] = (inputs[235]) | (inputs[80]);
    assign layer0_outputs[2688] = ~(inputs[65]) | (inputs[100]);
    assign layer0_outputs[2689] = (inputs[185]) ^ (inputs[106]);
    assign layer0_outputs[2690] = (inputs[146]) & ~(inputs[204]);
    assign layer0_outputs[2691] = 1'b1;
    assign layer0_outputs[2692] = (inputs[38]) & ~(inputs[199]);
    assign layer0_outputs[2693] = 1'b1;
    assign layer0_outputs[2694] = 1'b0;
    assign layer0_outputs[2695] = (inputs[228]) & ~(inputs[165]);
    assign layer0_outputs[2696] = (inputs[154]) & (inputs[82]);
    assign layer0_outputs[2697] = ~((inputs[67]) | (inputs[155]));
    assign layer0_outputs[2698] = (inputs[96]) & ~(inputs[7]);
    assign layer0_outputs[2699] = 1'b0;
    assign layer0_outputs[2700] = ~(inputs[231]) | (inputs[1]);
    assign layer0_outputs[2701] = ~((inputs[205]) | (inputs[181]));
    assign layer0_outputs[2702] = 1'b1;
    assign layer0_outputs[2703] = ~(inputs[133]);
    assign layer0_outputs[2704] = inputs[22];
    assign layer0_outputs[2705] = inputs[238];
    assign layer0_outputs[2706] = 1'b1;
    assign layer0_outputs[2707] = ~((inputs[204]) & (inputs[206]));
    assign layer0_outputs[2708] = (inputs[68]) ^ (inputs[3]);
    assign layer0_outputs[2709] = inputs[178];
    assign layer0_outputs[2710] = inputs[123];
    assign layer0_outputs[2711] = 1'b1;
    assign layer0_outputs[2712] = 1'b1;
    assign layer0_outputs[2713] = inputs[62];
    assign layer0_outputs[2714] = ~((inputs[181]) ^ (inputs[48]));
    assign layer0_outputs[2715] = (inputs[10]) & ~(inputs[90]);
    assign layer0_outputs[2716] = ~(inputs[133]) | (inputs[211]);
    assign layer0_outputs[2717] = (inputs[12]) & (inputs[43]);
    assign layer0_outputs[2718] = (inputs[239]) | (inputs[174]);
    assign layer0_outputs[2719] = 1'b1;
    assign layer0_outputs[2720] = 1'b1;
    assign layer0_outputs[2721] = inputs[242];
    assign layer0_outputs[2722] = ~(inputs[80]);
    assign layer0_outputs[2723] = inputs[235];
    assign layer0_outputs[2724] = ~((inputs[62]) & (inputs[232]));
    assign layer0_outputs[2725] = 1'b1;
    assign layer0_outputs[2726] = (inputs[32]) ^ (inputs[63]);
    assign layer0_outputs[2727] = (inputs[72]) & ~(inputs[209]);
    assign layer0_outputs[2728] = 1'b0;
    assign layer0_outputs[2729] = ~((inputs[229]) | (inputs[143]));
    assign layer0_outputs[2730] = ~(inputs[152]) | (inputs[176]);
    assign layer0_outputs[2731] = ~((inputs[132]) | (inputs[102]));
    assign layer0_outputs[2732] = 1'b0;
    assign layer0_outputs[2733] = ~((inputs[161]) | (inputs[254]));
    assign layer0_outputs[2734] = (inputs[177]) | (inputs[201]);
    assign layer0_outputs[2735] = 1'b1;
    assign layer0_outputs[2736] = (inputs[182]) & ~(inputs[112]);
    assign layer0_outputs[2737] = ~(inputs[239]) | (inputs[55]);
    assign layer0_outputs[2738] = ~(inputs[151]) | (inputs[57]);
    assign layer0_outputs[2739] = (inputs[73]) | (inputs[162]);
    assign layer0_outputs[2740] = inputs[111];
    assign layer0_outputs[2741] = ~(inputs[160]);
    assign layer0_outputs[2742] = ~((inputs[138]) ^ (inputs[84]));
    assign layer0_outputs[2743] = ~((inputs[141]) | (inputs[153]));
    assign layer0_outputs[2744] = (inputs[113]) & ~(inputs[113]);
    assign layer0_outputs[2745] = ~(inputs[76]);
    assign layer0_outputs[2746] = ~((inputs[209]) & (inputs[154]));
    assign layer0_outputs[2747] = (inputs[145]) ^ (inputs[228]);
    assign layer0_outputs[2748] = ~((inputs[72]) | (inputs[179]));
    assign layer0_outputs[2749] = inputs[33];
    assign layer0_outputs[2750] = (inputs[41]) & ~(inputs[184]);
    assign layer0_outputs[2751] = ~(inputs[186]) | (inputs[191]);
    assign layer0_outputs[2752] = 1'b1;
    assign layer0_outputs[2753] = inputs[187];
    assign layer0_outputs[2754] = ~((inputs[107]) & (inputs[148]));
    assign layer0_outputs[2755] = ~((inputs[138]) | (inputs[180]));
    assign layer0_outputs[2756] = (inputs[108]) & ~(inputs[27]);
    assign layer0_outputs[2757] = inputs[184];
    assign layer0_outputs[2758] = ~((inputs[17]) & (inputs[244]));
    assign layer0_outputs[2759] = 1'b1;
    assign layer0_outputs[2760] = (inputs[49]) ^ (inputs[4]);
    assign layer0_outputs[2761] = 1'b1;
    assign layer0_outputs[2762] = ~(inputs[74]) | (inputs[99]);
    assign layer0_outputs[2763] = ~(inputs[221]) | (inputs[97]);
    assign layer0_outputs[2764] = inputs[128];
    assign layer0_outputs[2765] = ~((inputs[30]) & (inputs[64]));
    assign layer0_outputs[2766] = ~((inputs[191]) & (inputs[57]));
    assign layer0_outputs[2767] = inputs[206];
    assign layer0_outputs[2768] = 1'b0;
    assign layer0_outputs[2769] = ~(inputs[172]) | (inputs[109]);
    assign layer0_outputs[2770] = ~((inputs[69]) & (inputs[83]));
    assign layer0_outputs[2771] = 1'b0;
    assign layer0_outputs[2772] = ~(inputs[255]) | (inputs[183]);
    assign layer0_outputs[2773] = ~(inputs[250]) | (inputs[110]);
    assign layer0_outputs[2774] = (inputs[47]) | (inputs[93]);
    assign layer0_outputs[2775] = ~((inputs[74]) & (inputs[14]));
    assign layer0_outputs[2776] = 1'b0;
    assign layer0_outputs[2777] = inputs[230];
    assign layer0_outputs[2778] = ~((inputs[212]) & (inputs[235]));
    assign layer0_outputs[2779] = ~((inputs[240]) ^ (inputs[183]));
    assign layer0_outputs[2780] = inputs[62];
    assign layer0_outputs[2781] = ~((inputs[217]) | (inputs[145]));
    assign layer0_outputs[2782] = 1'b1;
    assign layer0_outputs[2783] = (inputs[182]) & ~(inputs[54]);
    assign layer0_outputs[2784] = (inputs[122]) & ~(inputs[152]);
    assign layer0_outputs[2785] = ~(inputs[92]) | (inputs[192]);
    assign layer0_outputs[2786] = 1'b0;
    assign layer0_outputs[2787] = (inputs[19]) & (inputs[235]);
    assign layer0_outputs[2788] = ~(inputs[131]) | (inputs[87]);
    assign layer0_outputs[2789] = ~((inputs[135]) ^ (inputs[210]));
    assign layer0_outputs[2790] = ~(inputs[225]) | (inputs[184]);
    assign layer0_outputs[2791] = ~((inputs[7]) | (inputs[218]));
    assign layer0_outputs[2792] = ~(inputs[169]);
    assign layer0_outputs[2793] = (inputs[241]) & ~(inputs[241]);
    assign layer0_outputs[2794] = ~(inputs[166]) | (inputs[52]);
    assign layer0_outputs[2795] = (inputs[54]) & ~(inputs[149]);
    assign layer0_outputs[2796] = (inputs[200]) & ~(inputs[134]);
    assign layer0_outputs[2797] = ~((inputs[225]) | (inputs[98]));
    assign layer0_outputs[2798] = ~((inputs[211]) ^ (inputs[16]));
    assign layer0_outputs[2799] = (inputs[163]) | (inputs[176]);
    assign layer0_outputs[2800] = ~((inputs[155]) | (inputs[40]));
    assign layer0_outputs[2801] = (inputs[83]) & ~(inputs[26]);
    assign layer0_outputs[2802] = ~((inputs[96]) & (inputs[9]));
    assign layer0_outputs[2803] = (inputs[112]) & ~(inputs[237]);
    assign layer0_outputs[2804] = inputs[93];
    assign layer0_outputs[2805] = ~((inputs[143]) ^ (inputs[135]));
    assign layer0_outputs[2806] = ~(inputs[142]) | (inputs[173]);
    assign layer0_outputs[2807] = ~((inputs[206]) & (inputs[224]));
    assign layer0_outputs[2808] = 1'b0;
    assign layer0_outputs[2809] = (inputs[78]) | (inputs[38]);
    assign layer0_outputs[2810] = ~((inputs[96]) & (inputs[151]));
    assign layer0_outputs[2811] = ~(inputs[120]) | (inputs[240]);
    assign layer0_outputs[2812] = (inputs[78]) & ~(inputs[3]);
    assign layer0_outputs[2813] = inputs[34];
    assign layer0_outputs[2814] = inputs[183];
    assign layer0_outputs[2815] = ~(inputs[152]) | (inputs[134]);
    assign layer0_outputs[2816] = ~(inputs[184]) | (inputs[130]);
    assign layer0_outputs[2817] = ~(inputs[78]) | (inputs[51]);
    assign layer0_outputs[2818] = inputs[196];
    assign layer0_outputs[2819] = ~(inputs[108]);
    assign layer0_outputs[2820] = ~(inputs[170]);
    assign layer0_outputs[2821] = 1'b1;
    assign layer0_outputs[2822] = ~(inputs[217]);
    assign layer0_outputs[2823] = ~((inputs[211]) & (inputs[52]));
    assign layer0_outputs[2824] = inputs[179];
    assign layer0_outputs[2825] = 1'b1;
    assign layer0_outputs[2826] = (inputs[106]) ^ (inputs[126]);
    assign layer0_outputs[2827] = inputs[184];
    assign layer0_outputs[2828] = (inputs[78]) | (inputs[40]);
    assign layer0_outputs[2829] = (inputs[6]) | (inputs[31]);
    assign layer0_outputs[2830] = inputs[139];
    assign layer0_outputs[2831] = (inputs[194]) & ~(inputs[124]);
    assign layer0_outputs[2832] = (inputs[235]) | (inputs[2]);
    assign layer0_outputs[2833] = ~((inputs[199]) & (inputs[53]));
    assign layer0_outputs[2834] = (inputs[117]) & ~(inputs[202]);
    assign layer0_outputs[2835] = inputs[18];
    assign layer0_outputs[2836] = ~(inputs[141]);
    assign layer0_outputs[2837] = ~(inputs[40]) | (inputs[158]);
    assign layer0_outputs[2838] = inputs[124];
    assign layer0_outputs[2839] = ~(inputs[119]);
    assign layer0_outputs[2840] = ~((inputs[131]) | (inputs[98]));
    assign layer0_outputs[2841] = ~(inputs[184]) | (inputs[118]);
    assign layer0_outputs[2842] = (inputs[88]) & ~(inputs[175]);
    assign layer0_outputs[2843] = ~(inputs[109]) | (inputs[105]);
    assign layer0_outputs[2844] = ~(inputs[12]) | (inputs[67]);
    assign layer0_outputs[2845] = ~(inputs[141]) | (inputs[248]);
    assign layer0_outputs[2846] = ~(inputs[225]);
    assign layer0_outputs[2847] = inputs[155];
    assign layer0_outputs[2848] = 1'b0;
    assign layer0_outputs[2849] = 1'b1;
    assign layer0_outputs[2850] = inputs[116];
    assign layer0_outputs[2851] = ~(inputs[23]) | (inputs[108]);
    assign layer0_outputs[2852] = ~(inputs[114]);
    assign layer0_outputs[2853] = 1'b0;
    assign layer0_outputs[2854] = ~(inputs[92]);
    assign layer0_outputs[2855] = ~(inputs[38]);
    assign layer0_outputs[2856] = inputs[253];
    assign layer0_outputs[2857] = 1'b1;
    assign layer0_outputs[2858] = ~((inputs[131]) ^ (inputs[32]));
    assign layer0_outputs[2859] = ~(inputs[69]);
    assign layer0_outputs[2860] = (inputs[32]) & (inputs[70]);
    assign layer0_outputs[2861] = inputs[9];
    assign layer0_outputs[2862] = ~(inputs[162]);
    assign layer0_outputs[2863] = inputs[176];
    assign layer0_outputs[2864] = (inputs[168]) ^ (inputs[0]);
    assign layer0_outputs[2865] = ~(inputs[86]) | (inputs[58]);
    assign layer0_outputs[2866] = (inputs[10]) ^ (inputs[103]);
    assign layer0_outputs[2867] = ~(inputs[93]) | (inputs[107]);
    assign layer0_outputs[2868] = (inputs[0]) & (inputs[78]);
    assign layer0_outputs[2869] = ~((inputs[115]) & (inputs[177]));
    assign layer0_outputs[2870] = ~((inputs[8]) | (inputs[109]));
    assign layer0_outputs[2871] = ~(inputs[247]) | (inputs[207]);
    assign layer0_outputs[2872] = (inputs[115]) | (inputs[40]);
    assign layer0_outputs[2873] = ~(inputs[227]);
    assign layer0_outputs[2874] = (inputs[212]) & (inputs[224]);
    assign layer0_outputs[2875] = ~(inputs[59]) | (inputs[178]);
    assign layer0_outputs[2876] = (inputs[16]) | (inputs[52]);
    assign layer0_outputs[2877] = ~((inputs[202]) | (inputs[140]));
    assign layer0_outputs[2878] = ~((inputs[146]) | (inputs[22]));
    assign layer0_outputs[2879] = ~((inputs[174]) | (inputs[30]));
    assign layer0_outputs[2880] = ~((inputs[97]) & (inputs[43]));
    assign layer0_outputs[2881] = 1'b1;
    assign layer0_outputs[2882] = ~((inputs[198]) & (inputs[245]));
    assign layer0_outputs[2883] = (inputs[52]) | (inputs[16]);
    assign layer0_outputs[2884] = ~(inputs[18]) | (inputs[7]);
    assign layer0_outputs[2885] = ~((inputs[84]) | (inputs[217]));
    assign layer0_outputs[2886] = 1'b0;
    assign layer0_outputs[2887] = ~(inputs[44]);
    assign layer0_outputs[2888] = inputs[138];
    assign layer0_outputs[2889] = (inputs[234]) & ~(inputs[70]);
    assign layer0_outputs[2890] = (inputs[222]) & ~(inputs[176]);
    assign layer0_outputs[2891] = inputs[59];
    assign layer0_outputs[2892] = (inputs[226]) | (inputs[154]);
    assign layer0_outputs[2893] = (inputs[5]) & ~(inputs[48]);
    assign layer0_outputs[2894] = (inputs[63]) & (inputs[124]);
    assign layer0_outputs[2895] = ~(inputs[84]);
    assign layer0_outputs[2896] = ~(inputs[241]) | (inputs[249]);
    assign layer0_outputs[2897] = (inputs[213]) & ~(inputs[18]);
    assign layer0_outputs[2898] = (inputs[60]) & ~(inputs[239]);
    assign layer0_outputs[2899] = ~(inputs[221]) | (inputs[24]);
    assign layer0_outputs[2900] = (inputs[80]) ^ (inputs[95]);
    assign layer0_outputs[2901] = ~((inputs[94]) ^ (inputs[110]));
    assign layer0_outputs[2902] = 1'b0;
    assign layer0_outputs[2903] = (inputs[24]) | (inputs[33]);
    assign layer0_outputs[2904] = (inputs[98]) & ~(inputs[192]);
    assign layer0_outputs[2905] = 1'b0;
    assign layer0_outputs[2906] = (inputs[92]) | (inputs[80]);
    assign layer0_outputs[2907] = ~((inputs[189]) & (inputs[91]));
    assign layer0_outputs[2908] = inputs[214];
    assign layer0_outputs[2909] = inputs[146];
    assign layer0_outputs[2910] = 1'b1;
    assign layer0_outputs[2911] = 1'b1;
    assign layer0_outputs[2912] = inputs[123];
    assign layer0_outputs[2913] = ~(inputs[78]) | (inputs[86]);
    assign layer0_outputs[2914] = (inputs[154]) & ~(inputs[1]);
    assign layer0_outputs[2915] = ~(inputs[49]) | (inputs[193]);
    assign layer0_outputs[2916] = 1'b1;
    assign layer0_outputs[2917] = ~(inputs[97]) | (inputs[176]);
    assign layer0_outputs[2918] = ~(inputs[131]) | (inputs[234]);
    assign layer0_outputs[2919] = 1'b0;
    assign layer0_outputs[2920] = ~(inputs[178]);
    assign layer0_outputs[2921] = (inputs[142]) & ~(inputs[168]);
    assign layer0_outputs[2922] = ~(inputs[215]) | (inputs[205]);
    assign layer0_outputs[2923] = (inputs[203]) & ~(inputs[217]);
    assign layer0_outputs[2924] = ~((inputs[152]) ^ (inputs[191]));
    assign layer0_outputs[2925] = ~(inputs[79]) | (inputs[20]);
    assign layer0_outputs[2926] = 1'b0;
    assign layer0_outputs[2927] = inputs[156];
    assign layer0_outputs[2928] = inputs[132];
    assign layer0_outputs[2929] = 1'b1;
    assign layer0_outputs[2930] = (inputs[194]) | (inputs[198]);
    assign layer0_outputs[2931] = ~(inputs[66]);
    assign layer0_outputs[2932] = ~((inputs[6]) & (inputs[84]));
    assign layer0_outputs[2933] = inputs[206];
    assign layer0_outputs[2934] = (inputs[33]) & ~(inputs[84]);
    assign layer0_outputs[2935] = (inputs[82]) & ~(inputs[194]);
    assign layer0_outputs[2936] = (inputs[238]) & (inputs[123]);
    assign layer0_outputs[2937] = (inputs[197]) & ~(inputs[146]);
    assign layer0_outputs[2938] = inputs[151];
    assign layer0_outputs[2939] = 1'b0;
    assign layer0_outputs[2940] = ~((inputs[218]) & (inputs[70]));
    assign layer0_outputs[2941] = ~(inputs[11]) | (inputs[196]);
    assign layer0_outputs[2942] = (inputs[222]) ^ (inputs[40]);
    assign layer0_outputs[2943] = 1'b1;
    assign layer0_outputs[2944] = (inputs[229]) ^ (inputs[103]);
    assign layer0_outputs[2945] = ~(inputs[52]) | (inputs[227]);
    assign layer0_outputs[2946] = ~(inputs[153]) | (inputs[162]);
    assign layer0_outputs[2947] = (inputs[171]) & (inputs[147]);
    assign layer0_outputs[2948] = (inputs[11]) | (inputs[125]);
    assign layer0_outputs[2949] = (inputs[237]) & ~(inputs[95]);
    assign layer0_outputs[2950] = (inputs[95]) | (inputs[187]);
    assign layer0_outputs[2951] = ~(inputs[187]);
    assign layer0_outputs[2952] = (inputs[194]) & ~(inputs[32]);
    assign layer0_outputs[2953] = inputs[31];
    assign layer0_outputs[2954] = (inputs[230]) & (inputs[138]);
    assign layer0_outputs[2955] = (inputs[111]) ^ (inputs[203]);
    assign layer0_outputs[2956] = ~((inputs[213]) | (inputs[208]));
    assign layer0_outputs[2957] = 1'b0;
    assign layer0_outputs[2958] = (inputs[142]) ^ (inputs[223]);
    assign layer0_outputs[2959] = ~((inputs[95]) & (inputs[242]));
    assign layer0_outputs[2960] = inputs[150];
    assign layer0_outputs[2961] = ~(inputs[153]) | (inputs[208]);
    assign layer0_outputs[2962] = (inputs[20]) | (inputs[108]);
    assign layer0_outputs[2963] = (inputs[202]) ^ (inputs[69]);
    assign layer0_outputs[2964] = (inputs[95]) & ~(inputs[123]);
    assign layer0_outputs[2965] = 1'b0;
    assign layer0_outputs[2966] = inputs[21];
    assign layer0_outputs[2967] = (inputs[171]) & ~(inputs[25]);
    assign layer0_outputs[2968] = ~(inputs[197]);
    assign layer0_outputs[2969] = ~(inputs[56]) | (inputs[167]);
    assign layer0_outputs[2970] = inputs[150];
    assign layer0_outputs[2971] = (inputs[171]) | (inputs[116]);
    assign layer0_outputs[2972] = ~(inputs[61]);
    assign layer0_outputs[2973] = (inputs[133]) & ~(inputs[204]);
    assign layer0_outputs[2974] = (inputs[57]) | (inputs[249]);
    assign layer0_outputs[2975] = (inputs[9]) ^ (inputs[44]);
    assign layer0_outputs[2976] = ~((inputs[13]) ^ (inputs[181]));
    assign layer0_outputs[2977] = (inputs[201]) | (inputs[193]);
    assign layer0_outputs[2978] = (inputs[127]) ^ (inputs[152]);
    assign layer0_outputs[2979] = (inputs[90]) & ~(inputs[15]);
    assign layer0_outputs[2980] = ~((inputs[55]) | (inputs[186]));
    assign layer0_outputs[2981] = inputs[254];
    assign layer0_outputs[2982] = ~((inputs[232]) ^ (inputs[159]));
    assign layer0_outputs[2983] = 1'b0;
    assign layer0_outputs[2984] = (inputs[73]) & ~(inputs[15]);
    assign layer0_outputs[2985] = 1'b0;
    assign layer0_outputs[2986] = 1'b1;
    assign layer0_outputs[2987] = (inputs[143]) & (inputs[172]);
    assign layer0_outputs[2988] = ~(inputs[110]) | (inputs[88]);
    assign layer0_outputs[2989] = ~((inputs[140]) & (inputs[181]));
    assign layer0_outputs[2990] = (inputs[27]) ^ (inputs[88]);
    assign layer0_outputs[2991] = (inputs[76]) | (inputs[94]);
    assign layer0_outputs[2992] = ~(inputs[182]);
    assign layer0_outputs[2993] = ~(inputs[99]);
    assign layer0_outputs[2994] = ~((inputs[228]) | (inputs[105]));
    assign layer0_outputs[2995] = (inputs[195]) & ~(inputs[218]);
    assign layer0_outputs[2996] = 1'b0;
    assign layer0_outputs[2997] = ~((inputs[13]) ^ (inputs[25]));
    assign layer0_outputs[2998] = 1'b0;
    assign layer0_outputs[2999] = ~((inputs[190]) | (inputs[249]));
    assign layer0_outputs[3000] = inputs[206];
    assign layer0_outputs[3001] = ~(inputs[166]);
    assign layer0_outputs[3002] = ~(inputs[198]);
    assign layer0_outputs[3003] = ~(inputs[107]) | (inputs[175]);
    assign layer0_outputs[3004] = inputs[111];
    assign layer0_outputs[3005] = 1'b1;
    assign layer0_outputs[3006] = ~(inputs[204]);
    assign layer0_outputs[3007] = 1'b1;
    assign layer0_outputs[3008] = inputs[88];
    assign layer0_outputs[3009] = (inputs[137]) & (inputs[37]);
    assign layer0_outputs[3010] = 1'b1;
    assign layer0_outputs[3011] = 1'b0;
    assign layer0_outputs[3012] = (inputs[158]) & ~(inputs[93]);
    assign layer0_outputs[3013] = ~(inputs[18]);
    assign layer0_outputs[3014] = 1'b0;
    assign layer0_outputs[3015] = ~((inputs[173]) & (inputs[166]));
    assign layer0_outputs[3016] = (inputs[39]) & (inputs[185]);
    assign layer0_outputs[3017] = (inputs[211]) | (inputs[75]);
    assign layer0_outputs[3018] = ~((inputs[134]) ^ (inputs[176]));
    assign layer0_outputs[3019] = inputs[133];
    assign layer0_outputs[3020] = (inputs[29]) ^ (inputs[203]);
    assign layer0_outputs[3021] = ~(inputs[138]) | (inputs[96]);
    assign layer0_outputs[3022] = ~(inputs[124]);
    assign layer0_outputs[3023] = ~(inputs[147]);
    assign layer0_outputs[3024] = ~(inputs[131]);
    assign layer0_outputs[3025] = ~(inputs[0]) | (inputs[7]);
    assign layer0_outputs[3026] = inputs[44];
    assign layer0_outputs[3027] = (inputs[76]) | (inputs[146]);
    assign layer0_outputs[3028] = (inputs[230]) ^ (inputs[138]);
    assign layer0_outputs[3029] = 1'b1;
    assign layer0_outputs[3030] = inputs[103];
    assign layer0_outputs[3031] = (inputs[89]) & ~(inputs[131]);
    assign layer0_outputs[3032] = inputs[63];
    assign layer0_outputs[3033] = (inputs[12]) & ~(inputs[97]);
    assign layer0_outputs[3034] = ~((inputs[214]) | (inputs[207]));
    assign layer0_outputs[3035] = inputs[54];
    assign layer0_outputs[3036] = ~(inputs[167]) | (inputs[141]);
    assign layer0_outputs[3037] = inputs[228];
    assign layer0_outputs[3038] = ~(inputs[89]) | (inputs[120]);
    assign layer0_outputs[3039] = (inputs[119]) ^ (inputs[16]);
    assign layer0_outputs[3040] = (inputs[220]) & ~(inputs[196]);
    assign layer0_outputs[3041] = ~(inputs[153]);
    assign layer0_outputs[3042] = 1'b0;
    assign layer0_outputs[3043] = (inputs[195]) & ~(inputs[178]);
    assign layer0_outputs[3044] = (inputs[129]) ^ (inputs[29]);
    assign layer0_outputs[3045] = ~(inputs[124]) | (inputs[52]);
    assign layer0_outputs[3046] = inputs[232];
    assign layer0_outputs[3047] = ~(inputs[7]);
    assign layer0_outputs[3048] = ~(inputs[139]) | (inputs[90]);
    assign layer0_outputs[3049] = (inputs[54]) & ~(inputs[129]);
    assign layer0_outputs[3050] = ~(inputs[138]) | (inputs[54]);
    assign layer0_outputs[3051] = ~(inputs[114]) | (inputs[164]);
    assign layer0_outputs[3052] = 1'b1;
    assign layer0_outputs[3053] = ~((inputs[85]) | (inputs[15]));
    assign layer0_outputs[3054] = (inputs[226]) | (inputs[18]);
    assign layer0_outputs[3055] = ~((inputs[237]) & (inputs[208]));
    assign layer0_outputs[3056] = 1'b0;
    assign layer0_outputs[3057] = ~(inputs[154]) | (inputs[47]);
    assign layer0_outputs[3058] = (inputs[248]) & ~(inputs[29]);
    assign layer0_outputs[3059] = ~((inputs[106]) | (inputs[148]));
    assign layer0_outputs[3060] = inputs[111];
    assign layer0_outputs[3061] = ~(inputs[243]);
    assign layer0_outputs[3062] = 1'b0;
    assign layer0_outputs[3063] = ~(inputs[36]) | (inputs[146]);
    assign layer0_outputs[3064] = (inputs[180]) & ~(inputs[246]);
    assign layer0_outputs[3065] = ~(inputs[152]);
    assign layer0_outputs[3066] = (inputs[193]) & ~(inputs[71]);
    assign layer0_outputs[3067] = inputs[3];
    assign layer0_outputs[3068] = ~(inputs[117]);
    assign layer0_outputs[3069] = (inputs[127]) ^ (inputs[46]);
    assign layer0_outputs[3070] = ~(inputs[2]) | (inputs[229]);
    assign layer0_outputs[3071] = ~(inputs[84]) | (inputs[121]);
    assign layer0_outputs[3072] = ~((inputs[112]) | (inputs[121]));
    assign layer0_outputs[3073] = ~(inputs[228]);
    assign layer0_outputs[3074] = (inputs[128]) & ~(inputs[219]);
    assign layer0_outputs[3075] = ~(inputs[194]) | (inputs[41]);
    assign layer0_outputs[3076] = (inputs[168]) | (inputs[46]);
    assign layer0_outputs[3077] = (inputs[104]) & ~(inputs[48]);
    assign layer0_outputs[3078] = inputs[56];
    assign layer0_outputs[3079] = ~((inputs[130]) & (inputs[119]));
    assign layer0_outputs[3080] = ~(inputs[4]) | (inputs[188]);
    assign layer0_outputs[3081] = inputs[121];
    assign layer0_outputs[3082] = ~((inputs[62]) | (inputs[77]));
    assign layer0_outputs[3083] = 1'b0;
    assign layer0_outputs[3084] = (inputs[16]) & ~(inputs[14]);
    assign layer0_outputs[3085] = ~(inputs[186]) | (inputs[89]);
    assign layer0_outputs[3086] = ~((inputs[208]) ^ (inputs[238]));
    assign layer0_outputs[3087] = (inputs[88]) | (inputs[81]);
    assign layer0_outputs[3088] = 1'b1;
    assign layer0_outputs[3089] = (inputs[164]) | (inputs[38]);
    assign layer0_outputs[3090] = (inputs[64]) & (inputs[20]);
    assign layer0_outputs[3091] = (inputs[181]) & (inputs[82]);
    assign layer0_outputs[3092] = (inputs[176]) | (inputs[18]);
    assign layer0_outputs[3093] = (inputs[100]) & (inputs[195]);
    assign layer0_outputs[3094] = ~(inputs[77]);
    assign layer0_outputs[3095] = 1'b1;
    assign layer0_outputs[3096] = (inputs[211]) ^ (inputs[209]);
    assign layer0_outputs[3097] = ~(inputs[134]);
    assign layer0_outputs[3098] = 1'b0;
    assign layer0_outputs[3099] = (inputs[191]) & ~(inputs[189]);
    assign layer0_outputs[3100] = 1'b0;
    assign layer0_outputs[3101] = (inputs[223]) ^ (inputs[25]);
    assign layer0_outputs[3102] = (inputs[106]) | (inputs[207]);
    assign layer0_outputs[3103] = 1'b1;
    assign layer0_outputs[3104] = ~(inputs[18]);
    assign layer0_outputs[3105] = ~((inputs[19]) ^ (inputs[246]));
    assign layer0_outputs[3106] = inputs[163];
    assign layer0_outputs[3107] = (inputs[17]) & ~(inputs[34]);
    assign layer0_outputs[3108] = ~(inputs[51]);
    assign layer0_outputs[3109] = (inputs[11]) | (inputs[8]);
    assign layer0_outputs[3110] = 1'b1;
    assign layer0_outputs[3111] = ~(inputs[47]) | (inputs[22]);
    assign layer0_outputs[3112] = ~(inputs[21]) | (inputs[194]);
    assign layer0_outputs[3113] = (inputs[87]) & ~(inputs[172]);
    assign layer0_outputs[3114] = ~((inputs[245]) & (inputs[116]));
    assign layer0_outputs[3115] = (inputs[7]) | (inputs[145]);
    assign layer0_outputs[3116] = inputs[231];
    assign layer0_outputs[3117] = 1'b0;
    assign layer0_outputs[3118] = ~((inputs[129]) ^ (inputs[167]));
    assign layer0_outputs[3119] = inputs[138];
    assign layer0_outputs[3120] = (inputs[125]) | (inputs[104]);
    assign layer0_outputs[3121] = (inputs[91]) | (inputs[3]);
    assign layer0_outputs[3122] = ~(inputs[100]) | (inputs[16]);
    assign layer0_outputs[3123] = (inputs[29]) & ~(inputs[228]);
    assign layer0_outputs[3124] = inputs[144];
    assign layer0_outputs[3125] = ~((inputs[173]) | (inputs[190]));
    assign layer0_outputs[3126] = ~((inputs[205]) ^ (inputs[69]));
    assign layer0_outputs[3127] = ~((inputs[4]) & (inputs[113]));
    assign layer0_outputs[3128] = ~((inputs[61]) | (inputs[180]));
    assign layer0_outputs[3129] = ~(inputs[25]) | (inputs[51]);
    assign layer0_outputs[3130] = ~(inputs[80]) | (inputs[121]);
    assign layer0_outputs[3131] = ~((inputs[90]) | (inputs[212]));
    assign layer0_outputs[3132] = (inputs[115]) & (inputs[59]);
    assign layer0_outputs[3133] = inputs[70];
    assign layer0_outputs[3134] = ~((inputs[49]) | (inputs[243]));
    assign layer0_outputs[3135] = ~(inputs[221]);
    assign layer0_outputs[3136] = 1'b1;
    assign layer0_outputs[3137] = ~(inputs[104]);
    assign layer0_outputs[3138] = 1'b0;
    assign layer0_outputs[3139] = ~(inputs[246]);
    assign layer0_outputs[3140] = ~(inputs[30]) | (inputs[28]);
    assign layer0_outputs[3141] = ~((inputs[168]) & (inputs[154]));
    assign layer0_outputs[3142] = 1'b1;
    assign layer0_outputs[3143] = inputs[122];
    assign layer0_outputs[3144] = ~(inputs[52]);
    assign layer0_outputs[3145] = inputs[218];
    assign layer0_outputs[3146] = ~(inputs[63]);
    assign layer0_outputs[3147] = (inputs[230]) ^ (inputs[199]);
    assign layer0_outputs[3148] = (inputs[193]) & ~(inputs[223]);
    assign layer0_outputs[3149] = ~((inputs[6]) | (inputs[100]));
    assign layer0_outputs[3150] = (inputs[12]) ^ (inputs[190]);
    assign layer0_outputs[3151] = ~((inputs[127]) & (inputs[226]));
    assign layer0_outputs[3152] = ~(inputs[116]) | (inputs[188]);
    assign layer0_outputs[3153] = inputs[146];
    assign layer0_outputs[3154] = 1'b1;
    assign layer0_outputs[3155] = (inputs[178]) & ~(inputs[232]);
    assign layer0_outputs[3156] = ~(inputs[114]);
    assign layer0_outputs[3157] = 1'b0;
    assign layer0_outputs[3158] = 1'b1;
    assign layer0_outputs[3159] = ~((inputs[24]) | (inputs[113]));
    assign layer0_outputs[3160] = (inputs[193]) & ~(inputs[5]);
    assign layer0_outputs[3161] = (inputs[220]) ^ (inputs[137]);
    assign layer0_outputs[3162] = (inputs[190]) | (inputs[159]);
    assign layer0_outputs[3163] = (inputs[112]) & (inputs[197]);
    assign layer0_outputs[3164] = ~(inputs[176]);
    assign layer0_outputs[3165] = 1'b1;
    assign layer0_outputs[3166] = ~((inputs[66]) & (inputs[196]));
    assign layer0_outputs[3167] = 1'b0;
    assign layer0_outputs[3168] = (inputs[245]) & ~(inputs[41]);
    assign layer0_outputs[3169] = inputs[121];
    assign layer0_outputs[3170] = ~((inputs[181]) | (inputs[77]));
    assign layer0_outputs[3171] = ~(inputs[173]);
    assign layer0_outputs[3172] = ~(inputs[214]) | (inputs[112]);
    assign layer0_outputs[3173] = ~((inputs[91]) | (inputs[90]));
    assign layer0_outputs[3174] = inputs[91];
    assign layer0_outputs[3175] = 1'b1;
    assign layer0_outputs[3176] = ~((inputs[64]) | (inputs[134]));
    assign layer0_outputs[3177] = ~(inputs[85]) | (inputs[239]);
    assign layer0_outputs[3178] = 1'b1;
    assign layer0_outputs[3179] = (inputs[78]) & ~(inputs[243]);
    assign layer0_outputs[3180] = ~((inputs[239]) | (inputs[211]));
    assign layer0_outputs[3181] = ~(inputs[35]);
    assign layer0_outputs[3182] = 1'b0;
    assign layer0_outputs[3183] = ~((inputs[223]) & (inputs[177]));
    assign layer0_outputs[3184] = 1'b0;
    assign layer0_outputs[3185] = (inputs[67]) | (inputs[214]);
    assign layer0_outputs[3186] = (inputs[255]) & ~(inputs[160]);
    assign layer0_outputs[3187] = ~(inputs[116]);
    assign layer0_outputs[3188] = ~(inputs[7]) | (inputs[26]);
    assign layer0_outputs[3189] = ~(inputs[16]);
    assign layer0_outputs[3190] = ~((inputs[112]) & (inputs[244]));
    assign layer0_outputs[3191] = inputs[187];
    assign layer0_outputs[3192] = 1'b1;
    assign layer0_outputs[3193] = ~(inputs[112]) | (inputs[31]);
    assign layer0_outputs[3194] = (inputs[206]) & ~(inputs[172]);
    assign layer0_outputs[3195] = ~((inputs[219]) | (inputs[180]));
    assign layer0_outputs[3196] = 1'b1;
    assign layer0_outputs[3197] = ~(inputs[106]) | (inputs[75]);
    assign layer0_outputs[3198] = 1'b1;
    assign layer0_outputs[3199] = ~(inputs[129]) | (inputs[98]);
    assign layer0_outputs[3200] = 1'b0;
    assign layer0_outputs[3201] = (inputs[181]) & ~(inputs[100]);
    assign layer0_outputs[3202] = ~(inputs[227]);
    assign layer0_outputs[3203] = 1'b0;
    assign layer0_outputs[3204] = ~(inputs[167]);
    assign layer0_outputs[3205] = ~(inputs[177]);
    assign layer0_outputs[3206] = (inputs[187]) & ~(inputs[200]);
    assign layer0_outputs[3207] = ~((inputs[116]) | (inputs[140]));
    assign layer0_outputs[3208] = ~(inputs[197]) | (inputs[221]);
    assign layer0_outputs[3209] = ~(inputs[34]);
    assign layer0_outputs[3210] = ~(inputs[204]);
    assign layer0_outputs[3211] = (inputs[255]) & ~(inputs[22]);
    assign layer0_outputs[3212] = ~((inputs[16]) | (inputs[120]));
    assign layer0_outputs[3213] = ~((inputs[131]) ^ (inputs[202]));
    assign layer0_outputs[3214] = (inputs[139]) & ~(inputs[145]);
    assign layer0_outputs[3215] = 1'b1;
    assign layer0_outputs[3216] = (inputs[121]) & (inputs[216]);
    assign layer0_outputs[3217] = 1'b0;
    assign layer0_outputs[3218] = ~(inputs[74]) | (inputs[78]);
    assign layer0_outputs[3219] = ~(inputs[197]) | (inputs[235]);
    assign layer0_outputs[3220] = (inputs[153]) & ~(inputs[11]);
    assign layer0_outputs[3221] = (inputs[202]) | (inputs[40]);
    assign layer0_outputs[3222] = (inputs[54]) ^ (inputs[92]);
    assign layer0_outputs[3223] = inputs[188];
    assign layer0_outputs[3224] = ~((inputs[38]) & (inputs[143]));
    assign layer0_outputs[3225] = inputs[52];
    assign layer0_outputs[3226] = (inputs[229]) ^ (inputs[112]);
    assign layer0_outputs[3227] = inputs[140];
    assign layer0_outputs[3228] = 1'b1;
    assign layer0_outputs[3229] = 1'b1;
    assign layer0_outputs[3230] = ~(inputs[17]);
    assign layer0_outputs[3231] = ~(inputs[125]);
    assign layer0_outputs[3232] = (inputs[166]) | (inputs[189]);
    assign layer0_outputs[3233] = ~(inputs[144]);
    assign layer0_outputs[3234] = inputs[134];
    assign layer0_outputs[3235] = ~(inputs[147]);
    assign layer0_outputs[3236] = (inputs[12]) & ~(inputs[237]);
    assign layer0_outputs[3237] = ~(inputs[67]) | (inputs[27]);
    assign layer0_outputs[3238] = ~(inputs[154]) | (inputs[78]);
    assign layer0_outputs[3239] = 1'b0;
    assign layer0_outputs[3240] = ~(inputs[105]);
    assign layer0_outputs[3241] = ~(inputs[179]) | (inputs[250]);
    assign layer0_outputs[3242] = ~(inputs[112]) | (inputs[73]);
    assign layer0_outputs[3243] = (inputs[58]) & ~(inputs[199]);
    assign layer0_outputs[3244] = (inputs[55]) & ~(inputs[16]);
    assign layer0_outputs[3245] = ~((inputs[8]) | (inputs[83]));
    assign layer0_outputs[3246] = ~(inputs[164]);
    assign layer0_outputs[3247] = ~(inputs[25]) | (inputs[210]);
    assign layer0_outputs[3248] = 1'b1;
    assign layer0_outputs[3249] = inputs[167];
    assign layer0_outputs[3250] = inputs[81];
    assign layer0_outputs[3251] = ~((inputs[147]) | (inputs[116]));
    assign layer0_outputs[3252] = 1'b0;
    assign layer0_outputs[3253] = inputs[99];
    assign layer0_outputs[3254] = (inputs[230]) & ~(inputs[139]);
    assign layer0_outputs[3255] = ~((inputs[18]) & (inputs[80]));
    assign layer0_outputs[3256] = ~(inputs[112]);
    assign layer0_outputs[3257] = ~(inputs[148]);
    assign layer0_outputs[3258] = ~((inputs[156]) & (inputs[164]));
    assign layer0_outputs[3259] = ~(inputs[230]);
    assign layer0_outputs[3260] = 1'b0;
    assign layer0_outputs[3261] = (inputs[99]) & ~(inputs[8]);
    assign layer0_outputs[3262] = ~(inputs[33]);
    assign layer0_outputs[3263] = inputs[102];
    assign layer0_outputs[3264] = (inputs[209]) | (inputs[207]);
    assign layer0_outputs[3265] = 1'b1;
    assign layer0_outputs[3266] = ~((inputs[98]) ^ (inputs[103]));
    assign layer0_outputs[3267] = ~(inputs[14]);
    assign layer0_outputs[3268] = ~(inputs[122]) | (inputs[141]);
    assign layer0_outputs[3269] = inputs[9];
    assign layer0_outputs[3270] = (inputs[12]) & (inputs[0]);
    assign layer0_outputs[3271] = inputs[214];
    assign layer0_outputs[3272] = ~(inputs[52]) | (inputs[254]);
    assign layer0_outputs[3273] = (inputs[239]) & ~(inputs[160]);
    assign layer0_outputs[3274] = ~((inputs[208]) & (inputs[255]));
    assign layer0_outputs[3275] = (inputs[24]) & (inputs[103]);
    assign layer0_outputs[3276] = ~((inputs[233]) | (inputs[60]));
    assign layer0_outputs[3277] = ~(inputs[132]) | (inputs[88]);
    assign layer0_outputs[3278] = (inputs[133]) & ~(inputs[231]);
    assign layer0_outputs[3279] = ~((inputs[28]) | (inputs[114]));
    assign layer0_outputs[3280] = ~((inputs[230]) | (inputs[46]));
    assign layer0_outputs[3281] = (inputs[37]) & ~(inputs[6]);
    assign layer0_outputs[3282] = ~((inputs[175]) | (inputs[163]));
    assign layer0_outputs[3283] = ~(inputs[26]) | (inputs[16]);
    assign layer0_outputs[3284] = ~(inputs[20]);
    assign layer0_outputs[3285] = ~((inputs[111]) ^ (inputs[106]));
    assign layer0_outputs[3286] = (inputs[128]) & ~(inputs[242]);
    assign layer0_outputs[3287] = inputs[246];
    assign layer0_outputs[3288] = ~(inputs[105]) | (inputs[241]);
    assign layer0_outputs[3289] = 1'b1;
    assign layer0_outputs[3290] = ~(inputs[142]) | (inputs[255]);
    assign layer0_outputs[3291] = (inputs[179]) & ~(inputs[235]);
    assign layer0_outputs[3292] = (inputs[155]) | (inputs[120]);
    assign layer0_outputs[3293] = inputs[243];
    assign layer0_outputs[3294] = 1'b1;
    assign layer0_outputs[3295] = 1'b1;
    assign layer0_outputs[3296] = 1'b1;
    assign layer0_outputs[3297] = 1'b1;
    assign layer0_outputs[3298] = ~((inputs[183]) & (inputs[155]));
    assign layer0_outputs[3299] = (inputs[63]) & ~(inputs[111]);
    assign layer0_outputs[3300] = ~(inputs[34]);
    assign layer0_outputs[3301] = (inputs[184]) & (inputs[186]);
    assign layer0_outputs[3302] = (inputs[135]) & ~(inputs[196]);
    assign layer0_outputs[3303] = (inputs[250]) ^ (inputs[24]);
    assign layer0_outputs[3304] = ~(inputs[177]) | (inputs[245]);
    assign layer0_outputs[3305] = ~(inputs[132]);
    assign layer0_outputs[3306] = inputs[184];
    assign layer0_outputs[3307] = (inputs[158]) & (inputs[162]);
    assign layer0_outputs[3308] = (inputs[180]) & ~(inputs[232]);
    assign layer0_outputs[3309] = (inputs[102]) | (inputs[49]);
    assign layer0_outputs[3310] = 1'b0;
    assign layer0_outputs[3311] = inputs[162];
    assign layer0_outputs[3312] = ~(inputs[157]) | (inputs[199]);
    assign layer0_outputs[3313] = ~((inputs[119]) ^ (inputs[250]));
    assign layer0_outputs[3314] = inputs[153];
    assign layer0_outputs[3315] = inputs[89];
    assign layer0_outputs[3316] = ~(inputs[250]) | (inputs[207]);
    assign layer0_outputs[3317] = inputs[116];
    assign layer0_outputs[3318] = ~((inputs[173]) & (inputs[9]));
    assign layer0_outputs[3319] = inputs[88];
    assign layer0_outputs[3320] = (inputs[67]) ^ (inputs[126]);
    assign layer0_outputs[3321] = (inputs[82]) & ~(inputs[5]);
    assign layer0_outputs[3322] = (inputs[170]) & ~(inputs[19]);
    assign layer0_outputs[3323] = ~(inputs[94]);
    assign layer0_outputs[3324] = 1'b1;
    assign layer0_outputs[3325] = (inputs[205]) | (inputs[248]);
    assign layer0_outputs[3326] = ~(inputs[70]) | (inputs[228]);
    assign layer0_outputs[3327] = 1'b1;
    assign layer0_outputs[3328] = 1'b0;
    assign layer0_outputs[3329] = ~(inputs[39]);
    assign layer0_outputs[3330] = ~((inputs[108]) | (inputs[152]));
    assign layer0_outputs[3331] = ~((inputs[190]) | (inputs[131]));
    assign layer0_outputs[3332] = ~(inputs[107]) | (inputs[22]);
    assign layer0_outputs[3333] = ~(inputs[68]) | (inputs[79]);
    assign layer0_outputs[3334] = (inputs[32]) | (inputs[185]);
    assign layer0_outputs[3335] = inputs[9];
    assign layer0_outputs[3336] = 1'b0;
    assign layer0_outputs[3337] = ~(inputs[225]);
    assign layer0_outputs[3338] = ~((inputs[231]) ^ (inputs[115]));
    assign layer0_outputs[3339] = ~(inputs[226]);
    assign layer0_outputs[3340] = ~((inputs[85]) | (inputs[219]));
    assign layer0_outputs[3341] = inputs[209];
    assign layer0_outputs[3342] = inputs[63];
    assign layer0_outputs[3343] = inputs[153];
    assign layer0_outputs[3344] = (inputs[25]) & (inputs[55]);
    assign layer0_outputs[3345] = ~((inputs[27]) | (inputs[57]));
    assign layer0_outputs[3346] = 1'b1;
    assign layer0_outputs[3347] = inputs[207];
    assign layer0_outputs[3348] = (inputs[19]) ^ (inputs[19]);
    assign layer0_outputs[3349] = (inputs[37]) ^ (inputs[77]);
    assign layer0_outputs[3350] = (inputs[31]) ^ (inputs[114]);
    assign layer0_outputs[3351] = ~((inputs[75]) & (inputs[36]));
    assign layer0_outputs[3352] = 1'b1;
    assign layer0_outputs[3353] = ~((inputs[2]) | (inputs[129]));
    assign layer0_outputs[3354] = 1'b0;
    assign layer0_outputs[3355] = ~(inputs[30]);
    assign layer0_outputs[3356] = ~((inputs[241]) | (inputs[212]));
    assign layer0_outputs[3357] = (inputs[81]) & (inputs[114]);
    assign layer0_outputs[3358] = 1'b1;
    assign layer0_outputs[3359] = 1'b0;
    assign layer0_outputs[3360] = (inputs[193]) | (inputs[160]);
    assign layer0_outputs[3361] = inputs[218];
    assign layer0_outputs[3362] = ~((inputs[210]) & (inputs[99]));
    assign layer0_outputs[3363] = ~(inputs[162]) | (inputs[97]);
    assign layer0_outputs[3364] = ~(inputs[174]);
    assign layer0_outputs[3365] = (inputs[32]) & ~(inputs[251]);
    assign layer0_outputs[3366] = ~(inputs[19]) | (inputs[135]);
    assign layer0_outputs[3367] = 1'b1;
    assign layer0_outputs[3368] = (inputs[15]) & ~(inputs[140]);
    assign layer0_outputs[3369] = ~(inputs[196]);
    assign layer0_outputs[3370] = ~((inputs[51]) ^ (inputs[245]));
    assign layer0_outputs[3371] = ~((inputs[132]) ^ (inputs[240]));
    assign layer0_outputs[3372] = ~(inputs[161]) | (inputs[220]);
    assign layer0_outputs[3373] = (inputs[244]) & ~(inputs[209]);
    assign layer0_outputs[3374] = (inputs[180]) | (inputs[170]);
    assign layer0_outputs[3375] = 1'b1;
    assign layer0_outputs[3376] = ~(inputs[222]);
    assign layer0_outputs[3377] = ~((inputs[20]) ^ (inputs[97]));
    assign layer0_outputs[3378] = (inputs[72]) & (inputs[121]);
    assign layer0_outputs[3379] = (inputs[130]) | (inputs[82]);
    assign layer0_outputs[3380] = ~(inputs[48]) | (inputs[76]);
    assign layer0_outputs[3381] = ~((inputs[190]) | (inputs[58]));
    assign layer0_outputs[3382] = 1'b1;
    assign layer0_outputs[3383] = 1'b1;
    assign layer0_outputs[3384] = 1'b1;
    assign layer0_outputs[3385] = 1'b0;
    assign layer0_outputs[3386] = (inputs[1]) & ~(inputs[249]);
    assign layer0_outputs[3387] = 1'b1;
    assign layer0_outputs[3388] = ~(inputs[250]) | (inputs[22]);
    assign layer0_outputs[3389] = ~(inputs[24]) | (inputs[10]);
    assign layer0_outputs[3390] = (inputs[80]) & (inputs[109]);
    assign layer0_outputs[3391] = 1'b1;
    assign layer0_outputs[3392] = (inputs[92]) & ~(inputs[210]);
    assign layer0_outputs[3393] = ~((inputs[3]) ^ (inputs[241]));
    assign layer0_outputs[3394] = ~(inputs[6]);
    assign layer0_outputs[3395] = ~((inputs[78]) | (inputs[84]));
    assign layer0_outputs[3396] = (inputs[177]) | (inputs[199]);
    assign layer0_outputs[3397] = ~((inputs[5]) ^ (inputs[233]));
    assign layer0_outputs[3398] = inputs[36];
    assign layer0_outputs[3399] = ~((inputs[130]) | (inputs[23]));
    assign layer0_outputs[3400] = (inputs[53]) & ~(inputs[131]);
    assign layer0_outputs[3401] = inputs[102];
    assign layer0_outputs[3402] = ~(inputs[75]);
    assign layer0_outputs[3403] = ~(inputs[74]);
    assign layer0_outputs[3404] = ~(inputs[66]) | (inputs[178]);
    assign layer0_outputs[3405] = (inputs[135]) ^ (inputs[32]);
    assign layer0_outputs[3406] = (inputs[174]) ^ (inputs[178]);
    assign layer0_outputs[3407] = ~((inputs[223]) & (inputs[2]));
    assign layer0_outputs[3408] = ~(inputs[236]);
    assign layer0_outputs[3409] = ~((inputs[115]) & (inputs[96]));
    assign layer0_outputs[3410] = (inputs[56]) ^ (inputs[174]);
    assign layer0_outputs[3411] = ~(inputs[3]) | (inputs[42]);
    assign layer0_outputs[3412] = inputs[146];
    assign layer0_outputs[3413] = ~(inputs[5]);
    assign layer0_outputs[3414] = inputs[52];
    assign layer0_outputs[3415] = ~((inputs[13]) & (inputs[153]));
    assign layer0_outputs[3416] = (inputs[58]) ^ (inputs[194]);
    assign layer0_outputs[3417] = ~(inputs[23]);
    assign layer0_outputs[3418] = ~(inputs[108]) | (inputs[88]);
    assign layer0_outputs[3419] = (inputs[236]) | (inputs[186]);
    assign layer0_outputs[3420] = ~(inputs[133]);
    assign layer0_outputs[3421] = inputs[100];
    assign layer0_outputs[3422] = inputs[174];
    assign layer0_outputs[3423] = 1'b1;
    assign layer0_outputs[3424] = ~(inputs[171]) | (inputs[179]);
    assign layer0_outputs[3425] = 1'b0;
    assign layer0_outputs[3426] = ~(inputs[187]);
    assign layer0_outputs[3427] = ~((inputs[115]) | (inputs[221]));
    assign layer0_outputs[3428] = (inputs[151]) & ~(inputs[13]);
    assign layer0_outputs[3429] = inputs[84];
    assign layer0_outputs[3430] = (inputs[155]) & ~(inputs[92]);
    assign layer0_outputs[3431] = 1'b0;
    assign layer0_outputs[3432] = (inputs[233]) & ~(inputs[13]);
    assign layer0_outputs[3433] = inputs[76];
    assign layer0_outputs[3434] = (inputs[150]) ^ (inputs[208]);
    assign layer0_outputs[3435] = (inputs[202]) | (inputs[217]);
    assign layer0_outputs[3436] = ~((inputs[2]) | (inputs[27]));
    assign layer0_outputs[3437] = inputs[128];
    assign layer0_outputs[3438] = inputs[124];
    assign layer0_outputs[3439] = ~(inputs[251]) | (inputs[192]);
    assign layer0_outputs[3440] = (inputs[125]) & ~(inputs[229]);
    assign layer0_outputs[3441] = inputs[146];
    assign layer0_outputs[3442] = ~(inputs[75]);
    assign layer0_outputs[3443] = ~(inputs[117]) | (inputs[36]);
    assign layer0_outputs[3444] = (inputs[50]) & (inputs[43]);
    assign layer0_outputs[3445] = ~(inputs[245]);
    assign layer0_outputs[3446] = inputs[243];
    assign layer0_outputs[3447] = ~(inputs[198]) | (inputs[203]);
    assign layer0_outputs[3448] = ~((inputs[207]) & (inputs[146]));
    assign layer0_outputs[3449] = ~(inputs[137]) | (inputs[138]);
    assign layer0_outputs[3450] = ~((inputs[57]) & (inputs[82]));
    assign layer0_outputs[3451] = inputs[175];
    assign layer0_outputs[3452] = ~((inputs[30]) | (inputs[167]));
    assign layer0_outputs[3453] = (inputs[21]) | (inputs[1]);
    assign layer0_outputs[3454] = 1'b0;
    assign layer0_outputs[3455] = (inputs[156]) ^ (inputs[134]);
    assign layer0_outputs[3456] = ~(inputs[136]) | (inputs[99]);
    assign layer0_outputs[3457] = (inputs[214]) | (inputs[248]);
    assign layer0_outputs[3458] = ~((inputs[30]) | (inputs[31]));
    assign layer0_outputs[3459] = 1'b1;
    assign layer0_outputs[3460] = (inputs[111]) ^ (inputs[72]);
    assign layer0_outputs[3461] = 1'b0;
    assign layer0_outputs[3462] = 1'b0;
    assign layer0_outputs[3463] = ~((inputs[177]) & (inputs[111]));
    assign layer0_outputs[3464] = ~((inputs[42]) ^ (inputs[212]));
    assign layer0_outputs[3465] = 1'b0;
    assign layer0_outputs[3466] = (inputs[209]) & ~(inputs[70]);
    assign layer0_outputs[3467] = ~((inputs[229]) & (inputs[219]));
    assign layer0_outputs[3468] = ~(inputs[47]);
    assign layer0_outputs[3469] = (inputs[113]) | (inputs[87]);
    assign layer0_outputs[3470] = (inputs[40]) & ~(inputs[194]);
    assign layer0_outputs[3471] = ~(inputs[72]) | (inputs[67]);
    assign layer0_outputs[3472] = ~((inputs[183]) | (inputs[127]));
    assign layer0_outputs[3473] = ~(inputs[202]);
    assign layer0_outputs[3474] = ~(inputs[169]);
    assign layer0_outputs[3475] = inputs[40];
    assign layer0_outputs[3476] = 1'b0;
    assign layer0_outputs[3477] = (inputs[199]) | (inputs[174]);
    assign layer0_outputs[3478] = (inputs[222]) | (inputs[202]);
    assign layer0_outputs[3479] = ~((inputs[217]) & (inputs[182]));
    assign layer0_outputs[3480] = inputs[145];
    assign layer0_outputs[3481] = (inputs[214]) | (inputs[226]);
    assign layer0_outputs[3482] = (inputs[175]) & (inputs[221]);
    assign layer0_outputs[3483] = ~(inputs[241]) | (inputs[132]);
    assign layer0_outputs[3484] = (inputs[118]) & ~(inputs[133]);
    assign layer0_outputs[3485] = ~((inputs[15]) | (inputs[207]));
    assign layer0_outputs[3486] = (inputs[126]) & (inputs[38]);
    assign layer0_outputs[3487] = (inputs[232]) & (inputs[216]);
    assign layer0_outputs[3488] = ~(inputs[191]) | (inputs[70]);
    assign layer0_outputs[3489] = 1'b1;
    assign layer0_outputs[3490] = 1'b1;
    assign layer0_outputs[3491] = ~((inputs[230]) | (inputs[116]));
    assign layer0_outputs[3492] = ~((inputs[200]) & (inputs[130]));
    assign layer0_outputs[3493] = ~((inputs[171]) & (inputs[108]));
    assign layer0_outputs[3494] = (inputs[237]) | (inputs[116]);
    assign layer0_outputs[3495] = (inputs[242]) | (inputs[32]);
    assign layer0_outputs[3496] = (inputs[53]) | (inputs[193]);
    assign layer0_outputs[3497] = inputs[208];
    assign layer0_outputs[3498] = ~(inputs[2]) | (inputs[8]);
    assign layer0_outputs[3499] = 1'b0;
    assign layer0_outputs[3500] = 1'b0;
    assign layer0_outputs[3501] = (inputs[236]) & ~(inputs[142]);
    assign layer0_outputs[3502] = (inputs[246]) | (inputs[165]);
    assign layer0_outputs[3503] = (inputs[24]) & ~(inputs[218]);
    assign layer0_outputs[3504] = ~(inputs[247]);
    assign layer0_outputs[3505] = ~(inputs[241]) | (inputs[64]);
    assign layer0_outputs[3506] = 1'b0;
    assign layer0_outputs[3507] = ~(inputs[50]) | (inputs[244]);
    assign layer0_outputs[3508] = (inputs[141]) & ~(inputs[165]);
    assign layer0_outputs[3509] = (inputs[43]) | (inputs[76]);
    assign layer0_outputs[3510] = inputs[18];
    assign layer0_outputs[3511] = ~((inputs[105]) | (inputs[48]));
    assign layer0_outputs[3512] = inputs[9];
    assign layer0_outputs[3513] = ~((inputs[97]) | (inputs[71]));
    assign layer0_outputs[3514] = ~(inputs[86]);
    assign layer0_outputs[3515] = (inputs[80]) & ~(inputs[16]);
    assign layer0_outputs[3516] = (inputs[246]) & ~(inputs[40]);
    assign layer0_outputs[3517] = inputs[61];
    assign layer0_outputs[3518] = ~((inputs[30]) ^ (inputs[65]));
    assign layer0_outputs[3519] = ~(inputs[225]) | (inputs[99]);
    assign layer0_outputs[3520] = ~((inputs[2]) ^ (inputs[204]));
    assign layer0_outputs[3521] = 1'b1;
    assign layer0_outputs[3522] = ~(inputs[53]) | (inputs[23]);
    assign layer0_outputs[3523] = ~(inputs[20]) | (inputs[162]);
    assign layer0_outputs[3524] = (inputs[4]) | (inputs[142]);
    assign layer0_outputs[3525] = (inputs[140]) | (inputs[44]);
    assign layer0_outputs[3526] = 1'b0;
    assign layer0_outputs[3527] = 1'b1;
    assign layer0_outputs[3528] = ~(inputs[43]) | (inputs[99]);
    assign layer0_outputs[3529] = (inputs[179]) ^ (inputs[157]);
    assign layer0_outputs[3530] = (inputs[245]) ^ (inputs[209]);
    assign layer0_outputs[3531] = ~(inputs[232]);
    assign layer0_outputs[3532] = inputs[208];
    assign layer0_outputs[3533] = (inputs[77]) & (inputs[99]);
    assign layer0_outputs[3534] = (inputs[253]) & (inputs[111]);
    assign layer0_outputs[3535] = ~(inputs[171]) | (inputs[47]);
    assign layer0_outputs[3536] = (inputs[161]) & ~(inputs[23]);
    assign layer0_outputs[3537] = ~(inputs[126]) | (inputs[160]);
    assign layer0_outputs[3538] = ~((inputs[37]) & (inputs[216]));
    assign layer0_outputs[3539] = ~(inputs[137]) | (inputs[203]);
    assign layer0_outputs[3540] = (inputs[50]) | (inputs[160]);
    assign layer0_outputs[3541] = ~((inputs[159]) | (inputs[38]));
    assign layer0_outputs[3542] = (inputs[222]) | (inputs[218]);
    assign layer0_outputs[3543] = (inputs[118]) | (inputs[154]);
    assign layer0_outputs[3544] = ~((inputs[61]) ^ (inputs[88]));
    assign layer0_outputs[3545] = ~(inputs[176]);
    assign layer0_outputs[3546] = ~(inputs[241]) | (inputs[134]);
    assign layer0_outputs[3547] = (inputs[166]) & ~(inputs[245]);
    assign layer0_outputs[3548] = inputs[207];
    assign layer0_outputs[3549] = 1'b0;
    assign layer0_outputs[3550] = ~(inputs[77]);
    assign layer0_outputs[3551] = ~((inputs[154]) & (inputs[223]));
    assign layer0_outputs[3552] = ~(inputs[189]);
    assign layer0_outputs[3553] = ~(inputs[138]) | (inputs[113]);
    assign layer0_outputs[3554] = ~(inputs[11]);
    assign layer0_outputs[3555] = inputs[27];
    assign layer0_outputs[3556] = ~((inputs[224]) ^ (inputs[29]));
    assign layer0_outputs[3557] = 1'b1;
    assign layer0_outputs[3558] = inputs[38];
    assign layer0_outputs[3559] = (inputs[28]) | (inputs[6]);
    assign layer0_outputs[3560] = 1'b1;
    assign layer0_outputs[3561] = ~((inputs[28]) | (inputs[150]));
    assign layer0_outputs[3562] = ~((inputs[171]) | (inputs[161]));
    assign layer0_outputs[3563] = ~((inputs[195]) | (inputs[96]));
    assign layer0_outputs[3564] = (inputs[141]) & (inputs[7]);
    assign layer0_outputs[3565] = (inputs[204]) & ~(inputs[217]);
    assign layer0_outputs[3566] = ~((inputs[101]) | (inputs[250]));
    assign layer0_outputs[3567] = inputs[196];
    assign layer0_outputs[3568] = 1'b1;
    assign layer0_outputs[3569] = ~(inputs[77]);
    assign layer0_outputs[3570] = (inputs[192]) & (inputs[143]);
    assign layer0_outputs[3571] = (inputs[147]) & ~(inputs[110]);
    assign layer0_outputs[3572] = inputs[238];
    assign layer0_outputs[3573] = 1'b0;
    assign layer0_outputs[3574] = (inputs[146]) | (inputs[154]);
    assign layer0_outputs[3575] = ~(inputs[43]) | (inputs[248]);
    assign layer0_outputs[3576] = (inputs[29]) ^ (inputs[29]);
    assign layer0_outputs[3577] = 1'b1;
    assign layer0_outputs[3578] = inputs[38];
    assign layer0_outputs[3579] = (inputs[132]) & (inputs[30]);
    assign layer0_outputs[3580] = ~((inputs[159]) ^ (inputs[109]));
    assign layer0_outputs[3581] = (inputs[217]) | (inputs[66]);
    assign layer0_outputs[3582] = inputs[128];
    assign layer0_outputs[3583] = inputs[19];
    assign layer0_outputs[3584] = (inputs[166]) & ~(inputs[151]);
    assign layer0_outputs[3585] = (inputs[145]) & (inputs[212]);
    assign layer0_outputs[3586] = ~(inputs[156]) | (inputs[16]);
    assign layer0_outputs[3587] = ~(inputs[153]) | (inputs[217]);
    assign layer0_outputs[3588] = ~(inputs[120]) | (inputs[94]);
    assign layer0_outputs[3589] = (inputs[199]) & ~(inputs[176]);
    assign layer0_outputs[3590] = inputs[197];
    assign layer0_outputs[3591] = ~(inputs[233]);
    assign layer0_outputs[3592] = inputs[188];
    assign layer0_outputs[3593] = (inputs[159]) | (inputs[205]);
    assign layer0_outputs[3594] = ~(inputs[136]) | (inputs[160]);
    assign layer0_outputs[3595] = (inputs[49]) & (inputs[155]);
    assign layer0_outputs[3596] = ~((inputs[235]) | (inputs[89]));
    assign layer0_outputs[3597] = ~((inputs[167]) | (inputs[94]));
    assign layer0_outputs[3598] = 1'b0;
    assign layer0_outputs[3599] = ~(inputs[235]) | (inputs[128]);
    assign layer0_outputs[3600] = (inputs[222]) & ~(inputs[130]);
    assign layer0_outputs[3601] = ~((inputs[120]) ^ (inputs[30]));
    assign layer0_outputs[3602] = (inputs[86]) & ~(inputs[37]);
    assign layer0_outputs[3603] = ~((inputs[54]) | (inputs[204]));
    assign layer0_outputs[3604] = (inputs[79]) | (inputs[57]);
    assign layer0_outputs[3605] = ~(inputs[140]) | (inputs[247]);
    assign layer0_outputs[3606] = ~(inputs[1]) | (inputs[87]);
    assign layer0_outputs[3607] = ~(inputs[10]);
    assign layer0_outputs[3608] = ~(inputs[255]);
    assign layer0_outputs[3609] = ~(inputs[133]) | (inputs[96]);
    assign layer0_outputs[3610] = (inputs[24]) & ~(inputs[225]);
    assign layer0_outputs[3611] = inputs[232];
    assign layer0_outputs[3612] = ~(inputs[119]);
    assign layer0_outputs[3613] = ~((inputs[85]) ^ (inputs[6]));
    assign layer0_outputs[3614] = (inputs[78]) & ~(inputs[255]);
    assign layer0_outputs[3615] = ~((inputs[176]) | (inputs[150]));
    assign layer0_outputs[3616] = ~(inputs[221]);
    assign layer0_outputs[3617] = (inputs[3]) & ~(inputs[117]);
    assign layer0_outputs[3618] = (inputs[11]) & ~(inputs[57]);
    assign layer0_outputs[3619] = ~((inputs[225]) & (inputs[32]));
    assign layer0_outputs[3620] = 1'b0;
    assign layer0_outputs[3621] = (inputs[44]) & ~(inputs[249]);
    assign layer0_outputs[3622] = ~(inputs[17]);
    assign layer0_outputs[3623] = 1'b0;
    assign layer0_outputs[3624] = ~((inputs[9]) & (inputs[46]));
    assign layer0_outputs[3625] = ~((inputs[245]) | (inputs[145]));
    assign layer0_outputs[3626] = ~(inputs[92]) | (inputs[224]);
    assign layer0_outputs[3627] = inputs[113];
    assign layer0_outputs[3628] = ~(inputs[0]) | (inputs[68]);
    assign layer0_outputs[3629] = ~(inputs[69]);
    assign layer0_outputs[3630] = (inputs[1]) & (inputs[50]);
    assign layer0_outputs[3631] = ~(inputs[223]);
    assign layer0_outputs[3632] = ~(inputs[195]) | (inputs[40]);
    assign layer0_outputs[3633] = 1'b0;
    assign layer0_outputs[3634] = 1'b0;
    assign layer0_outputs[3635] = (inputs[142]) & ~(inputs[39]);
    assign layer0_outputs[3636] = (inputs[73]) | (inputs[240]);
    assign layer0_outputs[3637] = (inputs[157]) & ~(inputs[249]);
    assign layer0_outputs[3638] = ~(inputs[76]);
    assign layer0_outputs[3639] = ~(inputs[76]) | (inputs[125]);
    assign layer0_outputs[3640] = ~(inputs[181]);
    assign layer0_outputs[3641] = ~(inputs[138]);
    assign layer0_outputs[3642] = ~(inputs[28]);
    assign layer0_outputs[3643] = ~((inputs[114]) | (inputs[24]));
    assign layer0_outputs[3644] = (inputs[227]) & ~(inputs[246]);
    assign layer0_outputs[3645] = ~((inputs[214]) | (inputs[154]));
    assign layer0_outputs[3646] = (inputs[48]) ^ (inputs[141]);
    assign layer0_outputs[3647] = (inputs[246]) ^ (inputs[164]);
    assign layer0_outputs[3648] = (inputs[167]) & ~(inputs[133]);
    assign layer0_outputs[3649] = ~((inputs[124]) & (inputs[247]));
    assign layer0_outputs[3650] = ~((inputs[129]) & (inputs[103]));
    assign layer0_outputs[3651] = (inputs[128]) ^ (inputs[11]);
    assign layer0_outputs[3652] = (inputs[153]) | (inputs[77]);
    assign layer0_outputs[3653] = ~((inputs[105]) ^ (inputs[104]));
    assign layer0_outputs[3654] = ~(inputs[108]);
    assign layer0_outputs[3655] = ~(inputs[113]) | (inputs[0]);
    assign layer0_outputs[3656] = inputs[137];
    assign layer0_outputs[3657] = (inputs[116]) & (inputs[48]);
    assign layer0_outputs[3658] = inputs[45];
    assign layer0_outputs[3659] = ~(inputs[55]) | (inputs[155]);
    assign layer0_outputs[3660] = ~(inputs[24]);
    assign layer0_outputs[3661] = 1'b0;
    assign layer0_outputs[3662] = ~(inputs[235]);
    assign layer0_outputs[3663] = ~((inputs[84]) | (inputs[173]));
    assign layer0_outputs[3664] = ~(inputs[109]);
    assign layer0_outputs[3665] = (inputs[84]) & (inputs[195]);
    assign layer0_outputs[3666] = ~(inputs[73]) | (inputs[166]);
    assign layer0_outputs[3667] = (inputs[204]) | (inputs[187]);
    assign layer0_outputs[3668] = ~((inputs[37]) | (inputs[120]));
    assign layer0_outputs[3669] = ~((inputs[172]) ^ (inputs[243]));
    assign layer0_outputs[3670] = (inputs[88]) & ~(inputs[45]);
    assign layer0_outputs[3671] = 1'b0;
    assign layer0_outputs[3672] = ~(inputs[111]);
    assign layer0_outputs[3673] = inputs[120];
    assign layer0_outputs[3674] = inputs[215];
    assign layer0_outputs[3675] = ~(inputs[47]) | (inputs[118]);
    assign layer0_outputs[3676] = inputs[241];
    assign layer0_outputs[3677] = 1'b1;
    assign layer0_outputs[3678] = 1'b1;
    assign layer0_outputs[3679] = ~(inputs[245]);
    assign layer0_outputs[3680] = inputs[72];
    assign layer0_outputs[3681] = ~(inputs[30]);
    assign layer0_outputs[3682] = inputs[139];
    assign layer0_outputs[3683] = (inputs[104]) & ~(inputs[138]);
    assign layer0_outputs[3684] = inputs[120];
    assign layer0_outputs[3685] = ~((inputs[122]) & (inputs[59]));
    assign layer0_outputs[3686] = ~(inputs[95]);
    assign layer0_outputs[3687] = ~(inputs[156]) | (inputs[224]);
    assign layer0_outputs[3688] = (inputs[14]) | (inputs[150]);
    assign layer0_outputs[3689] = (inputs[124]) & ~(inputs[202]);
    assign layer0_outputs[3690] = ~((inputs[238]) | (inputs[25]));
    assign layer0_outputs[3691] = (inputs[114]) & ~(inputs[133]);
    assign layer0_outputs[3692] = (inputs[160]) & (inputs[101]);
    assign layer0_outputs[3693] = ~((inputs[33]) ^ (inputs[108]));
    assign layer0_outputs[3694] = inputs[143];
    assign layer0_outputs[3695] = 1'b1;
    assign layer0_outputs[3696] = (inputs[152]) & (inputs[122]);
    assign layer0_outputs[3697] = inputs[140];
    assign layer0_outputs[3698] = (inputs[194]) & (inputs[23]);
    assign layer0_outputs[3699] = ~((inputs[168]) | (inputs[26]));
    assign layer0_outputs[3700] = ~(inputs[204]) | (inputs[3]);
    assign layer0_outputs[3701] = (inputs[179]) ^ (inputs[36]);
    assign layer0_outputs[3702] = inputs[247];
    assign layer0_outputs[3703] = 1'b0;
    assign layer0_outputs[3704] = ~(inputs[58]);
    assign layer0_outputs[3705] = inputs[197];
    assign layer0_outputs[3706] = inputs[119];
    assign layer0_outputs[3707] = 1'b0;
    assign layer0_outputs[3708] = inputs[247];
    assign layer0_outputs[3709] = ~((inputs[190]) | (inputs[224]));
    assign layer0_outputs[3710] = ~(inputs[193]) | (inputs[67]);
    assign layer0_outputs[3711] = ~((inputs[0]) | (inputs[80]));
    assign layer0_outputs[3712] = ~((inputs[121]) & (inputs[139]));
    assign layer0_outputs[3713] = 1'b1;
    assign layer0_outputs[3714] = (inputs[84]) & ~(inputs[172]);
    assign layer0_outputs[3715] = (inputs[13]) & (inputs[144]);
    assign layer0_outputs[3716] = (inputs[105]) ^ (inputs[182]);
    assign layer0_outputs[3717] = (inputs[227]) & ~(inputs[79]);
    assign layer0_outputs[3718] = ~(inputs[111]) | (inputs[39]);
    assign layer0_outputs[3719] = inputs[172];
    assign layer0_outputs[3720] = ~((inputs[103]) | (inputs[187]));
    assign layer0_outputs[3721] = ~(inputs[59]);
    assign layer0_outputs[3722] = ~((inputs[77]) & (inputs[12]));
    assign layer0_outputs[3723] = inputs[89];
    assign layer0_outputs[3724] = ~((inputs[181]) | (inputs[2]));
    assign layer0_outputs[3725] = ~((inputs[181]) | (inputs[222]));
    assign layer0_outputs[3726] = ~(inputs[135]);
    assign layer0_outputs[3727] = ~(inputs[119]);
    assign layer0_outputs[3728] = inputs[190];
    assign layer0_outputs[3729] = (inputs[48]) & (inputs[40]);
    assign layer0_outputs[3730] = (inputs[58]) & (inputs[222]);
    assign layer0_outputs[3731] = ~((inputs[232]) ^ (inputs[127]));
    assign layer0_outputs[3732] = (inputs[132]) & ~(inputs[202]);
    assign layer0_outputs[3733] = inputs[175];
    assign layer0_outputs[3734] = ~(inputs[215]);
    assign layer0_outputs[3735] = ~(inputs[189]);
    assign layer0_outputs[3736] = (inputs[155]) & ~(inputs[16]);
    assign layer0_outputs[3737] = (inputs[226]) & (inputs[42]);
    assign layer0_outputs[3738] = ~(inputs[185]);
    assign layer0_outputs[3739] = inputs[148];
    assign layer0_outputs[3740] = ~(inputs[62]) | (inputs[224]);
    assign layer0_outputs[3741] = inputs[90];
    assign layer0_outputs[3742] = (inputs[241]) & (inputs[103]);
    assign layer0_outputs[3743] = inputs[207];
    assign layer0_outputs[3744] = (inputs[133]) & ~(inputs[114]);
    assign layer0_outputs[3745] = 1'b0;
    assign layer0_outputs[3746] = ~(inputs[252]) | (inputs[135]);
    assign layer0_outputs[3747] = ~((inputs[135]) ^ (inputs[20]));
    assign layer0_outputs[3748] = ~(inputs[32]) | (inputs[52]);
    assign layer0_outputs[3749] = (inputs[206]) ^ (inputs[185]);
    assign layer0_outputs[3750] = inputs[104];
    assign layer0_outputs[3751] = 1'b0;
    assign layer0_outputs[3752] = inputs[72];
    assign layer0_outputs[3753] = (inputs[4]) | (inputs[157]);
    assign layer0_outputs[3754] = ~((inputs[146]) & (inputs[112]));
    assign layer0_outputs[3755] = 1'b1;
    assign layer0_outputs[3756] = ~(inputs[157]);
    assign layer0_outputs[3757] = 1'b1;
    assign layer0_outputs[3758] = (inputs[246]) & ~(inputs[56]);
    assign layer0_outputs[3759] = ~((inputs[241]) & (inputs[110]));
    assign layer0_outputs[3760] = ~((inputs[95]) & (inputs[71]));
    assign layer0_outputs[3761] = inputs[209];
    assign layer0_outputs[3762] = ~((inputs[147]) | (inputs[146]));
    assign layer0_outputs[3763] = ~(inputs[35]) | (inputs[50]);
    assign layer0_outputs[3764] = (inputs[213]) ^ (inputs[114]);
    assign layer0_outputs[3765] = ~((inputs[197]) & (inputs[102]));
    assign layer0_outputs[3766] = (inputs[58]) ^ (inputs[16]);
    assign layer0_outputs[3767] = inputs[80];
    assign layer0_outputs[3768] = (inputs[26]) | (inputs[108]);
    assign layer0_outputs[3769] = (inputs[24]) & ~(inputs[205]);
    assign layer0_outputs[3770] = 1'b1;
    assign layer0_outputs[3771] = ~(inputs[100]);
    assign layer0_outputs[3772] = ~(inputs[246]);
    assign layer0_outputs[3773] = 1'b1;
    assign layer0_outputs[3774] = ~(inputs[212]) | (inputs[220]);
    assign layer0_outputs[3775] = ~(inputs[63]) | (inputs[61]);
    assign layer0_outputs[3776] = ~(inputs[141]) | (inputs[171]);
    assign layer0_outputs[3777] = ~(inputs[209]) | (inputs[205]);
    assign layer0_outputs[3778] = ~(inputs[11]);
    assign layer0_outputs[3779] = ~(inputs[203]);
    assign layer0_outputs[3780] = inputs[238];
    assign layer0_outputs[3781] = ~(inputs[248]) | (inputs[127]);
    assign layer0_outputs[3782] = (inputs[22]) & (inputs[124]);
    assign layer0_outputs[3783] = ~(inputs[245]) | (inputs[145]);
    assign layer0_outputs[3784] = 1'b0;
    assign layer0_outputs[3785] = (inputs[229]) & ~(inputs[93]);
    assign layer0_outputs[3786] = ~(inputs[184]) | (inputs[130]);
    assign layer0_outputs[3787] = inputs[47];
    assign layer0_outputs[3788] = ~((inputs[97]) | (inputs[124]));
    assign layer0_outputs[3789] = ~(inputs[36]) | (inputs[28]);
    assign layer0_outputs[3790] = ~((inputs[225]) | (inputs[61]));
    assign layer0_outputs[3791] = inputs[107];
    assign layer0_outputs[3792] = (inputs[101]) & (inputs[188]);
    assign layer0_outputs[3793] = (inputs[210]) & (inputs[100]);
    assign layer0_outputs[3794] = ~(inputs[117]) | (inputs[210]);
    assign layer0_outputs[3795] = ~((inputs[178]) & (inputs[148]));
    assign layer0_outputs[3796] = (inputs[138]) & ~(inputs[94]);
    assign layer0_outputs[3797] = inputs[176];
    assign layer0_outputs[3798] = ~(inputs[33]) | (inputs[54]);
    assign layer0_outputs[3799] = inputs[248];
    assign layer0_outputs[3800] = ~(inputs[194]) | (inputs[28]);
    assign layer0_outputs[3801] = ~((inputs[114]) ^ (inputs[206]));
    assign layer0_outputs[3802] = (inputs[164]) & ~(inputs[112]);
    assign layer0_outputs[3803] = ~(inputs[161]);
    assign layer0_outputs[3804] = ~(inputs[201]) | (inputs[16]);
    assign layer0_outputs[3805] = (inputs[176]) | (inputs[236]);
    assign layer0_outputs[3806] = ~(inputs[168]);
    assign layer0_outputs[3807] = (inputs[23]) & ~(inputs[243]);
    assign layer0_outputs[3808] = 1'b1;
    assign layer0_outputs[3809] = ~((inputs[114]) ^ (inputs[8]));
    assign layer0_outputs[3810] = ~(inputs[238]);
    assign layer0_outputs[3811] = ~(inputs[229]) | (inputs[154]);
    assign layer0_outputs[3812] = ~(inputs[91]);
    assign layer0_outputs[3813] = ~((inputs[237]) & (inputs[226]));
    assign layer0_outputs[3814] = ~(inputs[60]) | (inputs[151]);
    assign layer0_outputs[3815] = 1'b0;
    assign layer0_outputs[3816] = ~((inputs[26]) ^ (inputs[132]));
    assign layer0_outputs[3817] = (inputs[43]) | (inputs[254]);
    assign layer0_outputs[3818] = 1'b0;
    assign layer0_outputs[3819] = ~(inputs[80]);
    assign layer0_outputs[3820] = ~(inputs[15]) | (inputs[158]);
    assign layer0_outputs[3821] = ~((inputs[234]) | (inputs[96]));
    assign layer0_outputs[3822] = (inputs[11]) ^ (inputs[226]);
    assign layer0_outputs[3823] = ~((inputs[199]) & (inputs[150]));
    assign layer0_outputs[3824] = ~(inputs[65]);
    assign layer0_outputs[3825] = (inputs[247]) | (inputs[183]);
    assign layer0_outputs[3826] = ~((inputs[247]) | (inputs[127]));
    assign layer0_outputs[3827] = ~(inputs[255]);
    assign layer0_outputs[3828] = ~(inputs[128]) | (inputs[139]);
    assign layer0_outputs[3829] = (inputs[155]) & ~(inputs[241]);
    assign layer0_outputs[3830] = (inputs[136]) | (inputs[52]);
    assign layer0_outputs[3831] = ~((inputs[96]) | (inputs[22]));
    assign layer0_outputs[3832] = 1'b0;
    assign layer0_outputs[3833] = 1'b1;
    assign layer0_outputs[3834] = ~(inputs[245]) | (inputs[154]);
    assign layer0_outputs[3835] = ~((inputs[192]) & (inputs[59]));
    assign layer0_outputs[3836] = ~(inputs[220]) | (inputs[149]);
    assign layer0_outputs[3837] = (inputs[38]) & (inputs[190]);
    assign layer0_outputs[3838] = (inputs[190]) | (inputs[88]);
    assign layer0_outputs[3839] = (inputs[239]) | (inputs[61]);
    assign layer0_outputs[3840] = ~(inputs[7]);
    assign layer0_outputs[3841] = ~(inputs[120]);
    assign layer0_outputs[3842] = ~((inputs[227]) | (inputs[182]));
    assign layer0_outputs[3843] = ~((inputs[234]) & (inputs[141]));
    assign layer0_outputs[3844] = (inputs[104]) & ~(inputs[159]);
    assign layer0_outputs[3845] = (inputs[2]) & ~(inputs[185]);
    assign layer0_outputs[3846] = ~((inputs[165]) | (inputs[230]));
    assign layer0_outputs[3847] = 1'b1;
    assign layer0_outputs[3848] = ~(inputs[157]);
    assign layer0_outputs[3849] = (inputs[147]) | (inputs[176]);
    assign layer0_outputs[3850] = (inputs[36]) & ~(inputs[233]);
    assign layer0_outputs[3851] = ~(inputs[215]);
    assign layer0_outputs[3852] = (inputs[216]) & ~(inputs[42]);
    assign layer0_outputs[3853] = 1'b0;
    assign layer0_outputs[3854] = ~(inputs[136]);
    assign layer0_outputs[3855] = ~((inputs[107]) | (inputs[81]));
    assign layer0_outputs[3856] = ~(inputs[30]) | (inputs[156]);
    assign layer0_outputs[3857] = ~((inputs[173]) ^ (inputs[1]));
    assign layer0_outputs[3858] = 1'b0;
    assign layer0_outputs[3859] = inputs[114];
    assign layer0_outputs[3860] = ~(inputs[144]) | (inputs[84]);
    assign layer0_outputs[3861] = inputs[233];
    assign layer0_outputs[3862] = inputs[123];
    assign layer0_outputs[3863] = (inputs[92]) & ~(inputs[63]);
    assign layer0_outputs[3864] = (inputs[210]) & ~(inputs[109]);
    assign layer0_outputs[3865] = 1'b0;
    assign layer0_outputs[3866] = ~(inputs[99]);
    assign layer0_outputs[3867] = ~(inputs[23]);
    assign layer0_outputs[3868] = ~(inputs[118]) | (inputs[73]);
    assign layer0_outputs[3869] = 1'b0;
    assign layer0_outputs[3870] = 1'b1;
    assign layer0_outputs[3871] = (inputs[6]) ^ (inputs[192]);
    assign layer0_outputs[3872] = inputs[157];
    assign layer0_outputs[3873] = ~(inputs[18]);
    assign layer0_outputs[3874] = (inputs[4]) & ~(inputs[91]);
    assign layer0_outputs[3875] = 1'b1;
    assign layer0_outputs[3876] = ~(inputs[18]);
    assign layer0_outputs[3877] = 1'b0;
    assign layer0_outputs[3878] = ~(inputs[28]) | (inputs[109]);
    assign layer0_outputs[3879] = (inputs[132]) & (inputs[124]);
    assign layer0_outputs[3880] = inputs[122];
    assign layer0_outputs[3881] = ~((inputs[33]) & (inputs[218]));
    assign layer0_outputs[3882] = (inputs[1]) | (inputs[254]);
    assign layer0_outputs[3883] = ~(inputs[70]) | (inputs[17]);
    assign layer0_outputs[3884] = 1'b1;
    assign layer0_outputs[3885] = 1'b1;
    assign layer0_outputs[3886] = (inputs[33]) | (inputs[120]);
    assign layer0_outputs[3887] = 1'b0;
    assign layer0_outputs[3888] = ~(inputs[250]) | (inputs[76]);
    assign layer0_outputs[3889] = ~(inputs[236]);
    assign layer0_outputs[3890] = (inputs[196]) & ~(inputs[27]);
    assign layer0_outputs[3891] = (inputs[99]) | (inputs[100]);
    assign layer0_outputs[3892] = 1'b1;
    assign layer0_outputs[3893] = ~((inputs[241]) | (inputs[117]));
    assign layer0_outputs[3894] = (inputs[65]) & ~(inputs[49]);
    assign layer0_outputs[3895] = ~(inputs[219]) | (inputs[217]);
    assign layer0_outputs[3896] = ~(inputs[254]);
    assign layer0_outputs[3897] = 1'b0;
    assign layer0_outputs[3898] = ~((inputs[177]) ^ (inputs[226]));
    assign layer0_outputs[3899] = ~(inputs[27]) | (inputs[89]);
    assign layer0_outputs[3900] = ~((inputs[144]) | (inputs[118]));
    assign layer0_outputs[3901] = inputs[119];
    assign layer0_outputs[3902] = 1'b1;
    assign layer0_outputs[3903] = ~(inputs[27]) | (inputs[56]);
    assign layer0_outputs[3904] = ~(inputs[167]) | (inputs[50]);
    assign layer0_outputs[3905] = (inputs[41]) ^ (inputs[72]);
    assign layer0_outputs[3906] = ~(inputs[85]) | (inputs[171]);
    assign layer0_outputs[3907] = ~(inputs[197]);
    assign layer0_outputs[3908] = inputs[230];
    assign layer0_outputs[3909] = inputs[95];
    assign layer0_outputs[3910] = ~(inputs[3]) | (inputs[87]);
    assign layer0_outputs[3911] = 1'b0;
    assign layer0_outputs[3912] = ~((inputs[41]) & (inputs[214]));
    assign layer0_outputs[3913] = ~(inputs[182]);
    assign layer0_outputs[3914] = (inputs[89]) & ~(inputs[31]);
    assign layer0_outputs[3915] = ~(inputs[193]);
    assign layer0_outputs[3916] = 1'b0;
    assign layer0_outputs[3917] = ~((inputs[91]) ^ (inputs[78]));
    assign layer0_outputs[3918] = (inputs[71]) & (inputs[3]);
    assign layer0_outputs[3919] = (inputs[229]) | (inputs[179]);
    assign layer0_outputs[3920] = ~((inputs[64]) | (inputs[147]));
    assign layer0_outputs[3921] = ~(inputs[130]);
    assign layer0_outputs[3922] = ~((inputs[97]) & (inputs[181]));
    assign layer0_outputs[3923] = (inputs[93]) | (inputs[83]);
    assign layer0_outputs[3924] = inputs[208];
    assign layer0_outputs[3925] = ~(inputs[168]) | (inputs[76]);
    assign layer0_outputs[3926] = (inputs[183]) | (inputs[115]);
    assign layer0_outputs[3927] = (inputs[78]) & ~(inputs[46]);
    assign layer0_outputs[3928] = ~(inputs[104]) | (inputs[57]);
    assign layer0_outputs[3929] = ~((inputs[161]) ^ (inputs[132]));
    assign layer0_outputs[3930] = ~((inputs[224]) & (inputs[234]));
    assign layer0_outputs[3931] = ~((inputs[143]) | (inputs[99]));
    assign layer0_outputs[3932] = ~((inputs[195]) & (inputs[39]));
    assign layer0_outputs[3933] = inputs[225];
    assign layer0_outputs[3934] = (inputs[52]) & ~(inputs[160]);
    assign layer0_outputs[3935] = ~((inputs[101]) | (inputs[76]));
    assign layer0_outputs[3936] = ~(inputs[70]) | (inputs[24]);
    assign layer0_outputs[3937] = (inputs[160]) & (inputs[35]);
    assign layer0_outputs[3938] = inputs[113];
    assign layer0_outputs[3939] = ~(inputs[107]);
    assign layer0_outputs[3940] = inputs[216];
    assign layer0_outputs[3941] = ~((inputs[205]) | (inputs[115]));
    assign layer0_outputs[3942] = (inputs[202]) | (inputs[83]);
    assign layer0_outputs[3943] = ~(inputs[9]) | (inputs[214]);
    assign layer0_outputs[3944] = (inputs[254]) & ~(inputs[97]);
    assign layer0_outputs[3945] = inputs[215];
    assign layer0_outputs[3946] = (inputs[47]) | (inputs[225]);
    assign layer0_outputs[3947] = (inputs[26]) | (inputs[245]);
    assign layer0_outputs[3948] = ~((inputs[8]) ^ (inputs[179]));
    assign layer0_outputs[3949] = (inputs[191]) & ~(inputs[22]);
    assign layer0_outputs[3950] = (inputs[10]) & ~(inputs[234]);
    assign layer0_outputs[3951] = 1'b0;
    assign layer0_outputs[3952] = ~(inputs[26]) | (inputs[90]);
    assign layer0_outputs[3953] = ~(inputs[77]) | (inputs[170]);
    assign layer0_outputs[3954] = ~(inputs[226]);
    assign layer0_outputs[3955] = (inputs[52]) & ~(inputs[174]);
    assign layer0_outputs[3956] = (inputs[247]) ^ (inputs[75]);
    assign layer0_outputs[3957] = (inputs[57]) & ~(inputs[187]);
    assign layer0_outputs[3958] = 1'b0;
    assign layer0_outputs[3959] = ~(inputs[231]) | (inputs[138]);
    assign layer0_outputs[3960] = inputs[250];
    assign layer0_outputs[3961] = ~((inputs[244]) & (inputs[141]));
    assign layer0_outputs[3962] = ~((inputs[112]) ^ (inputs[70]));
    assign layer0_outputs[3963] = ~(inputs[210]) | (inputs[47]);
    assign layer0_outputs[3964] = ~((inputs[241]) | (inputs[178]));
    assign layer0_outputs[3965] = ~(inputs[25]) | (inputs[44]);
    assign layer0_outputs[3966] = (inputs[251]) & (inputs[212]);
    assign layer0_outputs[3967] = ~((inputs[163]) ^ (inputs[18]));
    assign layer0_outputs[3968] = 1'b0;
    assign layer0_outputs[3969] = ~((inputs[53]) ^ (inputs[241]));
    assign layer0_outputs[3970] = ~((inputs[242]) | (inputs[130]));
    assign layer0_outputs[3971] = ~(inputs[96]) | (inputs[144]);
    assign layer0_outputs[3972] = ~((inputs[38]) ^ (inputs[12]));
    assign layer0_outputs[3973] = ~((inputs[78]) ^ (inputs[157]));
    assign layer0_outputs[3974] = ~(inputs[244]);
    assign layer0_outputs[3975] = inputs[31];
    assign layer0_outputs[3976] = (inputs[182]) & ~(inputs[76]);
    assign layer0_outputs[3977] = inputs[171];
    assign layer0_outputs[3978] = (inputs[117]) | (inputs[140]);
    assign layer0_outputs[3979] = 1'b1;
    assign layer0_outputs[3980] = (inputs[157]) & ~(inputs[0]);
    assign layer0_outputs[3981] = ~(inputs[176]) | (inputs[153]);
    assign layer0_outputs[3982] = 1'b1;
    assign layer0_outputs[3983] = ~(inputs[203]) | (inputs[61]);
    assign layer0_outputs[3984] = (inputs[30]) & (inputs[225]);
    assign layer0_outputs[3985] = ~((inputs[187]) | (inputs[75]));
    assign layer0_outputs[3986] = ~(inputs[188]);
    assign layer0_outputs[3987] = ~(inputs[86]);
    assign layer0_outputs[3988] = inputs[174];
    assign layer0_outputs[3989] = ~((inputs[214]) | (inputs[68]));
    assign layer0_outputs[3990] = (inputs[168]) & (inputs[87]);
    assign layer0_outputs[3991] = ~(inputs[182]);
    assign layer0_outputs[3992] = (inputs[12]) & ~(inputs[238]);
    assign layer0_outputs[3993] = ~(inputs[247]) | (inputs[59]);
    assign layer0_outputs[3994] = (inputs[21]) & ~(inputs[80]);
    assign layer0_outputs[3995] = ~((inputs[253]) ^ (inputs[98]));
    assign layer0_outputs[3996] = inputs[206];
    assign layer0_outputs[3997] = inputs[27];
    assign layer0_outputs[3998] = ~(inputs[119]);
    assign layer0_outputs[3999] = (inputs[167]) & ~(inputs[229]);
    assign layer0_outputs[4000] = ~((inputs[139]) ^ (inputs[240]));
    assign layer0_outputs[4001] = ~((inputs[107]) ^ (inputs[142]));
    assign layer0_outputs[4002] = ~(inputs[72]);
    assign layer0_outputs[4003] = (inputs[74]) & ~(inputs[151]);
    assign layer0_outputs[4004] = 1'b1;
    assign layer0_outputs[4005] = 1'b1;
    assign layer0_outputs[4006] = (inputs[158]) & ~(inputs[113]);
    assign layer0_outputs[4007] = (inputs[7]) & ~(inputs[66]);
    assign layer0_outputs[4008] = (inputs[189]) ^ (inputs[51]);
    assign layer0_outputs[4009] = inputs[175];
    assign layer0_outputs[4010] = 1'b1;
    assign layer0_outputs[4011] = ~((inputs[69]) | (inputs[153]));
    assign layer0_outputs[4012] = ~(inputs[223]) | (inputs[124]);
    assign layer0_outputs[4013] = 1'b1;
    assign layer0_outputs[4014] = (inputs[77]) & ~(inputs[12]);
    assign layer0_outputs[4015] = (inputs[70]) ^ (inputs[158]);
    assign layer0_outputs[4016] = ~((inputs[95]) ^ (inputs[244]));
    assign layer0_outputs[4017] = ~(inputs[134]) | (inputs[37]);
    assign layer0_outputs[4018] = inputs[199];
    assign layer0_outputs[4019] = ~(inputs[189]) | (inputs[13]);
    assign layer0_outputs[4020] = (inputs[159]) & ~(inputs[251]);
    assign layer0_outputs[4021] = (inputs[149]) & ~(inputs[187]);
    assign layer0_outputs[4022] = ~(inputs[65]);
    assign layer0_outputs[4023] = inputs[45];
    assign layer0_outputs[4024] = (inputs[118]) & ~(inputs[240]);
    assign layer0_outputs[4025] = inputs[108];
    assign layer0_outputs[4026] = (inputs[163]) & (inputs[98]);
    assign layer0_outputs[4027] = 1'b1;
    assign layer0_outputs[4028] = ~(inputs[2]);
    assign layer0_outputs[4029] = inputs[199];
    assign layer0_outputs[4030] = (inputs[174]) & (inputs[126]);
    assign layer0_outputs[4031] = (inputs[231]) & ~(inputs[187]);
    assign layer0_outputs[4032] = ~(inputs[210]);
    assign layer0_outputs[4033] = 1'b1;
    assign layer0_outputs[4034] = (inputs[43]) ^ (inputs[93]);
    assign layer0_outputs[4035] = 1'b1;
    assign layer0_outputs[4036] = ~(inputs[136]) | (inputs[91]);
    assign layer0_outputs[4037] = inputs[129];
    assign layer0_outputs[4038] = (inputs[142]) & ~(inputs[33]);
    assign layer0_outputs[4039] = ~((inputs[91]) & (inputs[146]));
    assign layer0_outputs[4040] = inputs[141];
    assign layer0_outputs[4041] = ~(inputs[69]) | (inputs[56]);
    assign layer0_outputs[4042] = ~((inputs[14]) & (inputs[190]));
    assign layer0_outputs[4043] = (inputs[252]) & (inputs[179]);
    assign layer0_outputs[4044] = ~(inputs[232]);
    assign layer0_outputs[4045] = (inputs[45]) & (inputs[21]);
    assign layer0_outputs[4046] = (inputs[171]) & ~(inputs[84]);
    assign layer0_outputs[4047] = ~(inputs[251]);
    assign layer0_outputs[4048] = ~(inputs[142]);
    assign layer0_outputs[4049] = ~(inputs[143]) | (inputs[43]);
    assign layer0_outputs[4050] = inputs[14];
    assign layer0_outputs[4051] = (inputs[210]) & ~(inputs[159]);
    assign layer0_outputs[4052] = (inputs[66]) & (inputs[57]);
    assign layer0_outputs[4053] = (inputs[9]) & (inputs[95]);
    assign layer0_outputs[4054] = (inputs[147]) & ~(inputs[11]);
    assign layer0_outputs[4055] = ~(inputs[14]) | (inputs[222]);
    assign layer0_outputs[4056] = (inputs[29]) ^ (inputs[61]);
    assign layer0_outputs[4057] = ~(inputs[231]) | (inputs[55]);
    assign layer0_outputs[4058] = (inputs[228]) & ~(inputs[23]);
    assign layer0_outputs[4059] = 1'b1;
    assign layer0_outputs[4060] = ~((inputs[27]) ^ (inputs[216]));
    assign layer0_outputs[4061] = 1'b1;
    assign layer0_outputs[4062] = (inputs[245]) & (inputs[113]);
    assign layer0_outputs[4063] = ~((inputs[201]) | (inputs[60]));
    assign layer0_outputs[4064] = ~((inputs[199]) & (inputs[168]));
    assign layer0_outputs[4065] = ~(inputs[28]);
    assign layer0_outputs[4066] = (inputs[41]) | (inputs[163]);
    assign layer0_outputs[4067] = ~(inputs[11]);
    assign layer0_outputs[4068] = 1'b0;
    assign layer0_outputs[4069] = (inputs[1]) ^ (inputs[33]);
    assign layer0_outputs[4070] = inputs[46];
    assign layer0_outputs[4071] = 1'b0;
    assign layer0_outputs[4072] = ~(inputs[181]) | (inputs[212]);
    assign layer0_outputs[4073] = ~(inputs[147]);
    assign layer0_outputs[4074] = (inputs[114]) ^ (inputs[158]);
    assign layer0_outputs[4075] = ~(inputs[72]) | (inputs[50]);
    assign layer0_outputs[4076] = (inputs[63]) & ~(inputs[23]);
    assign layer0_outputs[4077] = inputs[2];
    assign layer0_outputs[4078] = ~(inputs[217]) | (inputs[255]);
    assign layer0_outputs[4079] = (inputs[192]) | (inputs[54]);
    assign layer0_outputs[4080] = ~(inputs[39]) | (inputs[174]);
    assign layer0_outputs[4081] = ~((inputs[3]) ^ (inputs[15]));
    assign layer0_outputs[4082] = ~((inputs[75]) | (inputs[204]));
    assign layer0_outputs[4083] = 1'b1;
    assign layer0_outputs[4084] = ~((inputs[198]) | (inputs[244]));
    assign layer0_outputs[4085] = ~(inputs[144]);
    assign layer0_outputs[4086] = ~(inputs[16]) | (inputs[11]);
    assign layer0_outputs[4087] = (inputs[21]) & (inputs[27]);
    assign layer0_outputs[4088] = ~((inputs[197]) ^ (inputs[77]));
    assign layer0_outputs[4089] = 1'b1;
    assign layer0_outputs[4090] = ~(inputs[56]);
    assign layer0_outputs[4091] = ~(inputs[253]);
    assign layer0_outputs[4092] = (inputs[43]) ^ (inputs[79]);
    assign layer0_outputs[4093] = inputs[122];
    assign layer0_outputs[4094] = 1'b1;
    assign layer0_outputs[4095] = (inputs[186]) & ~(inputs[84]);
    assign layer0_outputs[4096] = ~((inputs[231]) | (inputs[66]));
    assign layer0_outputs[4097] = 1'b0;
    assign layer0_outputs[4098] = ~((inputs[180]) ^ (inputs[191]));
    assign layer0_outputs[4099] = (inputs[79]) & ~(inputs[187]);
    assign layer0_outputs[4100] = ~((inputs[114]) & (inputs[31]));
    assign layer0_outputs[4101] = (inputs[92]) ^ (inputs[153]);
    assign layer0_outputs[4102] = 1'b1;
    assign layer0_outputs[4103] = ~((inputs[218]) ^ (inputs[159]));
    assign layer0_outputs[4104] = 1'b1;
    assign layer0_outputs[4105] = 1'b0;
    assign layer0_outputs[4106] = ~(inputs[45]);
    assign layer0_outputs[4107] = ~(inputs[247]) | (inputs[253]);
    assign layer0_outputs[4108] = inputs[237];
    assign layer0_outputs[4109] = (inputs[254]) & ~(inputs[144]);
    assign layer0_outputs[4110] = 1'b0;
    assign layer0_outputs[4111] = ~(inputs[91]);
    assign layer0_outputs[4112] = (inputs[192]) & ~(inputs[198]);
    assign layer0_outputs[4113] = ~(inputs[21]) | (inputs[255]);
    assign layer0_outputs[4114] = (inputs[66]) & ~(inputs[97]);
    assign layer0_outputs[4115] = ~(inputs[62]) | (inputs[29]);
    assign layer0_outputs[4116] = ~(inputs[87]) | (inputs[151]);
    assign layer0_outputs[4117] = (inputs[75]) | (inputs[242]);
    assign layer0_outputs[4118] = ~(inputs[131]);
    assign layer0_outputs[4119] = ~(inputs[57]);
    assign layer0_outputs[4120] = (inputs[51]) & ~(inputs[227]);
    assign layer0_outputs[4121] = inputs[167];
    assign layer0_outputs[4122] = (inputs[56]) & ~(inputs[230]);
    assign layer0_outputs[4123] = ~((inputs[251]) | (inputs[167]));
    assign layer0_outputs[4124] = (inputs[99]) & (inputs[184]);
    assign layer0_outputs[4125] = (inputs[157]) & (inputs[219]);
    assign layer0_outputs[4126] = inputs[97];
    assign layer0_outputs[4127] = (inputs[215]) ^ (inputs[253]);
    assign layer0_outputs[4128] = 1'b1;
    assign layer0_outputs[4129] = ~(inputs[118]);
    assign layer0_outputs[4130] = (inputs[14]) & (inputs[246]);
    assign layer0_outputs[4131] = (inputs[248]) & (inputs[124]);
    assign layer0_outputs[4132] = ~(inputs[96]) | (inputs[93]);
    assign layer0_outputs[4133] = inputs[117];
    assign layer0_outputs[4134] = ~(inputs[254]);
    assign layer0_outputs[4135] = 1'b0;
    assign layer0_outputs[4136] = 1'b1;
    assign layer0_outputs[4137] = ~((inputs[224]) & (inputs[253]));
    assign layer0_outputs[4138] = (inputs[137]) | (inputs[27]);
    assign layer0_outputs[4139] = ~(inputs[26]) | (inputs[155]);
    assign layer0_outputs[4140] = ~(inputs[180]);
    assign layer0_outputs[4141] = (inputs[236]) & ~(inputs[29]);
    assign layer0_outputs[4142] = 1'b1;
    assign layer0_outputs[4143] = ~((inputs[170]) & (inputs[44]));
    assign layer0_outputs[4144] = 1'b0;
    assign layer0_outputs[4145] = (inputs[195]) ^ (inputs[129]);
    assign layer0_outputs[4146] = ~(inputs[244]);
    assign layer0_outputs[4147] = inputs[16];
    assign layer0_outputs[4148] = 1'b0;
    assign layer0_outputs[4149] = (inputs[67]) & (inputs[10]);
    assign layer0_outputs[4150] = ~(inputs[149]) | (inputs[236]);
    assign layer0_outputs[4151] = inputs[236];
    assign layer0_outputs[4152] = (inputs[209]) & ~(inputs[128]);
    assign layer0_outputs[4153] = ~((inputs[7]) | (inputs[102]));
    assign layer0_outputs[4154] = ~((inputs[30]) & (inputs[44]));
    assign layer0_outputs[4155] = ~(inputs[149]);
    assign layer0_outputs[4156] = ~(inputs[230]);
    assign layer0_outputs[4157] = ~(inputs[243]);
    assign layer0_outputs[4158] = (inputs[183]) & (inputs[110]);
    assign layer0_outputs[4159] = inputs[150];
    assign layer0_outputs[4160] = ~((inputs[142]) | (inputs[151]));
    assign layer0_outputs[4161] = 1'b0;
    assign layer0_outputs[4162] = ~(inputs[104]) | (inputs[36]);
    assign layer0_outputs[4163] = (inputs[49]) | (inputs[236]);
    assign layer0_outputs[4164] = (inputs[159]) & (inputs[112]);
    assign layer0_outputs[4165] = (inputs[230]) & ~(inputs[188]);
    assign layer0_outputs[4166] = 1'b0;
    assign layer0_outputs[4167] = ~(inputs[102]);
    assign layer0_outputs[4168] = ~(inputs[174]);
    assign layer0_outputs[4169] = ~(inputs[58]);
    assign layer0_outputs[4170] = 1'b1;
    assign layer0_outputs[4171] = ~(inputs[83]) | (inputs[2]);
    assign layer0_outputs[4172] = ~(inputs[35]);
    assign layer0_outputs[4173] = (inputs[235]) & ~(inputs[135]);
    assign layer0_outputs[4174] = 1'b1;
    assign layer0_outputs[4175] = 1'b0;
    assign layer0_outputs[4176] = ~((inputs[80]) ^ (inputs[48]));
    assign layer0_outputs[4177] = ~(inputs[174]) | (inputs[70]);
    assign layer0_outputs[4178] = inputs[179];
    assign layer0_outputs[4179] = (inputs[192]) & (inputs[150]);
    assign layer0_outputs[4180] = inputs[27];
    assign layer0_outputs[4181] = inputs[161];
    assign layer0_outputs[4182] = (inputs[252]) & ~(inputs[151]);
    assign layer0_outputs[4183] = (inputs[82]) & ~(inputs[141]);
    assign layer0_outputs[4184] = ~((inputs[185]) & (inputs[237]));
    assign layer0_outputs[4185] = ~(inputs[240]) | (inputs[216]);
    assign layer0_outputs[4186] = ~(inputs[110]);
    assign layer0_outputs[4187] = inputs[250];
    assign layer0_outputs[4188] = 1'b0;
    assign layer0_outputs[4189] = ~(inputs[150]) | (inputs[66]);
    assign layer0_outputs[4190] = ~((inputs[182]) ^ (inputs[211]));
    assign layer0_outputs[4191] = 1'b0;
    assign layer0_outputs[4192] = inputs[214];
    assign layer0_outputs[4193] = ~(inputs[175]);
    assign layer0_outputs[4194] = ~(inputs[131]) | (inputs[39]);
    assign layer0_outputs[4195] = ~(inputs[146]);
    assign layer0_outputs[4196] = 1'b0;
    assign layer0_outputs[4197] = 1'b1;
    assign layer0_outputs[4198] = inputs[120];
    assign layer0_outputs[4199] = (inputs[165]) ^ (inputs[18]);
    assign layer0_outputs[4200] = ~(inputs[97]);
    assign layer0_outputs[4201] = ~(inputs[254]);
    assign layer0_outputs[4202] = ~(inputs[234]) | (inputs[206]);
    assign layer0_outputs[4203] = ~((inputs[199]) & (inputs[221]));
    assign layer0_outputs[4204] = inputs[231];
    assign layer0_outputs[4205] = ~(inputs[243]) | (inputs[242]);
    assign layer0_outputs[4206] = ~((inputs[138]) ^ (inputs[161]));
    assign layer0_outputs[4207] = ~(inputs[205]);
    assign layer0_outputs[4208] = ~((inputs[138]) | (inputs[52]));
    assign layer0_outputs[4209] = ~((inputs[45]) ^ (inputs[177]));
    assign layer0_outputs[4210] = ~((inputs[70]) | (inputs[16]));
    assign layer0_outputs[4211] = inputs[190];
    assign layer0_outputs[4212] = (inputs[96]) & ~(inputs[60]);
    assign layer0_outputs[4213] = (inputs[127]) ^ (inputs[55]);
    assign layer0_outputs[4214] = ~((inputs[82]) | (inputs[209]));
    assign layer0_outputs[4215] = (inputs[60]) | (inputs[230]);
    assign layer0_outputs[4216] = ~(inputs[17]) | (inputs[151]);
    assign layer0_outputs[4217] = (inputs[239]) & ~(inputs[112]);
    assign layer0_outputs[4218] = (inputs[97]) & ~(inputs[144]);
    assign layer0_outputs[4219] = ~(inputs[165]) | (inputs[28]);
    assign layer0_outputs[4220] = (inputs[98]) & (inputs[97]);
    assign layer0_outputs[4221] = inputs[148];
    assign layer0_outputs[4222] = inputs[13];
    assign layer0_outputs[4223] = 1'b0;
    assign layer0_outputs[4224] = 1'b1;
    assign layer0_outputs[4225] = ~(inputs[89]) | (inputs[97]);
    assign layer0_outputs[4226] = ~(inputs[123]) | (inputs[183]);
    assign layer0_outputs[4227] = ~((inputs[251]) ^ (inputs[220]));
    assign layer0_outputs[4228] = (inputs[121]) & (inputs[179]);
    assign layer0_outputs[4229] = 1'b0;
    assign layer0_outputs[4230] = ~(inputs[230]);
    assign layer0_outputs[4231] = inputs[103];
    assign layer0_outputs[4232] = inputs[117];
    assign layer0_outputs[4233] = (inputs[189]) ^ (inputs[21]);
    assign layer0_outputs[4234] = ~(inputs[212]) | (inputs[217]);
    assign layer0_outputs[4235] = ~((inputs[31]) ^ (inputs[236]));
    assign layer0_outputs[4236] = ~(inputs[43]) | (inputs[176]);
    assign layer0_outputs[4237] = ~((inputs[152]) | (inputs[28]));
    assign layer0_outputs[4238] = ~((inputs[124]) | (inputs[165]));
    assign layer0_outputs[4239] = 1'b0;
    assign layer0_outputs[4240] = ~((inputs[245]) & (inputs[16]));
    assign layer0_outputs[4241] = 1'b0;
    assign layer0_outputs[4242] = ~((inputs[3]) | (inputs[150]));
    assign layer0_outputs[4243] = inputs[245];
    assign layer0_outputs[4244] = ~(inputs[59]);
    assign layer0_outputs[4245] = (inputs[69]) | (inputs[197]);
    assign layer0_outputs[4246] = (inputs[163]) & ~(inputs[230]);
    assign layer0_outputs[4247] = ~(inputs[55]);
    assign layer0_outputs[4248] = ~((inputs[165]) | (inputs[20]));
    assign layer0_outputs[4249] = ~(inputs[22]) | (inputs[23]);
    assign layer0_outputs[4250] = ~(inputs[114]) | (inputs[200]);
    assign layer0_outputs[4251] = (inputs[67]) ^ (inputs[14]);
    assign layer0_outputs[4252] = ~((inputs[72]) | (inputs[9]));
    assign layer0_outputs[4253] = (inputs[148]) | (inputs[13]);
    assign layer0_outputs[4254] = (inputs[101]) | (inputs[12]);
    assign layer0_outputs[4255] = 1'b1;
    assign layer0_outputs[4256] = 1'b1;
    assign layer0_outputs[4257] = inputs[202];
    assign layer0_outputs[4258] = (inputs[201]) & ~(inputs[194]);
    assign layer0_outputs[4259] = ~((inputs[137]) | (inputs[26]));
    assign layer0_outputs[4260] = (inputs[148]) & ~(inputs[161]);
    assign layer0_outputs[4261] = (inputs[131]) ^ (inputs[223]);
    assign layer0_outputs[4262] = ~(inputs[140]);
    assign layer0_outputs[4263] = ~((inputs[224]) & (inputs[248]));
    assign layer0_outputs[4264] = ~((inputs[107]) & (inputs[114]));
    assign layer0_outputs[4265] = ~(inputs[144]);
    assign layer0_outputs[4266] = 1'b0;
    assign layer0_outputs[4267] = inputs[155];
    assign layer0_outputs[4268] = (inputs[28]) & ~(inputs[62]);
    assign layer0_outputs[4269] = (inputs[196]) | (inputs[44]);
    assign layer0_outputs[4270] = (inputs[213]) & ~(inputs[150]);
    assign layer0_outputs[4271] = ~((inputs[201]) | (inputs[119]));
    assign layer0_outputs[4272] = ~(inputs[77]) | (inputs[202]);
    assign layer0_outputs[4273] = ~((inputs[41]) ^ (inputs[63]));
    assign layer0_outputs[4274] = 1'b1;
    assign layer0_outputs[4275] = inputs[186];
    assign layer0_outputs[4276] = inputs[235];
    assign layer0_outputs[4277] = ~(inputs[170]);
    assign layer0_outputs[4278] = (inputs[186]) & ~(inputs[101]);
    assign layer0_outputs[4279] = (inputs[42]) ^ (inputs[173]);
    assign layer0_outputs[4280] = ~(inputs[106]);
    assign layer0_outputs[4281] = ~(inputs[148]) | (inputs[168]);
    assign layer0_outputs[4282] = inputs[235];
    assign layer0_outputs[4283] = 1'b0;
    assign layer0_outputs[4284] = ~((inputs[73]) & (inputs[22]));
    assign layer0_outputs[4285] = (inputs[153]) & ~(inputs[191]);
    assign layer0_outputs[4286] = ~((inputs[175]) & (inputs[3]));
    assign layer0_outputs[4287] = ~(inputs[179]) | (inputs[53]);
    assign layer0_outputs[4288] = ~(inputs[34]) | (inputs[59]);
    assign layer0_outputs[4289] = (inputs[117]) & ~(inputs[247]);
    assign layer0_outputs[4290] = (inputs[57]) ^ (inputs[175]);
    assign layer0_outputs[4291] = (inputs[29]) & ~(inputs[203]);
    assign layer0_outputs[4292] = 1'b0;
    assign layer0_outputs[4293] = ~(inputs[56]);
    assign layer0_outputs[4294] = (inputs[208]) | (inputs[11]);
    assign layer0_outputs[4295] = ~((inputs[98]) & (inputs[244]));
    assign layer0_outputs[4296] = ~(inputs[105]);
    assign layer0_outputs[4297] = (inputs[13]) | (inputs[15]);
    assign layer0_outputs[4298] = inputs[216];
    assign layer0_outputs[4299] = ~(inputs[16]);
    assign layer0_outputs[4300] = (inputs[51]) | (inputs[55]);
    assign layer0_outputs[4301] = ~((inputs[134]) | (inputs[130]));
    assign layer0_outputs[4302] = inputs[249];
    assign layer0_outputs[4303] = (inputs[182]) | (inputs[96]);
    assign layer0_outputs[4304] = ~((inputs[200]) & (inputs[135]));
    assign layer0_outputs[4305] = ~((inputs[232]) ^ (inputs[34]));
    assign layer0_outputs[4306] = ~(inputs[143]) | (inputs[226]);
    assign layer0_outputs[4307] = (inputs[34]) & (inputs[246]);
    assign layer0_outputs[4308] = (inputs[33]) & (inputs[26]);
    assign layer0_outputs[4309] = ~((inputs[131]) & (inputs[208]));
    assign layer0_outputs[4310] = inputs[18];
    assign layer0_outputs[4311] = 1'b0;
    assign layer0_outputs[4312] = ~(inputs[45]) | (inputs[148]);
    assign layer0_outputs[4313] = ~((inputs[160]) ^ (inputs[252]));
    assign layer0_outputs[4314] = inputs[241];
    assign layer0_outputs[4315] = ~(inputs[75]) | (inputs[201]);
    assign layer0_outputs[4316] = ~(inputs[49]);
    assign layer0_outputs[4317] = ~((inputs[104]) ^ (inputs[10]));
    assign layer0_outputs[4318] = (inputs[25]) & ~(inputs[30]);
    assign layer0_outputs[4319] = ~((inputs[83]) ^ (inputs[248]));
    assign layer0_outputs[4320] = 1'b1;
    assign layer0_outputs[4321] = 1'b0;
    assign layer0_outputs[4322] = inputs[5];
    assign layer0_outputs[4323] = ~(inputs[160]);
    assign layer0_outputs[4324] = (inputs[73]) | (inputs[250]);
    assign layer0_outputs[4325] = ~((inputs[139]) | (inputs[140]));
    assign layer0_outputs[4326] = ~(inputs[176]) | (inputs[130]);
    assign layer0_outputs[4327] = (inputs[234]) & (inputs[139]);
    assign layer0_outputs[4328] = inputs[140];
    assign layer0_outputs[4329] = (inputs[3]) & (inputs[220]);
    assign layer0_outputs[4330] = inputs[150];
    assign layer0_outputs[4331] = 1'b0;
    assign layer0_outputs[4332] = (inputs[9]) & ~(inputs[216]);
    assign layer0_outputs[4333] = ~(inputs[214]) | (inputs[206]);
    assign layer0_outputs[4334] = inputs[133];
    assign layer0_outputs[4335] = ~((inputs[208]) ^ (inputs[42]));
    assign layer0_outputs[4336] = 1'b0;
    assign layer0_outputs[4337] = (inputs[2]) & (inputs[65]);
    assign layer0_outputs[4338] = ~((inputs[145]) | (inputs[94]));
    assign layer0_outputs[4339] = ~(inputs[135]) | (inputs[146]);
    assign layer0_outputs[4340] = ~((inputs[112]) ^ (inputs[76]));
    assign layer0_outputs[4341] = (inputs[230]) & ~(inputs[37]);
    assign layer0_outputs[4342] = (inputs[17]) & (inputs[215]);
    assign layer0_outputs[4343] = (inputs[103]) & ~(inputs[97]);
    assign layer0_outputs[4344] = ~((inputs[74]) | (inputs[48]));
    assign layer0_outputs[4345] = inputs[53];
    assign layer0_outputs[4346] = ~(inputs[74]);
    assign layer0_outputs[4347] = ~((inputs[236]) ^ (inputs[58]));
    assign layer0_outputs[4348] = (inputs[151]) & ~(inputs[6]);
    assign layer0_outputs[4349] = (inputs[108]) | (inputs[171]);
    assign layer0_outputs[4350] = 1'b0;
    assign layer0_outputs[4351] = (inputs[11]) & ~(inputs[93]);
    assign layer0_outputs[4352] = (inputs[105]) & (inputs[183]);
    assign layer0_outputs[4353] = 1'b0;
    assign layer0_outputs[4354] = ~(inputs[183]) | (inputs[30]);
    assign layer0_outputs[4355] = (inputs[228]) & (inputs[200]);
    assign layer0_outputs[4356] = (inputs[175]) ^ (inputs[42]);
    assign layer0_outputs[4357] = ~(inputs[254]);
    assign layer0_outputs[4358] = ~(inputs[82]) | (inputs[139]);
    assign layer0_outputs[4359] = ~(inputs[77]);
    assign layer0_outputs[4360] = 1'b1;
    assign layer0_outputs[4361] = inputs[239];
    assign layer0_outputs[4362] = (inputs[188]) | (inputs[121]);
    assign layer0_outputs[4363] = (inputs[221]) & ~(inputs[22]);
    assign layer0_outputs[4364] = ~(inputs[179]) | (inputs[171]);
    assign layer0_outputs[4365] = (inputs[83]) & ~(inputs[141]);
    assign layer0_outputs[4366] = ~((inputs[132]) ^ (inputs[79]));
    assign layer0_outputs[4367] = inputs[167];
    assign layer0_outputs[4368] = (inputs[111]) & (inputs[234]);
    assign layer0_outputs[4369] = (inputs[12]) | (inputs[191]);
    assign layer0_outputs[4370] = (inputs[169]) & ~(inputs[240]);
    assign layer0_outputs[4371] = ~(inputs[148]) | (inputs[115]);
    assign layer0_outputs[4372] = (inputs[172]) & ~(inputs[136]);
    assign layer0_outputs[4373] = 1'b1;
    assign layer0_outputs[4374] = inputs[223];
    assign layer0_outputs[4375] = (inputs[180]) ^ (inputs[165]);
    assign layer0_outputs[4376] = inputs[214];
    assign layer0_outputs[4377] = inputs[208];
    assign layer0_outputs[4378] = (inputs[55]) & ~(inputs[144]);
    assign layer0_outputs[4379] = ~((inputs[11]) | (inputs[119]));
    assign layer0_outputs[4380] = ~(inputs[113]) | (inputs[66]);
    assign layer0_outputs[4381] = inputs[9];
    assign layer0_outputs[4382] = 1'b1;
    assign layer0_outputs[4383] = ~((inputs[233]) ^ (inputs[61]));
    assign layer0_outputs[4384] = ~(inputs[125]) | (inputs[242]);
    assign layer0_outputs[4385] = 1'b1;
    assign layer0_outputs[4386] = ~(inputs[123]);
    assign layer0_outputs[4387] = ~((inputs[247]) ^ (inputs[191]));
    assign layer0_outputs[4388] = ~((inputs[217]) & (inputs[162]));
    assign layer0_outputs[4389] = ~(inputs[165]);
    assign layer0_outputs[4390] = ~(inputs[118]) | (inputs[217]);
    assign layer0_outputs[4391] = ~(inputs[32]);
    assign layer0_outputs[4392] = (inputs[63]) | (inputs[227]);
    assign layer0_outputs[4393] = (inputs[214]) & ~(inputs[248]);
    assign layer0_outputs[4394] = ~((inputs[212]) ^ (inputs[127]));
    assign layer0_outputs[4395] = ~(inputs[184]) | (inputs[41]);
    assign layer0_outputs[4396] = (inputs[86]) ^ (inputs[213]);
    assign layer0_outputs[4397] = ~((inputs[128]) ^ (inputs[93]));
    assign layer0_outputs[4398] = inputs[193];
    assign layer0_outputs[4399] = (inputs[105]) & (inputs[183]);
    assign layer0_outputs[4400] = inputs[82];
    assign layer0_outputs[4401] = (inputs[196]) ^ (inputs[240]);
    assign layer0_outputs[4402] = (inputs[206]) & ~(inputs[229]);
    assign layer0_outputs[4403] = 1'b1;
    assign layer0_outputs[4404] = ~((inputs[121]) | (inputs[239]));
    assign layer0_outputs[4405] = 1'b1;
    assign layer0_outputs[4406] = ~((inputs[36]) & (inputs[59]));
    assign layer0_outputs[4407] = (inputs[169]) & ~(inputs[127]);
    assign layer0_outputs[4408] = ~(inputs[214]) | (inputs[82]);
    assign layer0_outputs[4409] = ~(inputs[159]);
    assign layer0_outputs[4410] = (inputs[255]) & ~(inputs[46]);
    assign layer0_outputs[4411] = inputs[23];
    assign layer0_outputs[4412] = 1'b1;
    assign layer0_outputs[4413] = ~(inputs[177]) | (inputs[253]);
    assign layer0_outputs[4414] = ~(inputs[152]) | (inputs[47]);
    assign layer0_outputs[4415] = 1'b0;
    assign layer0_outputs[4416] = (inputs[142]) & ~(inputs[228]);
    assign layer0_outputs[4417] = ~((inputs[9]) & (inputs[226]));
    assign layer0_outputs[4418] = inputs[228];
    assign layer0_outputs[4419] = inputs[81];
    assign layer0_outputs[4420] = ~(inputs[247]);
    assign layer0_outputs[4421] = (inputs[134]) ^ (inputs[10]);
    assign layer0_outputs[4422] = ~((inputs[135]) & (inputs[4]));
    assign layer0_outputs[4423] = (inputs[158]) & ~(inputs[147]);
    assign layer0_outputs[4424] = (inputs[168]) & ~(inputs[102]);
    assign layer0_outputs[4425] = inputs[24];
    assign layer0_outputs[4426] = ~(inputs[38]) | (inputs[191]);
    assign layer0_outputs[4427] = 1'b1;
    assign layer0_outputs[4428] = ~(inputs[234]);
    assign layer0_outputs[4429] = (inputs[116]) & ~(inputs[143]);
    assign layer0_outputs[4430] = 1'b0;
    assign layer0_outputs[4431] = (inputs[211]) & (inputs[208]);
    assign layer0_outputs[4432] = 1'b1;
    assign layer0_outputs[4433] = (inputs[92]) ^ (inputs[32]);
    assign layer0_outputs[4434] = (inputs[132]) ^ (inputs[188]);
    assign layer0_outputs[4435] = inputs[123];
    assign layer0_outputs[4436] = inputs[167];
    assign layer0_outputs[4437] = ~(inputs[17]);
    assign layer0_outputs[4438] = (inputs[79]) | (inputs[79]);
    assign layer0_outputs[4439] = ~(inputs[64]);
    assign layer0_outputs[4440] = ~(inputs[238]);
    assign layer0_outputs[4441] = inputs[176];
    assign layer0_outputs[4442] = (inputs[104]) & (inputs[72]);
    assign layer0_outputs[4443] = ~(inputs[228]) | (inputs[217]);
    assign layer0_outputs[4444] = (inputs[176]) | (inputs[206]);
    assign layer0_outputs[4445] = (inputs[225]) & ~(inputs[133]);
    assign layer0_outputs[4446] = (inputs[57]) ^ (inputs[237]);
    assign layer0_outputs[4447] = ~((inputs[16]) | (inputs[3]));
    assign layer0_outputs[4448] = (inputs[38]) & ~(inputs[133]);
    assign layer0_outputs[4449] = (inputs[34]) & ~(inputs[236]);
    assign layer0_outputs[4450] = ~(inputs[243]) | (inputs[2]);
    assign layer0_outputs[4451] = inputs[127];
    assign layer0_outputs[4452] = inputs[252];
    assign layer0_outputs[4453] = ~((inputs[200]) & (inputs[0]));
    assign layer0_outputs[4454] = (inputs[53]) & ~(inputs[158]);
    assign layer0_outputs[4455] = ~(inputs[41]);
    assign layer0_outputs[4456] = (inputs[201]) | (inputs[41]);
    assign layer0_outputs[4457] = ~((inputs[218]) | (inputs[75]));
    assign layer0_outputs[4458] = inputs[195];
    assign layer0_outputs[4459] = (inputs[135]) ^ (inputs[163]);
    assign layer0_outputs[4460] = ~(inputs[226]);
    assign layer0_outputs[4461] = (inputs[195]) & ~(inputs[15]);
    assign layer0_outputs[4462] = (inputs[71]) | (inputs[221]);
    assign layer0_outputs[4463] = ~((inputs[46]) ^ (inputs[77]));
    assign layer0_outputs[4464] = (inputs[57]) & (inputs[7]);
    assign layer0_outputs[4465] = ~(inputs[55]);
    assign layer0_outputs[4466] = (inputs[20]) & ~(inputs[140]);
    assign layer0_outputs[4467] = ~((inputs[202]) & (inputs[18]));
    assign layer0_outputs[4468] = (inputs[117]) | (inputs[149]);
    assign layer0_outputs[4469] = ~((inputs[49]) | (inputs[31]));
    assign layer0_outputs[4470] = ~((inputs[244]) & (inputs[37]));
    assign layer0_outputs[4471] = inputs[91];
    assign layer0_outputs[4472] = ~((inputs[145]) ^ (inputs[8]));
    assign layer0_outputs[4473] = 1'b0;
    assign layer0_outputs[4474] = (inputs[37]) & ~(inputs[124]);
    assign layer0_outputs[4475] = (inputs[213]) & (inputs[73]);
    assign layer0_outputs[4476] = ~((inputs[75]) & (inputs[224]));
    assign layer0_outputs[4477] = (inputs[70]) & (inputs[60]);
    assign layer0_outputs[4478] = (inputs[152]) & ~(inputs[223]);
    assign layer0_outputs[4479] = (inputs[163]) & ~(inputs[128]);
    assign layer0_outputs[4480] = 1'b0;
    assign layer0_outputs[4481] = inputs[79];
    assign layer0_outputs[4482] = 1'b0;
    assign layer0_outputs[4483] = ~((inputs[162]) & (inputs[129]));
    assign layer0_outputs[4484] = ~(inputs[223]);
    assign layer0_outputs[4485] = inputs[69];
    assign layer0_outputs[4486] = ~((inputs[128]) & (inputs[71]));
    assign layer0_outputs[4487] = ~((inputs[168]) | (inputs[222]));
    assign layer0_outputs[4488] = ~((inputs[208]) & (inputs[222]));
    assign layer0_outputs[4489] = ~(inputs[63]) | (inputs[219]);
    assign layer0_outputs[4490] = ~(inputs[196]) | (inputs[79]);
    assign layer0_outputs[4491] = ~(inputs[200]) | (inputs[18]);
    assign layer0_outputs[4492] = (inputs[251]) & ~(inputs[169]);
    assign layer0_outputs[4493] = ~((inputs[232]) ^ (inputs[123]));
    assign layer0_outputs[4494] = 1'b1;
    assign layer0_outputs[4495] = 1'b0;
    assign layer0_outputs[4496] = ~((inputs[85]) & (inputs[70]));
    assign layer0_outputs[4497] = ~(inputs[107]) | (inputs[211]);
    assign layer0_outputs[4498] = (inputs[115]) & (inputs[12]);
    assign layer0_outputs[4499] = (inputs[232]) & ~(inputs[227]);
    assign layer0_outputs[4500] = ~(inputs[206]) | (inputs[221]);
    assign layer0_outputs[4501] = ~((inputs[229]) & (inputs[108]));
    assign layer0_outputs[4502] = ~((inputs[53]) & (inputs[12]));
    assign layer0_outputs[4503] = ~((inputs[32]) ^ (inputs[87]));
    assign layer0_outputs[4504] = ~((inputs[186]) | (inputs[99]));
    assign layer0_outputs[4505] = inputs[33];
    assign layer0_outputs[4506] = (inputs[95]) & (inputs[74]);
    assign layer0_outputs[4507] = (inputs[210]) | (inputs[198]);
    assign layer0_outputs[4508] = (inputs[149]) & ~(inputs[235]);
    assign layer0_outputs[4509] = (inputs[235]) | (inputs[131]);
    assign layer0_outputs[4510] = inputs[15];
    assign layer0_outputs[4511] = (inputs[223]) & (inputs[206]);
    assign layer0_outputs[4512] = (inputs[149]) & ~(inputs[215]);
    assign layer0_outputs[4513] = (inputs[218]) | (inputs[30]);
    assign layer0_outputs[4514] = 1'b0;
    assign layer0_outputs[4515] = ~((inputs[254]) & (inputs[198]));
    assign layer0_outputs[4516] = inputs[158];
    assign layer0_outputs[4517] = (inputs[67]) & ~(inputs[0]);
    assign layer0_outputs[4518] = ~(inputs[18]) | (inputs[27]);
    assign layer0_outputs[4519] = (inputs[73]) & ~(inputs[214]);
    assign layer0_outputs[4520] = (inputs[89]) & ~(inputs[100]);
    assign layer0_outputs[4521] = (inputs[59]) ^ (inputs[194]);
    assign layer0_outputs[4522] = ~((inputs[63]) | (inputs[68]));
    assign layer0_outputs[4523] = ~(inputs[155]);
    assign layer0_outputs[4524] = 1'b0;
    assign layer0_outputs[4525] = (inputs[188]) ^ (inputs[155]);
    assign layer0_outputs[4526] = ~((inputs[144]) ^ (inputs[77]));
    assign layer0_outputs[4527] = (inputs[212]) & (inputs[32]);
    assign layer0_outputs[4528] = 1'b0;
    assign layer0_outputs[4529] = ~(inputs[139]);
    assign layer0_outputs[4530] = ~((inputs[216]) & (inputs[114]));
    assign layer0_outputs[4531] = ~((inputs[145]) ^ (inputs[21]));
    assign layer0_outputs[4532] = ~((inputs[176]) & (inputs[123]));
    assign layer0_outputs[4533] = 1'b1;
    assign layer0_outputs[4534] = (inputs[233]) & ~(inputs[93]);
    assign layer0_outputs[4535] = (inputs[89]) | (inputs[228]);
    assign layer0_outputs[4536] = ~(inputs[185]);
    assign layer0_outputs[4537] = ~((inputs[53]) ^ (inputs[126]));
    assign layer0_outputs[4538] = ~(inputs[120]) | (inputs[143]);
    assign layer0_outputs[4539] = inputs[119];
    assign layer0_outputs[4540] = (inputs[85]) & (inputs[62]);
    assign layer0_outputs[4541] = ~(inputs[35]);
    assign layer0_outputs[4542] = (inputs[104]) & ~(inputs[91]);
    assign layer0_outputs[4543] = 1'b1;
    assign layer0_outputs[4544] = inputs[67];
    assign layer0_outputs[4545] = ~(inputs[98]);
    assign layer0_outputs[4546] = (inputs[179]) & ~(inputs[245]);
    assign layer0_outputs[4547] = ~(inputs[210]);
    assign layer0_outputs[4548] = ~(inputs[25]) | (inputs[59]);
    assign layer0_outputs[4549] = (inputs[3]) & ~(inputs[158]);
    assign layer0_outputs[4550] = ~(inputs[181]);
    assign layer0_outputs[4551] = ~(inputs[127]);
    assign layer0_outputs[4552] = ~(inputs[152]);
    assign layer0_outputs[4553] = ~(inputs[65]);
    assign layer0_outputs[4554] = (inputs[232]) & ~(inputs[16]);
    assign layer0_outputs[4555] = ~((inputs[133]) | (inputs[225]));
    assign layer0_outputs[4556] = ~((inputs[251]) & (inputs[154]));
    assign layer0_outputs[4557] = 1'b0;
    assign layer0_outputs[4558] = inputs[131];
    assign layer0_outputs[4559] = ~((inputs[65]) | (inputs[14]));
    assign layer0_outputs[4560] = ~(inputs[23]) | (inputs[253]);
    assign layer0_outputs[4561] = 1'b0;
    assign layer0_outputs[4562] = inputs[140];
    assign layer0_outputs[4563] = (inputs[42]) ^ (inputs[250]);
    assign layer0_outputs[4564] = (inputs[106]) & ~(inputs[31]);
    assign layer0_outputs[4565] = ~(inputs[26]);
    assign layer0_outputs[4566] = inputs[203];
    assign layer0_outputs[4567] = 1'b0;
    assign layer0_outputs[4568] = inputs[183];
    assign layer0_outputs[4569] = (inputs[166]) & ~(inputs[71]);
    assign layer0_outputs[4570] = inputs[171];
    assign layer0_outputs[4571] = (inputs[111]) & ~(inputs[139]);
    assign layer0_outputs[4572] = 1'b0;
    assign layer0_outputs[4573] = 1'b0;
    assign layer0_outputs[4574] = (inputs[8]) | (inputs[36]);
    assign layer0_outputs[4575] = ~((inputs[101]) & (inputs[119]));
    assign layer0_outputs[4576] = ~((inputs[144]) ^ (inputs[232]));
    assign layer0_outputs[4577] = 1'b0;
    assign layer0_outputs[4578] = (inputs[207]) | (inputs[29]);
    assign layer0_outputs[4579] = ~((inputs[38]) | (inputs[245]));
    assign layer0_outputs[4580] = ~(inputs[86]) | (inputs[5]);
    assign layer0_outputs[4581] = ~(inputs[100]);
    assign layer0_outputs[4582] = ~(inputs[8]);
    assign layer0_outputs[4583] = ~((inputs[49]) & (inputs[0]));
    assign layer0_outputs[4584] = (inputs[42]) & ~(inputs[87]);
    assign layer0_outputs[4585] = ~((inputs[100]) & (inputs[120]));
    assign layer0_outputs[4586] = (inputs[205]) & ~(inputs[176]);
    assign layer0_outputs[4587] = (inputs[79]) | (inputs[174]);
    assign layer0_outputs[4588] = ~(inputs[132]);
    assign layer0_outputs[4589] = inputs[213];
    assign layer0_outputs[4590] = (inputs[54]) | (inputs[91]);
    assign layer0_outputs[4591] = (inputs[42]) & ~(inputs[242]);
    assign layer0_outputs[4592] = (inputs[69]) ^ (inputs[37]);
    assign layer0_outputs[4593] = (inputs[130]) | (inputs[89]);
    assign layer0_outputs[4594] = (inputs[23]) & ~(inputs[197]);
    assign layer0_outputs[4595] = ~(inputs[98]);
    assign layer0_outputs[4596] = 1'b0;
    assign layer0_outputs[4597] = inputs[85];
    assign layer0_outputs[4598] = (inputs[132]) ^ (inputs[126]);
    assign layer0_outputs[4599] = ~(inputs[74]);
    assign layer0_outputs[4600] = ~(inputs[1]);
    assign layer0_outputs[4601] = ~(inputs[55]);
    assign layer0_outputs[4602] = inputs[124];
    assign layer0_outputs[4603] = ~((inputs[143]) | (inputs[99]));
    assign layer0_outputs[4604] = inputs[28];
    assign layer0_outputs[4605] = ~((inputs[248]) ^ (inputs[242]));
    assign layer0_outputs[4606] = (inputs[99]) & (inputs[255]);
    assign layer0_outputs[4607] = (inputs[248]) & ~(inputs[156]);
    assign layer0_outputs[4608] = ~((inputs[181]) & (inputs[214]));
    assign layer0_outputs[4609] = (inputs[172]) & ~(inputs[89]);
    assign layer0_outputs[4610] = ~(inputs[30]) | (inputs[152]);
    assign layer0_outputs[4611] = (inputs[8]) & ~(inputs[40]);
    assign layer0_outputs[4612] = (inputs[8]) | (inputs[190]);
    assign layer0_outputs[4613] = ~((inputs[143]) ^ (inputs[7]));
    assign layer0_outputs[4614] = ~((inputs[236]) & (inputs[248]));
    assign layer0_outputs[4615] = inputs[255];
    assign layer0_outputs[4616] = inputs[141];
    assign layer0_outputs[4617] = ~(inputs[149]) | (inputs[194]);
    assign layer0_outputs[4618] = inputs[134];
    assign layer0_outputs[4619] = ~((inputs[226]) & (inputs[17]));
    assign layer0_outputs[4620] = ~((inputs[217]) | (inputs[59]));
    assign layer0_outputs[4621] = inputs[120];
    assign layer0_outputs[4622] = ~(inputs[111]);
    assign layer0_outputs[4623] = (inputs[201]) & ~(inputs[247]);
    assign layer0_outputs[4624] = (inputs[0]) & (inputs[210]);
    assign layer0_outputs[4625] = ~(inputs[157]) | (inputs[6]);
    assign layer0_outputs[4626] = (inputs[49]) & ~(inputs[232]);
    assign layer0_outputs[4627] = ~((inputs[75]) | (inputs[237]));
    assign layer0_outputs[4628] = ~(inputs[102]);
    assign layer0_outputs[4629] = ~(inputs[139]);
    assign layer0_outputs[4630] = 1'b0;
    assign layer0_outputs[4631] = ~(inputs[148]) | (inputs[208]);
    assign layer0_outputs[4632] = ~(inputs[190]) | (inputs[6]);
    assign layer0_outputs[4633] = ~(inputs[145]) | (inputs[35]);
    assign layer0_outputs[4634] = ~(inputs[149]) | (inputs[168]);
    assign layer0_outputs[4635] = ~(inputs[90]) | (inputs[45]);
    assign layer0_outputs[4636] = (inputs[84]) ^ (inputs[69]);
    assign layer0_outputs[4637] = ~((inputs[254]) ^ (inputs[164]));
    assign layer0_outputs[4638] = ~((inputs[60]) | (inputs[156]));
    assign layer0_outputs[4639] = (inputs[246]) | (inputs[50]);
    assign layer0_outputs[4640] = (inputs[50]) & ~(inputs[182]);
    assign layer0_outputs[4641] = 1'b1;
    assign layer0_outputs[4642] = 1'b1;
    assign layer0_outputs[4643] = ~(inputs[231]) | (inputs[41]);
    assign layer0_outputs[4644] = (inputs[1]) & ~(inputs[212]);
    assign layer0_outputs[4645] = (inputs[50]) | (inputs[134]);
    assign layer0_outputs[4646] = ~(inputs[189]) | (inputs[215]);
    assign layer0_outputs[4647] = (inputs[3]) & ~(inputs[100]);
    assign layer0_outputs[4648] = (inputs[249]) & ~(inputs[161]);
    assign layer0_outputs[4649] = 1'b1;
    assign layer0_outputs[4650] = ~((inputs[235]) & (inputs[194]));
    assign layer0_outputs[4651] = (inputs[142]) | (inputs[181]);
    assign layer0_outputs[4652] = ~((inputs[164]) ^ (inputs[22]));
    assign layer0_outputs[4653] = ~((inputs[175]) & (inputs[118]));
    assign layer0_outputs[4654] = inputs[244];
    assign layer0_outputs[4655] = inputs[59];
    assign layer0_outputs[4656] = ~(inputs[194]);
    assign layer0_outputs[4657] = (inputs[168]) & ~(inputs[127]);
    assign layer0_outputs[4658] = (inputs[90]) ^ (inputs[242]);
    assign layer0_outputs[4659] = ~((inputs[119]) | (inputs[0]));
    assign layer0_outputs[4660] = inputs[248];
    assign layer0_outputs[4661] = (inputs[227]) ^ (inputs[17]);
    assign layer0_outputs[4662] = inputs[97];
    assign layer0_outputs[4663] = inputs[212];
    assign layer0_outputs[4664] = (inputs[53]) | (inputs[57]);
    assign layer0_outputs[4665] = 1'b0;
    assign layer0_outputs[4666] = ~(inputs[7]);
    assign layer0_outputs[4667] = ~(inputs[51]);
    assign layer0_outputs[4668] = ~((inputs[250]) ^ (inputs[161]));
    assign layer0_outputs[4669] = ~((inputs[106]) | (inputs[18]));
    assign layer0_outputs[4670] = (inputs[150]) ^ (inputs[238]);
    assign layer0_outputs[4671] = ~(inputs[41]);
    assign layer0_outputs[4672] = (inputs[152]) & ~(inputs[255]);
    assign layer0_outputs[4673] = ~(inputs[137]) | (inputs[43]);
    assign layer0_outputs[4674] = ~(inputs[235]) | (inputs[78]);
    assign layer0_outputs[4675] = (inputs[63]) & (inputs[100]);
    assign layer0_outputs[4676] = ~(inputs[240]) | (inputs[125]);
    assign layer0_outputs[4677] = (inputs[221]) & ~(inputs[155]);
    assign layer0_outputs[4678] = ~(inputs[120]);
    assign layer0_outputs[4679] = ~((inputs[15]) & (inputs[23]));
    assign layer0_outputs[4680] = (inputs[35]) & ~(inputs[238]);
    assign layer0_outputs[4681] = inputs[108];
    assign layer0_outputs[4682] = ~(inputs[236]) | (inputs[57]);
    assign layer0_outputs[4683] = (inputs[213]) ^ (inputs[249]);
    assign layer0_outputs[4684] = ~(inputs[197]);
    assign layer0_outputs[4685] = 1'b0;
    assign layer0_outputs[4686] = inputs[36];
    assign layer0_outputs[4687] = ~(inputs[111]);
    assign layer0_outputs[4688] = 1'b0;
    assign layer0_outputs[4689] = ~((inputs[30]) | (inputs[224]));
    assign layer0_outputs[4690] = (inputs[166]) & ~(inputs[180]);
    assign layer0_outputs[4691] = ~((inputs[245]) ^ (inputs[86]));
    assign layer0_outputs[4692] = (inputs[111]) ^ (inputs[86]);
    assign layer0_outputs[4693] = 1'b1;
    assign layer0_outputs[4694] = (inputs[92]) ^ (inputs[144]);
    assign layer0_outputs[4695] = ~((inputs[0]) ^ (inputs[144]));
    assign layer0_outputs[4696] = inputs[152];
    assign layer0_outputs[4697] = 1'b0;
    assign layer0_outputs[4698] = ~(inputs[30]);
    assign layer0_outputs[4699] = (inputs[190]) ^ (inputs[139]);
    assign layer0_outputs[4700] = (inputs[197]) ^ (inputs[20]);
    assign layer0_outputs[4701] = 1'b1;
    assign layer0_outputs[4702] = ~(inputs[202]) | (inputs[69]);
    assign layer0_outputs[4703] = ~((inputs[120]) | (inputs[78]));
    assign layer0_outputs[4704] = ~((inputs[162]) | (inputs[55]));
    assign layer0_outputs[4705] = (inputs[90]) | (inputs[188]);
    assign layer0_outputs[4706] = (inputs[169]) | (inputs[140]);
    assign layer0_outputs[4707] = ~(inputs[25]);
    assign layer0_outputs[4708] = 1'b1;
    assign layer0_outputs[4709] = ~(inputs[93]) | (inputs[227]);
    assign layer0_outputs[4710] = 1'b0;
    assign layer0_outputs[4711] = inputs[23];
    assign layer0_outputs[4712] = (inputs[252]) & ~(inputs[139]);
    assign layer0_outputs[4713] = (inputs[19]) | (inputs[87]);
    assign layer0_outputs[4714] = ~(inputs[94]);
    assign layer0_outputs[4715] = (inputs[59]) & ~(inputs[11]);
    assign layer0_outputs[4716] = ~((inputs[104]) | (inputs[217]));
    assign layer0_outputs[4717] = 1'b0;
    assign layer0_outputs[4718] = (inputs[231]) & ~(inputs[101]);
    assign layer0_outputs[4719] = ~((inputs[219]) ^ (inputs[10]));
    assign layer0_outputs[4720] = (inputs[113]) | (inputs[66]);
    assign layer0_outputs[4721] = (inputs[114]) & (inputs[25]);
    assign layer0_outputs[4722] = (inputs[16]) & ~(inputs[254]);
    assign layer0_outputs[4723] = inputs[227];
    assign layer0_outputs[4724] = (inputs[8]) & ~(inputs[195]);
    assign layer0_outputs[4725] = (inputs[45]) & ~(inputs[252]);
    assign layer0_outputs[4726] = 1'b0;
    assign layer0_outputs[4727] = ~(inputs[51]) | (inputs[105]);
    assign layer0_outputs[4728] = inputs[191];
    assign layer0_outputs[4729] = 1'b1;
    assign layer0_outputs[4730] = ~(inputs[60]);
    assign layer0_outputs[4731] = ~((inputs[67]) & (inputs[128]));
    assign layer0_outputs[4732] = ~((inputs[218]) & (inputs[251]));
    assign layer0_outputs[4733] = 1'b1;
    assign layer0_outputs[4734] = ~(inputs[182]) | (inputs[130]);
    assign layer0_outputs[4735] = ~((inputs[240]) | (inputs[130]));
    assign layer0_outputs[4736] = (inputs[229]) ^ (inputs[44]);
    assign layer0_outputs[4737] = 1'b1;
    assign layer0_outputs[4738] = (inputs[174]) & (inputs[1]);
    assign layer0_outputs[4739] = (inputs[10]) | (inputs[120]);
    assign layer0_outputs[4740] = ~(inputs[64]) | (inputs[69]);
    assign layer0_outputs[4741] = ~(inputs[126]) | (inputs[96]);
    assign layer0_outputs[4742] = ~(inputs[177]);
    assign layer0_outputs[4743] = ~(inputs[138]) | (inputs[74]);
    assign layer0_outputs[4744] = 1'b0;
    assign layer0_outputs[4745] = (inputs[110]) ^ (inputs[19]);
    assign layer0_outputs[4746] = inputs[161];
    assign layer0_outputs[4747] = (inputs[51]) & (inputs[29]);
    assign layer0_outputs[4748] = ~((inputs[203]) | (inputs[196]));
    assign layer0_outputs[4749] = (inputs[118]) & ~(inputs[63]);
    assign layer0_outputs[4750] = (inputs[59]) & ~(inputs[209]);
    assign layer0_outputs[4751] = inputs[211];
    assign layer0_outputs[4752] = ~((inputs[6]) ^ (inputs[132]));
    assign layer0_outputs[4753] = (inputs[46]) ^ (inputs[62]);
    assign layer0_outputs[4754] = 1'b1;
    assign layer0_outputs[4755] = (inputs[159]) | (inputs[251]);
    assign layer0_outputs[4756] = ~((inputs[48]) & (inputs[128]));
    assign layer0_outputs[4757] = (inputs[124]) | (inputs[95]);
    assign layer0_outputs[4758] = (inputs[128]) & (inputs[138]);
    assign layer0_outputs[4759] = 1'b1;
    assign layer0_outputs[4760] = inputs[136];
    assign layer0_outputs[4761] = ~((inputs[26]) | (inputs[182]));
    assign layer0_outputs[4762] = ~(inputs[62]) | (inputs[173]);
    assign layer0_outputs[4763] = ~((inputs[206]) ^ (inputs[183]));
    assign layer0_outputs[4764] = ~(inputs[168]);
    assign layer0_outputs[4765] = (inputs[143]) | (inputs[168]);
    assign layer0_outputs[4766] = (inputs[213]) ^ (inputs[253]);
    assign layer0_outputs[4767] = ~(inputs[192]) | (inputs[35]);
    assign layer0_outputs[4768] = ~((inputs[142]) | (inputs[153]));
    assign layer0_outputs[4769] = inputs[247];
    assign layer0_outputs[4770] = inputs[167];
    assign layer0_outputs[4771] = ~((inputs[238]) & (inputs[40]));
    assign layer0_outputs[4772] = (inputs[136]) | (inputs[31]);
    assign layer0_outputs[4773] = (inputs[224]) & ~(inputs[172]);
    assign layer0_outputs[4774] = ~((inputs[75]) | (inputs[70]));
    assign layer0_outputs[4775] = ~(inputs[93]) | (inputs[144]);
    assign layer0_outputs[4776] = 1'b0;
    assign layer0_outputs[4777] = (inputs[178]) & ~(inputs[15]);
    assign layer0_outputs[4778] = (inputs[62]) & (inputs[244]);
    assign layer0_outputs[4779] = (inputs[122]) & ~(inputs[131]);
    assign layer0_outputs[4780] = 1'b0;
    assign layer0_outputs[4781] = inputs[206];
    assign layer0_outputs[4782] = ~(inputs[126]) | (inputs[76]);
    assign layer0_outputs[4783] = (inputs[117]) ^ (inputs[164]);
    assign layer0_outputs[4784] = ~((inputs[189]) & (inputs[70]));
    assign layer0_outputs[4785] = (inputs[15]) & (inputs[71]);
    assign layer0_outputs[4786] = (inputs[152]) ^ (inputs[226]);
    assign layer0_outputs[4787] = ~((inputs[152]) & (inputs[57]));
    assign layer0_outputs[4788] = 1'b0;
    assign layer0_outputs[4789] = 1'b1;
    assign layer0_outputs[4790] = ~(inputs[175]) | (inputs[2]);
    assign layer0_outputs[4791] = ~(inputs[48]) | (inputs[102]);
    assign layer0_outputs[4792] = (inputs[189]) & (inputs[105]);
    assign layer0_outputs[4793] = ~(inputs[96]);
    assign layer0_outputs[4794] = (inputs[131]) ^ (inputs[87]);
    assign layer0_outputs[4795] = 1'b0;
    assign layer0_outputs[4796] = inputs[183];
    assign layer0_outputs[4797] = (inputs[69]) & (inputs[144]);
    assign layer0_outputs[4798] = (inputs[77]) | (inputs[243]);
    assign layer0_outputs[4799] = 1'b0;
    assign layer0_outputs[4800] = 1'b1;
    assign layer0_outputs[4801] = (inputs[161]) ^ (inputs[107]);
    assign layer0_outputs[4802] = ~(inputs[105]);
    assign layer0_outputs[4803] = ~((inputs[11]) & (inputs[5]));
    assign layer0_outputs[4804] = 1'b0;
    assign layer0_outputs[4805] = inputs[247];
    assign layer0_outputs[4806] = (inputs[191]) | (inputs[185]);
    assign layer0_outputs[4807] = (inputs[207]) & ~(inputs[228]);
    assign layer0_outputs[4808] = ~(inputs[193]);
    assign layer0_outputs[4809] = ~(inputs[26]) | (inputs[248]);
    assign layer0_outputs[4810] = ~(inputs[81]);
    assign layer0_outputs[4811] = 1'b1;
    assign layer0_outputs[4812] = ~((inputs[9]) | (inputs[15]));
    assign layer0_outputs[4813] = inputs[136];
    assign layer0_outputs[4814] = (inputs[38]) | (inputs[149]);
    assign layer0_outputs[4815] = ~(inputs[12]);
    assign layer0_outputs[4816] = inputs[94];
    assign layer0_outputs[4817] = 1'b1;
    assign layer0_outputs[4818] = (inputs[88]) & ~(inputs[98]);
    assign layer0_outputs[4819] = inputs[244];
    assign layer0_outputs[4820] = 1'b0;
    assign layer0_outputs[4821] = inputs[195];
    assign layer0_outputs[4822] = ~((inputs[91]) | (inputs[104]));
    assign layer0_outputs[4823] = ~(inputs[201]) | (inputs[83]);
    assign layer0_outputs[4824] = (inputs[132]) | (inputs[84]);
    assign layer0_outputs[4825] = ~(inputs[117]);
    assign layer0_outputs[4826] = ~(inputs[32]) | (inputs[174]);
    assign layer0_outputs[4827] = (inputs[237]) ^ (inputs[84]);
    assign layer0_outputs[4828] = ~((inputs[216]) | (inputs[170]));
    assign layer0_outputs[4829] = ~((inputs[0]) | (inputs[118]));
    assign layer0_outputs[4830] = 1'b1;
    assign layer0_outputs[4831] = (inputs[146]) ^ (inputs[10]);
    assign layer0_outputs[4832] = 1'b0;
    assign layer0_outputs[4833] = ~(inputs[134]) | (inputs[127]);
    assign layer0_outputs[4834] = (inputs[255]) & ~(inputs[116]);
    assign layer0_outputs[4835] = ~(inputs[162]) | (inputs[235]);
    assign layer0_outputs[4836] = ~(inputs[247]);
    assign layer0_outputs[4837] = inputs[98];
    assign layer0_outputs[4838] = inputs[37];
    assign layer0_outputs[4839] = (inputs[242]) & ~(inputs[0]);
    assign layer0_outputs[4840] = ~(inputs[190]);
    assign layer0_outputs[4841] = inputs[71];
    assign layer0_outputs[4842] = ~((inputs[37]) ^ (inputs[28]));
    assign layer0_outputs[4843] = inputs[168];
    assign layer0_outputs[4844] = (inputs[122]) ^ (inputs[162]);
    assign layer0_outputs[4845] = ~((inputs[235]) | (inputs[52]));
    assign layer0_outputs[4846] = ~((inputs[116]) | (inputs[212]));
    assign layer0_outputs[4847] = ~(inputs[215]);
    assign layer0_outputs[4848] = ~(inputs[223]);
    assign layer0_outputs[4849] = 1'b0;
    assign layer0_outputs[4850] = ~(inputs[109]) | (inputs[28]);
    assign layer0_outputs[4851] = inputs[110];
    assign layer0_outputs[4852] = (inputs[33]) & ~(inputs[198]);
    assign layer0_outputs[4853] = inputs[13];
    assign layer0_outputs[4854] = inputs[109];
    assign layer0_outputs[4855] = ~(inputs[113]) | (inputs[208]);
    assign layer0_outputs[4856] = (inputs[98]) & ~(inputs[226]);
    assign layer0_outputs[4857] = ~(inputs[29]) | (inputs[46]);
    assign layer0_outputs[4858] = 1'b1;
    assign layer0_outputs[4859] = (inputs[240]) & (inputs[251]);
    assign layer0_outputs[4860] = (inputs[168]) & ~(inputs[15]);
    assign layer0_outputs[4861] = 1'b0;
    assign layer0_outputs[4862] = inputs[154];
    assign layer0_outputs[4863] = inputs[184];
    assign layer0_outputs[4864] = (inputs[123]) & ~(inputs[153]);
    assign layer0_outputs[4865] = ~((inputs[175]) | (inputs[212]));
    assign layer0_outputs[4866] = inputs[181];
    assign layer0_outputs[4867] = ~((inputs[65]) ^ (inputs[216]));
    assign layer0_outputs[4868] = ~(inputs[178]);
    assign layer0_outputs[4869] = ~((inputs[11]) | (inputs[138]));
    assign layer0_outputs[4870] = ~((inputs[165]) | (inputs[69]));
    assign layer0_outputs[4871] = (inputs[71]) & ~(inputs[124]);
    assign layer0_outputs[4872] = ~((inputs[94]) | (inputs[130]));
    assign layer0_outputs[4873] = ~(inputs[230]) | (inputs[172]);
    assign layer0_outputs[4874] = ~((inputs[37]) | (inputs[127]));
    assign layer0_outputs[4875] = ~(inputs[249]) | (inputs[151]);
    assign layer0_outputs[4876] = inputs[27];
    assign layer0_outputs[4877] = ~(inputs[221]) | (inputs[70]);
    assign layer0_outputs[4878] = 1'b0;
    assign layer0_outputs[4879] = inputs[56];
    assign layer0_outputs[4880] = (inputs[230]) & (inputs[42]);
    assign layer0_outputs[4881] = (inputs[213]) & ~(inputs[138]);
    assign layer0_outputs[4882] = ~((inputs[90]) | (inputs[207]));
    assign layer0_outputs[4883] = (inputs[242]) & ~(inputs[12]);
    assign layer0_outputs[4884] = (inputs[160]) ^ (inputs[90]);
    assign layer0_outputs[4885] = (inputs[231]) | (inputs[145]);
    assign layer0_outputs[4886] = (inputs[167]) & ~(inputs[5]);
    assign layer0_outputs[4887] = (inputs[129]) | (inputs[188]);
    assign layer0_outputs[4888] = inputs[140];
    assign layer0_outputs[4889] = ~(inputs[29]) | (inputs[62]);
    assign layer0_outputs[4890] = ~(inputs[117]);
    assign layer0_outputs[4891] = ~((inputs[3]) | (inputs[208]));
    assign layer0_outputs[4892] = ~((inputs[58]) | (inputs[41]));
    assign layer0_outputs[4893] = ~(inputs[85]) | (inputs[183]);
    assign layer0_outputs[4894] = ~(inputs[240]) | (inputs[155]);
    assign layer0_outputs[4895] = ~(inputs[205]);
    assign layer0_outputs[4896] = inputs[164];
    assign layer0_outputs[4897] = (inputs[122]) & (inputs[171]);
    assign layer0_outputs[4898] = ~(inputs[51]);
    assign layer0_outputs[4899] = ~(inputs[241]) | (inputs[116]);
    assign layer0_outputs[4900] = 1'b0;
    assign layer0_outputs[4901] = ~(inputs[194]);
    assign layer0_outputs[4902] = ~(inputs[81]) | (inputs[4]);
    assign layer0_outputs[4903] = 1'b0;
    assign layer0_outputs[4904] = 1'b0;
    assign layer0_outputs[4905] = inputs[243];
    assign layer0_outputs[4906] = (inputs[231]) ^ (inputs[253]);
    assign layer0_outputs[4907] = inputs[250];
    assign layer0_outputs[4908] = ~(inputs[187]);
    assign layer0_outputs[4909] = ~(inputs[227]);
    assign layer0_outputs[4910] = (inputs[234]) | (inputs[102]);
    assign layer0_outputs[4911] = inputs[127];
    assign layer0_outputs[4912] = ~(inputs[6]);
    assign layer0_outputs[4913] = (inputs[58]) & ~(inputs[207]);
    assign layer0_outputs[4914] = 1'b1;
    assign layer0_outputs[4915] = ~(inputs[68]);
    assign layer0_outputs[4916] = (inputs[163]) | (inputs[60]);
    assign layer0_outputs[4917] = (inputs[223]) & ~(inputs[159]);
    assign layer0_outputs[4918] = 1'b0;
    assign layer0_outputs[4919] = inputs[233];
    assign layer0_outputs[4920] = (inputs[140]) ^ (inputs[106]);
    assign layer0_outputs[4921] = inputs[232];
    assign layer0_outputs[4922] = (inputs[62]) ^ (inputs[58]);
    assign layer0_outputs[4923] = ~(inputs[67]);
    assign layer0_outputs[4924] = 1'b1;
    assign layer0_outputs[4925] = ~(inputs[174]) | (inputs[232]);
    assign layer0_outputs[4926] = ~((inputs[73]) & (inputs[26]));
    assign layer0_outputs[4927] = (inputs[69]) & (inputs[35]);
    assign layer0_outputs[4928] = ~((inputs[40]) | (inputs[37]));
    assign layer0_outputs[4929] = 1'b0;
    assign layer0_outputs[4930] = 1'b1;
    assign layer0_outputs[4931] = ~(inputs[107]) | (inputs[45]);
    assign layer0_outputs[4932] = 1'b0;
    assign layer0_outputs[4933] = (inputs[26]) & ~(inputs[92]);
    assign layer0_outputs[4934] = (inputs[191]) & ~(inputs[202]);
    assign layer0_outputs[4935] = ~(inputs[109]);
    assign layer0_outputs[4936] = ~((inputs[152]) & (inputs[9]));
    assign layer0_outputs[4937] = inputs[180];
    assign layer0_outputs[4938] = (inputs[139]) | (inputs[116]);
    assign layer0_outputs[4939] = inputs[157];
    assign layer0_outputs[4940] = ~((inputs[153]) | (inputs[131]));
    assign layer0_outputs[4941] = ~(inputs[29]) | (inputs[15]);
    assign layer0_outputs[4942] = ~(inputs[19]) | (inputs[137]);
    assign layer0_outputs[4943] = (inputs[240]) & ~(inputs[194]);
    assign layer0_outputs[4944] = (inputs[158]) | (inputs[209]);
    assign layer0_outputs[4945] = ~((inputs[107]) | (inputs[243]));
    assign layer0_outputs[4946] = ~(inputs[224]);
    assign layer0_outputs[4947] = (inputs[211]) | (inputs[114]);
    assign layer0_outputs[4948] = (inputs[108]) & ~(inputs[139]);
    assign layer0_outputs[4949] = ~((inputs[240]) ^ (inputs[74]));
    assign layer0_outputs[4950] = ~((inputs[226]) & (inputs[99]));
    assign layer0_outputs[4951] = (inputs[56]) & ~(inputs[14]);
    assign layer0_outputs[4952] = inputs[251];
    assign layer0_outputs[4953] = inputs[174];
    assign layer0_outputs[4954] = ~(inputs[3]);
    assign layer0_outputs[4955] = (inputs[118]) & ~(inputs[35]);
    assign layer0_outputs[4956] = inputs[109];
    assign layer0_outputs[4957] = 1'b0;
    assign layer0_outputs[4958] = inputs[131];
    assign layer0_outputs[4959] = ~((inputs[13]) ^ (inputs[234]));
    assign layer0_outputs[4960] = ~(inputs[53]) | (inputs[13]);
    assign layer0_outputs[4961] = ~(inputs[158]);
    assign layer0_outputs[4962] = inputs[191];
    assign layer0_outputs[4963] = ~((inputs[103]) & (inputs[21]));
    assign layer0_outputs[4964] = inputs[128];
    assign layer0_outputs[4965] = 1'b0;
    assign layer0_outputs[4966] = ~(inputs[198]);
    assign layer0_outputs[4967] = ~(inputs[231]) | (inputs[141]);
    assign layer0_outputs[4968] = ~(inputs[64]);
    assign layer0_outputs[4969] = (inputs[134]) & ~(inputs[223]);
    assign layer0_outputs[4970] = ~((inputs[238]) ^ (inputs[152]));
    assign layer0_outputs[4971] = inputs[107];
    assign layer0_outputs[4972] = ~((inputs[5]) & (inputs[200]));
    assign layer0_outputs[4973] = inputs[94];
    assign layer0_outputs[4974] = (inputs[134]) & ~(inputs[245]);
    assign layer0_outputs[4975] = ~((inputs[59]) ^ (inputs[187]));
    assign layer0_outputs[4976] = ~((inputs[117]) ^ (inputs[115]));
    assign layer0_outputs[4977] = 1'b0;
    assign layer0_outputs[4978] = inputs[48];
    assign layer0_outputs[4979] = 1'b1;
    assign layer0_outputs[4980] = (inputs[104]) & ~(inputs[229]);
    assign layer0_outputs[4981] = ~(inputs[130]);
    assign layer0_outputs[4982] = (inputs[245]) & ~(inputs[48]);
    assign layer0_outputs[4983] = (inputs[212]) & ~(inputs[114]);
    assign layer0_outputs[4984] = inputs[67];
    assign layer0_outputs[4985] = 1'b1;
    assign layer0_outputs[4986] = ~(inputs[36]);
    assign layer0_outputs[4987] = 1'b1;
    assign layer0_outputs[4988] = ~((inputs[226]) ^ (inputs[255]));
    assign layer0_outputs[4989] = 1'b1;
    assign layer0_outputs[4990] = (inputs[181]) & ~(inputs[244]);
    assign layer0_outputs[4991] = ~(inputs[138]);
    assign layer0_outputs[4992] = ~(inputs[251]) | (inputs[196]);
    assign layer0_outputs[4993] = (inputs[237]) & (inputs[221]);
    assign layer0_outputs[4994] = ~(inputs[162]) | (inputs[243]);
    assign layer0_outputs[4995] = inputs[68];
    assign layer0_outputs[4996] = ~((inputs[103]) & (inputs[254]));
    assign layer0_outputs[4997] = 1'b0;
    assign layer0_outputs[4998] = (inputs[238]) ^ (inputs[242]);
    assign layer0_outputs[4999] = 1'b1;
    assign layer0_outputs[5000] = ~(inputs[189]);
    assign layer0_outputs[5001] = (inputs[30]) ^ (inputs[175]);
    assign layer0_outputs[5002] = (inputs[159]) & (inputs[134]);
    assign layer0_outputs[5003] = inputs[10];
    assign layer0_outputs[5004] = (inputs[109]) & (inputs[53]);
    assign layer0_outputs[5005] = ~(inputs[179]);
    assign layer0_outputs[5006] = ~(inputs[236]);
    assign layer0_outputs[5007] = (inputs[62]) & ~(inputs[136]);
    assign layer0_outputs[5008] = 1'b1;
    assign layer0_outputs[5009] = inputs[173];
    assign layer0_outputs[5010] = inputs[240];
    assign layer0_outputs[5011] = 1'b1;
    assign layer0_outputs[5012] = (inputs[153]) & ~(inputs[209]);
    assign layer0_outputs[5013] = ~((inputs[73]) & (inputs[82]));
    assign layer0_outputs[5014] = (inputs[187]) & ~(inputs[123]);
    assign layer0_outputs[5015] = (inputs[226]) & ~(inputs[156]);
    assign layer0_outputs[5016] = ~((inputs[85]) ^ (inputs[126]));
    assign layer0_outputs[5017] = ~((inputs[86]) | (inputs[78]));
    assign layer0_outputs[5018] = inputs[145];
    assign layer0_outputs[5019] = (inputs[60]) & ~(inputs[83]);
    assign layer0_outputs[5020] = (inputs[43]) & ~(inputs[161]);
    assign layer0_outputs[5021] = inputs[12];
    assign layer0_outputs[5022] = inputs[226];
    assign layer0_outputs[5023] = (inputs[135]) & ~(inputs[236]);
    assign layer0_outputs[5024] = (inputs[134]) ^ (inputs[47]);
    assign layer0_outputs[5025] = (inputs[136]) & (inputs[29]);
    assign layer0_outputs[5026] = ~(inputs[27]) | (inputs[23]);
    assign layer0_outputs[5027] = inputs[189];
    assign layer0_outputs[5028] = ~((inputs[248]) | (inputs[79]));
    assign layer0_outputs[5029] = (inputs[28]) & ~(inputs[37]);
    assign layer0_outputs[5030] = 1'b0;
    assign layer0_outputs[5031] = inputs[189];
    assign layer0_outputs[5032] = inputs[27];
    assign layer0_outputs[5033] = (inputs[132]) ^ (inputs[64]);
    assign layer0_outputs[5034] = ~(inputs[61]);
    assign layer0_outputs[5035] = ~(inputs[122]);
    assign layer0_outputs[5036] = (inputs[240]) & ~(inputs[4]);
    assign layer0_outputs[5037] = inputs[114];
    assign layer0_outputs[5038] = (inputs[251]) & ~(inputs[254]);
    assign layer0_outputs[5039] = inputs[189];
    assign layer0_outputs[5040] = (inputs[222]) | (inputs[61]);
    assign layer0_outputs[5041] = ~(inputs[88]) | (inputs[124]);
    assign layer0_outputs[5042] = (inputs[106]) & ~(inputs[239]);
    assign layer0_outputs[5043] = (inputs[163]) | (inputs[18]);
    assign layer0_outputs[5044] = ~(inputs[65]) | (inputs[59]);
    assign layer0_outputs[5045] = 1'b0;
    assign layer0_outputs[5046] = ~((inputs[130]) | (inputs[137]));
    assign layer0_outputs[5047] = 1'b0;
    assign layer0_outputs[5048] = inputs[118];
    assign layer0_outputs[5049] = inputs[201];
    assign layer0_outputs[5050] = (inputs[36]) | (inputs[19]);
    assign layer0_outputs[5051] = (inputs[167]) & ~(inputs[62]);
    assign layer0_outputs[5052] = (inputs[34]) & (inputs[44]);
    assign layer0_outputs[5053] = ~(inputs[80]);
    assign layer0_outputs[5054] = 1'b0;
    assign layer0_outputs[5055] = (inputs[76]) ^ (inputs[240]);
    assign layer0_outputs[5056] = ~(inputs[128]);
    assign layer0_outputs[5057] = inputs[32];
    assign layer0_outputs[5058] = inputs[255];
    assign layer0_outputs[5059] = 1'b0;
    assign layer0_outputs[5060] = (inputs[46]) & ~(inputs[69]);
    assign layer0_outputs[5061] = 1'b0;
    assign layer0_outputs[5062] = inputs[139];
    assign layer0_outputs[5063] = 1'b1;
    assign layer0_outputs[5064] = inputs[16];
    assign layer0_outputs[5065] = (inputs[237]) & ~(inputs[35]);
    assign layer0_outputs[5066] = ~((inputs[56]) ^ (inputs[251]));
    assign layer0_outputs[5067] = ~(inputs[3]) | (inputs[63]);
    assign layer0_outputs[5068] = ~(inputs[207]);
    assign layer0_outputs[5069] = inputs[196];
    assign layer0_outputs[5070] = (inputs[233]) & ~(inputs[35]);
    assign layer0_outputs[5071] = ~(inputs[209]) | (inputs[20]);
    assign layer0_outputs[5072] = ~(inputs[90]) | (inputs[242]);
    assign layer0_outputs[5073] = 1'b1;
    assign layer0_outputs[5074] = 1'b1;
    assign layer0_outputs[5075] = 1'b1;
    assign layer0_outputs[5076] = (inputs[154]) & ~(inputs[96]);
    assign layer0_outputs[5077] = ~((inputs[26]) ^ (inputs[43]));
    assign layer0_outputs[5078] = 1'b1;
    assign layer0_outputs[5079] = (inputs[65]) & ~(inputs[108]);
    assign layer0_outputs[5080] = ~((inputs[245]) & (inputs[185]));
    assign layer0_outputs[5081] = (inputs[12]) & ~(inputs[162]);
    assign layer0_outputs[5082] = (inputs[42]) & ~(inputs[71]);
    assign layer0_outputs[5083] = (inputs[126]) ^ (inputs[4]);
    assign layer0_outputs[5084] = inputs[117];
    assign layer0_outputs[5085] = 1'b1;
    assign layer0_outputs[5086] = ~(inputs[175]);
    assign layer0_outputs[5087] = (inputs[142]) & (inputs[100]);
    assign layer0_outputs[5088] = 1'b1;
    assign layer0_outputs[5089] = inputs[79];
    assign layer0_outputs[5090] = ~(inputs[165]);
    assign layer0_outputs[5091] = 1'b1;
    assign layer0_outputs[5092] = ~(inputs[49]);
    assign layer0_outputs[5093] = inputs[231];
    assign layer0_outputs[5094] = inputs[22];
    assign layer0_outputs[5095] = ~(inputs[183]) | (inputs[84]);
    assign layer0_outputs[5096] = (inputs[184]) & (inputs[235]);
    assign layer0_outputs[5097] = inputs[148];
    assign layer0_outputs[5098] = inputs[43];
    assign layer0_outputs[5099] = (inputs[253]) & ~(inputs[242]);
    assign layer0_outputs[5100] = 1'b1;
    assign layer0_outputs[5101] = inputs[112];
    assign layer0_outputs[5102] = ~((inputs[20]) & (inputs[145]));
    assign layer0_outputs[5103] = ~(inputs[211]) | (inputs[197]);
    assign layer0_outputs[5104] = (inputs[209]) & ~(inputs[141]);
    assign layer0_outputs[5105] = ~(inputs[60]) | (inputs[111]);
    assign layer0_outputs[5106] = 1'b0;
    assign layer0_outputs[5107] = (inputs[0]) | (inputs[255]);
    assign layer0_outputs[5108] = ~((inputs[121]) ^ (inputs[151]));
    assign layer0_outputs[5109] = ~(inputs[248]);
    assign layer0_outputs[5110] = ~(inputs[20]);
    assign layer0_outputs[5111] = (inputs[220]) & ~(inputs[202]);
    assign layer0_outputs[5112] = (inputs[28]) & ~(inputs[6]);
    assign layer0_outputs[5113] = (inputs[77]) ^ (inputs[39]);
    assign layer0_outputs[5114] = ~((inputs[154]) ^ (inputs[217]));
    assign layer0_outputs[5115] = ~(inputs[129]);
    assign layer0_outputs[5116] = ~((inputs[137]) ^ (inputs[222]));
    assign layer0_outputs[5117] = ~(inputs[225]);
    assign layer0_outputs[5118] = (inputs[68]) & ~(inputs[88]);
    assign layer0_outputs[5119] = ~((inputs[53]) | (inputs[52]));
    assign layer1_outputs[0] = (layer0_outputs[2086]) & ~(layer0_outputs[3801]);
    assign layer1_outputs[1] = 1'b0;
    assign layer1_outputs[2] = ~(layer0_outputs[3206]) | (layer0_outputs[2915]);
    assign layer1_outputs[3] = ~(layer0_outputs[2884]) | (layer0_outputs[2120]);
    assign layer1_outputs[4] = layer0_outputs[2804];
    assign layer1_outputs[5] = (layer0_outputs[4697]) & (layer0_outputs[4011]);
    assign layer1_outputs[6] = layer0_outputs[2758];
    assign layer1_outputs[7] = 1'b0;
    assign layer1_outputs[8] = (layer0_outputs[3830]) | (layer0_outputs[1230]);
    assign layer1_outputs[9] = (layer0_outputs[262]) & ~(layer0_outputs[3706]);
    assign layer1_outputs[10] = 1'b0;
    assign layer1_outputs[11] = ~(layer0_outputs[1923]);
    assign layer1_outputs[12] = ~(layer0_outputs[2562]);
    assign layer1_outputs[13] = (layer0_outputs[3726]) & ~(layer0_outputs[3676]);
    assign layer1_outputs[14] = (layer0_outputs[3184]) & ~(layer0_outputs[582]);
    assign layer1_outputs[15] = 1'b1;
    assign layer1_outputs[16] = (layer0_outputs[3041]) | (layer0_outputs[2111]);
    assign layer1_outputs[17] = (layer0_outputs[3965]) & (layer0_outputs[4592]);
    assign layer1_outputs[18] = (layer0_outputs[2908]) ^ (layer0_outputs[4717]);
    assign layer1_outputs[19] = ~((layer0_outputs[2484]) | (layer0_outputs[4614]));
    assign layer1_outputs[20] = ~((layer0_outputs[3449]) & (layer0_outputs[716]));
    assign layer1_outputs[21] = 1'b0;
    assign layer1_outputs[22] = ~(layer0_outputs[2630]) | (layer0_outputs[3075]);
    assign layer1_outputs[23] = (layer0_outputs[209]) | (layer0_outputs[1846]);
    assign layer1_outputs[24] = (layer0_outputs[3901]) & ~(layer0_outputs[5033]);
    assign layer1_outputs[25] = (layer0_outputs[3572]) & ~(layer0_outputs[1204]);
    assign layer1_outputs[26] = ~(layer0_outputs[2993]) | (layer0_outputs[2493]);
    assign layer1_outputs[27] = (layer0_outputs[2334]) & (layer0_outputs[1365]);
    assign layer1_outputs[28] = (layer0_outputs[2289]) | (layer0_outputs[3259]);
    assign layer1_outputs[29] = 1'b0;
    assign layer1_outputs[30] = 1'b1;
    assign layer1_outputs[31] = 1'b1;
    assign layer1_outputs[32] = ~((layer0_outputs[2874]) & (layer0_outputs[117]));
    assign layer1_outputs[33] = (layer0_outputs[1181]) | (layer0_outputs[3197]);
    assign layer1_outputs[34] = ~(layer0_outputs[4336]) | (layer0_outputs[4207]);
    assign layer1_outputs[35] = 1'b1;
    assign layer1_outputs[36] = (layer0_outputs[4543]) | (layer0_outputs[0]);
    assign layer1_outputs[37] = (layer0_outputs[2152]) & ~(layer0_outputs[229]);
    assign layer1_outputs[38] = ~((layer0_outputs[822]) | (layer0_outputs[3490]));
    assign layer1_outputs[39] = 1'b1;
    assign layer1_outputs[40] = ~((layer0_outputs[4291]) & (layer0_outputs[953]));
    assign layer1_outputs[41] = (layer0_outputs[2138]) & ~(layer0_outputs[4269]);
    assign layer1_outputs[42] = ~((layer0_outputs[888]) & (layer0_outputs[3316]));
    assign layer1_outputs[43] = ~((layer0_outputs[1060]) | (layer0_outputs[4914]));
    assign layer1_outputs[44] = 1'b1;
    assign layer1_outputs[45] = ~((layer0_outputs[1542]) & (layer0_outputs[2981]));
    assign layer1_outputs[46] = (layer0_outputs[1857]) & (layer0_outputs[980]);
    assign layer1_outputs[47] = (layer0_outputs[5019]) ^ (layer0_outputs[2117]);
    assign layer1_outputs[48] = layer0_outputs[2398];
    assign layer1_outputs[49] = (layer0_outputs[5111]) & ~(layer0_outputs[4676]);
    assign layer1_outputs[50] = ~(layer0_outputs[2192]) | (layer0_outputs[3080]);
    assign layer1_outputs[51] = ~(layer0_outputs[3936]);
    assign layer1_outputs[52] = ~(layer0_outputs[465]);
    assign layer1_outputs[53] = 1'b0;
    assign layer1_outputs[54] = ~((layer0_outputs[2530]) | (layer0_outputs[2774]));
    assign layer1_outputs[55] = (layer0_outputs[2528]) & ~(layer0_outputs[642]);
    assign layer1_outputs[56] = ~((layer0_outputs[4848]) & (layer0_outputs[2948]));
    assign layer1_outputs[57] = (layer0_outputs[4420]) & ~(layer0_outputs[4271]);
    assign layer1_outputs[58] = ~(layer0_outputs[965]) | (layer0_outputs[1039]);
    assign layer1_outputs[59] = (layer0_outputs[1319]) & ~(layer0_outputs[71]);
    assign layer1_outputs[60] = (layer0_outputs[269]) | (layer0_outputs[4343]);
    assign layer1_outputs[61] = ~((layer0_outputs[1187]) ^ (layer0_outputs[4488]));
    assign layer1_outputs[62] = (layer0_outputs[908]) & (layer0_outputs[3614]);
    assign layer1_outputs[63] = ~(layer0_outputs[3558]);
    assign layer1_outputs[64] = (layer0_outputs[4922]) & (layer0_outputs[3300]);
    assign layer1_outputs[65] = (layer0_outputs[1762]) | (layer0_outputs[2148]);
    assign layer1_outputs[66] = 1'b1;
    assign layer1_outputs[67] = ~(layer0_outputs[1632]) | (layer0_outputs[2880]);
    assign layer1_outputs[68] = ~(layer0_outputs[3830]) | (layer0_outputs[3604]);
    assign layer1_outputs[69] = ~((layer0_outputs[670]) & (layer0_outputs[1832]));
    assign layer1_outputs[70] = ~(layer0_outputs[2162]) | (layer0_outputs[3500]);
    assign layer1_outputs[71] = ~(layer0_outputs[3734]);
    assign layer1_outputs[72] = 1'b0;
    assign layer1_outputs[73] = layer0_outputs[3738];
    assign layer1_outputs[74] = ~((layer0_outputs[947]) | (layer0_outputs[4945]));
    assign layer1_outputs[75] = ~((layer0_outputs[140]) & (layer0_outputs[4783]));
    assign layer1_outputs[76] = 1'b1;
    assign layer1_outputs[77] = layer0_outputs[4786];
    assign layer1_outputs[78] = layer0_outputs[2625];
    assign layer1_outputs[79] = ~(layer0_outputs[2013]);
    assign layer1_outputs[80] = (layer0_outputs[391]) | (layer0_outputs[2093]);
    assign layer1_outputs[81] = (layer0_outputs[1031]) | (layer0_outputs[1100]);
    assign layer1_outputs[82] = ~(layer0_outputs[296]);
    assign layer1_outputs[83] = 1'b0;
    assign layer1_outputs[84] = ~(layer0_outputs[4166]);
    assign layer1_outputs[85] = ~(layer0_outputs[2379]) | (layer0_outputs[1741]);
    assign layer1_outputs[86] = ~(layer0_outputs[2023]);
    assign layer1_outputs[87] = ~(layer0_outputs[5107]) | (layer0_outputs[4542]);
    assign layer1_outputs[88] = layer0_outputs[3034];
    assign layer1_outputs[89] = ~(layer0_outputs[4425]);
    assign layer1_outputs[90] = layer0_outputs[2769];
    assign layer1_outputs[91] = (layer0_outputs[3172]) | (layer0_outputs[5103]);
    assign layer1_outputs[92] = (layer0_outputs[4689]) | (layer0_outputs[2632]);
    assign layer1_outputs[93] = (layer0_outputs[3296]) | (layer0_outputs[4305]);
    assign layer1_outputs[94] = ~(layer0_outputs[453]);
    assign layer1_outputs[95] = ~((layer0_outputs[1125]) | (layer0_outputs[1758]));
    assign layer1_outputs[96] = (layer0_outputs[2056]) | (layer0_outputs[1673]);
    assign layer1_outputs[97] = 1'b1;
    assign layer1_outputs[98] = ~(layer0_outputs[4330]);
    assign layer1_outputs[99] = (layer0_outputs[142]) ^ (layer0_outputs[2271]);
    assign layer1_outputs[100] = layer0_outputs[3271];
    assign layer1_outputs[101] = layer0_outputs[351];
    assign layer1_outputs[102] = layer0_outputs[3752];
    assign layer1_outputs[103] = (layer0_outputs[2568]) | (layer0_outputs[1492]);
    assign layer1_outputs[104] = ~(layer0_outputs[4480]) | (layer0_outputs[1536]);
    assign layer1_outputs[105] = 1'b1;
    assign layer1_outputs[106] = layer0_outputs[1225];
    assign layer1_outputs[107] = layer0_outputs[422];
    assign layer1_outputs[108] = layer0_outputs[1002];
    assign layer1_outputs[109] = (layer0_outputs[2946]) | (layer0_outputs[4907]);
    assign layer1_outputs[110] = layer0_outputs[1211];
    assign layer1_outputs[111] = (layer0_outputs[2841]) & ~(layer0_outputs[1548]);
    assign layer1_outputs[112] = ~((layer0_outputs[4630]) ^ (layer0_outputs[3065]));
    assign layer1_outputs[113] = (layer0_outputs[2270]) & (layer0_outputs[1324]);
    assign layer1_outputs[114] = ~(layer0_outputs[4921]) | (layer0_outputs[2603]);
    assign layer1_outputs[115] = ~((layer0_outputs[3974]) | (layer0_outputs[779]));
    assign layer1_outputs[116] = ~(layer0_outputs[1604]);
    assign layer1_outputs[117] = 1'b1;
    assign layer1_outputs[118] = (layer0_outputs[1489]) | (layer0_outputs[3390]);
    assign layer1_outputs[119] = 1'b1;
    assign layer1_outputs[120] = (layer0_outputs[4388]) | (layer0_outputs[3108]);
    assign layer1_outputs[121] = 1'b0;
    assign layer1_outputs[122] = 1'b0;
    assign layer1_outputs[123] = ~((layer0_outputs[266]) ^ (layer0_outputs[62]));
    assign layer1_outputs[124] = (layer0_outputs[2669]) & (layer0_outputs[1017]);
    assign layer1_outputs[125] = ~(layer0_outputs[2201]) | (layer0_outputs[1874]);
    assign layer1_outputs[126] = ~((layer0_outputs[3278]) ^ (layer0_outputs[1179]));
    assign layer1_outputs[127] = ~((layer0_outputs[4680]) | (layer0_outputs[776]));
    assign layer1_outputs[128] = (layer0_outputs[3984]) & (layer0_outputs[2147]);
    assign layer1_outputs[129] = ~(layer0_outputs[3388]) | (layer0_outputs[374]);
    assign layer1_outputs[130] = (layer0_outputs[3896]) & ~(layer0_outputs[1183]);
    assign layer1_outputs[131] = (layer0_outputs[1173]) & ~(layer0_outputs[4442]);
    assign layer1_outputs[132] = ~((layer0_outputs[2857]) & (layer0_outputs[4910]));
    assign layer1_outputs[133] = 1'b0;
    assign layer1_outputs[134] = (layer0_outputs[919]) & (layer0_outputs[3332]);
    assign layer1_outputs[135] = (layer0_outputs[244]) & (layer0_outputs[869]);
    assign layer1_outputs[136] = ~((layer0_outputs[5117]) ^ (layer0_outputs[1545]));
    assign layer1_outputs[137] = (layer0_outputs[3373]) & (layer0_outputs[1992]);
    assign layer1_outputs[138] = 1'b1;
    assign layer1_outputs[139] = ~(layer0_outputs[4192]);
    assign layer1_outputs[140] = ~(layer0_outputs[4168]) | (layer0_outputs[340]);
    assign layer1_outputs[141] = ~(layer0_outputs[2383]);
    assign layer1_outputs[142] = ~(layer0_outputs[1429]);
    assign layer1_outputs[143] = (layer0_outputs[2183]) & ~(layer0_outputs[20]);
    assign layer1_outputs[144] = layer0_outputs[1972];
    assign layer1_outputs[145] = 1'b1;
    assign layer1_outputs[146] = ~((layer0_outputs[4465]) & (layer0_outputs[4535]));
    assign layer1_outputs[147] = 1'b0;
    assign layer1_outputs[148] = ~(layer0_outputs[2961]);
    assign layer1_outputs[149] = (layer0_outputs[4874]) & ~(layer0_outputs[1689]);
    assign layer1_outputs[150] = (layer0_outputs[353]) & ~(layer0_outputs[3183]);
    assign layer1_outputs[151] = layer0_outputs[1629];
    assign layer1_outputs[152] = 1'b1;
    assign layer1_outputs[153] = ~(layer0_outputs[612]) | (layer0_outputs[3120]);
    assign layer1_outputs[154] = (layer0_outputs[1903]) | (layer0_outputs[3875]);
    assign layer1_outputs[155] = layer0_outputs[3927];
    assign layer1_outputs[156] = (layer0_outputs[3407]) | (layer0_outputs[1162]);
    assign layer1_outputs[157] = 1'b0;
    assign layer1_outputs[158] = ~((layer0_outputs[4161]) & (layer0_outputs[1246]));
    assign layer1_outputs[159] = ~((layer0_outputs[2360]) & (layer0_outputs[4529]));
    assign layer1_outputs[160] = ~((layer0_outputs[426]) | (layer0_outputs[1653]));
    assign layer1_outputs[161] = layer0_outputs[3219];
    assign layer1_outputs[162] = (layer0_outputs[3003]) & ~(layer0_outputs[688]);
    assign layer1_outputs[163] = 1'b1;
    assign layer1_outputs[164] = 1'b0;
    assign layer1_outputs[165] = 1'b1;
    assign layer1_outputs[166] = 1'b1;
    assign layer1_outputs[167] = 1'b0;
    assign layer1_outputs[168] = layer0_outputs[1516];
    assign layer1_outputs[169] = ~(layer0_outputs[1609]);
    assign layer1_outputs[170] = ~(layer0_outputs[4451]);
    assign layer1_outputs[171] = ~((layer0_outputs[3073]) ^ (layer0_outputs[3339]));
    assign layer1_outputs[172] = 1'b0;
    assign layer1_outputs[173] = 1'b1;
    assign layer1_outputs[174] = 1'b0;
    assign layer1_outputs[175] = (layer0_outputs[432]) & ~(layer0_outputs[3893]);
    assign layer1_outputs[176] = ~((layer0_outputs[1724]) | (layer0_outputs[1586]));
    assign layer1_outputs[177] = layer0_outputs[1222];
    assign layer1_outputs[178] = (layer0_outputs[4015]) | (layer0_outputs[2801]);
    assign layer1_outputs[179] = (layer0_outputs[604]) & (layer0_outputs[96]);
    assign layer1_outputs[180] = 1'b1;
    assign layer1_outputs[181] = (layer0_outputs[3045]) | (layer0_outputs[5075]);
    assign layer1_outputs[182] = 1'b0;
    assign layer1_outputs[183] = ~(layer0_outputs[4171]) | (layer0_outputs[4725]);
    assign layer1_outputs[184] = (layer0_outputs[261]) & ~(layer0_outputs[3630]);
    assign layer1_outputs[185] = ~(layer0_outputs[3503]);
    assign layer1_outputs[186] = 1'b1;
    assign layer1_outputs[187] = (layer0_outputs[2767]) & ~(layer0_outputs[95]);
    assign layer1_outputs[188] = 1'b0;
    assign layer1_outputs[189] = (layer0_outputs[4388]) & (layer0_outputs[3570]);
    assign layer1_outputs[190] = ~(layer0_outputs[4351]) | (layer0_outputs[5063]);
    assign layer1_outputs[191] = ~((layer0_outputs[1185]) ^ (layer0_outputs[4083]));
    assign layer1_outputs[192] = ~((layer0_outputs[4607]) | (layer0_outputs[4571]));
    assign layer1_outputs[193] = layer0_outputs[3712];
    assign layer1_outputs[194] = ~((layer0_outputs[5072]) & (layer0_outputs[2245]));
    assign layer1_outputs[195] = ~((layer0_outputs[2876]) & (layer0_outputs[4007]));
    assign layer1_outputs[196] = 1'b1;
    assign layer1_outputs[197] = layer0_outputs[79];
    assign layer1_outputs[198] = 1'b0;
    assign layer1_outputs[199] = ~(layer0_outputs[3381]) | (layer0_outputs[2991]);
    assign layer1_outputs[200] = (layer0_outputs[3315]) ^ (layer0_outputs[493]);
    assign layer1_outputs[201] = ~(layer0_outputs[4669]);
    assign layer1_outputs[202] = layer0_outputs[1477];
    assign layer1_outputs[203] = layer0_outputs[4788];
    assign layer1_outputs[204] = (layer0_outputs[2776]) & ~(layer0_outputs[2766]);
    assign layer1_outputs[205] = 1'b1;
    assign layer1_outputs[206] = (layer0_outputs[4371]) & (layer0_outputs[121]);
    assign layer1_outputs[207] = 1'b0;
    assign layer1_outputs[208] = layer0_outputs[3427];
    assign layer1_outputs[209] = layer0_outputs[3422];
    assign layer1_outputs[210] = ~(layer0_outputs[3838]) | (layer0_outputs[251]);
    assign layer1_outputs[211] = layer0_outputs[433];
    assign layer1_outputs[212] = layer0_outputs[2635];
    assign layer1_outputs[213] = (layer0_outputs[2434]) | (layer0_outputs[1756]);
    assign layer1_outputs[214] = ~(layer0_outputs[4757]) | (layer0_outputs[2664]);
    assign layer1_outputs[215] = ~((layer0_outputs[4511]) | (layer0_outputs[3113]));
    assign layer1_outputs[216] = ~((layer0_outputs[148]) & (layer0_outputs[414]));
    assign layer1_outputs[217] = 1'b1;
    assign layer1_outputs[218] = (layer0_outputs[3452]) & (layer0_outputs[87]);
    assign layer1_outputs[219] = layer0_outputs[2912];
    assign layer1_outputs[220] = (layer0_outputs[5009]) & ~(layer0_outputs[4353]);
    assign layer1_outputs[221] = (layer0_outputs[3851]) | (layer0_outputs[349]);
    assign layer1_outputs[222] = layer0_outputs[4921];
    assign layer1_outputs[223] = ~(layer0_outputs[1559]) | (layer0_outputs[3700]);
    assign layer1_outputs[224] = 1'b0;
    assign layer1_outputs[225] = ~(layer0_outputs[3872]) | (layer0_outputs[3841]);
    assign layer1_outputs[226] = (layer0_outputs[4899]) & (layer0_outputs[3580]);
    assign layer1_outputs[227] = ~(layer0_outputs[559]);
    assign layer1_outputs[228] = ~((layer0_outputs[1104]) ^ (layer0_outputs[1413]));
    assign layer1_outputs[229] = layer0_outputs[3517];
    assign layer1_outputs[230] = layer0_outputs[3718];
    assign layer1_outputs[231] = (layer0_outputs[4530]) | (layer0_outputs[966]);
    assign layer1_outputs[232] = layer0_outputs[1173];
    assign layer1_outputs[233] = ~(layer0_outputs[4100]) | (layer0_outputs[3248]);
    assign layer1_outputs[234] = ~(layer0_outputs[4885]) | (layer0_outputs[1933]);
    assign layer1_outputs[235] = (layer0_outputs[2286]) & ~(layer0_outputs[228]);
    assign layer1_outputs[236] = layer0_outputs[4986];
    assign layer1_outputs[237] = ~(layer0_outputs[3221]);
    assign layer1_outputs[238] = ~(layer0_outputs[4121]);
    assign layer1_outputs[239] = ~((layer0_outputs[3304]) | (layer0_outputs[2498]));
    assign layer1_outputs[240] = (layer0_outputs[3541]) & (layer0_outputs[1887]);
    assign layer1_outputs[241] = ~(layer0_outputs[3040]) | (layer0_outputs[1318]);
    assign layer1_outputs[242] = (layer0_outputs[3876]) & (layer0_outputs[1264]);
    assign layer1_outputs[243] = (layer0_outputs[1111]) & (layer0_outputs[1886]);
    assign layer1_outputs[244] = ~(layer0_outputs[2168]);
    assign layer1_outputs[245] = ~((layer0_outputs[3387]) ^ (layer0_outputs[1949]));
    assign layer1_outputs[246] = layer0_outputs[2801];
    assign layer1_outputs[247] = layer0_outputs[3118];
    assign layer1_outputs[248] = ~((layer0_outputs[3493]) | (layer0_outputs[3622]));
    assign layer1_outputs[249] = ~((layer0_outputs[2871]) | (layer0_outputs[1394]));
    assign layer1_outputs[250] = (layer0_outputs[3005]) ^ (layer0_outputs[2079]);
    assign layer1_outputs[251] = ~(layer0_outputs[2202]) | (layer0_outputs[3141]);
    assign layer1_outputs[252] = ~(layer0_outputs[2762]) | (layer0_outputs[2488]);
    assign layer1_outputs[253] = ~((layer0_outputs[4596]) & (layer0_outputs[306]));
    assign layer1_outputs[254] = ~((layer0_outputs[4089]) | (layer0_outputs[9]));
    assign layer1_outputs[255] = layer0_outputs[652];
    assign layer1_outputs[256] = (layer0_outputs[2931]) & ~(layer0_outputs[3764]);
    assign layer1_outputs[257] = (layer0_outputs[808]) & (layer0_outputs[4269]);
    assign layer1_outputs[258] = layer0_outputs[559];
    assign layer1_outputs[259] = ~((layer0_outputs[4196]) & (layer0_outputs[3338]));
    assign layer1_outputs[260] = ~(layer0_outputs[4589]);
    assign layer1_outputs[261] = ~(layer0_outputs[2729]) | (layer0_outputs[1355]);
    assign layer1_outputs[262] = 1'b0;
    assign layer1_outputs[263] = ~(layer0_outputs[1701]);
    assign layer1_outputs[264] = (layer0_outputs[3599]) & (layer0_outputs[286]);
    assign layer1_outputs[265] = (layer0_outputs[1823]) & ~(layer0_outputs[1351]);
    assign layer1_outputs[266] = 1'b0;
    assign layer1_outputs[267] = 1'b0;
    assign layer1_outputs[268] = ~(layer0_outputs[3001]);
    assign layer1_outputs[269] = ~(layer0_outputs[1281]) | (layer0_outputs[542]);
    assign layer1_outputs[270] = ~(layer0_outputs[59]);
    assign layer1_outputs[271] = 1'b0;
    assign layer1_outputs[272] = ~((layer0_outputs[1608]) | (layer0_outputs[4257]));
    assign layer1_outputs[273] = layer0_outputs[2565];
    assign layer1_outputs[274] = ~((layer0_outputs[1796]) & (layer0_outputs[4264]));
    assign layer1_outputs[275] = layer0_outputs[1915];
    assign layer1_outputs[276] = 1'b0;
    assign layer1_outputs[277] = ~((layer0_outputs[1950]) & (layer0_outputs[3695]));
    assign layer1_outputs[278] = (layer0_outputs[4165]) & ~(layer0_outputs[1983]);
    assign layer1_outputs[279] = (layer0_outputs[265]) & ~(layer0_outputs[2474]);
    assign layer1_outputs[280] = 1'b0;
    assign layer1_outputs[281] = ~(layer0_outputs[4562]);
    assign layer1_outputs[282] = ~((layer0_outputs[2524]) & (layer0_outputs[843]));
    assign layer1_outputs[283] = (layer0_outputs[3149]) & (layer0_outputs[1068]);
    assign layer1_outputs[284] = (layer0_outputs[2898]) & (layer0_outputs[2787]);
    assign layer1_outputs[285] = layer0_outputs[1528];
    assign layer1_outputs[286] = ~((layer0_outputs[339]) | (layer0_outputs[3821]));
    assign layer1_outputs[287] = ~(layer0_outputs[114]) | (layer0_outputs[2881]);
    assign layer1_outputs[288] = 1'b0;
    assign layer1_outputs[289] = layer0_outputs[4538];
    assign layer1_outputs[290] = (layer0_outputs[4499]) | (layer0_outputs[301]);
    assign layer1_outputs[291] = (layer0_outputs[2967]) | (layer0_outputs[734]);
    assign layer1_outputs[292] = layer0_outputs[2596];
    assign layer1_outputs[293] = 1'b1;
    assign layer1_outputs[294] = layer0_outputs[1540];
    assign layer1_outputs[295] = ~(layer0_outputs[1233]) | (layer0_outputs[3479]);
    assign layer1_outputs[296] = (layer0_outputs[1628]) & ~(layer0_outputs[4710]);
    assign layer1_outputs[297] = (layer0_outputs[573]) ^ (layer0_outputs[67]);
    assign layer1_outputs[298] = (layer0_outputs[4062]) & ~(layer0_outputs[2589]);
    assign layer1_outputs[299] = layer0_outputs[1499];
    assign layer1_outputs[300] = 1'b1;
    assign layer1_outputs[301] = ~(layer0_outputs[592]);
    assign layer1_outputs[302] = ~((layer0_outputs[2838]) & (layer0_outputs[2741]));
    assign layer1_outputs[303] = (layer0_outputs[1363]) | (layer0_outputs[3739]);
    assign layer1_outputs[304] = 1'b1;
    assign layer1_outputs[305] = ~(layer0_outputs[3752]);
    assign layer1_outputs[306] = layer0_outputs[4664];
    assign layer1_outputs[307] = ~(layer0_outputs[4669]);
    assign layer1_outputs[308] = ~((layer0_outputs[4347]) & (layer0_outputs[2320]));
    assign layer1_outputs[309] = (layer0_outputs[3799]) & ~(layer0_outputs[1256]);
    assign layer1_outputs[310] = 1'b1;
    assign layer1_outputs[311] = ~(layer0_outputs[1194]) | (layer0_outputs[2738]);
    assign layer1_outputs[312] = ~(layer0_outputs[667]);
    assign layer1_outputs[313] = ~((layer0_outputs[1853]) ^ (layer0_outputs[4845]));
    assign layer1_outputs[314] = layer0_outputs[4701];
    assign layer1_outputs[315] = 1'b1;
    assign layer1_outputs[316] = ~((layer0_outputs[225]) & (layer0_outputs[898]));
    assign layer1_outputs[317] = (layer0_outputs[5081]) & (layer0_outputs[4849]);
    assign layer1_outputs[318] = 1'b0;
    assign layer1_outputs[319] = layer0_outputs[1086];
    assign layer1_outputs[320] = ~((layer0_outputs[2410]) | (layer0_outputs[4243]));
    assign layer1_outputs[321] = 1'b0;
    assign layer1_outputs[322] = (layer0_outputs[4922]) & ~(layer0_outputs[3136]);
    assign layer1_outputs[323] = layer0_outputs[4587];
    assign layer1_outputs[324] = ~((layer0_outputs[4433]) ^ (layer0_outputs[3243]));
    assign layer1_outputs[325] = ~((layer0_outputs[4281]) | (layer0_outputs[4287]));
    assign layer1_outputs[326] = 1'b0;
    assign layer1_outputs[327] = layer0_outputs[3277];
    assign layer1_outputs[328] = (layer0_outputs[3161]) & ~(layer0_outputs[3420]);
    assign layer1_outputs[329] = ~(layer0_outputs[3868]) | (layer0_outputs[4588]);
    assign layer1_outputs[330] = ~(layer0_outputs[971]);
    assign layer1_outputs[331] = (layer0_outputs[3604]) | (layer0_outputs[3438]);
    assign layer1_outputs[332] = (layer0_outputs[3952]) & ~(layer0_outputs[2753]);
    assign layer1_outputs[333] = layer0_outputs[2534];
    assign layer1_outputs[334] = 1'b1;
    assign layer1_outputs[335] = (layer0_outputs[1486]) ^ (layer0_outputs[556]);
    assign layer1_outputs[336] = (layer0_outputs[3610]) | (layer0_outputs[2426]);
    assign layer1_outputs[337] = ~((layer0_outputs[2091]) ^ (layer0_outputs[4234]));
    assign layer1_outputs[338] = ~((layer0_outputs[3552]) & (layer0_outputs[3469]));
    assign layer1_outputs[339] = ~(layer0_outputs[2984]) | (layer0_outputs[5057]);
    assign layer1_outputs[340] = ~(layer0_outputs[945]);
    assign layer1_outputs[341] = ~(layer0_outputs[864]);
    assign layer1_outputs[342] = ~((layer0_outputs[4635]) | (layer0_outputs[1427]));
    assign layer1_outputs[343] = ~((layer0_outputs[931]) | (layer0_outputs[1556]));
    assign layer1_outputs[344] = layer0_outputs[339];
    assign layer1_outputs[345] = 1'b0;
    assign layer1_outputs[346] = 1'b1;
    assign layer1_outputs[347] = ~(layer0_outputs[4573]);
    assign layer1_outputs[348] = 1'b0;
    assign layer1_outputs[349] = (layer0_outputs[1581]) & ~(layer0_outputs[4284]);
    assign layer1_outputs[350] = (layer0_outputs[2490]) & ~(layer0_outputs[1818]);
    assign layer1_outputs[351] = 1'b1;
    assign layer1_outputs[352] = (layer0_outputs[2704]) | (layer0_outputs[657]);
    assign layer1_outputs[353] = 1'b1;
    assign layer1_outputs[354] = ~((layer0_outputs[790]) ^ (layer0_outputs[3095]));
    assign layer1_outputs[355] = layer0_outputs[3905];
    assign layer1_outputs[356] = layer0_outputs[595];
    assign layer1_outputs[357] = ~(layer0_outputs[962]);
    assign layer1_outputs[358] = ~(layer0_outputs[2140]) | (layer0_outputs[1174]);
    assign layer1_outputs[359] = (layer0_outputs[423]) & (layer0_outputs[3962]);
    assign layer1_outputs[360] = (layer0_outputs[2385]) | (layer0_outputs[1517]);
    assign layer1_outputs[361] = 1'b1;
    assign layer1_outputs[362] = ~(layer0_outputs[4436]);
    assign layer1_outputs[363] = 1'b1;
    assign layer1_outputs[364] = ~((layer0_outputs[5102]) | (layer0_outputs[2345]));
    assign layer1_outputs[365] = ~((layer0_outputs[2537]) | (layer0_outputs[4242]));
    assign layer1_outputs[366] = layer0_outputs[1847];
    assign layer1_outputs[367] = ~(layer0_outputs[2504]) | (layer0_outputs[3582]);
    assign layer1_outputs[368] = ~(layer0_outputs[646]) | (layer0_outputs[4623]);
    assign layer1_outputs[369] = (layer0_outputs[468]) & (layer0_outputs[2176]);
    assign layer1_outputs[370] = 1'b1;
    assign layer1_outputs[371] = 1'b1;
    assign layer1_outputs[372] = layer0_outputs[1918];
    assign layer1_outputs[373] = (layer0_outputs[5029]) & ~(layer0_outputs[92]);
    assign layer1_outputs[374] = ~((layer0_outputs[1289]) & (layer0_outputs[4101]));
    assign layer1_outputs[375] = 1'b0;
    assign layer1_outputs[376] = ~((layer0_outputs[5073]) | (layer0_outputs[4714]));
    assign layer1_outputs[377] = ~((layer0_outputs[674]) ^ (layer0_outputs[3084]));
    assign layer1_outputs[378] = 1'b1;
    assign layer1_outputs[379] = layer0_outputs[2572];
    assign layer1_outputs[380] = (layer0_outputs[1350]) & ~(layer0_outputs[3363]);
    assign layer1_outputs[381] = ~(layer0_outputs[848]) | (layer0_outputs[388]);
    assign layer1_outputs[382] = 1'b1;
    assign layer1_outputs[383] = (layer0_outputs[3729]) & (layer0_outputs[4681]);
    assign layer1_outputs[384] = ~(layer0_outputs[5005]);
    assign layer1_outputs[385] = 1'b1;
    assign layer1_outputs[386] = ~((layer0_outputs[177]) & (layer0_outputs[3699]));
    assign layer1_outputs[387] = ~((layer0_outputs[2713]) & (layer0_outputs[1411]));
    assign layer1_outputs[388] = 1'b1;
    assign layer1_outputs[389] = layer0_outputs[2529];
    assign layer1_outputs[390] = (layer0_outputs[2030]) & ~(layer0_outputs[1496]);
    assign layer1_outputs[391] = ~(layer0_outputs[4851]);
    assign layer1_outputs[392] = ~(layer0_outputs[3128]);
    assign layer1_outputs[393] = (layer0_outputs[4467]) & ~(layer0_outputs[2522]);
    assign layer1_outputs[394] = 1'b0;
    assign layer1_outputs[395] = (layer0_outputs[1771]) & ~(layer0_outputs[1755]);
    assign layer1_outputs[396] = (layer0_outputs[3303]) & ~(layer0_outputs[3423]);
    assign layer1_outputs[397] = (layer0_outputs[3063]) | (layer0_outputs[3132]);
    assign layer1_outputs[398] = layer0_outputs[2877];
    assign layer1_outputs[399] = layer0_outputs[475];
    assign layer1_outputs[400] = 1'b1;
    assign layer1_outputs[401] = layer0_outputs[4018];
    assign layer1_outputs[402] = layer0_outputs[3017];
    assign layer1_outputs[403] = (layer0_outputs[2704]) & ~(layer0_outputs[3570]);
    assign layer1_outputs[404] = layer0_outputs[4945];
    assign layer1_outputs[405] = (layer0_outputs[3302]) & (layer0_outputs[3581]);
    assign layer1_outputs[406] = ~(layer0_outputs[3352]) | (layer0_outputs[3021]);
    assign layer1_outputs[407] = (layer0_outputs[3624]) & ~(layer0_outputs[1820]);
    assign layer1_outputs[408] = (layer0_outputs[4665]) & ~(layer0_outputs[529]);
    assign layer1_outputs[409] = ~((layer0_outputs[2776]) ^ (layer0_outputs[3560]));
    assign layer1_outputs[410] = ~(layer0_outputs[575]);
    assign layer1_outputs[411] = ~(layer0_outputs[1596]) | (layer0_outputs[5042]);
    assign layer1_outputs[412] = (layer0_outputs[1639]) & ~(layer0_outputs[4877]);
    assign layer1_outputs[413] = 1'b0;
    assign layer1_outputs[414] = (layer0_outputs[2417]) & (layer0_outputs[4315]);
    assign layer1_outputs[415] = (layer0_outputs[951]) & ~(layer0_outputs[5084]);
    assign layer1_outputs[416] = ~(layer0_outputs[300]);
    assign layer1_outputs[417] = ~((layer0_outputs[3970]) | (layer0_outputs[1584]));
    assign layer1_outputs[418] = 1'b1;
    assign layer1_outputs[419] = ~(layer0_outputs[3189]) | (layer0_outputs[5073]);
    assign layer1_outputs[420] = ~(layer0_outputs[230]) | (layer0_outputs[3052]);
    assign layer1_outputs[421] = (layer0_outputs[1356]) | (layer0_outputs[2470]);
    assign layer1_outputs[422] = (layer0_outputs[666]) ^ (layer0_outputs[1905]);
    assign layer1_outputs[423] = ~((layer0_outputs[2398]) & (layer0_outputs[1965]));
    assign layer1_outputs[424] = ~((layer0_outputs[1085]) & (layer0_outputs[2519]));
    assign layer1_outputs[425] = ~(layer0_outputs[4191]) | (layer0_outputs[11]);
    assign layer1_outputs[426] = layer0_outputs[4619];
    assign layer1_outputs[427] = 1'b0;
    assign layer1_outputs[428] = layer0_outputs[3569];
    assign layer1_outputs[429] = 1'b0;
    assign layer1_outputs[430] = (layer0_outputs[3232]) & ~(layer0_outputs[1901]);
    assign layer1_outputs[431] = ~(layer0_outputs[1128]) | (layer0_outputs[355]);
    assign layer1_outputs[432] = (layer0_outputs[4295]) & ~(layer0_outputs[3516]);
    assign layer1_outputs[433] = ~((layer0_outputs[509]) & (layer0_outputs[2673]));
    assign layer1_outputs[434] = ~((layer0_outputs[1241]) & (layer0_outputs[2840]));
    assign layer1_outputs[435] = ~(layer0_outputs[3828]);
    assign layer1_outputs[436] = ~((layer0_outputs[1692]) & (layer0_outputs[3689]));
    assign layer1_outputs[437] = (layer0_outputs[3497]) | (layer0_outputs[1428]);
    assign layer1_outputs[438] = ~((layer0_outputs[5083]) ^ (layer0_outputs[4423]));
    assign layer1_outputs[439] = ~((layer0_outputs[184]) & (layer0_outputs[343]));
    assign layer1_outputs[440] = ~(layer0_outputs[4620]);
    assign layer1_outputs[441] = (layer0_outputs[1134]) & ~(layer0_outputs[90]);
    assign layer1_outputs[442] = (layer0_outputs[160]) & ~(layer0_outputs[2948]);
    assign layer1_outputs[443] = (layer0_outputs[290]) & (layer0_outputs[3069]);
    assign layer1_outputs[444] = (layer0_outputs[3674]) & ~(layer0_outputs[5038]);
    assign layer1_outputs[445] = ~((layer0_outputs[791]) ^ (layer0_outputs[1586]));
    assign layer1_outputs[446] = 1'b0;
    assign layer1_outputs[447] = (layer0_outputs[3224]) | (layer0_outputs[3573]);
    assign layer1_outputs[448] = layer0_outputs[1228];
    assign layer1_outputs[449] = ~((layer0_outputs[4354]) & (layer0_outputs[4222]));
    assign layer1_outputs[450] = (layer0_outputs[1187]) | (layer0_outputs[4063]);
    assign layer1_outputs[451] = (layer0_outputs[1023]) & ~(layer0_outputs[4582]);
    assign layer1_outputs[452] = ~((layer0_outputs[2001]) & (layer0_outputs[313]));
    assign layer1_outputs[453] = (layer0_outputs[255]) & ~(layer0_outputs[342]);
    assign layer1_outputs[454] = (layer0_outputs[276]) ^ (layer0_outputs[4792]);
    assign layer1_outputs[455] = (layer0_outputs[3432]) & ~(layer0_outputs[2649]);
    assign layer1_outputs[456] = ~(layer0_outputs[4315]) | (layer0_outputs[1340]);
    assign layer1_outputs[457] = (layer0_outputs[347]) & ~(layer0_outputs[4553]);
    assign layer1_outputs[458] = ~(layer0_outputs[4180]);
    assign layer1_outputs[459] = (layer0_outputs[2285]) & ~(layer0_outputs[1004]);
    assign layer1_outputs[460] = ~((layer0_outputs[1349]) | (layer0_outputs[4456]));
    assign layer1_outputs[461] = ~((layer0_outputs[2383]) & (layer0_outputs[1916]));
    assign layer1_outputs[462] = ~(layer0_outputs[407]);
    assign layer1_outputs[463] = (layer0_outputs[3374]) & ~(layer0_outputs[907]);
    assign layer1_outputs[464] = layer0_outputs[1000];
    assign layer1_outputs[465] = 1'b0;
    assign layer1_outputs[466] = layer0_outputs[4478];
    assign layer1_outputs[467] = (layer0_outputs[2715]) | (layer0_outputs[2703]);
    assign layer1_outputs[468] = ~((layer0_outputs[2742]) & (layer0_outputs[3097]));
    assign layer1_outputs[469] = (layer0_outputs[3412]) & ~(layer0_outputs[4892]);
    assign layer1_outputs[470] = layer0_outputs[4078];
    assign layer1_outputs[471] = ~(layer0_outputs[72]);
    assign layer1_outputs[472] = layer0_outputs[1602];
    assign layer1_outputs[473] = (layer0_outputs[391]) | (layer0_outputs[1492]);
    assign layer1_outputs[474] = ~((layer0_outputs[3275]) | (layer0_outputs[1562]));
    assign layer1_outputs[475] = layer0_outputs[440];
    assign layer1_outputs[476] = layer0_outputs[5018];
    assign layer1_outputs[477] = ~(layer0_outputs[3288]) | (layer0_outputs[3381]);
    assign layer1_outputs[478] = ~(layer0_outputs[4253]);
    assign layer1_outputs[479] = 1'b1;
    assign layer1_outputs[480] = (layer0_outputs[2872]) & ~(layer0_outputs[684]);
    assign layer1_outputs[481] = (layer0_outputs[1165]) & (layer0_outputs[2584]);
    assign layer1_outputs[482] = (layer0_outputs[1899]) & (layer0_outputs[3562]);
    assign layer1_outputs[483] = ~((layer0_outputs[3127]) | (layer0_outputs[4107]));
    assign layer1_outputs[484] = (layer0_outputs[1191]) & (layer0_outputs[4016]);
    assign layer1_outputs[485] = 1'b1;
    assign layer1_outputs[486] = 1'b0;
    assign layer1_outputs[487] = layer0_outputs[1170];
    assign layer1_outputs[488] = 1'b1;
    assign layer1_outputs[489] = (layer0_outputs[3008]) ^ (layer0_outputs[4048]);
    assign layer1_outputs[490] = ~((layer0_outputs[4902]) & (layer0_outputs[1008]));
    assign layer1_outputs[491] = (layer0_outputs[3413]) & ~(layer0_outputs[3316]);
    assign layer1_outputs[492] = (layer0_outputs[3150]) & (layer0_outputs[874]);
    assign layer1_outputs[493] = (layer0_outputs[546]) & (layer0_outputs[2769]);
    assign layer1_outputs[494] = (layer0_outputs[1251]) & ~(layer0_outputs[4252]);
    assign layer1_outputs[495] = ~(layer0_outputs[2975]) | (layer0_outputs[4679]);
    assign layer1_outputs[496] = 1'b1;
    assign layer1_outputs[497] = ~(layer0_outputs[4604]) | (layer0_outputs[2530]);
    assign layer1_outputs[498] = (layer0_outputs[4558]) & (layer0_outputs[2303]);
    assign layer1_outputs[499] = ~(layer0_outputs[2288]) | (layer0_outputs[3904]);
    assign layer1_outputs[500] = ~(layer0_outputs[2727]);
    assign layer1_outputs[501] = ~(layer0_outputs[1109]);
    assign layer1_outputs[502] = ~(layer0_outputs[337]) | (layer0_outputs[3253]);
    assign layer1_outputs[503] = ~(layer0_outputs[1475]) | (layer0_outputs[3014]);
    assign layer1_outputs[504] = 1'b1;
    assign layer1_outputs[505] = 1'b1;
    assign layer1_outputs[506] = 1'b1;
    assign layer1_outputs[507] = ~((layer0_outputs[2014]) | (layer0_outputs[3883]));
    assign layer1_outputs[508] = layer0_outputs[546];
    assign layer1_outputs[509] = ~(layer0_outputs[3784]) | (layer0_outputs[4245]);
    assign layer1_outputs[510] = ~(layer0_outputs[691]) | (layer0_outputs[387]);
    assign layer1_outputs[511] = ~((layer0_outputs[2267]) | (layer0_outputs[2737]));
    assign layer1_outputs[512] = layer0_outputs[386];
    assign layer1_outputs[513] = ~(layer0_outputs[2708]);
    assign layer1_outputs[514] = 1'b0;
    assign layer1_outputs[515] = ~((layer0_outputs[2504]) | (layer0_outputs[4421]));
    assign layer1_outputs[516] = 1'b0;
    assign layer1_outputs[517] = ~(layer0_outputs[4397]);
    assign layer1_outputs[518] = (layer0_outputs[720]) | (layer0_outputs[179]);
    assign layer1_outputs[519] = ~(layer0_outputs[3266]);
    assign layer1_outputs[520] = ~((layer0_outputs[788]) & (layer0_outputs[3172]));
    assign layer1_outputs[521] = 1'b1;
    assign layer1_outputs[522] = ~(layer0_outputs[4581]) | (layer0_outputs[3085]);
    assign layer1_outputs[523] = ~(layer0_outputs[824]);
    assign layer1_outputs[524] = layer0_outputs[492];
    assign layer1_outputs[525] = layer0_outputs[4160];
    assign layer1_outputs[526] = ~((layer0_outputs[2047]) & (layer0_outputs[293]));
    assign layer1_outputs[527] = ~((layer0_outputs[3910]) ^ (layer0_outputs[4796]));
    assign layer1_outputs[528] = 1'b0;
    assign layer1_outputs[529] = layer0_outputs[1959];
    assign layer1_outputs[530] = ~(layer0_outputs[4152]) | (layer0_outputs[1932]);
    assign layer1_outputs[531] = (layer0_outputs[3749]) | (layer0_outputs[2777]);
    assign layer1_outputs[532] = 1'b0;
    assign layer1_outputs[533] = ~(layer0_outputs[760]);
    assign layer1_outputs[534] = layer0_outputs[1577];
    assign layer1_outputs[535] = layer0_outputs[3350];
    assign layer1_outputs[536] = (layer0_outputs[3022]) & ~(layer0_outputs[4787]);
    assign layer1_outputs[537] = ~(layer0_outputs[3287]) | (layer0_outputs[4490]);
    assign layer1_outputs[538] = (layer0_outputs[5044]) & ~(layer0_outputs[568]);
    assign layer1_outputs[539] = ~(layer0_outputs[2751]);
    assign layer1_outputs[540] = layer0_outputs[1652];
    assign layer1_outputs[541] = ~((layer0_outputs[1858]) & (layer0_outputs[4820]));
    assign layer1_outputs[542] = (layer0_outputs[413]) & ~(layer0_outputs[4630]);
    assign layer1_outputs[543] = (layer0_outputs[913]) & ~(layer0_outputs[1017]);
    assign layer1_outputs[544] = (layer0_outputs[873]) | (layer0_outputs[3017]);
    assign layer1_outputs[545] = ~((layer0_outputs[3777]) ^ (layer0_outputs[415]));
    assign layer1_outputs[546] = layer0_outputs[581];
    assign layer1_outputs[547] = (layer0_outputs[1162]) | (layer0_outputs[2690]);
    assign layer1_outputs[548] = ~((layer0_outputs[2550]) | (layer0_outputs[2289]));
    assign layer1_outputs[549] = 1'b0;
    assign layer1_outputs[550] = ~(layer0_outputs[4557]);
    assign layer1_outputs[551] = 1'b0;
    assign layer1_outputs[552] = (layer0_outputs[1079]) & (layer0_outputs[4648]);
    assign layer1_outputs[553] = ~(layer0_outputs[3154]) | (layer0_outputs[3625]);
    assign layer1_outputs[554] = ~(layer0_outputs[4000]) | (layer0_outputs[431]);
    assign layer1_outputs[555] = ~(layer0_outputs[4702]) | (layer0_outputs[2553]);
    assign layer1_outputs[556] = ~((layer0_outputs[1693]) & (layer0_outputs[3499]));
    assign layer1_outputs[557] = (layer0_outputs[57]) & ~(layer0_outputs[2958]);
    assign layer1_outputs[558] = ~((layer0_outputs[1567]) | (layer0_outputs[983]));
    assign layer1_outputs[559] = ~(layer0_outputs[1565]);
    assign layer1_outputs[560] = 1'b0;
    assign layer1_outputs[561] = ~(layer0_outputs[3205]);
    assign layer1_outputs[562] = 1'b0;
    assign layer1_outputs[563] = (layer0_outputs[1373]) & ~(layer0_outputs[242]);
    assign layer1_outputs[564] = 1'b0;
    assign layer1_outputs[565] = 1'b1;
    assign layer1_outputs[566] = 1'b1;
    assign layer1_outputs[567] = ~(layer0_outputs[690]);
    assign layer1_outputs[568] = 1'b1;
    assign layer1_outputs[569] = layer0_outputs[3524];
    assign layer1_outputs[570] = (layer0_outputs[1180]) | (layer0_outputs[1757]);
    assign layer1_outputs[571] = ~(layer0_outputs[3659]) | (layer0_outputs[1845]);
    assign layer1_outputs[572] = ~(layer0_outputs[2435]) | (layer0_outputs[1399]);
    assign layer1_outputs[573] = layer0_outputs[2403];
    assign layer1_outputs[574] = (layer0_outputs[2032]) & ~(layer0_outputs[3383]);
    assign layer1_outputs[575] = (layer0_outputs[3165]) | (layer0_outputs[1690]);
    assign layer1_outputs[576] = 1'b1;
    assign layer1_outputs[577] = layer0_outputs[275];
    assign layer1_outputs[578] = 1'b1;
    assign layer1_outputs[579] = (layer0_outputs[2578]) & (layer0_outputs[2560]);
    assign layer1_outputs[580] = ~(layer0_outputs[1910]);
    assign layer1_outputs[581] = (layer0_outputs[4560]) & ~(layer0_outputs[4866]);
    assign layer1_outputs[582] = ~(layer0_outputs[3934]);
    assign layer1_outputs[583] = ~(layer0_outputs[4389]);
    assign layer1_outputs[584] = (layer0_outputs[18]) & (layer0_outputs[637]);
    assign layer1_outputs[585] = ~(layer0_outputs[3736]);
    assign layer1_outputs[586] = ~(layer0_outputs[986]);
    assign layer1_outputs[587] = (layer0_outputs[4402]) | (layer0_outputs[1091]);
    assign layer1_outputs[588] = (layer0_outputs[1697]) & ~(layer0_outputs[1698]);
    assign layer1_outputs[589] = ~(layer0_outputs[1054]) | (layer0_outputs[1658]);
    assign layer1_outputs[590] = ~(layer0_outputs[3854]);
    assign layer1_outputs[591] = 1'b1;
    assign layer1_outputs[592] = layer0_outputs[983];
    assign layer1_outputs[593] = ~((layer0_outputs[573]) & (layer0_outputs[344]));
    assign layer1_outputs[594] = layer0_outputs[3038];
    assign layer1_outputs[595] = ~(layer0_outputs[4323]) | (layer0_outputs[4545]);
    assign layer1_outputs[596] = 1'b0;
    assign layer1_outputs[597] = ~(layer0_outputs[964]) | (layer0_outputs[3787]);
    assign layer1_outputs[598] = ~(layer0_outputs[3478]) | (layer0_outputs[3334]);
    assign layer1_outputs[599] = ~(layer0_outputs[3213]) | (layer0_outputs[4380]);
    assign layer1_outputs[600] = (layer0_outputs[61]) & (layer0_outputs[741]);
    assign layer1_outputs[601] = layer0_outputs[3823];
    assign layer1_outputs[602] = 1'b0;
    assign layer1_outputs[603] = layer0_outputs[3277];
    assign layer1_outputs[604] = 1'b0;
    assign layer1_outputs[605] = ~(layer0_outputs[4116]);
    assign layer1_outputs[606] = (layer0_outputs[3354]) & ~(layer0_outputs[3875]);
    assign layer1_outputs[607] = 1'b0;
    assign layer1_outputs[608] = ~(layer0_outputs[3386]) | (layer0_outputs[5030]);
    assign layer1_outputs[609] = ~(layer0_outputs[741]);
    assign layer1_outputs[610] = (layer0_outputs[3865]) & ~(layer0_outputs[1032]);
    assign layer1_outputs[611] = (layer0_outputs[2582]) & (layer0_outputs[3842]);
    assign layer1_outputs[612] = ~(layer0_outputs[3684]);
    assign layer1_outputs[613] = ~((layer0_outputs[1957]) | (layer0_outputs[3333]));
    assign layer1_outputs[614] = ~((layer0_outputs[4720]) | (layer0_outputs[2229]));
    assign layer1_outputs[615] = (layer0_outputs[1399]) & ~(layer0_outputs[4568]);
    assign layer1_outputs[616] = 1'b0;
    assign layer1_outputs[617] = (layer0_outputs[369]) ^ (layer0_outputs[4748]);
    assign layer1_outputs[618] = ~(layer0_outputs[2818]) | (layer0_outputs[2998]);
    assign layer1_outputs[619] = (layer0_outputs[1738]) & ~(layer0_outputs[2341]);
    assign layer1_outputs[620] = layer0_outputs[2844];
    assign layer1_outputs[621] = ~(layer0_outputs[4554]);
    assign layer1_outputs[622] = ~((layer0_outputs[1270]) & (layer0_outputs[701]));
    assign layer1_outputs[623] = layer0_outputs[1057];
    assign layer1_outputs[624] = (layer0_outputs[2500]) | (layer0_outputs[4794]);
    assign layer1_outputs[625] = 1'b1;
    assign layer1_outputs[626] = (layer0_outputs[748]) & ~(layer0_outputs[4834]);
    assign layer1_outputs[627] = ~((layer0_outputs[4944]) ^ (layer0_outputs[256]));
    assign layer1_outputs[628] = ~(layer0_outputs[4392]);
    assign layer1_outputs[629] = 1'b1;
    assign layer1_outputs[630] = ~(layer0_outputs[3113]) | (layer0_outputs[3860]);
    assign layer1_outputs[631] = 1'b1;
    assign layer1_outputs[632] = (layer0_outputs[4806]) & (layer0_outputs[2526]);
    assign layer1_outputs[633] = ~(layer0_outputs[204]);
    assign layer1_outputs[634] = ~(layer0_outputs[2555]);
    assign layer1_outputs[635] = 1'b1;
    assign layer1_outputs[636] = ~(layer0_outputs[3357]);
    assign layer1_outputs[637] = (layer0_outputs[2101]) & (layer0_outputs[4046]);
    assign layer1_outputs[638] = 1'b1;
    assign layer1_outputs[639] = layer0_outputs[3031];
    assign layer1_outputs[640] = ~(layer0_outputs[3027]);
    assign layer1_outputs[641] = ~(layer0_outputs[2789]);
    assign layer1_outputs[642] = 1'b0;
    assign layer1_outputs[643] = 1'b1;
    assign layer1_outputs[644] = ~((layer0_outputs[3564]) & (layer0_outputs[913]));
    assign layer1_outputs[645] = 1'b1;
    assign layer1_outputs[646] = (layer0_outputs[3869]) & (layer0_outputs[4863]);
    assign layer1_outputs[647] = 1'b0;
    assign layer1_outputs[648] = ~(layer0_outputs[4093]) | (layer0_outputs[2861]);
    assign layer1_outputs[649] = 1'b0;
    assign layer1_outputs[650] = ~(layer0_outputs[4963]);
    assign layer1_outputs[651] = layer0_outputs[3917];
    assign layer1_outputs[652] = (layer0_outputs[3822]) & ~(layer0_outputs[748]);
    assign layer1_outputs[653] = (layer0_outputs[1321]) | (layer0_outputs[4777]);
    assign layer1_outputs[654] = ~(layer0_outputs[4406]);
    assign layer1_outputs[655] = ~((layer0_outputs[189]) | (layer0_outputs[4135]));
    assign layer1_outputs[656] = (layer0_outputs[4403]) | (layer0_outputs[4386]);
    assign layer1_outputs[657] = ~(layer0_outputs[1804]) | (layer0_outputs[3554]);
    assign layer1_outputs[658] = 1'b0;
    assign layer1_outputs[659] = layer0_outputs[3935];
    assign layer1_outputs[660] = ~((layer0_outputs[1546]) & (layer0_outputs[268]));
    assign layer1_outputs[661] = (layer0_outputs[914]) & (layer0_outputs[4776]);
    assign layer1_outputs[662] = ~(layer0_outputs[1530]);
    assign layer1_outputs[663] = (layer0_outputs[1454]) | (layer0_outputs[4687]);
    assign layer1_outputs[664] = ~((layer0_outputs[665]) & (layer0_outputs[4524]));
    assign layer1_outputs[665] = (layer0_outputs[1047]) ^ (layer0_outputs[636]);
    assign layer1_outputs[666] = (layer0_outputs[2152]) & (layer0_outputs[1489]);
    assign layer1_outputs[667] = layer0_outputs[1254];
    assign layer1_outputs[668] = ~((layer0_outputs[5093]) & (layer0_outputs[1038]));
    assign layer1_outputs[669] = (layer0_outputs[4023]) | (layer0_outputs[686]);
    assign layer1_outputs[670] = layer0_outputs[1664];
    assign layer1_outputs[671] = ~(layer0_outputs[3742]) | (layer0_outputs[2940]);
    assign layer1_outputs[672] = ~(layer0_outputs[1276]);
    assign layer1_outputs[673] = (layer0_outputs[4966]) & (layer0_outputs[987]);
    assign layer1_outputs[674] = 1'b1;
    assign layer1_outputs[675] = (layer0_outputs[4071]) & (layer0_outputs[919]);
    assign layer1_outputs[676] = ~((layer0_outputs[4151]) | (layer0_outputs[4871]));
    assign layer1_outputs[677] = ~(layer0_outputs[4606]) | (layer0_outputs[2512]);
    assign layer1_outputs[678] = (layer0_outputs[1720]) & ~(layer0_outputs[3253]);
    assign layer1_outputs[679] = ~(layer0_outputs[2660]) | (layer0_outputs[2905]);
    assign layer1_outputs[680] = ~(layer0_outputs[3861]);
    assign layer1_outputs[681] = ~((layer0_outputs[2937]) ^ (layer0_outputs[4498]));
    assign layer1_outputs[682] = ~((layer0_outputs[1312]) & (layer0_outputs[2760]));
    assign layer1_outputs[683] = 1'b1;
    assign layer1_outputs[684] = ~((layer0_outputs[3048]) & (layer0_outputs[2976]));
    assign layer1_outputs[685] = layer0_outputs[4084];
    assign layer1_outputs[686] = layer0_outputs[3026];
    assign layer1_outputs[687] = ~((layer0_outputs[2421]) | (layer0_outputs[2608]));
    assign layer1_outputs[688] = ~((layer0_outputs[3368]) ^ (layer0_outputs[3439]));
    assign layer1_outputs[689] = (layer0_outputs[188]) | (layer0_outputs[705]);
    assign layer1_outputs[690] = ~(layer0_outputs[1280]) | (layer0_outputs[2706]);
    assign layer1_outputs[691] = (layer0_outputs[1403]) & ~(layer0_outputs[701]);
    assign layer1_outputs[692] = layer0_outputs[1319];
    assign layer1_outputs[693] = ~(layer0_outputs[3794]);
    assign layer1_outputs[694] = layer0_outputs[4821];
    assign layer1_outputs[695] = (layer0_outputs[1602]) ^ (layer0_outputs[2020]);
    assign layer1_outputs[696] = (layer0_outputs[5013]) | (layer0_outputs[380]);
    assign layer1_outputs[697] = 1'b1;
    assign layer1_outputs[698] = (layer0_outputs[1060]) & (layer0_outputs[3788]);
    assign layer1_outputs[699] = (layer0_outputs[578]) | (layer0_outputs[2638]);
    assign layer1_outputs[700] = 1'b0;
    assign layer1_outputs[701] = 1'b1;
    assign layer1_outputs[702] = (layer0_outputs[89]) & (layer0_outputs[3236]);
    assign layer1_outputs[703] = 1'b0;
    assign layer1_outputs[704] = 1'b0;
    assign layer1_outputs[705] = ~((layer0_outputs[639]) ^ (layer0_outputs[2253]));
    assign layer1_outputs[706] = 1'b0;
    assign layer1_outputs[707] = ~(layer0_outputs[992]) | (layer0_outputs[4365]);
    assign layer1_outputs[708] = ~(layer0_outputs[4931]) | (layer0_outputs[2747]);
    assign layer1_outputs[709] = (layer0_outputs[205]) & ~(layer0_outputs[4060]);
    assign layer1_outputs[710] = (layer0_outputs[2894]) & (layer0_outputs[4647]);
    assign layer1_outputs[711] = (layer0_outputs[4695]) & ~(layer0_outputs[4130]);
    assign layer1_outputs[712] = 1'b0;
    assign layer1_outputs[713] = (layer0_outputs[3833]) & ~(layer0_outputs[3790]);
    assign layer1_outputs[714] = ~((layer0_outputs[5106]) ^ (layer0_outputs[4602]));
    assign layer1_outputs[715] = ~(layer0_outputs[4928]) | (layer0_outputs[3464]);
    assign layer1_outputs[716] = ~((layer0_outputs[3944]) & (layer0_outputs[308]));
    assign layer1_outputs[717] = ~((layer0_outputs[3590]) | (layer0_outputs[1348]));
    assign layer1_outputs[718] = ~(layer0_outputs[1398]) | (layer0_outputs[2747]);
    assign layer1_outputs[719] = ~((layer0_outputs[4648]) ^ (layer0_outputs[3370]));
    assign layer1_outputs[720] = (layer0_outputs[3158]) & (layer0_outputs[3786]);
    assign layer1_outputs[721] = ~(layer0_outputs[5104]);
    assign layer1_outputs[722] = 1'b1;
    assign layer1_outputs[723] = ~(layer0_outputs[4120]) | (layer0_outputs[643]);
    assign layer1_outputs[724] = 1'b0;
    assign layer1_outputs[725] = ~((layer0_outputs[811]) & (layer0_outputs[4939]));
    assign layer1_outputs[726] = ~(layer0_outputs[4438]) | (layer0_outputs[4215]);
    assign layer1_outputs[727] = (layer0_outputs[1897]) ^ (layer0_outputs[1355]);
    assign layer1_outputs[728] = (layer0_outputs[3095]) & (layer0_outputs[1419]);
    assign layer1_outputs[729] = (layer0_outputs[4845]) & ~(layer0_outputs[1537]);
    assign layer1_outputs[730] = ~((layer0_outputs[4983]) & (layer0_outputs[2535]));
    assign layer1_outputs[731] = ~(layer0_outputs[1642]);
    assign layer1_outputs[732] = ~(layer0_outputs[1869]) | (layer0_outputs[3765]);
    assign layer1_outputs[733] = (layer0_outputs[5107]) & (layer0_outputs[4022]);
    assign layer1_outputs[734] = ~((layer0_outputs[3038]) ^ (layer0_outputs[309]));
    assign layer1_outputs[735] = 1'b1;
    assign layer1_outputs[736] = ~((layer0_outputs[4476]) & (layer0_outputs[1203]));
    assign layer1_outputs[737] = ~(layer0_outputs[479]) | (layer0_outputs[763]);
    assign layer1_outputs[738] = (layer0_outputs[1201]) ^ (layer0_outputs[1113]);
    assign layer1_outputs[739] = (layer0_outputs[5001]) & ~(layer0_outputs[3951]);
    assign layer1_outputs[740] = ~((layer0_outputs[2084]) | (layer0_outputs[3011]));
    assign layer1_outputs[741] = ~((layer0_outputs[3232]) & (layer0_outputs[2585]));
    assign layer1_outputs[742] = (layer0_outputs[316]) & ~(layer0_outputs[245]);
    assign layer1_outputs[743] = (layer0_outputs[2564]) & (layer0_outputs[442]);
    assign layer1_outputs[744] = (layer0_outputs[379]) ^ (layer0_outputs[3715]);
    assign layer1_outputs[745] = ~(layer0_outputs[2746]);
    assign layer1_outputs[746] = layer0_outputs[224];
    assign layer1_outputs[747] = ~((layer0_outputs[1904]) ^ (layer0_outputs[4902]));
    assign layer1_outputs[748] = (layer0_outputs[563]) & ~(layer0_outputs[4245]);
    assign layer1_outputs[749] = (layer0_outputs[1235]) & ~(layer0_outputs[715]);
    assign layer1_outputs[750] = 1'b0;
    assign layer1_outputs[751] = 1'b0;
    assign layer1_outputs[752] = (layer0_outputs[3273]) & ~(layer0_outputs[2712]);
    assign layer1_outputs[753] = ~(layer0_outputs[3556]);
    assign layer1_outputs[754] = ~(layer0_outputs[4065]);
    assign layer1_outputs[755] = layer0_outputs[2599];
    assign layer1_outputs[756] = ~((layer0_outputs[2445]) | (layer0_outputs[5003]));
    assign layer1_outputs[757] = (layer0_outputs[4743]) & ~(layer0_outputs[3905]);
    assign layer1_outputs[758] = (layer0_outputs[2141]) & ~(layer0_outputs[1729]);
    assign layer1_outputs[759] = ~(layer0_outputs[2391]) | (layer0_outputs[3212]);
    assign layer1_outputs[760] = (layer0_outputs[4763]) | (layer0_outputs[5071]);
    assign layer1_outputs[761] = (layer0_outputs[3932]) & ~(layer0_outputs[1337]);
    assign layer1_outputs[762] = ~(layer0_outputs[1458]) | (layer0_outputs[480]);
    assign layer1_outputs[763] = 1'b1;
    assign layer1_outputs[764] = 1'b1;
    assign layer1_outputs[765] = ~(layer0_outputs[1440]) | (layer0_outputs[4016]);
    assign layer1_outputs[766] = ~((layer0_outputs[4244]) & (layer0_outputs[4732]));
    assign layer1_outputs[767] = layer0_outputs[2461];
    assign layer1_outputs[768] = (layer0_outputs[3396]) & (layer0_outputs[1020]);
    assign layer1_outputs[769] = ~((layer0_outputs[912]) & (layer0_outputs[4917]));
    assign layer1_outputs[770] = (layer0_outputs[407]) & ~(layer0_outputs[4069]);
    assign layer1_outputs[771] = (layer0_outputs[2254]) & ~(layer0_outputs[2471]);
    assign layer1_outputs[772] = (layer0_outputs[3991]) & ~(layer0_outputs[4122]);
    assign layer1_outputs[773] = ~(layer0_outputs[979]);
    assign layer1_outputs[774] = ~(layer0_outputs[5016]);
    assign layer1_outputs[775] = ~((layer0_outputs[2558]) & (layer0_outputs[325]));
    assign layer1_outputs[776] = ~((layer0_outputs[4002]) & (layer0_outputs[2545]));
    assign layer1_outputs[777] = (layer0_outputs[5077]) & (layer0_outputs[198]);
    assign layer1_outputs[778] = 1'b1;
    assign layer1_outputs[779] = (layer0_outputs[4962]) & ~(layer0_outputs[1947]);
    assign layer1_outputs[780] = ~(layer0_outputs[4074]);
    assign layer1_outputs[781] = 1'b0;
    assign layer1_outputs[782] = (layer0_outputs[3153]) & ~(layer0_outputs[519]);
    assign layer1_outputs[783] = (layer0_outputs[550]) ^ (layer0_outputs[570]);
    assign layer1_outputs[784] = ~(layer0_outputs[3257]);
    assign layer1_outputs[785] = (layer0_outputs[522]) ^ (layer0_outputs[4064]);
    assign layer1_outputs[786] = layer0_outputs[3886];
    assign layer1_outputs[787] = ~((layer0_outputs[4374]) & (layer0_outputs[3098]));
    assign layer1_outputs[788] = 1'b1;
    assign layer1_outputs[789] = layer0_outputs[1500];
    assign layer1_outputs[790] = ~(layer0_outputs[594]) | (layer0_outputs[405]);
    assign layer1_outputs[791] = layer0_outputs[611];
    assign layer1_outputs[792] = 1'b0;
    assign layer1_outputs[793] = layer0_outputs[398];
    assign layer1_outputs[794] = ~((layer0_outputs[2966]) | (layer0_outputs[4990]));
    assign layer1_outputs[795] = ~(layer0_outputs[999]) | (layer0_outputs[4901]);
    assign layer1_outputs[796] = layer0_outputs[4292];
    assign layer1_outputs[797] = (layer0_outputs[4930]) | (layer0_outputs[1368]);
    assign layer1_outputs[798] = layer0_outputs[642];
    assign layer1_outputs[799] = (layer0_outputs[1257]) & ~(layer0_outputs[3326]);
    assign layer1_outputs[800] = (layer0_outputs[1909]) | (layer0_outputs[1708]);
    assign layer1_outputs[801] = ~((layer0_outputs[4387]) | (layer0_outputs[1553]));
    assign layer1_outputs[802] = (layer0_outputs[150]) & ~(layer0_outputs[1000]);
    assign layer1_outputs[803] = ~(layer0_outputs[3451]);
    assign layer1_outputs[804] = ~(layer0_outputs[33]) | (layer0_outputs[1500]);
    assign layer1_outputs[805] = 1'b0;
    assign layer1_outputs[806] = layer0_outputs[5043];
    assign layer1_outputs[807] = layer0_outputs[2356];
    assign layer1_outputs[808] = ~(layer0_outputs[2870]);
    assign layer1_outputs[809] = 1'b0;
    assign layer1_outputs[810] = ~(layer0_outputs[2903]);
    assign layer1_outputs[811] = (layer0_outputs[992]) | (layer0_outputs[139]);
    assign layer1_outputs[812] = layer0_outputs[2171];
    assign layer1_outputs[813] = ~((layer0_outputs[1615]) & (layer0_outputs[849]));
    assign layer1_outputs[814] = layer0_outputs[4252];
    assign layer1_outputs[815] = 1'b1;
    assign layer1_outputs[816] = ~((layer0_outputs[3308]) & (layer0_outputs[4967]));
    assign layer1_outputs[817] = ~((layer0_outputs[1372]) | (layer0_outputs[5069]));
    assign layer1_outputs[818] = ~(layer0_outputs[2594]);
    assign layer1_outputs[819] = layer0_outputs[1103];
    assign layer1_outputs[820] = (layer0_outputs[2218]) & ~(layer0_outputs[2933]);
    assign layer1_outputs[821] = (layer0_outputs[1467]) ^ (layer0_outputs[1652]);
    assign layer1_outputs[822] = ~(layer0_outputs[4951]);
    assign layer1_outputs[823] = 1'b1;
    assign layer1_outputs[824] = (layer0_outputs[2797]) ^ (layer0_outputs[2829]);
    assign layer1_outputs[825] = ~(layer0_outputs[1223]) | (layer0_outputs[4843]);
    assign layer1_outputs[826] = ~(layer0_outputs[3941]);
    assign layer1_outputs[827] = (layer0_outputs[4368]) & ~(layer0_outputs[2455]);
    assign layer1_outputs[828] = ~(layer0_outputs[384]);
    assign layer1_outputs[829] = ~(layer0_outputs[840]) | (layer0_outputs[1552]);
    assign layer1_outputs[830] = ~((layer0_outputs[2713]) & (layer0_outputs[4413]));
    assign layer1_outputs[831] = ~(layer0_outputs[3188]) | (layer0_outputs[182]);
    assign layer1_outputs[832] = ~(layer0_outputs[888]) | (layer0_outputs[4621]);
    assign layer1_outputs[833] = layer0_outputs[2786];
    assign layer1_outputs[834] = 1'b1;
    assign layer1_outputs[835] = layer0_outputs[205];
    assign layer1_outputs[836] = 1'b0;
    assign layer1_outputs[837] = ~((layer0_outputs[1753]) & (layer0_outputs[4788]));
    assign layer1_outputs[838] = layer0_outputs[2820];
    assign layer1_outputs[839] = (layer0_outputs[1171]) & ~(layer0_outputs[1702]);
    assign layer1_outputs[840] = ~(layer0_outputs[4118]);
    assign layer1_outputs[841] = ~(layer0_outputs[4253]);
    assign layer1_outputs[842] = (layer0_outputs[1926]) & (layer0_outputs[1799]);
    assign layer1_outputs[843] = ~(layer0_outputs[2768]) | (layer0_outputs[2541]);
    assign layer1_outputs[844] = (layer0_outputs[4973]) & ~(layer0_outputs[1434]);
    assign layer1_outputs[845] = (layer0_outputs[3505]) & ~(layer0_outputs[367]);
    assign layer1_outputs[846] = ~((layer0_outputs[3682]) | (layer0_outputs[1646]));
    assign layer1_outputs[847] = layer0_outputs[4864];
    assign layer1_outputs[848] = layer0_outputs[3223];
    assign layer1_outputs[849] = 1'b0;
    assign layer1_outputs[850] = layer0_outputs[1326];
    assign layer1_outputs[851] = (layer0_outputs[3200]) & ~(layer0_outputs[1965]);
    assign layer1_outputs[852] = 1'b0;
    assign layer1_outputs[853] = 1'b0;
    assign layer1_outputs[854] = ~((layer0_outputs[1343]) ^ (layer0_outputs[3105]));
    assign layer1_outputs[855] = ~((layer0_outputs[1484]) | (layer0_outputs[900]));
    assign layer1_outputs[856] = (layer0_outputs[4349]) | (layer0_outputs[2016]);
    assign layer1_outputs[857] = ~(layer0_outputs[4916]);
    assign layer1_outputs[858] = (layer0_outputs[1206]) | (layer0_outputs[3414]);
    assign layer1_outputs[859] = ~((layer0_outputs[4146]) ^ (layer0_outputs[1974]));
    assign layer1_outputs[860] = 1'b0;
    assign layer1_outputs[861] = 1'b1;
    assign layer1_outputs[862] = 1'b0;
    assign layer1_outputs[863] = layer0_outputs[1234];
    assign layer1_outputs[864] = ~(layer0_outputs[1932]) | (layer0_outputs[2179]);
    assign layer1_outputs[865] = layer0_outputs[3620];
    assign layer1_outputs[866] = 1'b0;
    assign layer1_outputs[867] = 1'b1;
    assign layer1_outputs[868] = 1'b1;
    assign layer1_outputs[869] = 1'b0;
    assign layer1_outputs[870] = layer0_outputs[3683];
    assign layer1_outputs[871] = ~(layer0_outputs[2349]) | (layer0_outputs[2351]);
    assign layer1_outputs[872] = 1'b0;
    assign layer1_outputs[873] = ~(layer0_outputs[1883]) | (layer0_outputs[2172]);
    assign layer1_outputs[874] = (layer0_outputs[2441]) & ~(layer0_outputs[3087]);
    assign layer1_outputs[875] = (layer0_outputs[48]) ^ (layer0_outputs[4984]);
    assign layer1_outputs[876] = ~(layer0_outputs[1393]);
    assign layer1_outputs[877] = (layer0_outputs[4311]) & ~(layer0_outputs[4132]);
    assign layer1_outputs[878] = 1'b1;
    assign layer1_outputs[879] = (layer0_outputs[1798]) & (layer0_outputs[3002]);
    assign layer1_outputs[880] = ~((layer0_outputs[3609]) & (layer0_outputs[4126]));
    assign layer1_outputs[881] = layer0_outputs[1753];
    assign layer1_outputs[882] = ~((layer0_outputs[2131]) | (layer0_outputs[3691]));
    assign layer1_outputs[883] = layer0_outputs[4526];
    assign layer1_outputs[884] = ~(layer0_outputs[299]);
    assign layer1_outputs[885] = ~(layer0_outputs[3520]) | (layer0_outputs[4479]);
    assign layer1_outputs[886] = layer0_outputs[1836];
    assign layer1_outputs[887] = layer0_outputs[1425];
    assign layer1_outputs[888] = (layer0_outputs[2125]) | (layer0_outputs[4331]);
    assign layer1_outputs[889] = (layer0_outputs[816]) & (layer0_outputs[4832]);
    assign layer1_outputs[890] = ~(layer0_outputs[4338]);
    assign layer1_outputs[891] = layer0_outputs[2805];
    assign layer1_outputs[892] = layer0_outputs[2751];
    assign layer1_outputs[893] = layer0_outputs[4917];
    assign layer1_outputs[894] = ~((layer0_outputs[3435]) | (layer0_outputs[764]));
    assign layer1_outputs[895] = ~(layer0_outputs[3330]) | (layer0_outputs[322]);
    assign layer1_outputs[896] = 1'b0;
    assign layer1_outputs[897] = ~((layer0_outputs[1948]) & (layer0_outputs[1885]));
    assign layer1_outputs[898] = 1'b0;
    assign layer1_outputs[899] = ~(layer0_outputs[4534]);
    assign layer1_outputs[900] = (layer0_outputs[4590]) & ~(layer0_outputs[3344]);
    assign layer1_outputs[901] = 1'b1;
    assign layer1_outputs[902] = (layer0_outputs[4956]) ^ (layer0_outputs[534]);
    assign layer1_outputs[903] = (layer0_outputs[3166]) | (layer0_outputs[4494]);
    assign layer1_outputs[904] = 1'b0;
    assign layer1_outputs[905] = 1'b0;
    assign layer1_outputs[906] = (layer0_outputs[921]) & ~(layer0_outputs[3574]);
    assign layer1_outputs[907] = ~(layer0_outputs[3628]);
    assign layer1_outputs[908] = ~((layer0_outputs[3084]) | (layer0_outputs[537]));
    assign layer1_outputs[909] = ~(layer0_outputs[4206]) | (layer0_outputs[1510]);
    assign layer1_outputs[910] = (layer0_outputs[942]) | (layer0_outputs[4864]);
    assign layer1_outputs[911] = (layer0_outputs[4504]) & ~(layer0_outputs[2812]);
    assign layer1_outputs[912] = layer0_outputs[3945];
    assign layer1_outputs[913] = 1'b1;
    assign layer1_outputs[914] = ~((layer0_outputs[520]) & (layer0_outputs[868]));
    assign layer1_outputs[915] = (layer0_outputs[4996]) & ~(layer0_outputs[2225]);
    assign layer1_outputs[916] = ~(layer0_outputs[982]);
    assign layer1_outputs[917] = ~((layer0_outputs[362]) ^ (layer0_outputs[4745]));
    assign layer1_outputs[918] = 1'b1;
    assign layer1_outputs[919] = (layer0_outputs[4264]) & ~(layer0_outputs[1332]);
    assign layer1_outputs[920] = ~(layer0_outputs[3630]);
    assign layer1_outputs[921] = ~(layer0_outputs[4955]) | (layer0_outputs[447]);
    assign layer1_outputs[922] = ~((layer0_outputs[3239]) & (layer0_outputs[1649]));
    assign layer1_outputs[923] = (layer0_outputs[1269]) & ~(layer0_outputs[1205]);
    assign layer1_outputs[924] = 1'b0;
    assign layer1_outputs[925] = (layer0_outputs[3598]) | (layer0_outputs[2015]);
    assign layer1_outputs[926] = 1'b1;
    assign layer1_outputs[927] = layer0_outputs[3144];
    assign layer1_outputs[928] = (layer0_outputs[2824]) & (layer0_outputs[1191]);
    assign layer1_outputs[929] = (layer0_outputs[488]) & ~(layer0_outputs[143]);
    assign layer1_outputs[930] = ~(layer0_outputs[2938]);
    assign layer1_outputs[931] = ~((layer0_outputs[1580]) | (layer0_outputs[3072]));
    assign layer1_outputs[932] = ~(layer0_outputs[1588]);
    assign layer1_outputs[933] = (layer0_outputs[1634]) & ~(layer0_outputs[3140]);
    assign layer1_outputs[934] = (layer0_outputs[5051]) & ~(layer0_outputs[3204]);
    assign layer1_outputs[935] = (layer0_outputs[4136]) & ~(layer0_outputs[1710]);
    assign layer1_outputs[936] = 1'b0;
    assign layer1_outputs[937] = ~(layer0_outputs[4409]);
    assign layer1_outputs[938] = ~(layer0_outputs[4542]);
    assign layer1_outputs[939] = ~(layer0_outputs[1994]) | (layer0_outputs[71]);
    assign layer1_outputs[940] = ~((layer0_outputs[2625]) & (layer0_outputs[1898]));
    assign layer1_outputs[941] = (layer0_outputs[2518]) | (layer0_outputs[1138]);
    assign layer1_outputs[942] = layer0_outputs[2139];
    assign layer1_outputs[943] = ~((layer0_outputs[3906]) | (layer0_outputs[2286]));
    assign layer1_outputs[944] = (layer0_outputs[901]) & (layer0_outputs[2587]);
    assign layer1_outputs[945] = (layer0_outputs[1616]) & ~(layer0_outputs[930]);
    assign layer1_outputs[946] = ~((layer0_outputs[4370]) | (layer0_outputs[4660]));
    assign layer1_outputs[947] = ~(layer0_outputs[1307]) | (layer0_outputs[4371]);
    assign layer1_outputs[948] = ~(layer0_outputs[2561]) | (layer0_outputs[1973]);
    assign layer1_outputs[949] = (layer0_outputs[4827]) ^ (layer0_outputs[2544]);
    assign layer1_outputs[950] = ~((layer0_outputs[3489]) | (layer0_outputs[4762]));
    assign layer1_outputs[951] = (layer0_outputs[2182]) | (layer0_outputs[1819]);
    assign layer1_outputs[952] = (layer0_outputs[2672]) & (layer0_outputs[1525]);
    assign layer1_outputs[953] = layer0_outputs[2006];
    assign layer1_outputs[954] = (layer0_outputs[1055]) & ~(layer0_outputs[101]);
    assign layer1_outputs[955] = ~(layer0_outputs[2092]);
    assign layer1_outputs[956] = ~((layer0_outputs[521]) ^ (layer0_outputs[5031]));
    assign layer1_outputs[957] = 1'b0;
    assign layer1_outputs[958] = (layer0_outputs[1155]) & ~(layer0_outputs[1984]);
    assign layer1_outputs[959] = layer0_outputs[1252];
    assign layer1_outputs[960] = ~(layer0_outputs[2085]) | (layer0_outputs[4099]);
    assign layer1_outputs[961] = ~(layer0_outputs[1738]) | (layer0_outputs[737]);
    assign layer1_outputs[962] = 1'b0;
    assign layer1_outputs[963] = ~((layer0_outputs[1585]) & (layer0_outputs[4473]));
    assign layer1_outputs[964] = (layer0_outputs[4629]) & ~(layer0_outputs[884]);
    assign layer1_outputs[965] = (layer0_outputs[4387]) | (layer0_outputs[2292]);
    assign layer1_outputs[966] = (layer0_outputs[81]) & ~(layer0_outputs[3150]);
    assign layer1_outputs[967] = (layer0_outputs[3853]) & (layer0_outputs[1106]);
    assign layer1_outputs[968] = (layer0_outputs[2740]) & (layer0_outputs[119]);
    assign layer1_outputs[969] = ~(layer0_outputs[4189]);
    assign layer1_outputs[970] = ~(layer0_outputs[4491]);
    assign layer1_outputs[971] = 1'b0;
    assign layer1_outputs[972] = layer0_outputs[3419];
    assign layer1_outputs[973] = ~((layer0_outputs[1478]) & (layer0_outputs[4868]));
    assign layer1_outputs[974] = ~(layer0_outputs[4860]);
    assign layer1_outputs[975] = ~((layer0_outputs[3740]) | (layer0_outputs[4785]));
    assign layer1_outputs[976] = ~((layer0_outputs[1468]) | (layer0_outputs[984]));
    assign layer1_outputs[977] = 1'b1;
    assign layer1_outputs[978] = ~(layer0_outputs[912]);
    assign layer1_outputs[979] = layer0_outputs[144];
    assign layer1_outputs[980] = (layer0_outputs[4410]) | (layer0_outputs[3205]);
    assign layer1_outputs[981] = (layer0_outputs[4225]) & ~(layer0_outputs[4265]);
    assign layer1_outputs[982] = ~(layer0_outputs[1601]) | (layer0_outputs[825]);
    assign layer1_outputs[983] = layer0_outputs[4463];
    assign layer1_outputs[984] = (layer0_outputs[1969]) & ~(layer0_outputs[812]);
    assign layer1_outputs[985] = ~(layer0_outputs[2038]);
    assign layer1_outputs[986] = ~(layer0_outputs[814]);
    assign layer1_outputs[987] = layer0_outputs[4459];
    assign layer1_outputs[988] = layer0_outputs[2539];
    assign layer1_outputs[989] = (layer0_outputs[2401]) & ~(layer0_outputs[3291]);
    assign layer1_outputs[990] = layer0_outputs[1242];
    assign layer1_outputs[991] = ~(layer0_outputs[3051]) | (layer0_outputs[2220]);
    assign layer1_outputs[992] = ~(layer0_outputs[2798]);
    assign layer1_outputs[993] = ~((layer0_outputs[317]) & (layer0_outputs[2611]));
    assign layer1_outputs[994] = layer0_outputs[4601];
    assign layer1_outputs[995] = ~((layer0_outputs[4847]) | (layer0_outputs[4924]));
    assign layer1_outputs[996] = (layer0_outputs[4482]) & ~(layer0_outputs[330]);
    assign layer1_outputs[997] = (layer0_outputs[2447]) & ~(layer0_outputs[1968]);
    assign layer1_outputs[998] = ~(layer0_outputs[2839]) | (layer0_outputs[2682]);
    assign layer1_outputs[999] = (layer0_outputs[2217]) & ~(layer0_outputs[2236]);
    assign layer1_outputs[1000] = ~(layer0_outputs[1843]) | (layer0_outputs[2070]);
    assign layer1_outputs[1001] = (layer0_outputs[431]) | (layer0_outputs[2542]);
    assign layer1_outputs[1002] = 1'b0;
    assign layer1_outputs[1003] = ~((layer0_outputs[4964]) & (layer0_outputs[2177]));
    assign layer1_outputs[1004] = ~(layer0_outputs[4919]) | (layer0_outputs[4081]);
    assign layer1_outputs[1005] = ~(layer0_outputs[2924]);
    assign layer1_outputs[1006] = 1'b0;
    assign layer1_outputs[1007] = ~(layer0_outputs[1927]);
    assign layer1_outputs[1008] = ~(layer0_outputs[1143]) | (layer0_outputs[1220]);
    assign layer1_outputs[1009] = ~((layer0_outputs[4384]) & (layer0_outputs[222]));
    assign layer1_outputs[1010] = (layer0_outputs[4101]) & ~(layer0_outputs[979]);
    assign layer1_outputs[1011] = 1'b1;
    assign layer1_outputs[1012] = ~((layer0_outputs[1094]) | (layer0_outputs[2907]));
    assign layer1_outputs[1013] = (layer0_outputs[429]) & ~(layer0_outputs[2883]);
    assign layer1_outputs[1014] = ~((layer0_outputs[215]) | (layer0_outputs[4608]));
    assign layer1_outputs[1015] = ~(layer0_outputs[5110]);
    assign layer1_outputs[1016] = layer0_outputs[412];
    assign layer1_outputs[1017] = (layer0_outputs[3368]) | (layer0_outputs[1587]);
    assign layer1_outputs[1018] = ~((layer0_outputs[4415]) ^ (layer0_outputs[1386]));
    assign layer1_outputs[1019] = ~((layer0_outputs[4699]) | (layer0_outputs[1505]));
    assign layer1_outputs[1020] = ~(layer0_outputs[2918]) | (layer0_outputs[2506]);
    assign layer1_outputs[1021] = ~((layer0_outputs[2879]) & (layer0_outputs[631]));
    assign layer1_outputs[1022] = (layer0_outputs[4909]) & (layer0_outputs[4149]);
    assign layer1_outputs[1023] = ~(layer0_outputs[2620]);
    assign layer1_outputs[1024] = ~(layer0_outputs[960]) | (layer0_outputs[801]);
    assign layer1_outputs[1025] = (layer0_outputs[33]) & ~(layer0_outputs[1937]);
    assign layer1_outputs[1026] = (layer0_outputs[1715]) & ~(layer0_outputs[2788]);
    assign layer1_outputs[1027] = 1'b0;
    assign layer1_outputs[1028] = (layer0_outputs[1789]) | (layer0_outputs[2899]);
    assign layer1_outputs[1029] = ~((layer0_outputs[3669]) ^ (layer0_outputs[2090]));
    assign layer1_outputs[1030] = ~((layer0_outputs[37]) | (layer0_outputs[1575]));
    assign layer1_outputs[1031] = ~(layer0_outputs[1428]) | (layer0_outputs[3815]);
    assign layer1_outputs[1032] = (layer0_outputs[1726]) & (layer0_outputs[851]);
    assign layer1_outputs[1033] = ~(layer0_outputs[556]) | (layer0_outputs[329]);
    assign layer1_outputs[1034] = (layer0_outputs[4027]) | (layer0_outputs[1435]);
    assign layer1_outputs[1035] = 1'b1;
    assign layer1_outputs[1036] = ~((layer0_outputs[3247]) | (layer0_outputs[755]));
    assign layer1_outputs[1037] = layer0_outputs[3559];
    assign layer1_outputs[1038] = (layer0_outputs[3308]) ^ (layer0_outputs[676]);
    assign layer1_outputs[1039] = layer0_outputs[1116];
    assign layer1_outputs[1040] = ~(layer0_outputs[4870]) | (layer0_outputs[5008]);
    assign layer1_outputs[1041] = ~(layer0_outputs[1019]) | (layer0_outputs[4507]);
    assign layer1_outputs[1042] = layer0_outputs[819];
    assign layer1_outputs[1043] = (layer0_outputs[4225]) & ~(layer0_outputs[3631]);
    assign layer1_outputs[1044] = layer0_outputs[1493];
    assign layer1_outputs[1045] = (layer0_outputs[3133]) | (layer0_outputs[402]);
    assign layer1_outputs[1046] = ~(layer0_outputs[328]) | (layer0_outputs[2078]);
    assign layer1_outputs[1047] = layer0_outputs[352];
    assign layer1_outputs[1048] = ~(layer0_outputs[4674]) | (layer0_outputs[3586]);
    assign layer1_outputs[1049] = layer0_outputs[4958];
    assign layer1_outputs[1050] = ~((layer0_outputs[999]) ^ (layer0_outputs[1841]));
    assign layer1_outputs[1051] = (layer0_outputs[1609]) & (layer0_outputs[3223]);
    assign layer1_outputs[1052] = (layer0_outputs[1604]) | (layer0_outputs[151]);
    assign layer1_outputs[1053] = ~(layer0_outputs[1370]) | (layer0_outputs[4417]);
    assign layer1_outputs[1054] = ~(layer0_outputs[1934]) | (layer0_outputs[540]);
    assign layer1_outputs[1055] = (layer0_outputs[2983]) & ~(layer0_outputs[201]);
    assign layer1_outputs[1056] = ~(layer0_outputs[3081]) | (layer0_outputs[211]);
    assign layer1_outputs[1057] = ~(layer0_outputs[3767]) | (layer0_outputs[101]);
    assign layer1_outputs[1058] = ~((layer0_outputs[2725]) & (layer0_outputs[2229]));
    assign layer1_outputs[1059] = layer0_outputs[4123];
    assign layer1_outputs[1060] = layer0_outputs[4551];
    assign layer1_outputs[1061] = ~(layer0_outputs[4182]) | (layer0_outputs[4606]);
    assign layer1_outputs[1062] = (layer0_outputs[485]) & (layer0_outputs[4872]);
    assign layer1_outputs[1063] = (layer0_outputs[4532]) & ~(layer0_outputs[1788]);
    assign layer1_outputs[1064] = (layer0_outputs[1574]) & (layer0_outputs[4063]);
    assign layer1_outputs[1065] = (layer0_outputs[930]) | (layer0_outputs[1076]);
    assign layer1_outputs[1066] = (layer0_outputs[443]) & ~(layer0_outputs[2216]);
    assign layer1_outputs[1067] = layer0_outputs[461];
    assign layer1_outputs[1068] = (layer0_outputs[4256]) | (layer0_outputs[4106]);
    assign layer1_outputs[1069] = (layer0_outputs[2118]) & ~(layer0_outputs[2647]);
    assign layer1_outputs[1070] = ~((layer0_outputs[2302]) ^ (layer0_outputs[4961]));
    assign layer1_outputs[1071] = 1'b0;
    assign layer1_outputs[1072] = ~(layer0_outputs[1565]) | (layer0_outputs[643]);
    assign layer1_outputs[1073] = (layer0_outputs[2147]) | (layer0_outputs[1147]);
    assign layer1_outputs[1074] = ~(layer0_outputs[3594]);
    assign layer1_outputs[1075] = ~(layer0_outputs[365]) | (layer0_outputs[1379]);
    assign layer1_outputs[1076] = ~((layer0_outputs[818]) & (layer0_outputs[3880]));
    assign layer1_outputs[1077] = ~((layer0_outputs[4356]) | (layer0_outputs[3789]));
    assign layer1_outputs[1078] = ~((layer0_outputs[3866]) | (layer0_outputs[5067]));
    assign layer1_outputs[1079] = 1'b1;
    assign layer1_outputs[1080] = ~((layer0_outputs[4161]) | (layer0_outputs[1003]));
    assign layer1_outputs[1081] = ~(layer0_outputs[2592]);
    assign layer1_outputs[1082] = ~(layer0_outputs[4214]);
    assign layer1_outputs[1083] = ~(layer0_outputs[4815]) | (layer0_outputs[2352]);
    assign layer1_outputs[1084] = ~((layer0_outputs[3912]) | (layer0_outputs[2516]));
    assign layer1_outputs[1085] = layer0_outputs[3249];
    assign layer1_outputs[1086] = ~(layer0_outputs[4761]);
    assign layer1_outputs[1087] = ~(layer0_outputs[4982]);
    assign layer1_outputs[1088] = ~(layer0_outputs[1687]) | (layer0_outputs[893]);
    assign layer1_outputs[1089] = (layer0_outputs[3399]) & ~(layer0_outputs[4220]);
    assign layer1_outputs[1090] = (layer0_outputs[755]) ^ (layer0_outputs[1410]);
    assign layer1_outputs[1091] = 1'b0;
    assign layer1_outputs[1092] = ~((layer0_outputs[4598]) & (layer0_outputs[885]));
    assign layer1_outputs[1093] = layer0_outputs[3081];
    assign layer1_outputs[1094] = 1'b0;
    assign layer1_outputs[1095] = (layer0_outputs[4993]) & ~(layer0_outputs[4744]);
    assign layer1_outputs[1096] = ~(layer0_outputs[2053]);
    assign layer1_outputs[1097] = layer0_outputs[2551];
    assign layer1_outputs[1098] = ~(layer0_outputs[4616]) | (layer0_outputs[254]);
    assign layer1_outputs[1099] = (layer0_outputs[1970]) & (layer0_outputs[14]);
    assign layer1_outputs[1100] = (layer0_outputs[2956]) ^ (layer0_outputs[4096]);
    assign layer1_outputs[1101] = (layer0_outputs[981]) & ~(layer0_outputs[4006]);
    assign layer1_outputs[1102] = ~(layer0_outputs[1619]);
    assign layer1_outputs[1103] = (layer0_outputs[111]) | (layer0_outputs[697]);
    assign layer1_outputs[1104] = (layer0_outputs[2617]) & ~(layer0_outputs[3891]);
    assign layer1_outputs[1105] = ~((layer0_outputs[4238]) & (layer0_outputs[3566]));
    assign layer1_outputs[1106] = (layer0_outputs[2639]) | (layer0_outputs[3536]);
    assign layer1_outputs[1107] = layer0_outputs[4113];
    assign layer1_outputs[1108] = layer0_outputs[2502];
    assign layer1_outputs[1109] = ~(layer0_outputs[4536]);
    assign layer1_outputs[1110] = ~(layer0_outputs[732]);
    assign layer1_outputs[1111] = (layer0_outputs[1372]) & ~(layer0_outputs[2634]);
    assign layer1_outputs[1112] = layer0_outputs[3433];
    assign layer1_outputs[1113] = layer0_outputs[4750];
    assign layer1_outputs[1114] = ~(layer0_outputs[2655]) | (layer0_outputs[4502]);
    assign layer1_outputs[1115] = layer0_outputs[1781];
    assign layer1_outputs[1116] = (layer0_outputs[3987]) & ~(layer0_outputs[2622]);
    assign layer1_outputs[1117] = (layer0_outputs[4726]) & ~(layer0_outputs[3813]);
    assign layer1_outputs[1118] = 1'b1;
    assign layer1_outputs[1119] = (layer0_outputs[1050]) & (layer0_outputs[2090]);
    assign layer1_outputs[1120] = layer0_outputs[3378];
    assign layer1_outputs[1121] = (layer0_outputs[524]) & ~(layer0_outputs[3473]);
    assign layer1_outputs[1122] = ~((layer0_outputs[1700]) & (layer0_outputs[5024]));
    assign layer1_outputs[1123] = (layer0_outputs[1308]) & ~(layer0_outputs[144]);
    assign layer1_outputs[1124] = ~((layer0_outputs[2106]) | (layer0_outputs[2249]));
    assign layer1_outputs[1125] = (layer0_outputs[561]) & (layer0_outputs[4887]);
    assign layer1_outputs[1126] = layer0_outputs[4651];
    assign layer1_outputs[1127] = ~(layer0_outputs[612]) | (layer0_outputs[4052]);
    assign layer1_outputs[1128] = ~((layer0_outputs[1840]) & (layer0_outputs[1320]));
    assign layer1_outputs[1129] = layer0_outputs[1092];
    assign layer1_outputs[1130] = ~((layer0_outputs[403]) | (layer0_outputs[4563]));
    assign layer1_outputs[1131] = 1'b1;
    assign layer1_outputs[1132] = 1'b0;
    assign layer1_outputs[1133] = 1'b1;
    assign layer1_outputs[1134] = (layer0_outputs[2715]) & (layer0_outputs[3042]);
    assign layer1_outputs[1135] = ~(layer0_outputs[1780]) | (layer0_outputs[2595]);
    assign layer1_outputs[1136] = layer0_outputs[5097];
    assign layer1_outputs[1137] = 1'b1;
    assign layer1_outputs[1138] = 1'b0;
    assign layer1_outputs[1139] = ~(layer0_outputs[4586]);
    assign layer1_outputs[1140] = (layer0_outputs[1996]) & ~(layer0_outputs[4608]);
    assign layer1_outputs[1141] = 1'b1;
    assign layer1_outputs[1142] = ~((layer0_outputs[3731]) | (layer0_outputs[4364]));
    assign layer1_outputs[1143] = (layer0_outputs[714]) | (layer0_outputs[1436]);
    assign layer1_outputs[1144] = ~((layer0_outputs[3454]) | (layer0_outputs[3064]));
    assign layer1_outputs[1145] = 1'b0;
    assign layer1_outputs[1146] = 1'b0;
    assign layer1_outputs[1147] = ~((layer0_outputs[1673]) | (layer0_outputs[897]));
    assign layer1_outputs[1148] = layer0_outputs[4568];
    assign layer1_outputs[1149] = 1'b1;
    assign layer1_outputs[1150] = 1'b0;
    assign layer1_outputs[1151] = layer0_outputs[1470];
    assign layer1_outputs[1152] = (layer0_outputs[496]) & ~(layer0_outputs[2397]);
    assign layer1_outputs[1153] = ~(layer0_outputs[1424]) | (layer0_outputs[5077]);
    assign layer1_outputs[1154] = (layer0_outputs[2654]) & ~(layer0_outputs[3953]);
    assign layer1_outputs[1155] = 1'b0;
    assign layer1_outputs[1156] = 1'b1;
    assign layer1_outputs[1157] = (layer0_outputs[1247]) | (layer0_outputs[2103]);
    assign layer1_outputs[1158] = ~(layer0_outputs[1923]) | (layer0_outputs[3004]);
    assign layer1_outputs[1159] = ~(layer0_outputs[1979]) | (layer0_outputs[4402]);
    assign layer1_outputs[1160] = (layer0_outputs[1520]) & ~(layer0_outputs[1699]);
    assign layer1_outputs[1161] = ~(layer0_outputs[96]);
    assign layer1_outputs[1162] = ~((layer0_outputs[5039]) & (layer0_outputs[3271]));
    assign layer1_outputs[1163] = ~(layer0_outputs[3724]);
    assign layer1_outputs[1164] = 1'b0;
    assign layer1_outputs[1165] = ~(layer0_outputs[1740]);
    assign layer1_outputs[1166] = 1'b0;
    assign layer1_outputs[1167] = (layer0_outputs[3943]) & ~(layer0_outputs[3520]);
    assign layer1_outputs[1168] = (layer0_outputs[1818]) & ~(layer0_outputs[3369]);
    assign layer1_outputs[1169] = ~(layer0_outputs[1169]) | (layer0_outputs[1991]);
    assign layer1_outputs[1170] = (layer0_outputs[1509]) & ~(layer0_outputs[1962]);
    assign layer1_outputs[1171] = layer0_outputs[458];
    assign layer1_outputs[1172] = layer0_outputs[4167];
    assign layer1_outputs[1173] = ~((layer0_outputs[1331]) | (layer0_outputs[1825]));
    assign layer1_outputs[1174] = (layer0_outputs[4400]) ^ (layer0_outputs[3807]);
    assign layer1_outputs[1175] = (layer0_outputs[3166]) & ~(layer0_outputs[2241]);
    assign layer1_outputs[1176] = (layer0_outputs[4566]) | (layer0_outputs[2668]);
    assign layer1_outputs[1177] = ~((layer0_outputs[3800]) | (layer0_outputs[2911]));
    assign layer1_outputs[1178] = (layer0_outputs[1440]) & ~(layer0_outputs[4857]);
    assign layer1_outputs[1179] = layer0_outputs[3916];
    assign layer1_outputs[1180] = layer0_outputs[3913];
    assign layer1_outputs[1181] = (layer0_outputs[2480]) & ~(layer0_outputs[3087]);
    assign layer1_outputs[1182] = ~(layer0_outputs[1606]) | (layer0_outputs[3195]);
    assign layer1_outputs[1183] = ~(layer0_outputs[4770]);
    assign layer1_outputs[1184] = ~(layer0_outputs[2093]) | (layer0_outputs[1601]);
    assign layer1_outputs[1185] = ~(layer0_outputs[185]) | (layer0_outputs[792]);
    assign layer1_outputs[1186] = 1'b0;
    assign layer1_outputs[1187] = (layer0_outputs[2081]) ^ (layer0_outputs[3003]);
    assign layer1_outputs[1188] = (layer0_outputs[5012]) | (layer0_outputs[867]);
    assign layer1_outputs[1189] = ~(layer0_outputs[4667]);
    assign layer1_outputs[1190] = 1'b0;
    assign layer1_outputs[1191] = layer0_outputs[1274];
    assign layer1_outputs[1192] = (layer0_outputs[1045]) & ~(layer0_outputs[4551]);
    assign layer1_outputs[1193] = (layer0_outputs[393]) & (layer0_outputs[2023]);
    assign layer1_outputs[1194] = ~(layer0_outputs[1144]);
    assign layer1_outputs[1195] = (layer0_outputs[3751]) & ~(layer0_outputs[4949]);
    assign layer1_outputs[1196] = layer0_outputs[2107];
    assign layer1_outputs[1197] = 1'b0;
    assign layer1_outputs[1198] = ~((layer0_outputs[3161]) ^ (layer0_outputs[1559]));
    assign layer1_outputs[1199] = (layer0_outputs[1370]) & ~(layer0_outputs[355]);
    assign layer1_outputs[1200] = ~((layer0_outputs[1576]) & (layer0_outputs[1066]));
    assign layer1_outputs[1201] = 1'b1;
    assign layer1_outputs[1202] = (layer0_outputs[890]) & (layer0_outputs[4842]);
    assign layer1_outputs[1203] = ~(layer0_outputs[1119]) | (layer0_outputs[459]);
    assign layer1_outputs[1204] = ~((layer0_outputs[2877]) & (layer0_outputs[3344]));
    assign layer1_outputs[1205] = 1'b1;
    assign layer1_outputs[1206] = layer0_outputs[3763];
    assign layer1_outputs[1207] = (layer0_outputs[3671]) | (layer0_outputs[1574]);
    assign layer1_outputs[1208] = 1'b0;
    assign layer1_outputs[1209] = ~(layer0_outputs[4221]);
    assign layer1_outputs[1210] = ~((layer0_outputs[2697]) | (layer0_outputs[3518]));
    assign layer1_outputs[1211] = (layer0_outputs[1724]) | (layer0_outputs[4598]);
    assign layer1_outputs[1212] = (layer0_outputs[4661]) & ~(layer0_outputs[2004]);
    assign layer1_outputs[1213] = (layer0_outputs[1093]) ^ (layer0_outputs[712]);
    assign layer1_outputs[1214] = ~((layer0_outputs[2395]) | (layer0_outputs[1026]));
    assign layer1_outputs[1215] = ~((layer0_outputs[4970]) ^ (layer0_outputs[1944]));
    assign layer1_outputs[1216] = ~(layer0_outputs[3108]);
    assign layer1_outputs[1217] = (layer0_outputs[4698]) & ~(layer0_outputs[528]);
    assign layer1_outputs[1218] = ~(layer0_outputs[4331]);
    assign layer1_outputs[1219] = ~(layer0_outputs[336]);
    assign layer1_outputs[1220] = 1'b0;
    assign layer1_outputs[1221] = ~((layer0_outputs[3356]) & (layer0_outputs[4379]));
    assign layer1_outputs[1222] = layer0_outputs[4618];
    assign layer1_outputs[1223] = layer0_outputs[3096];
    assign layer1_outputs[1224] = ~(layer0_outputs[2569]);
    assign layer1_outputs[1225] = ~(layer0_outputs[572]) | (layer0_outputs[21]);
    assign layer1_outputs[1226] = ~((layer0_outputs[1342]) | (layer0_outputs[1595]));
    assign layer1_outputs[1227] = (layer0_outputs[3356]) & ~(layer0_outputs[927]);
    assign layer1_outputs[1228] = (layer0_outputs[1358]) & (layer0_outputs[2847]);
    assign layer1_outputs[1229] = ~((layer0_outputs[373]) | (layer0_outputs[2798]));
    assign layer1_outputs[1230] = (layer0_outputs[998]) & (layer0_outputs[1598]);
    assign layer1_outputs[1231] = ~((layer0_outputs[4875]) & (layer0_outputs[3109]));
    assign layer1_outputs[1232] = ~((layer0_outputs[797]) & (layer0_outputs[1569]));
    assign layer1_outputs[1233] = 1'b0;
    assign layer1_outputs[1234] = 1'b1;
    assign layer1_outputs[1235] = (layer0_outputs[1027]) | (layer0_outputs[4671]);
    assign layer1_outputs[1236] = 1'b1;
    assign layer1_outputs[1237] = (layer0_outputs[2540]) | (layer0_outputs[2999]);
    assign layer1_outputs[1238] = ~(layer0_outputs[2667]);
    assign layer1_outputs[1239] = ~((layer0_outputs[3756]) & (layer0_outputs[2045]));
    assign layer1_outputs[1240] = 1'b1;
    assign layer1_outputs[1241] = ~((layer0_outputs[3888]) | (layer0_outputs[444]));
    assign layer1_outputs[1242] = ~((layer0_outputs[1457]) & (layer0_outputs[4423]));
    assign layer1_outputs[1243] = ~(layer0_outputs[2992]);
    assign layer1_outputs[1244] = ~(layer0_outputs[1661]);
    assign layer1_outputs[1245] = ~(layer0_outputs[2916]) | (layer0_outputs[345]);
    assign layer1_outputs[1246] = (layer0_outputs[1299]) & (layer0_outputs[1900]);
    assign layer1_outputs[1247] = layer0_outputs[313];
    assign layer1_outputs[1248] = layer0_outputs[3094];
    assign layer1_outputs[1249] = ~(layer0_outputs[372]) | (layer0_outputs[2285]);
    assign layer1_outputs[1250] = ~(layer0_outputs[273]);
    assign layer1_outputs[1251] = ~(layer0_outputs[784]);
    assign layer1_outputs[1252] = (layer0_outputs[4519]) & ~(layer0_outputs[1882]);
    assign layer1_outputs[1253] = 1'b0;
    assign layer1_outputs[1254] = ~(layer0_outputs[3434]) | (layer0_outputs[4682]);
    assign layer1_outputs[1255] = (layer0_outputs[308]) & ~(layer0_outputs[1624]);
    assign layer1_outputs[1256] = ~((layer0_outputs[3214]) | (layer0_outputs[1219]));
    assign layer1_outputs[1257] = (layer0_outputs[4596]) & ~(layer0_outputs[2799]);
    assign layer1_outputs[1258] = (layer0_outputs[3809]) | (layer0_outputs[5023]);
    assign layer1_outputs[1259] = ~((layer0_outputs[4250]) & (layer0_outputs[157]));
    assign layer1_outputs[1260] = (layer0_outputs[2351]) | (layer0_outputs[4458]);
    assign layer1_outputs[1261] = ~((layer0_outputs[3337]) & (layer0_outputs[4218]));
    assign layer1_outputs[1262] = ~(layer0_outputs[419]);
    assign layer1_outputs[1263] = (layer0_outputs[4438]) & ~(layer0_outputs[3364]);
    assign layer1_outputs[1264] = layer0_outputs[356];
    assign layer1_outputs[1265] = layer0_outputs[932];
    assign layer1_outputs[1266] = layer0_outputs[2342];
    assign layer1_outputs[1267] = (layer0_outputs[162]) & (layer0_outputs[74]);
    assign layer1_outputs[1268] = ~((layer0_outputs[4617]) & (layer0_outputs[3351]));
    assign layer1_outputs[1269] = ~(layer0_outputs[3975]) | (layer0_outputs[4875]);
    assign layer1_outputs[1270] = ~(layer0_outputs[3666]);
    assign layer1_outputs[1271] = (layer0_outputs[1396]) & ~(layer0_outputs[3825]);
    assign layer1_outputs[1272] = ~(layer0_outputs[248]) | (layer0_outputs[2130]);
    assign layer1_outputs[1273] = ~(layer0_outputs[2982]) | (layer0_outputs[870]);
    assign layer1_outputs[1274] = 1'b0;
    assign layer1_outputs[1275] = 1'b0;
    assign layer1_outputs[1276] = ~(layer0_outputs[1519]) | (layer0_outputs[3170]);
    assign layer1_outputs[1277] = ~(layer0_outputs[4574]);
    assign layer1_outputs[1278] = (layer0_outputs[2492]) ^ (layer0_outputs[1098]);
    assign layer1_outputs[1279] = 1'b1;
    assign layer1_outputs[1280] = ~(layer0_outputs[3791]) | (layer0_outputs[4422]);
    assign layer1_outputs[1281] = ~((layer0_outputs[421]) | (layer0_outputs[3983]));
    assign layer1_outputs[1282] = ~(layer0_outputs[3364]);
    assign layer1_outputs[1283] = (layer0_outputs[1286]) & ~(layer0_outputs[4076]);
    assign layer1_outputs[1284] = (layer0_outputs[3667]) & (layer0_outputs[3649]);
    assign layer1_outputs[1285] = ~((layer0_outputs[3491]) & (layer0_outputs[1314]));
    assign layer1_outputs[1286] = layer0_outputs[469];
    assign layer1_outputs[1287] = layer0_outputs[2730];
    assign layer1_outputs[1288] = layer0_outputs[4948];
    assign layer1_outputs[1289] = 1'b1;
    assign layer1_outputs[1290] = ~((layer0_outputs[2589]) | (layer0_outputs[619]));
    assign layer1_outputs[1291] = ~((layer0_outputs[4523]) | (layer0_outputs[2166]));
    assign layer1_outputs[1292] = ~((layer0_outputs[910]) & (layer0_outputs[821]));
    assign layer1_outputs[1293] = ~(layer0_outputs[1115]) | (layer0_outputs[4185]);
    assign layer1_outputs[1294] = layer0_outputs[693];
    assign layer1_outputs[1295] = ~(layer0_outputs[1814]);
    assign layer1_outputs[1296] = (layer0_outputs[1681]) ^ (layer0_outputs[1300]);
    assign layer1_outputs[1297] = ~(layer0_outputs[2633]);
    assign layer1_outputs[1298] = (layer0_outputs[4079]) & ~(layer0_outputs[3370]);
    assign layer1_outputs[1299] = layer0_outputs[2568];
    assign layer1_outputs[1300] = 1'b0;
    assign layer1_outputs[1301] = layer0_outputs[1233];
    assign layer1_outputs[1302] = (layer0_outputs[4734]) & ~(layer0_outputs[2794]);
    assign layer1_outputs[1303] = layer0_outputs[143];
    assign layer1_outputs[1304] = ~(layer0_outputs[3352]) | (layer0_outputs[1695]);
    assign layer1_outputs[1305] = (layer0_outputs[3058]) & (layer0_outputs[1323]);
    assign layer1_outputs[1306] = ~((layer0_outputs[4986]) | (layer0_outputs[4466]));
    assign layer1_outputs[1307] = ~(layer0_outputs[4995]) | (layer0_outputs[4081]);
    assign layer1_outputs[1308] = ~(layer0_outputs[1152]);
    assign layer1_outputs[1309] = (layer0_outputs[128]) & ~(layer0_outputs[4124]);
    assign layer1_outputs[1310] = (layer0_outputs[2378]) & (layer0_outputs[4886]);
    assign layer1_outputs[1311] = ~(layer0_outputs[1566]);
    assign layer1_outputs[1312] = ~((layer0_outputs[3494]) | (layer0_outputs[1218]));
    assign layer1_outputs[1313] = ~(layer0_outputs[2043]) | (layer0_outputs[4996]);
    assign layer1_outputs[1314] = ~((layer0_outputs[312]) ^ (layer0_outputs[1958]));
    assign layer1_outputs[1315] = (layer0_outputs[4664]) | (layer0_outputs[4782]);
    assign layer1_outputs[1316] = layer0_outputs[4847];
    assign layer1_outputs[1317] = 1'b1;
    assign layer1_outputs[1318] = ~(layer0_outputs[2981]) | (layer0_outputs[2745]);
    assign layer1_outputs[1319] = (layer0_outputs[178]) & (layer0_outputs[4204]);
    assign layer1_outputs[1320] = ~(layer0_outputs[1497]) | (layer0_outputs[1361]);
    assign layer1_outputs[1321] = layer0_outputs[1061];
    assign layer1_outputs[1322] = ~((layer0_outputs[3931]) ^ (layer0_outputs[2442]));
    assign layer1_outputs[1323] = 1'b0;
    assign layer1_outputs[1324] = layer0_outputs[2469];
    assign layer1_outputs[1325] = ~((layer0_outputs[295]) | (layer0_outputs[2216]));
    assign layer1_outputs[1326] = (layer0_outputs[3212]) | (layer0_outputs[4362]);
    assign layer1_outputs[1327] = ~(layer0_outputs[4366]);
    assign layer1_outputs[1328] = (layer0_outputs[5074]) | (layer0_outputs[2702]);
    assign layer1_outputs[1329] = ~(layer0_outputs[2210]);
    assign layer1_outputs[1330] = 1'b0;
    assign layer1_outputs[1331] = (layer0_outputs[1056]) | (layer0_outputs[2941]);
    assign layer1_outputs[1332] = (layer0_outputs[2139]) | (layer0_outputs[2362]);
    assign layer1_outputs[1333] = ~(layer0_outputs[1171]) | (layer0_outputs[1833]);
    assign layer1_outputs[1334] = 1'b1;
    assign layer1_outputs[1335] = (layer0_outputs[3365]) & (layer0_outputs[35]);
    assign layer1_outputs[1336] = layer0_outputs[3325];
    assign layer1_outputs[1337] = (layer0_outputs[3668]) & ~(layer0_outputs[1013]);
    assign layer1_outputs[1338] = 1'b1;
    assign layer1_outputs[1339] = (layer0_outputs[3819]) & ~(layer0_outputs[3330]);
    assign layer1_outputs[1340] = ~(layer0_outputs[3968]) | (layer0_outputs[4974]);
    assign layer1_outputs[1341] = (layer0_outputs[1090]) ^ (layer0_outputs[2311]);
    assign layer1_outputs[1342] = (layer0_outputs[743]) & ~(layer0_outputs[2626]);
    assign layer1_outputs[1343] = (layer0_outputs[4819]) & (layer0_outputs[2054]);
    assign layer1_outputs[1344] = 1'b0;
    assign layer1_outputs[1345] = ~(layer0_outputs[1543]) | (layer0_outputs[4111]);
    assign layer1_outputs[1346] = ~(layer0_outputs[1640]) | (layer0_outputs[220]);
    assign layer1_outputs[1347] = 1'b0;
    assign layer1_outputs[1348] = (layer0_outputs[4871]) & ~(layer0_outputs[2588]);
    assign layer1_outputs[1349] = ~((layer0_outputs[2544]) | (layer0_outputs[142]));
    assign layer1_outputs[1350] = ~((layer0_outputs[3860]) & (layer0_outputs[4066]));
    assign layer1_outputs[1351] = ~(layer0_outputs[2003]);
    assign layer1_outputs[1352] = (layer0_outputs[4749]) | (layer0_outputs[2165]);
    assign layer1_outputs[1353] = layer0_outputs[535];
    assign layer1_outputs[1354] = ~(layer0_outputs[4049]) | (layer0_outputs[2695]);
    assign layer1_outputs[1355] = (layer0_outputs[4427]) | (layer0_outputs[3503]);
    assign layer1_outputs[1356] = ~((layer0_outputs[3844]) | (layer0_outputs[3825]));
    assign layer1_outputs[1357] = ~((layer0_outputs[3707]) & (layer0_outputs[3762]));
    assign layer1_outputs[1358] = 1'b0;
    assign layer1_outputs[1359] = (layer0_outputs[4741]) & (layer0_outputs[47]);
    assign layer1_outputs[1360] = layer0_outputs[4622];
    assign layer1_outputs[1361] = 1'b0;
    assign layer1_outputs[1362] = ~(layer0_outputs[2499]);
    assign layer1_outputs[1363] = layer0_outputs[1378];
    assign layer1_outputs[1364] = (layer0_outputs[2415]) & (layer0_outputs[492]);
    assign layer1_outputs[1365] = (layer0_outputs[2370]) | (layer0_outputs[3114]);
    assign layer1_outputs[1366] = ~(layer0_outputs[728]) | (layer0_outputs[235]);
    assign layer1_outputs[1367] = ~(layer0_outputs[3416]);
    assign layer1_outputs[1368] = ~((layer0_outputs[4417]) ^ (layer0_outputs[685]));
    assign layer1_outputs[1369] = ~(layer0_outputs[2276]) | (layer0_outputs[3899]);
    assign layer1_outputs[1370] = (layer0_outputs[2256]) & ~(layer0_outputs[238]);
    assign layer1_outputs[1371] = (layer0_outputs[2077]) & ~(layer0_outputs[2115]);
    assign layer1_outputs[1372] = ~(layer0_outputs[3268]) | (layer0_outputs[2552]);
    assign layer1_outputs[1373] = (layer0_outputs[5016]) & ~(layer0_outputs[3571]);
    assign layer1_outputs[1374] = ~(layer0_outputs[4639]) | (layer0_outputs[341]);
    assign layer1_outputs[1375] = ~((layer0_outputs[1754]) ^ (layer0_outputs[28]));
    assign layer1_outputs[1376] = 1'b0;
    assign layer1_outputs[1377] = layer0_outputs[1189];
    assign layer1_outputs[1378] = (layer0_outputs[2837]) & ~(layer0_outputs[301]);
    assign layer1_outputs[1379] = ~((layer0_outputs[828]) & (layer0_outputs[5101]));
    assign layer1_outputs[1380] = ~((layer0_outputs[351]) & (layer0_outputs[3618]));
    assign layer1_outputs[1381] = (layer0_outputs[632]) & ~(layer0_outputs[3237]);
    assign layer1_outputs[1382] = (layer0_outputs[2376]) ^ (layer0_outputs[4826]);
    assign layer1_outputs[1383] = ~(layer0_outputs[1168]);
    assign layer1_outputs[1384] = ~(layer0_outputs[4777]);
    assign layer1_outputs[1385] = ~(layer0_outputs[1245]);
    assign layer1_outputs[1386] = 1'b1;
    assign layer1_outputs[1387] = 1'b1;
    assign layer1_outputs[1388] = 1'b0;
    assign layer1_outputs[1389] = ~(layer0_outputs[705]);
    assign layer1_outputs[1390] = (layer0_outputs[2245]) & ~(layer0_outputs[1847]);
    assign layer1_outputs[1391] = ~((layer0_outputs[4508]) & (layer0_outputs[181]));
    assign layer1_outputs[1392] = (layer0_outputs[2676]) & ~(layer0_outputs[1159]);
    assign layer1_outputs[1393] = 1'b0;
    assign layer1_outputs[1394] = ~((layer0_outputs[4455]) & (layer0_outputs[1763]));
    assign layer1_outputs[1395] = ~((layer0_outputs[1563]) & (layer0_outputs[1268]));
    assign layer1_outputs[1396] = ~(layer0_outputs[2839]) | (layer0_outputs[1743]);
    assign layer1_outputs[1397] = layer0_outputs[2711];
    assign layer1_outputs[1398] = (layer0_outputs[465]) | (layer0_outputs[1744]);
    assign layer1_outputs[1399] = (layer0_outputs[916]) & ~(layer0_outputs[4879]);
    assign layer1_outputs[1400] = (layer0_outputs[4164]) & (layer0_outputs[2952]);
    assign layer1_outputs[1401] = (layer0_outputs[3134]) & (layer0_outputs[1929]);
    assign layer1_outputs[1402] = layer0_outputs[1431];
    assign layer1_outputs[1403] = (layer0_outputs[1540]) ^ (layer0_outputs[300]);
    assign layer1_outputs[1404] = ~(layer0_outputs[4908]) | (layer0_outputs[1732]);
    assign layer1_outputs[1405] = ~((layer0_outputs[667]) | (layer0_outputs[3398]));
    assign layer1_outputs[1406] = 1'b0;
    assign layer1_outputs[1407] = 1'b1;
    assign layer1_outputs[1408] = (layer0_outputs[867]) & ~(layer0_outputs[1473]);
    assign layer1_outputs[1409] = layer0_outputs[4678];
    assign layer1_outputs[1410] = 1'b0;
    assign layer1_outputs[1411] = ~((layer0_outputs[1366]) & (layer0_outputs[3171]));
    assign layer1_outputs[1412] = ~(layer0_outputs[949]) | (layer0_outputs[88]);
    assign layer1_outputs[1413] = (layer0_outputs[1658]) & (layer0_outputs[2153]);
    assign layer1_outputs[1414] = 1'b1;
    assign layer1_outputs[1415] = 1'b1;
    assign layer1_outputs[1416] = 1'b1;
    assign layer1_outputs[1417] = ~(layer0_outputs[2365]);
    assign layer1_outputs[1418] = ~((layer0_outputs[1048]) & (layer0_outputs[4704]));
    assign layer1_outputs[1419] = 1'b0;
    assign layer1_outputs[1420] = layer0_outputs[1199];
    assign layer1_outputs[1421] = (layer0_outputs[903]) | (layer0_outputs[4644]);
    assign layer1_outputs[1422] = layer0_outputs[605];
    assign layer1_outputs[1423] = (layer0_outputs[1618]) | (layer0_outputs[1811]);
    assign layer1_outputs[1424] = ~(layer0_outputs[2487]);
    assign layer1_outputs[1425] = ~(layer0_outputs[3541]);
    assign layer1_outputs[1426] = ~((layer0_outputs[4556]) | (layer0_outputs[1359]));
    assign layer1_outputs[1427] = ~(layer0_outputs[3218]);
    assign layer1_outputs[1428] = (layer0_outputs[497]) & (layer0_outputs[4461]);
    assign layer1_outputs[1429] = ~(layer0_outputs[1105]) | (layer0_outputs[64]);
    assign layer1_outputs[1430] = ~((layer0_outputs[4140]) & (layer0_outputs[2208]));
    assign layer1_outputs[1431] = (layer0_outputs[95]) & ~(layer0_outputs[3834]);
    assign layer1_outputs[1432] = ~(layer0_outputs[2279]) | (layer0_outputs[3628]);
    assign layer1_outputs[1433] = (layer0_outputs[226]) & (layer0_outputs[2250]);
    assign layer1_outputs[1434] = ~((layer0_outputs[1953]) ^ (layer0_outputs[714]));
    assign layer1_outputs[1435] = ~(layer0_outputs[1246]) | (layer0_outputs[2561]);
    assign layer1_outputs[1436] = layer0_outputs[844];
    assign layer1_outputs[1437] = layer0_outputs[1392];
    assign layer1_outputs[1438] = ~(layer0_outputs[5116]) | (layer0_outputs[2311]);
    assign layer1_outputs[1439] = layer0_outputs[3016];
    assign layer1_outputs[1440] = (layer0_outputs[1768]) & ~(layer0_outputs[2326]);
    assign layer1_outputs[1441] = 1'b1;
    assign layer1_outputs[1442] = (layer0_outputs[2895]) & ~(layer0_outputs[1079]);
    assign layer1_outputs[1443] = ~((layer0_outputs[655]) ^ (layer0_outputs[4222]));
    assign layer1_outputs[1444] = ~((layer0_outputs[4645]) | (layer0_outputs[3646]));
    assign layer1_outputs[1445] = (layer0_outputs[4125]) & ~(layer0_outputs[1010]);
    assign layer1_outputs[1446] = 1'b0;
    assign layer1_outputs[1447] = 1'b1;
    assign layer1_outputs[1448] = 1'b1;
    assign layer1_outputs[1449] = ~(layer0_outputs[1215]);
    assign layer1_outputs[1450] = layer0_outputs[687];
    assign layer1_outputs[1451] = ~(layer0_outputs[4354]);
    assign layer1_outputs[1452] = layer0_outputs[2689];
    assign layer1_outputs[1453] = 1'b0;
    assign layer1_outputs[1454] = (layer0_outputs[514]) ^ (layer0_outputs[67]);
    assign layer1_outputs[1455] = ~(layer0_outputs[2122]) | (layer0_outputs[4554]);
    assign layer1_outputs[1456] = 1'b1;
    assign layer1_outputs[1457] = ~((layer0_outputs[2646]) | (layer0_outputs[2261]));
    assign layer1_outputs[1458] = ~(layer0_outputs[1227]) | (layer0_outputs[3584]);
    assign layer1_outputs[1459] = ~((layer0_outputs[1278]) | (layer0_outputs[4999]));
    assign layer1_outputs[1460] = (layer0_outputs[850]) | (layer0_outputs[5088]);
    assign layer1_outputs[1461] = (layer0_outputs[4394]) & (layer0_outputs[2474]);
    assign layer1_outputs[1462] = ~((layer0_outputs[191]) | (layer0_outputs[2359]));
    assign layer1_outputs[1463] = (layer0_outputs[3099]) & (layer0_outputs[2980]);
    assign layer1_outputs[1464] = ~(layer0_outputs[4853]);
    assign layer1_outputs[1465] = (layer0_outputs[1632]) & ~(layer0_outputs[3470]);
    assign layer1_outputs[1466] = (layer0_outputs[2813]) & ~(layer0_outputs[374]);
    assign layer1_outputs[1467] = layer0_outputs[1407];
    assign layer1_outputs[1468] = (layer0_outputs[2127]) & (layer0_outputs[858]);
    assign layer1_outputs[1469] = ~(layer0_outputs[4912]);
    assign layer1_outputs[1470] = ~(layer0_outputs[2483]) | (layer0_outputs[2997]);
    assign layer1_outputs[1471] = ~(layer0_outputs[1117]) | (layer0_outputs[1200]);
    assign layer1_outputs[1472] = (layer0_outputs[2966]) & (layer0_outputs[2344]);
    assign layer1_outputs[1473] = 1'b0;
    assign layer1_outputs[1474] = ~(layer0_outputs[2673]);
    assign layer1_outputs[1475] = (layer0_outputs[2323]) & (layer0_outputs[1505]);
    assign layer1_outputs[1476] = 1'b0;
    assign layer1_outputs[1477] = layer0_outputs[2517];
    assign layer1_outputs[1478] = ~((layer0_outputs[3807]) & (layer0_outputs[3889]));
    assign layer1_outputs[1479] = ~(layer0_outputs[2426]);
    assign layer1_outputs[1480] = 1'b1;
    assign layer1_outputs[1481] = ~((layer0_outputs[1714]) | (layer0_outputs[2355]));
    assign layer1_outputs[1482] = ~((layer0_outputs[2284]) | (layer0_outputs[4813]));
    assign layer1_outputs[1483] = (layer0_outputs[2531]) & (layer0_outputs[42]);
    assign layer1_outputs[1484] = 1'b1;
    assign layer1_outputs[1485] = ~(layer0_outputs[3147]) | (layer0_outputs[2438]);
    assign layer1_outputs[1486] = ~(layer0_outputs[2616]);
    assign layer1_outputs[1487] = ~(layer0_outputs[1224]);
    assign layer1_outputs[1488] = ~(layer0_outputs[3]);
    assign layer1_outputs[1489] = ~(layer0_outputs[4248]);
    assign layer1_outputs[1490] = 1'b0;
    assign layer1_outputs[1491] = (layer0_outputs[3020]) & ~(layer0_outputs[1436]);
    assign layer1_outputs[1492] = 1'b0;
    assign layer1_outputs[1493] = ~((layer0_outputs[3901]) & (layer0_outputs[929]));
    assign layer1_outputs[1494] = (layer0_outputs[1699]) & ~(layer0_outputs[2423]);
    assign layer1_outputs[1495] = ~((layer0_outputs[703]) | (layer0_outputs[879]));
    assign layer1_outputs[1496] = (layer0_outputs[4933]) & ~(layer0_outputs[190]);
    assign layer1_outputs[1497] = ~((layer0_outputs[362]) & (layer0_outputs[4711]));
    assign layer1_outputs[1498] = ~(layer0_outputs[2560]) | (layer0_outputs[29]);
    assign layer1_outputs[1499] = (layer0_outputs[2169]) & ~(layer0_outputs[2380]);
    assign layer1_outputs[1500] = ~(layer0_outputs[689]) | (layer0_outputs[1677]);
    assign layer1_outputs[1501] = (layer0_outputs[385]) & ~(layer0_outputs[1713]);
    assign layer1_outputs[1502] = (layer0_outputs[3446]) & (layer0_outputs[995]);
    assign layer1_outputs[1503] = (layer0_outputs[440]) & (layer0_outputs[86]);
    assign layer1_outputs[1504] = (layer0_outputs[1553]) & ~(layer0_outputs[154]);
    assign layer1_outputs[1505] = layer0_outputs[4706];
    assign layer1_outputs[1506] = (layer0_outputs[3623]) & (layer0_outputs[7]);
    assign layer1_outputs[1507] = ~(layer0_outputs[4156]) | (layer0_outputs[3238]);
    assign layer1_outputs[1508] = layer0_outputs[1874];
    assign layer1_outputs[1509] = 1'b0;
    assign layer1_outputs[1510] = ~(layer0_outputs[1719]) | (layer0_outputs[2280]);
    assign layer1_outputs[1511] = layer0_outputs[154];
    assign layer1_outputs[1512] = layer0_outputs[1];
    assign layer1_outputs[1513] = (layer0_outputs[3839]) & ~(layer0_outputs[4779]);
    assign layer1_outputs[1514] = ~((layer0_outputs[4978]) ^ (layer0_outputs[114]));
    assign layer1_outputs[1515] = (layer0_outputs[2098]) & (layer0_outputs[797]);
    assign layer1_outputs[1516] = layer0_outputs[2533];
    assign layer1_outputs[1517] = ~(layer0_outputs[4748]);
    assign layer1_outputs[1518] = (layer0_outputs[2306]) & ~(layer0_outputs[134]);
    assign layer1_outputs[1519] = layer0_outputs[2791];
    assign layer1_outputs[1520] = (layer0_outputs[3310]) & ~(layer0_outputs[3053]);
    assign layer1_outputs[1521] = ~(layer0_outputs[1163]);
    assign layer1_outputs[1522] = (layer0_outputs[4722]) | (layer0_outputs[3662]);
    assign layer1_outputs[1523] = layer0_outputs[2573];
    assign layer1_outputs[1524] = (layer0_outputs[2062]) & (layer0_outputs[793]);
    assign layer1_outputs[1525] = ~((layer0_outputs[2430]) | (layer0_outputs[4510]));
    assign layer1_outputs[1526] = (layer0_outputs[2507]) | (layer0_outputs[1524]);
    assign layer1_outputs[1527] = ~(layer0_outputs[4918]) | (layer0_outputs[3555]);
    assign layer1_outputs[1528] = ~((layer0_outputs[1102]) & (layer0_outputs[4872]));
    assign layer1_outputs[1529] = ~(layer0_outputs[3120]) | (layer0_outputs[896]);
    assign layer1_outputs[1530] = ~(layer0_outputs[2083]);
    assign layer1_outputs[1531] = (layer0_outputs[4908]) & (layer0_outputs[1365]);
    assign layer1_outputs[1532] = (layer0_outputs[1871]) & ~(layer0_outputs[3772]);
    assign layer1_outputs[1533] = ~((layer0_outputs[2048]) | (layer0_outputs[4524]));
    assign layer1_outputs[1534] = (layer0_outputs[3141]) & ~(layer0_outputs[4349]);
    assign layer1_outputs[1535] = ~(layer0_outputs[4044]);
    assign layer1_outputs[1536] = ~(layer0_outputs[4239]);
    assign layer1_outputs[1537] = 1'b1;
    assign layer1_outputs[1538] = (layer0_outputs[3958]) & ~(layer0_outputs[73]);
    assign layer1_outputs[1539] = ~(layer0_outputs[3039]) | (layer0_outputs[3998]);
    assign layer1_outputs[1540] = layer0_outputs[1218];
    assign layer1_outputs[1541] = ~((layer0_outputs[4391]) | (layer0_outputs[1800]));
    assign layer1_outputs[1542] = ~(layer0_outputs[3062]);
    assign layer1_outputs[1543] = (layer0_outputs[3226]) & (layer0_outputs[3653]);
    assign layer1_outputs[1544] = ~(layer0_outputs[1914]);
    assign layer1_outputs[1545] = (layer0_outputs[2185]) & ~(layer0_outputs[806]);
    assign layer1_outputs[1546] = ~((layer0_outputs[4389]) & (layer0_outputs[3690]));
    assign layer1_outputs[1547] = ~(layer0_outputs[2454]);
    assign layer1_outputs[1548] = 1'b1;
    assign layer1_outputs[1549] = ~((layer0_outputs[2407]) & (layer0_outputs[662]));
    assign layer1_outputs[1550] = ~(layer0_outputs[1732]);
    assign layer1_outputs[1551] = (layer0_outputs[238]) | (layer0_outputs[790]);
    assign layer1_outputs[1552] = ~(layer0_outputs[3615]);
    assign layer1_outputs[1553] = 1'b0;
    assign layer1_outputs[1554] = ~(layer0_outputs[4504]);
    assign layer1_outputs[1555] = 1'b1;
    assign layer1_outputs[1556] = ~(layer0_outputs[2858]);
    assign layer1_outputs[1557] = (layer0_outputs[3487]) & (layer0_outputs[4070]);
    assign layer1_outputs[1558] = ~(layer0_outputs[677]);
    assign layer1_outputs[1559] = ~(layer0_outputs[76]);
    assign layer1_outputs[1560] = (layer0_outputs[2260]) & ~(layer0_outputs[2802]);
    assign layer1_outputs[1561] = 1'b1;
    assign layer1_outputs[1562] = layer0_outputs[427];
    assign layer1_outputs[1563] = ~(layer0_outputs[4437]);
    assign layer1_outputs[1564] = (layer0_outputs[1656]) & ~(layer0_outputs[4538]);
    assign layer1_outputs[1565] = layer0_outputs[3956];
    assign layer1_outputs[1566] = 1'b1;
    assign layer1_outputs[1567] = 1'b0;
    assign layer1_outputs[1568] = 1'b1;
    assign layer1_outputs[1569] = ~(layer0_outputs[1892]);
    assign layer1_outputs[1570] = 1'b1;
    assign layer1_outputs[1571] = ~(layer0_outputs[3057]);
    assign layer1_outputs[1572] = ~((layer0_outputs[4335]) | (layer0_outputs[1767]));
    assign layer1_outputs[1573] = 1'b0;
    assign layer1_outputs[1574] = ~((layer0_outputs[3922]) ^ (layer0_outputs[2083]));
    assign layer1_outputs[1575] = ~(layer0_outputs[297]);
    assign layer1_outputs[1576] = (layer0_outputs[2836]) ^ (layer0_outputs[4493]);
    assign layer1_outputs[1577] = (layer0_outputs[3994]) & ~(layer0_outputs[892]);
    assign layer1_outputs[1578] = ~(layer0_outputs[3896]);
    assign layer1_outputs[1579] = ~((layer0_outputs[510]) & (layer0_outputs[1198]));
    assign layer1_outputs[1580] = 1'b0;
    assign layer1_outputs[1581] = ~(layer0_outputs[141]) | (layer0_outputs[601]);
    assign layer1_outputs[1582] = 1'b0;
    assign layer1_outputs[1583] = 1'b0;
    assign layer1_outputs[1584] = (layer0_outputs[56]) & ~(layer0_outputs[3775]);
    assign layer1_outputs[1585] = 1'b1;
    assign layer1_outputs[1586] = ~(layer0_outputs[352]) | (layer0_outputs[4158]);
    assign layer1_outputs[1587] = 1'b0;
    assign layer1_outputs[1588] = ~(layer0_outputs[2444]) | (layer0_outputs[2114]);
    assign layer1_outputs[1589] = 1'b0;
    assign layer1_outputs[1590] = ~((layer0_outputs[1406]) & (layer0_outputs[4943]));
    assign layer1_outputs[1591] = ~(layer0_outputs[3849]);
    assign layer1_outputs[1592] = ~((layer0_outputs[4035]) & (layer0_outputs[185]));
    assign layer1_outputs[1593] = 1'b1;
    assign layer1_outputs[1594] = layer0_outputs[5054];
    assign layer1_outputs[1595] = (layer0_outputs[1706]) & ~(layer0_outputs[338]);
    assign layer1_outputs[1596] = 1'b0;
    assign layer1_outputs[1597] = (layer0_outputs[109]) & ~(layer0_outputs[3306]);
    assign layer1_outputs[1598] = (layer0_outputs[1482]) & (layer0_outputs[2006]);
    assign layer1_outputs[1599] = (layer0_outputs[1705]) & ~(layer0_outputs[1751]);
    assign layer1_outputs[1600] = ~(layer0_outputs[4419]) | (layer0_outputs[97]);
    assign layer1_outputs[1601] = ~(layer0_outputs[610]);
    assign layer1_outputs[1602] = 1'b1;
    assign layer1_outputs[1603] = (layer0_outputs[5036]) & ~(layer0_outputs[1385]);
    assign layer1_outputs[1604] = 1'b0;
    assign layer1_outputs[1605] = layer0_outputs[2109];
    assign layer1_outputs[1606] = ~((layer0_outputs[1674]) | (layer0_outputs[3138]));
    assign layer1_outputs[1607] = (layer0_outputs[3098]) & ~(layer0_outputs[147]);
    assign layer1_outputs[1608] = ~((layer0_outputs[1253]) & (layer0_outputs[1745]));
    assign layer1_outputs[1609] = (layer0_outputs[439]) ^ (layer0_outputs[2291]);
    assign layer1_outputs[1610] = (layer0_outputs[2631]) | (layer0_outputs[1853]);
    assign layer1_outputs[1611] = ~(layer0_outputs[4044]) | (layer0_outputs[13]);
    assign layer1_outputs[1612] = ~((layer0_outputs[3994]) | (layer0_outputs[2842]));
    assign layer1_outputs[1613] = layer0_outputs[4045];
    assign layer1_outputs[1614] = ~(layer0_outputs[306]);
    assign layer1_outputs[1615] = ~((layer0_outputs[1394]) | (layer0_outputs[1792]));
    assign layer1_outputs[1616] = ~((layer0_outputs[2158]) ^ (layer0_outputs[4873]));
    assign layer1_outputs[1617] = (layer0_outputs[3535]) | (layer0_outputs[2889]);
    assign layer1_outputs[1618] = 1'b1;
    assign layer1_outputs[1619] = ~(layer0_outputs[3471]) | (layer0_outputs[4249]);
    assign layer1_outputs[1620] = layer0_outputs[3261];
    assign layer1_outputs[1621] = layer0_outputs[3859];
    assign layer1_outputs[1622] = (layer0_outputs[3907]) | (layer0_outputs[4488]);
    assign layer1_outputs[1623] = layer0_outputs[5090];
    assign layer1_outputs[1624] = (layer0_outputs[2374]) & ~(layer0_outputs[1512]);
    assign layer1_outputs[1625] = ~(layer0_outputs[812]) | (layer0_outputs[696]);
    assign layer1_outputs[1626] = 1'b1;
    assign layer1_outputs[1627] = ~((layer0_outputs[3948]) & (layer0_outputs[845]));
    assign layer1_outputs[1628] = (layer0_outputs[3207]) & ~(layer0_outputs[4955]);
    assign layer1_outputs[1629] = 1'b1;
    assign layer1_outputs[1630] = ~(layer0_outputs[2967]) | (layer0_outputs[1295]);
    assign layer1_outputs[1631] = ~(layer0_outputs[3682]);
    assign layer1_outputs[1632] = ~(layer0_outputs[2793]);
    assign layer1_outputs[1633] = layer0_outputs[3622];
    assign layer1_outputs[1634] = layer0_outputs[2543];
    assign layer1_outputs[1635] = 1'b0;
    assign layer1_outputs[1636] = ~(layer0_outputs[3043]);
    assign layer1_outputs[1637] = layer0_outputs[4361];
    assign layer1_outputs[1638] = (layer0_outputs[3230]) & (layer0_outputs[4414]);
    assign layer1_outputs[1639] = (layer0_outputs[4051]) & ~(layer0_outputs[2516]);
    assign layer1_outputs[1640] = 1'b0;
    assign layer1_outputs[1641] = ~((layer0_outputs[1924]) ^ (layer0_outputs[4873]));
    assign layer1_outputs[1642] = 1'b1;
    assign layer1_outputs[1643] = ~(layer0_outputs[504]) | (layer0_outputs[1053]);
    assign layer1_outputs[1644] = layer0_outputs[2731];
    assign layer1_outputs[1645] = ~(layer0_outputs[2732]) | (layer0_outputs[4867]);
    assign layer1_outputs[1646] = (layer0_outputs[2358]) & ~(layer0_outputs[3449]);
    assign layer1_outputs[1647] = ~(layer0_outputs[1129]);
    assign layer1_outputs[1648] = ~((layer0_outputs[1582]) & (layer0_outputs[3148]));
    assign layer1_outputs[1649] = ~(layer0_outputs[3720]);
    assign layer1_outputs[1650] = layer0_outputs[4372];
    assign layer1_outputs[1651] = (layer0_outputs[899]) & ~(layer0_outputs[1259]);
    assign layer1_outputs[1652] = layer0_outputs[4474];
    assign layer1_outputs[1653] = ~(layer0_outputs[3923]);
    assign layer1_outputs[1654] = ~(layer0_outputs[4477]);
    assign layer1_outputs[1655] = 1'b1;
    assign layer1_outputs[1656] = (layer0_outputs[1095]) & ~(layer0_outputs[472]);
    assign layer1_outputs[1657] = (layer0_outputs[5032]) & ~(layer0_outputs[4841]);
    assign layer1_outputs[1658] = (layer0_outputs[23]) & (layer0_outputs[1052]);
    assign layer1_outputs[1659] = ~(layer0_outputs[4896]);
    assign layer1_outputs[1660] = (layer0_outputs[4509]) ^ (layer0_outputs[1802]);
    assign layer1_outputs[1661] = (layer0_outputs[1849]) & (layer0_outputs[2324]);
    assign layer1_outputs[1662] = ~(layer0_outputs[2794]) | (layer0_outputs[2008]);
    assign layer1_outputs[1663] = ~(layer0_outputs[2895]) | (layer0_outputs[1179]);
    assign layer1_outputs[1664] = ~(layer0_outputs[1253]) | (layer0_outputs[2597]);
    assign layer1_outputs[1665] = (layer0_outputs[658]) & ~(layer0_outputs[686]);
    assign layer1_outputs[1666] = ~(layer0_outputs[4160]) | (layer0_outputs[4008]);
    assign layer1_outputs[1667] = (layer0_outputs[649]) & ~(layer0_outputs[2449]);
    assign layer1_outputs[1668] = (layer0_outputs[4211]) & (layer0_outputs[3583]);
    assign layer1_outputs[1669] = layer0_outputs[174];
    assign layer1_outputs[1670] = layer0_outputs[517];
    assign layer1_outputs[1671] = (layer0_outputs[4569]) & (layer0_outputs[2840]);
    assign layer1_outputs[1672] = (layer0_outputs[4380]) ^ (layer0_outputs[3771]);
    assign layer1_outputs[1673] = ~(layer0_outputs[2921]) | (layer0_outputs[1717]);
    assign layer1_outputs[1674] = ~((layer0_outputs[54]) | (layer0_outputs[2293]));
    assign layer1_outputs[1675] = ~(layer0_outputs[1375]) | (layer0_outputs[1127]);
    assign layer1_outputs[1676] = 1'b0;
    assign layer1_outputs[1677] = ~((layer0_outputs[1903]) | (layer0_outputs[68]));
    assign layer1_outputs[1678] = ~(layer0_outputs[3967]) | (layer0_outputs[813]);
    assign layer1_outputs[1679] = 1'b0;
    assign layer1_outputs[1680] = layer0_outputs[669];
    assign layer1_outputs[1681] = (layer0_outputs[2627]) & ~(layer0_outputs[4696]);
    assign layer1_outputs[1682] = ~(layer0_outputs[2875]);
    assign layer1_outputs[1683] = 1'b0;
    assign layer1_outputs[1684] = ~((layer0_outputs[1075]) | (layer0_outputs[2735]));
    assign layer1_outputs[1685] = 1'b1;
    assign layer1_outputs[1686] = ~(layer0_outputs[2042]) | (layer0_outputs[531]);
    assign layer1_outputs[1687] = ~(layer0_outputs[1009]) | (layer0_outputs[4258]);
    assign layer1_outputs[1688] = 1'b0;
    assign layer1_outputs[1689] = (layer0_outputs[5071]) & ~(layer0_outputs[547]);
    assign layer1_outputs[1690] = layer0_outputs[4930];
    assign layer1_outputs[1691] = ~((layer0_outputs[2273]) | (layer0_outputs[5037]));
    assign layer1_outputs[1692] = (layer0_outputs[1161]) & ~(layer0_outputs[207]);
    assign layer1_outputs[1693] = (layer0_outputs[3029]) & ~(layer0_outputs[3396]);
    assign layer1_outputs[1694] = 1'b0;
    assign layer1_outputs[1695] = ~((layer0_outputs[3071]) & (layer0_outputs[1352]));
    assign layer1_outputs[1696] = ~(layer0_outputs[655]) | (layer0_outputs[60]);
    assign layer1_outputs[1697] = ~(layer0_outputs[3796]);
    assign layer1_outputs[1698] = (layer0_outputs[3059]) & ~(layer0_outputs[3320]);
    assign layer1_outputs[1699] = ~(layer0_outputs[4652]);
    assign layer1_outputs[1700] = 1'b1;
    assign layer1_outputs[1701] = (layer0_outputs[3303]) & ~(layer0_outputs[1795]);
    assign layer1_outputs[1702] = layer0_outputs[1240];
    assign layer1_outputs[1703] = (layer0_outputs[4832]) & ~(layer0_outputs[1114]);
    assign layer1_outputs[1704] = ~(layer0_outputs[397]);
    assign layer1_outputs[1705] = ~(layer0_outputs[4317]) | (layer0_outputs[346]);
    assign layer1_outputs[1706] = layer0_outputs[4275];
    assign layer1_outputs[1707] = 1'b0;
    assign layer1_outputs[1708] = ~(layer0_outputs[3023]) | (layer0_outputs[4591]);
    assign layer1_outputs[1709] = (layer0_outputs[61]) & (layer0_outputs[3383]);
    assign layer1_outputs[1710] = (layer0_outputs[4638]) & ~(layer0_outputs[328]);
    assign layer1_outputs[1711] = ~((layer0_outputs[1942]) | (layer0_outputs[2899]));
    assign layer1_outputs[1712] = ~(layer0_outputs[853]) | (layer0_outputs[5069]);
    assign layer1_outputs[1713] = (layer0_outputs[899]) & ~(layer0_outputs[2033]);
    assign layer1_outputs[1714] = ~((layer0_outputs[944]) | (layer0_outputs[2852]));
    assign layer1_outputs[1715] = (layer0_outputs[3068]) & ~(layer0_outputs[735]);
    assign layer1_outputs[1716] = ~(layer0_outputs[2347]);
    assign layer1_outputs[1717] = ~(layer0_outputs[1527]) | (layer0_outputs[4375]);
    assign layer1_outputs[1718] = ~(layer0_outputs[4]) | (layer0_outputs[1495]);
    assign layer1_outputs[1719] = layer0_outputs[838];
    assign layer1_outputs[1720] = (layer0_outputs[4470]) & ~(layer0_outputs[1848]);
    assign layer1_outputs[1721] = (layer0_outputs[3448]) ^ (layer0_outputs[5018]);
    assign layer1_outputs[1722] = ~((layer0_outputs[1851]) & (layer0_outputs[2264]));
    assign layer1_outputs[1723] = ~(layer0_outputs[4640]) | (layer0_outputs[2265]);
    assign layer1_outputs[1724] = 1'b1;
    assign layer1_outputs[1725] = 1'b1;
    assign layer1_outputs[1726] = (layer0_outputs[803]) & (layer0_outputs[104]);
    assign layer1_outputs[1727] = 1'b0;
    assign layer1_outputs[1728] = 1'b1;
    assign layer1_outputs[1729] = (layer0_outputs[2638]) & ~(layer0_outputs[2953]);
    assign layer1_outputs[1730] = (layer0_outputs[5005]) & (layer0_outputs[4653]);
    assign layer1_outputs[1731] = 1'b1;
    assign layer1_outputs[1732] = ~(layer0_outputs[2024]);
    assign layer1_outputs[1733] = (layer0_outputs[5098]) | (layer0_outputs[4244]);
    assign layer1_outputs[1734] = 1'b0;
    assign layer1_outputs[1735] = 1'b0;
    assign layer1_outputs[1736] = 1'b0;
    assign layer1_outputs[1737] = layer0_outputs[5061];
    assign layer1_outputs[1738] = ~(layer0_outputs[3744]);
    assign layer1_outputs[1739] = (layer0_outputs[3671]) & (layer0_outputs[1490]);
    assign layer1_outputs[1740] = ~(layer0_outputs[2491]);
    assign layer1_outputs[1741] = layer0_outputs[20];
    assign layer1_outputs[1742] = (layer0_outputs[786]) | (layer0_outputs[2066]);
    assign layer1_outputs[1743] = ~(layer0_outputs[1196]) | (layer0_outputs[2297]);
    assign layer1_outputs[1744] = (layer0_outputs[464]) & ~(layer0_outputs[2367]);
    assign layer1_outputs[1745] = 1'b1;
    assign layer1_outputs[1746] = (layer0_outputs[1452]) & ~(layer0_outputs[565]);
    assign layer1_outputs[1747] = ~((layer0_outputs[2174]) | (layer0_outputs[4513]));
    assign layer1_outputs[1748] = (layer0_outputs[1242]) & ~(layer0_outputs[392]);
    assign layer1_outputs[1749] = layer0_outputs[2977];
    assign layer1_outputs[1750] = (layer0_outputs[3768]) & (layer0_outputs[1266]);
    assign layer1_outputs[1751] = ~(layer0_outputs[3911]) | (layer0_outputs[2960]);
    assign layer1_outputs[1752] = ~(layer0_outputs[3976]);
    assign layer1_outputs[1753] = 1'b1;
    assign layer1_outputs[1754] = (layer0_outputs[2463]) & (layer0_outputs[4615]);
    assign layer1_outputs[1755] = 1'b1;
    assign layer1_outputs[1756] = 1'b0;
    assign layer1_outputs[1757] = ~(layer0_outputs[710]) | (layer0_outputs[1072]);
    assign layer1_outputs[1758] = (layer0_outputs[4746]) & ~(layer0_outputs[1111]);
    assign layer1_outputs[1759] = layer0_outputs[224];
    assign layer1_outputs[1760] = ~((layer0_outputs[4270]) | (layer0_outputs[3107]));
    assign layer1_outputs[1761] = ~(layer0_outputs[1945]);
    assign layer1_outputs[1762] = 1'b0;
    assign layer1_outputs[1763] = (layer0_outputs[2613]) | (layer0_outputs[2385]);
    assign layer1_outputs[1764] = layer0_outputs[1643];
    assign layer1_outputs[1765] = ~(layer0_outputs[5036]) | (layer0_outputs[3824]);
    assign layer1_outputs[1766] = (layer0_outputs[272]) & ~(layer0_outputs[1464]);
    assign layer1_outputs[1767] = ~(layer0_outputs[4195]) | (layer0_outputs[2162]);
    assign layer1_outputs[1768] = (layer0_outputs[2759]) | (layer0_outputs[1040]);
    assign layer1_outputs[1769] = (layer0_outputs[3918]) & ~(layer0_outputs[3941]);
    assign layer1_outputs[1770] = layer0_outputs[4282];
    assign layer1_outputs[1771] = ~(layer0_outputs[2012]) | (layer0_outputs[1467]);
    assign layer1_outputs[1772] = layer0_outputs[3195];
    assign layer1_outputs[1773] = (layer0_outputs[531]) | (layer0_outputs[694]);
    assign layer1_outputs[1774] = ~(layer0_outputs[4807]) | (layer0_outputs[59]);
    assign layer1_outputs[1775] = ~(layer0_outputs[3496]);
    assign layer1_outputs[1776] = (layer0_outputs[3111]) | (layer0_outputs[2663]);
    assign layer1_outputs[1777] = 1'b0;
    assign layer1_outputs[1778] = (layer0_outputs[4439]) | (layer0_outputs[3736]);
    assign layer1_outputs[1779] = (layer0_outputs[428]) & ~(layer0_outputs[459]);
    assign layer1_outputs[1780] = ~(layer0_outputs[2610]);
    assign layer1_outputs[1781] = ~((layer0_outputs[2235]) & (layer0_outputs[1468]));
    assign layer1_outputs[1782] = ~(layer0_outputs[3984]) | (layer0_outputs[2151]);
    assign layer1_outputs[1783] = layer0_outputs[4485];
    assign layer1_outputs[1784] = ~(layer0_outputs[3908]) | (layer0_outputs[4385]);
    assign layer1_outputs[1785] = ~(layer0_outputs[2772]) | (layer0_outputs[3479]);
    assign layer1_outputs[1786] = 1'b1;
    assign layer1_outputs[1787] = 1'b1;
    assign layer1_outputs[1788] = (layer0_outputs[3431]) & ~(layer0_outputs[297]);
    assign layer1_outputs[1789] = ~(layer0_outputs[4824]);
    assign layer1_outputs[1790] = ~(layer0_outputs[2336]);
    assign layer1_outputs[1791] = layer0_outputs[1613];
    assign layer1_outputs[1792] = ~(layer0_outputs[4098]);
    assign layer1_outputs[1793] = layer0_outputs[848];
    assign layer1_outputs[1794] = ~(layer0_outputs[3474]);
    assign layer1_outputs[1795] = layer0_outputs[3250];
    assign layer1_outputs[1796] = ~(layer0_outputs[1969]);
    assign layer1_outputs[1797] = 1'b1;
    assign layer1_outputs[1798] = (layer0_outputs[4486]) ^ (layer0_outputs[4213]);
    assign layer1_outputs[1799] = ~(layer0_outputs[3059]);
    assign layer1_outputs[1800] = (layer0_outputs[3792]) & (layer0_outputs[5002]);
    assign layer1_outputs[1801] = (layer0_outputs[2550]) & ~(layer0_outputs[2]);
    assign layer1_outputs[1802] = layer0_outputs[3795];
    assign layer1_outputs[1803] = (layer0_outputs[1132]) & ~(layer0_outputs[3485]);
    assign layer1_outputs[1804] = ~((layer0_outputs[4472]) ^ (layer0_outputs[1338]));
    assign layer1_outputs[1805] = (layer0_outputs[927]) & ~(layer0_outputs[4398]);
    assign layer1_outputs[1806] = (layer0_outputs[243]) & ~(layer0_outputs[1544]);
    assign layer1_outputs[1807] = ~((layer0_outputs[2845]) & (layer0_outputs[2466]));
    assign layer1_outputs[1808] = (layer0_outputs[1552]) & ~(layer0_outputs[4347]);
    assign layer1_outputs[1809] = ~(layer0_outputs[1607]);
    assign layer1_outputs[1810] = (layer0_outputs[2494]) & (layer0_outputs[1978]);
    assign layer1_outputs[1811] = (layer0_outputs[3547]) & ~(layer0_outputs[1251]);
    assign layer1_outputs[1812] = 1'b0;
    assign layer1_outputs[1813] = (layer0_outputs[1931]) & ~(layer0_outputs[1380]);
    assign layer1_outputs[1814] = 1'b0;
    assign layer1_outputs[1815] = layer0_outputs[3496];
    assign layer1_outputs[1816] = layer0_outputs[2143];
    assign layer1_outputs[1817] = (layer0_outputs[1671]) & ~(layer0_outputs[925]);
    assign layer1_outputs[1818] = layer0_outputs[3077];
    assign layer1_outputs[1819] = ~(layer0_outputs[1779]);
    assign layer1_outputs[1820] = (layer0_outputs[4512]) ^ (layer0_outputs[4065]);
    assign layer1_outputs[1821] = (layer0_outputs[507]) ^ (layer0_outputs[3887]);
    assign layer1_outputs[1822] = ~((layer0_outputs[2119]) & (layer0_outputs[1888]));
    assign layer1_outputs[1823] = (layer0_outputs[3714]) & ~(layer0_outputs[3508]);
    assign layer1_outputs[1824] = ~(layer0_outputs[4017]);
    assign layer1_outputs[1825] = ~(layer0_outputs[2246]) | (layer0_outputs[1252]);
    assign layer1_outputs[1826] = ~((layer0_outputs[1243]) & (layer0_outputs[2943]));
    assign layer1_outputs[1827] = 1'b1;
    assign layer1_outputs[1828] = 1'b0;
    assign layer1_outputs[1829] = ~(layer0_outputs[3505]);
    assign layer1_outputs[1830] = (layer0_outputs[990]) & ~(layer0_outputs[2375]);
    assign layer1_outputs[1831] = layer0_outputs[2166];
    assign layer1_outputs[1832] = ~(layer0_outputs[1974]) | (layer0_outputs[3646]);
    assign layer1_outputs[1833] = layer0_outputs[3852];
    assign layer1_outputs[1834] = ~((layer0_outputs[2965]) ^ (layer0_outputs[3612]));
    assign layer1_outputs[1835] = 1'b1;
    assign layer1_outputs[1836] = layer0_outputs[1087];
    assign layer1_outputs[1837] = 1'b0;
    assign layer1_outputs[1838] = ~(layer0_outputs[2161]);
    assign layer1_outputs[1839] = (layer0_outputs[3078]) | (layer0_outputs[1730]);
    assign layer1_outputs[1840] = (layer0_outputs[3472]) & (layer0_outputs[909]);
    assign layer1_outputs[1841] = ~(layer0_outputs[3949]);
    assign layer1_outputs[1842] = (layer0_outputs[1664]) & ~(layer0_outputs[2927]);
    assign layer1_outputs[1843] = ~((layer0_outputs[268]) ^ (layer0_outputs[4039]));
    assign layer1_outputs[1844] = (layer0_outputs[3191]) ^ (layer0_outputs[1096]);
    assign layer1_outputs[1845] = 1'b1;
    assign layer1_outputs[1846] = 1'b0;
    assign layer1_outputs[1847] = (layer0_outputs[1655]) | (layer0_outputs[1487]);
    assign layer1_outputs[1848] = (layer0_outputs[3242]) & ~(layer0_outputs[2633]);
    assign layer1_outputs[1849] = 1'b0;
    assign layer1_outputs[1850] = layer0_outputs[3621];
    assign layer1_outputs[1851] = layer0_outputs[3601];
    assign layer1_outputs[1852] = ~((layer0_outputs[3569]) & (layer0_outputs[3443]));
    assign layer1_outputs[1853] = (layer0_outputs[917]) & ~(layer0_outputs[2102]);
    assign layer1_outputs[1854] = 1'b0;
    assign layer1_outputs[1855] = (layer0_outputs[3591]) & (layer0_outputs[112]);
    assign layer1_outputs[1856] = (layer0_outputs[4572]) & ~(layer0_outputs[1285]);
    assign layer1_outputs[1857] = ~(layer0_outputs[2065]);
    assign layer1_outputs[1858] = layer0_outputs[4637];
    assign layer1_outputs[1859] = ~(layer0_outputs[1596]);
    assign layer1_outputs[1860] = ~(layer0_outputs[4348]);
    assign layer1_outputs[1861] = layer0_outputs[3104];
    assign layer1_outputs[1862] = 1'b0;
    assign layer1_outputs[1863] = layer0_outputs[2236];
    assign layer1_outputs[1864] = 1'b0;
    assign layer1_outputs[1865] = (layer0_outputs[1812]) ^ (layer0_outputs[904]);
    assign layer1_outputs[1866] = (layer0_outputs[1235]) & ~(layer0_outputs[3116]);
    assign layer1_outputs[1867] = ~((layer0_outputs[3849]) ^ (layer0_outputs[2618]));
    assign layer1_outputs[1868] = 1'b0;
    assign layer1_outputs[1869] = layer0_outputs[2965];
    assign layer1_outputs[1870] = layer0_outputs[3965];
    assign layer1_outputs[1871] = layer0_outputs[47];
    assign layer1_outputs[1872] = 1'b1;
    assign layer1_outputs[1873] = ~((layer0_outputs[2403]) ^ (layer0_outputs[598]));
    assign layer1_outputs[1874] = (layer0_outputs[2618]) & (layer0_outputs[2897]);
    assign layer1_outputs[1875] = ~(layer0_outputs[5096]) | (layer0_outputs[2503]);
    assign layer1_outputs[1876] = ~((layer0_outputs[4746]) & (layer0_outputs[406]));
    assign layer1_outputs[1877] = (layer0_outputs[4806]) | (layer0_outputs[161]);
    assign layer1_outputs[1878] = (layer0_outputs[4992]) ^ (layer0_outputs[4005]);
    assign layer1_outputs[1879] = (layer0_outputs[621]) & (layer0_outputs[4276]);
    assign layer1_outputs[1880] = (layer0_outputs[2288]) & (layer0_outputs[2912]);
    assign layer1_outputs[1881] = 1'b0;
    assign layer1_outputs[1882] = (layer0_outputs[3874]) & (layer0_outputs[4635]);
    assign layer1_outputs[1883] = ~((layer0_outputs[2661]) | (layer0_outputs[882]));
    assign layer1_outputs[1884] = layer0_outputs[2314];
    assign layer1_outputs[1885] = (layer0_outputs[1855]) & ~(layer0_outputs[5098]);
    assign layer1_outputs[1886] = layer0_outputs[1493];
    assign layer1_outputs[1887] = ~(layer0_outputs[3030]);
    assign layer1_outputs[1888] = 1'b1;
    assign layer1_outputs[1889] = (layer0_outputs[2003]) & ~(layer0_outputs[4743]);
    assign layer1_outputs[1890] = (layer0_outputs[3440]) & ~(layer0_outputs[4728]);
    assign layer1_outputs[1891] = ~(layer0_outputs[937]) | (layer0_outputs[3946]);
    assign layer1_outputs[1892] = ~(layer0_outputs[1306]);
    assign layer1_outputs[1893] = 1'b1;
    assign layer1_outputs[1894] = ~(layer0_outputs[4494]);
    assign layer1_outputs[1895] = ~(layer0_outputs[3055]);
    assign layer1_outputs[1896] = 1'b1;
    assign layer1_outputs[1897] = ~((layer0_outputs[1709]) & (layer0_outputs[2450]));
    assign layer1_outputs[1898] = ~(layer0_outputs[2734]);
    assign layer1_outputs[1899] = (layer0_outputs[2209]) & (layer0_outputs[553]);
    assign layer1_outputs[1900] = (layer0_outputs[2924]) & ~(layer0_outputs[3526]);
    assign layer1_outputs[1901] = (layer0_outputs[159]) & (layer0_outputs[279]);
    assign layer1_outputs[1902] = ~(layer0_outputs[1630]);
    assign layer1_outputs[1903] = layer0_outputs[1480];
    assign layer1_outputs[1904] = ~(layer0_outputs[2339]);
    assign layer1_outputs[1905] = 1'b0;
    assign layer1_outputs[1906] = 1'b1;
    assign layer1_outputs[1907] = ~(layer0_outputs[1525]) | (layer0_outputs[1648]);
    assign layer1_outputs[1908] = ~(layer0_outputs[2507]) | (layer0_outputs[2228]);
    assign layer1_outputs[1909] = (layer0_outputs[3723]) & ~(layer0_outputs[1821]);
    assign layer1_outputs[1910] = (layer0_outputs[5034]) & (layer0_outputs[1263]);
    assign layer1_outputs[1911] = ~(layer0_outputs[2567]) | (layer0_outputs[3624]);
    assign layer1_outputs[1912] = 1'b1;
    assign layer1_outputs[1913] = (layer0_outputs[1626]) & ~(layer0_outputs[1783]);
    assign layer1_outputs[1914] = ~((layer0_outputs[2988]) ^ (layer0_outputs[3292]));
    assign layer1_outputs[1915] = ~((layer0_outputs[3377]) | (layer0_outputs[1280]));
    assign layer1_outputs[1916] = (layer0_outputs[1644]) & (layer0_outputs[2335]);
    assign layer1_outputs[1917] = ~(layer0_outputs[2106]) | (layer0_outputs[3137]);
    assign layer1_outputs[1918] = 1'b0;
    assign layer1_outputs[1919] = layer0_outputs[318];
    assign layer1_outputs[1920] = (layer0_outputs[2200]) & ~(layer0_outputs[1364]);
    assign layer1_outputs[1921] = ~((layer0_outputs[4708]) & (layer0_outputs[2146]));
    assign layer1_outputs[1922] = (layer0_outputs[1331]) | (layer0_outputs[3256]);
    assign layer1_outputs[1923] = (layer0_outputs[4969]) & ~(layer0_outputs[1385]);
    assign layer1_outputs[1924] = ~(layer0_outputs[4014]) | (layer0_outputs[4134]);
    assign layer1_outputs[1925] = ~(layer0_outputs[125]);
    assign layer1_outputs[1926] = (layer0_outputs[1414]) | (layer0_outputs[1478]);
    assign layer1_outputs[1927] = ~(layer0_outputs[446]) | (layer0_outputs[2803]);
    assign layer1_outputs[1928] = (layer0_outputs[4082]) & ~(layer0_outputs[1719]);
    assign layer1_outputs[1929] = 1'b1;
    assign layer1_outputs[1930] = ~(layer0_outputs[2276]) | (layer0_outputs[1522]);
    assign layer1_outputs[1931] = 1'b1;
    assign layer1_outputs[1932] = layer0_outputs[3720];
    assign layer1_outputs[1933] = 1'b1;
    assign layer1_outputs[1934] = (layer0_outputs[2508]) ^ (layer0_outputs[3781]);
    assign layer1_outputs[1935] = 1'b0;
    assign layer1_outputs[1936] = ~(layer0_outputs[470]) | (layer0_outputs[4193]);
    assign layer1_outputs[1937] = ~(layer0_outputs[1169]) | (layer0_outputs[1071]);
    assign layer1_outputs[1938] = 1'b1;
    assign layer1_outputs[1939] = ~(layer0_outputs[2479]) | (layer0_outputs[3007]);
    assign layer1_outputs[1940] = ~((layer0_outputs[4162]) & (layer0_outputs[4153]));
    assign layer1_outputs[1941] = (layer0_outputs[29]) & ~(layer0_outputs[2954]);
    assign layer1_outputs[1942] = ~((layer0_outputs[22]) | (layer0_outputs[498]));
    assign layer1_outputs[1943] = 1'b0;
    assign layer1_outputs[1944] = ~(layer0_outputs[5039]) | (layer0_outputs[3771]);
    assign layer1_outputs[1945] = ~(layer0_outputs[2585]);
    assign layer1_outputs[1946] = ~(layer0_outputs[103]);
    assign layer1_outputs[1947] = (layer0_outputs[3637]) & (layer0_outputs[442]);
    assign layer1_outputs[1948] = 1'b0;
    assign layer1_outputs[1949] = ~(layer0_outputs[4302]) | (layer0_outputs[5043]);
    assign layer1_outputs[1950] = ~(layer0_outputs[4905]) | (layer0_outputs[527]);
    assign layer1_outputs[1951] = 1'b0;
    assign layer1_outputs[1952] = (layer0_outputs[5105]) & (layer0_outputs[357]);
    assign layer1_outputs[1953] = ~((layer0_outputs[4183]) & (layer0_outputs[5067]));
    assign layer1_outputs[1954] = 1'b0;
    assign layer1_outputs[1955] = ~((layer0_outputs[2784]) & (layer0_outputs[1324]));
    assign layer1_outputs[1956] = (layer0_outputs[2340]) & ~(layer0_outputs[4060]);
    assign layer1_outputs[1957] = 1'b1;
    assign layer1_outputs[1958] = ~(layer0_outputs[1354]) | (layer0_outputs[4202]);
    assign layer1_outputs[1959] = (layer0_outputs[4107]) | (layer0_outputs[4833]);
    assign layer1_outputs[1960] = (layer0_outputs[1074]) & ~(layer0_outputs[212]);
    assign layer1_outputs[1961] = layer0_outputs[4075];
    assign layer1_outputs[1962] = ~(layer0_outputs[1678]) | (layer0_outputs[3835]);
    assign layer1_outputs[1963] = layer0_outputs[234];
    assign layer1_outputs[1964] = ~((layer0_outputs[4531]) & (layer0_outputs[3609]));
    assign layer1_outputs[1965] = (layer0_outputs[3483]) | (layer0_outputs[4653]);
    assign layer1_outputs[1966] = ~(layer0_outputs[3298]) | (layer0_outputs[149]);
    assign layer1_outputs[1967] = (layer0_outputs[3155]) & ~(layer0_outputs[2364]);
    assign layer1_outputs[1968] = ~(layer0_outputs[4626]) | (layer0_outputs[2996]);
    assign layer1_outputs[1969] = layer0_outputs[3426];
    assign layer1_outputs[1970] = 1'b1;
    assign layer1_outputs[1971] = ~((layer0_outputs[3443]) & (layer0_outputs[2817]));
    assign layer1_outputs[1972] = ~(layer0_outputs[3864]) | (layer0_outputs[627]);
    assign layer1_outputs[1973] = ~(layer0_outputs[1809]);
    assign layer1_outputs[1974] = ~(layer0_outputs[2069]);
    assign layer1_outputs[1975] = (layer0_outputs[2416]) & (layer0_outputs[2733]);
    assign layer1_outputs[1976] = layer0_outputs[1188];
    assign layer1_outputs[1977] = (layer0_outputs[3691]) ^ (layer0_outputs[2019]);
    assign layer1_outputs[1978] = (layer0_outputs[4870]) & ~(layer0_outputs[784]);
    assign layer1_outputs[1979] = ~(layer0_outputs[2823]) | (layer0_outputs[1966]);
    assign layer1_outputs[1980] = layer0_outputs[3229];
    assign layer1_outputs[1981] = ~((layer0_outputs[3850]) ^ (layer0_outputs[2061]));
    assign layer1_outputs[1982] = ~(layer0_outputs[1459]) | (layer0_outputs[1344]);
    assign layer1_outputs[1983] = 1'b0;
    assign layer1_outputs[1984] = 1'b0;
    assign layer1_outputs[1985] = (layer0_outputs[3776]) | (layer0_outputs[3403]);
    assign layer1_outputs[1986] = layer0_outputs[4211];
    assign layer1_outputs[1987] = ~((layer0_outputs[2995]) & (layer0_outputs[4924]));
    assign layer1_outputs[1988] = layer0_outputs[3193];
    assign layer1_outputs[1989] = layer0_outputs[4248];
    assign layer1_outputs[1990] = layer0_outputs[1862];
    assign layer1_outputs[1991] = ~(layer0_outputs[1978]) | (layer0_outputs[3667]);
    assign layer1_outputs[1992] = ~((layer0_outputs[2594]) & (layer0_outputs[1224]));
    assign layer1_outputs[1993] = ~(layer0_outputs[830]) | (layer0_outputs[1290]);
    assign layer1_outputs[1994] = 1'b0;
    assign layer1_outputs[1995] = layer0_outputs[472];
    assign layer1_outputs[1996] = ~(layer0_outputs[4673]) | (layer0_outputs[3955]);
    assign layer1_outputs[1997] = ~((layer0_outputs[1871]) | (layer0_outputs[2337]));
    assign layer1_outputs[1998] = ~(layer0_outputs[35]) | (layer0_outputs[2987]);
    assign layer1_outputs[1999] = (layer0_outputs[1197]) & ~(layer0_outputs[609]);
    assign layer1_outputs[2000] = layer0_outputs[46];
    assign layer1_outputs[2001] = (layer0_outputs[2698]) & ~(layer0_outputs[5078]);
    assign layer1_outputs[2002] = 1'b0;
    assign layer1_outputs[2003] = layer0_outputs[630];
    assign layer1_outputs[2004] = ~((layer0_outputs[3302]) & (layer0_outputs[1930]));
    assign layer1_outputs[2005] = (layer0_outputs[4587]) & ~(layer0_outputs[2336]);
    assign layer1_outputs[2006] = (layer0_outputs[3669]) & ~(layer0_outputs[3259]);
    assign layer1_outputs[2007] = (layer0_outputs[1177]) & ~(layer0_outputs[9]);
    assign layer1_outputs[2008] = 1'b1;
    assign layer1_outputs[2009] = 1'b1;
    assign layer1_outputs[2010] = layer0_outputs[3629];
    assign layer1_outputs[2011] = ~(layer0_outputs[4569]);
    assign layer1_outputs[2012] = 1'b0;
    assign layer1_outputs[2013] = (layer0_outputs[1236]) & ~(layer0_outputs[3346]);
    assign layer1_outputs[2014] = ~((layer0_outputs[3703]) & (layer0_outputs[4736]));
    assign layer1_outputs[2015] = layer0_outputs[1549];
    assign layer1_outputs[2016] = (layer0_outputs[4235]) & (layer0_outputs[2978]);
    assign layer1_outputs[2017] = (layer0_outputs[203]) & ~(layer0_outputs[1451]);
    assign layer1_outputs[2018] = ~(layer0_outputs[4783]);
    assign layer1_outputs[2019] = 1'b1;
    assign layer1_outputs[2020] = ~((layer0_outputs[626]) & (layer0_outputs[131]));
    assign layer1_outputs[2021] = (layer0_outputs[3660]) | (layer0_outputs[2707]);
    assign layer1_outputs[2022] = 1'b1;
    assign layer1_outputs[2023] = (layer0_outputs[567]) & ~(layer0_outputs[805]);
    assign layer1_outputs[2024] = ~((layer0_outputs[724]) & (layer0_outputs[3824]));
    assign layer1_outputs[2025] = ~(layer0_outputs[4233]);
    assign layer1_outputs[2026] = ~(layer0_outputs[682]);
    assign layer1_outputs[2027] = layer0_outputs[1474];
    assign layer1_outputs[2028] = (layer0_outputs[1438]) & ~(layer0_outputs[3919]);
    assign layer1_outputs[2029] = ~((layer0_outputs[1597]) | (layer0_outputs[1655]));
    assign layer1_outputs[2030] = ~(layer0_outputs[590]) | (layer0_outputs[2348]);
    assign layer1_outputs[2031] = 1'b1;
    assign layer1_outputs[2032] = 1'b1;
    assign layer1_outputs[2033] = 1'b0;
    assign layer1_outputs[2034] = ~((layer0_outputs[256]) | (layer0_outputs[278]));
    assign layer1_outputs[2035] = (layer0_outputs[2343]) | (layer0_outputs[4877]);
    assign layer1_outputs[2036] = ~(layer0_outputs[1929]);
    assign layer1_outputs[2037] = (layer0_outputs[3417]) & (layer0_outputs[3456]);
    assign layer1_outputs[2038] = (layer0_outputs[2848]) & ~(layer0_outputs[4197]);
    assign layer1_outputs[2039] = ~(layer0_outputs[5028]) | (layer0_outputs[1921]);
    assign layer1_outputs[2040] = ~((layer0_outputs[2230]) | (layer0_outputs[1495]));
    assign layer1_outputs[2041] = (layer0_outputs[4685]) & ~(layer0_outputs[5063]);
    assign layer1_outputs[2042] = 1'b1;
    assign layer1_outputs[2043] = ~((layer0_outputs[2440]) | (layer0_outputs[2915]));
    assign layer1_outputs[2044] = (layer0_outputs[3460]) & ~(layer0_outputs[2829]);
    assign layer1_outputs[2045] = ~(layer0_outputs[871]);
    assign layer1_outputs[2046] = ~((layer0_outputs[4687]) | (layer0_outputs[226]));
    assign layer1_outputs[2047] = ~((layer0_outputs[4341]) & (layer0_outputs[2945]));
    assign layer1_outputs[2048] = (layer0_outputs[1600]) & (layer0_outputs[4953]);
    assign layer1_outputs[2049] = (layer0_outputs[4289]) ^ (layer0_outputs[1733]);
    assign layer1_outputs[2050] = ~(layer0_outputs[4431]) | (layer0_outputs[918]);
    assign layer1_outputs[2051] = ~((layer0_outputs[1774]) | (layer0_outputs[3603]));
    assign layer1_outputs[2052] = layer0_outputs[4237];
    assign layer1_outputs[2053] = 1'b1;
    assign layer1_outputs[2054] = layer0_outputs[5003];
    assign layer1_outputs[2055] = 1'b1;
    assign layer1_outputs[2056] = 1'b1;
    assign layer1_outputs[2057] = (layer0_outputs[2813]) & ~(layer0_outputs[4719]);
    assign layer1_outputs[2058] = layer0_outputs[1223];
    assign layer1_outputs[2059] = (layer0_outputs[3988]) & ~(layer0_outputs[3157]);
    assign layer1_outputs[2060] = 1'b1;
    assign layer1_outputs[2061] = ~(layer0_outputs[2010]);
    assign layer1_outputs[2062] = (layer0_outputs[4333]) & (layer0_outputs[251]);
    assign layer1_outputs[2063] = ~(layer0_outputs[4925]) | (layer0_outputs[208]);
    assign layer1_outputs[2064] = ~((layer0_outputs[1098]) & (layer0_outputs[3702]));
    assign layer1_outputs[2065] = ~((layer0_outputs[681]) ^ (layer0_outputs[2654]));
    assign layer1_outputs[2066] = (layer0_outputs[129]) & ~(layer0_outputs[3855]);
    assign layer1_outputs[2067] = ~((layer0_outputs[1765]) ^ (layer0_outputs[4610]));
    assign layer1_outputs[2068] = ~((layer0_outputs[2496]) | (layer0_outputs[246]));
    assign layer1_outputs[2069] = ~((layer0_outputs[2741]) ^ (layer0_outputs[847]));
    assign layer1_outputs[2070] = 1'b0;
    assign layer1_outputs[2071] = (layer0_outputs[2796]) & (layer0_outputs[673]);
    assign layer1_outputs[2072] = ~((layer0_outputs[3411]) | (layer0_outputs[2517]));
    assign layer1_outputs[2073] = ~((layer0_outputs[825]) & (layer0_outputs[2122]));
    assign layer1_outputs[2074] = ~((layer0_outputs[804]) & (layer0_outputs[4463]));
    assign layer1_outputs[2075] = 1'b1;
    assign layer1_outputs[2076] = 1'b1;
    assign layer1_outputs[2077] = 1'b0;
    assign layer1_outputs[2078] = ~(layer0_outputs[2392]);
    assign layer1_outputs[2079] = 1'b1;
    assign layer1_outputs[2080] = ~((layer0_outputs[3511]) | (layer0_outputs[793]));
    assign layer1_outputs[2081] = layer0_outputs[213];
    assign layer1_outputs[2082] = ~(layer0_outputs[4270]) | (layer0_outputs[2584]);
    assign layer1_outputs[2083] = (layer0_outputs[167]) & (layer0_outputs[2552]);
    assign layer1_outputs[2084] = layer0_outputs[140];
    assign layer1_outputs[2085] = ~(layer0_outputs[4965]);
    assign layer1_outputs[2086] = 1'b1;
    assign layer1_outputs[2087] = (layer0_outputs[5014]) & ~(layer0_outputs[2630]);
    assign layer1_outputs[2088] = layer0_outputs[962];
    assign layer1_outputs[2089] = 1'b0;
    assign layer1_outputs[2090] = ~(layer0_outputs[3897]) | (layer0_outputs[2223]);
    assign layer1_outputs[2091] = ~(layer0_outputs[817]);
    assign layer1_outputs[2092] = layer0_outputs[1393];
    assign layer1_outputs[2093] = ~(layer0_outputs[386]);
    assign layer1_outputs[2094] = ~(layer0_outputs[3920]) | (layer0_outputs[3043]);
    assign layer1_outputs[2095] = 1'b0;
    assign layer1_outputs[2096] = 1'b0;
    assign layer1_outputs[2097] = layer0_outputs[3036];
    assign layer1_outputs[2098] = ~(layer0_outputs[2404]) | (layer0_outputs[1352]);
    assign layer1_outputs[2099] = ~(layer0_outputs[3687]);
    assign layer1_outputs[2100] = ~((layer0_outputs[2299]) & (layer0_outputs[3311]));
    assign layer1_outputs[2101] = (layer0_outputs[2082]) ^ (layer0_outputs[3654]);
    assign layer1_outputs[2102] = ~(layer0_outputs[3970]) | (layer0_outputs[1761]);
    assign layer1_outputs[2103] = ~(layer0_outputs[2368]);
    assign layer1_outputs[2104] = (layer0_outputs[639]) | (layer0_outputs[4053]);
    assign layer1_outputs[2105] = layer0_outputs[2546];
    assign layer1_outputs[2106] = ~((layer0_outputs[768]) | (layer0_outputs[586]));
    assign layer1_outputs[2107] = layer0_outputs[1760];
    assign layer1_outputs[2108] = ~(layer0_outputs[2757]);
    assign layer1_outputs[2109] = ~(layer0_outputs[1893]) | (layer0_outputs[1405]);
    assign layer1_outputs[2110] = (layer0_outputs[3710]) & ~(layer0_outputs[1804]);
    assign layer1_outputs[2111] = (layer0_outputs[118]) | (layer0_outputs[4487]);
    assign layer1_outputs[2112] = ~((layer0_outputs[2699]) & (layer0_outputs[946]));
    assign layer1_outputs[2113] = ~(layer0_outputs[774]);
    assign layer1_outputs[2114] = ~((layer0_outputs[3512]) & (layer0_outputs[3730]));
    assign layer1_outputs[2115] = 1'b1;
    assign layer1_outputs[2116] = ~((layer0_outputs[4116]) & (layer0_outputs[2944]));
    assign layer1_outputs[2117] = ~(layer0_outputs[1472]) | (layer0_outputs[1297]);
    assign layer1_outputs[2118] = ~((layer0_outputs[1782]) | (layer0_outputs[2192]));
    assign layer1_outputs[2119] = ~((layer0_outputs[4894]) | (layer0_outputs[1051]));
    assign layer1_outputs[2120] = (layer0_outputs[1066]) & ~(layer0_outputs[3998]);
    assign layer1_outputs[2121] = ~(layer0_outputs[1102]) | (layer0_outputs[2018]);
    assign layer1_outputs[2122] = ~(layer0_outputs[3725]);
    assign layer1_outputs[2123] = (layer0_outputs[3616]) | (layer0_outputs[2513]);
    assign layer1_outputs[2124] = ~((layer0_outputs[4207]) & (layer0_outputs[3750]));
    assign layer1_outputs[2125] = ~(layer0_outputs[4691]) | (layer0_outputs[670]);
    assign layer1_outputs[2126] = (layer0_outputs[604]) ^ (layer0_outputs[2939]);
    assign layer1_outputs[2127] = (layer0_outputs[3981]) | (layer0_outputs[789]);
    assign layer1_outputs[2128] = layer0_outputs[2199];
    assign layer1_outputs[2129] = layer0_outputs[2178];
    assign layer1_outputs[2130] = ~(layer0_outputs[4658]);
    assign layer1_outputs[2131] = 1'b0;
    assign layer1_outputs[2132] = layer0_outputs[445];
    assign layer1_outputs[2133] = layer0_outputs[3194];
    assign layer1_outputs[2134] = ~(layer0_outputs[1990]);
    assign layer1_outputs[2135] = ~(layer0_outputs[2784]) | (layer0_outputs[648]);
    assign layer1_outputs[2136] = 1'b1;
    assign layer1_outputs[2137] = ~(layer0_outputs[2556]) | (layer0_outputs[5049]);
    assign layer1_outputs[2138] = 1'b1;
    assign layer1_outputs[2139] = (layer0_outputs[1461]) | (layer0_outputs[4047]);
    assign layer1_outputs[2140] = ~((layer0_outputs[3495]) | (layer0_outputs[505]));
    assign layer1_outputs[2141] = 1'b1;
    assign layer1_outputs[2142] = layer0_outputs[871];
    assign layer1_outputs[2143] = layer0_outputs[707];
    assign layer1_outputs[2144] = ~(layer0_outputs[3533]) | (layer0_outputs[423]);
    assign layer1_outputs[2145] = 1'b0;
    assign layer1_outputs[2146] = 1'b1;
    assign layer1_outputs[2147] = layer0_outputs[3385];
    assign layer1_outputs[2148] = (layer0_outputs[2739]) ^ (layer0_outputs[769]);
    assign layer1_outputs[2149] = ~(layer0_outputs[4287]) | (layer0_outputs[4038]);
    assign layer1_outputs[2150] = 1'b1;
    assign layer1_outputs[2151] = ~(layer0_outputs[4774]);
    assign layer1_outputs[2152] = ~(layer0_outputs[3643]);
    assign layer1_outputs[2153] = ~((layer0_outputs[1875]) & (layer0_outputs[460]));
    assign layer1_outputs[2154] = (layer0_outputs[4913]) & ~(layer0_outputs[4092]);
    assign layer1_outputs[2155] = (layer0_outputs[4959]) ^ (layer0_outputs[4770]);
    assign layer1_outputs[2156] = ~(layer0_outputs[753]) | (layer0_outputs[2752]);
    assign layer1_outputs[2157] = (layer0_outputs[3394]) & ~(layer0_outputs[2307]);
    assign layer1_outputs[2158] = ~(layer0_outputs[3721]);
    assign layer1_outputs[2159] = ~(layer0_outputs[5007]) | (layer0_outputs[4989]);
    assign layer1_outputs[2160] = ~(layer0_outputs[281]);
    assign layer1_outputs[2161] = ~(layer0_outputs[707]);
    assign layer1_outputs[2162] = ~((layer0_outputs[4724]) & (layer0_outputs[2181]));
    assign layer1_outputs[2163] = ~((layer0_outputs[108]) & (layer0_outputs[4424]));
    assign layer1_outputs[2164] = ~((layer0_outputs[2241]) | (layer0_outputs[287]));
    assign layer1_outputs[2165] = 1'b0;
    assign layer1_outputs[2166] = (layer0_outputs[777]) & ~(layer0_outputs[1199]);
    assign layer1_outputs[2167] = (layer0_outputs[2716]) & ~(layer0_outputs[4938]);
    assign layer1_outputs[2168] = ~(layer0_outputs[18]) | (layer0_outputs[2642]);
    assign layer1_outputs[2169] = ~(layer0_outputs[229]);
    assign layer1_outputs[2170] = 1'b0;
    assign layer1_outputs[2171] = (layer0_outputs[4564]) | (layer0_outputs[2779]);
    assign layer1_outputs[2172] = ~(layer0_outputs[78]) | (layer0_outputs[3]);
    assign layer1_outputs[2173] = ~((layer0_outputs[2281]) | (layer0_outputs[2429]));
    assign layer1_outputs[2174] = ~(layer0_outputs[1268]) | (layer0_outputs[4552]);
    assign layer1_outputs[2175] = ~((layer0_outputs[4644]) & (layer0_outputs[1582]));
    assign layer1_outputs[2176] = ~((layer0_outputs[1217]) & (layer0_outputs[1742]));
    assign layer1_outputs[2177] = (layer0_outputs[4384]) & ~(layer0_outputs[3582]);
    assign layer1_outputs[2178] = (layer0_outputs[3683]) & ~(layer0_outputs[4407]);
    assign layer1_outputs[2179] = (layer0_outputs[943]) & (layer0_outputs[2489]);
    assign layer1_outputs[2180] = ~(layer0_outputs[863]);
    assign layer1_outputs[2181] = (layer0_outputs[22]) ^ (layer0_outputs[4992]);
    assign layer1_outputs[2182] = ~(layer0_outputs[3477]);
    assign layer1_outputs[2183] = ~(layer0_outputs[168]) | (layer0_outputs[750]);
    assign layer1_outputs[2184] = (layer0_outputs[916]) | (layer0_outputs[2865]);
    assign layer1_outputs[2185] = (layer0_outputs[2502]) & ~(layer0_outputs[3322]);
    assign layer1_outputs[2186] = (layer0_outputs[3990]) & ~(layer0_outputs[2576]);
    assign layer1_outputs[2187] = ~(layer0_outputs[876]) | (layer0_outputs[911]);
    assign layer1_outputs[2188] = layer0_outputs[2849];
    assign layer1_outputs[2189] = (layer0_outputs[1935]) & (layer0_outputs[969]);
    assign layer1_outputs[2190] = ~(layer0_outputs[4577]) | (layer0_outputs[4961]);
    assign layer1_outputs[2191] = 1'b1;
    assign layer1_outputs[2192] = layer0_outputs[3434];
    assign layer1_outputs[2193] = 1'b0;
    assign layer1_outputs[2194] = ~(layer0_outputs[2826]) | (layer0_outputs[1261]);
    assign layer1_outputs[2195] = ~(layer0_outputs[2598]) | (layer0_outputs[3953]);
    assign layer1_outputs[2196] = ~((layer0_outputs[5048]) & (layer0_outputs[1764]));
    assign layer1_outputs[2197] = ~((layer0_outputs[1712]) ^ (layer0_outputs[2547]));
    assign layer1_outputs[2198] = 1'b1;
    assign layer1_outputs[2199] = 1'b0;
    assign layer1_outputs[2200] = ~(layer0_outputs[3008]) | (layer0_outputs[153]);
    assign layer1_outputs[2201] = ~(layer0_outputs[722]) | (layer0_outputs[4865]);
    assign layer1_outputs[2202] = (layer0_outputs[3915]) | (layer0_outputs[2726]);
    assign layer1_outputs[2203] = 1'b0;
    assign layer1_outputs[2204] = ~((layer0_outputs[4892]) & (layer0_outputs[1208]));
    assign layer1_outputs[2205] = 1'b1;
    assign layer1_outputs[2206] = (layer0_outputs[1546]) & (layer0_outputs[593]);
    assign layer1_outputs[2207] = (layer0_outputs[5046]) & ~(layer0_outputs[2686]);
    assign layer1_outputs[2208] = 1'b1;
    assign layer1_outputs[2209] = ~(layer0_outputs[3365]) | (layer0_outputs[4489]);
    assign layer1_outputs[2210] = layer0_outputs[1850];
    assign layer1_outputs[2211] = ~((layer0_outputs[1680]) & (layer0_outputs[2300]));
    assign layer1_outputs[2212] = (layer0_outputs[2554]) | (layer0_outputs[152]);
    assign layer1_outputs[2213] = ~(layer0_outputs[887]) | (layer0_outputs[5085]);
    assign layer1_outputs[2214] = ~(layer0_outputs[1680]) | (layer0_outputs[4221]);
    assign layer1_outputs[2215] = (layer0_outputs[2707]) | (layer0_outputs[4138]);
    assign layer1_outputs[2216] = 1'b0;
    assign layer1_outputs[2217] = ~((layer0_outputs[4030]) & (layer0_outputs[400]));
    assign layer1_outputs[2218] = ~((layer0_outputs[5095]) | (layer0_outputs[4627]));
    assign layer1_outputs[2219] = 1'b0;
    assign layer1_outputs[2220] = ~(layer0_outputs[1178]);
    assign layer1_outputs[2221] = ~(layer0_outputs[585]);
    assign layer1_outputs[2222] = (layer0_outputs[2923]) & ~(layer0_outputs[4277]);
    assign layer1_outputs[2223] = ~(layer0_outputs[1080]);
    assign layer1_outputs[2224] = (layer0_outputs[2846]) & ~(layer0_outputs[1993]);
    assign layer1_outputs[2225] = (layer0_outputs[1005]) & ~(layer0_outputs[4229]);
    assign layer1_outputs[2226] = layer0_outputs[2957];
    assign layer1_outputs[2227] = (layer0_outputs[4784]) & ~(layer0_outputs[483]);
    assign layer1_outputs[2228] = ~((layer0_outputs[1588]) & (layer0_outputs[1108]));
    assign layer1_outputs[2229] = 1'b0;
    assign layer1_outputs[2230] = ~(layer0_outputs[4517]) | (layer0_outputs[1498]);
    assign layer1_outputs[2231] = ~(layer0_outputs[4711]) | (layer0_outputs[3906]);
    assign layer1_outputs[2232] = 1'b0;
    assign layer1_outputs[2233] = (layer0_outputs[2848]) & ~(layer0_outputs[591]);
    assign layer1_outputs[2234] = 1'b1;
    assign layer1_outputs[2235] = ~((layer0_outputs[1290]) | (layer0_outputs[2988]));
    assign layer1_outputs[2236] = ~((layer0_outputs[3288]) | (layer0_outputs[2243]));
    assign layer1_outputs[2237] = (layer0_outputs[2391]) & ~(layer0_outputs[1272]);
    assign layer1_outputs[2238] = 1'b0;
    assign layer1_outputs[2239] = 1'b0;
    assign layer1_outputs[2240] = 1'b0;
    assign layer1_outputs[2241] = ~(layer0_outputs[3182]);
    assign layer1_outputs[2242] = (layer0_outputs[4507]) & (layer0_outputs[3385]);
    assign layer1_outputs[2243] = ~((layer0_outputs[4055]) & (layer0_outputs[1275]));
    assign layer1_outputs[2244] = layer0_outputs[3940];
    assign layer1_outputs[2245] = 1'b0;
    assign layer1_outputs[2246] = ~((layer0_outputs[3296]) | (layer0_outputs[948]));
    assign layer1_outputs[2247] = ~(layer0_outputs[4073]) | (layer0_outputs[3498]);
    assign layer1_outputs[2248] = (layer0_outputs[2920]) & (layer0_outputs[2500]);
    assign layer1_outputs[2249] = ~(layer0_outputs[2097]) | (layer0_outputs[3210]);
    assign layer1_outputs[2250] = 1'b1;
    assign layer1_outputs[2251] = layer0_outputs[3563];
    assign layer1_outputs[2252] = ~((layer0_outputs[478]) | (layer0_outputs[4904]));
    assign layer1_outputs[2253] = ~((layer0_outputs[2346]) & (layer0_outputs[1053]));
    assign layer1_outputs[2254] = layer0_outputs[3934];
    assign layer1_outputs[2255] = layer0_outputs[4208];
    assign layer1_outputs[2256] = ~((layer0_outputs[3251]) | (layer0_outputs[1322]));
    assign layer1_outputs[2257] = (layer0_outputs[1952]) & ~(layer0_outputs[113]);
    assign layer1_outputs[2258] = (layer0_outputs[1835]) | (layer0_outputs[4800]);
    assign layer1_outputs[2259] = ~((layer0_outputs[3481]) | (layer0_outputs[1567]));
    assign layer1_outputs[2260] = (layer0_outputs[4559]) | (layer0_outputs[4037]);
    assign layer1_outputs[2261] = ~((layer0_outputs[2413]) | (layer0_outputs[4440]));
    assign layer1_outputs[2262] = (layer0_outputs[1778]) & ~(layer0_outputs[4798]);
    assign layer1_outputs[2263] = layer0_outputs[2141];
    assign layer1_outputs[2264] = (layer0_outputs[3746]) & ~(layer0_outputs[4238]);
    assign layer1_outputs[2265] = layer0_outputs[3285];
    assign layer1_outputs[2266] = ~(layer0_outputs[3658]) | (layer0_outputs[2481]);
    assign layer1_outputs[2267] = ~((layer0_outputs[4373]) ^ (layer0_outputs[4769]));
    assign layer1_outputs[2268] = ~(layer0_outputs[941]);
    assign layer1_outputs[2269] = ~((layer0_outputs[1347]) & (layer0_outputs[1912]));
    assign layer1_outputs[2270] = ~(layer0_outputs[646]) | (layer0_outputs[1124]);
    assign layer1_outputs[2271] = (layer0_outputs[4452]) & ~(layer0_outputs[920]);
    assign layer1_outputs[2272] = 1'b1;
    assign layer1_outputs[2273] = (layer0_outputs[3852]) & ~(layer0_outputs[1131]);
    assign layer1_outputs[2274] = ~((layer0_outputs[1870]) | (layer0_outputs[1995]));
    assign layer1_outputs[2275] = ~((layer0_outputs[3599]) ^ (layer0_outputs[1442]));
    assign layer1_outputs[2276] = ~(layer0_outputs[5076]);
    assign layer1_outputs[2277] = (layer0_outputs[1263]) & (layer0_outputs[4603]);
    assign layer1_outputs[2278] = 1'b1;
    assign layer1_outputs[2279] = ~(layer0_outputs[4257]) | (layer0_outputs[4523]);
    assign layer1_outputs[2280] = ~(layer0_outputs[981]) | (layer0_outputs[4876]);
    assign layer1_outputs[2281] = layer0_outputs[928];
    assign layer1_outputs[2282] = layer0_outputs[4279];
    assign layer1_outputs[2283] = ~(layer0_outputs[1769]);
    assign layer1_outputs[2284] = ~(layer0_outputs[4807]);
    assign layer1_outputs[2285] = (layer0_outputs[4739]) & (layer0_outputs[856]);
    assign layer1_outputs[2286] = 1'b1;
    assign layer1_outputs[2287] = (layer0_outputs[2909]) & ~(layer0_outputs[2250]);
    assign layer1_outputs[2288] = ~(layer0_outputs[2551]);
    assign layer1_outputs[2289] = ~(layer0_outputs[1797]);
    assign layer1_outputs[2290] = (layer0_outputs[5068]) & ~(layer0_outputs[1367]);
    assign layer1_outputs[2291] = ~(layer0_outputs[3943]) | (layer0_outputs[698]);
    assign layer1_outputs[2292] = (layer0_outputs[233]) | (layer0_outputs[45]);
    assign layer1_outputs[2293] = layer0_outputs[3831];
    assign layer1_outputs[2294] = ~(layer0_outputs[1209]);
    assign layer1_outputs[2295] = ~(layer0_outputs[4980]) | (layer0_outputs[2513]);
    assign layer1_outputs[2296] = ~(layer0_outputs[1239]);
    assign layer1_outputs[2297] = layer0_outputs[908];
    assign layer1_outputs[2298] = ~(layer0_outputs[2620]);
    assign layer1_outputs[2299] = ~((layer0_outputs[2045]) ^ (layer0_outputs[2482]));
    assign layer1_outputs[2300] = (layer0_outputs[3985]) & (layer0_outputs[4522]);
    assign layer1_outputs[2301] = 1'b0;
    assign layer1_outputs[2302] = ~((layer0_outputs[4178]) | (layer0_outputs[3190]));
    assign layer1_outputs[2303] = (layer0_outputs[2025]) & ~(layer0_outputs[1861]);
    assign layer1_outputs[2304] = 1'b0;
    assign layer1_outputs[2305] = layer0_outputs[4001];
    assign layer1_outputs[2306] = ~((layer0_outputs[3580]) & (layer0_outputs[4340]));
    assign layer1_outputs[2307] = (layer0_outputs[3395]) ^ (layer0_outputs[1430]);
    assign layer1_outputs[2308] = 1'b0;
    assign layer1_outputs[2309] = ~(layer0_outputs[3661]);
    assign layer1_outputs[2310] = (layer0_outputs[3436]) & ~(layer0_outputs[3065]);
    assign layer1_outputs[2311] = 1'b0;
    assign layer1_outputs[2312] = (layer0_outputs[4166]) & ~(layer0_outputs[3267]);
    assign layer1_outputs[2313] = (layer0_outputs[1328]) | (layer0_outputs[4869]);
    assign layer1_outputs[2314] = ~((layer0_outputs[2951]) & (layer0_outputs[3194]));
    assign layer1_outputs[2315] = (layer0_outputs[815]) & ~(layer0_outputs[2566]);
    assign layer1_outputs[2316] = ~((layer0_outputs[2278]) & (layer0_outputs[543]));
    assign layer1_outputs[2317] = (layer0_outputs[1112]) & (layer0_outputs[4718]);
    assign layer1_outputs[2318] = layer0_outputs[4444];
    assign layer1_outputs[2319] = (layer0_outputs[3053]) & (layer0_outputs[253]);
    assign layer1_outputs[2320] = ~((layer0_outputs[2358]) & (layer0_outputs[4367]));
    assign layer1_outputs[2321] = 1'b0;
    assign layer1_outputs[2322] = ~((layer0_outputs[4771]) | (layer0_outputs[3348]));
    assign layer1_outputs[2323] = ~(layer0_outputs[1997]) | (layer0_outputs[1216]);
    assign layer1_outputs[2324] = layer0_outputs[1156];
    assign layer1_outputs[2325] = ~(layer0_outputs[2717]) | (layer0_outputs[4028]);
    assign layer1_outputs[2326] = ~((layer0_outputs[3961]) | (layer0_outputs[1074]));
    assign layer1_outputs[2327] = 1'b0;
    assign layer1_outputs[2328] = ~((layer0_outputs[4975]) & (layer0_outputs[1858]));
    assign layer1_outputs[2329] = layer0_outputs[4216];
    assign layer1_outputs[2330] = (layer0_outputs[1084]) & ~(layer0_outputs[2810]);
    assign layer1_outputs[2331] = (layer0_outputs[4131]) & ~(layer0_outputs[1778]);
    assign layer1_outputs[2332] = ~(layer0_outputs[4991]);
    assign layer1_outputs[2333] = layer0_outputs[2161];
    assign layer1_outputs[2334] = (layer0_outputs[1636]) & (layer0_outputs[288]);
    assign layer1_outputs[2335] = (layer0_outputs[1203]) & ~(layer0_outputs[3748]);
    assign layer1_outputs[2336] = 1'b0;
    assign layer1_outputs[2337] = 1'b1;
    assign layer1_outputs[2338] = 1'b1;
    assign layer1_outputs[2339] = (layer0_outputs[2425]) & (layer0_outputs[38]);
    assign layer1_outputs[2340] = ~((layer0_outputs[3119]) ^ (layer0_outputs[4887]));
    assign layer1_outputs[2341] = layer0_outputs[1193];
    assign layer1_outputs[2342] = 1'b0;
    assign layer1_outputs[2343] = ~((layer0_outputs[3996]) & (layer0_outputs[2294]));
    assign layer1_outputs[2344] = ~((layer0_outputs[5112]) | (layer0_outputs[695]));
    assign layer1_outputs[2345] = 1'b1;
    assign layer1_outputs[2346] = layer0_outputs[1721];
    assign layer1_outputs[2347] = ~((layer0_outputs[729]) ^ (layer0_outputs[893]));
    assign layer1_outputs[2348] = (layer0_outputs[4250]) | (layer0_outputs[1278]);
    assign layer1_outputs[2349] = ~(layer0_outputs[2950]) | (layer0_outputs[4024]);
    assign layer1_outputs[2350] = (layer0_outputs[1534]) ^ (layer0_outputs[3939]);
    assign layer1_outputs[2351] = (layer0_outputs[1167]) & (layer0_outputs[1573]);
    assign layer1_outputs[2352] = ~(layer0_outputs[3409]);
    assign layer1_outputs[2353] = (layer0_outputs[1603]) | (layer0_outputs[758]);
    assign layer1_outputs[2354] = (layer0_outputs[3657]) & ~(layer0_outputs[1920]);
    assign layer1_outputs[2355] = (layer0_outputs[5027]) & ~(layer0_outputs[820]);
    assign layer1_outputs[2356] = layer0_outputs[2450];
    assign layer1_outputs[2357] = ~((layer0_outputs[1167]) | (layer0_outputs[5026]));
    assign layer1_outputs[2358] = (layer0_outputs[31]) & ~(layer0_outputs[2424]);
    assign layer1_outputs[2359] = (layer0_outputs[1292]) & (layer0_outputs[3117]);
    assign layer1_outputs[2360] = ~((layer0_outputs[3125]) & (layer0_outputs[4692]));
    assign layer1_outputs[2361] = ~(layer0_outputs[3627]);
    assign layer1_outputs[2362] = ~((layer0_outputs[4224]) & (layer0_outputs[1299]));
    assign layer1_outputs[2363] = (layer0_outputs[5055]) & (layer0_outputs[310]);
    assign layer1_outputs[2364] = layer0_outputs[27];
    assign layer1_outputs[2365] = 1'b0;
    assign layer1_outputs[2366] = ~((layer0_outputs[720]) & (layer0_outputs[4110]));
    assign layer1_outputs[2367] = ~(layer0_outputs[3429]) | (layer0_outputs[3006]);
    assign layer1_outputs[2368] = ~(layer0_outputs[4348]) | (layer0_outputs[216]);
    assign layer1_outputs[2369] = layer0_outputs[2635];
    assign layer1_outputs[2370] = 1'b0;
    assign layer1_outputs[2371] = (layer0_outputs[4838]) & ~(layer0_outputs[3074]);
    assign layer1_outputs[2372] = ~(layer0_outputs[3716]);
    assign layer1_outputs[2373] = 1'b1;
    assign layer1_outputs[2374] = ~(layer0_outputs[3360]) | (layer0_outputs[94]);
    assign layer1_outputs[2375] = (layer0_outputs[4448]) & ~(layer0_outputs[1889]);
    assign layer1_outputs[2376] = ~(layer0_outputs[5025]);
    assign layer1_outputs[2377] = (layer0_outputs[3696]) & ~(layer0_outputs[5074]);
    assign layer1_outputs[2378] = ~((layer0_outputs[865]) & (layer0_outputs[3684]));
    assign layer1_outputs[2379] = ~(layer0_outputs[316]);
    assign layer1_outputs[2380] = (layer0_outputs[3766]) | (layer0_outputs[475]);
    assign layer1_outputs[2381] = ~((layer0_outputs[2088]) & (layer0_outputs[583]));
    assign layer1_outputs[2382] = ~(layer0_outputs[692]);
    assign layer1_outputs[2383] = ~(layer0_outputs[2011]) | (layer0_outputs[3269]);
    assign layer1_outputs[2384] = (layer0_outputs[2736]) & ~(layer0_outputs[3708]);
    assign layer1_outputs[2385] = layer0_outputs[4298];
    assign layer1_outputs[2386] = (layer0_outputs[4441]) | (layer0_outputs[2621]);
    assign layer1_outputs[2387] = ~((layer0_outputs[2015]) | (layer0_outputs[1071]));
    assign layer1_outputs[2388] = ~(layer0_outputs[2342]);
    assign layer1_outputs[2389] = (layer0_outputs[2156]) & ~(layer0_outputs[250]);
    assign layer1_outputs[2390] = layer0_outputs[264];
    assign layer1_outputs[2391] = 1'b0;
    assign layer1_outputs[2392] = 1'b0;
    assign layer1_outputs[2393] = ~(layer0_outputs[4745]);
    assign layer1_outputs[2394] = ~((layer0_outputs[1826]) & (layer0_outputs[887]));
    assign layer1_outputs[2395] = ~(layer0_outputs[2744]) | (layer0_outputs[1797]);
    assign layer1_outputs[2396] = layer0_outputs[3576];
    assign layer1_outputs[2397] = ~((layer0_outputs[500]) | (layer0_outputs[4578]));
    assign layer1_outputs[2398] = ~(layer0_outputs[1568]);
    assign layer1_outputs[2399] = ~(layer0_outputs[5050]);
    assign layer1_outputs[2400] = 1'b0;
    assign layer1_outputs[2401] = (layer0_outputs[740]) & ~(layer0_outputs[3504]);
    assign layer1_outputs[2402] = ~(layer0_outputs[3888]) | (layer0_outputs[3885]);
    assign layer1_outputs[2403] = (layer0_outputs[2485]) & (layer0_outputs[3579]);
    assign layer1_outputs[2404] = ~((layer0_outputs[850]) & (layer0_outputs[2515]));
    assign layer1_outputs[2405] = ~(layer0_outputs[2333]);
    assign layer1_outputs[2406] = ~(layer0_outputs[2540]);
    assign layer1_outputs[2407] = (layer0_outputs[2524]) & ~(layer0_outputs[1793]);
    assign layer1_outputs[2408] = layer0_outputs[1250];
    assign layer1_outputs[2409] = ~((layer0_outputs[1371]) | (layer0_outputs[1570]));
    assign layer1_outputs[2410] = (layer0_outputs[3711]) & (layer0_outputs[4370]);
    assign layer1_outputs[2411] = (layer0_outputs[242]) ^ (layer0_outputs[4612]);
    assign layer1_outputs[2412] = layer0_outputs[609];
    assign layer1_outputs[2413] = (layer0_outputs[689]) & ~(layer0_outputs[1390]);
    assign layer1_outputs[2414] = 1'b0;
    assign layer1_outputs[2415] = 1'b1;
    assign layer1_outputs[2416] = ~(layer0_outputs[671]);
    assign layer1_outputs[2417] = layer0_outputs[834];
    assign layer1_outputs[2418] = layer0_outputs[4448];
    assign layer1_outputs[2419] = ~(layer0_outputs[4618]);
    assign layer1_outputs[2420] = ~(layer0_outputs[4184]) | (layer0_outputs[278]);
    assign layer1_outputs[2421] = ~(layer0_outputs[3293]) | (layer0_outputs[3299]);
    assign layer1_outputs[2422] = layer0_outputs[721];
    assign layer1_outputs[2423] = 1'b1;
    assign layer1_outputs[2424] = (layer0_outputs[2534]) & ~(layer0_outputs[4661]);
    assign layer1_outputs[2425] = ~((layer0_outputs[2573]) & (layer0_outputs[4888]));
    assign layer1_outputs[2426] = ~(layer0_outputs[4812]) | (layer0_outputs[2864]);
    assign layer1_outputs[2427] = ~((layer0_outputs[1636]) ^ (layer0_outputs[1891]));
    assign layer1_outputs[2428] = 1'b0;
    assign layer1_outputs[2429] = (layer0_outputs[3446]) & (layer0_outputs[2996]);
    assign layer1_outputs[2430] = ~((layer0_outputs[2845]) ^ (layer0_outputs[5001]));
    assign layer1_outputs[2431] = ~((layer0_outputs[3542]) | (layer0_outputs[4646]));
    assign layer1_outputs[2432] = layer0_outputs[3644];
    assign layer1_outputs[2433] = ~((layer0_outputs[2951]) ^ (layer0_outputs[2824]));
    assign layer1_outputs[2434] = (layer0_outputs[4223]) & (layer0_outputs[106]);
    assign layer1_outputs[2435] = 1'b0;
    assign layer1_outputs[2436] = layer0_outputs[4075];
    assign layer1_outputs[2437] = 1'b1;
    assign layer1_outputs[2438] = ~(layer0_outputs[3732]);
    assign layer1_outputs[2439] = (layer0_outputs[1849]) & ~(layer0_outputs[2051]);
    assign layer1_outputs[2440] = ~((layer0_outputs[4792]) | (layer0_outputs[4678]));
    assign layer1_outputs[2441] = layer0_outputs[3455];
    assign layer1_outputs[2442] = 1'b1;
    assign layer1_outputs[2443] = ~((layer0_outputs[4547]) | (layer0_outputs[4522]));
    assign layer1_outputs[2444] = ~((layer0_outputs[1688]) & (layer0_outputs[2004]));
    assign layer1_outputs[2445] = 1'b1;
    assign layer1_outputs[2446] = (layer0_outputs[1776]) & ~(layer0_outputs[3759]);
    assign layer1_outputs[2447] = (layer0_outputs[4839]) & (layer0_outputs[4977]);
    assign layer1_outputs[2448] = layer0_outputs[517];
    assign layer1_outputs[2449] = (layer0_outputs[1112]) | (layer0_outputs[1931]);
    assign layer1_outputs[2450] = 1'b0;
    assign layer1_outputs[2451] = layer0_outputs[2319];
    assign layer1_outputs[2452] = 1'b0;
    assign layer1_outputs[2453] = ~(layer0_outputs[4]) | (layer0_outputs[3103]);
    assign layer1_outputs[2454] = ~((layer0_outputs[2527]) | (layer0_outputs[2104]));
    assign layer1_outputs[2455] = ~(layer0_outputs[3063]);
    assign layer1_outputs[2456] = ~(layer0_outputs[3926]);
    assign layer1_outputs[2457] = ~((layer0_outputs[4701]) & (layer0_outputs[3009]));
    assign layer1_outputs[2458] = ~(layer0_outputs[1064]);
    assign layer1_outputs[2459] = ~((layer0_outputs[1341]) | (layer0_outputs[5002]));
    assign layer1_outputs[2460] = 1'b1;
    assign layer1_outputs[2461] = 1'b1;
    assign layer1_outputs[2462] = ~(layer0_outputs[991]);
    assign layer1_outputs[2463] = (layer0_outputs[4262]) | (layer0_outputs[2221]);
    assign layer1_outputs[2464] = ~((layer0_outputs[708]) | (layer0_outputs[566]));
    assign layer1_outputs[2465] = ~(layer0_outputs[1622]) | (layer0_outputs[216]);
    assign layer1_outputs[2466] = ~(layer0_outputs[4465]);
    assign layer1_outputs[2467] = ~(layer0_outputs[3419]);
    assign layer1_outputs[2468] = (layer0_outputs[487]) & ~(layer0_outputs[5118]);
    assign layer1_outputs[2469] = (layer0_outputs[838]) | (layer0_outputs[4844]);
    assign layer1_outputs[2470] = layer0_outputs[211];
    assign layer1_outputs[2471] = (layer0_outputs[1371]) & ~(layer0_outputs[2542]);
    assign layer1_outputs[2472] = layer0_outputs[3116];
    assign layer1_outputs[2473] = (layer0_outputs[293]) | (layer0_outputs[2670]);
    assign layer1_outputs[2474] = layer0_outputs[164];
    assign layer1_outputs[2475] = ~(layer0_outputs[4624]);
    assign layer1_outputs[2476] = ~((layer0_outputs[2765]) | (layer0_outputs[3650]));
    assign layer1_outputs[2477] = (layer0_outputs[1149]) & ~(layer0_outputs[1943]);
    assign layer1_outputs[2478] = ~(layer0_outputs[2808]);
    assign layer1_outputs[2479] = ~(layer0_outputs[1840]) | (layer0_outputs[558]);
    assign layer1_outputs[2480] = ~((layer0_outputs[1791]) | (layer0_outputs[638]));
    assign layer1_outputs[2481] = (layer0_outputs[418]) & ~(layer0_outputs[1226]);
    assign layer1_outputs[2482] = ~((layer0_outputs[2124]) & (layer0_outputs[1739]));
    assign layer1_outputs[2483] = 1'b1;
    assign layer1_outputs[2484] = ~(layer0_outputs[1820]) | (layer0_outputs[2095]);
    assign layer1_outputs[2485] = (layer0_outputs[456]) & ~(layer0_outputs[1766]);
    assign layer1_outputs[2486] = (layer0_outputs[679]) & (layer0_outputs[3019]);
    assign layer1_outputs[2487] = ~(layer0_outputs[4672]) | (layer0_outputs[3217]);
    assign layer1_outputs[2488] = ~((layer0_outputs[809]) & (layer0_outputs[2705]));
    assign layer1_outputs[2489] = ~(layer0_outputs[208]) | (layer0_outputs[3204]);
    assign layer1_outputs[2490] = ~(layer0_outputs[767]);
    assign layer1_outputs[2491] = ~(layer0_outputs[51]);
    assign layer1_outputs[2492] = ~(layer0_outputs[684]);
    assign layer1_outputs[2493] = ~((layer0_outputs[1736]) | (layer0_outputs[1407]));
    assign layer1_outputs[2494] = layer0_outputs[2800];
    assign layer1_outputs[2495] = (layer0_outputs[3802]) & ~(layer0_outputs[2168]);
    assign layer1_outputs[2496] = ~((layer0_outputs[107]) | (layer0_outputs[3975]));
    assign layer1_outputs[2497] = ~(layer0_outputs[858]);
    assign layer1_outputs[2498] = ~(layer0_outputs[855]);
    assign layer1_outputs[2499] = 1'b1;
    assign layer1_outputs[2500] = (layer0_outputs[449]) & ~(layer0_outputs[2123]);
    assign layer1_outputs[2501] = ~(layer0_outputs[2234]) | (layer0_outputs[3960]);
    assign layer1_outputs[2502] = 1'b1;
    assign layer1_outputs[2503] = 1'b1;
    assign layer1_outputs[2504] = 1'b0;
    assign layer1_outputs[2505] = 1'b1;
    assign layer1_outputs[2506] = (layer0_outputs[1073]) | (layer0_outputs[4271]);
    assign layer1_outputs[2507] = ~(layer0_outputs[4056]);
    assign layer1_outputs[2508] = 1'b1;
    assign layer1_outputs[2509] = ~(layer0_outputs[4260]) | (layer0_outputs[998]);
    assign layer1_outputs[2510] = (layer0_outputs[4869]) & (layer0_outputs[2052]);
    assign layer1_outputs[2511] = ~(layer0_outputs[3562]);
    assign layer1_outputs[2512] = 1'b0;
    assign layer1_outputs[2513] = ~((layer0_outputs[976]) & (layer0_outputs[1749]));
    assign layer1_outputs[2514] = ~((layer0_outputs[3972]) | (layer0_outputs[2837]));
    assign layer1_outputs[2515] = (layer0_outputs[2323]) & ~(layer0_outputs[83]);
    assign layer1_outputs[2516] = (layer0_outputs[2075]) | (layer0_outputs[1827]);
    assign layer1_outputs[2517] = 1'b0;
    assign layer1_outputs[2518] = ~((layer0_outputs[2193]) | (layer0_outputs[4893]));
    assign layer1_outputs[2519] = ~((layer0_outputs[3049]) | (layer0_outputs[1846]));
    assign layer1_outputs[2520] = layer0_outputs[178];
    assign layer1_outputs[2521] = 1'b0;
    assign layer1_outputs[2522] = ~(layer0_outputs[4704]);
    assign layer1_outputs[2523] = layer0_outputs[5042];
    assign layer1_outputs[2524] = ~((layer0_outputs[4326]) | (layer0_outputs[227]));
    assign layer1_outputs[2525] = ~(layer0_outputs[1317]);
    assign layer1_outputs[2526] = 1'b0;
    assign layer1_outputs[2527] = ~(layer0_outputs[2362]);
    assign layer1_outputs[2528] = (layer0_outputs[2586]) & ~(layer0_outputs[578]);
    assign layer1_outputs[2529] = ~(layer0_outputs[622]);
    assign layer1_outputs[2530] = ~((layer0_outputs[1259]) ^ (layer0_outputs[1896]));
    assign layer1_outputs[2531] = 1'b0;
    assign layer1_outputs[2532] = (layer0_outputs[3135]) & (layer0_outputs[606]);
    assign layer1_outputs[2533] = (layer0_outputs[4933]) ^ (layer0_outputs[1838]);
    assign layer1_outputs[2534] = 1'b1;
    assign layer1_outputs[2535] = ~(layer0_outputs[209]);
    assign layer1_outputs[2536] = 1'b1;
    assign layer1_outputs[2537] = (layer0_outputs[3932]) & (layer0_outputs[3697]);
    assign layer1_outputs[2538] = (layer0_outputs[3214]) & ~(layer0_outputs[2606]);
    assign layer1_outputs[2539] = (layer0_outputs[1003]) & (layer0_outputs[803]);
    assign layer1_outputs[2540] = (layer0_outputs[4310]) & ~(layer0_outputs[2324]);
    assign layer1_outputs[2541] = (layer0_outputs[2860]) & ~(layer0_outputs[1815]);
    assign layer1_outputs[2542] = ~(layer0_outputs[3927]) | (layer0_outputs[2581]);
    assign layer1_outputs[2543] = 1'b1;
    assign layer1_outputs[2544] = (layer0_outputs[1667]) | (layer0_outputs[1118]);
    assign layer1_outputs[2545] = (layer0_outputs[530]) & (layer0_outputs[5047]);
    assign layer1_outputs[2546] = 1'b0;
    assign layer1_outputs[2547] = ~((layer0_outputs[2549]) | (layer0_outputs[1831]));
    assign layer1_outputs[2548] = ~(layer0_outputs[1590]);
    assign layer1_outputs[2549] = ~((layer0_outputs[2795]) | (layer0_outputs[2365]));
    assign layer1_outputs[2550] = 1'b0;
    assign layer1_outputs[2551] = ~(layer0_outputs[3115]) | (layer0_outputs[3556]);
    assign layer1_outputs[2552] = (layer0_outputs[1378]) & (layer0_outputs[2073]);
    assign layer1_outputs[2553] = layer0_outputs[512];
    assign layer1_outputs[2554] = (layer0_outputs[736]) & ~(layer0_outputs[811]);
    assign layer1_outputs[2555] = (layer0_outputs[2971]) & ~(layer0_outputs[1765]);
    assign layer1_outputs[2556] = 1'b0;
    assign layer1_outputs[2557] = (layer0_outputs[2259]) & (layer0_outputs[4117]);
    assign layer1_outputs[2558] = layer0_outputs[4576];
    assign layer1_outputs[2559] = (layer0_outputs[264]) & ~(layer0_outputs[3602]);
    assign layer1_outputs[2560] = (layer0_outputs[1215]) ^ (layer0_outputs[4288]);
    assign layer1_outputs[2561] = ~(layer0_outputs[1313]);
    assign layer1_outputs[2562] = (layer0_outputs[267]) | (layer0_outputs[4240]);
    assign layer1_outputs[2563] = ~((layer0_outputs[1919]) | (layer0_outputs[3358]));
    assign layer1_outputs[2564] = ~(layer0_outputs[752]);
    assign layer1_outputs[2565] = ~(layer0_outputs[783]);
    assign layer1_outputs[2566] = ~(layer0_outputs[1805]) | (layer0_outputs[4013]);
    assign layer1_outputs[2567] = ~(layer0_outputs[2132]);
    assign layer1_outputs[2568] = ~((layer0_outputs[1578]) & (layer0_outputs[3822]));
    assign layer1_outputs[2569] = (layer0_outputs[536]) & (layer0_outputs[2600]);
    assign layer1_outputs[2570] = ~(layer0_outputs[3641]) | (layer0_outputs[3728]);
    assign layer1_outputs[2571] = ~((layer0_outputs[4941]) | (layer0_outputs[1387]));
    assign layer1_outputs[2572] = layer0_outputs[1514];
    assign layer1_outputs[2573] = ~(layer0_outputs[3925]);
    assign layer1_outputs[2574] = (layer0_outputs[2639]) & (layer0_outputs[1210]);
    assign layer1_outputs[2575] = ~((layer0_outputs[5056]) | (layer0_outputs[4487]));
    assign layer1_outputs[2576] = layer0_outputs[2159];
    assign layer1_outputs[2577] = ~(layer0_outputs[3264]);
    assign layer1_outputs[2578] = ~((layer0_outputs[3486]) | (layer0_outputs[4338]));
    assign layer1_outputs[2579] = (layer0_outputs[2145]) & ~(layer0_outputs[2404]);
    assign layer1_outputs[2580] = (layer0_outputs[3864]) & ~(layer0_outputs[4209]);
    assign layer1_outputs[2581] = ~(layer0_outputs[2531]);
    assign layer1_outputs[2582] = (layer0_outputs[2765]) & ~(layer0_outputs[223]);
    assign layer1_outputs[2583] = ~(layer0_outputs[1532]) | (layer0_outputs[3803]);
    assign layer1_outputs[2584] = (layer0_outputs[3050]) | (layer0_outputs[2795]);
    assign layer1_outputs[2585] = ~((layer0_outputs[4127]) & (layer0_outputs[3217]));
    assign layer1_outputs[2586] = (layer0_outputs[2170]) & ~(layer0_outputs[1674]);
    assign layer1_outputs[2587] = ~(layer0_outputs[3681]);
    assign layer1_outputs[2588] = (layer0_outputs[2199]) & ~(layer0_outputs[5031]);
    assign layer1_outputs[2589] = 1'b1;
    assign layer1_outputs[2590] = (layer0_outputs[3045]) & (layer0_outputs[4263]);
    assign layer1_outputs[2591] = (layer0_outputs[2722]) ^ (layer0_outputs[1787]);
    assign layer1_outputs[2592] = ~(layer0_outputs[17]) | (layer0_outputs[2739]);
    assign layer1_outputs[2593] = layer0_outputs[4566];
    assign layer1_outputs[2594] = 1'b1;
    assign layer1_outputs[2595] = layer0_outputs[3314];
    assign layer1_outputs[2596] = (layer0_outputs[2131]) & ~(layer0_outputs[2716]);
    assign layer1_outputs[2597] = ~(layer0_outputs[906]);
    assign layer1_outputs[2598] = ~(layer0_outputs[3848]);
    assign layer1_outputs[2599] = ~((layer0_outputs[4201]) & (layer0_outputs[2858]));
    assign layer1_outputs[2600] = (layer0_outputs[3146]) & (layer0_outputs[336]);
    assign layer1_outputs[2601] = (layer0_outputs[2970]) & (layer0_outputs[929]);
    assign layer1_outputs[2602] = layer0_outputs[3137];
    assign layer1_outputs[2603] = (layer0_outputs[2946]) ^ (layer0_outputs[2196]);
    assign layer1_outputs[2604] = ~(layer0_outputs[3198]);
    assign layer1_outputs[2605] = ~((layer0_outputs[1611]) | (layer0_outputs[3142]));
    assign layer1_outputs[2606] = (layer0_outputs[2104]) & (layer0_outputs[2275]);
    assign layer1_outputs[2607] = 1'b1;
    assign layer1_outputs[2608] = 1'b0;
    assign layer1_outputs[2609] = layer0_outputs[4237];
    assign layer1_outputs[2610] = layer0_outputs[66];
    assign layer1_outputs[2611] = 1'b1;
    assign layer1_outputs[2612] = ~(layer0_outputs[2041]) | (layer0_outputs[1083]);
    assign layer1_outputs[2613] = layer0_outputs[3526];
    assign layer1_outputs[2614] = (layer0_outputs[3438]) & ~(layer0_outputs[4452]);
    assign layer1_outputs[2615] = (layer0_outputs[1537]) & ~(layer0_outputs[2412]);
    assign layer1_outputs[2616] = (layer0_outputs[4188]) & ~(layer0_outputs[5011]);
    assign layer1_outputs[2617] = layer0_outputs[319];
    assign layer1_outputs[2618] = ~(layer0_outputs[4997]) | (layer0_outputs[4294]);
    assign layer1_outputs[2619] = ~(layer0_outputs[3118]);
    assign layer1_outputs[2620] = ~((layer0_outputs[706]) & (layer0_outputs[3313]));
    assign layer1_outputs[2621] = (layer0_outputs[5000]) | (layer0_outputs[1592]);
    assign layer1_outputs[2622] = ~(layer0_outputs[3666]);
    assign layer1_outputs[2623] = 1'b0;
    assign layer1_outputs[2624] = ~((layer0_outputs[4715]) & (layer0_outputs[4040]));
    assign layer1_outputs[2625] = (layer0_outputs[2563]) ^ (layer0_outputs[4585]);
    assign layer1_outputs[2626] = (layer0_outputs[917]) & ~(layer0_outputs[1543]);
    assign layer1_outputs[2627] = ~(layer0_outputs[3942]) | (layer0_outputs[3312]);
    assign layer1_outputs[2628] = 1'b1;
    assign layer1_outputs[2629] = ~(layer0_outputs[2755]) | (layer0_outputs[1423]);
    assign layer1_outputs[2630] = ~(layer0_outputs[452]);
    assign layer1_outputs[2631] = ~(layer0_outputs[1456]) | (layer0_outputs[1384]);
    assign layer1_outputs[2632] = 1'b0;
    assign layer1_outputs[2633] = (layer0_outputs[1339]) & (layer0_outputs[4010]);
    assign layer1_outputs[2634] = layer0_outputs[4895];
    assign layer1_outputs[2635] = ~(layer0_outputs[897]);
    assign layer1_outputs[2636] = 1'b1;
    assign layer1_outputs[2637] = layer0_outputs[1409];
    assign layer1_outputs[2638] = (layer0_outputs[2677]) | (layer0_outputs[3507]);
    assign layer1_outputs[2639] = 1'b1;
    assign layer1_outputs[2640] = (layer0_outputs[2059]) & (layer0_outputs[3557]);
    assign layer1_outputs[2641] = layer0_outputs[4386];
    assign layer1_outputs[2642] = 1'b1;
    assign layer1_outputs[2643] = ~((layer0_outputs[3451]) & (layer0_outputs[948]));
    assign layer1_outputs[2644] = 1'b0;
    assign layer1_outputs[2645] = (layer0_outputs[2554]) ^ (layer0_outputs[2543]);
    assign layer1_outputs[2646] = layer0_outputs[2920];
    assign layer1_outputs[2647] = ~((layer0_outputs[1416]) & (layer0_outputs[3182]));
    assign layer1_outputs[2648] = 1'b1;
    assign layer1_outputs[2649] = (layer0_outputs[2497]) | (layer0_outputs[2890]);
    assign layer1_outputs[2650] = (layer0_outputs[357]) & ~(layer0_outputs[3879]);
    assign layer1_outputs[2651] = (layer0_outputs[975]) | (layer0_outputs[792]);
    assign layer1_outputs[2652] = (layer0_outputs[3519]) & (layer0_outputs[4292]);
    assign layer1_outputs[2653] = (layer0_outputs[2687]) & ~(layer0_outputs[3980]);
    assign layer1_outputs[2654] = 1'b1;
    assign layer1_outputs[2655] = ~((layer0_outputs[524]) & (layer0_outputs[3540]));
    assign layer1_outputs[2656] = (layer0_outputs[1812]) & ~(layer0_outputs[1706]);
    assign layer1_outputs[2657] = ~(layer0_outputs[4339]) | (layer0_outputs[5027]);
    assign layer1_outputs[2658] = ~(layer0_outputs[2897]);
    assign layer1_outputs[2659] = ~(layer0_outputs[513]);
    assign layer1_outputs[2660] = (layer0_outputs[1284]) & ~(layer0_outputs[2213]);
    assign layer1_outputs[2661] = (layer0_outputs[3290]) ^ (layer0_outputs[617]);
    assign layer1_outputs[2662] = ~((layer0_outputs[1348]) & (layer0_outputs[4322]));
    assign layer1_outputs[2663] = ~((layer0_outputs[1129]) & (layer0_outputs[4404]));
    assign layer1_outputs[2664] = ~(layer0_outputs[4021]) | (layer0_outputs[4312]);
    assign layer1_outputs[2665] = ~(layer0_outputs[822]) | (layer0_outputs[2790]);
    assign layer1_outputs[2666] = 1'b0;
    assign layer1_outputs[2667] = 1'b1;
    assign layer1_outputs[2668] = ~(layer0_outputs[3169]) | (layer0_outputs[3516]);
    assign layer1_outputs[2669] = ~(layer0_outputs[1598]) | (layer0_outputs[137]);
    assign layer1_outputs[2670] = layer0_outputs[3731];
    assign layer1_outputs[2671] = ~((layer0_outputs[4279]) ^ (layer0_outputs[2619]));
    assign layer1_outputs[2672] = ~((layer0_outputs[2]) & (layer0_outputs[614]));
    assign layer1_outputs[2673] = ~((layer0_outputs[2160]) | (layer0_outputs[4204]));
    assign layer1_outputs[2674] = (layer0_outputs[4447]) & (layer0_outputs[3783]);
    assign layer1_outputs[2675] = layer0_outputs[846];
    assign layer1_outputs[2676] = ~((layer0_outputs[112]) | (layer0_outputs[4690]));
    assign layer1_outputs[2677] = ~(layer0_outputs[4150]) | (layer0_outputs[2722]);
    assign layer1_outputs[2678] = layer0_outputs[3000];
    assign layer1_outputs[2679] = ~(layer0_outputs[4105]) | (layer0_outputs[4766]);
    assign layer1_outputs[2680] = ~(layer0_outputs[3190]) | (layer0_outputs[765]);
    assign layer1_outputs[2681] = (layer0_outputs[3169]) | (layer0_outputs[1110]);
    assign layer1_outputs[2682] = 1'b1;
    assign layer1_outputs[2683] = (layer0_outputs[587]) & (layer0_outputs[5066]);
    assign layer1_outputs[2684] = ~(layer0_outputs[2337]);
    assign layer1_outputs[2685] = ~(layer0_outputs[461]) | (layer0_outputs[4316]);
    assign layer1_outputs[2686] = (layer0_outputs[3447]) | (layer0_outputs[4830]);
    assign layer1_outputs[2687] = ~(layer0_outputs[4516]);
    assign layer1_outputs[2688] = ~((layer0_outputs[2325]) | (layer0_outputs[1256]));
    assign layer1_outputs[2689] = (layer0_outputs[2727]) & (layer0_outputs[2135]);
    assign layer1_outputs[2690] = ~((layer0_outputs[716]) | (layer0_outputs[3246]));
    assign layer1_outputs[2691] = ~((layer0_outputs[3027]) & (layer0_outputs[2420]));
    assign layer1_outputs[2692] = 1'b1;
    assign layer1_outputs[2693] = ~(layer0_outputs[1323]);
    assign layer1_outputs[2694] = (layer0_outputs[4456]) & (layer0_outputs[3254]);
    assign layer1_outputs[2695] = 1'b1;
    assign layer1_outputs[2696] = ~(layer0_outputs[3151]) | (layer0_outputs[1902]);
    assign layer1_outputs[2697] = (layer0_outputs[1550]) & ~(layer0_outputs[2270]);
    assign layer1_outputs[2698] = ~(layer0_outputs[2163]) | (layer0_outputs[4427]);
    assign layer1_outputs[2699] = ~(layer0_outputs[3001]);
    assign layer1_outputs[2700] = (layer0_outputs[1400]) & (layer0_outputs[4767]);
    assign layer1_outputs[2701] = ~((layer0_outputs[3913]) | (layer0_outputs[2604]));
    assign layer1_outputs[2702] = layer0_outputs[399];
    assign layer1_outputs[2703] = (layer0_outputs[3075]) & ~(layer0_outputs[1109]);
    assign layer1_outputs[2704] = layer0_outputs[3585];
    assign layer1_outputs[2705] = (layer0_outputs[3121]) | (layer0_outputs[151]);
    assign layer1_outputs[2706] = layer0_outputs[3198];
    assign layer1_outputs[2707] = ~(layer0_outputs[4041]);
    assign layer1_outputs[2708] = ~(layer0_outputs[3571]);
    assign layer1_outputs[2709] = (layer0_outputs[1133]) ^ (layer0_outputs[1772]);
    assign layer1_outputs[2710] = layer0_outputs[3044];
    assign layer1_outputs[2711] = layer0_outputs[1614];
    assign layer1_outputs[2712] = layer0_outputs[2384];
    assign layer1_outputs[2713] = 1'b0;
    assign layer1_outputs[2714] = ~(layer0_outputs[1184]);
    assign layer1_outputs[2715] = (layer0_outputs[4686]) ^ (layer0_outputs[2198]);
    assign layer1_outputs[2716] = layer0_outputs[754];
    assign layer1_outputs[2717] = ~(layer0_outputs[304]);
    assign layer1_outputs[2718] = ~((layer0_outputs[1865]) ^ (layer0_outputs[2186]));
    assign layer1_outputs[2719] = (layer0_outputs[4646]) & ~(layer0_outputs[2313]);
    assign layer1_outputs[2720] = (layer0_outputs[3912]) & (layer0_outputs[1157]);
    assign layer1_outputs[2721] = 1'b0;
    assign layer1_outputs[2722] = 1'b0;
    assign layer1_outputs[2723] = 1'b0;
    assign layer1_outputs[2724] = 1'b1;
    assign layer1_outputs[2725] = ~((layer0_outputs[2191]) | (layer0_outputs[51]));
    assign layer1_outputs[2726] = (layer0_outputs[4749]) | (layer0_outputs[2476]);
    assign layer1_outputs[2727] = 1'b1;
    assign layer1_outputs[2728] = (layer0_outputs[3076]) & (layer0_outputs[3064]);
    assign layer1_outputs[2729] = ~((layer0_outputs[1679]) | (layer0_outputs[2719]));
    assign layer1_outputs[2730] = (layer0_outputs[4102]) & (layer0_outputs[5037]);
    assign layer1_outputs[2731] = ~(layer0_outputs[4341]) | (layer0_outputs[522]);
    assign layer1_outputs[2732] = ~((layer0_outputs[4307]) & (layer0_outputs[4947]));
    assign layer1_outputs[2733] = (layer0_outputs[2367]) ^ (layer0_outputs[3007]);
    assign layer1_outputs[2734] = ~((layer0_outputs[3502]) | (layer0_outputs[287]));
    assign layer1_outputs[2735] = layer0_outputs[580];
    assign layer1_outputs[2736] = 1'b1;
    assign layer1_outputs[2737] = 1'b1;
    assign layer1_outputs[2738] = ~((layer0_outputs[1231]) | (layer0_outputs[4435]));
    assign layer1_outputs[2739] = ~((layer0_outputs[80]) | (layer0_outputs[4570]));
    assign layer1_outputs[2740] = (layer0_outputs[4550]) & (layer0_outputs[1513]);
    assign layer1_outputs[2741] = (layer0_outputs[2115]) & (layer0_outputs[4480]);
    assign layer1_outputs[2742] = ~(layer0_outputs[237]) | (layer0_outputs[870]);
    assign layer1_outputs[2743] = (layer0_outputs[2361]) & (layer0_outputs[2501]);
    assign layer1_outputs[2744] = (layer0_outputs[2828]) & ~(layer0_outputs[4593]);
    assign layer1_outputs[2745] = layer0_outputs[1322];
    assign layer1_outputs[2746] = (layer0_outputs[1563]) & ~(layer0_outputs[768]);
    assign layer1_outputs[2747] = (layer0_outputs[607]) & ~(layer0_outputs[1292]);
    assign layer1_outputs[2748] = (layer0_outputs[4319]) | (layer0_outputs[32]);
    assign layer1_outputs[2749] = (layer0_outputs[2763]) ^ (layer0_outputs[2292]);
    assign layer1_outputs[2750] = (layer0_outputs[3245]) | (layer0_outputs[70]);
    assign layer1_outputs[2751] = ~(layer0_outputs[1050]) | (layer0_outputs[2999]);
    assign layer1_outputs[2752] = (layer0_outputs[594]) & (layer0_outputs[4140]);
    assign layer1_outputs[2753] = (layer0_outputs[2121]) & ~(layer0_outputs[173]);
    assign layer1_outputs[2754] = (layer0_outputs[3405]) & (layer0_outputs[2036]);
    assign layer1_outputs[2755] = (layer0_outputs[326]) & ~(layer0_outputs[2671]);
    assign layer1_outputs[2756] = (layer0_outputs[348]) | (layer0_outputs[3361]);
    assign layer1_outputs[2757] = ~(layer0_outputs[2343]);
    assign layer1_outputs[2758] = 1'b0;
    assign layer1_outputs[2759] = ~((layer0_outputs[448]) & (layer0_outputs[94]));
    assign layer1_outputs[2760] = 1'b1;
    assign layer1_outputs[2761] = ~((layer0_outputs[3926]) & (layer0_outputs[8]));
    assign layer1_outputs[2762] = 1'b1;
    assign layer1_outputs[2763] = 1'b0;
    assign layer1_outputs[2764] = ~((layer0_outputs[516]) | (layer0_outputs[4078]));
    assign layer1_outputs[2765] = (layer0_outputs[2487]) | (layer0_outputs[2641]);
    assign layer1_outputs[2766] = ~((layer0_outputs[1057]) & (layer0_outputs[1188]));
    assign layer1_outputs[2767] = ~(layer0_outputs[3983]);
    assign layer1_outputs[2768] = ~(layer0_outputs[2990]) | (layer0_outputs[2822]);
    assign layer1_outputs[2769] = ~(layer0_outputs[2178]) | (layer0_outputs[451]);
    assign layer1_outputs[2770] = layer0_outputs[933];
    assign layer1_outputs[2771] = ~(layer0_outputs[4328]);
    assign layer1_outputs[2772] = (layer0_outputs[16]) & ~(layer0_outputs[4291]);
    assign layer1_outputs[2773] = ~(layer0_outputs[65]) | (layer0_outputs[4718]);
    assign layer1_outputs[2774] = layer0_outputs[1880];
    assign layer1_outputs[2775] = (layer0_outputs[118]) | (layer0_outputs[1593]);
    assign layer1_outputs[2776] = (layer0_outputs[2464]) | (layer0_outputs[2373]);
    assign layer1_outputs[2777] = (layer0_outputs[3185]) | (layer0_outputs[4320]);
    assign layer1_outputs[2778] = (layer0_outputs[128]) | (layer0_outputs[1672]);
    assign layer1_outputs[2779] = layer0_outputs[395];
    assign layer1_outputs[2780] = 1'b0;
    assign layer1_outputs[2781] = 1'b1;
    assign layer1_outputs[2782] = layer0_outputs[1770];
    assign layer1_outputs[2783] = ~(layer0_outputs[2643]) | (layer0_outputs[1630]);
    assign layer1_outputs[2784] = ~(layer0_outputs[975]);
    assign layer1_outputs[2785] = layer0_outputs[3546];
    assign layer1_outputs[2786] = (layer0_outputs[1380]) & (layer0_outputs[1414]);
    assign layer1_outputs[2787] = ~((layer0_outputs[4860]) & (layer0_outputs[1707]));
    assign layer1_outputs[2788] = layer0_outputs[1410];
    assign layer1_outputs[2789] = ~(layer0_outputs[4346]) | (layer0_outputs[3018]);
    assign layer1_outputs[2790] = (layer0_outputs[3670]) & ~(layer0_outputs[1759]);
    assign layer1_outputs[2791] = ~((layer0_outputs[3813]) & (layer0_outputs[2958]));
    assign layer1_outputs[2792] = (layer0_outputs[2762]) | (layer0_outputs[2785]);
    assign layer1_outputs[2793] = (layer0_outputs[4764]) & (layer0_outputs[2264]);
    assign layer1_outputs[2794] = ~(layer0_outputs[4024]) | (layer0_outputs[3287]);
    assign layer1_outputs[2795] = ~(layer0_outputs[464]) | (layer0_outputs[3990]);
    assign layer1_outputs[2796] = ~(layer0_outputs[497]);
    assign layer1_outputs[2797] = ~(layer0_outputs[3634]) | (layer0_outputs[2148]);
    assign layer1_outputs[2798] = ~(layer0_outputs[4751]);
    assign layer1_outputs[2799] = (layer0_outputs[1240]) | (layer0_outputs[2348]);
    assign layer1_outputs[2800] = 1'b0;
    assign layer1_outputs[2801] = ~(layer0_outputs[3057]);
    assign layer1_outputs[2802] = ~((layer0_outputs[1742]) | (layer0_outputs[3800]));
    assign layer1_outputs[2803] = (layer0_outputs[3031]) & ~(layer0_outputs[4901]);
    assign layer1_outputs[2804] = ~(layer0_outputs[3237]) | (layer0_outputs[1981]);
    assign layer1_outputs[2805] = ~((layer0_outputs[2898]) & (layer0_outputs[2239]));
    assign layer1_outputs[2806] = ~((layer0_outputs[378]) & (layer0_outputs[331]));
    assign layer1_outputs[2807] = (layer0_outputs[2679]) ^ (layer0_outputs[3439]);
    assign layer1_outputs[2808] = 1'b0;
    assign layer1_outputs[2809] = ~(layer0_outputs[4738]) | (layer0_outputs[4130]);
    assign layer1_outputs[2810] = ~((layer0_outputs[550]) ^ (layer0_outputs[4058]));
    assign layer1_outputs[2811] = (layer0_outputs[1330]) & ~(layer0_outputs[2891]);
    assign layer1_outputs[2812] = layer0_outputs[1036];
    assign layer1_outputs[2813] = (layer0_outputs[162]) & ~(layer0_outputs[64]);
    assign layer1_outputs[2814] = ~(layer0_outputs[1120]);
    assign layer1_outputs[2815] = ~(layer0_outputs[3206]);
    assign layer1_outputs[2816] = ~((layer0_outputs[680]) | (layer0_outputs[2676]));
    assign layer1_outputs[2817] = (layer0_outputs[885]) & ~(layer0_outputs[2691]);
    assign layer1_outputs[2818] = ~(layer0_outputs[2669]);
    assign layer1_outputs[2819] = (layer0_outputs[437]) | (layer0_outputs[4383]);
    assign layer1_outputs[2820] = (layer0_outputs[2683]) | (layer0_outputs[2144]);
    assign layer1_outputs[2821] = ~((layer0_outputs[2164]) & (layer0_outputs[3634]));
    assign layer1_outputs[2822] = layer0_outputs[1293];
    assign layer1_outputs[2823] = layer0_outputs[659];
    assign layer1_outputs[2824] = ~(layer0_outputs[3645]) | (layer0_outputs[1485]);
    assign layer1_outputs[2825] = ~(layer0_outputs[1213]);
    assign layer1_outputs[2826] = (layer0_outputs[2903]) & ~(layer0_outputs[1065]);
    assign layer1_outputs[2827] = layer0_outputs[1249];
    assign layer1_outputs[2828] = ~(layer0_outputs[1444]) | (layer0_outputs[4261]);
    assign layer1_outputs[2829] = 1'b0;
    assign layer1_outputs[2830] = (layer0_outputs[2252]) ^ (layer0_outputs[5083]);
    assign layer1_outputs[2831] = ~(layer0_outputs[1395]);
    assign layer1_outputs[2832] = layer0_outputs[485];
    assign layer1_outputs[2833] = (layer0_outputs[1415]) & ~(layer0_outputs[1209]);
    assign layer1_outputs[2834] = layer0_outputs[4703];
    assign layer1_outputs[2835] = 1'b0;
    assign layer1_outputs[2836] = ~(layer0_outputs[4987]);
    assign layer1_outputs[2837] = layer0_outputs[657];
    assign layer1_outputs[2838] = layer0_outputs[3201];
    assign layer1_outputs[2839] = (layer0_outputs[1557]) & ~(layer0_outputs[958]);
    assign layer1_outputs[2840] = (layer0_outputs[3854]) & (layer0_outputs[3974]);
    assign layer1_outputs[2841] = ~(layer0_outputs[4281]);
    assign layer1_outputs[2842] = 1'b0;
    assign layer1_outputs[2843] = layer0_outputs[3343];
    assign layer1_outputs[2844] = ~((layer0_outputs[200]) & (layer0_outputs[3598]));
    assign layer1_outputs[2845] = (layer0_outputs[4056]) & (layer0_outputs[4360]);
    assign layer1_outputs[2846] = ~((layer0_outputs[2703]) | (layer0_outputs[2962]));
    assign layer1_outputs[2847] = ~(layer0_outputs[1829]) | (layer0_outputs[4458]);
    assign layer1_outputs[2848] = ~((layer0_outputs[1868]) & (layer0_outputs[3529]));
    assign layer1_outputs[2849] = 1'b0;
    assign layer1_outputs[2850] = ~((layer0_outputs[5038]) ^ (layer0_outputs[3861]));
    assign layer1_outputs[2851] = 1'b0;
    assign layer1_outputs[2852] = ~(layer0_outputs[3069]);
    assign layer1_outputs[2853] = ~(layer0_outputs[3410]);
    assign layer1_outputs[2854] = ~(layer0_outputs[2414]) | (layer0_outputs[1660]);
    assign layer1_outputs[2855] = (layer0_outputs[86]) ^ (layer0_outputs[416]);
    assign layer1_outputs[2856] = (layer0_outputs[3405]) | (layer0_outputs[934]);
    assign layer1_outputs[2857] = (layer0_outputs[4817]) | (layer0_outputs[1675]);
    assign layer1_outputs[2858] = ~(layer0_outputs[996]) | (layer0_outputs[4985]);
    assign layer1_outputs[2859] = 1'b1;
    assign layer1_outputs[2860] = (layer0_outputs[2238]) | (layer0_outputs[1130]);
    assign layer1_outputs[2861] = ~(layer0_outputs[2545]);
    assign layer1_outputs[2862] = ~(layer0_outputs[248]) | (layer0_outputs[3294]);
    assign layer1_outputs[2863] = ~(layer0_outputs[3863]);
    assign layer1_outputs[2864] = (layer0_outputs[976]) & ~(layer0_outputs[1177]);
    assign layer1_outputs[2865] = 1'b0;
    assign layer1_outputs[2866] = layer0_outputs[4936];
    assign layer1_outputs[2867] = ~((layer0_outputs[511]) & (layer0_outputs[4656]));
    assign layer1_outputs[2868] = ~(layer0_outputs[3763]) | (layer0_outputs[1809]);
    assign layer1_outputs[2869] = ~((layer0_outputs[580]) | (layer0_outputs[4169]));
    assign layer1_outputs[2870] = 1'b1;
    assign layer1_outputs[2871] = ~(layer0_outputs[4246]);
    assign layer1_outputs[2872] = 1'b1;
    assign layer1_outputs[2873] = (layer0_outputs[4478]) & ~(layer0_outputs[2901]);
    assign layer1_outputs[2874] = (layer0_outputs[4109]) ^ (layer0_outputs[221]);
    assign layer1_outputs[2875] = ~(layer0_outputs[1561]);
    assign layer1_outputs[2876] = ~(layer0_outputs[3371]);
    assign layer1_outputs[2877] = 1'b1;
    assign layer1_outputs[2878] = (layer0_outputs[4057]) & ~(layer0_outputs[2789]);
    assign layer1_outputs[2879] = 1'b1;
    assign layer1_outputs[2880] = (layer0_outputs[5007]) & (layer0_outputs[2740]);
    assign layer1_outputs[2881] = ~((layer0_outputs[5062]) | (layer0_outputs[640]));
    assign layer1_outputs[2882] = ~(layer0_outputs[3644]) | (layer0_outputs[2293]);
    assign layer1_outputs[2883] = 1'b0;
    assign layer1_outputs[2884] = (layer0_outputs[894]) & ~(layer0_outputs[1715]);
    assign layer1_outputs[2885] = 1'b0;
    assign layer1_outputs[2886] = (layer0_outputs[298]) & ~(layer0_outputs[2849]);
    assign layer1_outputs[2887] = (layer0_outputs[1052]) ^ (layer0_outputs[1155]);
    assign layer1_outputs[2888] = (layer0_outputs[2180]) | (layer0_outputs[3273]);
    assign layer1_outputs[2889] = (layer0_outputs[2381]) & (layer0_outputs[3220]);
    assign layer1_outputs[2890] = (layer0_outputs[2756]) | (layer0_outputs[1415]);
    assign layer1_outputs[2891] = ~(layer0_outputs[2366]);
    assign layer1_outputs[2892] = ~((layer0_outputs[14]) | (layer0_outputs[776]));
    assign layer1_outputs[2893] = ~(layer0_outputs[830]);
    assign layer1_outputs[2894] = (layer0_outputs[2922]) & ~(layer0_outputs[393]);
    assign layer1_outputs[2895] = (layer0_outputs[1041]) & (layer0_outputs[3286]);
    assign layer1_outputs[2896] = 1'b1;
    assign layer1_outputs[2897] = layer0_outputs[1108];
    assign layer1_outputs[2898] = layer0_outputs[2595];
    assign layer1_outputs[2899] = 1'b1;
    assign layer1_outputs[2900] = 1'b1;
    assign layer1_outputs[2901] = ~(layer0_outputs[1064]) | (layer0_outputs[1386]);
    assign layer1_outputs[2902] = ~((layer0_outputs[70]) | (layer0_outputs[1217]));
    assign layer1_outputs[2903] = 1'b1;
    assign layer1_outputs[2904] = (layer0_outputs[4957]) & ~(layer0_outputs[1522]);
    assign layer1_outputs[2905] = 1'b0;
    assign layer1_outputs[2906] = ~(layer0_outputs[2726]) | (layer0_outputs[4405]);
    assign layer1_outputs[2907] = 1'b0;
    assign layer1_outputs[2908] = (layer0_outputs[4072]) & (layer0_outputs[2615]);
    assign layer1_outputs[2909] = (layer0_outputs[1316]) & ~(layer0_outputs[3315]);
    assign layer1_outputs[2910] = ~(layer0_outputs[4308]) | (layer0_outputs[2126]);
    assign layer1_outputs[2911] = (layer0_outputs[486]) & ~(layer0_outputs[1472]);
    assign layer1_outputs[2912] = (layer0_outputs[938]) & ~(layer0_outputs[3654]);
    assign layer1_outputs[2913] = 1'b0;
    assign layer1_outputs[2914] = layer0_outputs[3144];
    assign layer1_outputs[2915] = ~(layer0_outputs[1554]);
    assign layer1_outputs[2916] = ~(layer0_outputs[2299]);
    assign layer1_outputs[2917] = ~(layer0_outputs[3016]);
    assign layer1_outputs[2918] = (layer0_outputs[4285]) & (layer0_outputs[219]);
    assign layer1_outputs[2919] = ~(layer0_outputs[4008]) | (layer0_outputs[4534]);
    assign layer1_outputs[2920] = (layer0_outputs[3510]) & ~(layer0_outputs[255]);
    assign layer1_outputs[2921] = (layer0_outputs[1357]) & ~(layer0_outputs[2215]);
    assign layer1_outputs[2922] = ~(layer0_outputs[198]) | (layer0_outputs[1952]);
    assign layer1_outputs[2923] = ~(layer0_outputs[1814]) | (layer0_outputs[833]);
    assign layer1_outputs[2924] = 1'b1;
    assign layer1_outputs[2925] = 1'b0;
    assign layer1_outputs[2926] = ~(layer0_outputs[4243]);
    assign layer1_outputs[2927] = layer0_outputs[3400];
    assign layer1_outputs[2928] = ~(layer0_outputs[4691]);
    assign layer1_outputs[2929] = (layer0_outputs[294]) & (layer0_outputs[3115]);
    assign layer1_outputs[2930] = (layer0_outputs[3834]) & ~(layer0_outputs[943]);
    assign layer1_outputs[2931] = layer0_outputs[1739];
    assign layer1_outputs[2932] = ~(layer0_outputs[3246]);
    assign layer1_outputs[2933] = layer0_outputs[2420];
    assign layer1_outputs[2934] = (layer0_outputs[523]) & ~(layer0_outputs[2611]);
    assign layer1_outputs[2935] = ~(layer0_outputs[4859]) | (layer0_outputs[1145]);
    assign layer1_outputs[2936] = ~((layer0_outputs[1955]) ^ (layer0_outputs[1076]));
    assign layer1_outputs[2937] = 1'b1;
    assign layer1_outputs[2938] = (layer0_outputs[245]) & (layer0_outputs[1641]);
    assign layer1_outputs[2939] = ~(layer0_outputs[3772]) | (layer0_outputs[510]);
    assign layer1_outputs[2940] = (layer0_outputs[1687]) & ~(layer0_outputs[1222]);
    assign layer1_outputs[2941] = (layer0_outputs[2258]) | (layer0_outputs[2484]);
    assign layer1_outputs[2942] = ~(layer0_outputs[813]) | (layer0_outputs[2417]);
    assign layer1_outputs[2943] = (layer0_outputs[736]) & ~(layer0_outputs[1610]);
    assign layer1_outputs[2944] = 1'b0;
    assign layer1_outputs[2945] = layer0_outputs[2867];
    assign layer1_outputs[2946] = ~((layer0_outputs[3988]) & (layer0_outputs[4406]));
    assign layer1_outputs[2947] = (layer0_outputs[2052]) | (layer0_outputs[309]);
    assign layer1_outputs[2948] = ~(layer0_outputs[3692]) | (layer0_outputs[2623]);
    assign layer1_outputs[2949] = 1'b1;
    assign layer1_outputs[2950] = (layer0_outputs[2976]) | (layer0_outputs[1212]);
    assign layer1_outputs[2951] = ~((layer0_outputs[4274]) | (layer0_outputs[4716]));
    assign layer1_outputs[2952] = (layer0_outputs[4074]) & ~(layer0_outputs[3145]);
    assign layer1_outputs[2953] = (layer0_outputs[3117]) | (layer0_outputs[1665]);
    assign layer1_outputs[2954] = layer0_outputs[1115];
    assign layer1_outputs[2955] = ~((layer0_outputs[4184]) | (layer0_outputs[839]));
    assign layer1_outputs[2956] = ~(layer0_outputs[3071]);
    assign layer1_outputs[2957] = ~(layer0_outputs[3724]) | (layer0_outputs[2512]);
    assign layer1_outputs[2958] = layer0_outputs[3101];
    assign layer1_outputs[2959] = (layer0_outputs[3096]) & ~(layer0_outputs[3180]);
    assign layer1_outputs[2960] = (layer0_outputs[3917]) | (layer0_outputs[4741]);
    assign layer1_outputs[2961] = ~(layer0_outputs[3227]);
    assign layer1_outputs[2962] = ~(layer0_outputs[3705]) | (layer0_outputs[4318]);
    assign layer1_outputs[2963] = ~(layer0_outputs[4003]) | (layer0_outputs[1798]);
    assign layer1_outputs[2964] = ~(layer0_outputs[2207]) | (layer0_outputs[3029]);
    assign layer1_outputs[2965] = 1'b1;
    assign layer1_outputs[2966] = 1'b1;
    assign layer1_outputs[2967] = 1'b1;
    assign layer1_outputs[2968] = (layer0_outputs[4097]) & ~(layer0_outputs[4651]);
    assign layer1_outputs[2969] = (layer0_outputs[2674]) & (layer0_outputs[4662]);
    assign layer1_outputs[2970] = ~(layer0_outputs[600]) | (layer0_outputs[1659]);
    assign layer1_outputs[2971] = (layer0_outputs[3018]) & (layer0_outputs[3462]);
    assign layer1_outputs[2972] = ~((layer0_outputs[3632]) & (layer0_outputs[4978]));
    assign layer1_outputs[2973] = (layer0_outputs[1125]) & ~(layer0_outputs[4316]);
    assign layer1_outputs[2974] = (layer0_outputs[401]) & (layer0_outputs[3440]);
    assign layer1_outputs[2975] = ~((layer0_outputs[4393]) & (layer0_outputs[4187]));
    assign layer1_outputs[2976] = ~(layer0_outputs[4709]);
    assign layer1_outputs[2977] = ~(layer0_outputs[2193]) | (layer0_outputs[2390]);
    assign layer1_outputs[2978] = ~((layer0_outputs[2393]) & (layer0_outputs[555]));
    assign layer1_outputs[2979] = layer0_outputs[3367];
    assign layer1_outputs[2980] = 1'b1;
    assign layer1_outputs[2981] = ~(layer0_outputs[2372]);
    assign layer1_outputs[2982] = (layer0_outputs[4408]) | (layer0_outputs[3868]);
    assign layer1_outputs[2983] = (layer0_outputs[2109]) | (layer0_outputs[5078]);
    assign layer1_outputs[2984] = (layer0_outputs[2693]) & ~(layer0_outputs[730]);
    assign layer1_outputs[2985] = (layer0_outputs[2047]) & (layer0_outputs[3967]);
    assign layer1_outputs[2986] = 1'b1;
    assign layer1_outputs[2987] = 1'b1;
    assign layer1_outputs[2988] = ~(layer0_outputs[3341]);
    assign layer1_outputs[2989] = 1'b1;
    assign layer1_outputs[2990] = (layer0_outputs[2645]) & (layer0_outputs[3760]);
    assign layer1_outputs[2991] = (layer0_outputs[1714]) | (layer0_outputs[3765]);
    assign layer1_outputs[2992] = ~(layer0_outputs[2165]);
    assign layer1_outputs[2993] = ~(layer0_outputs[3924]) | (layer0_outputs[5021]);
    assign layer1_outputs[2994] = layer0_outputs[1873];
    assign layer1_outputs[2995] = 1'b0;
    assign layer1_outputs[2996] = (layer0_outputs[3345]) & ~(layer0_outputs[4459]);
    assign layer1_outputs[2997] = ~(layer0_outputs[2058]);
    assign layer1_outputs[2998] = (layer0_outputs[2273]) ^ (layer0_outputs[2447]);
    assign layer1_outputs[2999] = (layer0_outputs[494]) & ~(layer0_outputs[2388]);
    assign layer1_outputs[3000] = 1'b1;
    assign layer1_outputs[3001] = ~(layer0_outputs[2049]);
    assign layer1_outputs[3002] = (layer0_outputs[2964]) & ~(layer0_outputs[1585]);
    assign layer1_outputs[3003] = (layer0_outputs[4029]) & ~(layer0_outputs[4863]);
    assign layer1_outputs[3004] = layer0_outputs[2680];
    assign layer1_outputs[3005] = ~(layer0_outputs[869]) | (layer0_outputs[4363]);
    assign layer1_outputs[3006] = (layer0_outputs[3745]) & ~(layer0_outputs[1650]);
    assign layer1_outputs[3007] = (layer0_outputs[540]) ^ (layer0_outputs[2799]);
    assign layer1_outputs[3008] = (layer0_outputs[3946]) & ~(layer0_outputs[3733]);
    assign layer1_outputs[3009] = (layer0_outputs[1984]) & ~(layer0_outputs[641]);
    assign layer1_outputs[3010] = (layer0_outputs[1897]) & (layer0_outputs[3627]);
    assign layer1_outputs[3011] = 1'b0;
    assign layer1_outputs[3012] = 1'b0;
    assign layer1_outputs[3013] = 1'b1;
    assign layer1_outputs[3014] = layer0_outputs[105];
    assign layer1_outputs[3015] = (layer0_outputs[1473]) | (layer0_outputs[827]);
    assign layer1_outputs[3016] = (layer0_outputs[1515]) ^ (layer0_outputs[1121]);
    assign layer1_outputs[3017] = 1'b0;
    assign layer1_outputs[3018] = 1'b0;
    assign layer1_outputs[3019] = 1'b1;
    assign layer1_outputs[3020] = ~((layer0_outputs[2071]) & (layer0_outputs[284]));
    assign layer1_outputs[3021] = 1'b1;
    assign layer1_outputs[3022] = (layer0_outputs[3805]) & ~(layer0_outputs[1628]);
    assign layer1_outputs[3023] = ~((layer0_outputs[2325]) | (layer0_outputs[3753]));
    assign layer1_outputs[3024] = ~((layer0_outputs[4668]) | (layer0_outputs[2665]));
    assign layer1_outputs[3025] = ~((layer0_outputs[3857]) & (layer0_outputs[2061]));
    assign layer1_outputs[3026] = (layer0_outputs[4508]) | (layer0_outputs[2648]);
    assign layer1_outputs[3027] = (layer0_outputs[1639]) & (layer0_outputs[1513]);
    assign layer1_outputs[3028] = ~(layer0_outputs[1014]);
    assign layer1_outputs[3029] = (layer0_outputs[658]) | (layer0_outputs[2040]);
    assign layer1_outputs[3030] = ~(layer0_outputs[4376]) | (layer0_outputs[2825]);
    assign layer1_outputs[3031] = ~(layer0_outputs[1747]) | (layer0_outputs[92]);
    assign layer1_outputs[3032] = ~((layer0_outputs[395]) | (layer0_outputs[1669]));
    assign layer1_outputs[3033] = (layer0_outputs[4148]) & ~(layer0_outputs[2495]);
    assign layer1_outputs[3034] = ~(layer0_outputs[4780]);
    assign layer1_outputs[3035] = ~(layer0_outputs[2425]) | (layer0_outputs[4753]);
    assign layer1_outputs[3036] = (layer0_outputs[2960]) & (layer0_outputs[5092]);
    assign layer1_outputs[3037] = (layer0_outputs[4914]) ^ (layer0_outputs[24]);
    assign layer1_outputs[3038] = (layer0_outputs[2196]) & ~(layer0_outputs[820]);
    assign layer1_outputs[3039] = ~(layer0_outputs[2574]) | (layer0_outputs[1983]);
    assign layer1_outputs[3040] = ~((layer0_outputs[4260]) | (layer0_outputs[2553]));
    assign layer1_outputs[3041] = ~((layer0_outputs[176]) | (layer0_outputs[1959]));
    assign layer1_outputs[3042] = ~((layer0_outputs[3855]) | (layer0_outputs[5115]));
    assign layer1_outputs[3043] = ~((layer0_outputs[382]) | (layer0_outputs[2318]));
    assign layer1_outputs[3044] = 1'b1;
    assign layer1_outputs[3045] = 1'b0;
    assign layer1_outputs[3046] = 1'b0;
    assign layer1_outputs[3047] = 1'b1;
    assign layer1_outputs[3048] = ~(layer0_outputs[3274]);
    assign layer1_outputs[3049] = ~(layer0_outputs[1491]);
    assign layer1_outputs[3050] = ~(layer0_outputs[2246]) | (layer0_outputs[2477]);
    assign layer1_outputs[3051] = ~(layer0_outputs[4906]);
    assign layer1_outputs[3052] = ~((layer0_outputs[4350]) & (layer0_outputs[311]));
    assign layer1_outputs[3053] = ~((layer0_outputs[5114]) & (layer0_outputs[1510]));
    assign layer1_outputs[3054] = ~((layer0_outputs[3995]) | (layer0_outputs[2957]));
    assign layer1_outputs[3055] = layer0_outputs[145];
    assign layer1_outputs[3056] = ~((layer0_outputs[3252]) & (layer0_outputs[1831]));
    assign layer1_outputs[3057] = layer0_outputs[3329];
    assign layer1_outputs[3058] = ~(layer0_outputs[2874]) | (layer0_outputs[971]);
    assign layer1_outputs[3059] = ~(layer0_outputs[3773]);
    assign layer1_outputs[3060] = (layer0_outputs[2034]) | (layer0_outputs[3595]);
    assign layer1_outputs[3061] = (layer0_outputs[4205]) ^ (layer0_outputs[2968]);
    assign layer1_outputs[3062] = ~(layer0_outputs[3637]);
    assign layer1_outputs[3063] = ~(layer0_outputs[396]);
    assign layer1_outputs[3064] = ~(layer0_outputs[3947]) | (layer0_outputs[747]);
    assign layer1_outputs[3065] = ~(layer0_outputs[3475]);
    assign layer1_outputs[3066] = layer0_outputs[851];
    assign layer1_outputs[3067] = ~(layer0_outputs[1432]);
    assign layer1_outputs[3068] = ~(layer0_outputs[1156]);
    assign layer1_outputs[3069] = (layer0_outputs[2407]) ^ (layer0_outputs[4731]);
    assign layer1_outputs[3070] = 1'b1;
    assign layer1_outputs[3071] = (layer0_outputs[4719]) & ~(layer0_outputs[215]);
    assign layer1_outputs[3072] = 1'b0;
    assign layer1_outputs[3073] = layer0_outputs[5095];
    assign layer1_outputs[3074] = 1'b0;
    assign layer1_outputs[3075] = layer0_outputs[368];
    assign layer1_outputs[3076] = 1'b0;
    assign layer1_outputs[3077] = (layer0_outputs[498]) & (layer0_outputs[1330]);
    assign layer1_outputs[3078] = ~((layer0_outputs[382]) & (layer0_outputs[1989]));
    assign layer1_outputs[3079] = (layer0_outputs[4679]) & ~(layer0_outputs[4154]);
    assign layer1_outputs[3080] = (layer0_outputs[1077]) | (layer0_outputs[2396]);
    assign layer1_outputs[3081] = layer0_outputs[1140];
    assign layer1_outputs[3082] = ~(layer0_outputs[2736]) | (layer0_outputs[350]);
    assign layer1_outputs[3083] = ~(layer0_outputs[2396]);
    assign layer1_outputs[3084] = ~(layer0_outputs[765]);
    assign layer1_outputs[3085] = 1'b0;
    assign layer1_outputs[3086] = ~(layer0_outputs[3251]);
    assign layer1_outputs[3087] = (layer0_outputs[1149]) ^ (layer0_outputs[5064]);
    assign layer1_outputs[3088] = (layer0_outputs[2928]) & ~(layer0_outputs[1672]);
    assign layer1_outputs[3089] = (layer0_outputs[2539]) & ~(layer0_outputs[4937]);
    assign layer1_outputs[3090] = ~(layer0_outputs[3046]);
    assign layer1_outputs[3091] = layer0_outputs[4671];
    assign layer1_outputs[3092] = ~(layer0_outputs[1939]) | (layer0_outputs[894]);
    assign layer1_outputs[3093] = layer0_outputs[1408];
    assign layer1_outputs[3094] = layer0_outputs[2997];
    assign layer1_outputs[3095] = ~(layer0_outputs[539]);
    assign layer1_outputs[3096] = ~(layer0_outputs[963]);
    assign layer1_outputs[3097] = ~(layer0_outputs[4369]);
    assign layer1_outputs[3098] = ~(layer0_outputs[829]);
    assign layer1_outputs[3099] = (layer0_outputs[1397]) & ~(layer0_outputs[3973]);
    assign layer1_outputs[3100] = ~(layer0_outputs[4927]);
    assign layer1_outputs[3101] = ~(layer0_outputs[2919]) | (layer0_outputs[2219]);
    assign layer1_outputs[3102] = ~(layer0_outputs[1087]) | (layer0_outputs[727]);
    assign layer1_outputs[3103] = ~(layer0_outputs[2750]) | (layer0_outputs[3551]);
    assign layer1_outputs[3104] = ~(layer0_outputs[189]) | (layer0_outputs[1822]);
    assign layer1_outputs[3105] = 1'b1;
    assign layer1_outputs[3106] = 1'b1;
    assign layer1_outputs[3107] = layer0_outputs[4518];
    assign layer1_outputs[3108] = (layer0_outputs[3392]) & (layer0_outputs[4170]);
    assign layer1_outputs[3109] = ~((layer0_outputs[4868]) ^ (layer0_outputs[3306]));
    assign layer1_outputs[3110] = ~(layer0_outputs[4591]) | (layer0_outputs[767]);
    assign layer1_outputs[3111] = (layer0_outputs[206]) & ~(layer0_outputs[327]);
    assign layer1_outputs[3112] = layer0_outputs[3012];
    assign layer1_outputs[3113] = ~(layer0_outputs[2596]) | (layer0_outputs[1035]);
    assign layer1_outputs[3114] = (layer0_outputs[1279]) & (layer0_outputs[854]);
    assign layer1_outputs[3115] = (layer0_outputs[3295]) & ~(layer0_outputs[3424]);
    assign layer1_outputs[3116] = ~(layer0_outputs[1430]);
    assign layer1_outputs[3117] = layer0_outputs[4853];
    assign layer1_outputs[3118] = (layer0_outputs[2975]) ^ (layer0_outputs[4805]);
    assign layer1_outputs[3119] = (layer0_outputs[200]) & ~(layer0_outputs[4162]);
    assign layer1_outputs[3120] = 1'b0;
    assign layer1_outputs[3121] = ~((layer0_outputs[3372]) | (layer0_outputs[3186]));
    assign layer1_outputs[3122] = ~(layer0_outputs[2744]);
    assign layer1_outputs[3123] = 1'b1;
    assign layer1_outputs[3124] = 1'b1;
    assign layer1_outputs[3125] = (layer0_outputs[257]) & ~(layer0_outputs[3130]);
    assign layer1_outputs[3126] = layer0_outputs[4127];
    assign layer1_outputs[3127] = layer0_outputs[4273];
    assign layer1_outputs[3128] = ~((layer0_outputs[589]) | (layer0_outputs[3677]));
    assign layer1_outputs[3129] = (layer0_outputs[1382]) | (layer0_outputs[3538]);
    assign layer1_outputs[3130] = 1'b1;
    assign layer1_outputs[3131] = (layer0_outputs[5050]) & ~(layer0_outputs[3638]);
    assign layer1_outputs[3132] = (layer0_outputs[3709]) & (layer0_outputs[4259]);
    assign layer1_outputs[3133] = ~(layer0_outputs[1090]);
    assign layer1_outputs[3134] = (layer0_outputs[4289]) & (layer0_outputs[2499]);
    assign layer1_outputs[3135] = (layer0_outputs[4405]) & (layer0_outputs[4525]);
    assign layer1_outputs[3136] = layer0_outputs[1449];
    assign layer1_outputs[3137] = ~(layer0_outputs[2930]) | (layer0_outputs[1594]);
    assign layer1_outputs[3138] = ~((layer0_outputs[849]) & (layer0_outputs[2755]));
    assign layer1_outputs[3139] = ~(layer0_outputs[4050]);
    assign layer1_outputs[3140] = (layer0_outputs[5104]) ^ (layer0_outputs[4086]);
    assign layer1_outputs[3141] = (layer0_outputs[2137]) & ~(layer0_outputs[2321]);
    assign layer1_outputs[3142] = layer0_outputs[2065];
    assign layer1_outputs[3143] = ~(layer0_outputs[3704]);
    assign layer1_outputs[3144] = (layer0_outputs[4038]) & ~(layer0_outputs[1708]);
    assign layer1_outputs[3145] = (layer0_outputs[1009]) | (layer0_outputs[2515]);
    assign layer1_outputs[3146] = 1'b0;
    assign layer1_outputs[3147] = ~((layer0_outputs[1600]) | (layer0_outputs[1558]));
    assign layer1_outputs[3148] = (layer0_outputs[3188]) & (layer0_outputs[3871]);
    assign layer1_outputs[3149] = (layer0_outputs[1556]) | (layer0_outputs[289]);
    assign layer1_outputs[3150] = layer0_outputs[1995];
    assign layer1_outputs[3151] = (layer0_outputs[1214]) & ~(layer0_outputs[4064]);
    assign layer1_outputs[3152] = ~(layer0_outputs[4548]) | (layer0_outputs[1152]);
    assign layer1_outputs[3153] = 1'b1;
    assign layer1_outputs[3154] = ~((layer0_outputs[641]) | (layer0_outputs[337]));
    assign layer1_outputs[3155] = 1'b0;
    assign layer1_outputs[3156] = ~((layer0_outputs[2841]) & (layer0_outputs[1043]));
    assign layer1_outputs[3157] = ~(layer0_outputs[3331]);
    assign layer1_outputs[3158] = ~(layer0_outputs[4475]);
    assign layer1_outputs[3159] = layer0_outputs[4451];
    assign layer1_outputs[3160] = ~(layer0_outputs[4735]) | (layer0_outputs[3882]);
    assign layer1_outputs[3161] = ~((layer0_outputs[1879]) | (layer0_outputs[2567]));
    assign layer1_outputs[3162] = layer0_outputs[3525];
    assign layer1_outputs[3163] = (layer0_outputs[3999]) & ~(layer0_outputs[708]);
    assign layer1_outputs[3164] = ~(layer0_outputs[1819]);
    assign layer1_outputs[3165] = (layer0_outputs[3470]) & ~(layer0_outputs[1534]);
    assign layer1_outputs[3166] = (layer0_outputs[512]) & (layer0_outputs[4311]);
    assign layer1_outputs[3167] = 1'b1;
    assign layer1_outputs[3168] = (layer0_outputs[1808]) & ~(layer0_outputs[2750]);
    assign layer1_outputs[3169] = ~(layer0_outputs[4043]);
    assign layer1_outputs[3170] = ~(layer0_outputs[3333]);
    assign layer1_outputs[3171] = ~((layer0_outputs[566]) & (layer0_outputs[585]));
    assign layer1_outputs[3172] = ~(layer0_outputs[2465]);
    assign layer1_outputs[3173] = (layer0_outputs[1294]) & (layer0_outputs[4159]);
    assign layer1_outputs[3174] = (layer0_outputs[3688]) & ~(layer0_outputs[4256]);
    assign layer1_outputs[3175] = (layer0_outputs[1786]) & (layer0_outputs[4119]);
    assign layer1_outputs[3176] = ~((layer0_outputs[3645]) | (layer0_outputs[1047]));
    assign layer1_outputs[3177] = layer0_outputs[3334];
    assign layer1_outputs[3178] = ~((layer0_outputs[4816]) & (layer0_outputs[1117]));
    assign layer1_outputs[3179] = layer0_outputs[4822];
    assign layer1_outputs[3180] = 1'b0;
    assign layer1_outputs[3181] = 1'b0;
    assign layer1_outputs[3182] = layer0_outputs[1447];
    assign layer1_outputs[3183] = ~(layer0_outputs[2607]);
    assign layer1_outputs[3184] = (layer0_outputs[2304]) | (layer0_outputs[4544]);
    assign layer1_outputs[3185] = ~((layer0_outputs[2688]) & (layer0_outputs[2072]));
    assign layer1_outputs[3186] = ~((layer0_outputs[2601]) | (layer0_outputs[1693]));
    assign layer1_outputs[3187] = layer0_outputs[1135];
    assign layer1_outputs[3188] = ~((layer0_outputs[4699]) | (layer0_outputs[1573]));
    assign layer1_outputs[3189] = ~(layer0_outputs[3944]) | (layer0_outputs[2559]);
    assign layer1_outputs[3190] = layer0_outputs[1727];
    assign layer1_outputs[3191] = layer0_outputs[2274];
    assign layer1_outputs[3192] = ~(layer0_outputs[133]) | (layer0_outputs[4546]);
    assign layer1_outputs[3193] = layer0_outputs[823];
    assign layer1_outputs[3194] = (layer0_outputs[771]) & ~(layer0_outputs[1633]);
    assign layer1_outputs[3195] = (layer0_outputs[2624]) & ~(layer0_outputs[1688]);
    assign layer1_outputs[3196] = layer0_outputs[4396];
    assign layer1_outputs[3197] = layer0_outputs[249];
    assign layer1_outputs[3198] = layer0_outputs[2783];
    assign layer1_outputs[3199] = (layer0_outputs[1935]) & (layer0_outputs[3929]);
    assign layer1_outputs[3200] = ~((layer0_outputs[3874]) & (layer0_outputs[5019]));
    assign layer1_outputs[3201] = (layer0_outputs[490]) & (layer0_outputs[2698]);
    assign layer1_outputs[3202] = ~(layer0_outputs[3910]) | (layer0_outputs[1654]);
    assign layer1_outputs[3203] = layer0_outputs[633];
    assign layer1_outputs[3204] = ~((layer0_outputs[3515]) ^ (layer0_outputs[712]));
    assign layer1_outputs[3205] = ~((layer0_outputs[4645]) & (layer0_outputs[1758]));
    assign layer1_outputs[3206] = (layer0_outputs[1909]) | (layer0_outputs[1334]);
    assign layer1_outputs[3207] = (layer0_outputs[3513]) ^ (layer0_outputs[3555]);
    assign layer1_outputs[3208] = layer0_outputs[473];
    assign layer1_outputs[3209] = ~((layer0_outputs[1433]) & (layer0_outputs[4181]));
    assign layer1_outputs[3210] = 1'b1;
    assign layer1_outputs[3211] = 1'b0;
    assign layer1_outputs[3212] = layer0_outputs[4759];
    assign layer1_outputs[3213] = (layer0_outputs[1465]) & (layer0_outputs[2483]);
    assign layer1_outputs[3214] = ~((layer0_outputs[758]) | (layer0_outputs[883]));
    assign layer1_outputs[3215] = (layer0_outputs[2913]) & ~(layer0_outputs[4809]);
    assign layer1_outputs[3216] = layer0_outputs[2644];
    assign layer1_outputs[3217] = layer0_outputs[1195];
    assign layer1_outputs[3218] = layer0_outputs[4490];
    assign layer1_outputs[3219] = ~(layer0_outputs[3651]);
    assign layer1_outputs[3220] = 1'b1;
    assign layer1_outputs[3221] = layer0_outputs[2234];
    assign layer1_outputs[3222] = layer0_outputs[2494];
    assign layer1_outputs[3223] = (layer0_outputs[2454]) | (layer0_outputs[4484]);
    assign layer1_outputs[3224] = layer0_outputs[1311];
    assign layer1_outputs[3225] = 1'b0;
    assign layer1_outputs[3226] = ~(layer0_outputs[619]) | (layer0_outputs[2796]);
    assign layer1_outputs[3227] = ~(layer0_outputs[1011]);
    assign layer1_outputs[3228] = ~(layer0_outputs[302]) | (layer0_outputs[1734]);
    assign layer1_outputs[3229] = 1'b0;
    assign layer1_outputs[3230] = ~(layer0_outputs[2636]) | (layer0_outputs[3952]);
    assign layer1_outputs[3231] = 1'b0;
    assign layer1_outputs[3232] = layer0_outputs[2592];
    assign layer1_outputs[3233] = ~(layer0_outputs[4850]);
    assign layer1_outputs[3234] = ~(layer0_outputs[3593]) | (layer0_outputs[1533]);
    assign layer1_outputs[3235] = 1'b0;
    assign layer1_outputs[3236] = ~(layer0_outputs[4111]) | (layer0_outputs[2804]);
    assign layer1_outputs[3237] = ~((layer0_outputs[291]) | (layer0_outputs[478]));
    assign layer1_outputs[3238] = 1'b0;
    assign layer1_outputs[3239] = layer0_outputs[4340];
    assign layer1_outputs[3240] = (layer0_outputs[997]) | (layer0_outputs[1279]);
    assign layer1_outputs[3241] = ~((layer0_outputs[265]) | (layer0_outputs[955]));
    assign layer1_outputs[3242] = layer0_outputs[2458];
    assign layer1_outputs[3243] = (layer0_outputs[3737]) & (layer0_outputs[1022]);
    assign layer1_outputs[3244] = ~(layer0_outputs[3114]) | (layer0_outputs[504]);
    assign layer1_outputs[3245] = ~(layer0_outputs[3530]) | (layer0_outputs[85]);
    assign layer1_outputs[3246] = ~((layer0_outputs[4171]) ^ (layer0_outputs[3355]));
    assign layer1_outputs[3247] = (layer0_outputs[2749]) & (layer0_outputs[4178]);
    assign layer1_outputs[3248] = ~(layer0_outputs[1613]) | (layer0_outputs[77]);
    assign layer1_outputs[3249] = (layer0_outputs[367]) & ~(layer0_outputs[506]);
    assign layer1_outputs[3250] = ~((layer0_outputs[4993]) | (layer0_outputs[155]));
    assign layer1_outputs[3251] = (layer0_outputs[1257]) & ~(layer0_outputs[961]);
    assign layer1_outputs[3252] = ~((layer0_outputs[495]) & (layer0_outputs[3461]));
    assign layer1_outputs[3253] = (layer0_outputs[3145]) & ~(layer0_outputs[1591]);
    assign layer1_outputs[3254] = (layer0_outputs[3076]) | (layer0_outputs[1692]);
    assign layer1_outputs[3255] = ~(layer0_outputs[2971]);
    assign layer1_outputs[3256] = (layer0_outputs[3778]) & ~(layer0_outputs[1181]);
    assign layer1_outputs[3257] = ~(layer0_outputs[832]) | (layer0_outputs[4468]);
    assign layer1_outputs[3258] = (layer0_outputs[1801]) & ~(layer0_outputs[1185]);
    assign layer1_outputs[3259] = ~(layer0_outputs[1142]);
    assign layer1_outputs[3260] = (layer0_outputs[346]) & ~(layer0_outputs[4998]);
    assign layer1_outputs[3261] = 1'b1;
    assign layer1_outputs[3262] = ~((layer0_outputs[3840]) & (layer0_outputs[1746]));
    assign layer1_outputs[3263] = layer0_outputs[1184];
    assign layer1_outputs[3264] = layer0_outputs[1852];
    assign layer1_outputs[3265] = layer0_outputs[880];
    assign layer1_outputs[3266] = layer0_outputs[113];
    assign layer1_outputs[3267] = ~(layer0_outputs[3021]) | (layer0_outputs[217]);
    assign layer1_outputs[3268] = ~((layer0_outputs[3335]) & (layer0_outputs[1817]));
    assign layer1_outputs[3269] = ~(layer0_outputs[3324]) | (layer0_outputs[15]);
    assign layer1_outputs[3270] = ~(layer0_outputs[1144]);
    assign layer1_outputs[3271] = (layer0_outputs[2627]) & ~(layer0_outputs[4040]);
    assign layer1_outputs[3272] = 1'b1;
    assign layer1_outputs[3273] = ~((layer0_outputs[484]) | (layer0_outputs[4411]));
    assign layer1_outputs[3274] = 1'b1;
    assign layer1_outputs[3275] = layer0_outputs[661];
    assign layer1_outputs[3276] = ~(layer0_outputs[4201]) | (layer0_outputs[554]);
    assign layer1_outputs[3277] = (layer0_outputs[5060]) & ~(layer0_outputs[4641]);
    assign layer1_outputs[3278] = (layer0_outputs[1518]) | (layer0_outputs[2206]);
    assign layer1_outputs[3279] = ~(layer0_outputs[4181]);
    assign layer1_outputs[3280] = ~(layer0_outputs[3160]) | (layer0_outputs[4090]);
    assign layer1_outputs[3281] = (layer0_outputs[5006]) | (layer0_outputs[1741]);
    assign layer1_outputs[3282] = (layer0_outputs[390]) & (layer0_outputs[2697]);
    assign layer1_outputs[3283] = 1'b0;
    assign layer1_outputs[3284] = (layer0_outputs[3999]) & (layer0_outputs[4460]);
    assign layer1_outputs[3285] = (layer0_outputs[186]) | (layer0_outputs[2884]);
    assign layer1_outputs[3286] = ~((layer0_outputs[690]) ^ (layer0_outputs[2933]));
    assign layer1_outputs[3287] = layer0_outputs[4865];
    assign layer1_outputs[3288] = ~((layer0_outputs[1271]) | (layer0_outputs[2759]));
    assign layer1_outputs[3289] = ~((layer0_outputs[1161]) | (layer0_outputs[3441]));
    assign layer1_outputs[3290] = ~(layer0_outputs[1707]) | (layer0_outputs[2070]);
    assign layer1_outputs[3291] = (layer0_outputs[1662]) & ~(layer0_outputs[4809]);
    assign layer1_outputs[3292] = ~(layer0_outputs[438]);
    assign layer1_outputs[3293] = (layer0_outputs[1988]) & (layer0_outputs[1868]);
    assign layer1_outputs[3294] = (layer0_outputs[450]) & ~(layer0_outputs[570]);
    assign layer1_outputs[3295] = (layer0_outputs[3846]) | (layer0_outputs[3799]);
    assign layer1_outputs[3296] = (layer0_outputs[558]) & ~(layer0_outputs[4559]);
    assign layer1_outputs[3297] = layer0_outputs[4054];
    assign layer1_outputs[3298] = ~((layer0_outputs[868]) | (layer0_outputs[3768]));
    assign layer1_outputs[3299] = layer0_outputs[4726];
    assign layer1_outputs[3300] = (layer0_outputs[4805]) & ~(layer0_outputs[4187]);
    assign layer1_outputs[3301] = 1'b1;
    assign layer1_outputs[3302] = (layer0_outputs[907]) & ~(layer0_outputs[775]);
    assign layer1_outputs[3303] = (layer0_outputs[3741]) & (layer0_outputs[3122]);
    assign layer1_outputs[3304] = 1'b1;
    assign layer1_outputs[3305] = (layer0_outputs[3175]) | (layer0_outputs[436]);
    assign layer1_outputs[3306] = (layer0_outputs[288]) & (layer0_outputs[491]);
    assign layer1_outputs[3307] = ~(layer0_outputs[3241]) | (layer0_outputs[4716]);
    assign layer1_outputs[3308] = ~(layer0_outputs[3278]);
    assign layer1_outputs[3309] = 1'b0;
    assign layer1_outputs[3310] = layer0_outputs[1569];
    assign layer1_outputs[3311] = ~(layer0_outputs[2046]) | (layer0_outputs[2164]);
    assign layer1_outputs[3312] = ~(layer0_outputs[1174]);
    assign layer1_outputs[3313] = ~(layer0_outputs[2648]) | (layer0_outputs[2456]);
    assign layer1_outputs[3314] = ~(layer0_outputs[3937]) | (layer0_outputs[3533]);
    assign layer1_outputs[3315] = ~(layer0_outputs[886]) | (layer0_outputs[3399]);
    assign layer1_outputs[3316] = 1'b0;
    assign layer1_outputs[3317] = (layer0_outputs[1033]) & (layer0_outputs[1835]);
    assign layer1_outputs[3318] = (layer0_outputs[1067]) & ~(layer0_outputs[4481]);
    assign layer1_outputs[3319] = (layer0_outputs[3395]) & (layer0_outputs[923]);
    assign layer1_outputs[3320] = 1'b1;
    assign layer1_outputs[3321] = (layer0_outputs[530]) & ~(layer0_outputs[1997]);
    assign layer1_outputs[3322] = 1'b1;
    assign layer1_outputs[3323] = (layer0_outputs[602]) ^ (layer0_outputs[3759]);
    assign layer1_outputs[3324] = ~(layer0_outputs[3532]);
    assign layer1_outputs[3325] = (layer0_outputs[3392]) | (layer0_outputs[3455]);
    assign layer1_outputs[3326] = ~(layer0_outputs[3234]);
    assign layer1_outputs[3327] = ~(layer0_outputs[2379]);
    assign layer1_outputs[3328] = layer0_outputs[4001];
    assign layer1_outputs[3329] = ~(layer0_outputs[1016]) | (layer0_outputs[1302]);
    assign layer1_outputs[3330] = (layer0_outputs[2520]) | (layer0_outputs[644]);
    assign layer1_outputs[3331] = 1'b1;
    assign layer1_outputs[3332] = ~((layer0_outputs[4167]) | (layer0_outputs[1985]));
    assign layer1_outputs[3333] = (layer0_outputs[184]) & (layer0_outputs[1834]);
    assign layer1_outputs[3334] = ~(layer0_outputs[3948]) | (layer0_outputs[1062]);
    assign layer1_outputs[3335] = layer0_outputs[2082];
    assign layer1_outputs[3336] = (layer0_outputs[1844]) & ~(layer0_outputs[3739]);
    assign layer1_outputs[3337] = ~((layer0_outputs[325]) & (layer0_outputs[282]));
    assign layer1_outputs[3338] = ~(layer0_outputs[1784]);
    assign layer1_outputs[3339] = ~(layer0_outputs[4570]);
    assign layer1_outputs[3340] = ~((layer0_outputs[3482]) ^ (layer0_outputs[34]));
    assign layer1_outputs[3341] = layer0_outputs[3189];
    assign layer1_outputs[3342] = ~(layer0_outputs[4118]);
    assign layer1_outputs[3343] = (layer0_outputs[1795]) & ~(layer0_outputs[4836]);
    assign layer1_outputs[3344] = ~((layer0_outputs[1328]) & (layer0_outputs[1237]));
    assign layer1_outputs[3345] = ~(layer0_outputs[458]);
    assign layer1_outputs[3346] = (layer0_outputs[3279]) & (layer0_outputs[4228]);
    assign layer1_outputs[3347] = layer0_outputs[632];
    assign layer1_outputs[3348] = 1'b0;
    assign layer1_outputs[3349] = ~(layer0_outputs[3821]) | (layer0_outputs[1681]);
    assign layer1_outputs[3350] = ~((layer0_outputs[2659]) & (layer0_outputs[3266]));
    assign layer1_outputs[3351] = 1'b0;
    assign layer1_outputs[3352] = (layer0_outputs[3067]) & ~(layer0_outputs[1981]);
    assign layer1_outputs[3353] = ~((layer0_outputs[2714]) | (layer0_outputs[3350]));
    assign layer1_outputs[3354] = ~(layer0_outputs[2374]) | (layer0_outputs[713]);
    assign layer1_outputs[3355] = ~((layer0_outputs[2312]) | (layer0_outputs[4734]));
    assign layer1_outputs[3356] = (layer0_outputs[1806]) & ~(layer0_outputs[625]);
    assign layer1_outputs[3357] = ~((layer0_outputs[3235]) | (layer0_outputs[4725]));
    assign layer1_outputs[3358] = layer0_outputs[3812];
    assign layer1_outputs[3359] = layer0_outputs[2269];
    assign layer1_outputs[3360] = (layer0_outputs[2603]) & ~(layer0_outputs[876]);
    assign layer1_outputs[3361] = ~(layer0_outputs[804]) | (layer0_outputs[3301]);
    assign layer1_outputs[3362] = ~(layer0_outputs[2655]) | (layer0_outputs[2593]);
    assign layer1_outputs[3363] = (layer0_outputs[4890]) & ~(layer0_outputs[4462]);
    assign layer1_outputs[3364] = ~(layer0_outputs[739]);
    assign layer1_outputs[3365] = (layer0_outputs[4141]) & ~(layer0_outputs[1949]);
    assign layer1_outputs[3366] = ~(layer0_outputs[262]);
    assign layer1_outputs[3367] = ~(layer0_outputs[1967]) | (layer0_outputs[625]);
    assign layer1_outputs[3368] = layer0_outputs[4033];
    assign layer1_outputs[3369] = layer0_outputs[4367];
    assign layer1_outputs[3370] = ~(layer0_outputs[4938]);
    assign layer1_outputs[3371] = 1'b0;
    assign layer1_outputs[3372] = (layer0_outputs[1702]) & ~(layer0_outputs[1936]);
    assign layer1_outputs[3373] = ~((layer0_outputs[1821]) & (layer0_outputs[42]));
    assign layer1_outputs[3374] = ~(layer0_outputs[603]) | (layer0_outputs[3458]);
    assign layer1_outputs[3375] = ~((layer0_outputs[1677]) | (layer0_outputs[4236]));
    assign layer1_outputs[3376] = ~((layer0_outputs[223]) & (layer0_outputs[4325]));
    assign layer1_outputs[3377] = 1'b1;
    assign layer1_outputs[3378] = ~(layer0_outputs[2522]) | (layer0_outputs[2194]);
    assign layer1_outputs[3379] = layer0_outputs[4335];
    assign layer1_outputs[3380] = 1'b0;
    assign layer1_outputs[3381] = ~(layer0_outputs[3605]);
    assign layer1_outputs[3382] = (layer0_outputs[3960]) ^ (layer0_outputs[3732]);
    assign layer1_outputs[3383] = 1'b1;
    assign layer1_outputs[3384] = 1'b1;
    assign layer1_outputs[3385] = ~((layer0_outputs[673]) | (layer0_outputs[84]));
    assign layer1_outputs[3386] = ~(layer0_outputs[3638]) | (layer0_outputs[1494]);
    assign layer1_outputs[3387] = 1'b0;
    assign layer1_outputs[3388] = ~(layer0_outputs[2213]) | (layer0_outputs[2224]);
    assign layer1_outputs[3389] = layer0_outputs[695];
    assign layer1_outputs[3390] = ~(layer0_outputs[2701]) | (layer0_outputs[247]);
    assign layer1_outputs[3391] = (layer0_outputs[158]) & ~(layer0_outputs[1354]);
    assign layer1_outputs[3392] = ~(layer0_outputs[4192]) | (layer0_outputs[3986]);
    assign layer1_outputs[3393] = (layer0_outputs[2059]) & (layer0_outputs[1922]);
    assign layer1_outputs[3394] = (layer0_outputs[926]) & (layer0_outputs[2710]);
    assign layer1_outputs[3395] = layer0_outputs[590];
    assign layer1_outputs[3396] = ~(layer0_outputs[2743]);
    assign layer1_outputs[3397] = ~(layer0_outputs[1554]);
    assign layer1_outputs[3398] = ~((layer0_outputs[4597]) | (layer0_outputs[366]));
    assign layer1_outputs[3399] = ~(layer0_outputs[1528]);
    assign layer1_outputs[3400] = layer0_outputs[3649];
    assign layer1_outputs[3401] = (layer0_outputs[683]) | (layer0_outputs[4255]);
    assign layer1_outputs[3402] = (layer0_outputs[536]) & (layer0_outputs[2852]);
    assign layer1_outputs[3403] = 1'b0;
    assign layer1_outputs[3404] = (layer0_outputs[4659]) & (layer0_outputs[2479]);
    assign layer1_outputs[3405] = 1'b1;
    assign layer1_outputs[3406] = ~(layer0_outputs[2856]) | (layer0_outputs[3521]);
    assign layer1_outputs[3407] = (layer0_outputs[4603]) ^ (layer0_outputs[2056]);
    assign layer1_outputs[3408] = (layer0_outputs[100]) | (layer0_outputs[3299]);
    assign layer1_outputs[3409] = ~(layer0_outputs[3070]);
    assign layer1_outputs[3410] = ~(layer0_outputs[2822]);
    assign layer1_outputs[3411] = ~(layer0_outputs[972]);
    assign layer1_outputs[3412] = (layer0_outputs[4794]) & ~(layer0_outputs[2428]);
    assign layer1_outputs[3413] = ~((layer0_outputs[4939]) ^ (layer0_outputs[993]));
    assign layer1_outputs[3414] = ~(layer0_outputs[107]);
    assign layer1_outputs[3415] = ~(layer0_outputs[4147]) | (layer0_outputs[4889]);
    assign layer1_outputs[3416] = 1'b1;
    assign layer1_outputs[3417] = (layer0_outputs[902]) ^ (layer0_outputs[505]);
    assign layer1_outputs[3418] = (layer0_outputs[3950]) & ~(layer0_outputs[4920]);
    assign layer1_outputs[3419] = 1'b1;
    assign layer1_outputs[3420] = ~((layer0_outputs[4994]) | (layer0_outputs[763]));
    assign layer1_outputs[3421] = (layer0_outputs[2973]) & ~(layer0_outputs[2242]);
    assign layer1_outputs[3422] = (layer0_outputs[3400]) & (layer0_outputs[1274]);
    assign layer1_outputs[3423] = ~((layer0_outputs[1362]) | (layer0_outputs[4802]));
    assign layer1_outputs[3424] = layer0_outputs[4714];
    assign layer1_outputs[3425] = ~(layer0_outputs[3106]);
    assign layer1_outputs[3426] = ~(layer0_outputs[2700]) | (layer0_outputs[3465]);
    assign layer1_outputs[3427] = 1'b0;
    assign layer1_outputs[3428] = 1'b0;
    assign layer1_outputs[3429] = 1'b1;
    assign layer1_outputs[3430] = ~((layer0_outputs[1670]) & (layer0_outputs[2701]));
    assign layer1_outputs[3431] = 1'b1;
    assign layer1_outputs[3432] = layer0_outputs[4273];
    assign layer1_outputs[3433] = 1'b1;
    assign layer1_outputs[3434] = layer0_outputs[1647];
    assign layer1_outputs[3435] = ~(layer0_outputs[3245]) | (layer0_outputs[4376]);
    assign layer1_outputs[3436] = (layer0_outputs[1938]) & ~(layer0_outputs[6]);
    assign layer1_outputs[3437] = ~((layer0_outputs[4128]) & (layer0_outputs[3517]));
    assign layer1_outputs[3438] = ~(layer0_outputs[662]);
    assign layer1_outputs[3439] = ~((layer0_outputs[49]) & (layer0_outputs[1986]));
    assign layer1_outputs[3440] = ~(layer0_outputs[1226]) | (layer0_outputs[1122]);
    assign layer1_outputs[3441] = ~(layer0_outputs[1042]);
    assign layer1_outputs[3442] = 1'b0;
    assign layer1_outputs[3443] = ~((layer0_outputs[4496]) ^ (layer0_outputs[862]));
    assign layer1_outputs[3444] = (layer0_outputs[1760]) | (layer0_outputs[620]);
    assign layer1_outputs[3445] = (layer0_outputs[1788]) & ~(layer0_outputs[2067]);
    assign layer1_outputs[3446] = layer0_outputs[3180];
    assign layer1_outputs[3447] = 1'b1;
    assign layer1_outputs[3448] = 1'b0;
    assign layer1_outputs[3449] = ~(layer0_outputs[1479]) | (layer0_outputs[58]);
    assign layer1_outputs[3450] = ~(layer0_outputs[1398]) | (layer0_outputs[3174]);
    assign layer1_outputs[3451] = 1'b1;
    assign layer1_outputs[3452] = ~(layer0_outputs[1627]);
    assign layer1_outputs[3453] = ~(layer0_outputs[4954]) | (layer0_outputs[1750]);
    assign layer1_outputs[3454] = (layer0_outputs[726]) & ~(layer0_outputs[1061]);
    assign layer1_outputs[3455] = 1'b0;
    assign layer1_outputs[3456] = 1'b0;
    assign layer1_outputs[3457] = ~(layer0_outputs[2378]) | (layer0_outputs[236]);
    assign layer1_outputs[3458] = (layer0_outputs[171]) & (layer0_outputs[4392]);
    assign layer1_outputs[3459] = ~(layer0_outputs[1624]);
    assign layer1_outputs[3460] = (layer0_outputs[2392]) & ~(layer0_outputs[5040]);
    assign layer1_outputs[3461] = layer0_outputs[2176];
    assign layer1_outputs[3462] = ~((layer0_outputs[3586]) | (layer0_outputs[1022]));
    assign layer1_outputs[3463] = (layer0_outputs[1722]) & ~(layer0_outputs[4133]);
    assign layer1_outputs[3464] = layer0_outputs[3276];
    assign layer1_outputs[3465] = ~(layer0_outputs[4268]) | (layer0_outputs[4444]);
    assign layer1_outputs[3466] = ~(layer0_outputs[4449]) | (layer0_outputs[4175]);
    assign layer1_outputs[3467] = 1'b1;
    assign layer1_outputs[3468] = ~((layer0_outputs[77]) & (layer0_outputs[2525]));
    assign layer1_outputs[3469] = ~(layer0_outputs[4497]) | (layer0_outputs[260]);
    assign layer1_outputs[3470] = (layer0_outputs[789]) & ~(layer0_outputs[4234]);
    assign layer1_outputs[3471] = layer0_outputs[2847];
    assign layer1_outputs[3472] = ~(layer0_outputs[2217]);
    assign layer1_outputs[3473] = ~(layer0_outputs[2632]) | (layer0_outputs[240]);
    assign layer1_outputs[3474] = (layer0_outputs[218]) | (layer0_outputs[2044]);
    assign layer1_outputs[3475] = ~(layer0_outputs[1198]) | (layer0_outputs[420]);
    assign layer1_outputs[3476] = ~(layer0_outputs[1075]) | (layer0_outputs[3359]);
    assign layer1_outputs[3477] = ~(layer0_outputs[3793]) | (layer0_outputs[3605]);
    assign layer1_outputs[3478] = (layer0_outputs[4593]) & (layer0_outputs[3082]);
    assign layer1_outputs[3479] = (layer0_outputs[4070]) & ~(layer0_outputs[4119]);
    assign layer1_outputs[3480] = ~(layer0_outputs[4229]);
    assign layer1_outputs[3481] = layer0_outputs[4489];
    assign layer1_outputs[3482] = 1'b1;
    assign layer1_outputs[3483] = ~(layer0_outputs[2764]) | (layer0_outputs[3437]);
    assign layer1_outputs[3484] = 1'b0;
    assign layer1_outputs[3485] = (layer0_outputs[3196]) | (layer0_outputs[5021]);
    assign layer1_outputs[3486] = ~((layer0_outputs[1877]) & (layer0_outputs[731]));
    assign layer1_outputs[3487] = layer0_outputs[2048];
    assign layer1_outputs[3488] = (layer0_outputs[6]) ^ (layer0_outputs[687]);
    assign layer1_outputs[3489] = (layer0_outputs[1046]) | (layer0_outputs[3102]);
    assign layer1_outputs[3490] = ~((layer0_outputs[3015]) & (layer0_outputs[1159]));
    assign layer1_outputs[3491] = (layer0_outputs[4846]) | (layer0_outputs[274]);
    assign layer1_outputs[3492] = layer0_outputs[2445];
    assign layer1_outputs[3493] = 1'b0;
    assign layer1_outputs[3494] = (layer0_outputs[4067]) & ~(layer0_outputs[4768]);
    assign layer1_outputs[3495] = layer0_outputs[333];
    assign layer1_outputs[3496] = 1'b0;
    assign layer1_outputs[3497] = (layer0_outputs[1157]) & ~(layer0_outputs[4210]);
    assign layer1_outputs[3498] = (layer0_outputs[1862]) & ~(layer0_outputs[2287]);
    assign layer1_outputs[3499] = (layer0_outputs[4276]) & ~(layer0_outputs[4588]);
    assign layer1_outputs[3500] = (layer0_outputs[354]) & ~(layer0_outputs[3473]);
    assign layer1_outputs[3501] = 1'b0;
    assign layer1_outputs[3502] = (layer0_outputs[3222]) & ~(layer0_outputs[2947]);
    assign layer1_outputs[3503] = 1'b0;
    assign layer1_outputs[3504] = ~(layer0_outputs[1446]) | (layer0_outputs[3464]);
    assign layer1_outputs[3505] = ~((layer0_outputs[533]) & (layer0_outputs[4562]));
    assign layer1_outputs[3506] = ~(layer0_outputs[4469]) | (layer0_outputs[2007]);
    assign layer1_outputs[3507] = ~(layer0_outputs[2481]) | (layer0_outputs[2623]);
    assign layer1_outputs[3508] = 1'b0;
    assign layer1_outputs[3509] = (layer0_outputs[1445]) | (layer0_outputs[3613]);
    assign layer1_outputs[3510] = layer0_outputs[2887];
    assign layer1_outputs[3511] = ~((layer0_outputs[4831]) & (layer0_outputs[3430]));
    assign layer1_outputs[3512] = (layer0_outputs[2386]) & ~(layer0_outputs[1021]);
    assign layer1_outputs[3513] = ~((layer0_outputs[3013]) | (layer0_outputs[1448]));
    assign layer1_outputs[3514] = layer0_outputs[4103];
    assign layer1_outputs[3515] = ~((layer0_outputs[2334]) & (layer0_outputs[4650]));
    assign layer1_outputs[3516] = 1'b1;
    assign layer1_outputs[3517] = (layer0_outputs[4932]) & ~(layer0_outputs[3878]);
    assign layer1_outputs[3518] = (layer0_outputs[2035]) & ~(layer0_outputs[463]);
    assign layer1_outputs[3519] = ~(layer0_outputs[3407]) | (layer0_outputs[4739]);
    assign layer1_outputs[3520] = (layer0_outputs[4505]) & ~(layer0_outputs[781]);
    assign layer1_outputs[3521] = ~((layer0_outputs[3639]) ^ (layer0_outputs[373]));
    assign layer1_outputs[3522] = ~(layer0_outputs[4177]) | (layer0_outputs[4923]);
    assign layer1_outputs[3523] = (layer0_outputs[55]) & (layer0_outputs[4900]);
    assign layer1_outputs[3524] = ~(layer0_outputs[1313]);
    assign layer1_outputs[3525] = 1'b1;
    assign layer1_outputs[3526] = layer0_outputs[3338];
    assign layer1_outputs[3527] = 1'b0;
    assign layer1_outputs[3528] = ~((layer0_outputs[3597]) & (layer0_outputs[1041]));
    assign layer1_outputs[3529] = (layer0_outputs[1303]) | (layer0_outputs[3672]);
    assign layer1_outputs[3530] = ~(layer0_outputs[1190]);
    assign layer1_outputs[3531] = ~((layer0_outputs[3457]) & (layer0_outputs[1038]));
    assign layer1_outputs[3532] = ~(layer0_outputs[2979]);
    assign layer1_outputs[3533] = (layer0_outputs[4174]) & ~(layer0_outputs[4176]);
    assign layer1_outputs[3534] = (layer0_outputs[2267]) & ~(layer0_outputs[4889]);
    assign layer1_outputs[3535] = layer0_outputs[1625];
    assign layer1_outputs[3536] = 1'b0;
    assign layer1_outputs[3537] = (layer0_outputs[3389]) & (layer0_outputs[4956]);
    assign layer1_outputs[3538] = ~(layer0_outputs[4979]) | (layer0_outputs[4825]);
    assign layer1_outputs[3539] = layer0_outputs[4793];
    assign layer1_outputs[3540] = ~(layer0_outputs[4535]);
    assign layer1_outputs[3541] = (layer0_outputs[1802]) & ~(layer0_outputs[4634]);
    assign layer1_outputs[3542] = ~(layer0_outputs[3131]) | (layer0_outputs[1442]);
    assign layer1_outputs[3543] = ~(layer0_outputs[2814]);
    assign layer1_outputs[3544] = layer0_outputs[4537];
    assign layer1_outputs[3545] = layer0_outputs[4772];
    assign layer1_outputs[3546] = ~(layer0_outputs[4565]) | (layer0_outputs[3596]);
    assign layer1_outputs[3547] = (layer0_outputs[2255]) & ~(layer0_outputs[3663]);
    assign layer1_outputs[3548] = ~(layer0_outputs[3662]) | (layer0_outputs[1037]);
    assign layer1_outputs[3549] = 1'b1;
    assign layer1_outputs[3550] = ~(layer0_outputs[2462]) | (layer0_outputs[2843]);
    assign layer1_outputs[3551] = 1'b1;
    assign layer1_outputs[3552] = ~(layer0_outputs[1860]) | (layer0_outputs[4310]);
    assign layer1_outputs[3553] = ~(layer0_outputs[110]) | (layer0_outputs[3058]);
    assign layer1_outputs[3554] = ~((layer0_outputs[2506]) | (layer0_outputs[4047]));
    assign layer1_outputs[3555] = (layer0_outputs[3693]) | (layer0_outputs[2973]);
    assign layer1_outputs[3556] = layer0_outputs[392];
    assign layer1_outputs[3557] = ~(layer0_outputs[1911]) | (layer0_outputs[1293]);
    assign layer1_outputs[3558] = layer0_outputs[3925];
    assign layer1_outputs[3559] = (layer0_outputs[4674]) & ~(layer0_outputs[3878]);
    assign layer1_outputs[3560] = 1'b1;
    assign layer1_outputs[3561] = (layer0_outputs[49]) & ~(layer0_outputs[1722]);
    assign layer1_outputs[3562] = (layer0_outputs[2757]) & ~(layer0_outputs[1148]);
    assign layer1_outputs[3563] = ~((layer0_outputs[411]) | (layer0_outputs[3179]));
    assign layer1_outputs[3564] = (layer0_outputs[2079]) | (layer0_outputs[3701]);
    assign layer1_outputs[3565] = 1'b0;
    assign layer1_outputs[3566] = ~(layer0_outputs[2439]);
    assign layer1_outputs[3567] = layer0_outputs[925];
    assign layer1_outputs[3568] = (layer0_outputs[3618]) | (layer0_outputs[4621]);
    assign layer1_outputs[3569] = (layer0_outputs[4383]) | (layer0_outputs[3545]);
    assign layer1_outputs[3570] = 1'b1;
    assign layer1_outputs[3571] = ~(layer0_outputs[800]);
    assign layer1_outputs[3572] = ~((layer0_outputs[664]) ^ (layer0_outputs[1805]));
    assign layer1_outputs[3573] = ~((layer0_outputs[1447]) ^ (layer0_outputs[428]));
    assign layer1_outputs[3574] = ~(layer0_outputs[2072]);
    assign layer1_outputs[3575] = ~((layer0_outputs[836]) & (layer0_outputs[2478]));
    assign layer1_outputs[3576] = ~(layer0_outputs[4752]);
    assign layer1_outputs[3577] = (layer0_outputs[3162]) | (layer0_outputs[837]);
    assign layer1_outputs[3578] = 1'b1;
    assign layer1_outputs[3579] = (layer0_outputs[5089]) & ~(layer0_outputs[3713]);
    assign layer1_outputs[3580] = (layer0_outputs[1036]) & ~(layer0_outputs[4246]);
    assign layer1_outputs[3581] = (layer0_outputs[1508]) & ~(layer0_outputs[284]);
    assign layer1_outputs[3582] = ~(layer0_outputs[2037]);
    assign layer1_outputs[3583] = layer0_outputs[4578];
    assign layer1_outputs[3584] = 1'b1;
    assign layer1_outputs[3585] = layer0_outputs[2771];
    assign layer1_outputs[3586] = ~((layer0_outputs[3091]) | (layer0_outputs[321]));
    assign layer1_outputs[3587] = layer0_outputs[508];
    assign layer1_outputs[3588] = ~((layer0_outputs[1376]) | (layer0_outputs[560]));
    assign layer1_outputs[3589] = (layer0_outputs[3408]) | (layer0_outputs[3899]);
    assign layer1_outputs[3590] = ~(layer0_outputs[965]) | (layer0_outputs[4059]);
    assign layer1_outputs[3591] = layer0_outputs[487];
    assign layer1_outputs[3592] = ~(layer0_outputs[2240]) | (layer0_outputs[1561]);
    assign layer1_outputs[3593] = layer0_outputs[4143];
    assign layer1_outputs[3594] = ~((layer0_outputs[4855]) ^ (layer0_outputs[4622]));
    assign layer1_outputs[3595] = layer0_outputs[1921];
    assign layer1_outputs[3596] = ~(layer0_outputs[694]) | (layer0_outputs[633]);
    assign layer1_outputs[3597] = ~(layer0_outputs[1848]) | (layer0_outputs[1940]);
    assign layer1_outputs[3598] = 1'b0;
    assign layer1_outputs[3599] = (layer0_outputs[4122]) ^ (layer0_outputs[2370]);
    assign layer1_outputs[3600] = (layer0_outputs[2095]) & (layer0_outputs[2758]);
    assign layer1_outputs[3601] = ~((layer0_outputs[1662]) & (layer0_outputs[4796]));
    assign layer1_outputs[3602] = 1'b0;
    assign layer1_outputs[3603] = 1'b1;
    assign layer1_outputs[3604] = 1'b0;
    assign layer1_outputs[3605] = ~(layer0_outputs[2092]);
    assign layer1_outputs[3606] = ~((layer0_outputs[3321]) & (layer0_outputs[1304]));
    assign layer1_outputs[3607] = (layer0_outputs[4527]) & (layer0_outputs[5081]);
    assign layer1_outputs[3608] = layer0_outputs[2469];
    assign layer1_outputs[3609] = ~(layer0_outputs[4958]);
    assign layer1_outputs[3610] = layer0_outputs[807];
    assign layer1_outputs[3611] = ~(layer0_outputs[3729]) | (layer0_outputs[618]);
    assign layer1_outputs[3612] = (layer0_outputs[2473]) | (layer0_outputs[2938]);
    assign layer1_outputs[3613] = ~(layer0_outputs[5099]);
    assign layer1_outputs[3614] = ~((layer0_outputs[3836]) | (layer0_outputs[4447]));
    assign layer1_outputs[3615] = 1'b1;
    assign layer1_outputs[3616] = 1'b1;
    assign layer1_outputs[3617] = layer0_outputs[5008];
    assign layer1_outputs[3618] = (layer0_outputs[3611]) & (layer0_outputs[4810]);
    assign layer1_outputs[3619] = ~((layer0_outputs[1856]) | (layer0_outputs[5119]));
    assign layer1_outputs[3620] = layer0_outputs[5116];
    assign layer1_outputs[3621] = layer0_outputs[5058];
    assign layer1_outputs[3622] = (layer0_outputs[928]) | (layer0_outputs[1444]);
    assign layer1_outputs[3623] = layer0_outputs[2662];
    assign layer1_outputs[3624] = 1'b1;
    assign layer1_outputs[3625] = ~(layer0_outputs[4586]) | (layer0_outputs[3202]);
    assign layer1_outputs[3626] = ~((layer0_outputs[4284]) ^ (layer0_outputs[4144]));
    assign layer1_outputs[3627] = ~(layer0_outputs[1547]);
    assign layer1_outputs[3628] = ~(layer0_outputs[3982]);
    assign layer1_outputs[3629] = layer0_outputs[1975];
    assign layer1_outputs[3630] = (layer0_outputs[1207]) & ~(layer0_outputs[4374]);
    assign layer1_outputs[3631] = (layer0_outputs[4579]) & ~(layer0_outputs[4051]);
    assign layer1_outputs[3632] = (layer0_outputs[1641]) & (layer0_outputs[1310]);
    assign layer1_outputs[3633] = layer0_outputs[4280];
    assign layer1_outputs[3634] = layer0_outputs[2352];
    assign layer1_outputs[3635] = ~(layer0_outputs[421]) | (layer0_outputs[637]);
    assign layer1_outputs[3636] = layer0_outputs[3073];
    assign layer1_outputs[3637] = layer0_outputs[4700];
    assign layer1_outputs[3638] = (layer0_outputs[2232]) & ~(layer0_outputs[4251]);
    assign layer1_outputs[3639] = ~(layer0_outputs[439]);
    assign layer1_outputs[3640] = 1'b1;
    assign layer1_outputs[3641] = ~(layer0_outputs[2219]);
    assign layer1_outputs[3642] = 1'b0;
    assign layer1_outputs[3643] = (layer0_outputs[409]) & ~(layer0_outputs[3463]);
    assign layer1_outputs[3644] = ~((layer0_outputs[3340]) | (layer0_outputs[3056]));
    assign layer1_outputs[3645] = layer0_outputs[4684];
    assign layer1_outputs[3646] = ~((layer0_outputs[4219]) & (layer0_outputs[1481]));
    assign layer1_outputs[3647] = (layer0_outputs[1863]) | (layer0_outputs[2994]);
    assign layer1_outputs[3648] = ~((layer0_outputs[4329]) | (layer0_outputs[2643]));
    assign layer1_outputs[3649] = layer0_outputs[359];
    assign layer1_outputs[3650] = 1'b0;
    assign layer1_outputs[3651] = (layer0_outputs[666]) & ~(layer0_outputs[2885]);
    assign layer1_outputs[3652] = layer0_outputs[631];
    assign layer1_outputs[3653] = (layer0_outputs[4500]) ^ (layer0_outputs[2027]);
    assign layer1_outputs[3654] = layer0_outputs[2136];
    assign layer1_outputs[3655] = (layer0_outputs[1441]) | (layer0_outputs[1107]);
    assign layer1_outputs[3656] = layer0_outputs[4148];
    assign layer1_outputs[3657] = 1'b0;
    assign layer1_outputs[3658] = ~(layer0_outputs[2854]) | (layer0_outputs[452]);
    assign layer1_outputs[3659] = (layer0_outputs[5045]) & ~(layer0_outputs[2836]);
    assign layer1_outputs[3660] = ~((layer0_outputs[3567]) ^ (layer0_outputs[2116]));
    assign layer1_outputs[3661] = ~(layer0_outputs[1891]) | (layer0_outputs[4395]);
    assign layer1_outputs[3662] = ~(layer0_outputs[2693]) | (layer0_outputs[1471]);
    assign layer1_outputs[3663] = layer0_outputs[4920];
    assign layer1_outputs[3664] = ~(layer0_outputs[3508]) | (layer0_outputs[4226]);
    assign layer1_outputs[3665] = ~(layer0_outputs[4572]) | (layer0_outputs[1466]);
    assign layer1_outputs[3666] = ~((layer0_outputs[4903]) & (layer0_outputs[610]));
    assign layer1_outputs[3667] = (layer0_outputs[2834]) & ~(layer0_outputs[1870]);
    assign layer1_outputs[3668] = 1'b1;
    assign layer1_outputs[3669] = ~(layer0_outputs[75]);
    assign layer1_outputs[3670] = ~(layer0_outputs[2332]) | (layer0_outputs[97]);
    assign layer1_outputs[3671] = (layer0_outputs[3664]) | (layer0_outputs[1813]);
    assign layer1_outputs[3672] = 1'b1;
    assign layer1_outputs[3673] = (layer0_outputs[83]) & ~(layer0_outputs[3201]);
    assign layer1_outputs[3674] = ~(layer0_outputs[1466]);
    assign layer1_outputs[3675] = ~((layer0_outputs[1635]) & (layer0_outputs[87]));
    assign layer1_outputs[3676] = layer0_outputs[307];
    assign layer1_outputs[3677] = ~(layer0_outputs[863]);
    assign layer1_outputs[3678] = (layer0_outputs[3991]) & ~(layer0_outputs[2133]);
    assign layer1_outputs[3679] = ~(layer0_outputs[2446]) | (layer0_outputs[4774]);
    assign layer1_outputs[3680] = ~(layer0_outputs[4886]);
    assign layer1_outputs[3681] = ~((layer0_outputs[3779]) & (layer0_outputs[4940]));
    assign layer1_outputs[3682] = ~(layer0_outputs[4097]) | (layer0_outputs[807]);
    assign layer1_outputs[3683] = 1'b0;
    assign layer1_outputs[3684] = ~(layer0_outputs[649]);
    assign layer1_outputs[3685] = ~(layer0_outputs[1749]);
    assign layer1_outputs[3686] = (layer0_outputs[2510]) | (layer0_outputs[749]);
    assign layer1_outputs[3687] = layer0_outputs[4017];
    assign layer1_outputs[3688] = (layer0_outputs[2721]) & ~(layer0_outputs[3006]);
    assign layer1_outputs[3689] = 1'b1;
    assign layer1_outputs[3690] = ~(layer0_outputs[2022]) | (layer0_outputs[837]);
    assign layer1_outputs[3691] = layer0_outputs[4818];
    assign layer1_outputs[3692] = ~((layer0_outputs[569]) | (layer0_outputs[3134]));
    assign layer1_outputs[3693] = ~(layer0_outputs[3234]);
    assign layer1_outputs[3694] = ~(layer0_outputs[3750]);
    assign layer1_outputs[3695] = layer0_outputs[5033];
    assign layer1_outputs[3696] = (layer0_outputs[856]) & ~(layer0_outputs[1150]);
    assign layer1_outputs[3697] = (layer0_outputs[4433]) & ~(layer0_outputs[4840]);
    assign layer1_outputs[3698] = (layer0_outputs[978]) & ~(layer0_outputs[4137]);
    assign layer1_outputs[3699] = layer0_outputs[4882];
    assign layer1_outputs[3700] = ~((layer0_outputs[2395]) | (layer0_outputs[3677]));
    assign layer1_outputs[3701] = ~(layer0_outputs[905]) | (layer0_outputs[2806]);
    assign layer1_outputs[3702] = ~(layer0_outputs[810]) | (layer0_outputs[2564]);
    assign layer1_outputs[3703] = ~(layer0_outputs[4314]) | (layer0_outputs[1683]);
    assign layer1_outputs[3704] = (layer0_outputs[419]) & (layer0_outputs[314]);
    assign layer1_outputs[3705] = 1'b0;
    assign layer1_outputs[3706] = (layer0_outputs[5]) ^ (layer0_outputs[4503]);
    assign layer1_outputs[3707] = (layer0_outputs[3500]) & (layer0_outputs[711]);
    assign layer1_outputs[3708] = ~((layer0_outputs[2406]) | (layer0_outputs[4723]));
    assign layer1_outputs[3709] = ~((layer0_outputs[877]) ^ (layer0_outputs[878]));
    assign layer1_outputs[3710] = layer0_outputs[1420];
    assign layer1_outputs[3711] = 1'b0;
    assign layer1_outputs[3712] = ~(layer0_outputs[5051]) | (layer0_outputs[4404]);
    assign layer1_outputs[3713] = (layer0_outputs[3847]) & ~(layer0_outputs[814]);
    assign layer1_outputs[3714] = ~((layer0_outputs[2248]) | (layer0_outputs[3037]));
    assign layer1_outputs[3715] = layer0_outputs[653];
    assign layer1_outputs[3716] = (layer0_outputs[2461]) | (layer0_outputs[2260]);
    assign layer1_outputs[3717] = ~(layer0_outputs[3880]) | (layer0_outputs[1040]);
    assign layer1_outputs[3718] = ~((layer0_outputs[3360]) & (layer0_outputs[2315]));
    assign layer1_outputs[3719] = (layer0_outputs[1170]) & ~(layer0_outputs[730]);
    assign layer1_outputs[3720] = ~(layer0_outputs[4884]);
    assign layer1_outputs[3721] = (layer0_outputs[1908]) & (layer0_outputs[4345]);
    assign layer1_outputs[3722] = layer0_outputs[3187];
    assign layer1_outputs[3723] = ~(layer0_outputs[3054]);
    assign layer1_outputs[3724] = (layer0_outputs[4536]) & ~(layer0_outputs[541]);
    assign layer1_outputs[3725] = layer0_outputs[1914];
    assign layer1_outputs[3726] = ~(layer0_outputs[4419]) | (layer0_outputs[4968]);
    assign layer1_outputs[3727] = ~(layer0_outputs[4096]) | (layer0_outputs[2892]);
    assign layer1_outputs[3728] = ~(layer0_outputs[2309]) | (layer0_outputs[1521]);
    assign layer1_outputs[3729] = ~((layer0_outputs[1283]) ^ (layer0_outputs[1339]));
    assign layer1_outputs[3730] = (layer0_outputs[3726]) & (layer0_outputs[2614]);
    assign layer1_outputs[3731] = layer0_outputs[640];
    assign layer1_outputs[3732] = (layer0_outputs[2328]) & ~(layer0_outputs[2439]);
    assign layer1_outputs[3733] = ~(layer0_outputs[384]);
    assign layer1_outputs[3734] = layer0_outputs[389];
    assign layer1_outputs[3735] = 1'b0;
    assign layer1_outputs[3736] = ~(layer0_outputs[1395]) | (layer0_outputs[3035]);
    assign layer1_outputs[3737] = (layer0_outputs[1701]) & (layer0_outputs[4202]);
    assign layer1_outputs[3738] = layer0_outputs[826];
    assign layer1_outputs[3739] = ~(layer0_outputs[3460]);
    assign layer1_outputs[3740] = (layer0_outputs[430]) & ~(layer0_outputs[3723]);
    assign layer1_outputs[3741] = layer0_outputs[1085];
    assign layer1_outputs[3742] = ~((layer0_outputs[2031]) & (layer0_outputs[953]));
    assign layer1_outputs[3743] = layer0_outputs[3428];
    assign layer1_outputs[3744] = layer0_outputs[2390];
    assign layer1_outputs[3745] = ~(layer0_outputs[4628]);
    assign layer1_outputs[3746] = ~(layer0_outputs[1311]) | (layer0_outputs[1469]);
    assign layer1_outputs[3747] = ~(layer0_outputs[1010]);
    assign layer1_outputs[3748] = layer0_outputs[3270];
    assign layer1_outputs[3749] = ~((layer0_outputs[2613]) ^ (layer0_outputs[99]));
    assign layer1_outputs[3750] = ~(layer0_outputs[3177]);
    assign layer1_outputs[3751] = ~((layer0_outputs[2900]) & (layer0_outputs[3495]));
    assign layer1_outputs[3752] = (layer0_outputs[2136]) & (layer0_outputs[2742]);
    assign layer1_outputs[3753] = 1'b1;
    assign layer1_outputs[3754] = 1'b1;
    assign layer1_outputs[3755] = 1'b1;
    assign layer1_outputs[3756] = ~((layer0_outputs[1560]) & (layer0_outputs[2614]));
    assign layer1_outputs[3757] = layer0_outputs[2815];
    assign layer1_outputs[3758] = ~(layer0_outputs[4861]);
    assign layer1_outputs[3759] = ~(layer0_outputs[39]);
    assign layer1_outputs[3760] = ~((layer0_outputs[4059]) | (layer0_outputs[4858]));
    assign layer1_outputs[3761] = ~((layer0_outputs[4302]) | (layer0_outputs[709]));
    assign layer1_outputs[3762] = 1'b0;
    assign layer1_outputs[3763] = ~(layer0_outputs[1541]);
    assign layer1_outputs[3764] = (layer0_outputs[3066]) & ~(layer0_outputs[2381]);
    assign layer1_outputs[3765] = ~(layer0_outputs[2793]) | (layer0_outputs[1205]);
    assign layer1_outputs[3766] = 1'b1;
    assign layer1_outputs[3767] = ~(layer0_outputs[4378]) | (layer0_outputs[4108]);
    assign layer1_outputs[3768] = (layer0_outputs[715]) | (layer0_outputs[171]);
    assign layer1_outputs[3769] = (layer0_outputs[2671]) & ~(layer0_outputs[1435]);
    assign layer1_outputs[3770] = 1'b0;
    assign layer1_outputs[3771] = (layer0_outputs[3846]) & ~(layer0_outputs[4829]);
    assign layer1_outputs[3772] = ~(layer0_outputs[2532]);
    assign layer1_outputs[3773] = ~(layer0_outputs[4652]) | (layer0_outputs[1731]);
    assign layer1_outputs[3774] = (layer0_outputs[2854]) | (layer0_outputs[429]);
    assign layer1_outputs[3775] = ~((layer0_outputs[3025]) & (layer0_outputs[4552]));
    assign layer1_outputs[3776] = (layer0_outputs[2203]) & (layer0_outputs[1297]);
    assign layer1_outputs[3777] = ~(layer0_outputs[4426]);
    assign layer1_outputs[3778] = ~((layer0_outputs[1067]) ^ (layer0_outputs[1418]));
    assign layer1_outputs[3779] = layer0_outputs[3324];
    assign layer1_outputs[3780] = layer0_outputs[2313];
    assign layer1_outputs[3781] = ~(layer0_outputs[2437]);
    assign layer1_outputs[3782] = ~((layer0_outputs[411]) | (layer0_outputs[2826]));
    assign layer1_outputs[3783] = (layer0_outputs[996]) & (layer0_outputs[3606]);
    assign layer1_outputs[3784] = ~(layer0_outputs[3393]);
    assign layer1_outputs[3785] = 1'b0;
    assign layer1_outputs[3786] = (layer0_outputs[733]) | (layer0_outputs[3026]);
    assign layer1_outputs[3787] = (layer0_outputs[2360]) & ~(layer0_outputs[5082]);
    assign layer1_outputs[3788] = layer0_outputs[182];
    assign layer1_outputs[3789] = ~((layer0_outputs[3977]) ^ (layer0_outputs[614]));
    assign layer1_outputs[3790] = layer0_outputs[4152];
    assign layer1_outputs[3791] = (layer0_outputs[864]) & ~(layer0_outputs[4498]);
    assign layer1_outputs[3792] = ~((layer0_outputs[2306]) | (layer0_outputs[842]));
    assign layer1_outputs[3793] = ~(layer0_outputs[656]) | (layer0_outputs[2968]);
    assign layer1_outputs[3794] = ~(layer0_outputs[995]) | (layer0_outputs[2558]);
    assign layer1_outputs[3795] = (layer0_outputs[2415]) | (layer0_outputs[2195]);
    assign layer1_outputs[3796] = ~(layer0_outputs[2811]);
    assign layer1_outputs[3797] = 1'b0;
    assign layer1_outputs[3798] = (layer0_outputs[4602]) & ~(layer0_outputs[2959]);
    assign layer1_outputs[3799] = ~((layer0_outputs[4827]) & (layer0_outputs[3272]));
    assign layer1_outputs[3800] = ~((layer0_outputs[4940]) ^ (layer0_outputs[2855]));
    assign layer1_outputs[3801] = ~(layer0_outputs[5023]);
    assign layer1_outputs[3802] = layer0_outputs[4132];
    assign layer1_outputs[3803] = ~(layer0_outputs[4616]);
    assign layer1_outputs[3804] = ~(layer0_outputs[842]) | (layer0_outputs[2068]);
    assign layer1_outputs[3805] = 1'b0;
    assign layer1_outputs[3806] = ~((layer0_outputs[4998]) | (layer0_outputs[4768]));
    assign layer1_outputs[3807] = ~(layer0_outputs[3928]) | (layer0_outputs[3870]);
    assign layer1_outputs[3808] = ~((layer0_outputs[2685]) & (layer0_outputs[193]));
    assign layer1_outputs[3809] = ~(layer0_outputs[824]) | (layer0_outputs[1591]);
    assign layer1_outputs[3810] = ~(layer0_outputs[2709]);
    assign layer1_outputs[3811] = (layer0_outputs[2904]) | (layer0_outputs[2569]);
    assign layer1_outputs[3812] = ~(layer0_outputs[2184]) | (layer0_outputs[4306]);
    assign layer1_outputs[3813] = ~(layer0_outputs[217]);
    assign layer1_outputs[3814] = (layer0_outputs[2901]) & ~(layer0_outputs[3592]);
    assign layer1_outputs[3815] = ~(layer0_outputs[2956]);
    assign layer1_outputs[3816] = (layer0_outputs[3668]) & (layer0_outputs[2932]);
    assign layer1_outputs[3817] = layer0_outputs[1080];
    assign layer1_outputs[3818] = ~(layer0_outputs[388]) | (layer0_outputs[3068]);
    assign layer1_outputs[3819] = (layer0_outputs[3196]) & ~(layer0_outputs[744]);
    assign layer1_outputs[3820] = layer0_outputs[1101];
    assign layer1_outputs[3821] = layer0_outputs[1958];
    assign layer1_outputs[3822] = (layer0_outputs[3094]) & ~(layer0_outputs[1432]);
    assign layer1_outputs[3823] = (layer0_outputs[3829]) & ~(layer0_outputs[3712]);
    assign layer1_outputs[3824] = 1'b0;
    assign layer1_outputs[3825] = ~((layer0_outputs[1427]) | (layer0_outputs[4138]));
    assign layer1_outputs[3826] = 1'b1;
    assign layer1_outputs[3827] = ~(layer0_outputs[2590]);
    assign layer1_outputs[3828] = 1'b1;
    assign layer1_outputs[3829] = layer0_outputs[3459];
    assign layer1_outputs[3830] = (layer0_outputs[1599]) & ~(layer0_outputs[2696]);
    assign layer1_outputs[3831] = (layer0_outputs[1406]) & ~(layer0_outputs[4318]);
    assign layer1_outputs[3832] = (layer0_outputs[743]) & ~(layer0_outputs[1455]);
    assign layer1_outputs[3833] = 1'b1;
    assign layer1_outputs[3834] = layer0_outputs[3097];
    assign layer1_outputs[3835] = ~((layer0_outputs[1576]) & (layer0_outputs[425]));
    assign layer1_outputs[3836] = layer0_outputs[69];
    assign layer1_outputs[3837] = 1'b0;
    assign layer1_outputs[3838] = ~((layer0_outputs[320]) & (layer0_outputs[906]));
    assign layer1_outputs[3839] = ~((layer0_outputs[3964]) | (layer0_outputs[3413]));
    assign layer1_outputs[3840] = 1'b1;
    assign layer1_outputs[3841] = ~((layer0_outputs[4095]) ^ (layer0_outputs[3789]));
    assign layer1_outputs[3842] = (layer0_outputs[4108]) & ~(layer0_outputs[4466]);
    assign layer1_outputs[3843] = ~((layer0_outputs[3761]) & (layer0_outputs[1723]));
    assign layer1_outputs[3844] = (layer0_outputs[4737]) & ~(layer0_outputs[1502]);
    assign layer1_outputs[3845] = (layer0_outputs[4509]) | (layer0_outputs[3785]);
    assign layer1_outputs[3846] = 1'b0;
    assign layer1_outputs[3847] = ~((layer0_outputs[4290]) | (layer0_outputs[4563]));
    assign layer1_outputs[3848] = layer0_outputs[1686];
    assign layer1_outputs[3849] = ~(layer0_outputs[2078]) | (layer0_outputs[840]);
    assign layer1_outputs[3850] = layer0_outputs[4999];
    assign layer1_outputs[3851] = 1'b1;
    assign layer1_outputs[3852] = 1'b0;
    assign layer1_outputs[3853] = 1'b0;
    assign layer1_outputs[3854] = layer0_outputs[3924];
    assign layer1_outputs[3855] = ~(layer0_outputs[4684]);
    assign layer1_outputs[3856] = ~(layer0_outputs[2335]);
    assign layer1_outputs[3857] = layer0_outputs[3565];
    assign layer1_outputs[3858] = (layer0_outputs[4050]) & ~(layer0_outputs[3047]);
    assign layer1_outputs[3859] = (layer0_outputs[2748]) & (layer0_outputs[471]);
    assign layer1_outputs[3860] = layer0_outputs[954];
    assign layer1_outputs[3861] = layer0_outputs[3139];
    assign layer1_outputs[3862] = layer0_outputs[1618];
    assign layer1_outputs[3863] = 1'b1;
    assign layer1_outputs[3864] = (layer0_outputs[2088]) & (layer0_outputs[4970]);
    assign layer1_outputs[3865] = (layer0_outputs[1803]) & (layer0_outputs[138]);
    assign layer1_outputs[3866] = ~((layer0_outputs[2434]) | (layer0_outputs[3304]));
    assign layer1_outputs[3867] = 1'b0;
    assign layer1_outputs[3868] = ~(layer0_outputs[2828]);
    assign layer1_outputs[3869] = (layer0_outputs[3269]) | (layer0_outputs[1006]);
    assign layer1_outputs[3870] = (layer0_outputs[3995]) | (layer0_outputs[3284]);
    assign layer1_outputs[3871] = 1'b1;
    assign layer1_outputs[3872] = layer0_outputs[4034];
    assign layer1_outputs[3873] = ~((layer0_outputs[1056]) & (layer0_outputs[2448]));
    assign layer1_outputs[3874] = (layer0_outputs[3755]) | (layer0_outputs[2357]);
    assign layer1_outputs[3875] = (layer0_outputs[3841]) & ~(layer0_outputs[2322]);
    assign layer1_outputs[3876] = 1'b1;
    assign layer1_outputs[3877] = (layer0_outputs[369]) & (layer0_outputs[1731]);
    assign layer1_outputs[3878] = ~(layer0_outputs[1225]) | (layer0_outputs[405]);
    assign layer1_outputs[3879] = (layer0_outputs[4571]) & (layer0_outputs[2214]);
    assign layer1_outputs[3880] = ~((layer0_outputs[4157]) | (layer0_outputs[3959]));
    assign layer1_outputs[3881] = ~(layer0_outputs[3122]) | (layer0_outputs[1261]);
    assign layer1_outputs[3882] = ~((layer0_outputs[104]) & (layer0_outputs[4481]));
    assign layer1_outputs[3883] = layer0_outputs[4753];
    assign layer1_outputs[3884] = 1'b0;
    assign layer1_outputs[3885] = (layer0_outputs[2113]) | (layer0_outputs[2470]);
    assign layer1_outputs[3886] = 1'b0;
    assign layer1_outputs[3887] = ~((layer0_outputs[4346]) & (layer0_outputs[1913]));
    assign layer1_outputs[3888] = layer0_outputs[4334];
    assign layer1_outputs[3889] = (layer0_outputs[3531]) & ~(layer0_outputs[23]);
    assign layer1_outputs[3890] = (layer0_outputs[4031]) & ~(layer0_outputs[1518]);
    assign layer1_outputs[3891] = ~(layer0_outputs[1028]);
    assign layer1_outputs[3892] = ~((layer0_outputs[3493]) | (layer0_outputs[116]));
    assign layer1_outputs[3893] = layer0_outputs[4960];
    assign layer1_outputs[3894] = ~(layer0_outputs[4421]);
    assign layer1_outputs[3895] = (layer0_outputs[3226]) ^ (layer0_outputs[5047]);
    assign layer1_outputs[3896] = layer0_outputs[3727];
    assign layer1_outputs[3897] = ~(layer0_outputs[4953]);
    assign layer1_outputs[3898] = (layer0_outputs[361]) & ~(layer0_outputs[4143]);
    assign layer1_outputs[3899] = layer0_outputs[543];
    assign layer1_outputs[3900] = ~(layer0_outputs[4350]);
    assign layer1_outputs[3901] = (layer0_outputs[3292]) & ~(layer0_outputs[3971]);
    assign layer1_outputs[3902] = ~((layer0_outputs[4727]) | (layer0_outputs[1843]));
    assign layer1_outputs[3903] = ~(layer0_outputs[2111]);
    assign layer1_outputs[3904] = ~((layer0_outputs[2939]) & (layer0_outputs[3347]));
    assign layer1_outputs[3905] = ~(layer0_outputs[68]) | (layer0_outputs[1920]);
    assign layer1_outputs[3906] = (layer0_outputs[4657]) ^ (layer0_outputs[663]);
    assign layer1_outputs[3907] = 1'b1;
    assign layer1_outputs[3908] = ~(layer0_outputs[4440]);
    assign layer1_outputs[3909] = ~(layer0_outputs[2754]) | (layer0_outputs[1743]);
    assign layer1_outputs[3910] = 1'b1;
    assign layer1_outputs[3911] = (layer0_outputs[32]) | (layer0_outputs[54]);
    assign layer1_outputs[3912] = 1'b1;
    assign layer1_outputs[3913] = ~(layer0_outputs[3892]);
    assign layer1_outputs[3914] = (layer0_outputs[3471]) | (layer0_outputs[2446]);
    assign layer1_outputs[3915] = ~((layer0_outputs[4232]) & (layer0_outputs[2472]));
    assign layer1_outputs[3916] = (layer0_outputs[3143]) | (layer0_outputs[3980]);
    assign layer1_outputs[3917] = layer0_outputs[2022];
    assign layer1_outputs[3918] = ~(layer0_outputs[4605]) | (layer0_outputs[3480]);
    assign layer1_outputs[3919] = ~(layer0_outputs[680]) | (layer0_outputs[2514]);
    assign layer1_outputs[3920] = ~((layer0_outputs[2301]) & (layer0_outputs[2077]));
    assign layer1_outputs[3921] = ~(layer0_outputs[172]);
    assign layer1_outputs[3922] = (layer0_outputs[3124]) & ~(layer0_outputs[4226]);
    assign layer1_outputs[3923] = ~((layer0_outputs[4476]) | (layer0_outputs[4856]));
    assign layer1_outputs[3924] = (layer0_outputs[3024]) ^ (layer0_outputs[4172]);
    assign layer1_outputs[3925] = (layer0_outputs[4321]) & ~(layer0_outputs[2123]);
    assign layer1_outputs[3926] = ~(layer0_outputs[2233]) | (layer0_outputs[2896]);
    assign layer1_outputs[3927] = ~((layer0_outputs[3639]) | (layer0_outputs[3033]));
    assign layer1_outputs[3928] = ~(layer0_outputs[1367]);
    assign layer1_outputs[3929] = layer0_outputs[1784];
    assign layer1_outputs[3930] = 1'b0;
    assign layer1_outputs[3931] = 1'b0;
    assign layer1_outputs[3932] = ~((layer0_outputs[2429]) | (layer0_outputs[3323]));
    assign layer1_outputs[3933] = 1'b1;
    assign layer1_outputs[3934] = ~((layer0_outputs[4848]) & (layer0_outputs[569]));
    assign layer1_outputs[3935] = ~((layer0_outputs[2130]) | (layer0_outputs[3981]));
    assign layer1_outputs[3936] = ~(layer0_outputs[576]) | (layer0_outputs[4497]);
    assign layer1_outputs[3937] = ~(layer0_outputs[4337]) | (layer0_outputs[3811]);
    assign layer1_outputs[3938] = layer0_outputs[4183];
    assign layer1_outputs[3939] = (layer0_outputs[2953]) ^ (layer0_outputs[2935]);
    assign layer1_outputs[3940] = (layer0_outputs[4333]) & ~(layer0_outputs[3719]);
    assign layer1_outputs[3941] = (layer0_outputs[2862]) & (layer0_outputs[2038]);
    assign layer1_outputs[3942] = layer0_outputs[127];
    assign layer1_outputs[3943] = ~((layer0_outputs[1439]) | (layer0_outputs[1062]));
    assign layer1_outputs[3944] = ~((layer0_outputs[3049]) & (layer0_outputs[4852]));
    assign layer1_outputs[3945] = ~((layer0_outputs[920]) & (layer0_outputs[3539]));
    assign layer1_outputs[3946] = 1'b0;
    assign layer1_outputs[3947] = layer0_outputs[2616];
    assign layer1_outputs[3948] = ~((layer0_outputs[2978]) & (layer0_outputs[693]));
    assign layer1_outputs[3949] = ~(layer0_outputs[4205]) | (layer0_outputs[360]);
    assign layer1_outputs[3950] = (layer0_outputs[3323]) & (layer0_outputs[1589]);
    assign layer1_outputs[3951] = ~(layer0_outputs[740]);
    assign layer1_outputs[3952] = 1'b0;
    assign layer1_outputs[3953] = (layer0_outputs[1300]) & (layer0_outputs[2663]);
    assign layer1_outputs[3954] = ~(layer0_outputs[2659]);
    assign layer1_outputs[3955] = ~(layer0_outputs[1307]);
    assign layer1_outputs[3956] = (layer0_outputs[2990]) & (layer0_outputs[3305]);
    assign layer1_outputs[3957] = ~((layer0_outputs[832]) & (layer0_outputs[4172]));
    assign layer1_outputs[3958] = 1'b1;
    assign layer1_outputs[3959] = ~((layer0_outputs[1998]) | (layer0_outputs[1128]));
    assign layer1_outputs[3960] = (layer0_outputs[1538]) & ~(layer0_outputs[1659]);
    assign layer1_outputs[3961] = ~((layer0_outputs[2170]) & (layer0_outputs[3559]));
    assign layer1_outputs[3962] = (layer0_outputs[2211]) & ~(layer0_outputs[4816]);
    assign layer1_outputs[3963] = 1'b1;
    assign layer1_outputs[3964] = ~((layer0_outputs[2421]) ^ (layer0_outputs[3504]));
    assign layer1_outputs[3965] = ~((layer0_outputs[3651]) ^ (layer0_outputs[3197]));
    assign layer1_outputs[3966] = ~(layer0_outputs[966]);
    assign layer1_outputs[3967] = ~(layer0_outputs[4995]);
    assign layer1_outputs[3968] = (layer0_outputs[3132]) & ~(layer0_outputs[4673]);
    assign layer1_outputs[3969] = ~(layer0_outputs[3551]);
    assign layer1_outputs[3970] = ~((layer0_outputs[3181]) | (layer0_outputs[721]));
    assign layer1_outputs[3971] = (layer0_outputs[3452]) & ~(layer0_outputs[799]);
    assign layer1_outputs[3972] = ~(layer0_outputs[613]);
    assign layer1_outputs[3973] = ~(layer0_outputs[2112]);
    assign layer1_outputs[3974] = (layer0_outputs[2098]) & ~(layer0_outputs[2637]);
    assign layer1_outputs[3975] = 1'b0;
    assign layer1_outputs[3976] = ~((layer0_outputs[1627]) | (layer0_outputs[3140]));
    assign layer1_outputs[3977] = ~(layer0_outputs[1906]);
    assign layer1_outputs[3978] = ~(layer0_outputs[2883]);
    assign layer1_outputs[3979] = ~(layer0_outputs[1775]) | (layer0_outputs[1018]);
    assign layer1_outputs[3980] = (layer0_outputs[4991]) | (layer0_outputs[3705]);
    assign layer1_outputs[3981] = 1'b0;
    assign layer1_outputs[3982] = ~(layer0_outputs[5065]) | (layer0_outputs[2869]);
    assign layer1_outputs[3983] = (layer0_outputs[4744]) & ~(layer0_outputs[4426]);
    assign layer1_outputs[3984] = (layer0_outputs[1383]) & ~(layer0_outputs[2700]);
    assign layer1_outputs[3985] = (layer0_outputs[2864]) & (layer0_outputs[4709]);
    assign layer1_outputs[3986] = ~(layer0_outputs[2605]) | (layer0_outputs[4450]);
    assign layer1_outputs[3987] = (layer0_outputs[835]) & ~(layer0_outputs[3762]);
    assign layer1_outputs[3988] = ~(layer0_outputs[400]);
    assign layer1_outputs[3989] = ~((layer0_outputs[1748]) & (layer0_outputs[1594]));
    assign layer1_outputs[3990] = (layer0_outputs[5059]) & ~(layer0_outputs[3607]);
    assign layer1_outputs[3991] = ~(layer0_outputs[3066]) | (layer0_outputs[2761]);
    assign layer1_outputs[3992] = (layer0_outputs[76]) & ~(layer0_outputs[4782]);
    assign layer1_outputs[3993] = layer0_outputs[3791];
    assign layer1_outputs[3994] = layer0_outputs[218];
    assign layer1_outputs[3995] = ~(layer0_outputs[60]) | (layer0_outputs[3620]);
    assign layer1_outputs[3996] = (layer0_outputs[788]) | (layer0_outputs[3317]);
    assign layer1_outputs[3997] = (layer0_outputs[547]) & ~(layer0_outputs[2019]);
    assign layer1_outputs[3998] = ~(layer0_outputs[438]) | (layer0_outputs[4549]);
    assign layer1_outputs[3999] = ~(layer0_outputs[4553]) | (layer0_outputs[1987]);
    assign layer1_outputs[4000] = (layer0_outputs[935]) & ~(layer0_outputs[286]);
    assign layer1_outputs[4001] = ~((layer0_outputs[935]) ^ (layer0_outputs[481]));
    assign layer1_outputs[4002] = (layer0_outputs[2242]) & ~(layer0_outputs[1895]);
    assign layer1_outputs[4003] = layer0_outputs[4149];
    assign layer1_outputs[4004] = layer0_outputs[3187];
    assign layer1_outputs[4005] = (layer0_outputs[4400]) & ~(layer0_outputs[956]);
    assign layer1_outputs[4006] = (layer0_outputs[1599]) & ~(layer0_outputs[2339]);
    assign layer1_outputs[4007] = ~(layer0_outputs[486]) | (layer0_outputs[4154]);
    assign layer1_outputs[4008] = (layer0_outputs[2786]) & ~(layer0_outputs[2327]);
    assign layer1_outputs[4009] = 1'b0;
    assign layer1_outputs[4010] = ~((layer0_outputs[4685]) & (layer0_outputs[2303]));
    assign layer1_outputs[4011] = 1'b0;
    assign layer1_outputs[4012] = ~(layer0_outputs[1288]) | (layer0_outputs[4576]);
    assign layer1_outputs[4013] = ~(layer0_outputs[4297]) | (layer0_outputs[3136]);
    assign layer1_outputs[4014] = (layer0_outputs[4842]) ^ (layer0_outputs[2112]);
    assign layer1_outputs[4015] = ~((layer0_outputs[3640]) & (layer0_outputs[2505]));
    assign layer1_outputs[4016] = 1'b0;
    assign layer1_outputs[4017] = ~((layer0_outputs[780]) | (layer0_outputs[3567]));
    assign layer1_outputs[4018] = ~((layer0_outputs[501]) & (layer0_outputs[1666]));
    assign layer1_outputs[4019] = (layer0_outputs[3331]) & ~(layer0_outputs[4170]);
    assign layer1_outputs[4020] = (layer0_outputs[4014]) | (layer0_outputs[4468]);
    assign layer1_outputs[4021] = ~(layer0_outputs[3535]);
    assign layer1_outputs[4022] = (layer0_outputs[1250]) & ~(layer0_outputs[2363]);
    assign layer1_outputs[4023] = (layer0_outputs[3143]) & (layer0_outputs[4840]);
    assign layer1_outputs[4024] = (layer0_outputs[5075]) | (layer0_outputs[5113]);
    assign layer1_outputs[4025] = 1'b1;
    assign layer1_outputs[4026] = ~(layer0_outputs[3222]);
    assign layer1_outputs[4027] = ~(layer0_outputs[794]);
    assign layer1_outputs[4028] = (layer0_outputs[4754]) | (layer0_outputs[700]);
    assign layer1_outputs[4029] = ~(layer0_outputs[2608]);
    assign layer1_outputs[4030] = 1'b0;
    assign layer1_outputs[4031] = ~(layer0_outputs[2464]) | (layer0_outputs[2452]);
    assign layer1_outputs[4032] = ~(layer0_outputs[4231]) | (layer0_outputs[4343]);
    assign layer1_outputs[4033] = ~((layer0_outputs[2074]) ^ (layer0_outputs[2679]));
    assign layer1_outputs[4034] = ~((layer0_outputs[4434]) | (layer0_outputs[2074]));
    assign layer1_outputs[4035] = ~((layer0_outputs[2035]) & (layer0_outputs[340]));
    assign layer1_outputs[4036] = ~(layer0_outputs[4486]) | (layer0_outputs[258]);
    assign layer1_outputs[4037] = ~(layer0_outputs[770]);
    assign layer1_outputs[4038] = (layer0_outputs[2021]) & ~(layer0_outputs[1452]);
    assign layer1_outputs[4039] = (layer0_outputs[2243]) | (layer0_outputs[2708]);
    assign layer1_outputs[4040] = 1'b0;
    assign layer1_outputs[4041] = ~(layer0_outputs[2233]) | (layer0_outputs[3746]);
    assign layer1_outputs[4042] = 1'b0;
    assign layer1_outputs[4043] = (layer0_outputs[3280]) & (layer0_outputs[1685]);
    assign layer1_outputs[4044] = 1'b1;
    assign layer1_outputs[4045] = ~((layer0_outputs[762]) | (layer0_outputs[4979]));
    assign layer1_outputs[4046] = 1'b0;
    assign layer1_outputs[4047] = (layer0_outputs[2819]) | (layer0_outputs[206]);
    assign layer1_outputs[4048] = ~((layer0_outputs[4599]) & (layer0_outputs[1971]));
    assign layer1_outputs[4049] = ~(layer0_outputs[3005]);
    assign layer1_outputs[4050] = 1'b0;
    assign layer1_outputs[4051] = 1'b0;
    assign layer1_outputs[4052] = 1'b0;
    assign layer1_outputs[4053] = layer0_outputs[1073];
    assign layer1_outputs[4054] = ~((layer0_outputs[3920]) | (layer0_outputs[1987]));
    assign layer1_outputs[4055] = layer0_outputs[115];
    assign layer1_outputs[4056] = 1'b0;
    assign layer1_outputs[4057] = (layer0_outputs[4526]) & (layer0_outputs[4823]);
    assign layer1_outputs[4058] = ~((layer0_outputs[4020]) & (layer0_outputs[3619]));
    assign layer1_outputs[4059] = ~(layer0_outputs[3478]);
    assign layer1_outputs[4060] = ~((layer0_outputs[4707]) | (layer0_outputs[660]));
    assign layer1_outputs[4061] = ~(layer0_outputs[648]);
    assign layer1_outputs[4062] = ~((layer0_outputs[4076]) | (layer0_outputs[3430]));
    assign layer1_outputs[4063] = (layer0_outputs[678]) & ~(layer0_outputs[2599]);
    assign layer1_outputs[4064] = 1'b1;
    assign layer1_outputs[4065] = (layer0_outputs[3635]) & ~(layer0_outputs[4396]);
    assign layer1_outputs[4066] = ~(layer0_outputs[2723]);
    assign layer1_outputs[4067] = layer0_outputs[4952];
    assign layer1_outputs[4068] = ~((layer0_outputs[4186]) ^ (layer0_outputs[4309]));
    assign layer1_outputs[4069] = ~((layer0_outputs[3935]) | (layer0_outputs[2075]));
    assign layer1_outputs[4070] = ~(layer0_outputs[1695]) | (layer0_outputs[4308]);
    assign layer1_outputs[4071] = ~(layer0_outputs[4247]);
    assign layer1_outputs[4072] = ~(layer0_outputs[4155]);
    assign layer1_outputs[4073] = (layer0_outputs[4764]) & (layer0_outputs[1838]);
    assign layer1_outputs[4074] = layer0_outputs[4520];
    assign layer1_outputs[4075] = 1'b0;
    assign layer1_outputs[4076] = 1'b0;
    assign layer1_outputs[4077] = (layer0_outputs[3028]) & ~(layer0_outputs[3325]);
    assign layer1_outputs[4078] = 1'b1;
    assign layer1_outputs[4079] = ~(layer0_outputs[3281]);
    assign layer1_outputs[4080] = (layer0_outputs[4372]) & ~(layer0_outputs[1857]);
    assign layer1_outputs[4081] = (layer0_outputs[4200]) & (layer0_outputs[3561]);
    assign layer1_outputs[4082] = (layer0_outputs[4775]) & ~(layer0_outputs[4730]);
    assign layer1_outputs[4083] = layer0_outputs[4412];
    assign layer1_outputs[4084] = 1'b1;
    assign layer1_outputs[4085] = 1'b1;
    assign layer1_outputs[4086] = ~((layer0_outputs[4153]) | (layer0_outputs[1789]));
    assign layer1_outputs[4087] = ~(layer0_outputs[1934]);
    assign layer1_outputs[4088] = (layer0_outputs[1872]) & ~(layer0_outputs[2842]);
    assign layer1_outputs[4089] = (layer0_outputs[2419]) & ~(layer0_outputs[1620]);
    assign layer1_outputs[4090] = 1'b1;
    assign layer1_outputs[4091] = ~((layer0_outputs[1012]) | (layer0_outputs[977]));
    assign layer1_outputs[4092] = 1'b1;
    assign layer1_outputs[4093] = ~(layer0_outputs[4520]);
    assign layer1_outputs[4094] = (layer0_outputs[1277]) & ~(layer0_outputs[882]);
    assign layer1_outputs[4095] = ~((layer0_outputs[1575]) | (layer0_outputs[1770]));
    assign layer1_outputs[4096] = (layer0_outputs[3933]) ^ (layer0_outputs[2108]);
    assign layer1_outputs[4097] = ~(layer0_outputs[2443]) | (layer0_outputs[441]);
    assign layer1_outputs[4098] = ~(layer0_outputs[379]) | (layer0_outputs[2171]);
    assign layer1_outputs[4099] = ~(layer0_outputs[1013]);
    assign layer1_outputs[4100] = 1'b0;
    assign layer1_outputs[4101] = ~((layer0_outputs[3838]) & (layer0_outputs[1119]));
    assign layer1_outputs[4102] = layer0_outputs[4501];
    assign layer1_outputs[4103] = ~((layer0_outputs[4567]) ^ (layer0_outputs[2725]));
    assign layer1_outputs[4104] = (layer0_outputs[2444]) & (layer0_outputs[4947]);
    assign layer1_outputs[4105] = 1'b0;
    assign layer1_outputs[4106] = (layer0_outputs[2816]) ^ (layer0_outputs[2309]);
    assign layer1_outputs[4107] = ~(layer0_outputs[1132]) | (layer0_outputs[50]);
    assign layer1_outputs[4108] = ~(layer0_outputs[3955]) | (layer0_outputs[4784]);
    assign layer1_outputs[4109] = layer0_outputs[2057];
    assign layer1_outputs[4110] = (layer0_outputs[4642]) & ~(layer0_outputs[1610]);
    assign layer1_outputs[4111] = (layer0_outputs[5110]) ^ (layer0_outputs[2892]);
    assign layer1_outputs[4112] = layer0_outputs[3584];
    assign layer1_outputs[4113] = layer0_outputs[4969];
    assign layer1_outputs[4114] = ~(layer0_outputs[1977]) | (layer0_outputs[3037]);
    assign layer1_outputs[4115] = 1'b1;
    assign layer1_outputs[4116] = 1'b0;
    assign layer1_outputs[4117] = (layer0_outputs[4441]) & (layer0_outputs[2646]);
    assign layer1_outputs[4118] = (layer0_outputs[1961]) & ~(layer0_outputs[4300]);
    assign layer1_outputs[4119] = ~(layer0_outputs[2855]);
    assign layer1_outputs[4120] = ~(layer0_outputs[2029]) | (layer0_outputs[3621]);
    assign layer1_outputs[4121] = ~(layer0_outputs[2628]);
    assign layer1_outputs[4122] = 1'b0;
    assign layer1_outputs[4123] = layer0_outputs[2868];
    assign layer1_outputs[4124] = 1'b0;
    assign layer1_outputs[4125] = 1'b0;
    assign layer1_outputs[4126] = (layer0_outputs[2097]) & ~(layer0_outputs[3777]);
    assign layer1_outputs[4127] = 1'b0;
    assign layer1_outputs[4128] = ~((layer0_outputs[5032]) | (layer0_outputs[2341]));
    assign layer1_outputs[4129] = ~((layer0_outputs[650]) & (layer0_outputs[1332]));
    assign layer1_outputs[4130] = ~((layer0_outputs[1924]) & (layer0_outputs[3664]));
    assign layer1_outputs[4131] = 1'b0;
    assign layer1_outputs[4132] = layer0_outputs[3652];
    assign layer1_outputs[4133] = ~(layer0_outputs[3519]);
    assign layer1_outputs[4134] = ~((layer0_outputs[4683]) | (layer0_outputs[3340]));
    assign layer1_outputs[4135] = ~(layer0_outputs[4607]) | (layer0_outputs[4385]);
    assign layer1_outputs[4136] = 1'b0;
    assign layer1_outputs[4137] = (layer0_outputs[2886]) & ~(layer0_outputs[404]);
    assign layer1_outputs[4138] = ~((layer0_outputs[3866]) | (layer0_outputs[1285]));
    assign layer1_outputs[4139] = layer0_outputs[2333];
    assign layer1_outputs[4140] = layer0_outputs[1317];
    assign layer1_outputs[4141] = ~(layer0_outputs[589]);
    assign layer1_outputs[4142] = layer0_outputs[1383];
    assign layer1_outputs[4143] = (layer0_outputs[1682]) & (layer0_outputs[2435]);
    assign layer1_outputs[4144] = 1'b1;
    assign layer1_outputs[4145] = ~(layer0_outputs[3072]);
    assign layer1_outputs[4146] = ~(layer0_outputs[1166]);
    assign layer1_outputs[4147] = ~((layer0_outputs[3945]) | (layer0_outputs[677]));
    assign layer1_outputs[4148] = ~(layer0_outputs[2521]);
    assign layer1_outputs[4149] = ~((layer0_outputs[1764]) & (layer0_outputs[5108]));
    assign layer1_outputs[4150] = ~((layer0_outputs[166]) & (layer0_outputs[1859]));
    assign layer1_outputs[4151] = (layer0_outputs[990]) ^ (layer0_outputs[1893]);
    assign layer1_outputs[4152] = (layer0_outputs[219]) & ~(layer0_outputs[2977]);
    assign layer1_outputs[4153] = (layer0_outputs[3851]) & ~(layer0_outputs[4558]);
    assign layer1_outputs[4154] = ~(layer0_outputs[2800]) | (layer0_outputs[1034]);
    assign layer1_outputs[4155] = layer0_outputs[809];
    assign layer1_outputs[4156] = ~((layer0_outputs[4574]) & (layer0_outputs[4484]));
    assign layer1_outputs[4157] = layer0_outputs[2149];
    assign layer1_outputs[4158] = 1'b1;
    assign layer1_outputs[4159] = ~((layer0_outputs[1882]) & (layer0_outputs[2405]));
    assign layer1_outputs[4160] = (layer0_outputs[994]) & ~(layer0_outputs[2002]);
    assign layer1_outputs[4161] = ~(layer0_outputs[607]);
    assign layer1_outputs[4162] = ~(layer0_outputs[4736]) | (layer0_outputs[2586]);
    assign layer1_outputs[4163] = layer0_outputs[2188];
    assign layer1_outputs[4164] = 1'b0;
    assign layer1_outputs[4165] = 1'b0;
    assign layer1_outputs[4166] = ~(layer0_outputs[3675]) | (layer0_outputs[4638]);
    assign layer1_outputs[4167] = ~(layer0_outputs[4755]) | (layer0_outputs[410]);
    assign layer1_outputs[4168] = layer0_outputs[2033];
    assign layer1_outputs[4169] = ~(layer0_outputs[1325]) | (layer0_outputs[4597]);
    assign layer1_outputs[4170] = layer0_outputs[4061];
    assign layer1_outputs[4171] = layer0_outputs[3256];
    assign layer1_outputs[4172] = (layer0_outputs[1044]) & ~(layer0_outputs[3826]);
    assign layer1_outputs[4173] = (layer0_outputs[84]) & ~(layer0_outputs[4434]);
    assign layer1_outputs[4174] = layer0_outputs[3457];
    assign layer1_outputs[4175] = layer0_outputs[1593];
    assign layer1_outputs[4176] = layer0_outputs[2060];
    assign layer1_outputs[4177] = 1'b0;
    assign layer1_outputs[4178] = ~((layer0_outputs[4442]) & (layer0_outputs[4758]));
    assign layer1_outputs[4179] = (layer0_outputs[3790]) & ~(layer0_outputs[1391]);
    assign layer1_outputs[4180] = (layer0_outputs[571]) & (layer0_outputs[3749]);
    assign layer1_outputs[4181] = (layer0_outputs[1027]) & ~(layer0_outputs[1068]);
    assign layer1_outputs[4182] = layer0_outputs[2127];
    assign layer1_outputs[4183] = ~(layer0_outputs[2684]) | (layer0_outputs[4330]);
    assign layer1_outputs[4184] = ~(layer0_outputs[4855]) | (layer0_outputs[915]);
    assign layer1_outputs[4185] = 1'b1;
    assign layer1_outputs[4186] = (layer0_outputs[75]) ^ (layer0_outputs[2039]);
    assign layer1_outputs[4187] = (layer0_outputs[4966]) & (layer0_outputs[994]);
    assign layer1_outputs[4188] = (layer0_outputs[4694]) & ~(layer0_outputs[5012]);
    assign layer1_outputs[4189] = 1'b0;
    assign layer1_outputs[4190] = ~(layer0_outputs[2252]) | (layer0_outputs[4899]);
    assign layer1_outputs[4191] = 1'b1;
    assign layer1_outputs[4192] = ~(layer0_outputs[1718]);
    assign layer1_outputs[4193] = ~((layer0_outputs[1754]) & (layer0_outputs[4555]));
    assign layer1_outputs[4194] = layer0_outputs[2473];
    assign layer1_outputs[4195] = ~(layer0_outputs[3747]);
    assign layer1_outputs[4196] = (layer0_outputs[3283]) | (layer0_outputs[469]);
    assign layer1_outputs[4197] = ~((layer0_outputs[1621]) | (layer0_outputs[1961]));
    assign layer1_outputs[4198] = ~(layer0_outputs[4626]) | (layer0_outputs[653]);
    assign layer1_outputs[4199] = layer0_outputs[4765];
    assign layer1_outputs[4200] = ~(layer0_outputs[1663]);
    assign layer1_outputs[4201] = ~((layer0_outputs[2377]) ^ (layer0_outputs[4712]));
    assign layer1_outputs[4202] = (layer0_outputs[4457]) & (layer0_outputs[2818]);
    assign layer1_outputs[4203] = (layer0_outputs[3191]) | (layer0_outputs[2844]);
    assign layer1_outputs[4204] = (layer0_outputs[4159]) & ~(layer0_outputs[947]);
    assign layer1_outputs[4205] = 1'b1;
    assign layer1_outputs[4206] = ~(layer0_outputs[2678]);
    assign layer1_outputs[4207] = layer0_outputs[4313];
    assign layer1_outputs[4208] = (layer0_outputs[4609]) & (layer0_outputs[146]);
    assign layer1_outputs[4209] = ~((layer0_outputs[3871]) | (layer0_outputs[4659]));
    assign layer1_outputs[4210] = 1'b0;
    assign layer1_outputs[4211] = ~((layer0_outputs[2913]) ^ (layer0_outputs[2159]));
    assign layer1_outputs[4212] = (layer0_outputs[4907]) & ~(layer0_outputs[4332]);
    assign layer1_outputs[4213] = (layer0_outputs[3321]) & ~(layer0_outputs[3032]);
    assign layer1_outputs[4214] = (layer0_outputs[4549]) & ~(layer0_outputs[1837]);
    assign layer1_outputs[4215] = layer0_outputs[3688];
    assign layer1_outputs[4216] = ~((layer0_outputs[3694]) ^ (layer0_outputs[2422]));
    assign layer1_outputs[4217] = ~(layer0_outputs[3992]) | (layer0_outputs[324]);
    assign layer1_outputs[4218] = ~((layer0_outputs[3670]) & (layer0_outputs[744]));
    assign layer1_outputs[4219] = (layer0_outputs[285]) ^ (layer0_outputs[1671]);
    assign layer1_outputs[4220] = ~(layer0_outputs[467]);
    assign layer1_outputs[4221] = ~(layer0_outputs[4755]) | (layer0_outputs[1530]);
    assign layer1_outputs[4222] = (layer0_outputs[764]) & (layer0_outputs[4804]);
    assign layer1_outputs[4223] = 1'b1;
    assign layer1_outputs[4224] = ~(layer0_outputs[3348]) | (layer0_outputs[791]);
    assign layer1_outputs[4225] = layer0_outputs[3082];
    assign layer1_outputs[4226] = layer0_outputs[4976];
    assign layer1_outputs[4227] = (layer0_outputs[285]) & ~(layer0_outputs[4680]);
    assign layer1_outputs[4228] = (layer0_outputs[989]) & ~(layer0_outputs[2050]);
    assign layer1_outputs[4229] = ~(layer0_outputs[2133]);
    assign layer1_outputs[4230] = ~((layer0_outputs[4968]) | (layer0_outputs[3213]));
    assign layer1_outputs[4231] = ~(layer0_outputs[5041]);
    assign layer1_outputs[4232] = ~(layer0_outputs[3697]);
    assign layer1_outputs[4233] = (layer0_outputs[2498]) & (layer0_outputs[2330]);
    assign layer1_outputs[4234] = (layer0_outputs[4114]) & ~(layer0_outputs[4890]);
    assign layer1_outputs[4235] = ~(layer0_outputs[2772]);
    assign layer1_outputs[4236] = ~(layer0_outputs[4278]);
    assign layer1_outputs[4237] = ~(layer0_outputs[2277]) | (layer0_outputs[852]);
    assign layer1_outputs[4238] = ~(layer0_outputs[795]);
    assign layer1_outputs[4239] = layer0_outputs[2319];
    assign layer1_outputs[4240] = 1'b1;
    assign layer1_outputs[4241] = ~(layer0_outputs[2222]) | (layer0_outputs[5061]);
    assign layer1_outputs[4242] = ~(layer0_outputs[5035]);
    assign layer1_outputs[4243] = layer0_outputs[4919];
    assign layer1_outputs[4244] = ~((layer0_outputs[1403]) ^ (layer0_outputs[2511]));
    assign layer1_outputs[4245] = ~(layer0_outputs[3848]);
    assign layer1_outputs[4246] = (layer0_outputs[2380]) & ~(layer0_outputs[627]);
    assign layer1_outputs[4247] = ~(layer0_outputs[668]);
    assign layer1_outputs[4248] = (layer0_outputs[636]) & ~(layer0_outputs[3509]);
    assign layer1_outputs[4249] = (layer0_outputs[3862]) | (layer0_outputs[3309]);
    assign layer1_outputs[4250] = ~(layer0_outputs[1265]) | (layer0_outputs[2859]);
    assign layer1_outputs[4251] = layer0_outputs[2820];
    assign layer1_outputs[4252] = ~(layer0_outputs[1825]) | (layer0_outputs[344]);
    assign layer1_outputs[4253] = layer0_outputs[1851];
    assign layer1_outputs[4254] = ~(layer0_outputs[2792]);
    assign layer1_outputs[4255] = 1'b1;
    assign layer1_outputs[4256] = ~(layer0_outputs[3997]) | (layer0_outputs[4717]);
    assign layer1_outputs[4257] = (layer0_outputs[1520]) & ~(layer0_outputs[3585]);
    assign layer1_outputs[4258] = (layer0_outputs[754]) | (layer0_outputs[3085]);
    assign layer1_outputs[4259] = ~((layer0_outputs[2200]) | (layer0_outputs[3844]));
    assign layer1_outputs[4260] = layer0_outputs[1329];
    assign layer1_outputs[4261] = ~(layer0_outputs[779]) | (layer0_outputs[3892]);
    assign layer1_outputs[4262] = (layer0_outputs[4485]) & (layer0_outputs[746]);
    assign layer1_outputs[4263] = (layer0_outputs[2099]) | (layer0_outputs[815]);
    assign layer1_outputs[4264] = 1'b1;
    assign layer1_outputs[4265] = (layer0_outputs[3989]) & (layer0_outputs[444]);
    assign layer1_outputs[4266] = ~(layer0_outputs[4897]);
    assign layer1_outputs[4267] = ~((layer0_outputs[496]) | (layer0_outputs[5117]));
    assign layer1_outputs[4268] = (layer0_outputs[3522]) & ~(layer0_outputs[1229]);
    assign layer1_outputs[4269] = (layer0_outputs[3046]) & ~(layer0_outputs[2989]);
    assign layer1_outputs[4270] = layer0_outputs[2579];
    assign layer1_outputs[4271] = (layer0_outputs[4517]) & (layer0_outputs[334]);
    assign layer1_outputs[4272] = ~(layer0_outputs[1907]);
    assign layer1_outputs[4273] = ~(layer0_outputs[1541]);
    assign layer1_outputs[4274] = layer0_outputs[4317];
    assign layer1_outputs[4275] = 1'b0;
    assign layer1_outputs[4276] = (layer0_outputs[4325]) | (layer0_outputs[4666]);
    assign layer1_outputs[4277] = ~(layer0_outputs[3390]);
    assign layer1_outputs[4278] = ~(layer0_outputs[1501]) | (layer0_outputs[434]);
    assign layer1_outputs[4279] = 1'b0;
    assign layer1_outputs[4280] = layer0_outputs[3345];
    assign layer1_outputs[4281] = layer0_outputs[3919];
    assign layer1_outputs[4282] = ~(layer0_outputs[599]);
    assign layer1_outputs[4283] = 1'b1;
    assign layer1_outputs[4284] = 1'b1;
    assign layer1_outputs[4285] = ~(layer0_outputs[1100]);
    assign layer1_outputs[4286] = 1'b1;
    assign layer1_outputs[4287] = ~((layer0_outputs[2557]) & (layer0_outputs[1021]));
    assign layer1_outputs[4288] = ~((layer0_outputs[1729]) | (layer0_outputs[967]));
    assign layer1_outputs[4289] = ~(layer0_outputs[3548]) | (layer0_outputs[260]);
    assign layer1_outputs[4290] = (layer0_outputs[5079]) & ~(layer0_outputs[315]);
    assign layer1_outputs[4291] = ~(layer0_outputs[1963]);
    assign layer1_outputs[4292] = layer0_outputs[1001];
    assign layer1_outputs[4293] = layer0_outputs[1755];
    assign layer1_outputs[4294] = (layer0_outputs[2030]) | (layer0_outputs[1153]);
    assign layer1_outputs[4295] = layer0_outputs[4655];
    assign layer1_outputs[4296] = layer0_outputs[3420];
    assign layer1_outputs[4297] = (layer0_outputs[1069]) & ~(layer0_outputs[1508]);
    assign layer1_outputs[4298] = ~((layer0_outputs[1816]) ^ (layer0_outputs[2433]));
    assign layer1_outputs[4299] = ~(layer0_outputs[4381]) | (layer0_outputs[2790]);
    assign layer1_outputs[4300] = ~(layer0_outputs[1612]) | (layer0_outputs[4625]);
    assign layer1_outputs[4301] = (layer0_outputs[1813]) & ~(layer0_outputs[3258]);
    assign layer1_outputs[4302] = ~(layer0_outputs[4446]);
    assign layer1_outputs[4303] = ~(layer0_outputs[2436]);
    assign layer1_outputs[4304] = (layer0_outputs[1615]) & (layer0_outputs[3474]);
    assign layer1_outputs[4305] = layer0_outputs[2579];
    assign layer1_outputs[4306] = (layer0_outputs[942]) & ~(layer0_outputs[4818]);
    assign layer1_outputs[4307] = ~(layer0_outputs[3468]) | (layer0_outputs[2120]);
    assign layer1_outputs[4308] = 1'b1;
    assign layer1_outputs[4309] = ~(layer0_outputs[2902]);
    assign layer1_outputs[4310] = (layer0_outputs[3898]) & (layer0_outputs[1876]);
    assign layer1_outputs[4311] = (layer0_outputs[3462]) & (layer0_outputs[1723]);
    assign layer1_outputs[4312] = (layer0_outputs[4642]) & ~(layer0_outputs[474]);
    assign layer1_outputs[4313] = layer0_outputs[782];
    assign layer1_outputs[4314] = (layer0_outputs[4071]) & ~(layer0_outputs[3013]);
    assign layer1_outputs[4315] = layer0_outputs[1417];
    assign layer1_outputs[4316] = ~((layer0_outputs[2482]) ^ (layer0_outputs[3942]));
    assign layer1_outputs[4317] = layer0_outputs[3039];
    assign layer1_outputs[4318] = ~(layer0_outputs[3547]) | (layer0_outputs[1287]);
    assign layer1_outputs[4319] = ~(layer0_outputs[3647]);
    assign layer1_outputs[4320] = ~((layer0_outputs[1194]) & (layer0_outputs[4926]));
    assign layer1_outputs[4321] = ~((layer0_outputs[136]) | (layer0_outputs[41]));
    assign layer1_outputs[4322] = layer0_outputs[1782];
    assign layer1_outputs[4323] = 1'b1;
    assign layer1_outputs[4324] = ~(layer0_outputs[1927]);
    assign layer1_outputs[4325] = ~((layer0_outputs[1265]) | (layer0_outputs[4249]));
    assign layer1_outputs[4326] = ~(layer0_outputs[2728]);
    assign layer1_outputs[4327] = 1'b1;
    assign layer1_outputs[4328] = ~(layer0_outputs[2418]) | (layer0_outputs[5086]);
    assign layer1_outputs[4329] = (layer0_outputs[3661]) | (layer0_outputs[2248]);
    assign layer1_outputs[4330] = ~((layer0_outputs[2556]) & (layer0_outputs[4516]));
    assign layer1_outputs[4331] = ~(layer0_outputs[1509]) | (layer0_outputs[710]);
    assign layer1_outputs[4332] = ~(layer0_outputs[2347]);
    assign layer1_outputs[4333] = 1'b0;
    assign layer1_outputs[4334] = ~(layer0_outputs[2980]) | (layer0_outputs[3484]);
    assign layer1_outputs[4335] = (layer0_outputs[3648]) & ~(layer0_outputs[826]);
    assign layer1_outputs[4336] = (layer0_outputs[2893]) & ~(layer0_outputs[4676]);
    assign layer1_outputs[4337] = 1'b1;
    assign layer1_outputs[4338] = ~(layer0_outputs[3123]) | (layer0_outputs[432]);
    assign layer1_outputs[4339] = layer0_outputs[1088];
    assign layer1_outputs[4340] = layer0_outputs[3747];
    assign layer1_outputs[4341] = ~(layer0_outputs[4904]) | (layer0_outputs[4085]);
    assign layer1_outputs[4342] = ~((layer0_outputs[3641]) & (layer0_outputs[923]));
    assign layer1_outputs[4343] = ~((layer0_outputs[266]) | (layer0_outputs[3366]));
    assign layer1_outputs[4344] = (layer0_outputs[1828]) & (layer0_outputs[449]);
    assign layer1_outputs[4345] = (layer0_outputs[2262]) | (layer0_outputs[3939]);
    assign layer1_outputs[4346] = ~((layer0_outputs[163]) | (layer0_outputs[1392]));
    assign layer1_outputs[4347] = 1'b1;
    assign layer1_outputs[4348] = layer0_outputs[1230];
    assign layer1_outputs[4349] = (layer0_outputs[3055]) | (layer0_outputs[3819]);
    assign layer1_outputs[4350] = ~((layer0_outputs[926]) & (layer0_outputs[48]));
    assign layer1_outputs[4351] = ~((layer0_outputs[4977]) & (layer0_outputs[4533]));
    assign layer1_outputs[4352] = 1'b0;
    assign layer1_outputs[4353] = layer0_outputs[3427];
    assign layer1_outputs[4354] = ~(layer0_outputs[4147]) | (layer0_outputs[1287]);
    assign layer1_outputs[4355] = ~(layer0_outputs[4898]) | (layer0_outputs[4378]);
    assign layer1_outputs[4356] = 1'b1;
    assign layer1_outputs[4357] = (layer0_outputs[988]) & ~(layer0_outputs[810]);
    assign layer1_outputs[4358] = (layer0_outputs[443]) & ~(layer0_outputs[4692]);
    assign layer1_outputs[4359] = ~((layer0_outputs[4290]) | (layer0_outputs[380]));
    assign layer1_outputs[4360] = (layer0_outputs[4215]) & ~(layer0_outputs[2865]);
    assign layer1_outputs[4361] = (layer0_outputs[4195]) & ~(layer0_outputs[987]);
    assign layer1_outputs[4362] = 1'b1;
    assign layer1_outputs[4363] = ~(layer0_outputs[5068]) | (layer0_outputs[4640]);
    assign layer1_outputs[4364] = ~((layer0_outputs[2332]) ^ (layer0_outputs[3512]));
    assign layer1_outputs[4365] = (layer0_outputs[4247]) | (layer0_outputs[3966]);
    assign layer1_outputs[4366] = ~(layer0_outputs[5113]);
    assign layer1_outputs[4367] = 1'b0;
    assign layer1_outputs[4368] = layer0_outputs[1619];
    assign layer1_outputs[4369] = ~(layer0_outputs[2602]);
    assign layer1_outputs[4370] = ~(layer0_outputs[2160]);
    assign layer1_outputs[4371] = ~(layer0_outputs[4950]);
    assign layer1_outputs[4372] = ~(layer0_outputs[3587]) | (layer0_outputs[1603]);
    assign layer1_outputs[4373] = (layer0_outputs[2779]) & (layer0_outputs[43]);
    assign layer1_outputs[4374] = ~(layer0_outputs[371]) | (layer0_outputs[1107]);
    assign layer1_outputs[4375] = layer0_outputs[1535];
    assign layer1_outputs[4376] = (layer0_outputs[4781]) | (layer0_outputs[4529]);
    assign layer1_outputs[4377] = ~((layer0_outputs[3358]) | (layer0_outputs[1670]));
    assign layer1_outputs[4378] = ~(layer0_outputs[5091]) | (layer0_outputs[4286]);
    assign layer1_outputs[4379] = ~(layer0_outputs[4393]);
    assign layer1_outputs[4380] = ~(layer0_outputs[1583]);
    assign layer1_outputs[4381] = ~(layer0_outputs[1342]);
    assign layer1_outputs[4382] = (layer0_outputs[1793]) | (layer0_outputs[4013]);
    assign layer1_outputs[4383] = layer0_outputs[1197];
    assign layer1_outputs[4384] = layer0_outputs[1711];
    assign layer1_outputs[4385] = ~((layer0_outputs[3964]) | (layer0_outputs[1470]));
    assign layer1_outputs[4386] = ~((layer0_outputs[1919]) | (layer0_outputs[1232]));
    assign layer1_outputs[4387] = ~(layer0_outputs[2096]) | (layer0_outputs[1412]);
    assign layer1_outputs[4388] = ~((layer0_outputs[3890]) & (layer0_outputs[3706]));
    assign layer1_outputs[4389] = (layer0_outputs[3088]) & (layer0_outputs[1096]);
    assign layer1_outputs[4390] = layer0_outputs[1555];
    assign layer1_outputs[4391] = layer0_outputs[2314];
    assign layer1_outputs[4392] = layer0_outputs[4697];
    assign layer1_outputs[4393] = ~((layer0_outputs[4789]) | (layer0_outputs[1694]));
    assign layer1_outputs[4394] = (layer0_outputs[626]) | (layer0_outputs[1351]);
    assign layer1_outputs[4395] = layer0_outputs[2819];
    assign layer1_outputs[4396] = ~((layer0_outputs[25]) | (layer0_outputs[1083]));
    assign layer1_outputs[4397] = ~(layer0_outputs[3578]);
    assign layer1_outputs[4398] = ~(layer0_outputs[4368]) | (layer0_outputs[579]);
    assign layer1_outputs[4399] = (layer0_outputs[480]) & ~(layer0_outputs[616]);
    assign layer1_outputs[4400] = layer0_outputs[2891];
    assign layer1_outputs[4401] = 1'b0;
    assign layer1_outputs[4402] = ~(layer0_outputs[2809]) | (layer0_outputs[117]);
    assign layer1_outputs[4403] = (layer0_outputs[358]) & ~(layer0_outputs[207]);
    assign layer1_outputs[4404] = (layer0_outputs[1951]) | (layer0_outputs[482]);
    assign layer1_outputs[4405] = ~((layer0_outputs[1315]) ^ (layer0_outputs[5086]));
    assign layer1_outputs[4406] = 1'b1;
    assign layer1_outputs[4407] = ~(layer0_outputs[161]) | (layer0_outputs[3262]);
    assign layer1_outputs[4408] = ~((layer0_outputs[3537]) ^ (layer0_outputs[3947]));
    assign layer1_outputs[4409] = ~(layer0_outputs[3264]);
    assign layer1_outputs[4410] = (layer0_outputs[1166]) | (layer0_outputs[1999]);
    assign layer1_outputs[4411] = 1'b0;
    assign layer1_outputs[4412] = layer0_outputs[2661];
    assign layer1_outputs[4413] = ~(layer0_outputs[2692]) | (layer0_outputs[3151]);
    assign layer1_outputs[4414] = layer0_outputs[4163];
    assign layer1_outputs[4415] = 1'b0;
    assign layer1_outputs[4416] = 1'b1;
    assign layer1_outputs[4417] = (layer0_outputs[2647]) & (layer0_outputs[1506]);
    assign layer1_outputs[4418] = (layer0_outputs[4467]) & (layer0_outputs[1549]);
    assign layer1_outputs[4419] = 1'b0;
    assign layer1_outputs[4420] = (layer0_outputs[1996]) & ~(layer0_outputs[1968]);
    assign layer1_outputs[4421] = (layer0_outputs[4935]) & ~(layer0_outputs[1327]);
    assign layer1_outputs[4422] = (layer0_outputs[99]) & ~(layer0_outputs[303]);
    assign layer1_outputs[4423] = ~((layer0_outputs[977]) | (layer0_outputs[4934]));
    assign layer1_outputs[4424] = ~(layer0_outputs[1450]);
    assign layer1_outputs[4425] = ~(layer0_outputs[3176]) | (layer0_outputs[1796]);
    assign layer1_outputs[4426] = ~(layer0_outputs[305]) | (layer0_outputs[2830]);
    assign layer1_outputs[4427] = 1'b0;
    assign layer1_outputs[4428] = ~((layer0_outputs[2868]) & (layer0_outputs[742]));
    assign layer1_outputs[4429] = ~(layer0_outputs[3914]);
    assign layer1_outputs[4430] = ~(layer0_outputs[381]);
    assign layer1_outputs[4431] = layer0_outputs[2211];
    assign layer1_outputs[4432] = ~(layer0_outputs[709]);
    assign layer1_outputs[4433] = (layer0_outputs[1953]) ^ (layer0_outputs[2983]);
    assign layer1_outputs[4434] = 1'b1;
    assign layer1_outputs[4435] = ~((layer0_outputs[1940]) & (layer0_outputs[1353]));
    assign layer1_outputs[4436] = (layer0_outputs[1136]) & ~(layer0_outputs[4491]);
    assign layer1_outputs[4437] = (layer0_outputs[445]) & (layer0_outputs[4867]);
    assign layer1_outputs[4438] = (layer0_outputs[2959]) & ~(layer0_outputs[2223]);
    assign layer1_outputs[4439] = layer0_outputs[1409];
    assign layer1_outputs[4440] = (layer0_outputs[2084]) ^ (layer0_outputs[725]);
    assign layer1_outputs[4441] = ~(layer0_outputs[2382]) | (layer0_outputs[3963]);
    assign layer1_outputs[4442] = (layer0_outputs[4334]) | (layer0_outputs[698]);
    assign layer1_outputs[4443] = ~((layer0_outputs[1907]) & (layer0_outputs[2738]));
    assign layer1_outputs[4444] = ~((layer0_outputs[1906]) & (layer0_outputs[1644]));
    assign layer1_outputs[4445] = (layer0_outputs[1973]) & (layer0_outputs[3157]);
    assign layer1_outputs[4446] = 1'b0;
    assign layer1_outputs[4447] = (layer0_outputs[4088]) | (layer0_outputs[4828]);
    assign layer1_outputs[4448] = (layer0_outputs[126]) & (layer0_outputs[2468]);
    assign layer1_outputs[4449] = 1'b1;
    assign layer1_outputs[4450] = ~((layer0_outputs[565]) ^ (layer0_outputs[574]));
    assign layer1_outputs[4451] = (layer0_outputs[4145]) & (layer0_outputs[122]);
    assign layer1_outputs[4452] = (layer0_outputs[81]) ^ (layer0_outputs[2774]);
    assign layer1_outputs[4453] = layer0_outputs[2597];
    assign layer1_outputs[4454] = ~((layer0_outputs[2756]) | (layer0_outputs[4115]));
    assign layer1_outputs[4455] = (layer0_outputs[3079]) & (layer0_outputs[3719]);
    assign layer1_outputs[4456] = layer0_outputs[258];
    assign layer1_outputs[4457] = layer0_outputs[909];
    assign layer1_outputs[4458] = ~(layer0_outputs[4436]) | (layer0_outputs[1915]);
    assign layer1_outputs[4459] = ~((layer0_outputs[1854]) & (layer0_outputs[3511]));
    assign layer1_outputs[4460] = ~(layer0_outputs[4121]);
    assign layer1_outputs[4461] = ~(layer0_outputs[1890]);
    assign layer1_outputs[4462] = layer0_outputs[3349];
    assign layer1_outputs[4463] = (layer0_outputs[875]) & (layer0_outputs[4825]);
    assign layer1_outputs[4464] = (layer0_outputs[5025]) & (layer0_outputs[551]);
    assign layer1_outputs[4465] = (layer0_outputs[1622]) | (layer0_outputs[4179]);
    assign layer1_outputs[4466] = ~((layer0_outputs[1463]) | (layer0_outputs[877]));
    assign layer1_outputs[4467] = (layer0_outputs[3228]) | (layer0_outputs[571]);
    assign layer1_outputs[4468] = ~(layer0_outputs[82]);
    assign layer1_outputs[4469] = ~(layer0_outputs[2525]);
    assign layer1_outputs[4470] = (layer0_outputs[3867]) & ~(layer0_outputs[4592]);
    assign layer1_outputs[4471] = ~(layer0_outputs[4415]) | (layer0_outputs[1991]);
    assign layer1_outputs[4472] = 1'b1;
    assign layer1_outputs[4473] = layer0_outputs[2437];
    assign layer1_outputs[4474] = (layer0_outputs[1464]) & (layer0_outputs[4342]);
    assign layer1_outputs[4475] = layer0_outputs[3805];
    assign layer1_outputs[4476] = ~((layer0_outputs[2284]) & (layer0_outputs[155]));
    assign layer1_outputs[4477] = ~((layer0_outputs[1668]) & (layer0_outputs[4629]));
    assign layer1_outputs[4478] = ~((layer0_outputs[2409]) & (layer0_outputs[4019]));
    assign layer1_outputs[4479] = (layer0_outputs[4657]) & ~(layer0_outputs[1864]);
    assign layer1_outputs[4480] = ~((layer0_outputs[3650]) & (layer0_outputs[187]));
    assign layer1_outputs[4481] = layer0_outputs[4134];
    assign layer1_outputs[4482] = ~(layer0_outputs[2227]) | (layer0_outputs[2602]);
    assign layer1_outputs[4483] = (layer0_outputs[4944]) | (layer0_outputs[5093]);
    assign layer1_outputs[4484] = 1'b0;
    assign layer1_outputs[4485] = ~(layer0_outputs[1808]);
    assign layer1_outputs[4486] = 1'b1;
    assign layer1_outputs[4487] = 1'b0;
    assign layer1_outputs[4488] = ~(layer0_outputs[2526]);
    assign layer1_outputs[4489] = (layer0_outputs[3744]) & ~(layer0_outputs[4636]);
    assign layer1_outputs[4490] = ~(layer0_outputs[1462]) | (layer0_outputs[1091]);
    assign layer1_outputs[4491] = ~(layer0_outputs[3553]);
    assign layer1_outputs[4492] = 1'b0;
    assign layer1_outputs[4493] = ~(layer0_outputs[4647]);
    assign layer1_outputs[4494] = layer0_outputs[131];
    assign layer1_outputs[4495] = ~(layer0_outputs[3176]) | (layer0_outputs[4515]);
    assign layer1_outputs[4496] = ~(layer0_outputs[1918]) | (layer0_outputs[4700]);
    assign layer1_outputs[4497] = ~(layer0_outputs[1581]) | (layer0_outputs[2144]);
    assign layer1_outputs[4498] = 1'b1;
    assign layer1_outputs[4499] = ~(layer0_outputs[3244]);
    assign layer1_outputs[4500] = (layer0_outputs[4894]) & (layer0_outputs[2057]);
    assign layer1_outputs[4501] = (layer0_outputs[139]) & (layer0_outputs[1899]);
    assign layer1_outputs[4502] = ~(layer0_outputs[2885]) | (layer0_outputs[2202]);
    assign layer1_outputs[4503] = (layer0_outputs[3112]) & ~(layer0_outputs[900]);
    assign layer1_outputs[4504] = ~(layer0_outputs[435]) | (layer0_outputs[4773]);
    assign layer1_outputs[4505] = ~((layer0_outputs[3431]) | (layer0_outputs[4301]));
    assign layer1_outputs[4506] = layer0_outputs[3249];
    assign layer1_outputs[4507] = (layer0_outputs[5094]) & ~(layer0_outputs[3817]);
    assign layer1_outputs[4508] = ~((layer0_outputs[911]) & (layer0_outputs[494]));
    assign layer1_outputs[4509] = ~(layer0_outputs[2811]);
    assign layer1_outputs[4510] = (layer0_outputs[4599]) ^ (layer0_outputs[3817]);
    assign layer1_outputs[4511] = 1'b0;
    assign layer1_outputs[4512] = ~((layer0_outputs[230]) & (layer0_outputs[237]));
    assign layer1_outputs[4513] = ~(layer0_outputs[2909]) | (layer0_outputs[729]);
    assign layer1_outputs[4514] = layer0_outputs[1480];
    assign layer1_outputs[4515] = layer0_outputs[2116];
    assign layer1_outputs[4516] = ~((layer0_outputs[4937]) | (layer0_outputs[1499]));
    assign layer1_outputs[4517] = layer0_outputs[581];
    assign layer1_outputs[4518] = (layer0_outputs[50]) & ~(layer0_outputs[2962]);
    assign layer1_outputs[4519] = ~((layer0_outputs[436]) & (layer0_outputs[2459]));
    assign layer1_outputs[4520] = (layer0_outputs[3011]) & ~(layer0_outputs[4094]);
    assign layer1_outputs[4521] = layer0_outputs[2665];
    assign layer1_outputs[4522] = ~(layer0_outputs[3563]) | (layer0_outputs[1130]);
    assign layer1_outputs[4523] = (layer0_outputs[542]) & (layer0_outputs[2210]);
    assign layer1_outputs[4524] = 1'b0;
    assign layer1_outputs[4525] = layer0_outputs[4690];
    assign layer1_outputs[4526] = (layer0_outputs[1190]) & ~(layer0_outputs[4740]);
    assign layer1_outputs[4527] = (layer0_outputs[127]) & ~(layer0_outputs[1700]);
    assign layer1_outputs[4528] = ~(layer0_outputs[2994]);
    assign layer1_outputs[4529] = ~(layer0_outputs[4850]) | (layer0_outputs[5119]);
    assign layer1_outputs[4530] = (layer0_outputs[2931]) & ~(layer0_outputs[3701]);
    assign layer1_outputs[4531] = ~(layer0_outputs[659]);
    assign layer1_outputs[4532] = layer0_outputs[2731];
    assign layer1_outputs[4533] = ~(layer0_outputs[2878]);
    assign layer1_outputs[4534] = ~(layer0_outputs[2940]) | (layer0_outputs[3125]);
    assign layer1_outputs[4535] = layer0_outputs[1502];
    assign layer1_outputs[4536] = ~((layer0_outputs[4200]) & (layer0_outputs[4837]));
    assign layer1_outputs[4537] = ~(layer0_outputs[2781]);
    assign layer1_outputs[4538] = (layer0_outputs[3979]) | (layer0_outputs[4401]);
    assign layer1_outputs[4539] = 1'b0;
    assign layer1_outputs[4540] = ~(layer0_outputs[1172]) | (layer0_outputs[2514]);
    assign layer1_outputs[4541] = (layer0_outputs[2427]) | (layer0_outputs[4811]);
    assign layer1_outputs[4542] = (layer0_outputs[2866]) & ~(layer0_outputs[1675]);
    assign layer1_outputs[4543] = ~(layer0_outputs[1207]);
    assign layer1_outputs[4544] = ~(layer0_outputs[401]);
    assign layer1_outputs[4545] = layer0_outputs[1512];
    assign layer1_outputs[4546] = ~(layer0_outputs[3152]);
    assign layer1_outputs[4547] = ~((layer0_outputs[130]) ^ (layer0_outputs[1621]));
    assign layer1_outputs[4548] = (layer0_outputs[3047]) | (layer0_outputs[2135]);
    assign layer1_outputs[4549] = 1'b0;
    assign layer1_outputs[4550] = ~(layer0_outputs[2428]);
    assign layer1_outputs[4551] = ~(layer0_outputs[1310]);
    assign layer1_outputs[4552] = ~((layer0_outputs[1633]) | (layer0_outputs[2696]));
    assign layer1_outputs[4553] = ~(layer0_outputs[4654]);
    assign layer1_outputs[4554] = (layer0_outputs[3757]) | (layer0_outputs[1617]);
    assign layer1_outputs[4555] = ~(layer0_outputs[796]) | (layer0_outputs[1826]);
    assign layer1_outputs[4556] = 1'b0;
    assign layer1_outputs[4557] = (layer0_outputs[2402]) | (layer0_outputs[5087]);
    assign layer1_outputs[4558] = layer0_outputs[2338];
    assign layer1_outputs[4559] = ~((layer0_outputs[4357]) & (layer0_outputs[3842]));
    assign layer1_outputs[4560] = ~((layer0_outputs[2063]) & (layer0_outputs[3225]));
    assign layer1_outputs[4561] = layer0_outputs[4639];
    assign layer1_outputs[4562] = ~(layer0_outputs[1964]) | (layer0_outputs[2329]);
    assign layer1_outputs[4563] = 1'b0;
    assign layer1_outputs[4564] = ~(layer0_outputs[170]);
    assign layer1_outputs[4565] = ~((layer0_outputs[3283]) | (layer0_outputs[1001]));
    assign layer1_outputs[4566] = (layer0_outputs[4461]) ^ (layer0_outputs[4472]);
    assign layer1_outputs[4567] = ~(layer0_outputs[4129]);
    assign layer1_outputs[4568] = ~(layer0_outputs[2989]);
    assign layer1_outputs[4569] = 1'b1;
    assign layer1_outputs[4570] = ~(layer0_outputs[3404]);
    assign layer1_outputs[4571] = ~((layer0_outputs[2291]) | (layer0_outputs[1168]));
    assign layer1_outputs[4572] = 1'b1;
    assign layer1_outputs[4573] = 1'b1;
    assign layer1_outputs[4574] = layer0_outputs[1316];
    assign layer1_outputs[4575] = (layer0_outputs[3231]) | (layer0_outputs[3523]);
    assign layer1_outputs[4576] = ~(layer0_outputs[2034]) | (layer0_outputs[119]);
    assign layer1_outputs[4577] = ~(layer0_outputs[1532]) | (layer0_outputs[728]);
    assign layer1_outputs[4578] = ~(layer0_outputs[1526]) | (layer0_outputs[3362]);
    assign layer1_outputs[4579] = ~((layer0_outputs[4306]) | (layer0_outputs[4994]));
    assign layer1_outputs[4580] = layer0_outputs[993];
    assign layer1_outputs[4581] = ~(layer0_outputs[3543]) | (layer0_outputs[110]);
    assign layer1_outputs[4582] = layer0_outputs[4145];
    assign layer1_outputs[4583] = ~(layer0_outputs[4897]) | (layer0_outputs[4342]);
    assign layer1_outputs[4584] = ~(layer0_outputs[414]);
    assign layer1_outputs[4585] = (layer0_outputs[675]) & ~(layer0_outputs[985]);
    assign layer1_outputs[4586] = 1'b1;
    assign layer1_outputs[4587] = (layer0_outputs[4230]) | (layer0_outputs[3454]);
    assign layer1_outputs[4588] = layer0_outputs[366];
    assign layer1_outputs[4589] = (layer0_outputs[91]) & ~(layer0_outputs[3923]);
    assign layer1_outputs[4590] = ~((layer0_outputs[3282]) & (layer0_outputs[332]));
    assign layer1_outputs[4591] = ~((layer0_outputs[3415]) | (layer0_outputs[706]));
    assign layer1_outputs[4592] = ~(layer0_outputs[3588]);
    assign layer1_outputs[4593] = ~((layer0_outputs[5040]) | (layer0_outputs[499]));
    assign layer1_outputs[4594] = ~(layer0_outputs[1029]);
    assign layer1_outputs[4595] = ~(layer0_outputs[950]) | (layer0_outputs[2926]);
    assign layer1_outputs[4596] = ~(layer0_outputs[895]);
    assign layer1_outputs[4597] = ~(layer0_outputs[2184]);
    assign layer1_outputs[4598] = (layer0_outputs[1273]) & ~(layer0_outputs[2621]);
    assign layer1_outputs[4599] = ~(layer0_outputs[4747]) | (layer0_outputs[124]);
    assign layer1_outputs[4600] = ~(layer0_outputs[1665]) | (layer0_outputs[4190]);
    assign layer1_outputs[4601] = ~(layer0_outputs[4705]);
    assign layer1_outputs[4602] = ~(layer0_outputs[4828]) | (layer0_outputs[2723]);
    assign layer1_outputs[4603] = 1'b0;
    assign layer1_outputs[4604] = (layer0_outputs[2046]) & ~(layer0_outputs[3833]);
    assign layer1_outputs[4605] = 1'b1;
    assign layer1_outputs[4606] = ~((layer0_outputs[2320]) ^ (layer0_outputs[196]));
    assign layer1_outputs[4607] = ~(layer0_outputs[2687]) | (layer0_outputs[664]);
    assign layer1_outputs[4608] = ~((layer0_outputs[4139]) & (layer0_outputs[3244]));
    assign layer1_outputs[4609] = (layer0_outputs[4194]) & ~(layer0_outputs[4358]);
    assign layer1_outputs[4610] = ~(layer0_outputs[3371]) | (layer0_outputs[1105]);
    assign layer1_outputs[4611] = ~(layer0_outputs[4835]);
    assign layer1_outputs[4612] = ~(layer0_outputs[3748]) | (layer0_outputs[4359]);
    assign layer1_outputs[4613] = ~(layer0_outputs[3538]);
    assign layer1_outputs[4614] = (layer0_outputs[2080]) | (layer0_outputs[132]);
    assign layer1_outputs[4615] = 1'b1;
    assign layer1_outputs[4616] = (layer0_outputs[762]) & ~(layer0_outputs[3679]);
    assign layer1_outputs[4617] = ~(layer0_outputs[4670]);
    assign layer1_outputs[4618] = ~((layer0_outputs[3814]) | (layer0_outputs[2974]));
    assign layer1_outputs[4619] = ~(layer0_outputs[4275]) | (layer0_outputs[1964]);
    assign layer1_outputs[4620] = 1'b0;
    assign layer1_outputs[4621] = ~((layer0_outputs[806]) ^ (layer0_outputs[2244]));
    assign layer1_outputs[4622] = (layer0_outputs[4305]) & ~(layer0_outputs[4025]);
    assign layer1_outputs[4623] = ~(layer0_outputs[3680]);
    assign layer1_outputs[4624] = 1'b0;
    assign layer1_outputs[4625] = layer0_outputs[1298];
    assign layer1_outputs[4626] = (layer0_outputs[40]) & (layer0_outputs[3816]);
    assign layer1_outputs[4627] = (layer0_outputs[2942]) | (layer0_outputs[2100]);
    assign layer1_outputs[4628] = 1'b0;
    assign layer1_outputs[4629] = (layer0_outputs[4231]) & ~(layer0_outputs[378]);
    assign layer1_outputs[4630] = (layer0_outputs[4915]) & ~(layer0_outputs[3291]);
    assign layer1_outputs[4631] = ~(layer0_outputs[1134]);
    assign layer1_outputs[4632] = layer0_outputs[1589];
    assign layer1_outputs[4633] = layer0_outputs[279];
    assign layer1_outputs[4634] = (layer0_outputs[2231]) | (layer0_outputs[359]);
    assign layer1_outputs[4635] = 1'b0;
    assign layer1_outputs[4636] = 1'b0;
    assign layer1_outputs[4637] = (layer0_outputs[2433]) & ~(layer0_outputs[4366]);
    assign layer1_outputs[4638] = (layer0_outputs[170]) & ~(layer0_outputs[1730]);
    assign layer1_outputs[4639] = (layer0_outputs[1004]) & (layer0_outputs[4665]);
    assign layer1_outputs[4640] = ~((layer0_outputs[1676]) & (layer0_outputs[1329]));
    assign layer1_outputs[4641] = 1'b1;
    assign layer1_outputs[4642] = ~((layer0_outputs[1824]) & (layer0_outputs[1709]));
    assign layer1_outputs[4643] = layer0_outputs[4831];
    assign layer1_outputs[4644] = ~((layer0_outputs[4293]) | (layer0_outputs[350]));
    assign layer1_outputs[4645] = ~(layer0_outputs[1070]);
    assign layer1_outputs[4646] = (layer0_outputs[299]) & ~(layer0_outputs[4095]);
    assign layer1_outputs[4647] = layer0_outputs[3636];
    assign layer1_outputs[4648] = ~(layer0_outputs[2010]);
    assign layer1_outputs[4649] = ~((layer0_outputs[3179]) & (layer0_outputs[3279]));
    assign layer1_outputs[4650] = (layer0_outputs[4808]) & ~(layer0_outputs[3626]);
    assign layer1_outputs[4651] = ~((layer0_outputs[4414]) | (layer0_outputs[1234]));
    assign layer1_outputs[4652] = ~(layer0_outputs[2511]);
    assign layer1_outputs[4653] = ~(layer0_outputs[3101]) | (layer0_outputs[4198]);
    assign layer1_outputs[4654] = ~((layer0_outputs[2272]) & (layer0_outputs[1496]));
    assign layer1_outputs[4655] = ~(layer0_outputs[608]) | (layer0_outputs[3591]);
    assign layer1_outputs[4656] = (layer0_outputs[4767]) | (layer0_outputs[2186]);
    assign layer1_outputs[4657] = layer0_outputs[356];
    assign layer1_outputs[4658] = (layer0_outputs[2427]) | (layer0_outputs[4169]);
    assign layer1_outputs[4659] = (layer0_outputs[463]) | (layer0_outputs[1422]);
    assign layer1_outputs[4660] = ~(layer0_outputs[1298]);
    assign layer1_outputs[4661] = layer0_outputs[3375];
    assign layer1_outputs[4662] = (layer0_outputs[1227]) & (layer0_outputs[2890]);
    assign layer1_outputs[4663] = (layer0_outputs[375]) & (layer0_outputs[2371]);
    assign layer1_outputs[4664] = ~((layer0_outputs[778]) | (layer0_outputs[434]));
    assign layer1_outputs[4665] = (layer0_outputs[2307]) & ~(layer0_outputs[3156]);
    assign layer1_outputs[4666] = ~((layer0_outputs[2274]) ^ (layer0_outputs[3501]));
    assign layer1_outputs[4667] = ~(layer0_outputs[135]) | (layer0_outputs[5082]);
    assign layer1_outputs[4668] = ~((layer0_outputs[1651]) & (layer0_outputs[4712]));
    assign layer1_outputs[4669] = ~((layer0_outputs[1054]) | (layer0_outputs[3523]));
    assign layer1_outputs[4670] = ~((layer0_outputs[1402]) & (layer0_outputs[3853]));
    assign layer1_outputs[4671] = layer0_outputs[915];
    assign layer1_outputs[4672] = ~((layer0_outputs[3355]) | (layer0_outputs[4053]));
    assign layer1_outputs[4673] = (layer0_outputs[1471]) & (layer0_outputs[3721]);
    assign layer1_outputs[4674] = layer0_outputs[661];
    assign layer1_outputs[4675] = ~(layer0_outputs[3298]);
    assign layer1_outputs[4676] = ~(layer0_outputs[2356]);
    assign layer1_outputs[4677] = ~(layer0_outputs[4623]);
    assign layer1_outputs[4678] = ~((layer0_outputs[116]) & (layer0_outputs[2986]));
    assign layer1_outputs[4679] = 1'b0;
    assign layer1_outputs[4680] = (layer0_outputs[2262]) & ~(layer0_outputs[1294]);
    assign layer1_outputs[4681] = layer0_outputs[4401];
    assign layer1_outputs[4682] = (layer0_outputs[3820]) | (layer0_outputs[3382]);
    assign layer1_outputs[4683] = 1'b0;
    assign layer1_outputs[4684] = ~(layer0_outputs[98]);
    assign layer1_outputs[4685] = layer0_outputs[3366];
    assign layer1_outputs[4686] = ~((layer0_outputs[1016]) & (layer0_outputs[4656]));
    assign layer1_outputs[4687] = (layer0_outputs[26]) & ~(layer0_outputs[2128]);
    assign layer1_outputs[4688] = layer0_outputs[952];
    assign layer1_outputs[4689] = ~((layer0_outputs[1597]) & (layer0_outputs[1836]));
    assign layer1_outputs[4690] = (layer0_outputs[5014]) | (layer0_outputs[1856]);
    assign layer1_outputs[4691] = ~(layer0_outputs[3743]);
    assign layer1_outputs[4692] = ~((layer0_outputs[2208]) | (layer0_outputs[1258]));
    assign layer1_outputs[4693] = 1'b0;
    assign layer1_outputs[4694] = (layer0_outputs[4285]) & ~(layer0_outputs[1063]);
    assign layer1_outputs[4695] = ~(layer0_outputs[2215]) | (layer0_outputs[3798]);
    assign layer1_outputs[4696] = 1'b0;
    assign layer1_outputs[4697] = ~(layer0_outputs[598]) | (layer0_outputs[914]);
    assign layer1_outputs[4698] = (layer0_outputs[2406]) & ~(layer0_outputs[717]);
    assign layer1_outputs[4699] = ~((layer0_outputs[4564]) | (layer0_outputs[2376]));
    assign layer1_outputs[4700] = 1'b1;
    assign layer1_outputs[4701] = ~(layer0_outputs[1884]);
    assign layer1_outputs[4702] = 1'b0;
    assign layer1_outputs[4703] = (layer0_outputs[2110]) & (layer0_outputs[4545]);
    assign layer1_outputs[4704] = ~((layer0_outputs[1221]) & (layer0_outputs[1901]));
    assign layer1_outputs[4705] = ~(layer0_outputs[2187]) | (layer0_outputs[2150]);
    assign layer1_outputs[4706] = ~(layer0_outputs[3089]);
    assign layer1_outputs[4707] = ~((layer0_outputs[2728]) & (layer0_outputs[2528]));
    assign layer1_outputs[4708] = ~(layer0_outputs[4814]);
    assign layer1_outputs[4709] = ~((layer0_outputs[3803]) & (layer0_outputs[1866]));
    assign layer1_outputs[4710] = ~(layer0_outputs[3282]) | (layer0_outputs[2562]);
    assign layer1_outputs[4711] = (layer0_outputs[153]) ^ (layer0_outputs[2961]);
    assign layer1_outputs[4712] = (layer0_outputs[21]) & (layer0_outputs[4760]);
    assign layer1_outputs[4713] = (layer0_outputs[3714]) & ~(layer0_outputs[4199]);
    assign layer1_outputs[4714] = (layer0_outputs[2763]) & (layer0_outputs[2467]);
    assign layer1_outputs[4715] = ~(layer0_outputs[2987]) | (layer0_outputs[672]);
    assign layer1_outputs[4716] = 1'b0;
    assign layer1_outputs[4717] = ~(layer0_outputs[3224]) | (layer0_outputs[105]);
    assign layer1_outputs[4718] = 1'b0;
    assign layer1_outputs[4719] = ~(layer0_outputs[1291]);
    assign layer1_outputs[4720] = (layer0_outputs[3433]) & ~(layer0_outputs[3673]);
    assign layer1_outputs[4721] = ~(layer0_outputs[371]) | (layer0_outputs[2101]);
    assign layer1_outputs[4722] = ~(layer0_outputs[2601]) | (layer0_outputs[2548]);
    assign layer1_outputs[4723] = layer0_outputs[4129];
    assign layer1_outputs[4724] = (layer0_outputs[3210]) & ~(layer0_outputs[3514]);
    assign layer1_outputs[4725] = ~((layer0_outputs[4004]) & (layer0_outputs[1485]));
    assign layer1_outputs[4726] = ~(layer0_outputs[2889]) | (layer0_outputs[4960]);
    assign layer1_outputs[4727] = ~(layer0_outputs[3138]);
    assign layer1_outputs[4728] = ~(layer0_outputs[2005]);
    assign layer1_outputs[4729] = (layer0_outputs[310]) & ~(layer0_outputs[4457]);
    assign layer1_outputs[4730] = ~((layer0_outputs[4157]) & (layer0_outputs[3674]));
    assign layer1_outputs[4731] = ~(layer0_outputs[1614]) | (layer0_outputs[1116]);
    assign layer1_outputs[4732] = ~(layer0_outputs[4199]) | (layer0_outputs[3676]);
    assign layer1_outputs[4733] = (layer0_outputs[2775]) | (layer0_outputs[4735]);
    assign layer1_outputs[4734] = (layer0_outputs[3359]) & ~(layer0_outputs[403]);
    assign layer1_outputs[4735] = ~((layer0_outputs[1120]) & (layer0_outputs[1773]));
    assign layer1_outputs[4736] = (layer0_outputs[1387]) | (layer0_outputs[3391]);
    assign layer1_outputs[4737] = (layer0_outputs[3036]) & (layer0_outputs[3314]);
    assign layer1_outputs[4738] = (layer0_outputs[4418]) & ~(layer0_outputs[1998]);
    assign layer1_outputs[4739] = layer0_outputs[1200];
    assign layer1_outputs[4740] = ~((layer0_outputs[4589]) & (layer0_outputs[1301]));
    assign layer1_outputs[4741] = 1'b0;
    assign layer1_outputs[4742] = (layer0_outputs[4667]) & ~(layer0_outputs[1794]);
    assign layer1_outputs[4743] = ~(layer0_outputs[3806]) | (layer0_outputs[416]);
    assign layer1_outputs[4744] = 1'b0;
    assign layer1_outputs[4745] = (layer0_outputs[3737]) & ~(layer0_outputs[2695]);
    assign layer1_outputs[4746] = ~(layer0_outputs[618]);
    assign layer1_outputs[4747] = layer0_outputs[2937];
    assign layer1_outputs[4748] = 1'b1;
    assign layer1_outputs[4749] = layer0_outputs[3313];
    assign layer1_outputs[4750] = 1'b1;
    assign layer1_outputs[4751] = ~(layer0_outputs[2181]);
    assign layer1_outputs[4752] = ~(layer0_outputs[4048]) | (layer0_outputs[1443]);
    assign layer1_outputs[4753] = ~(layer0_outputs[2372]);
    assign layer1_outputs[4754] = (layer0_outputs[3042]) | (layer0_outputs[3836]);
    assign layer1_outputs[4755] = ~(layer0_outputs[4115]);
    assign layer1_outputs[4756] = 1'b1;
    assign layer1_outputs[4757] = (layer0_outputs[4636]) & (layer0_outputs[1186]);
    assign layer1_outputs[4758] = ~((layer0_outputs[413]) & (layer0_outputs[1775]));
    assign layer1_outputs[4759] = ~(layer0_outputs[1612]) | (layer0_outputs[704]);
    assign layer1_outputs[4760] = 1'b1;
    assign layer1_outputs[4761] = layer0_outputs[521];
    assign layer1_outputs[4762] = layer0_outputs[406];
    assign layer1_outputs[4763] = ~(layer0_outputs[123]);
    assign layer1_outputs[4764] = (layer0_outputs[945]) ^ (layer0_outputs[3453]);
    assign layer1_outputs[4765] = ~(layer0_outputs[678]);
    assign layer1_outputs[4766] = ~(layer0_outputs[551]) | (layer0_outputs[2805]);
    assign layer1_outputs[4767] = ~((layer0_outputs[2797]) ^ (layer0_outputs[4080]));
    assign layer1_outputs[4768] = ~(layer0_outputs[4583]) | (layer0_outputs[1606]);
    assign layer1_outputs[4769] = 1'b0;
    assign layer1_outputs[4770] = ~((layer0_outputs[997]) & (layer0_outputs[2081]));
    assign layer1_outputs[4771] = (layer0_outputs[3575]) | (layer0_outputs[4066]);
    assign layer1_outputs[4772] = layer0_outputs[1153];
    assign layer1_outputs[4773] = ~((layer0_outputs[3130]) & (layer0_outputs[1033]));
    assign layer1_outputs[4774] = layer0_outputs[1517];
    assign layer1_outputs[4775] = (layer0_outputs[3640]) & ~(layer0_outputs[5087]);
    assign layer1_outputs[4776] = 1'b0;
    assign layer1_outputs[4777] = 1'b1;
    assign layer1_outputs[4778] = layer0_outputs[1678];
    assign layer1_outputs[4779] = (layer0_outputs[3552]) | (layer0_outputs[4754]);
    assign layer1_outputs[4780] = ~(layer0_outputs[3135]);
    assign layer1_outputs[4781] = (layer0_outputs[4861]) & ~(layer0_outputs[548]);
    assign layer1_outputs[4782] = 1'b0;
    assign layer1_outputs[4783] = layer0_outputs[3463];
    assign layer1_outputs[4784] = (layer0_outputs[4677]) | (layer0_outputs[4403]);
    assign layer1_outputs[4785] = ~(layer0_outputs[1461]);
    assign layer1_outputs[4786] = ~(layer0_outputs[676]);
    assign layer1_outputs[4787] = ~((layer0_outputs[2073]) | (layer0_outputs[1954]));
    assign layer1_outputs[4788] = (layer0_outputs[3000]) | (layer0_outputs[3426]);
    assign layer1_outputs[4789] = layer0_outputs[3498];
    assign layer1_outputs[4790] = ~(layer0_outputs[1374]) | (layer0_outputs[4926]);
    assign layer1_outputs[4791] = (layer0_outputs[645]) & (layer0_outputs[5054]);
    assign layer1_outputs[4792] = 1'b1;
    assign layer1_outputs[4793] = 1'b0;
    assign layer1_outputs[4794] = ~(layer0_outputs[2418]) | (layer0_outputs[4546]);
    assign layer1_outputs[4795] = layer0_outputs[1231];
    assign layer1_outputs[4796] = (layer0_outputs[781]) | (layer0_outputs[1985]);
    assign layer1_outputs[4797] = (layer0_outputs[4186]) & ~(layer0_outputs[1942]);
    assign layer1_outputs[4798] = (layer0_outputs[3566]) & ~(layer0_outputs[2154]);
    assign layer1_outputs[4799] = layer0_outputs[4631];
    assign layer1_outputs[4800] = (layer0_outputs[2344]) & ~(layer0_outputs[4929]);
    assign layer1_outputs[4801] = 1'b1;
    assign layer1_outputs[4802] = ~((layer0_outputs[1441]) | (layer0_outputs[1503]));
    assign layer1_outputs[4803] = ~(layer0_outputs[4369]) | (layer0_outputs[2129]);
    assign layer1_outputs[4804] = ~(layer0_outputs[479]) | (layer0_outputs[2194]);
    assign layer1_outputs[4805] = ~(layer0_outputs[615]);
    assign layer1_outputs[4806] = (layer0_outputs[3911]) & ~(layer0_outputs[3642]);
    assign layer1_outputs[4807] = layer0_outputs[2177];
    assign layer1_outputs[4808] = 1'b0;
    assign layer1_outputs[4809] = layer0_outputs[4471];
    assign layer1_outputs[4810] = ~(layer0_outputs[665]);
    assign layer1_outputs[4811] = 1'b0;
    assign layer1_outputs[4812] = (layer0_outputs[1260]) & (layer0_outputs[2612]);
    assign layer1_outputs[4813] = ~((layer0_outputs[4948]) ^ (layer0_outputs[4543]));
    assign layer1_outputs[4814] = ~(layer0_outputs[3589]) | (layer0_outputs[1580]);
    assign layer1_outputs[4815] = (layer0_outputs[4632]) & ~(layer0_outputs[4072]);
    assign layer1_outputs[4816] = layer0_outputs[3977];
    assign layer1_outputs[4817] = (layer0_outputs[4117]) ^ (layer0_outputs[2835]);
    assign layer1_outputs[4818] = ~((layer0_outputs[437]) & (layer0_outputs[5]));
    assign layer1_outputs[4819] = ~((layer0_outputs[1751]) ^ (layer0_outputs[2201]));
    assign layer1_outputs[4820] = 1'b1;
    assign layer1_outputs[4821] = 1'b1;
    assign layer1_outputs[4822] = (layer0_outputs[3397]) | (layer0_outputs[974]);
    assign layer1_outputs[4823] = 1'b1;
    assign layer1_outputs[4824] = ~(layer0_outputs[241]);
    assign layer1_outputs[4825] = 1'b1;
    assign layer1_outputs[4826] = 1'b0;
    assign layer1_outputs[4827] = 1'b0;
    assign layer1_outputs[4828] = 1'b0;
    assign layer1_outputs[4829] = ~((layer0_outputs[959]) ^ (layer0_outputs[2863]));
    assign layer1_outputs[4830] = ~(layer0_outputs[4203]);
    assign layer1_outputs[4831] = 1'b0;
    assign layer1_outputs[4832] = 1'b1;
    assign layer1_outputs[4833] = ~((layer0_outputs[1305]) & (layer0_outputs[617]));
    assign layer1_outputs[4834] = 1'b0;
    assign layer1_outputs[4835] = 1'b1;
    assign layer1_outputs[4836] = ~(layer0_outputs[4808]) | (layer0_outputs[4309]);
    assign layer1_outputs[4837] = (layer0_outputs[1237]) & ~(layer0_outputs[55]);
    assign layer1_outputs[4838] = layer0_outputs[199];
    assign layer1_outputs[4839] = ~(layer0_outputs[760]);
    assign layer1_outputs[4840] = ~(layer0_outputs[4826]) | (layer0_outputs[939]);
    assign layer1_outputs[4841] = ~(layer0_outputs[3730]);
    assign layer1_outputs[4842] = ~(layer0_outputs[4303]) | (layer0_outputs[2699]);
    assign layer1_outputs[4843] = layer0_outputs[24];
    assign layer1_outputs[4844] = 1'b1;
    assign layer1_outputs[4845] = ~((layer0_outputs[785]) ^ (layer0_outputs[2605]));
    assign layer1_outputs[4846] = 1'b0;
    assign layer1_outputs[4847] = (layer0_outputs[1736]) & ~(layer0_outputs[1446]);
    assign layer1_outputs[4848] = ~(layer0_outputs[2100]) | (layer0_outputs[2894]);
    assign layer1_outputs[4849] = (layer0_outputs[4026]) & ~(layer0_outputs[3578]);
    assign layer1_outputs[4850] = ~((layer0_outputs[483]) & (layer0_outputs[4474]));
    assign layer1_outputs[4851] = ~(layer0_outputs[1086]);
    assign layer1_outputs[4852] = (layer0_outputs[1704]) | (layer0_outputs[4670]);
    assign layer1_outputs[4853] = 1'b1;
    assign layer1_outputs[4854] = 1'b0;
    assign layer1_outputs[4855] = ~(layer0_outputs[4012]) | (layer0_outputs[3041]);
    assign layer1_outputs[4856] = (layer0_outputs[4432]) | (layer0_outputs[2870]);
    assign layer1_outputs[4857] = 1'b0;
    assign layer1_outputs[4858] = ~(layer0_outputs[3389]) | (layer0_outputs[1463]);
    assign layer1_outputs[4859] = ~((layer0_outputs[1860]) | (layer0_outputs[1281]));
    assign layer1_outputs[4860] = layer0_outputs[3207];
    assign layer1_outputs[4861] = 1'b0;
    assign layer1_outputs[4862] = (layer0_outputs[1734]) & ~(layer0_outputs[4539]);
    assign layer1_outputs[4863] = ~(layer0_outputs[1347]) | (layer0_outputs[2397]);
    assign layer1_outputs[4864] = ~((layer0_outputs[1175]) & (layer0_outputs[2832]));
    assign layer1_outputs[4865] = 1'b0;
    assign layer1_outputs[4866] = 1'b1;
    assign layer1_outputs[4867] = ~(layer0_outputs[1314]) | (layer0_outputs[2935]);
    assign layer1_outputs[4868] = ~(layer0_outputs[4500]) | (layer0_outputs[2005]);
    assign layer1_outputs[4869] = ~((layer0_outputs[4567]) & (layer0_outputs[404]));
    assign layer1_outputs[4870] = 1'b1;
    assign layer1_outputs[4871] = 1'b1;
    assign layer1_outputs[4872] = ~((layer0_outputs[3524]) | (layer0_outputs[1262]));
    assign layer1_outputs[4873] = (layer0_outputs[1694]) & (layer0_outputs[4931]);
    assign layer1_outputs[4874] = 1'b1;
    assign layer1_outputs[4875] = 1'b1;
    assign layer1_outputs[4876] = 1'b0;
    assign layer1_outputs[4877] = layer0_outputs[3735];
    assign layer1_outputs[4878] = layer0_outputs[448];
    assign layer1_outputs[4879] = (layer0_outputs[3104]) & (layer0_outputs[4092]);
    assign layer1_outputs[4880] = ~(layer0_outputs[3351]);
    assign layer1_outputs[4881] = ~(layer0_outputs[737]) | (layer0_outputs[2317]);
    assign layer1_outputs[4882] = layer0_outputs[365];
    assign layer1_outputs[4883] = 1'b1;
    assign layer1_outputs[4884] = ~((layer0_outputs[4023]) ^ (layer0_outputs[1356]));
    assign layer1_outputs[4885] = ~(layer0_outputs[2710]) | (layer0_outputs[1608]);
    assign layer1_outputs[4886] = (layer0_outputs[1895]) & (layer0_outputs[4109]);
    assign layer1_outputs[4887] = (layer0_outputs[3921]) & ~(layer0_outputs[1936]);
    assign layer1_outputs[4888] = ~((layer0_outputs[727]) | (layer0_outputs[2331]));
    assign layer1_outputs[4889] = layer0_outputs[2424];
    assign layer1_outputs[4890] = 1'b1;
    assign layer1_outputs[4891] = ~(layer0_outputs[250]) | (layer0_outputs[69]);
    assign layer1_outputs[4892] = (layer0_outputs[447]) & (layer0_outputs[4927]);
    assign layer1_outputs[4893] = (layer0_outputs[835]) & (layer0_outputs[3568]);
    assign layer1_outputs[4894] = ~(layer0_outputs[4614]);
    assign layer1_outputs[4895] = ~(layer0_outputs[1864]);
    assign layer1_outputs[4896] = (layer0_outputs[4822]) & ~(layer0_outputs[2304]);
    assign layer1_outputs[4897] = 1'b0;
    assign layer1_outputs[4898] = ~(layer0_outputs[3897]);
    assign layer1_outputs[4899] = ~((layer0_outputs[387]) ^ (layer0_outputs[4216]));
    assign layer1_outputs[4900] = ~(layer0_outputs[1059]);
    assign layer1_outputs[4901] = 1'b0;
    assign layer1_outputs[4902] = layer0_outputs[453];
    assign layer1_outputs[4903] = (layer0_outputs[583]) & (layer0_outputs[3090]);
    assign layer1_outputs[4904] = layer0_outputs[2791];
    assign layer1_outputs[4905] = ~(layer0_outputs[984]) | (layer0_outputs[4006]);
    assign layer1_outputs[4906] = 1'b1;
    assign layer1_outputs[4907] = ~(layer0_outputs[2629]);
    assign layer1_outputs[4908] = (layer0_outputs[3816]) | (layer0_outputs[1396]);
    assign layer1_outputs[4909] = 1'b1;
    assign layer1_outputs[4910] = layer0_outputs[4000];
    assign layer1_outputs[4911] = ~(layer0_outputs[3178]);
    assign layer1_outputs[4912] = layer0_outputs[2922];
    assign layer1_outputs[4913] = 1'b0;
    assign layer1_outputs[4914] = layer0_outputs[4033];
    assign layer1_outputs[4915] = 1'b0;
    assign layer1_outputs[4916] = ~((layer0_outputs[1960]) & (layer0_outputs[808]));
    assign layer1_outputs[4917] = ~(layer0_outputs[2992]);
    assign layer1_outputs[4918] = 1'b0;
    assign layer1_outputs[4919] = layer0_outputs[2814];
    assign layer1_outputs[4920] = ~((layer0_outputs[89]) & (layer0_outputs[168]));
    assign layer1_outputs[4921] = layer0_outputs[2565];
    assign layer1_outputs[4922] = (layer0_outputs[2566]) & ~(layer0_outputs[159]);
    assign layer1_outputs[4923] = ~((layer0_outputs[3808]) | (layer0_outputs[2910]));
    assign layer1_outputs[4924] = 1'b0;
    assign layer1_outputs[4925] = (layer0_outputs[1676]) & ~(layer0_outputs[4324]);
    assign layer1_outputs[4926] = ~((layer0_outputs[5092]) | (layer0_outputs[2021]));
    assign layer1_outputs[4927] = (layer0_outputs[2666]) & (layer0_outputs[4077]);
    assign layer1_outputs[4928] = 1'b0;
    assign layer1_outputs[4929] = layer0_outputs[2689];
    assign layer1_outputs[4930] = ~(layer0_outputs[2888]);
    assign layer1_outputs[4931] = ~((layer0_outputs[5053]) | (layer0_outputs[772]));
    assign layer1_outputs[4932] = (layer0_outputs[477]) & (layer0_outputs[1271]);
    assign layer1_outputs[4933] = ~(layer0_outputs[1661]);
    assign layer1_outputs[4934] = ~(layer0_outputs[5100]);
    assign layer1_outputs[4935] = (layer0_outputs[3626]) & (layer0_outputs[1306]);
    assign layer1_outputs[4936] = ~(layer0_outputs[1683]) | (layer0_outputs[2287]);
    assign layer1_outputs[4937] = layer0_outputs[3758];
    assign layer1_outputs[4938] = ~(layer0_outputs[1419]);
    assign layer1_outputs[4939] = (layer0_outputs[2770]) & (layer0_outputs[2266]);
    assign layer1_outputs[4940] = ~(layer0_outputs[1122]);
    assign layer1_outputs[4941] = 1'b0;
    assign layer1_outputs[4942] = ~((layer0_outputs[1945]) | (layer0_outputs[759]));
    assign layer1_outputs[4943] = 1'b0;
    assign layer1_outputs[4944] = ~((layer0_outputs[586]) | (layer0_outputs[3369]));
    assign layer1_outputs[4945] = (layer0_outputs[3402]) & ~(layer0_outputs[3461]);
    assign layer1_outputs[4946] = ~((layer0_outputs[891]) & (layer0_outputs[1759]));
    assign layer1_outputs[4947] = (layer0_outputs[731]) | (layer0_outputs[3710]);
    assign layer1_outputs[4948] = layer0_outputs[1910];
    assign layer1_outputs[4949] = ~(layer0_outputs[4730]) | (layer0_outputs[3139]);
    assign layer1_outputs[4950] = (layer0_outputs[562]) | (layer0_outputs[455]);
    assign layer1_outputs[4951] = ~(layer0_outputs[1873]) | (layer0_outputs[2674]);
    assign layer1_outputs[4952] = ~((layer0_outputs[775]) | (layer0_outputs[1616]));
    assign layer1_outputs[4953] = (layer0_outputs[3202]) & ~(layer0_outputs[3909]);
    assign layer1_outputs[4954] = ~((layer0_outputs[523]) & (layer0_outputs[2817]));
    assign layer1_outputs[4955] = (layer0_outputs[5106]) | (layer0_outputs[5017]);
    assign layer1_outputs[4956] = (layer0_outputs[1544]) & ~(layer0_outputs[1830]);
    assign layer1_outputs[4957] = ~(layer0_outputs[787]);
    assign layer1_outputs[4958] = 1'b1;
    assign layer1_outputs[4959] = (layer0_outputs[2296]) ^ (layer0_outputs[1216]);
    assign layer1_outputs[4960] = layer0_outputs[5017];
    assign layer1_outputs[4961] = ~(layer0_outputs[3886]);
    assign layer1_outputs[4962] = ~(layer0_outputs[4672]);
    assign layer1_outputs[4963] = ~((layer0_outputs[2753]) & (layer0_outputs[141]));
    assign layer1_outputs[4964] = layer0_outputs[2338];
    assign layer1_outputs[4965] = ~(layer0_outputs[16]) | (layer0_outputs[4430]);
    assign layer1_outputs[4966] = (layer0_outputs[4896]) | (layer0_outputs[1031]);
    assign layer1_outputs[4967] = 1'b0;
    assign layer1_outputs[4968] = (layer0_outputs[212]) & ~(layer0_outputs[2020]);
    assign layer1_outputs[4969] = 1'b0;
    assign layer1_outputs[4970] = ~(layer0_outputs[3616]);
    assign layer1_outputs[4971] = ~((layer0_outputs[891]) | (layer0_outputs[507]));
    assign layer1_outputs[4972] = 1'b1;
    assign layer1_outputs[4973] = 1'b1;
    assign layer1_outputs[4974] = ~((layer0_outputs[1774]) ^ (layer0_outputs[1623]));
    assign layer1_outputs[4975] = ~(layer0_outputs[603]) | (layer0_outputs[759]);
    assign layer1_outputs[4976] = ~(layer0_outputs[102]);
    assign layer1_outputs[4977] = 1'b1;
    assign layer1_outputs[4978] = (layer0_outputs[2277]) | (layer0_outputs[4580]);
    assign layer1_outputs[4979] = layer0_outputs[3625];
    assign layer1_outputs[4980] = ~(layer0_outputs[4761]);
    assign layer1_outputs[4981] = (layer0_outputs[1165]) & (layer0_outputs[150]);
    assign layer1_outputs[4982] = 1'b1;
    assign layer1_outputs[4983] = (layer0_outputs[3831]) | (layer0_outputs[1304]);
    assign layer1_outputs[4984] = ~(layer0_outputs[4319]);
    assign layer1_outputs[4985] = ~(layer0_outputs[3380]) | (layer0_outputs[2495]);
    assign layer1_outputs[4986] = ~(layer0_outputs[197]);
    assign layer1_outputs[4987] = (layer0_outputs[3537]) & ~(layer0_outputs[221]);
    assign layer1_outputs[4988] = layer0_outputs[2583];
    assign layer1_outputs[4989] = layer0_outputs[1391];
    assign layer1_outputs[4990] = ~((layer0_outputs[2488]) | (layer0_outputs[3374]));
    assign layer1_outputs[4991] = ~(layer0_outputs[2936]);
    assign layer1_outputs[4992] = ~(layer0_outputs[4820]);
    assign layer1_outputs[4993] = ~(layer0_outputs[4874]);
    assign layer1_outputs[4994] = ~((layer0_outputs[3236]) | (layer0_outputs[2316]));
    assign layer1_outputs[4995] = layer0_outputs[2231];
    assign layer1_outputs[4996] = ~(layer0_outputs[5072]) | (layer0_outputs[2906]);
    assign layer1_outputs[4997] = (layer0_outputs[1459]) & (layer0_outputs[3534]);
    assign layer1_outputs[4998] = ~(layer0_outputs[4758]);
    assign layer1_outputs[4999] = ~((layer0_outputs[587]) | (layer0_outputs[3129]));
    assign layer1_outputs[5000] = ~(layer0_outputs[1975]);
    assign layer1_outputs[5001] = (layer0_outputs[4046]) & ~(layer0_outputs[2185]);
    assign layer1_outputs[5002] = (layer0_outputs[4416]) ^ (layer0_outputs[1568]);
    assign layer1_outputs[5003] = ~((layer0_outputs[2712]) | (layer0_outputs[1397]));
    assign layer1_outputs[5004] = layer0_outputs[2538];
    assign layer1_outputs[5005] = (layer0_outputs[2458]) & (layer0_outputs[3558]);
    assign layer1_outputs[5006] = (layer0_outputs[918]) & (layer0_outputs[3257]);
    assign layer1_outputs[5007] = (layer0_outputs[495]) & ~(layer0_outputs[3633]);
    assign layer1_outputs[5008] = (layer0_outputs[450]) & ~(layer0_outputs[1458]);
    assign layer1_outputs[5009] = (layer0_outputs[620]) & ~(layer0_outputs[3319]);
    assign layer1_outputs[5010] = ~((layer0_outputs[4236]) ^ (layer0_outputs[961]));
    assign layer1_outputs[5011] = 1'b1;
    assign layer1_outputs[5012] = 1'b1;
    assign layer1_outputs[5013] = 1'b1;
    assign layer1_outputs[5014] = ~(layer0_outputs[4786]);
    assign layer1_outputs[5015] = ~((layer0_outputs[3698]) & (layer0_outputs[2442]));
    assign layer1_outputs[5016] = layer0_outputs[2305];
    assign layer1_outputs[5017] = (layer0_outputs[1126]) | (layer0_outputs[4882]);
    assign layer1_outputs[5018] = (layer0_outputs[1879]) & (layer0_outputs[624]);
    assign layer1_outputs[5019] = ~(layer0_outputs[2179]);
    assign layer1_outputs[5020] = 1'b0;
    assign layer1_outputs[5021] = (layer0_outputs[2668]) & ~(layer0_outputs[3690]);
    assign layer1_outputs[5022] = (layer0_outputs[1607]) | (layer0_outputs[457]);
    assign layer1_outputs[5023] = ~((layer0_outputs[4360]) | (layer0_outputs[4925]));
    assign layer1_outputs[5024] = (layer0_outputs[4165]) & ~(layer0_outputs[3442]);
    assign layer1_outputs[5025] = (layer0_outputs[4703]) | (layer0_outputs[903]);
    assign layer1_outputs[5026] = (layer0_outputs[628]) & ~(layer0_outputs[4446]);
    assign layer1_outputs[5027] = (layer0_outputs[130]) & (layer0_outputs[2460]);
    assign layer1_outputs[5028] = ~(layer0_outputs[1827]) | (layer0_outputs[2510]);
    assign layer1_outputs[5029] = layer0_outputs[2049];
    assign layer1_outputs[5030] = (layer0_outputs[3401]) & ~(layer0_outputs[786]);
    assign layer1_outputs[5031] = (layer0_outputs[2717]) & ~(layer0_outputs[802]);
    assign layer1_outputs[5032] = (layer0_outputs[1638]) & (layer0_outputs[751]);
    assign layer1_outputs[5033] = (layer0_outputs[1210]) & ~(layer0_outputs[787]);
    assign layer1_outputs[5034] = ~((layer0_outputs[3092]) | (layer0_outputs[4155]));
    assign layer1_outputs[5035] = layer0_outputs[4073];
    assign layer1_outputs[5036] = ~(layer0_outputs[3343]) | (layer0_outputs[2729]);
    assign layer1_outputs[5037] = layer0_outputs[3544];
    assign layer1_outputs[5038] = layer0_outputs[4713];
    assign layer1_outputs[5039] = 1'b0;
    assign layer1_outputs[5040] = (layer0_outputs[3743]) & (layer0_outputs[4604]);
    assign layer1_outputs[5041] = (layer0_outputs[3124]) | (layer0_outputs[2156]);
    assign layer1_outputs[5042] = ~((layer0_outputs[4432]) | (layer0_outputs[2340]));
    assign layer1_outputs[5043] = layer0_outputs[1025];
    assign layer1_outputs[5044] = ~((layer0_outputs[672]) | (layer0_outputs[4539]));
    assign layer1_outputs[5045] = ~((layer0_outputs[1424]) | (layer0_outputs[1081]));
    assign layer1_outputs[5046] = (layer0_outputs[3751]) & ~(layer0_outputs[2947]);
    assign layer1_outputs[5047] = layer0_outputs[1752];
    assign layer1_outputs[5048] = ~(layer0_outputs[2297]);
    assign layer1_outputs[5049] = ~((layer0_outputs[3260]) & (layer0_outputs[1839]));
    assign layer1_outputs[5050] = 1'b0;
    assign layer1_outputs[5051] = ~((layer0_outputs[4846]) ^ (layer0_outputs[1829]));
    assign layer1_outputs[5052] = (layer0_outputs[3574]) | (layer0_outputs[132]);
    assign layer1_outputs[5053] = ~((layer0_outputs[862]) | (layer0_outputs[269]));
    assign layer1_outputs[5054] = (layer0_outputs[4649]) & ~(layer0_outputs[4757]);
    assign layer1_outputs[5055] = layer0_outputs[10];
    assign layer1_outputs[5056] = layer0_outputs[2322];
    assign layer1_outputs[5057] = (layer0_outputs[1696]) & (layer0_outputs[3320]);
    assign layer1_outputs[5058] = layer0_outputs[2683];
    assign layer1_outputs[5059] = ~(layer0_outputs[3173]);
    assign layer1_outputs[5060] = (layer0_outputs[4151]) ^ (layer0_outputs[668]);
    assign layer1_outputs[5061] = ~((layer0_outputs[3240]) & (layer0_outputs[3862]));
    assign layer1_outputs[5062] = (layer0_outputs[385]) & ~(layer0_outputs[3089]);
    assign layer1_outputs[5063] = 1'b1;
    assign layer1_outputs[5064] = 1'b1;
    assign layer1_outputs[5065] = layer0_outputs[1082];
    assign layer1_outputs[5066] = (layer0_outputs[1684]) & ~(layer0_outputs[1160]);
    assign layer1_outputs[5067] = ~(layer0_outputs[4261]);
    assign layer1_outputs[5068] = ~(layer0_outputs[2389]) | (layer0_outputs[2491]);
    assign layer1_outputs[5069] = (layer0_outputs[3832]) & ~(layer0_outputs[1193]);
    assign layer1_outputs[5070] = ~(layer0_outputs[3908]);
    assign layer1_outputs[5071] = (layer0_outputs[1550]) & ~(layer0_outputs[179]);
    assign layer1_outputs[5072] = 1'b1;
    assign layer1_outputs[5073] = ~((layer0_outputs[2985]) & (layer0_outputs[197]));
    assign layer1_outputs[5074] = ~(layer0_outputs[277]) | (layer0_outputs[4382]);
    assign layer1_outputs[5075] = ~(layer0_outputs[647]);
    assign layer1_outputs[5076] = ~((layer0_outputs[629]) & (layer0_outputs[846]));
    assign layer1_outputs[5077] = layer0_outputs[165];
    assign layer1_outputs[5078] = (layer0_outputs[1570]) & (layer0_outputs[136]);
    assign layer1_outputs[5079] = (layer0_outputs[3339]) | (layer0_outputs[4483]);
    assign layer1_outputs[5080] = (layer0_outputs[2457]) & ~(layer0_outputs[4913]);
    assign layer1_outputs[5081] = (layer0_outputs[4856]) & (layer0_outputs[526]);
    assign layer1_outputs[5082] = ~(layer0_outputs[2218]) | (layer0_outputs[2536]);
    assign layer1_outputs[5083] = 1'b1;
    assign layer1_outputs[5084] = layer0_outputs[3149];
    assign layer1_outputs[5085] = ~(layer0_outputs[3978]);
    assign layer1_outputs[5086] = 1'b1;
    assign layer1_outputs[5087] = ~(layer0_outputs[1746]);
    assign layer1_outputs[5088] = ~(layer0_outputs[3318]) | (layer0_outputs[2457]);
    assign layer1_outputs[5089] = (layer0_outputs[2085]) & ~(layer0_outputs[3379]);
    assign layer1_outputs[5090] = ~((layer0_outputs[2651]) & (layer0_outputs[3216]));
    assign layer1_outputs[5091] = (layer0_outputs[4361]) & ~(layer0_outputs[2329]);
    assign layer1_outputs[5092] = ~((layer0_outputs[482]) ^ (layer0_outputs[2831]));
    assign layer1_outputs[5093] = (layer0_outputs[430]) & ~(layer0_outputs[2230]);
    assign layer1_outputs[5094] = (layer0_outputs[861]) & (layer0_outputs[2060]);
    assign layer1_outputs[5095] = layer0_outputs[2970];
    assign layer1_outputs[5096] = ~(layer0_outputs[4742]);
    assign layer1_outputs[5097] = layer0_outputs[1791];
    assign layer1_outputs[5098] = (layer0_outputs[3850]) & ~(layer0_outputs[121]);
    assign layer1_outputs[5099] = layer0_outputs[1908];
    assign layer1_outputs[5100] = ~(layer0_outputs[3872]) | (layer0_outputs[2807]);
    assign layer1_outputs[5101] = 1'b0;
    assign layer1_outputs[5102] = (layer0_outputs[1834]) & ~(layer0_outputs[4627]);
    assign layer1_outputs[5103] = 1'b1;
    assign layer1_outputs[5104] = (layer0_outputs[699]) & ~(layer0_outputs[4212]);
    assign layer1_outputs[5105] = layer0_outputs[3889];
    assign layer1_outputs[5106] = (layer0_outputs[2037]) & ~(layer0_outputs[2400]);
    assign layer1_outputs[5107] = (layer0_outputs[691]) & (layer0_outputs[2559]);
    assign layer1_outputs[5108] = ~((layer0_outputs[3218]) | (layer0_outputs[2375]));
    assign layer1_outputs[5109] = 1'b0;
    assign layer1_outputs[5110] = ~((layer0_outputs[817]) | (layer0_outputs[2767]));
    assign layer1_outputs[5111] = layer0_outputs[187];
    assign layer1_outputs[5112] = 1'b1;
    assign layer1_outputs[5113] = ~((layer0_outputs[5064]) ^ (layer0_outputs[924]));
    assign layer1_outputs[5114] = layer0_outputs[1247];
    assign layer1_outputs[5115] = ~((layer0_outputs[3404]) | (layer0_outputs[180]));
    assign layer1_outputs[5116] = 1'b1;
    assign layer1_outputs[5117] = ~(layer0_outputs[4180]);
    assign layer1_outputs[5118] = 1'b0;
    assign layer1_outputs[5119] = ~(layer0_outputs[3421]) | (layer0_outputs[4814]);
    assign layer2_outputs[0] = ~((layer1_outputs[4728]) & (layer1_outputs[5085]));
    assign layer2_outputs[1] = (layer1_outputs[581]) & ~(layer1_outputs[3177]);
    assign layer2_outputs[2] = ~(layer1_outputs[1384]) | (layer1_outputs[5043]);
    assign layer2_outputs[3] = ~(layer1_outputs[4076]);
    assign layer2_outputs[4] = ~((layer1_outputs[1855]) | (layer1_outputs[1065]));
    assign layer2_outputs[5] = ~(layer1_outputs[354]);
    assign layer2_outputs[6] = ~(layer1_outputs[1089]) | (layer1_outputs[2129]);
    assign layer2_outputs[7] = (layer1_outputs[288]) & (layer1_outputs[1166]);
    assign layer2_outputs[8] = 1'b0;
    assign layer2_outputs[9] = layer1_outputs[1398];
    assign layer2_outputs[10] = ~(layer1_outputs[686]);
    assign layer2_outputs[11] = layer1_outputs[3179];
    assign layer2_outputs[12] = 1'b1;
    assign layer2_outputs[13] = ~(layer1_outputs[4101]);
    assign layer2_outputs[14] = ~((layer1_outputs[1111]) & (layer1_outputs[1798]));
    assign layer2_outputs[15] = ~(layer1_outputs[2510]) | (layer1_outputs[4915]);
    assign layer2_outputs[16] = ~(layer1_outputs[237]) | (layer1_outputs[3561]);
    assign layer2_outputs[17] = 1'b0;
    assign layer2_outputs[18] = layer1_outputs[4193];
    assign layer2_outputs[19] = (layer1_outputs[393]) & ~(layer1_outputs[193]);
    assign layer2_outputs[20] = ~(layer1_outputs[132]);
    assign layer2_outputs[21] = ~((layer1_outputs[4371]) | (layer1_outputs[3400]));
    assign layer2_outputs[22] = ~(layer1_outputs[1221]);
    assign layer2_outputs[23] = layer1_outputs[2484];
    assign layer2_outputs[24] = 1'b0;
    assign layer2_outputs[25] = ~(layer1_outputs[3328]);
    assign layer2_outputs[26] = layer1_outputs[50];
    assign layer2_outputs[27] = (layer1_outputs[4804]) | (layer1_outputs[2639]);
    assign layer2_outputs[28] = ~((layer1_outputs[2939]) ^ (layer1_outputs[4305]));
    assign layer2_outputs[29] = ~(layer1_outputs[472]);
    assign layer2_outputs[30] = layer1_outputs[3532];
    assign layer2_outputs[31] = ~(layer1_outputs[929]);
    assign layer2_outputs[32] = (layer1_outputs[3601]) & (layer1_outputs[4602]);
    assign layer2_outputs[33] = ~(layer1_outputs[1529]);
    assign layer2_outputs[34] = ~((layer1_outputs[2637]) & (layer1_outputs[3842]));
    assign layer2_outputs[35] = (layer1_outputs[1392]) & (layer1_outputs[1853]);
    assign layer2_outputs[36] = ~((layer1_outputs[1447]) | (layer1_outputs[4032]));
    assign layer2_outputs[37] = (layer1_outputs[1230]) & ~(layer1_outputs[5006]);
    assign layer2_outputs[38] = layer1_outputs[1112];
    assign layer2_outputs[39] = layer1_outputs[5004];
    assign layer2_outputs[40] = ~((layer1_outputs[4282]) | (layer1_outputs[1291]));
    assign layer2_outputs[41] = ~(layer1_outputs[2741]) | (layer1_outputs[4044]);
    assign layer2_outputs[42] = ~(layer1_outputs[3342]);
    assign layer2_outputs[43] = 1'b0;
    assign layer2_outputs[44] = 1'b0;
    assign layer2_outputs[45] = layer1_outputs[4845];
    assign layer2_outputs[46] = layer1_outputs[3150];
    assign layer2_outputs[47] = ~(layer1_outputs[862]) | (layer1_outputs[3114]);
    assign layer2_outputs[48] = 1'b0;
    assign layer2_outputs[49] = ~(layer1_outputs[2851]) | (layer1_outputs[2815]);
    assign layer2_outputs[50] = (layer1_outputs[514]) & ~(layer1_outputs[3703]);
    assign layer2_outputs[51] = (layer1_outputs[3316]) & ~(layer1_outputs[4948]);
    assign layer2_outputs[52] = ~(layer1_outputs[1187]) | (layer1_outputs[2050]);
    assign layer2_outputs[53] = layer1_outputs[1209];
    assign layer2_outputs[54] = ~((layer1_outputs[3674]) & (layer1_outputs[1497]));
    assign layer2_outputs[55] = ~((layer1_outputs[2989]) | (layer1_outputs[1269]));
    assign layer2_outputs[56] = (layer1_outputs[1646]) & (layer1_outputs[2290]);
    assign layer2_outputs[57] = (layer1_outputs[2840]) & ~(layer1_outputs[4257]);
    assign layer2_outputs[58] = layer1_outputs[4310];
    assign layer2_outputs[59] = layer1_outputs[3774];
    assign layer2_outputs[60] = (layer1_outputs[239]) & ~(layer1_outputs[3123]);
    assign layer2_outputs[61] = layer1_outputs[4851];
    assign layer2_outputs[62] = ~(layer1_outputs[3210]) | (layer1_outputs[1437]);
    assign layer2_outputs[63] = ~((layer1_outputs[1930]) | (layer1_outputs[2266]));
    assign layer2_outputs[64] = (layer1_outputs[864]) | (layer1_outputs[2642]);
    assign layer2_outputs[65] = ~((layer1_outputs[5096]) & (layer1_outputs[1318]));
    assign layer2_outputs[66] = 1'b1;
    assign layer2_outputs[67] = (layer1_outputs[4944]) & ~(layer1_outputs[4354]);
    assign layer2_outputs[68] = ~((layer1_outputs[2713]) & (layer1_outputs[1575]));
    assign layer2_outputs[69] = (layer1_outputs[3275]) & (layer1_outputs[4923]);
    assign layer2_outputs[70] = ~((layer1_outputs[3181]) & (layer1_outputs[781]));
    assign layer2_outputs[71] = (layer1_outputs[2025]) & ~(layer1_outputs[1017]);
    assign layer2_outputs[72] = ~(layer1_outputs[2619]);
    assign layer2_outputs[73] = (layer1_outputs[1252]) & (layer1_outputs[2723]);
    assign layer2_outputs[74] = ~(layer1_outputs[4896]);
    assign layer2_outputs[75] = layer1_outputs[1956];
    assign layer2_outputs[76] = layer1_outputs[4078];
    assign layer2_outputs[77] = (layer1_outputs[4404]) | (layer1_outputs[238]);
    assign layer2_outputs[78] = ~(layer1_outputs[1587]);
    assign layer2_outputs[79] = (layer1_outputs[3084]) ^ (layer1_outputs[4954]);
    assign layer2_outputs[80] = ~(layer1_outputs[1657]) | (layer1_outputs[4245]);
    assign layer2_outputs[81] = layer1_outputs[3815];
    assign layer2_outputs[82] = layer1_outputs[2954];
    assign layer2_outputs[83] = layer1_outputs[2711];
    assign layer2_outputs[84] = 1'b1;
    assign layer2_outputs[85] = 1'b1;
    assign layer2_outputs[86] = ~(layer1_outputs[1829]);
    assign layer2_outputs[87] = (layer1_outputs[5002]) & ~(layer1_outputs[2141]);
    assign layer2_outputs[88] = (layer1_outputs[3413]) & ~(layer1_outputs[4884]);
    assign layer2_outputs[89] = layer1_outputs[4981];
    assign layer2_outputs[90] = ~(layer1_outputs[675]);
    assign layer2_outputs[91] = 1'b1;
    assign layer2_outputs[92] = 1'b0;
    assign layer2_outputs[93] = ~(layer1_outputs[3202]);
    assign layer2_outputs[94] = 1'b1;
    assign layer2_outputs[95] = ~(layer1_outputs[3908]) | (layer1_outputs[1750]);
    assign layer2_outputs[96] = ~(layer1_outputs[3442]);
    assign layer2_outputs[97] = (layer1_outputs[2993]) | (layer1_outputs[4733]);
    assign layer2_outputs[98] = ~((layer1_outputs[1021]) | (layer1_outputs[3979]));
    assign layer2_outputs[99] = (layer1_outputs[4900]) & (layer1_outputs[3657]);
    assign layer2_outputs[100] = ~(layer1_outputs[3648]);
    assign layer2_outputs[101] = (layer1_outputs[3481]) & ~(layer1_outputs[1832]);
    assign layer2_outputs[102] = ~(layer1_outputs[4745]) | (layer1_outputs[4061]);
    assign layer2_outputs[103] = ~((layer1_outputs[843]) & (layer1_outputs[4049]));
    assign layer2_outputs[104] = ~(layer1_outputs[1885]);
    assign layer2_outputs[105] = ~(layer1_outputs[4447]) | (layer1_outputs[3208]);
    assign layer2_outputs[106] = layer1_outputs[2921];
    assign layer2_outputs[107] = ~(layer1_outputs[899]);
    assign layer2_outputs[108] = (layer1_outputs[4881]) & ~(layer1_outputs[3089]);
    assign layer2_outputs[109] = ~(layer1_outputs[4456]) | (layer1_outputs[3516]);
    assign layer2_outputs[110] = 1'b0;
    assign layer2_outputs[111] = 1'b0;
    assign layer2_outputs[112] = ~(layer1_outputs[1866]) | (layer1_outputs[3223]);
    assign layer2_outputs[113] = 1'b1;
    assign layer2_outputs[114] = ~(layer1_outputs[4364]);
    assign layer2_outputs[115] = ~((layer1_outputs[424]) & (layer1_outputs[2898]));
    assign layer2_outputs[116] = layer1_outputs[197];
    assign layer2_outputs[117] = 1'b1;
    assign layer2_outputs[118] = layer1_outputs[4858];
    assign layer2_outputs[119] = ~(layer1_outputs[98]) | (layer1_outputs[3312]);
    assign layer2_outputs[120] = 1'b0;
    assign layer2_outputs[121] = layer1_outputs[4907];
    assign layer2_outputs[122] = layer1_outputs[3585];
    assign layer2_outputs[123] = ~(layer1_outputs[951]) | (layer1_outputs[4726]);
    assign layer2_outputs[124] = ~(layer1_outputs[1086]) | (layer1_outputs[484]);
    assign layer2_outputs[125] = 1'b1;
    assign layer2_outputs[126] = layer1_outputs[2204];
    assign layer2_outputs[127] = ~(layer1_outputs[682]) | (layer1_outputs[2757]);
    assign layer2_outputs[128] = ~(layer1_outputs[3474]);
    assign layer2_outputs[129] = ~((layer1_outputs[4978]) & (layer1_outputs[848]));
    assign layer2_outputs[130] = layer1_outputs[829];
    assign layer2_outputs[131] = (layer1_outputs[188]) & ~(layer1_outputs[346]);
    assign layer2_outputs[132] = ~((layer1_outputs[3788]) | (layer1_outputs[3853]));
    assign layer2_outputs[133] = ~(layer1_outputs[2372]);
    assign layer2_outputs[134] = ~(layer1_outputs[339]);
    assign layer2_outputs[135] = 1'b1;
    assign layer2_outputs[136] = (layer1_outputs[2064]) | (layer1_outputs[4698]);
    assign layer2_outputs[137] = layer1_outputs[2076];
    assign layer2_outputs[138] = (layer1_outputs[2013]) ^ (layer1_outputs[3543]);
    assign layer2_outputs[139] = ~(layer1_outputs[1005]);
    assign layer2_outputs[140] = 1'b0;
    assign layer2_outputs[141] = ~((layer1_outputs[118]) | (layer1_outputs[4279]));
    assign layer2_outputs[142] = 1'b1;
    assign layer2_outputs[143] = ~(layer1_outputs[4581]);
    assign layer2_outputs[144] = (layer1_outputs[1164]) | (layer1_outputs[3142]);
    assign layer2_outputs[145] = ~((layer1_outputs[596]) & (layer1_outputs[262]));
    assign layer2_outputs[146] = ~(layer1_outputs[2153]);
    assign layer2_outputs[147] = ~(layer1_outputs[481]) | (layer1_outputs[4534]);
    assign layer2_outputs[148] = 1'b1;
    assign layer2_outputs[149] = (layer1_outputs[845]) | (layer1_outputs[4842]);
    assign layer2_outputs[150] = ~(layer1_outputs[2602]);
    assign layer2_outputs[151] = layer1_outputs[4259];
    assign layer2_outputs[152] = ~((layer1_outputs[3984]) | (layer1_outputs[2105]));
    assign layer2_outputs[153] = ~(layer1_outputs[4546]);
    assign layer2_outputs[154] = layer1_outputs[1267];
    assign layer2_outputs[155] = ~((layer1_outputs[4400]) ^ (layer1_outputs[1589]));
    assign layer2_outputs[156] = (layer1_outputs[695]) ^ (layer1_outputs[4846]);
    assign layer2_outputs[157] = layer1_outputs[2277];
    assign layer2_outputs[158] = layer1_outputs[3236];
    assign layer2_outputs[159] = (layer1_outputs[2919]) | (layer1_outputs[2258]);
    assign layer2_outputs[160] = layer1_outputs[1356];
    assign layer2_outputs[161] = (layer1_outputs[161]) & ~(layer1_outputs[2343]);
    assign layer2_outputs[162] = 1'b0;
    assign layer2_outputs[163] = ~(layer1_outputs[1140]) | (layer1_outputs[4495]);
    assign layer2_outputs[164] = ~(layer1_outputs[4472]);
    assign layer2_outputs[165] = (layer1_outputs[4624]) & (layer1_outputs[4707]);
    assign layer2_outputs[166] = (layer1_outputs[454]) & (layer1_outputs[2404]);
    assign layer2_outputs[167] = layer1_outputs[294];
    assign layer2_outputs[168] = ~(layer1_outputs[2802]) | (layer1_outputs[343]);
    assign layer2_outputs[169] = layer1_outputs[693];
    assign layer2_outputs[170] = 1'b0;
    assign layer2_outputs[171] = ~(layer1_outputs[2443]);
    assign layer2_outputs[172] = (layer1_outputs[875]) & (layer1_outputs[4678]);
    assign layer2_outputs[173] = (layer1_outputs[4690]) & ~(layer1_outputs[369]);
    assign layer2_outputs[174] = ~((layer1_outputs[996]) | (layer1_outputs[75]));
    assign layer2_outputs[175] = (layer1_outputs[4276]) & (layer1_outputs[4470]);
    assign layer2_outputs[176] = (layer1_outputs[1881]) & ~(layer1_outputs[4317]);
    assign layer2_outputs[177] = ~((layer1_outputs[3491]) & (layer1_outputs[1010]));
    assign layer2_outputs[178] = ~((layer1_outputs[4237]) | (layer1_outputs[203]));
    assign layer2_outputs[179] = ~((layer1_outputs[854]) & (layer1_outputs[2329]));
    assign layer2_outputs[180] = (layer1_outputs[4391]) & (layer1_outputs[127]);
    assign layer2_outputs[181] = ~((layer1_outputs[4418]) | (layer1_outputs[1851]));
    assign layer2_outputs[182] = ~(layer1_outputs[3329]) | (layer1_outputs[4429]);
    assign layer2_outputs[183] = layer1_outputs[89];
    assign layer2_outputs[184] = 1'b0;
    assign layer2_outputs[185] = ~(layer1_outputs[1350]);
    assign layer2_outputs[186] = (layer1_outputs[1208]) & ~(layer1_outputs[3614]);
    assign layer2_outputs[187] = 1'b0;
    assign layer2_outputs[188] = (layer1_outputs[3562]) & (layer1_outputs[375]);
    assign layer2_outputs[189] = ~(layer1_outputs[1677]) | (layer1_outputs[3833]);
    assign layer2_outputs[190] = ~(layer1_outputs[2599]);
    assign layer2_outputs[191] = ~((layer1_outputs[1615]) | (layer1_outputs[468]));
    assign layer2_outputs[192] = (layer1_outputs[4010]) & ~(layer1_outputs[1536]);
    assign layer2_outputs[193] = ~(layer1_outputs[2473]);
    assign layer2_outputs[194] = ~(layer1_outputs[4479]) | (layer1_outputs[4039]);
    assign layer2_outputs[195] = layer1_outputs[2873];
    assign layer2_outputs[196] = (layer1_outputs[1595]) & ~(layer1_outputs[4358]);
    assign layer2_outputs[197] = 1'b1;
    assign layer2_outputs[198] = 1'b1;
    assign layer2_outputs[199] = ~(layer1_outputs[881]);
    assign layer2_outputs[200] = (layer1_outputs[635]) & (layer1_outputs[2916]);
    assign layer2_outputs[201] = ~((layer1_outputs[48]) & (layer1_outputs[14]));
    assign layer2_outputs[202] = (layer1_outputs[791]) ^ (layer1_outputs[2982]);
    assign layer2_outputs[203] = ~(layer1_outputs[3131]) | (layer1_outputs[4634]);
    assign layer2_outputs[204] = (layer1_outputs[1475]) | (layer1_outputs[2760]);
    assign layer2_outputs[205] = ~((layer1_outputs[3337]) & (layer1_outputs[3438]));
    assign layer2_outputs[206] = 1'b1;
    assign layer2_outputs[207] = ~(layer1_outputs[144]) | (layer1_outputs[4082]);
    assign layer2_outputs[208] = ~(layer1_outputs[4164]) | (layer1_outputs[24]);
    assign layer2_outputs[209] = ~((layer1_outputs[3157]) & (layer1_outputs[1102]));
    assign layer2_outputs[210] = 1'b0;
    assign layer2_outputs[211] = (layer1_outputs[4873]) & (layer1_outputs[3324]);
    assign layer2_outputs[212] = ~((layer1_outputs[1390]) | (layer1_outputs[1248]));
    assign layer2_outputs[213] = layer1_outputs[990];
    assign layer2_outputs[214] = ~((layer1_outputs[2626]) & (layer1_outputs[2880]));
    assign layer2_outputs[215] = 1'b1;
    assign layer2_outputs[216] = ~(layer1_outputs[3518]);
    assign layer2_outputs[217] = ~(layer1_outputs[2255]);
    assign layer2_outputs[218] = ~(layer1_outputs[1001]);
    assign layer2_outputs[219] = (layer1_outputs[1212]) & ~(layer1_outputs[4170]);
    assign layer2_outputs[220] = ~((layer1_outputs[3730]) | (layer1_outputs[3885]));
    assign layer2_outputs[221] = 1'b0;
    assign layer2_outputs[222] = ~(layer1_outputs[2299]);
    assign layer2_outputs[223] = (layer1_outputs[2517]) & (layer1_outputs[2554]);
    assign layer2_outputs[224] = ~(layer1_outputs[4243]) | (layer1_outputs[2459]);
    assign layer2_outputs[225] = ~(layer1_outputs[1789]);
    assign layer2_outputs[226] = ~(layer1_outputs[4576]) | (layer1_outputs[2737]);
    assign layer2_outputs[227] = ~(layer1_outputs[1813]) | (layer1_outputs[928]);
    assign layer2_outputs[228] = ~(layer1_outputs[2703]);
    assign layer2_outputs[229] = (layer1_outputs[2886]) | (layer1_outputs[4982]);
    assign layer2_outputs[230] = ~(layer1_outputs[4995]) | (layer1_outputs[3034]);
    assign layer2_outputs[231] = ~(layer1_outputs[919]) | (layer1_outputs[1148]);
    assign layer2_outputs[232] = 1'b0;
    assign layer2_outputs[233] = ~(layer1_outputs[969]);
    assign layer2_outputs[234] = layer1_outputs[57];
    assign layer2_outputs[235] = (layer1_outputs[3104]) | (layer1_outputs[2562]);
    assign layer2_outputs[236] = layer1_outputs[620];
    assign layer2_outputs[237] = 1'b1;
    assign layer2_outputs[238] = layer1_outputs[3227];
    assign layer2_outputs[239] = (layer1_outputs[4600]) | (layer1_outputs[1543]);
    assign layer2_outputs[240] = ~(layer1_outputs[2173]);
    assign layer2_outputs[241] = ~((layer1_outputs[1577]) | (layer1_outputs[2685]));
    assign layer2_outputs[242] = ~(layer1_outputs[4815]);
    assign layer2_outputs[243] = (layer1_outputs[4360]) & (layer1_outputs[1110]);
    assign layer2_outputs[244] = 1'b1;
    assign layer2_outputs[245] = ~(layer1_outputs[3963]) | (layer1_outputs[1618]);
    assign layer2_outputs[246] = ~(layer1_outputs[618]) | (layer1_outputs[804]);
    assign layer2_outputs[247] = ~((layer1_outputs[3809]) | (layer1_outputs[2978]));
    assign layer2_outputs[248] = (layer1_outputs[3556]) & (layer1_outputs[3476]);
    assign layer2_outputs[249] = ~(layer1_outputs[4660]);
    assign layer2_outputs[250] = (layer1_outputs[4381]) & ~(layer1_outputs[4700]);
    assign layer2_outputs[251] = ~(layer1_outputs[4747]) | (layer1_outputs[1606]);
    assign layer2_outputs[252] = 1'b0;
    assign layer2_outputs[253] = ~(layer1_outputs[3913]);
    assign layer2_outputs[254] = ~(layer1_outputs[2185]) | (layer1_outputs[1638]);
    assign layer2_outputs[255] = ~(layer1_outputs[4269]) | (layer1_outputs[576]);
    assign layer2_outputs[256] = ~(layer1_outputs[4340]);
    assign layer2_outputs[257] = ~(layer1_outputs[1749]);
    assign layer2_outputs[258] = (layer1_outputs[2304]) & ~(layer1_outputs[3374]);
    assign layer2_outputs[259] = ~((layer1_outputs[2198]) | (layer1_outputs[593]));
    assign layer2_outputs[260] = (layer1_outputs[1882]) | (layer1_outputs[1250]);
    assign layer2_outputs[261] = ~(layer1_outputs[1385]);
    assign layer2_outputs[262] = ~((layer1_outputs[3478]) | (layer1_outputs[395]));
    assign layer2_outputs[263] = (layer1_outputs[2318]) | (layer1_outputs[2084]);
    assign layer2_outputs[264] = ~(layer1_outputs[3960]) | (layer1_outputs[4144]);
    assign layer2_outputs[265] = ~((layer1_outputs[2253]) | (layer1_outputs[250]));
    assign layer2_outputs[266] = ~(layer1_outputs[801]) | (layer1_outputs[2042]);
    assign layer2_outputs[267] = (layer1_outputs[3693]) | (layer1_outputs[1922]);
    assign layer2_outputs[268] = (layer1_outputs[3787]) & ~(layer1_outputs[2166]);
    assign layer2_outputs[269] = (layer1_outputs[3398]) & ~(layer1_outputs[1486]);
    assign layer2_outputs[270] = ~(layer1_outputs[2426]);
    assign layer2_outputs[271] = ~(layer1_outputs[1756]) | (layer1_outputs[4739]);
    assign layer2_outputs[272] = (layer1_outputs[3367]) & (layer1_outputs[2910]);
    assign layer2_outputs[273] = ~(layer1_outputs[155]);
    assign layer2_outputs[274] = (layer1_outputs[3682]) & ~(layer1_outputs[3432]);
    assign layer2_outputs[275] = ~((layer1_outputs[3757]) | (layer1_outputs[4475]));
    assign layer2_outputs[276] = (layer1_outputs[309]) & ~(layer1_outputs[3186]);
    assign layer2_outputs[277] = ~((layer1_outputs[678]) & (layer1_outputs[764]));
    assign layer2_outputs[278] = ~((layer1_outputs[5038]) | (layer1_outputs[3365]));
    assign layer2_outputs[279] = ~(layer1_outputs[2247]) | (layer1_outputs[2011]);
    assign layer2_outputs[280] = ~(layer1_outputs[1409]) | (layer1_outputs[139]);
    assign layer2_outputs[281] = ~(layer1_outputs[4060]) | (layer1_outputs[2690]);
    assign layer2_outputs[282] = ~(layer1_outputs[2998]);
    assign layer2_outputs[283] = ~(layer1_outputs[585]);
    assign layer2_outputs[284] = ~(layer1_outputs[4922]);
    assign layer2_outputs[285] = 1'b1;
    assign layer2_outputs[286] = ~(layer1_outputs[3172]) | (layer1_outputs[1003]);
    assign layer2_outputs[287] = ~(layer1_outputs[1840]) | (layer1_outputs[1114]);
    assign layer2_outputs[288] = 1'b1;
    assign layer2_outputs[289] = ~(layer1_outputs[1906]) | (layer1_outputs[3563]);
    assign layer2_outputs[290] = layer1_outputs[1435];
    assign layer2_outputs[291] = layer1_outputs[2881];
    assign layer2_outputs[292] = ~(layer1_outputs[3160]);
    assign layer2_outputs[293] = ~(layer1_outputs[2836]) | (layer1_outputs[598]);
    assign layer2_outputs[294] = layer1_outputs[4935];
    assign layer2_outputs[295] = ~(layer1_outputs[742]) | (layer1_outputs[4969]);
    assign layer2_outputs[296] = layer1_outputs[1848];
    assign layer2_outputs[297] = (layer1_outputs[1419]) & ~(layer1_outputs[4078]);
    assign layer2_outputs[298] = layer1_outputs[1601];
    assign layer2_outputs[299] = ~((layer1_outputs[344]) | (layer1_outputs[9]));
    assign layer2_outputs[300] = layer1_outputs[2614];
    assign layer2_outputs[301] = ~(layer1_outputs[1243]);
    assign layer2_outputs[302] = layer1_outputs[962];
    assign layer2_outputs[303] = (layer1_outputs[40]) | (layer1_outputs[878]);
    assign layer2_outputs[304] = (layer1_outputs[217]) | (layer1_outputs[2947]);
    assign layer2_outputs[305] = 1'b0;
    assign layer2_outputs[306] = ~((layer1_outputs[1836]) & (layer1_outputs[1606]));
    assign layer2_outputs[307] = ~(layer1_outputs[2785]);
    assign layer2_outputs[308] = layer1_outputs[2212];
    assign layer2_outputs[309] = 1'b0;
    assign layer2_outputs[310] = ~(layer1_outputs[366]) | (layer1_outputs[4917]);
    assign layer2_outputs[311] = ~(layer1_outputs[2701]);
    assign layer2_outputs[312] = (layer1_outputs[3450]) | (layer1_outputs[3547]);
    assign layer2_outputs[313] = ~(layer1_outputs[1706]) | (layer1_outputs[2636]);
    assign layer2_outputs[314] = 1'b0;
    assign layer2_outputs[315] = (layer1_outputs[1801]) ^ (layer1_outputs[1957]);
    assign layer2_outputs[316] = 1'b1;
    assign layer2_outputs[317] = (layer1_outputs[483]) | (layer1_outputs[1910]);
    assign layer2_outputs[318] = ~(layer1_outputs[4561]);
    assign layer2_outputs[319] = ~((layer1_outputs[2178]) | (layer1_outputs[1036]));
    assign layer2_outputs[320] = (layer1_outputs[4644]) | (layer1_outputs[890]);
    assign layer2_outputs[321] = 1'b1;
    assign layer2_outputs[322] = ~(layer1_outputs[551]) | (layer1_outputs[3709]);
    assign layer2_outputs[323] = 1'b1;
    assign layer2_outputs[324] = ~((layer1_outputs[1235]) | (layer1_outputs[2507]));
    assign layer2_outputs[325] = ~(layer1_outputs[4081]);
    assign layer2_outputs[326] = layer1_outputs[3372];
    assign layer2_outputs[327] = (layer1_outputs[1302]) & ~(layer1_outputs[1539]);
    assign layer2_outputs[328] = ~(layer1_outputs[4752]);
    assign layer2_outputs[329] = ~(layer1_outputs[4930]) | (layer1_outputs[2304]);
    assign layer2_outputs[330] = ~((layer1_outputs[887]) | (layer1_outputs[3232]));
    assign layer2_outputs[331] = layer1_outputs[4195];
    assign layer2_outputs[332] = layer1_outputs[2390];
    assign layer2_outputs[333] = (layer1_outputs[832]) | (layer1_outputs[3855]);
    assign layer2_outputs[334] = ~(layer1_outputs[841]) | (layer1_outputs[1121]);
    assign layer2_outputs[335] = (layer1_outputs[1739]) | (layer1_outputs[2879]);
    assign layer2_outputs[336] = ~((layer1_outputs[1717]) | (layer1_outputs[883]));
    assign layer2_outputs[337] = ~(layer1_outputs[4916]) | (layer1_outputs[3309]);
    assign layer2_outputs[338] = ~(layer1_outputs[3338]);
    assign layer2_outputs[339] = layer1_outputs[585];
    assign layer2_outputs[340] = layer1_outputs[4257];
    assign layer2_outputs[341] = ~(layer1_outputs[1353]) | (layer1_outputs[3795]);
    assign layer2_outputs[342] = layer1_outputs[4868];
    assign layer2_outputs[343] = ~(layer1_outputs[3691]) | (layer1_outputs[1027]);
    assign layer2_outputs[344] = ~((layer1_outputs[4681]) | (layer1_outputs[1058]));
    assign layer2_outputs[345] = (layer1_outputs[3242]) & ~(layer1_outputs[3335]);
    assign layer2_outputs[346] = layer1_outputs[3029];
    assign layer2_outputs[347] = ~(layer1_outputs[3896]) | (layer1_outputs[2630]);
    assign layer2_outputs[348] = ~((layer1_outputs[1757]) | (layer1_outputs[478]));
    assign layer2_outputs[349] = 1'b0;
    assign layer2_outputs[350] = ~((layer1_outputs[1535]) & (layer1_outputs[2309]));
    assign layer2_outputs[351] = ~((layer1_outputs[1858]) & (layer1_outputs[459]));
    assign layer2_outputs[352] = ~((layer1_outputs[3609]) ^ (layer1_outputs[958]));
    assign layer2_outputs[353] = (layer1_outputs[1284]) & ~(layer1_outputs[3496]);
    assign layer2_outputs[354] = ~(layer1_outputs[3298]);
    assign layer2_outputs[355] = ~((layer1_outputs[1868]) | (layer1_outputs[2766]));
    assign layer2_outputs[356] = ~(layer1_outputs[3868]) | (layer1_outputs[4412]);
    assign layer2_outputs[357] = (layer1_outputs[3211]) & ~(layer1_outputs[1795]);
    assign layer2_outputs[358] = 1'b1;
    assign layer2_outputs[359] = (layer1_outputs[3229]) & (layer1_outputs[4778]);
    assign layer2_outputs[360] = ~((layer1_outputs[4256]) | (layer1_outputs[416]));
    assign layer2_outputs[361] = ~((layer1_outputs[2391]) & (layer1_outputs[1901]));
    assign layer2_outputs[362] = layer1_outputs[858];
    assign layer2_outputs[363] = layer1_outputs[3495];
    assign layer2_outputs[364] = ~((layer1_outputs[5110]) & (layer1_outputs[3174]));
    assign layer2_outputs[365] = ~(layer1_outputs[3696]);
    assign layer2_outputs[366] = layer1_outputs[2489];
    assign layer2_outputs[367] = ~((layer1_outputs[2076]) & (layer1_outputs[4611]));
    assign layer2_outputs[368] = ~(layer1_outputs[4436]);
    assign layer2_outputs[369] = (layer1_outputs[358]) | (layer1_outputs[873]);
    assign layer2_outputs[370] = ~(layer1_outputs[1964]);
    assign layer2_outputs[371] = 1'b0;
    assign layer2_outputs[372] = ~(layer1_outputs[241]);
    assign layer2_outputs[373] = 1'b0;
    assign layer2_outputs[374] = 1'b0;
    assign layer2_outputs[375] = ~(layer1_outputs[3791]) | (layer1_outputs[445]);
    assign layer2_outputs[376] = ~(layer1_outputs[1837]) | (layer1_outputs[1967]);
    assign layer2_outputs[377] = ~((layer1_outputs[286]) | (layer1_outputs[2585]));
    assign layer2_outputs[378] = ~(layer1_outputs[205]);
    assign layer2_outputs[379] = (layer1_outputs[2531]) & ~(layer1_outputs[4196]);
    assign layer2_outputs[380] = 1'b0;
    assign layer2_outputs[381] = 1'b0;
    assign layer2_outputs[382] = ~((layer1_outputs[1285]) | (layer1_outputs[3927]));
    assign layer2_outputs[383] = layer1_outputs[4877];
    assign layer2_outputs[384] = layer1_outputs[698];
    assign layer2_outputs[385] = layer1_outputs[3494];
    assign layer2_outputs[386] = layer1_outputs[1123];
    assign layer2_outputs[387] = layer1_outputs[2493];
    assign layer2_outputs[388] = ~((layer1_outputs[4765]) & (layer1_outputs[2275]));
    assign layer2_outputs[389] = ~(layer1_outputs[917]) | (layer1_outputs[905]);
    assign layer2_outputs[390] = layer1_outputs[1772];
    assign layer2_outputs[391] = (layer1_outputs[1258]) & ~(layer1_outputs[2930]);
    assign layer2_outputs[392] = (layer1_outputs[2239]) ^ (layer1_outputs[5085]);
    assign layer2_outputs[393] = 1'b0;
    assign layer2_outputs[394] = ~(layer1_outputs[3721]);
    assign layer2_outputs[395] = ~(layer1_outputs[4594]) | (layer1_outputs[3735]);
    assign layer2_outputs[396] = 1'b1;
    assign layer2_outputs[397] = ~(layer1_outputs[4312]) | (layer1_outputs[2346]);
    assign layer2_outputs[398] = ~(layer1_outputs[885]) | (layer1_outputs[1895]);
    assign layer2_outputs[399] = layer1_outputs[197];
    assign layer2_outputs[400] = ~(layer1_outputs[4525]);
    assign layer2_outputs[401] = ~((layer1_outputs[244]) & (layer1_outputs[2225]));
    assign layer2_outputs[402] = ~((layer1_outputs[4512]) | (layer1_outputs[1819]));
    assign layer2_outputs[403] = (layer1_outputs[3734]) & (layer1_outputs[1376]);
    assign layer2_outputs[404] = (layer1_outputs[1100]) ^ (layer1_outputs[1088]);
    assign layer2_outputs[405] = ~((layer1_outputs[211]) ^ (layer1_outputs[1231]));
    assign layer2_outputs[406] = layer1_outputs[3027];
    assign layer2_outputs[407] = 1'b1;
    assign layer2_outputs[408] = 1'b0;
    assign layer2_outputs[409] = ~(layer1_outputs[2122]) | (layer1_outputs[4229]);
    assign layer2_outputs[410] = ~(layer1_outputs[4159]) | (layer1_outputs[858]);
    assign layer2_outputs[411] = (layer1_outputs[4398]) | (layer1_outputs[486]);
    assign layer2_outputs[412] = (layer1_outputs[258]) & ~(layer1_outputs[1093]);
    assign layer2_outputs[413] = ~((layer1_outputs[214]) | (layer1_outputs[429]));
    assign layer2_outputs[414] = (layer1_outputs[2443]) & ~(layer1_outputs[1625]);
    assign layer2_outputs[415] = (layer1_outputs[1091]) & ~(layer1_outputs[2463]);
    assign layer2_outputs[416] = layer1_outputs[140];
    assign layer2_outputs[417] = (layer1_outputs[1708]) & ~(layer1_outputs[2057]);
    assign layer2_outputs[418] = ~(layer1_outputs[4798]);
    assign layer2_outputs[419] = ~(layer1_outputs[4746]);
    assign layer2_outputs[420] = ~(layer1_outputs[4679]) | (layer1_outputs[1072]);
    assign layer2_outputs[421] = ~(layer1_outputs[4415]);
    assign layer2_outputs[422] = layer1_outputs[4274];
    assign layer2_outputs[423] = ~(layer1_outputs[662]) | (layer1_outputs[1196]);
    assign layer2_outputs[424] = (layer1_outputs[3581]) & ~(layer1_outputs[2669]);
    assign layer2_outputs[425] = (layer1_outputs[4515]) & (layer1_outputs[5115]);
    assign layer2_outputs[426] = ~(layer1_outputs[3577]);
    assign layer2_outputs[427] = (layer1_outputs[2705]) ^ (layer1_outputs[2497]);
    assign layer2_outputs[428] = ~((layer1_outputs[679]) & (layer1_outputs[4755]));
    assign layer2_outputs[429] = ~(layer1_outputs[4220]);
    assign layer2_outputs[430] = ~(layer1_outputs[3159]);
    assign layer2_outputs[431] = layer1_outputs[4111];
    assign layer2_outputs[432] = layer1_outputs[4];
    assign layer2_outputs[433] = ~(layer1_outputs[646]) | (layer1_outputs[4518]);
    assign layer2_outputs[434] = ~(layer1_outputs[2966]);
    assign layer2_outputs[435] = (layer1_outputs[5008]) & (layer1_outputs[2292]);
    assign layer2_outputs[436] = ~((layer1_outputs[4437]) & (layer1_outputs[560]));
    assign layer2_outputs[437] = ~(layer1_outputs[1279]);
    assign layer2_outputs[438] = ~(layer1_outputs[2569]);
    assign layer2_outputs[439] = (layer1_outputs[2476]) & ~(layer1_outputs[4413]);
    assign layer2_outputs[440] = 1'b0;
    assign layer2_outputs[441] = ~(layer1_outputs[4000]) | (layer1_outputs[42]);
    assign layer2_outputs[442] = layer1_outputs[411];
    assign layer2_outputs[443] = 1'b0;
    assign layer2_outputs[444] = ~((layer1_outputs[1758]) | (layer1_outputs[4938]));
    assign layer2_outputs[445] = 1'b0;
    assign layer2_outputs[446] = ~(layer1_outputs[416]);
    assign layer2_outputs[447] = ~(layer1_outputs[2169]);
    assign layer2_outputs[448] = ~(layer1_outputs[3409]);
    assign layer2_outputs[449] = ~(layer1_outputs[449]);
    assign layer2_outputs[450] = ~(layer1_outputs[2659]);
    assign layer2_outputs[451] = ~((layer1_outputs[2330]) & (layer1_outputs[5113]));
    assign layer2_outputs[452] = layer1_outputs[4081];
    assign layer2_outputs[453] = ~(layer1_outputs[55]) | (layer1_outputs[3652]);
    assign layer2_outputs[454] = ~(layer1_outputs[2022]) | (layer1_outputs[3209]);
    assign layer2_outputs[455] = ~(layer1_outputs[3543]) | (layer1_outputs[37]);
    assign layer2_outputs[456] = (layer1_outputs[4036]) & (layer1_outputs[3488]);
    assign layer2_outputs[457] = ~(layer1_outputs[4120]);
    assign layer2_outputs[458] = (layer1_outputs[670]) & ~(layer1_outputs[3851]);
    assign layer2_outputs[459] = (layer1_outputs[4516]) & ~(layer1_outputs[3637]);
    assign layer2_outputs[460] = ~((layer1_outputs[1877]) & (layer1_outputs[4232]));
    assign layer2_outputs[461] = ~((layer1_outputs[3602]) & (layer1_outputs[2801]));
    assign layer2_outputs[462] = layer1_outputs[2351];
    assign layer2_outputs[463] = (layer1_outputs[2396]) & ~(layer1_outputs[4535]);
    assign layer2_outputs[464] = (layer1_outputs[1104]) & ~(layer1_outputs[223]);
    assign layer2_outputs[465] = layer1_outputs[3297];
    assign layer2_outputs[466] = layer1_outputs[756];
    assign layer2_outputs[467] = 1'b1;
    assign layer2_outputs[468] = ~((layer1_outputs[1421]) & (layer1_outputs[4952]));
    assign layer2_outputs[469] = ~(layer1_outputs[3935]);
    assign layer2_outputs[470] = (layer1_outputs[4363]) & ~(layer1_outputs[3021]);
    assign layer2_outputs[471] = (layer1_outputs[2430]) | (layer1_outputs[4915]);
    assign layer2_outputs[472] = (layer1_outputs[4959]) & ~(layer1_outputs[2629]);
    assign layer2_outputs[473] = (layer1_outputs[1050]) & ~(layer1_outputs[998]);
    assign layer2_outputs[474] = layer1_outputs[3881];
    assign layer2_outputs[475] = layer1_outputs[2784];
    assign layer2_outputs[476] = layer1_outputs[2119];
    assign layer2_outputs[477] = layer1_outputs[4870];
    assign layer2_outputs[478] = (layer1_outputs[2452]) & ~(layer1_outputs[2986]);
    assign layer2_outputs[479] = ~((layer1_outputs[5074]) & (layer1_outputs[1388]));
    assign layer2_outputs[480] = 1'b0;
    assign layer2_outputs[481] = ~(layer1_outputs[2707]) | (layer1_outputs[1418]);
    assign layer2_outputs[482] = 1'b1;
    assign layer2_outputs[483] = ~(layer1_outputs[2061]);
    assign layer2_outputs[484] = ~(layer1_outputs[331]) | (layer1_outputs[4056]);
    assign layer2_outputs[485] = (layer1_outputs[1507]) & ~(layer1_outputs[3016]);
    assign layer2_outputs[486] = ~(layer1_outputs[4275]);
    assign layer2_outputs[487] = ~((layer1_outputs[3375]) & (layer1_outputs[72]));
    assign layer2_outputs[488] = 1'b0;
    assign layer2_outputs[489] = (layer1_outputs[51]) | (layer1_outputs[1425]);
    assign layer2_outputs[490] = layer1_outputs[4189];
    assign layer2_outputs[491] = ~((layer1_outputs[3225]) | (layer1_outputs[4782]));
    assign layer2_outputs[492] = (layer1_outputs[816]) & ~(layer1_outputs[128]);
    assign layer2_outputs[493] = layer1_outputs[2951];
    assign layer2_outputs[494] = (layer1_outputs[922]) | (layer1_outputs[2947]);
    assign layer2_outputs[495] = (layer1_outputs[1525]) | (layer1_outputs[2116]);
    assign layer2_outputs[496] = 1'b0;
    assign layer2_outputs[497] = (layer1_outputs[3117]) & ~(layer1_outputs[3978]);
    assign layer2_outputs[498] = (layer1_outputs[1160]) & ~(layer1_outputs[1319]);
    assign layer2_outputs[499] = (layer1_outputs[696]) & (layer1_outputs[2244]);
    assign layer2_outputs[500] = (layer1_outputs[4585]) & ~(layer1_outputs[4107]);
    assign layer2_outputs[501] = (layer1_outputs[4708]) & ~(layer1_outputs[4179]);
    assign layer2_outputs[502] = (layer1_outputs[4466]) & (layer1_outputs[4470]);
    assign layer2_outputs[503] = (layer1_outputs[1577]) & ~(layer1_outputs[385]);
    assign layer2_outputs[504] = ~(layer1_outputs[1673]);
    assign layer2_outputs[505] = (layer1_outputs[4878]) | (layer1_outputs[881]);
    assign layer2_outputs[506] = ~((layer1_outputs[5045]) & (layer1_outputs[2570]));
    assign layer2_outputs[507] = ~(layer1_outputs[4181]);
    assign layer2_outputs[508] = (layer1_outputs[5026]) & ~(layer1_outputs[872]);
    assign layer2_outputs[509] = 1'b0;
    assign layer2_outputs[510] = (layer1_outputs[4753]) & ~(layer1_outputs[1834]);
    assign layer2_outputs[511] = ~((layer1_outputs[4339]) & (layer1_outputs[1283]));
    assign layer2_outputs[512] = (layer1_outputs[1558]) & ~(layer1_outputs[2037]);
    assign layer2_outputs[513] = (layer1_outputs[1413]) & ~(layer1_outputs[3761]);
    assign layer2_outputs[514] = ~(layer1_outputs[99]);
    assign layer2_outputs[515] = 1'b1;
    assign layer2_outputs[516] = ~((layer1_outputs[1639]) & (layer1_outputs[4160]));
    assign layer2_outputs[517] = ~(layer1_outputs[3123]);
    assign layer2_outputs[518] = ~(layer1_outputs[5053]);
    assign layer2_outputs[519] = (layer1_outputs[82]) & ~(layer1_outputs[4370]);
    assign layer2_outputs[520] = (layer1_outputs[2209]) & (layer1_outputs[48]);
    assign layer2_outputs[521] = (layer1_outputs[4026]) | (layer1_outputs[3101]);
    assign layer2_outputs[522] = 1'b0;
    assign layer2_outputs[523] = (layer1_outputs[2128]) & ~(layer1_outputs[1358]);
    assign layer2_outputs[524] = ~(layer1_outputs[38]);
    assign layer2_outputs[525] = layer1_outputs[5000];
    assign layer2_outputs[526] = ~((layer1_outputs[2091]) & (layer1_outputs[1842]));
    assign layer2_outputs[527] = layer1_outputs[3663];
    assign layer2_outputs[528] = ~((layer1_outputs[2202]) | (layer1_outputs[2249]));
    assign layer2_outputs[529] = 1'b0;
    assign layer2_outputs[530] = 1'b0;
    assign layer2_outputs[531] = ~(layer1_outputs[676]);
    assign layer2_outputs[532] = ~(layer1_outputs[2495]);
    assign layer2_outputs[533] = ~(layer1_outputs[4172]);
    assign layer2_outputs[534] = 1'b0;
    assign layer2_outputs[535] = (layer1_outputs[3162]) & ~(layer1_outputs[922]);
    assign layer2_outputs[536] = ~(layer1_outputs[842]);
    assign layer2_outputs[537] = (layer1_outputs[1319]) & ~(layer1_outputs[3307]);
    assign layer2_outputs[538] = (layer1_outputs[1704]) | (layer1_outputs[4235]);
    assign layer2_outputs[539] = ~(layer1_outputs[2725]) | (layer1_outputs[2079]);
    assign layer2_outputs[540] = ~(layer1_outputs[1643]) | (layer1_outputs[4793]);
    assign layer2_outputs[541] = ~((layer1_outputs[2349]) & (layer1_outputs[4941]));
    assign layer2_outputs[542] = layer1_outputs[4764];
    assign layer2_outputs[543] = ~(layer1_outputs[1128]);
    assign layer2_outputs[544] = ~((layer1_outputs[3574]) | (layer1_outputs[3609]));
    assign layer2_outputs[545] = 1'b0;
    assign layer2_outputs[546] = layer1_outputs[2339];
    assign layer2_outputs[547] = (layer1_outputs[985]) | (layer1_outputs[3499]);
    assign layer2_outputs[548] = (layer1_outputs[3572]) & ~(layer1_outputs[2062]);
    assign layer2_outputs[549] = ~((layer1_outputs[4622]) ^ (layer1_outputs[1701]));
    assign layer2_outputs[550] = layer1_outputs[2595];
    assign layer2_outputs[551] = ~(layer1_outputs[1479]);
    assign layer2_outputs[552] = ~(layer1_outputs[839]);
    assign layer2_outputs[553] = (layer1_outputs[1017]) & ~(layer1_outputs[4884]);
    assign layer2_outputs[554] = layer1_outputs[2715];
    assign layer2_outputs[555] = layer1_outputs[1389];
    assign layer2_outputs[556] = ~((layer1_outputs[3387]) & (layer1_outputs[4484]));
    assign layer2_outputs[557] = ~((layer1_outputs[426]) | (layer1_outputs[591]));
    assign layer2_outputs[558] = ~(layer1_outputs[2059]);
    assign layer2_outputs[559] = (layer1_outputs[1489]) | (layer1_outputs[4180]);
    assign layer2_outputs[560] = ~(layer1_outputs[936]) | (layer1_outputs[2208]);
    assign layer2_outputs[561] = (layer1_outputs[4571]) & ~(layer1_outputs[3696]);
    assign layer2_outputs[562] = layer1_outputs[2276];
    assign layer2_outputs[563] = 1'b1;
    assign layer2_outputs[564] = layer1_outputs[4197];
    assign layer2_outputs[565] = ~((layer1_outputs[1576]) | (layer1_outputs[3044]));
    assign layer2_outputs[566] = ~((layer1_outputs[4798]) | (layer1_outputs[1731]));
    assign layer2_outputs[567] = ~((layer1_outputs[180]) ^ (layer1_outputs[670]));
    assign layer2_outputs[568] = ~(layer1_outputs[1146]) | (layer1_outputs[381]);
    assign layer2_outputs[569] = layer1_outputs[882];
    assign layer2_outputs[570] = ~(layer1_outputs[1848]);
    assign layer2_outputs[571] = ~(layer1_outputs[824]);
    assign layer2_outputs[572] = 1'b1;
    assign layer2_outputs[573] = (layer1_outputs[4714]) & (layer1_outputs[3214]);
    assign layer2_outputs[574] = ~((layer1_outputs[680]) & (layer1_outputs[948]));
    assign layer2_outputs[575] = ~(layer1_outputs[1549]);
    assign layer2_outputs[576] = ~((layer1_outputs[2635]) & (layer1_outputs[4022]));
    assign layer2_outputs[577] = (layer1_outputs[2014]) & ~(layer1_outputs[877]);
    assign layer2_outputs[578] = ~(layer1_outputs[4002]);
    assign layer2_outputs[579] = ~(layer1_outputs[2115]) | (layer1_outputs[3278]);
    assign layer2_outputs[580] = ~(layer1_outputs[3068]) | (layer1_outputs[2681]);
    assign layer2_outputs[581] = (layer1_outputs[3987]) & ~(layer1_outputs[3995]);
    assign layer2_outputs[582] = ~((layer1_outputs[1279]) & (layer1_outputs[2044]));
    assign layer2_outputs[583] = (layer1_outputs[3370]) | (layer1_outputs[2180]);
    assign layer2_outputs[584] = ~(layer1_outputs[1310]);
    assign layer2_outputs[585] = ~((layer1_outputs[5037]) & (layer1_outputs[57]));
    assign layer2_outputs[586] = ~((layer1_outputs[1893]) | (layer1_outputs[105]));
    assign layer2_outputs[587] = (layer1_outputs[3207]) & ~(layer1_outputs[1260]);
    assign layer2_outputs[588] = ~(layer1_outputs[2388]);
    assign layer2_outputs[589] = ~((layer1_outputs[210]) ^ (layer1_outputs[3118]));
    assign layer2_outputs[590] = ~((layer1_outputs[1857]) ^ (layer1_outputs[1929]));
    assign layer2_outputs[591] = (layer1_outputs[2511]) & (layer1_outputs[1373]);
    assign layer2_outputs[592] = (layer1_outputs[421]) ^ (layer1_outputs[3243]);
    assign layer2_outputs[593] = 1'b1;
    assign layer2_outputs[594] = ~(layer1_outputs[1786]);
    assign layer2_outputs[595] = ~((layer1_outputs[2421]) | (layer1_outputs[3986]));
    assign layer2_outputs[596] = ~((layer1_outputs[1195]) | (layer1_outputs[3408]));
    assign layer2_outputs[597] = (layer1_outputs[3426]) & (layer1_outputs[2249]);
    assign layer2_outputs[598] = (layer1_outputs[3234]) ^ (layer1_outputs[3810]);
    assign layer2_outputs[599] = ~(layer1_outputs[1467]) | (layer1_outputs[2757]);
    assign layer2_outputs[600] = ~(layer1_outputs[4976]);
    assign layer2_outputs[601] = (layer1_outputs[3173]) & ~(layer1_outputs[4622]);
    assign layer2_outputs[602] = (layer1_outputs[509]) & ~(layer1_outputs[4332]);
    assign layer2_outputs[603] = ~(layer1_outputs[2060]);
    assign layer2_outputs[604] = (layer1_outputs[1179]) & ~(layer1_outputs[4405]);
    assign layer2_outputs[605] = 1'b1;
    assign layer2_outputs[606] = 1'b0;
    assign layer2_outputs[607] = layer1_outputs[2154];
    assign layer2_outputs[608] = layer1_outputs[540];
    assign layer2_outputs[609] = ~(layer1_outputs[639]);
    assign layer2_outputs[610] = (layer1_outputs[919]) | (layer1_outputs[1087]);
    assign layer2_outputs[611] = ~(layer1_outputs[3891]);
    assign layer2_outputs[612] = 1'b0;
    assign layer2_outputs[613] = ~((layer1_outputs[1835]) ^ (layer1_outputs[4168]));
    assign layer2_outputs[614] = (layer1_outputs[2218]) & ~(layer1_outputs[2395]);
    assign layer2_outputs[615] = (layer1_outputs[3136]) & (layer1_outputs[1418]);
    assign layer2_outputs[616] = (layer1_outputs[2106]) & (layer1_outputs[268]);
    assign layer2_outputs[617] = (layer1_outputs[3988]) & ~(layer1_outputs[4214]);
    assign layer2_outputs[618] = (layer1_outputs[2136]) | (layer1_outputs[988]);
    assign layer2_outputs[619] = layer1_outputs[1215];
    assign layer2_outputs[620] = layer1_outputs[218];
    assign layer2_outputs[621] = (layer1_outputs[652]) & ~(layer1_outputs[1837]);
    assign layer2_outputs[622] = ~(layer1_outputs[1767]) | (layer1_outputs[600]);
    assign layer2_outputs[623] = layer1_outputs[2834];
    assign layer2_outputs[624] = ~(layer1_outputs[2888]);
    assign layer2_outputs[625] = layer1_outputs[200];
    assign layer2_outputs[626] = layer1_outputs[4625];
    assign layer2_outputs[627] = layer1_outputs[923];
    assign layer2_outputs[628] = ~((layer1_outputs[3874]) | (layer1_outputs[4641]));
    assign layer2_outputs[629] = ~(layer1_outputs[1457]);
    assign layer2_outputs[630] = layer1_outputs[2799];
    assign layer2_outputs[631] = layer1_outputs[3452];
    assign layer2_outputs[632] = ~(layer1_outputs[835]);
    assign layer2_outputs[633] = 1'b0;
    assign layer2_outputs[634] = 1'b1;
    assign layer2_outputs[635] = (layer1_outputs[498]) & ~(layer1_outputs[3012]);
    assign layer2_outputs[636] = (layer1_outputs[3729]) | (layer1_outputs[1204]);
    assign layer2_outputs[637] = ~((layer1_outputs[342]) & (layer1_outputs[4222]));
    assign layer2_outputs[638] = ~((layer1_outputs[413]) & (layer1_outputs[2222]));
    assign layer2_outputs[639] = ~(layer1_outputs[1783]) | (layer1_outputs[1335]);
    assign layer2_outputs[640] = 1'b0;
    assign layer2_outputs[641] = layer1_outputs[382];
    assign layer2_outputs[642] = ~((layer1_outputs[2051]) ^ (layer1_outputs[4795]));
    assign layer2_outputs[643] = ~((layer1_outputs[1641]) | (layer1_outputs[1436]));
    assign layer2_outputs[644] = (layer1_outputs[4349]) | (layer1_outputs[2042]);
    assign layer2_outputs[645] = ~(layer1_outputs[4153]) | (layer1_outputs[3749]);
    assign layer2_outputs[646] = ~(layer1_outputs[2108]);
    assign layer2_outputs[647] = (layer1_outputs[4560]) & ~(layer1_outputs[1191]);
    assign layer2_outputs[648] = layer1_outputs[4496];
    assign layer2_outputs[649] = (layer1_outputs[4147]) & ~(layer1_outputs[2435]);
    assign layer2_outputs[650] = ~(layer1_outputs[4031]);
    assign layer2_outputs[651] = ~((layer1_outputs[4336]) ^ (layer1_outputs[1384]));
    assign layer2_outputs[652] = ~(layer1_outputs[1136]) | (layer1_outputs[5103]);
    assign layer2_outputs[653] = layer1_outputs[1294];
    assign layer2_outputs[654] = ~(layer1_outputs[4708]);
    assign layer2_outputs[655] = 1'b1;
    assign layer2_outputs[656] = ~((layer1_outputs[2180]) & (layer1_outputs[1504]));
    assign layer2_outputs[657] = ~(layer1_outputs[3820]);
    assign layer2_outputs[658] = 1'b1;
    assign layer2_outputs[659] = 1'b0;
    assign layer2_outputs[660] = (layer1_outputs[4128]) & ~(layer1_outputs[2061]);
    assign layer2_outputs[661] = 1'b1;
    assign layer2_outputs[662] = ~(layer1_outputs[77]);
    assign layer2_outputs[663] = (layer1_outputs[3859]) & ~(layer1_outputs[2618]);
    assign layer2_outputs[664] = ~((layer1_outputs[4548]) ^ (layer1_outputs[4647]));
    assign layer2_outputs[665] = (layer1_outputs[3738]) & ~(layer1_outputs[1307]);
    assign layer2_outputs[666] = (layer1_outputs[4071]) | (layer1_outputs[4109]);
    assign layer2_outputs[667] = ~(layer1_outputs[3267]) | (layer1_outputs[4512]);
    assign layer2_outputs[668] = 1'b1;
    assign layer2_outputs[669] = 1'b0;
    assign layer2_outputs[670] = (layer1_outputs[1553]) & ~(layer1_outputs[593]);
    assign layer2_outputs[671] = layer1_outputs[3198];
    assign layer2_outputs[672] = 1'b1;
    assign layer2_outputs[673] = (layer1_outputs[1533]) & ~(layer1_outputs[2266]);
    assign layer2_outputs[674] = (layer1_outputs[3149]) & (layer1_outputs[1773]);
    assign layer2_outputs[675] = 1'b0;
    assign layer2_outputs[676] = (layer1_outputs[2109]) & ~(layer1_outputs[1111]);
    assign layer2_outputs[677] = (layer1_outputs[2005]) | (layer1_outputs[3938]);
    assign layer2_outputs[678] = 1'b0;
    assign layer2_outputs[679] = ~(layer1_outputs[2576]) | (layer1_outputs[2568]);
    assign layer2_outputs[680] = 1'b0;
    assign layer2_outputs[681] = layer1_outputs[4954];
    assign layer2_outputs[682] = ~((layer1_outputs[2679]) & (layer1_outputs[4277]));
    assign layer2_outputs[683] = (layer1_outputs[4705]) & (layer1_outputs[1556]);
    assign layer2_outputs[684] = ~(layer1_outputs[948]);
    assign layer2_outputs[685] = 1'b0;
    assign layer2_outputs[686] = layer1_outputs[1252];
    assign layer2_outputs[687] = ~(layer1_outputs[4579]) | (layer1_outputs[3660]);
    assign layer2_outputs[688] = layer1_outputs[829];
    assign layer2_outputs[689] = ~(layer1_outputs[1528]);
    assign layer2_outputs[690] = layer1_outputs[1124];
    assign layer2_outputs[691] = ~((layer1_outputs[3934]) ^ (layer1_outputs[2674]));
    assign layer2_outputs[692] = layer1_outputs[4021];
    assign layer2_outputs[693] = ~(layer1_outputs[1574]) | (layer1_outputs[4644]);
    assign layer2_outputs[694] = (layer1_outputs[2339]) & ~(layer1_outputs[4128]);
    assign layer2_outputs[695] = ~(layer1_outputs[176]) | (layer1_outputs[2614]);
    assign layer2_outputs[696] = ~(layer1_outputs[2225]) | (layer1_outputs[2946]);
    assign layer2_outputs[697] = ~(layer1_outputs[3803]);
    assign layer2_outputs[698] = 1'b0;
    assign layer2_outputs[699] = ~(layer1_outputs[666]) | (layer1_outputs[226]);
    assign layer2_outputs[700] = 1'b0;
    assign layer2_outputs[701] = layer1_outputs[4595];
    assign layer2_outputs[702] = ~((layer1_outputs[124]) | (layer1_outputs[3376]));
    assign layer2_outputs[703] = 1'b1;
    assign layer2_outputs[704] = (layer1_outputs[572]) & (layer1_outputs[3007]);
    assign layer2_outputs[705] = (layer1_outputs[4480]) & ~(layer1_outputs[4453]);
    assign layer2_outputs[706] = 1'b0;
    assign layer2_outputs[707] = layer1_outputs[4334];
    assign layer2_outputs[708] = ~((layer1_outputs[4491]) & (layer1_outputs[3566]));
    assign layer2_outputs[709] = ~((layer1_outputs[2532]) | (layer1_outputs[1854]));
    assign layer2_outputs[710] = ~(layer1_outputs[5054]);
    assign layer2_outputs[711] = layer1_outputs[4317];
    assign layer2_outputs[712] = ~(layer1_outputs[3289]) | (layer1_outputs[1863]);
    assign layer2_outputs[713] = (layer1_outputs[685]) & (layer1_outputs[4922]);
    assign layer2_outputs[714] = layer1_outputs[1164];
    assign layer2_outputs[715] = ~((layer1_outputs[4620]) & (layer1_outputs[3059]));
    assign layer2_outputs[716] = ~((layer1_outputs[4781]) & (layer1_outputs[4408]));
    assign layer2_outputs[717] = 1'b0;
    assign layer2_outputs[718] = 1'b0;
    assign layer2_outputs[719] = layer1_outputs[4408];
    assign layer2_outputs[720] = layer1_outputs[907];
    assign layer2_outputs[721] = layer1_outputs[65];
    assign layer2_outputs[722] = layer1_outputs[1412];
    assign layer2_outputs[723] = ~(layer1_outputs[397]);
    assign layer2_outputs[724] = (layer1_outputs[3434]) & ~(layer1_outputs[86]);
    assign layer2_outputs[725] = layer1_outputs[4657];
    assign layer2_outputs[726] = ~((layer1_outputs[3534]) & (layer1_outputs[1557]));
    assign layer2_outputs[727] = layer1_outputs[2440];
    assign layer2_outputs[728] = ~(layer1_outputs[4741]) | (layer1_outputs[158]);
    assign layer2_outputs[729] = 1'b1;
    assign layer2_outputs[730] = (layer1_outputs[2792]) | (layer1_outputs[1276]);
    assign layer2_outputs[731] = 1'b1;
    assign layer2_outputs[732] = (layer1_outputs[2501]) & ~(layer1_outputs[3745]);
    assign layer2_outputs[733] = ~(layer1_outputs[4794]) | (layer1_outputs[4394]);
    assign layer2_outputs[734] = layer1_outputs[329];
    assign layer2_outputs[735] = layer1_outputs[2333];
    assign layer2_outputs[736] = 1'b1;
    assign layer2_outputs[737] = ~(layer1_outputs[1421]);
    assign layer2_outputs[738] = ~((layer1_outputs[3900]) | (layer1_outputs[1386]));
    assign layer2_outputs[739] = (layer1_outputs[1735]) | (layer1_outputs[382]);
    assign layer2_outputs[740] = layer1_outputs[3774];
    assign layer2_outputs[741] = 1'b0;
    assign layer2_outputs[742] = ~(layer1_outputs[480]);
    assign layer2_outputs[743] = 1'b0;
    assign layer2_outputs[744] = ~(layer1_outputs[669]);
    assign layer2_outputs[745] = ~((layer1_outputs[4838]) | (layer1_outputs[718]));
    assign layer2_outputs[746] = ~((layer1_outputs[2230]) & (layer1_outputs[4425]));
    assign layer2_outputs[747] = ~(layer1_outputs[477]) | (layer1_outputs[1369]);
    assign layer2_outputs[748] = ~(layer1_outputs[4400]) | (layer1_outputs[425]);
    assign layer2_outputs[749] = ~((layer1_outputs[1918]) & (layer1_outputs[1637]));
    assign layer2_outputs[750] = (layer1_outputs[2509]) | (layer1_outputs[3754]);
    assign layer2_outputs[751] = layer1_outputs[1649];
    assign layer2_outputs[752] = ~((layer1_outputs[1566]) | (layer1_outputs[138]));
    assign layer2_outputs[753] = 1'b0;
    assign layer2_outputs[754] = ~(layer1_outputs[3308]);
    assign layer2_outputs[755] = ~(layer1_outputs[3435]);
    assign layer2_outputs[756] = layer1_outputs[2003];
    assign layer2_outputs[757] = ~((layer1_outputs[995]) | (layer1_outputs[2453]));
    assign layer2_outputs[758] = ~(layer1_outputs[1535]) | (layer1_outputs[1452]);
    assign layer2_outputs[759] = ~((layer1_outputs[1689]) ^ (layer1_outputs[469]));
    assign layer2_outputs[760] = (layer1_outputs[4316]) | (layer1_outputs[2660]);
    assign layer2_outputs[761] = ~(layer1_outputs[3526]);
    assign layer2_outputs[762] = layer1_outputs[367];
    assign layer2_outputs[763] = layer1_outputs[3545];
    assign layer2_outputs[764] = layer1_outputs[1628];
    assign layer2_outputs[765] = layer1_outputs[2937];
    assign layer2_outputs[766] = ~(layer1_outputs[1708]) | (layer1_outputs[618]);
    assign layer2_outputs[767] = ~(layer1_outputs[588]) | (layer1_outputs[4018]);
    assign layer2_outputs[768] = ~((layer1_outputs[2341]) & (layer1_outputs[4458]));
    assign layer2_outputs[769] = (layer1_outputs[1172]) & (layer1_outputs[4242]);
    assign layer2_outputs[770] = ~(layer1_outputs[4630]) | (layer1_outputs[4989]);
    assign layer2_outputs[771] = layer1_outputs[3035];
    assign layer2_outputs[772] = 1'b0;
    assign layer2_outputs[773] = (layer1_outputs[609]) & ~(layer1_outputs[2892]);
    assign layer2_outputs[774] = ~((layer1_outputs[5060]) & (layer1_outputs[4695]));
    assign layer2_outputs[775] = 1'b1;
    assign layer2_outputs[776] = ~(layer1_outputs[4666]) | (layer1_outputs[936]);
    assign layer2_outputs[777] = layer1_outputs[978];
    assign layer2_outputs[778] = (layer1_outputs[849]) & ~(layer1_outputs[3406]);
    assign layer2_outputs[779] = layer1_outputs[1096];
    assign layer2_outputs[780] = ~((layer1_outputs[4073]) & (layer1_outputs[496]));
    assign layer2_outputs[781] = ~(layer1_outputs[2221]) | (layer1_outputs[4640]);
    assign layer2_outputs[782] = (layer1_outputs[959]) | (layer1_outputs[4770]);
    assign layer2_outputs[783] = layer1_outputs[2080];
    assign layer2_outputs[784] = ~(layer1_outputs[79]) | (layer1_outputs[4249]);
    assign layer2_outputs[785] = ~((layer1_outputs[5017]) | (layer1_outputs[4664]));
    assign layer2_outputs[786] = (layer1_outputs[2779]) ^ (layer1_outputs[869]);
    assign layer2_outputs[787] = layer1_outputs[3256];
    assign layer2_outputs[788] = ~((layer1_outputs[4334]) & (layer1_outputs[290]));
    assign layer2_outputs[789] = 1'b1;
    assign layer2_outputs[790] = layer1_outputs[148];
    assign layer2_outputs[791] = layer1_outputs[2124];
    assign layer2_outputs[792] = layer1_outputs[2411];
    assign layer2_outputs[793] = ~((layer1_outputs[2913]) ^ (layer1_outputs[5036]));
    assign layer2_outputs[794] = ~(layer1_outputs[4029]) | (layer1_outputs[3709]);
    assign layer2_outputs[795] = (layer1_outputs[2141]) & ~(layer1_outputs[4399]);
    assign layer2_outputs[796] = 1'b1;
    assign layer2_outputs[797] = (layer1_outputs[3649]) & (layer1_outputs[3663]);
    assign layer2_outputs[798] = 1'b1;
    assign layer2_outputs[799] = ~((layer1_outputs[4154]) | (layer1_outputs[3363]));
    assign layer2_outputs[800] = ~((layer1_outputs[3377]) | (layer1_outputs[1447]));
    assign layer2_outputs[801] = ~(layer1_outputs[4718]) | (layer1_outputs[1456]);
    assign layer2_outputs[802] = layer1_outputs[3510];
    assign layer2_outputs[803] = ~(layer1_outputs[171]);
    assign layer2_outputs[804] = 1'b0;
    assign layer2_outputs[805] = ~(layer1_outputs[7]) | (layer1_outputs[3567]);
    assign layer2_outputs[806] = ~(layer1_outputs[3651]);
    assign layer2_outputs[807] = ~((layer1_outputs[1561]) | (layer1_outputs[4337]));
    assign layer2_outputs[808] = (layer1_outputs[517]) | (layer1_outputs[3249]);
    assign layer2_outputs[809] = ~(layer1_outputs[4844]) | (layer1_outputs[4658]);
    assign layer2_outputs[810] = ~((layer1_outputs[832]) & (layer1_outputs[3499]));
    assign layer2_outputs[811] = (layer1_outputs[4857]) & (layer1_outputs[3740]);
    assign layer2_outputs[812] = (layer1_outputs[4826]) & ~(layer1_outputs[3140]);
    assign layer2_outputs[813] = layer1_outputs[2161];
    assign layer2_outputs[814] = (layer1_outputs[4533]) & (layer1_outputs[4936]);
    assign layer2_outputs[815] = 1'b1;
    assign layer2_outputs[816] = (layer1_outputs[3947]) & ~(layer1_outputs[2640]);
    assign layer2_outputs[817] = (layer1_outputs[4986]) & ~(layer1_outputs[3586]);
    assign layer2_outputs[818] = ~(layer1_outputs[3618]) | (layer1_outputs[315]);
    assign layer2_outputs[819] = 1'b1;
    assign layer2_outputs[820] = layer1_outputs[1695];
    assign layer2_outputs[821] = 1'b1;
    assign layer2_outputs[822] = ~(layer1_outputs[3385]);
    assign layer2_outputs[823] = ~((layer1_outputs[4090]) | (layer1_outputs[4262]));
    assign layer2_outputs[824] = ~((layer1_outputs[2364]) | (layer1_outputs[4959]));
    assign layer2_outputs[825] = 1'b1;
    assign layer2_outputs[826] = (layer1_outputs[266]) & ~(layer1_outputs[1272]);
    assign layer2_outputs[827] = ~((layer1_outputs[1364]) & (layer1_outputs[838]));
    assign layer2_outputs[828] = layer1_outputs[8];
    assign layer2_outputs[829] = ~(layer1_outputs[3705]);
    assign layer2_outputs[830] = layer1_outputs[4968];
    assign layer2_outputs[831] = ~(layer1_outputs[5089]);
    assign layer2_outputs[832] = layer1_outputs[1878];
    assign layer2_outputs[833] = ~(layer1_outputs[1349]);
    assign layer2_outputs[834] = ~(layer1_outputs[3240]);
    assign layer2_outputs[835] = ~(layer1_outputs[1316]) | (layer1_outputs[1323]);
    assign layer2_outputs[836] = ~(layer1_outputs[1884]);
    assign layer2_outputs[837] = layer1_outputs[687];
    assign layer2_outputs[838] = ~(layer1_outputs[63]) | (layer1_outputs[2289]);
    assign layer2_outputs[839] = (layer1_outputs[580]) & ~(layer1_outputs[994]);
    assign layer2_outputs[840] = ~(layer1_outputs[770]);
    assign layer2_outputs[841] = 1'b0;
    assign layer2_outputs[842] = ~((layer1_outputs[1031]) | (layer1_outputs[3864]));
    assign layer2_outputs[843] = layer1_outputs[4103];
    assign layer2_outputs[844] = 1'b1;
    assign layer2_outputs[845] = layer1_outputs[4834];
    assign layer2_outputs[846] = layer1_outputs[694];
    assign layer2_outputs[847] = 1'b0;
    assign layer2_outputs[848] = ~(layer1_outputs[904]);
    assign layer2_outputs[849] = (layer1_outputs[448]) & (layer1_outputs[1490]);
    assign layer2_outputs[850] = ~(layer1_outputs[579]);
    assign layer2_outputs[851] = (layer1_outputs[4709]) | (layer1_outputs[2182]);
    assign layer2_outputs[852] = ~(layer1_outputs[4568]) | (layer1_outputs[2986]);
    assign layer2_outputs[853] = layer1_outputs[3248];
    assign layer2_outputs[854] = ~((layer1_outputs[3374]) | (layer1_outputs[4712]));
    assign layer2_outputs[855] = ~(layer1_outputs[4017]);
    assign layer2_outputs[856] = (layer1_outputs[77]) | (layer1_outputs[2107]);
    assign layer2_outputs[857] = ~((layer1_outputs[5069]) | (layer1_outputs[1424]));
    assign layer2_outputs[858] = ~((layer1_outputs[4454]) & (layer1_outputs[4205]));
    assign layer2_outputs[859] = (layer1_outputs[4171]) | (layer1_outputs[1827]);
    assign layer2_outputs[860] = ~(layer1_outputs[3038]) | (layer1_outputs[4684]);
    assign layer2_outputs[861] = ~(layer1_outputs[5111]);
    assign layer2_outputs[862] = (layer1_outputs[1229]) & (layer1_outputs[1656]);
    assign layer2_outputs[863] = ~(layer1_outputs[2657]);
    assign layer2_outputs[864] = (layer1_outputs[3914]) & (layer1_outputs[4740]);
    assign layer2_outputs[865] = ~((layer1_outputs[190]) ^ (layer1_outputs[4156]));
    assign layer2_outputs[866] = layer1_outputs[4236];
    assign layer2_outputs[867] = layer1_outputs[4991];
    assign layer2_outputs[868] = ~((layer1_outputs[41]) | (layer1_outputs[4057]));
    assign layer2_outputs[869] = 1'b0;
    assign layer2_outputs[870] = layer1_outputs[2096];
    assign layer2_outputs[871] = (layer1_outputs[3814]) & ~(layer1_outputs[2098]);
    assign layer2_outputs[872] = ~(layer1_outputs[1803]) | (layer1_outputs[3305]);
    assign layer2_outputs[873] = (layer1_outputs[1159]) & ~(layer1_outputs[4499]);
    assign layer2_outputs[874] = (layer1_outputs[1355]) ^ (layer1_outputs[868]);
    assign layer2_outputs[875] = 1'b1;
    assign layer2_outputs[876] = 1'b1;
    assign layer2_outputs[877] = ~(layer1_outputs[3808]) | (layer1_outputs[434]);
    assign layer2_outputs[878] = (layer1_outputs[4373]) & ~(layer1_outputs[2687]);
    assign layer2_outputs[879] = (layer1_outputs[4524]) ^ (layer1_outputs[161]);
    assign layer2_outputs[880] = 1'b1;
    assign layer2_outputs[881] = ~((layer1_outputs[3473]) | (layer1_outputs[3106]));
    assign layer2_outputs[882] = ~(layer1_outputs[5011]);
    assign layer2_outputs[883] = ~(layer1_outputs[1511]);
    assign layer2_outputs[884] = 1'b0;
    assign layer2_outputs[885] = ~((layer1_outputs[5083]) | (layer1_outputs[2466]));
    assign layer2_outputs[886] = layer1_outputs[558];
    assign layer2_outputs[887] = ~(layer1_outputs[2401]) | (layer1_outputs[1784]);
    assign layer2_outputs[888] = 1'b0;
    assign layer2_outputs[889] = 1'b1;
    assign layer2_outputs[890] = (layer1_outputs[535]) & ~(layer1_outputs[5076]);
    assign layer2_outputs[891] = layer1_outputs[1149];
    assign layer2_outputs[892] = layer1_outputs[3591];
    assign layer2_outputs[893] = (layer1_outputs[3201]) & (layer1_outputs[2974]);
    assign layer2_outputs[894] = ~(layer1_outputs[3994]);
    assign layer2_outputs[895] = layer1_outputs[584];
    assign layer2_outputs[896] = ~(layer1_outputs[944]) | (layer1_outputs[4009]);
    assign layer2_outputs[897] = (layer1_outputs[2273]) | (layer1_outputs[1363]);
    assign layer2_outputs[898] = ~((layer1_outputs[3078]) | (layer1_outputs[467]));
    assign layer2_outputs[899] = ~((layer1_outputs[1344]) & (layer1_outputs[1651]));
    assign layer2_outputs[900] = (layer1_outputs[249]) & ~(layer1_outputs[1888]);
    assign layer2_outputs[901] = layer1_outputs[485];
    assign layer2_outputs[902] = (layer1_outputs[3666]) & (layer1_outputs[345]);
    assign layer2_outputs[903] = ~(layer1_outputs[4679]);
    assign layer2_outputs[904] = (layer1_outputs[328]) & ~(layer1_outputs[1062]);
    assign layer2_outputs[905] = ~(layer1_outputs[2446]) | (layer1_outputs[608]);
    assign layer2_outputs[906] = ~(layer1_outputs[2507]) | (layer1_outputs[4898]);
    assign layer2_outputs[907] = 1'b1;
    assign layer2_outputs[908] = 1'b1;
    assign layer2_outputs[909] = ~(layer1_outputs[1299]);
    assign layer2_outputs[910] = ~(layer1_outputs[1833]);
    assign layer2_outputs[911] = (layer1_outputs[677]) ^ (layer1_outputs[4184]);
    assign layer2_outputs[912] = ~(layer1_outputs[3498]);
    assign layer2_outputs[913] = (layer1_outputs[3484]) & ~(layer1_outputs[3254]);
    assign layer2_outputs[914] = ~((layer1_outputs[1500]) ^ (layer1_outputs[2125]));
    assign layer2_outputs[915] = (layer1_outputs[3574]) & ~(layer1_outputs[4557]);
    assign layer2_outputs[916] = layer1_outputs[786];
    assign layer2_outputs[917] = layer1_outputs[2385];
    assign layer2_outputs[918] = ~((layer1_outputs[330]) & (layer1_outputs[345]));
    assign layer2_outputs[919] = layer1_outputs[4673];
    assign layer2_outputs[920] = ~((layer1_outputs[3281]) ^ (layer1_outputs[3940]));
    assign layer2_outputs[921] = (layer1_outputs[276]) & ~(layer1_outputs[4402]);
    assign layer2_outputs[922] = ~(layer1_outputs[2430]);
    assign layer2_outputs[923] = (layer1_outputs[3497]) & ~(layer1_outputs[1920]);
    assign layer2_outputs[924] = ~((layer1_outputs[4377]) & (layer1_outputs[3161]));
    assign layer2_outputs[925] = (layer1_outputs[263]) & ~(layer1_outputs[4561]);
    assign layer2_outputs[926] = ~(layer1_outputs[1818]) | (layer1_outputs[2539]);
    assign layer2_outputs[927] = 1'b0;
    assign layer2_outputs[928] = (layer1_outputs[3415]) | (layer1_outputs[599]);
    assign layer2_outputs[929] = (layer1_outputs[1969]) & ~(layer1_outputs[615]);
    assign layer2_outputs[930] = (layer1_outputs[1754]) & (layer1_outputs[351]);
    assign layer2_outputs[931] = (layer1_outputs[886]) | (layer1_outputs[4536]);
    assign layer2_outputs[932] = layer1_outputs[1599];
    assign layer2_outputs[933] = ~((layer1_outputs[1272]) ^ (layer1_outputs[1732]));
    assign layer2_outputs[934] = ~(layer1_outputs[1170]) | (layer1_outputs[1998]);
    assign layer2_outputs[935] = layer1_outputs[1071];
    assign layer2_outputs[936] = layer1_outputs[2412];
    assign layer2_outputs[937] = ~(layer1_outputs[4446]) | (layer1_outputs[3542]);
    assign layer2_outputs[938] = ~(layer1_outputs[3228]);
    assign layer2_outputs[939] = 1'b0;
    assign layer2_outputs[940] = ~(layer1_outputs[1670]);
    assign layer2_outputs[941] = (layer1_outputs[2465]) & (layer1_outputs[2049]);
    assign layer2_outputs[942] = layer1_outputs[2194];
    assign layer2_outputs[943] = (layer1_outputs[4811]) & ~(layer1_outputs[244]);
    assign layer2_outputs[944] = layer1_outputs[1640];
    assign layer2_outputs[945] = layer1_outputs[938];
    assign layer2_outputs[946] = ~(layer1_outputs[3369]) | (layer1_outputs[1372]);
    assign layer2_outputs[947] = layer1_outputs[222];
    assign layer2_outputs[948] = ~(layer1_outputs[4489]) | (layer1_outputs[1753]);
    assign layer2_outputs[949] = ~((layer1_outputs[4927]) | (layer1_outputs[2962]));
    assign layer2_outputs[950] = ~(layer1_outputs[3502]);
    assign layer2_outputs[951] = (layer1_outputs[4932]) | (layer1_outputs[5065]);
    assign layer2_outputs[952] = ~(layer1_outputs[206]);
    assign layer2_outputs[953] = (layer1_outputs[1966]) & (layer1_outputs[1664]);
    assign layer2_outputs[954] = layer1_outputs[1054];
    assign layer2_outputs[955] = ~(layer1_outputs[364]) | (layer1_outputs[3360]);
    assign layer2_outputs[956] = (layer1_outputs[1473]) & ~(layer1_outputs[4216]);
    assign layer2_outputs[957] = ~(layer1_outputs[4764]) | (layer1_outputs[2735]);
    assign layer2_outputs[958] = layer1_outputs[3894];
    assign layer2_outputs[959] = ~((layer1_outputs[1603]) & (layer1_outputs[132]));
    assign layer2_outputs[960] = (layer1_outputs[25]) & ~(layer1_outputs[1718]);
    assign layer2_outputs[961] = 1'b1;
    assign layer2_outputs[962] = ~(layer1_outputs[2558]);
    assign layer2_outputs[963] = layer1_outputs[4650];
    assign layer2_outputs[964] = ~((layer1_outputs[1844]) ^ (layer1_outputs[1374]));
    assign layer2_outputs[965] = layer1_outputs[3502];
    assign layer2_outputs[966] = ~(layer1_outputs[4809]) | (layer1_outputs[1076]);
    assign layer2_outputs[967] = 1'b0;
    assign layer2_outputs[968] = (layer1_outputs[3588]) & ~(layer1_outputs[30]);
    assign layer2_outputs[969] = (layer1_outputs[4179]) & (layer1_outputs[4105]);
    assign layer2_outputs[970] = (layer1_outputs[1935]) & ~(layer1_outputs[701]);
    assign layer2_outputs[971] = 1'b0;
    assign layer2_outputs[972] = (layer1_outputs[2457]) & ~(layer1_outputs[4303]);
    assign layer2_outputs[973] = ~((layer1_outputs[259]) & (layer1_outputs[3719]));
    assign layer2_outputs[974] = (layer1_outputs[1163]) | (layer1_outputs[2283]);
    assign layer2_outputs[975] = (layer1_outputs[1895]) & ~(layer1_outputs[2638]);
    assign layer2_outputs[976] = ~(layer1_outputs[4359]) | (layer1_outputs[2157]);
    assign layer2_outputs[977] = ~(layer1_outputs[3134]) | (layer1_outputs[2948]);
    assign layer2_outputs[978] = (layer1_outputs[1952]) & (layer1_outputs[3498]);
    assign layer2_outputs[979] = ~(layer1_outputs[5062]);
    assign layer2_outputs[980] = ~(layer1_outputs[2052]) | (layer1_outputs[602]);
    assign layer2_outputs[981] = ~(layer1_outputs[2949]);
    assign layer2_outputs[982] = ~(layer1_outputs[3245]);
    assign layer2_outputs[983] = ~(layer1_outputs[1987]) | (layer1_outputs[3956]);
    assign layer2_outputs[984] = 1'b0;
    assign layer2_outputs[985] = ~((layer1_outputs[1404]) | (layer1_outputs[1247]));
    assign layer2_outputs[986] = (layer1_outputs[4183]) | (layer1_outputs[1800]);
    assign layer2_outputs[987] = ~(layer1_outputs[1362]);
    assign layer2_outputs[988] = (layer1_outputs[1181]) & ~(layer1_outputs[951]);
    assign layer2_outputs[989] = 1'b1;
    assign layer2_outputs[990] = 1'b0;
    assign layer2_outputs[991] = ~(layer1_outputs[1049]);
    assign layer2_outputs[992] = ~(layer1_outputs[5117]);
    assign layer2_outputs[993] = ~(layer1_outputs[2609]);
    assign layer2_outputs[994] = (layer1_outputs[4325]) & (layer1_outputs[2889]);
    assign layer2_outputs[995] = ~(layer1_outputs[2352]) | (layer1_outputs[795]);
    assign layer2_outputs[996] = (layer1_outputs[1440]) | (layer1_outputs[1903]);
    assign layer2_outputs[997] = ~(layer1_outputs[4111]) | (layer1_outputs[3025]);
    assign layer2_outputs[998] = ~(layer1_outputs[2850]);
    assign layer2_outputs[999] = 1'b1;
    assign layer2_outputs[1000] = ~(layer1_outputs[2004]);
    assign layer2_outputs[1001] = (layer1_outputs[3661]) | (layer1_outputs[3954]);
    assign layer2_outputs[1002] = ~((layer1_outputs[5064]) | (layer1_outputs[4323]));
    assign layer2_outputs[1003] = ~(layer1_outputs[2316]);
    assign layer2_outputs[1004] = layer1_outputs[4280];
    assign layer2_outputs[1005] = layer1_outputs[473];
    assign layer2_outputs[1006] = (layer1_outputs[2655]) ^ (layer1_outputs[2470]);
    assign layer2_outputs[1007] = (layer1_outputs[2546]) & ~(layer1_outputs[1028]);
    assign layer2_outputs[1008] = (layer1_outputs[16]) | (layer1_outputs[2978]);
    assign layer2_outputs[1009] = (layer1_outputs[4115]) & (layer1_outputs[3559]);
    assign layer2_outputs[1010] = ~(layer1_outputs[3270]);
    assign layer2_outputs[1011] = (layer1_outputs[3615]) & ~(layer1_outputs[4476]);
    assign layer2_outputs[1012] = ~(layer1_outputs[4211]) | (layer1_outputs[1093]);
    assign layer2_outputs[1013] = ~(layer1_outputs[1668]) | (layer1_outputs[2462]);
    assign layer2_outputs[1014] = 1'b1;
    assign layer2_outputs[1015] = ~((layer1_outputs[1228]) & (layer1_outputs[4247]));
    assign layer2_outputs[1016] = (layer1_outputs[2213]) & ~(layer1_outputs[2197]);
    assign layer2_outputs[1017] = 1'b1;
    assign layer2_outputs[1018] = layer1_outputs[816];
    assign layer2_outputs[1019] = 1'b1;
    assign layer2_outputs[1020] = layer1_outputs[333];
    assign layer2_outputs[1021] = ~(layer1_outputs[3266]) | (layer1_outputs[3466]);
    assign layer2_outputs[1022] = layer1_outputs[249];
    assign layer2_outputs[1023] = ~(layer1_outputs[4457]) | (layer1_outputs[3051]);
    assign layer2_outputs[1024] = (layer1_outputs[4864]) & ~(layer1_outputs[4079]);
    assign layer2_outputs[1025] = ~(layer1_outputs[941]);
    assign layer2_outputs[1026] = layer1_outputs[673];
    assign layer2_outputs[1027] = ~((layer1_outputs[814]) & (layer1_outputs[4150]));
    assign layer2_outputs[1028] = 1'b0;
    assign layer2_outputs[1029] = (layer1_outputs[4043]) & ~(layer1_outputs[1383]);
    assign layer2_outputs[1030] = ~(layer1_outputs[2647]) | (layer1_outputs[2823]);
    assign layer2_outputs[1031] = ~(layer1_outputs[3081]);
    assign layer2_outputs[1032] = ~(layer1_outputs[241]) | (layer1_outputs[2323]);
    assign layer2_outputs[1033] = ~(layer1_outputs[3687]);
    assign layer2_outputs[1034] = layer1_outputs[2876];
    assign layer2_outputs[1035] = ~(layer1_outputs[359]);
    assign layer2_outputs[1036] = ~(layer1_outputs[4937]);
    assign layer2_outputs[1037] = ~(layer1_outputs[760]) | (layer1_outputs[283]);
    assign layer2_outputs[1038] = (layer1_outputs[2481]) & ~(layer1_outputs[351]);
    assign layer2_outputs[1039] = 1'b1;
    assign layer2_outputs[1040] = ~((layer1_outputs[4459]) | (layer1_outputs[1980]));
    assign layer2_outputs[1041] = ~(layer1_outputs[5113]);
    assign layer2_outputs[1042] = ~((layer1_outputs[4058]) & (layer1_outputs[18]));
    assign layer2_outputs[1043] = ~(layer1_outputs[4794]);
    assign layer2_outputs[1044] = (layer1_outputs[1392]) & (layer1_outputs[2829]);
    assign layer2_outputs[1045] = ~((layer1_outputs[4411]) & (layer1_outputs[5]));
    assign layer2_outputs[1046] = ~(layer1_outputs[4070]);
    assign layer2_outputs[1047] = ~((layer1_outputs[2263]) | (layer1_outputs[470]));
    assign layer2_outputs[1048] = (layer1_outputs[761]) & (layer1_outputs[3070]);
    assign layer2_outputs[1049] = (layer1_outputs[2851]) & (layer1_outputs[2005]);
    assign layer2_outputs[1050] = (layer1_outputs[1308]) & ~(layer1_outputs[3156]);
    assign layer2_outputs[1051] = layer1_outputs[4921];
    assign layer2_outputs[1052] = ~((layer1_outputs[3357]) | (layer1_outputs[1498]));
    assign layer2_outputs[1053] = (layer1_outputs[3037]) | (layer1_outputs[719]);
    assign layer2_outputs[1054] = ~((layer1_outputs[2854]) & (layer1_outputs[2171]));
    assign layer2_outputs[1055] = ~(layer1_outputs[2482]);
    assign layer2_outputs[1056] = 1'b1;
    assign layer2_outputs[1057] = layer1_outputs[3133];
    assign layer2_outputs[1058] = ~((layer1_outputs[4686]) | (layer1_outputs[399]));
    assign layer2_outputs[1059] = ~(layer1_outputs[2991]);
    assign layer2_outputs[1060] = layer1_outputs[4104];
    assign layer2_outputs[1061] = (layer1_outputs[3095]) | (layer1_outputs[1051]);
    assign layer2_outputs[1062] = (layer1_outputs[607]) & (layer1_outputs[147]);
    assign layer2_outputs[1063] = 1'b0;
    assign layer2_outputs[1064] = 1'b1;
    assign layer2_outputs[1065] = 1'b1;
    assign layer2_outputs[1066] = ~(layer1_outputs[238]);
    assign layer2_outputs[1067] = (layer1_outputs[4424]) | (layer1_outputs[1571]);
    assign layer2_outputs[1068] = ~(layer1_outputs[766]);
    assign layer2_outputs[1069] = ~((layer1_outputs[4384]) | (layer1_outputs[2765]));
    assign layer2_outputs[1070] = ~((layer1_outputs[2727]) & (layer1_outputs[3947]));
    assign layer2_outputs[1071] = ~((layer1_outputs[5106]) & (layer1_outputs[4230]));
    assign layer2_outputs[1072] = 1'b0;
    assign layer2_outputs[1073] = (layer1_outputs[3678]) & ~(layer1_outputs[2172]);
    assign layer2_outputs[1074] = ~((layer1_outputs[1721]) & (layer1_outputs[874]));
    assign layer2_outputs[1075] = ~(layer1_outputs[4439]);
    assign layer2_outputs[1076] = ~((layer1_outputs[4865]) | (layer1_outputs[1204]));
    assign layer2_outputs[1077] = ~((layer1_outputs[1900]) | (layer1_outputs[2884]));
    assign layer2_outputs[1078] = ~((layer1_outputs[1675]) & (layer1_outputs[2717]));
    assign layer2_outputs[1079] = ~((layer1_outputs[2401]) & (layer1_outputs[4727]));
    assign layer2_outputs[1080] = (layer1_outputs[4045]) & ~(layer1_outputs[1537]);
    assign layer2_outputs[1081] = ~(layer1_outputs[2743]) | (layer1_outputs[932]);
    assign layer2_outputs[1082] = (layer1_outputs[64]) | (layer1_outputs[306]);
    assign layer2_outputs[1083] = ~((layer1_outputs[2945]) ^ (layer1_outputs[2472]));
    assign layer2_outputs[1084] = ~((layer1_outputs[2475]) | (layer1_outputs[4148]));
    assign layer2_outputs[1085] = ~((layer1_outputs[1312]) & (layer1_outputs[2424]));
    assign layer2_outputs[1086] = ~(layer1_outputs[2124]) | (layer1_outputs[1941]);
    assign layer2_outputs[1087] = layer1_outputs[2739];
    assign layer2_outputs[1088] = ~(layer1_outputs[1974]);
    assign layer2_outputs[1089] = ~(layer1_outputs[3771]);
    assign layer2_outputs[1090] = layer1_outputs[3722];
    assign layer2_outputs[1091] = ~(layer1_outputs[807]) | (layer1_outputs[4200]);
    assign layer2_outputs[1092] = ~(layer1_outputs[379]);
    assign layer2_outputs[1093] = (layer1_outputs[378]) & (layer1_outputs[1515]);
    assign layer2_outputs[1094] = 1'b0;
    assign layer2_outputs[1095] = (layer1_outputs[571]) ^ (layer1_outputs[1523]);
    assign layer2_outputs[1096] = ~(layer1_outputs[4204]) | (layer1_outputs[1250]);
    assign layer2_outputs[1097] = ~(layer1_outputs[1701]) | (layer1_outputs[4953]);
    assign layer2_outputs[1098] = ~(layer1_outputs[4651]);
    assign layer2_outputs[1099] = layer1_outputs[1730];
    assign layer2_outputs[1100] = 1'b0;
    assign layer2_outputs[1101] = ~((layer1_outputs[1924]) | (layer1_outputs[35]));
    assign layer2_outputs[1102] = ~((layer1_outputs[935]) | (layer1_outputs[3014]));
    assign layer2_outputs[1103] = ~((layer1_outputs[393]) & (layer1_outputs[1073]));
    assign layer2_outputs[1104] = ~((layer1_outputs[410]) & (layer1_outputs[1007]));
    assign layer2_outputs[1105] = ~((layer1_outputs[2981]) | (layer1_outputs[3048]));
    assign layer2_outputs[1106] = layer1_outputs[1276];
    assign layer2_outputs[1107] = ~((layer1_outputs[2928]) ^ (layer1_outputs[114]));
    assign layer2_outputs[1108] = ~(layer1_outputs[1014]);
    assign layer2_outputs[1109] = (layer1_outputs[1460]) | (layer1_outputs[1063]);
    assign layer2_outputs[1110] = (layer1_outputs[2834]) & ~(layer1_outputs[3022]);
    assign layer2_outputs[1111] = (layer1_outputs[3715]) & ~(layer1_outputs[2564]);
    assign layer2_outputs[1112] = layer1_outputs[756];
    assign layer2_outputs[1113] = (layer1_outputs[3647]) & ~(layer1_outputs[2868]);
    assign layer2_outputs[1114] = (layer1_outputs[4532]) & (layer1_outputs[4055]);
    assign layer2_outputs[1115] = layer1_outputs[417];
    assign layer2_outputs[1116] = ~((layer1_outputs[748]) & (layer1_outputs[3368]));
    assign layer2_outputs[1117] = 1'b1;
    assign layer2_outputs[1118] = (layer1_outputs[3949]) & (layer1_outputs[4337]);
    assign layer2_outputs[1119] = ~(layer1_outputs[4563]) | (layer1_outputs[4973]);
    assign layer2_outputs[1120] = (layer1_outputs[2839]) & (layer1_outputs[3645]);
    assign layer2_outputs[1121] = ~((layer1_outputs[1850]) & (layer1_outputs[2419]));
    assign layer2_outputs[1122] = ~((layer1_outputs[5107]) & (layer1_outputs[463]));
    assign layer2_outputs[1123] = layer1_outputs[4985];
    assign layer2_outputs[1124] = ~(layer1_outputs[2140]) | (layer1_outputs[3793]);
    assign layer2_outputs[1125] = ~(layer1_outputs[1481]);
    assign layer2_outputs[1126] = (layer1_outputs[3282]) & ~(layer1_outputs[1434]);
    assign layer2_outputs[1127] = ~(layer1_outputs[830]);
    assign layer2_outputs[1128] = ~(layer1_outputs[3907]) | (layer1_outputs[4540]);
    assign layer2_outputs[1129] = (layer1_outputs[4509]) & ~(layer1_outputs[3729]);
    assign layer2_outputs[1130] = 1'b0;
    assign layer2_outputs[1131] = layer1_outputs[3830];
    assign layer2_outputs[1132] = (layer1_outputs[3343]) & ~(layer1_outputs[23]);
    assign layer2_outputs[1133] = (layer1_outputs[1469]) & ~(layer1_outputs[2347]);
    assign layer2_outputs[1134] = 1'b0;
    assign layer2_outputs[1135] = (layer1_outputs[443]) ^ (layer1_outputs[4924]);
    assign layer2_outputs[1136] = 1'b1;
    assign layer2_outputs[1137] = 1'b0;
    assign layer2_outputs[1138] = layer1_outputs[1136];
    assign layer2_outputs[1139] = ~((layer1_outputs[2952]) & (layer1_outputs[2418]));
    assign layer2_outputs[1140] = ~(layer1_outputs[3917]) | (layer1_outputs[4719]);
    assign layer2_outputs[1141] = (layer1_outputs[4087]) & ~(layer1_outputs[357]);
    assign layer2_outputs[1142] = layer1_outputs[1747];
    assign layer2_outputs[1143] = 1'b0;
    assign layer2_outputs[1144] = 1'b1;
    assign layer2_outputs[1145] = ~(layer1_outputs[206]);
    assign layer2_outputs[1146] = ~(layer1_outputs[3463]);
    assign layer2_outputs[1147] = ~(layer1_outputs[333]);
    assign layer2_outputs[1148] = ~(layer1_outputs[4438]) | (layer1_outputs[1092]);
    assign layer2_outputs[1149] = 1'b1;
    assign layer2_outputs[1150] = ~(layer1_outputs[33]) | (layer1_outputs[667]);
    assign layer2_outputs[1151] = ~(layer1_outputs[817]) | (layer1_outputs[3758]);
    assign layer2_outputs[1152] = ~((layer1_outputs[2869]) & (layer1_outputs[1743]));
    assign layer2_outputs[1153] = ~(layer1_outputs[5014]) | (layer1_outputs[726]);
    assign layer2_outputs[1154] = ~((layer1_outputs[1202]) & (layer1_outputs[2719]));
    assign layer2_outputs[1155] = (layer1_outputs[665]) | (layer1_outputs[1082]);
    assign layer2_outputs[1156] = ~((layer1_outputs[1720]) | (layer1_outputs[4194]));
    assign layer2_outputs[1157] = layer1_outputs[4861];
    assign layer2_outputs[1158] = layer1_outputs[4430];
    assign layer2_outputs[1159] = (layer1_outputs[3464]) ^ (layer1_outputs[3069]);
    assign layer2_outputs[1160] = ~((layer1_outputs[1934]) | (layer1_outputs[2276]));
    assign layer2_outputs[1161] = (layer1_outputs[1722]) | (layer1_outputs[4113]);
    assign layer2_outputs[1162] = ~(layer1_outputs[2448]);
    assign layer2_outputs[1163] = 1'b0;
    assign layer2_outputs[1164] = layer1_outputs[3887];
    assign layer2_outputs[1165] = (layer1_outputs[4702]) | (layer1_outputs[269]);
    assign layer2_outputs[1166] = ~(layer1_outputs[2960]);
    assign layer2_outputs[1167] = (layer1_outputs[2555]) ^ (layer1_outputs[2342]);
    assign layer2_outputs[1168] = ~(layer1_outputs[818]) | (layer1_outputs[547]);
    assign layer2_outputs[1169] = (layer1_outputs[110]) & ~(layer1_outputs[614]);
    assign layer2_outputs[1170] = ~((layer1_outputs[2075]) | (layer1_outputs[1097]));
    assign layer2_outputs[1171] = ~((layer1_outputs[3627]) | (layer1_outputs[4808]));
    assign layer2_outputs[1172] = ~(layer1_outputs[1190]) | (layer1_outputs[3212]);
    assign layer2_outputs[1173] = layer1_outputs[178];
    assign layer2_outputs[1174] = ~(layer1_outputs[1620]);
    assign layer2_outputs[1175] = ~(layer1_outputs[2915]);
    assign layer2_outputs[1176] = ~((layer1_outputs[3629]) & (layer1_outputs[3493]));
    assign layer2_outputs[1177] = ~(layer1_outputs[1817]) | (layer1_outputs[1875]);
    assign layer2_outputs[1178] = layer1_outputs[3422];
    assign layer2_outputs[1179] = (layer1_outputs[4214]) & ~(layer1_outputs[2977]);
    assign layer2_outputs[1180] = ~(layer1_outputs[2699]);
    assign layer2_outputs[1181] = ~(layer1_outputs[3188]) | (layer1_outputs[1383]);
    assign layer2_outputs[1182] = ~(layer1_outputs[2991]);
    assign layer2_outputs[1183] = (layer1_outputs[1351]) | (layer1_outputs[3036]);
    assign layer2_outputs[1184] = ~(layer1_outputs[1719]) | (layer1_outputs[1098]);
    assign layer2_outputs[1185] = ~(layer1_outputs[4145]);
    assign layer2_outputs[1186] = ~(layer1_outputs[111]);
    assign layer2_outputs[1187] = ~(layer1_outputs[5021]);
    assign layer2_outputs[1188] = ~(layer1_outputs[776]);
    assign layer2_outputs[1189] = layer1_outputs[1126];
    assign layer2_outputs[1190] = ~(layer1_outputs[1238]) | (layer1_outputs[3631]);
    assign layer2_outputs[1191] = layer1_outputs[4103];
    assign layer2_outputs[1192] = ~(layer1_outputs[3929]) | (layer1_outputs[3885]);
    assign layer2_outputs[1193] = ~(layer1_outputs[4100]);
    assign layer2_outputs[1194] = layer1_outputs[1112];
    assign layer2_outputs[1195] = ~(layer1_outputs[3641]) | (layer1_outputs[39]);
    assign layer2_outputs[1196] = (layer1_outputs[2821]) | (layer1_outputs[4481]);
    assign layer2_outputs[1197] = ~(layer1_outputs[4302]) | (layer1_outputs[573]);
    assign layer2_outputs[1198] = (layer1_outputs[1825]) & ~(layer1_outputs[23]);
    assign layer2_outputs[1199] = ~((layer1_outputs[2672]) & (layer1_outputs[4837]));
    assign layer2_outputs[1200] = (layer1_outputs[1583]) & ~(layer1_outputs[1286]);
    assign layer2_outputs[1201] = (layer1_outputs[1657]) & ~(layer1_outputs[4854]);
    assign layer2_outputs[1202] = ~(layer1_outputs[3618]) | (layer1_outputs[1939]);
    assign layer2_outputs[1203] = (layer1_outputs[1145]) & (layer1_outputs[439]);
    assign layer2_outputs[1204] = layer1_outputs[4498];
    assign layer2_outputs[1205] = layer1_outputs[71];
    assign layer2_outputs[1206] = 1'b1;
    assign layer2_outputs[1207] = ~((layer1_outputs[3514]) | (layer1_outputs[4482]));
    assign layer2_outputs[1208] = 1'b0;
    assign layer2_outputs[1209] = 1'b1;
    assign layer2_outputs[1210] = (layer1_outputs[1207]) & ~(layer1_outputs[71]);
    assign layer2_outputs[1211] = (layer1_outputs[814]) | (layer1_outputs[4571]);
    assign layer2_outputs[1212] = ~(layer1_outputs[4674]) | (layer1_outputs[1245]);
    assign layer2_outputs[1213] = ~((layer1_outputs[5084]) | (layer1_outputs[4094]));
    assign layer2_outputs[1214] = 1'b0;
    assign layer2_outputs[1215] = (layer1_outputs[2480]) & ~(layer1_outputs[2541]);
    assign layer2_outputs[1216] = 1'b1;
    assign layer2_outputs[1217] = (layer1_outputs[151]) & (layer1_outputs[1553]);
    assign layer2_outputs[1218] = ~(layer1_outputs[681]) | (layer1_outputs[2611]);
    assign layer2_outputs[1219] = ~(layer1_outputs[3476]) | (layer1_outputs[4940]);
    assign layer2_outputs[1220] = 1'b1;
    assign layer2_outputs[1221] = (layer1_outputs[370]) & ~(layer1_outputs[1197]);
    assign layer2_outputs[1222] = ~(layer1_outputs[2837]);
    assign layer2_outputs[1223] = 1'b0;
    assign layer2_outputs[1224] = ~(layer1_outputs[1868]);
    assign layer2_outputs[1225] = layer1_outputs[2887];
    assign layer2_outputs[1226] = (layer1_outputs[1545]) & (layer1_outputs[1132]);
    assign layer2_outputs[1227] = ~(layer1_outputs[2397]);
    assign layer2_outputs[1228] = ~((layer1_outputs[3596]) | (layer1_outputs[1972]));
    assign layer2_outputs[1229] = (layer1_outputs[1515]) & (layer1_outputs[596]);
    assign layer2_outputs[1230] = 1'b0;
    assign layer2_outputs[1231] = ~(layer1_outputs[4866]);
    assign layer2_outputs[1232] = layer1_outputs[3025];
    assign layer2_outputs[1233] = (layer1_outputs[2427]) & (layer1_outputs[1288]);
    assign layer2_outputs[1234] = ~(layer1_outputs[555]);
    assign layer2_outputs[1235] = 1'b0;
    assign layer2_outputs[1236] = 1'b0;
    assign layer2_outputs[1237] = layer1_outputs[2318];
    assign layer2_outputs[1238] = ~(layer1_outputs[3576]);
    assign layer2_outputs[1239] = 1'b0;
    assign layer2_outputs[1240] = layer1_outputs[3797];
    assign layer2_outputs[1241] = ~(layer1_outputs[1644]);
    assign layer2_outputs[1242] = ~((layer1_outputs[4272]) ^ (layer1_outputs[3424]));
    assign layer2_outputs[1243] = (layer1_outputs[3617]) | (layer1_outputs[1034]);
    assign layer2_outputs[1244] = ~(layer1_outputs[1698]);
    assign layer2_outputs[1245] = layer1_outputs[1681];
    assign layer2_outputs[1246] = ~((layer1_outputs[3883]) | (layer1_outputs[5000]));
    assign layer2_outputs[1247] = ~(layer1_outputs[4465]);
    assign layer2_outputs[1248] = (layer1_outputs[2146]) & (layer1_outputs[2720]);
    assign layer2_outputs[1249] = ~((layer1_outputs[2016]) | (layer1_outputs[3638]));
    assign layer2_outputs[1250] = (layer1_outputs[3805]) & ~(layer1_outputs[1765]);
    assign layer2_outputs[1251] = (layer1_outputs[1988]) | (layer1_outputs[4779]);
    assign layer2_outputs[1252] = (layer1_outputs[5109]) & ~(layer1_outputs[946]);
    assign layer2_outputs[1253] = ~((layer1_outputs[2436]) | (layer1_outputs[3291]));
    assign layer2_outputs[1254] = layer1_outputs[1243];
    assign layer2_outputs[1255] = (layer1_outputs[2810]) | (layer1_outputs[4077]);
    assign layer2_outputs[1256] = 1'b0;
    assign layer2_outputs[1257] = (layer1_outputs[4748]) & ~(layer1_outputs[1459]);
    assign layer2_outputs[1258] = 1'b1;
    assign layer2_outputs[1259] = ~((layer1_outputs[363]) ^ (layer1_outputs[2300]));
    assign layer2_outputs[1260] = (layer1_outputs[565]) | (layer1_outputs[3035]);
    assign layer2_outputs[1261] = (layer1_outputs[4773]) ^ (layer1_outputs[1189]);
    assign layer2_outputs[1262] = ~(layer1_outputs[4114]) | (layer1_outputs[1063]);
    assign layer2_outputs[1263] = ~((layer1_outputs[3006]) & (layer1_outputs[2732]));
    assign layer2_outputs[1264] = 1'b0;
    assign layer2_outputs[1265] = layer1_outputs[3817];
    assign layer2_outputs[1266] = layer1_outputs[2782];
    assign layer2_outputs[1267] = ~((layer1_outputs[2145]) & (layer1_outputs[679]));
    assign layer2_outputs[1268] = ~(layer1_outputs[404]);
    assign layer2_outputs[1269] = ~(layer1_outputs[2101]);
    assign layer2_outputs[1270] = (layer1_outputs[3354]) & ~(layer1_outputs[1706]);
    assign layer2_outputs[1271] = ~((layer1_outputs[955]) | (layer1_outputs[4879]));
    assign layer2_outputs[1272] = ~(layer1_outputs[4411]) | (layer1_outputs[3004]);
    assign layer2_outputs[1273] = 1'b1;
    assign layer2_outputs[1274] = (layer1_outputs[723]) & ~(layer1_outputs[2590]);
    assign layer2_outputs[1275] = (layer1_outputs[4075]) & ~(layer1_outputs[3770]);
    assign layer2_outputs[1276] = ~((layer1_outputs[4213]) ^ (layer1_outputs[1832]));
    assign layer2_outputs[1277] = ~((layer1_outputs[1673]) | (layer1_outputs[4586]));
    assign layer2_outputs[1278] = 1'b1;
    assign layer2_outputs[1279] = ~(layer1_outputs[373]) | (layer1_outputs[1287]);
    assign layer2_outputs[1280] = ~(layer1_outputs[3265]) | (layer1_outputs[1024]);
    assign layer2_outputs[1281] = (layer1_outputs[100]) ^ (layer1_outputs[1677]);
    assign layer2_outputs[1282] = 1'b1;
    assign layer2_outputs[1283] = layer1_outputs[3327];
    assign layer2_outputs[1284] = ~(layer1_outputs[515]);
    assign layer2_outputs[1285] = ~((layer1_outputs[2895]) & (layer1_outputs[1130]));
    assign layer2_outputs[1286] = (layer1_outputs[1712]) & ~(layer1_outputs[728]);
    assign layer2_outputs[1287] = layer1_outputs[4397];
    assign layer2_outputs[1288] = 1'b0;
    assign layer2_outputs[1289] = layer1_outputs[4445];
    assign layer2_outputs[1290] = layer1_outputs[2311];
    assign layer2_outputs[1291] = layer1_outputs[1297];
    assign layer2_outputs[1292] = ~(layer1_outputs[691]);
    assign layer2_outputs[1293] = ~(layer1_outputs[1401]);
    assign layer2_outputs[1294] = 1'b0;
    assign layer2_outputs[1295] = layer1_outputs[1054];
    assign layer2_outputs[1296] = ~(layer1_outputs[4318]) | (layer1_outputs[3965]);
    assign layer2_outputs[1297] = ~(layer1_outputs[2767]) | (layer1_outputs[4026]);
    assign layer2_outputs[1298] = layer1_outputs[3086];
    assign layer2_outputs[1299] = ~((layer1_outputs[2082]) ^ (layer1_outputs[85]));
    assign layer2_outputs[1300] = (layer1_outputs[3606]) & ~(layer1_outputs[404]);
    assign layer2_outputs[1301] = (layer1_outputs[627]) & ~(layer1_outputs[3437]);
    assign layer2_outputs[1302] = layer1_outputs[5013];
    assign layer2_outputs[1303] = ~((layer1_outputs[2095]) & (layer1_outputs[3581]));
    assign layer2_outputs[1304] = (layer1_outputs[772]) | (layer1_outputs[3853]);
    assign layer2_outputs[1305] = (layer1_outputs[3313]) | (layer1_outputs[3628]);
    assign layer2_outputs[1306] = (layer1_outputs[3165]) & ~(layer1_outputs[1959]);
    assign layer2_outputs[1307] = (layer1_outputs[2995]) ^ (layer1_outputs[4803]);
    assign layer2_outputs[1308] = (layer1_outputs[1049]) | (layer1_outputs[3714]);
    assign layer2_outputs[1309] = ~((layer1_outputs[3006]) | (layer1_outputs[1328]));
    assign layer2_outputs[1310] = ~((layer1_outputs[3143]) | (layer1_outputs[4829]));
    assign layer2_outputs[1311] = ~(layer1_outputs[4772]);
    assign layer2_outputs[1312] = ~(layer1_outputs[2423]) | (layer1_outputs[947]);
    assign layer2_outputs[1313] = (layer1_outputs[2831]) | (layer1_outputs[594]);
    assign layer2_outputs[1314] = ~(layer1_outputs[4603]) | (layer1_outputs[2135]);
    assign layer2_outputs[1315] = ~(layer1_outputs[4800]);
    assign layer2_outputs[1316] = 1'b1;
    assign layer2_outputs[1317] = (layer1_outputs[3752]) & ~(layer1_outputs[4736]);
    assign layer2_outputs[1318] = (layer1_outputs[3451]) | (layer1_outputs[737]);
    assign layer2_outputs[1319] = ~((layer1_outputs[451]) ^ (layer1_outputs[728]));
    assign layer2_outputs[1320] = ~(layer1_outputs[3799]);
    assign layer2_outputs[1321] = ~((layer1_outputs[4047]) & (layer1_outputs[961]));
    assign layer2_outputs[1322] = layer1_outputs[2738];
    assign layer2_outputs[1323] = (layer1_outputs[2710]) & (layer1_outputs[2892]);
    assign layer2_outputs[1324] = layer1_outputs[3507];
    assign layer2_outputs[1325] = (layer1_outputs[495]) | (layer1_outputs[2920]);
    assign layer2_outputs[1326] = (layer1_outputs[653]) & (layer1_outputs[2089]);
    assign layer2_outputs[1327] = (layer1_outputs[414]) & (layer1_outputs[2220]);
    assign layer2_outputs[1328] = 1'b0;
    assign layer2_outputs[1329] = ~(layer1_outputs[3127]);
    assign layer2_outputs[1330] = ~(layer1_outputs[2940]);
    assign layer2_outputs[1331] = ~((layer1_outputs[1894]) ^ (layer1_outputs[2147]));
    assign layer2_outputs[1332] = layer1_outputs[2003];
    assign layer2_outputs[1333] = layer1_outputs[2078];
    assign layer2_outputs[1334] = (layer1_outputs[1155]) & ~(layer1_outputs[4614]);
    assign layer2_outputs[1335] = (layer1_outputs[934]) & ~(layer1_outputs[2578]);
    assign layer2_outputs[1336] = ~(layer1_outputs[2446]);
    assign layer2_outputs[1337] = ~((layer1_outputs[223]) & (layer1_outputs[4882]));
    assign layer2_outputs[1338] = ~((layer1_outputs[1306]) ^ (layer1_outputs[3054]));
    assign layer2_outputs[1339] = ~(layer1_outputs[4669]) | (layer1_outputs[388]);
    assign layer2_outputs[1340] = (layer1_outputs[4680]) | (layer1_outputs[3828]);
    assign layer2_outputs[1341] = (layer1_outputs[3281]) | (layer1_outputs[2043]);
    assign layer2_outputs[1342] = (layer1_outputs[1617]) & (layer1_outputs[274]);
    assign layer2_outputs[1343] = (layer1_outputs[3088]) & (layer1_outputs[3425]);
    assign layer2_outputs[1344] = ~(layer1_outputs[1662]);
    assign layer2_outputs[1345] = ~((layer1_outputs[4734]) ^ (layer1_outputs[3831]));
    assign layer2_outputs[1346] = layer1_outputs[4731];
    assign layer2_outputs[1347] = (layer1_outputs[691]) & ~(layer1_outputs[58]);
    assign layer2_outputs[1348] = layer1_outputs[1601];
    assign layer2_outputs[1349] = 1'b0;
    assign layer2_outputs[1350] = 1'b0;
    assign layer2_outputs[1351] = 1'b0;
    assign layer2_outputs[1352] = ~(layer1_outputs[1271]) | (layer1_outputs[156]);
    assign layer2_outputs[1353] = ~(layer1_outputs[3326]);
    assign layer2_outputs[1354] = ~(layer1_outputs[2969]);
    assign layer2_outputs[1355] = ~((layer1_outputs[2029]) & (layer1_outputs[2257]));
    assign layer2_outputs[1356] = (layer1_outputs[974]) & ~(layer1_outputs[2100]);
    assign layer2_outputs[1357] = ~((layer1_outputs[1745]) | (layer1_outputs[697]));
    assign layer2_outputs[1358] = ~(layer1_outputs[2248]);
    assign layer2_outputs[1359] = (layer1_outputs[1461]) & ~(layer1_outputs[1156]);
    assign layer2_outputs[1360] = ~((layer1_outputs[2127]) | (layer1_outputs[3219]));
    assign layer2_outputs[1361] = (layer1_outputs[4581]) | (layer1_outputs[4724]);
    assign layer2_outputs[1362] = (layer1_outputs[1213]) | (layer1_outputs[1743]);
    assign layer2_outputs[1363] = ~(layer1_outputs[2653]) | (layer1_outputs[4348]);
    assign layer2_outputs[1364] = 1'b1;
    assign layer2_outputs[1365] = ~(layer1_outputs[3027]) | (layer1_outputs[3751]);
    assign layer2_outputs[1366] = ~(layer1_outputs[5047]) | (layer1_outputs[4304]);
    assign layer2_outputs[1367] = (layer1_outputs[144]) & ~(layer1_outputs[1910]);
    assign layer2_outputs[1368] = (layer1_outputs[2792]) & ~(layer1_outputs[3951]);
    assign layer2_outputs[1369] = layer1_outputs[4004];
    assign layer2_outputs[1370] = (layer1_outputs[296]) | (layer1_outputs[4905]);
    assign layer2_outputs[1371] = ~((layer1_outputs[4979]) | (layer1_outputs[3039]));
    assign layer2_outputs[1372] = ~(layer1_outputs[3962]);
    assign layer2_outputs[1373] = (layer1_outputs[5077]) | (layer1_outputs[5114]);
    assign layer2_outputs[1374] = ~((layer1_outputs[739]) | (layer1_outputs[3675]));
    assign layer2_outputs[1375] = (layer1_outputs[1203]) & (layer1_outputs[1554]);
    assign layer2_outputs[1376] = (layer1_outputs[1842]) & ~(layer1_outputs[2845]);
    assign layer2_outputs[1377] = 1'b0;
    assign layer2_outputs[1378] = layer1_outputs[5020];
    assign layer2_outputs[1379] = 1'b1;
    assign layer2_outputs[1380] = ~(layer1_outputs[4135]) | (layer1_outputs[2790]);
    assign layer2_outputs[1381] = ~(layer1_outputs[2635]) | (layer1_outputs[4594]);
    assign layer2_outputs[1382] = ~((layer1_outputs[1878]) & (layer1_outputs[583]));
    assign layer2_outputs[1383] = ~((layer1_outputs[205]) | (layer1_outputs[2423]));
    assign layer2_outputs[1384] = 1'b1;
    assign layer2_outputs[1385] = layer1_outputs[4209];
    assign layer2_outputs[1386] = (layer1_outputs[3318]) & ~(layer1_outputs[4654]);
    assign layer2_outputs[1387] = ~(layer1_outputs[1000]);
    assign layer2_outputs[1388] = (layer1_outputs[3613]) | (layer1_outputs[2361]);
    assign layer2_outputs[1389] = ~((layer1_outputs[1052]) & (layer1_outputs[4155]));
    assign layer2_outputs[1390] = ~(layer1_outputs[2897]);
    assign layer2_outputs[1391] = layer1_outputs[2980];
    assign layer2_outputs[1392] = (layer1_outputs[4621]) & ~(layer1_outputs[891]);
    assign layer2_outputs[1393] = layer1_outputs[2132];
    assign layer2_outputs[1394] = ~(layer1_outputs[2409]);
    assign layer2_outputs[1395] = ~(layer1_outputs[2215]);
    assign layer2_outputs[1396] = 1'b0;
    assign layer2_outputs[1397] = ~((layer1_outputs[4102]) | (layer1_outputs[2592]));
    assign layer2_outputs[1398] = (layer1_outputs[299]) & ~(layer1_outputs[3653]);
    assign layer2_outputs[1399] = (layer1_outputs[2703]) ^ (layer1_outputs[2944]);
    assign layer2_outputs[1400] = 1'b1;
    assign layer2_outputs[1401] = (layer1_outputs[1138]) & (layer1_outputs[1263]);
    assign layer2_outputs[1402] = (layer1_outputs[1861]) ^ (layer1_outputs[788]);
    assign layer2_outputs[1403] = layer1_outputs[311];
    assign layer2_outputs[1404] = ~(layer1_outputs[3128]);
    assign layer2_outputs[1405] = layer1_outputs[4136];
    assign layer2_outputs[1406] = ~(layer1_outputs[612]) | (layer1_outputs[2825]);
    assign layer2_outputs[1407] = (layer1_outputs[3154]) & ~(layer1_outputs[2381]);
    assign layer2_outputs[1408] = (layer1_outputs[1055]) & ~(layer1_outputs[1464]);
    assign layer2_outputs[1409] = 1'b0;
    assign layer2_outputs[1410] = (layer1_outputs[215]) & ~(layer1_outputs[812]);
    assign layer2_outputs[1411] = 1'b1;
    assign layer2_outputs[1412] = ~(layer1_outputs[1178]) | (layer1_outputs[3175]);
    assign layer2_outputs[1413] = ~(layer1_outputs[3743]);
    assign layer2_outputs[1414] = ~(layer1_outputs[3465]) | (layer1_outputs[1963]);
    assign layer2_outputs[1415] = ~(layer1_outputs[979]);
    assign layer2_outputs[1416] = 1'b0;
    assign layer2_outputs[1417] = ~(layer1_outputs[532]) | (layer1_outputs[1521]);
    assign layer2_outputs[1418] = (layer1_outputs[1503]) & ~(layer1_outputs[1080]);
    assign layer2_outputs[1419] = ~((layer1_outputs[1854]) & (layer1_outputs[13]));
    assign layer2_outputs[1420] = 1'b1;
    assign layer2_outputs[1421] = ~(layer1_outputs[2958]);
    assign layer2_outputs[1422] = ~(layer1_outputs[825]);
    assign layer2_outputs[1423] = (layer1_outputs[376]) & (layer1_outputs[3642]);
    assign layer2_outputs[1424] = (layer1_outputs[4544]) & ~(layer1_outputs[3366]);
    assign layer2_outputs[1425] = (layer1_outputs[3323]) & ~(layer1_outputs[2121]);
    assign layer2_outputs[1426] = (layer1_outputs[1921]) & ~(layer1_outputs[2254]);
    assign layer2_outputs[1427] = 1'b1;
    assign layer2_outputs[1428] = ~((layer1_outputs[4142]) ^ (layer1_outputs[282]));
    assign layer2_outputs[1429] = ~(layer1_outputs[1762]) | (layer1_outputs[1580]);
    assign layer2_outputs[1430] = 1'b1;
    assign layer2_outputs[1431] = ~(layer1_outputs[4438]) | (layer1_outputs[4443]);
    assign layer2_outputs[1432] = ~(layer1_outputs[3405]);
    assign layer2_outputs[1433] = 1'b0;
    assign layer2_outputs[1434] = ~(layer1_outputs[2311]) | (layer1_outputs[5012]);
    assign layer2_outputs[1435] = (layer1_outputs[4379]) | (layer1_outputs[1720]);
    assign layer2_outputs[1436] = ~(layer1_outputs[1660]);
    assign layer2_outputs[1437] = (layer1_outputs[482]) & ~(layer1_outputs[1626]);
    assign layer2_outputs[1438] = ~(layer1_outputs[718]);
    assign layer2_outputs[1439] = 1'b1;
    assign layer2_outputs[1440] = ~(layer1_outputs[3420]) | (layer1_outputs[3840]);
    assign layer2_outputs[1441] = layer1_outputs[153];
    assign layer2_outputs[1442] = ~((layer1_outputs[4136]) & (layer1_outputs[1043]));
    assign layer2_outputs[1443] = ~(layer1_outputs[4501]);
    assign layer2_outputs[1444] = 1'b0;
    assign layer2_outputs[1445] = layer1_outputs[2733];
    assign layer2_outputs[1446] = ~(layer1_outputs[794]);
    assign layer2_outputs[1447] = ~((layer1_outputs[1407]) ^ (layer1_outputs[2227]));
    assign layer2_outputs[1448] = 1'b1;
    assign layer2_outputs[1449] = (layer1_outputs[285]) & (layer1_outputs[588]);
    assign layer2_outputs[1450] = ~(layer1_outputs[2253]) | (layer1_outputs[458]);
    assign layer2_outputs[1451] = ~(layer1_outputs[2973]);
    assign layer2_outputs[1452] = ~((layer1_outputs[4098]) | (layer1_outputs[2040]));
    assign layer2_outputs[1453] = (layer1_outputs[3337]) | (layer1_outputs[2918]);
    assign layer2_outputs[1454] = ~(layer1_outputs[4491]);
    assign layer2_outputs[1455] = 1'b0;
    assign layer2_outputs[1456] = ~(layer1_outputs[1892]);
    assign layer2_outputs[1457] = layer1_outputs[4639];
    assign layer2_outputs[1458] = 1'b1;
    assign layer2_outputs[1459] = layer1_outputs[183];
    assign layer2_outputs[1460] = ~((layer1_outputs[2382]) & (layer1_outputs[4725]));
    assign layer2_outputs[1461] = (layer1_outputs[2775]) & (layer1_outputs[4796]);
    assign layer2_outputs[1462] = ~(layer1_outputs[1587]) | (layer1_outputs[1985]);
    assign layer2_outputs[1463] = (layer1_outputs[4065]) & ~(layer1_outputs[4434]);
    assign layer2_outputs[1464] = layer1_outputs[2417];
    assign layer2_outputs[1465] = (layer1_outputs[4462]) & ~(layer1_outputs[2984]);
    assign layer2_outputs[1466] = ~(layer1_outputs[2274]);
    assign layer2_outputs[1467] = layer1_outputs[3280];
    assign layer2_outputs[1468] = (layer1_outputs[647]) & ~(layer1_outputs[1919]);
    assign layer2_outputs[1469] = ~(layer1_outputs[1605]);
    assign layer2_outputs[1470] = ~((layer1_outputs[4862]) | (layer1_outputs[2380]));
    assign layer2_outputs[1471] = ~(layer1_outputs[3411]) | (layer1_outputs[729]);
    assign layer2_outputs[1472] = ~(layer1_outputs[2856]);
    assign layer2_outputs[1473] = ~(layer1_outputs[2065]);
    assign layer2_outputs[1474] = ~((layer1_outputs[4709]) & (layer1_outputs[4199]));
    assign layer2_outputs[1475] = layer1_outputs[2571];
    assign layer2_outputs[1476] = (layer1_outputs[2685]) ^ (layer1_outputs[5059]);
    assign layer2_outputs[1477] = layer1_outputs[1198];
    assign layer2_outputs[1478] = ~(layer1_outputs[2024]) | (layer1_outputs[2406]);
    assign layer2_outputs[1479] = 1'b1;
    assign layer2_outputs[1480] = 1'b1;
    assign layer2_outputs[1481] = (layer1_outputs[3531]) | (layer1_outputs[3443]);
    assign layer2_outputs[1482] = (layer1_outputs[103]) | (layer1_outputs[4891]);
    assign layer2_outputs[1483] = (layer1_outputs[465]) & (layer1_outputs[2989]);
    assign layer2_outputs[1484] = (layer1_outputs[1405]) & ~(layer1_outputs[4756]);
    assign layer2_outputs[1485] = ~(layer1_outputs[2695]) | (layer1_outputs[3223]);
    assign layer2_outputs[1486] = ~(layer1_outputs[4996]);
    assign layer2_outputs[1487] = (layer1_outputs[4336]) & (layer1_outputs[678]);
    assign layer2_outputs[1488] = layer1_outputs[1004];
    assign layer2_outputs[1489] = ~((layer1_outputs[3763]) & (layer1_outputs[2086]));
    assign layer2_outputs[1490] = ~((layer1_outputs[2587]) | (layer1_outputs[4529]));
    assign layer2_outputs[1491] = (layer1_outputs[1117]) & ~(layer1_outputs[1827]);
    assign layer2_outputs[1492] = layer1_outputs[1529];
    assign layer2_outputs[1493] = layer1_outputs[4076];
    assign layer2_outputs[1494] = layer1_outputs[4181];
    assign layer2_outputs[1495] = (layer1_outputs[866]) & (layer1_outputs[2400]);
    assign layer2_outputs[1496] = layer1_outputs[3517];
    assign layer2_outputs[1497] = (layer1_outputs[1707]) & (layer1_outputs[2218]);
    assign layer2_outputs[1498] = (layer1_outputs[4914]) & ~(layer1_outputs[770]);
    assign layer2_outputs[1499] = ~(layer1_outputs[2994]);
    assign layer2_outputs[1500] = 1'b1;
    assign layer2_outputs[1501] = (layer1_outputs[2702]) & (layer1_outputs[3902]);
    assign layer2_outputs[1502] = (layer1_outputs[237]) | (layer1_outputs[4464]);
    assign layer2_outputs[1503] = 1'b1;
    assign layer2_outputs[1504] = 1'b1;
    assign layer2_outputs[1505] = layer1_outputs[1680];
    assign layer2_outputs[1506] = 1'b0;
    assign layer2_outputs[1507] = ~(layer1_outputs[4460]);
    assign layer2_outputs[1508] = ~(layer1_outputs[4540]) | (layer1_outputs[4646]);
    assign layer2_outputs[1509] = ~((layer1_outputs[2522]) | (layer1_outputs[4974]));
    assign layer2_outputs[1510] = layer1_outputs[3621];
    assign layer2_outputs[1511] = layer1_outputs[1312];
    assign layer2_outputs[1512] = 1'b0;
    assign layer2_outputs[1513] = ~(layer1_outputs[1158]) | (layer1_outputs[1675]);
    assign layer2_outputs[1514] = ~(layer1_outputs[794]);
    assign layer2_outputs[1515] = (layer1_outputs[3188]) & ~(layer1_outputs[1142]);
    assign layer2_outputs[1516] = layer1_outputs[2559];
    assign layer2_outputs[1517] = 1'b0;
    assign layer2_outputs[1518] = layer1_outputs[4875];
    assign layer2_outputs[1519] = (layer1_outputs[24]) & (layer1_outputs[628]);
    assign layer2_outputs[1520] = ~(layer1_outputs[2414]) | (layer1_outputs[3511]);
    assign layer2_outputs[1521] = (layer1_outputs[2505]) | (layer1_outputs[1847]);
    assign layer2_outputs[1522] = 1'b0;
    assign layer2_outputs[1523] = ~(layer1_outputs[3939]) | (layer1_outputs[2425]);
    assign layer2_outputs[1524] = ~(layer1_outputs[3630]);
    assign layer2_outputs[1525] = 1'b1;
    assign layer2_outputs[1526] = 1'b1;
    assign layer2_outputs[1527] = 1'b1;
    assign layer2_outputs[1528] = (layer1_outputs[648]) | (layer1_outputs[1284]);
    assign layer2_outputs[1529] = 1'b1;
    assign layer2_outputs[1530] = ~(layer1_outputs[3836]);
    assign layer2_outputs[1531] = (layer1_outputs[914]) | (layer1_outputs[1616]);
    assign layer2_outputs[1532] = ~((layer1_outputs[2868]) & (layer1_outputs[1934]));
    assign layer2_outputs[1533] = ~((layer1_outputs[684]) & (layer1_outputs[3278]));
    assign layer2_outputs[1534] = 1'b0;
    assign layer2_outputs[1535] = layer1_outputs[3135];
    assign layer2_outputs[1536] = ~((layer1_outputs[4929]) & (layer1_outputs[4880]));
    assign layer2_outputs[1537] = ~((layer1_outputs[4938]) ^ (layer1_outputs[2766]));
    assign layer2_outputs[1538] = 1'b1;
    assign layer2_outputs[1539] = layer1_outputs[1547];
    assign layer2_outputs[1540] = 1'b0;
    assign layer2_outputs[1541] = layer1_outputs[4274];
    assign layer2_outputs[1542] = ~(layer1_outputs[3040]);
    assign layer2_outputs[1543] = ~(layer1_outputs[3931]) | (layer1_outputs[2232]);
    assign layer2_outputs[1544] = layer1_outputs[3028];
    assign layer2_outputs[1545] = 1'b1;
    assign layer2_outputs[1546] = 1'b1;
    assign layer2_outputs[1547] = (layer1_outputs[1750]) ^ (layer1_outputs[2857]);
    assign layer2_outputs[1548] = ~((layer1_outputs[1454]) & (layer1_outputs[2694]));
    assign layer2_outputs[1549] = (layer1_outputs[4573]) & ~(layer1_outputs[3822]);
    assign layer2_outputs[1550] = ~(layer1_outputs[4269]) | (layer1_outputs[657]);
    assign layer2_outputs[1551] = ~((layer1_outputs[817]) & (layer1_outputs[2688]));
    assign layer2_outputs[1552] = layer1_outputs[2917];
    assign layer2_outputs[1553] = (layer1_outputs[2039]) & (layer1_outputs[3713]);
    assign layer2_outputs[1554] = ~(layer1_outputs[4810]);
    assign layer2_outputs[1555] = ~((layer1_outputs[5049]) ^ (layer1_outputs[2579]));
    assign layer2_outputs[1556] = ~(layer1_outputs[3221]);
    assign layer2_outputs[1557] = (layer1_outputs[4694]) & ~(layer1_outputs[3375]);
    assign layer2_outputs[1558] = (layer1_outputs[4019]) & ~(layer1_outputs[2191]);
    assign layer2_outputs[1559] = (layer1_outputs[1417]) | (layer1_outputs[1153]);
    assign layer2_outputs[1560] = layer1_outputs[2539];
    assign layer2_outputs[1561] = 1'b0;
    assign layer2_outputs[1562] = (layer1_outputs[242]) & ~(layer1_outputs[2940]);
    assign layer2_outputs[1563] = (layer1_outputs[466]) & (layer1_outputs[5073]);
    assign layer2_outputs[1564] = layer1_outputs[1444];
    assign layer2_outputs[1565] = 1'b0;
    assign layer2_outputs[1566] = ~(layer1_outputs[532]);
    assign layer2_outputs[1567] = layer1_outputs[2898];
    assign layer2_outputs[1568] = layer1_outputs[533];
    assign layer2_outputs[1569] = (layer1_outputs[937]) & (layer1_outputs[1274]);
    assign layer2_outputs[1570] = ~(layer1_outputs[4096]) | (layer1_outputs[4755]);
    assign layer2_outputs[1571] = ~(layer1_outputs[3185]);
    assign layer2_outputs[1572] = ~(layer1_outputs[1377]);
    assign layer2_outputs[1573] = layer1_outputs[3430];
    assign layer2_outputs[1574] = ~(layer1_outputs[369]) | (layer1_outputs[669]);
    assign layer2_outputs[1575] = ~(layer1_outputs[1304]);
    assign layer2_outputs[1576] = 1'b1;
    assign layer2_outputs[1577] = layer1_outputs[1984];
    assign layer2_outputs[1578] = layer1_outputs[1234];
    assign layer2_outputs[1579] = layer1_outputs[5075];
    assign layer2_outputs[1580] = 1'b1;
    assign layer2_outputs[1581] = ~(layer1_outputs[1802]) | (layer1_outputs[3766]);
    assign layer2_outputs[1582] = ~(layer1_outputs[2726]);
    assign layer2_outputs[1583] = ~((layer1_outputs[4017]) & (layer1_outputs[2751]));
    assign layer2_outputs[1584] = layer1_outputs[96];
    assign layer2_outputs[1585] = layer1_outputs[4458];
    assign layer2_outputs[1586] = ~(layer1_outputs[4116]) | (layer1_outputs[4856]);
    assign layer2_outputs[1587] = ~((layer1_outputs[4712]) | (layer1_outputs[1552]));
    assign layer2_outputs[1588] = layer1_outputs[2302];
    assign layer2_outputs[1589] = (layer1_outputs[3600]) & (layer1_outputs[3765]);
    assign layer2_outputs[1590] = layer1_outputs[3579];
    assign layer2_outputs[1591] = ~((layer1_outputs[2709]) | (layer1_outputs[589]));
    assign layer2_outputs[1592] = ~(layer1_outputs[2432]) | (layer1_outputs[1562]);
    assign layer2_outputs[1593] = ~(layer1_outputs[3353]);
    assign layer2_outputs[1594] = ~(layer1_outputs[3956]) | (layer1_outputs[4451]);
    assign layer2_outputs[1595] = 1'b0;
    assign layer2_outputs[1596] = layer1_outputs[2128];
    assign layer2_outputs[1597] = layer1_outputs[1519];
    assign layer2_outputs[1598] = layer1_outputs[704];
    assign layer2_outputs[1599] = ~(layer1_outputs[1511]);
    assign layer2_outputs[1600] = 1'b0;
    assign layer2_outputs[1601] = ~(layer1_outputs[2332]);
    assign layer2_outputs[1602] = 1'b0;
    assign layer2_outputs[1603] = layer1_outputs[1505];
    assign layer2_outputs[1604] = (layer1_outputs[387]) ^ (layer1_outputs[247]);
    assign layer2_outputs[1605] = (layer1_outputs[3494]) | (layer1_outputs[209]);
    assign layer2_outputs[1606] = (layer1_outputs[3]) | (layer1_outputs[116]);
    assign layer2_outputs[1607] = ~(layer1_outputs[3101]);
    assign layer2_outputs[1608] = ~((layer1_outputs[4397]) | (layer1_outputs[4600]));
    assign layer2_outputs[1609] = ~(layer1_outputs[2359]) | (layer1_outputs[2356]);
    assign layer2_outputs[1610] = ~(layer1_outputs[324]) | (layer1_outputs[2387]);
    assign layer2_outputs[1611] = layer1_outputs[5025];
    assign layer2_outputs[1612] = ~(layer1_outputs[1838]) | (layer1_outputs[652]);
    assign layer2_outputs[1613] = ~(layer1_outputs[963]) | (layer1_outputs[3723]);
    assign layer2_outputs[1614] = 1'b0;
    assign layer2_outputs[1615] = (layer1_outputs[359]) | (layer1_outputs[1144]);
    assign layer2_outputs[1616] = (layer1_outputs[871]) ^ (layer1_outputs[2333]);
    assign layer2_outputs[1617] = 1'b0;
    assign layer2_outputs[1618] = (layer1_outputs[2845]) & ~(layer1_outputs[4203]);
    assign layer2_outputs[1619] = (layer1_outputs[3632]) ^ (layer1_outputs[1994]);
    assign layer2_outputs[1620] = (layer1_outputs[1540]) & ~(layer1_outputs[2144]);
    assign layer2_outputs[1621] = (layer1_outputs[4245]) | (layer1_outputs[4291]);
    assign layer2_outputs[1622] = (layer1_outputs[4587]) & ~(layer1_outputs[26]);
    assign layer2_outputs[1623] = ~(layer1_outputs[4617]) | (layer1_outputs[1603]);
    assign layer2_outputs[1624] = (layer1_outputs[2882]) | (layer1_outputs[432]);
    assign layer2_outputs[1625] = layer1_outputs[1477];
    assign layer2_outputs[1626] = (layer1_outputs[4770]) & ~(layer1_outputs[327]);
    assign layer2_outputs[1627] = ~((layer1_outputs[4246]) | (layer1_outputs[3432]));
    assign layer2_outputs[1628] = 1'b0;
    assign layer2_outputs[1629] = ~(layer1_outputs[902]);
    assign layer2_outputs[1630] = ~(layer1_outputs[4485]) | (layer1_outputs[1011]);
    assign layer2_outputs[1631] = (layer1_outputs[4949]) & ~(layer1_outputs[2794]);
    assign layer2_outputs[1632] = ~(layer1_outputs[2962]);
    assign layer2_outputs[1633] = ~((layer1_outputs[3252]) | (layer1_outputs[377]));
    assign layer2_outputs[1634] = ~(layer1_outputs[2738]) | (layer1_outputs[1185]);
    assign layer2_outputs[1635] = (layer1_outputs[3289]) & (layer1_outputs[649]);
    assign layer2_outputs[1636] = ~(layer1_outputs[1796]);
    assign layer2_outputs[1637] = 1'b1;
    assign layer2_outputs[1638] = 1'b0;
    assign layer2_outputs[1639] = ~((layer1_outputs[3551]) | (layer1_outputs[5107]));
    assign layer2_outputs[1640] = ~(layer1_outputs[1805]) | (layer1_outputs[2264]);
    assign layer2_outputs[1641] = 1'b0;
    assign layer2_outputs[1642] = ~(layer1_outputs[3066]);
    assign layer2_outputs[1643] = (layer1_outputs[1185]) | (layer1_outputs[1841]);
    assign layer2_outputs[1644] = layer1_outputs[3736];
    assign layer2_outputs[1645] = 1'b1;
    assign layer2_outputs[1646] = 1'b1;
    assign layer2_outputs[1647] = (layer1_outputs[4127]) & (layer1_outputs[4857]);
    assign layer2_outputs[1648] = layer1_outputs[2021];
    assign layer2_outputs[1649] = ~((layer1_outputs[2880]) & (layer1_outputs[877]));
    assign layer2_outputs[1650] = (layer1_outputs[2909]) & ~(layer1_outputs[1542]);
    assign layer2_outputs[1651] = 1'b0;
    assign layer2_outputs[1652] = (layer1_outputs[176]) & (layer1_outputs[1727]);
    assign layer2_outputs[1653] = ~(layer1_outputs[3257]);
    assign layer2_outputs[1654] = ~((layer1_outputs[1154]) | (layer1_outputs[1973]));
    assign layer2_outputs[1655] = ~(layer1_outputs[3060]) | (layer1_outputs[3710]);
    assign layer2_outputs[1656] = (layer1_outputs[914]) | (layer1_outputs[504]);
    assign layer2_outputs[1657] = (layer1_outputs[2992]) | (layer1_outputs[4435]);
    assign layer2_outputs[1658] = layer1_outputs[5095];
    assign layer2_outputs[1659] = (layer1_outputs[2838]) ^ (layer1_outputs[2758]);
    assign layer2_outputs[1660] = ~((layer1_outputs[4509]) | (layer1_outputs[4550]));
    assign layer2_outputs[1661] = ~(layer1_outputs[1345]);
    assign layer2_outputs[1662] = (layer1_outputs[751]) & ~(layer1_outputs[3473]);
    assign layer2_outputs[1663] = (layer1_outputs[301]) & ~(layer1_outputs[1492]);
    assign layer2_outputs[1664] = 1'b0;
    assign layer2_outputs[1665] = 1'b1;
    assign layer2_outputs[1666] = layer1_outputs[3882];
    assign layer2_outputs[1667] = ~(layer1_outputs[3444]);
    assign layer2_outputs[1668] = ~(layer1_outputs[4701]) | (layer1_outputs[2286]);
    assign layer2_outputs[1669] = layer1_outputs[3404];
    assign layer2_outputs[1670] = 1'b1;
    assign layer2_outputs[1671] = ~((layer1_outputs[419]) | (layer1_outputs[3029]));
    assign layer2_outputs[1672] = ~(layer1_outputs[3909]);
    assign layer2_outputs[1673] = (layer1_outputs[3634]) | (layer1_outputs[623]);
    assign layer2_outputs[1674] = (layer1_outputs[1019]) & (layer1_outputs[113]);
    assign layer2_outputs[1675] = 1'b0;
    assign layer2_outputs[1676] = ~(layer1_outputs[4590]) | (layer1_outputs[1674]);
    assign layer2_outputs[1677] = ~((layer1_outputs[3053]) | (layer1_outputs[2908]));
    assign layer2_outputs[1678] = ~(layer1_outputs[3731]) | (layer1_outputs[461]);
    assign layer2_outputs[1679] = (layer1_outputs[2518]) & ~(layer1_outputs[3672]);
    assign layer2_outputs[1680] = ~(layer1_outputs[4463]);
    assign layer2_outputs[1681] = (layer1_outputs[2889]) | (layer1_outputs[4424]);
    assign layer2_outputs[1682] = ~(layer1_outputs[3775]) | (layer1_outputs[2964]);
    assign layer2_outputs[1683] = layer1_outputs[3649];
    assign layer2_outputs[1684] = ~(layer1_outputs[2520]);
    assign layer2_outputs[1685] = ~(layer1_outputs[4285]);
    assign layer2_outputs[1686] = ~((layer1_outputs[2093]) & (layer1_outputs[1471]));
    assign layer2_outputs[1687] = layer1_outputs[3010];
    assign layer2_outputs[1688] = ~((layer1_outputs[1988]) & (layer1_outputs[3206]));
    assign layer2_outputs[1689] = ~(layer1_outputs[3164]) | (layer1_outputs[1070]);
    assign layer2_outputs[1690] = (layer1_outputs[4419]) & ~(layer1_outputs[3779]);
    assign layer2_outputs[1691] = ~(layer1_outputs[840]);
    assign layer2_outputs[1692] = (layer1_outputs[2529]) & ~(layer1_outputs[2458]);
    assign layer2_outputs[1693] = (layer1_outputs[836]) & ~(layer1_outputs[797]);
    assign layer2_outputs[1694] = (layer1_outputs[3099]) & ~(layer1_outputs[4796]);
    assign layer2_outputs[1695] = ~(layer1_outputs[3260]) | (layer1_outputs[1391]);
    assign layer2_outputs[1696] = ~((layer1_outputs[1510]) ^ (layer1_outputs[2176]));
    assign layer2_outputs[1697] = 1'b1;
    assign layer2_outputs[1698] = ~(layer1_outputs[4994]) | (layer1_outputs[474]);
    assign layer2_outputs[1699] = ~(layer1_outputs[538]);
    assign layer2_outputs[1700] = (layer1_outputs[426]) | (layer1_outputs[2883]);
    assign layer2_outputs[1701] = 1'b1;
    assign layer2_outputs[1702] = ~(layer1_outputs[2667]) | (layer1_outputs[3195]);
    assign layer2_outputs[1703] = ~(layer1_outputs[1449]) | (layer1_outputs[3829]);
    assign layer2_outputs[1704] = ~(layer1_outputs[1193]) | (layer1_outputs[2900]);
    assign layer2_outputs[1705] = (layer1_outputs[4177]) & ~(layer1_outputs[5041]);
    assign layer2_outputs[1706] = ~(layer1_outputs[1304]);
    assign layer2_outputs[1707] = ~(layer1_outputs[4093]) | (layer1_outputs[3445]);
    assign layer2_outputs[1708] = ~(layer1_outputs[2943]) | (layer1_outputs[3767]);
    assign layer2_outputs[1709] = ~(layer1_outputs[3704]) | (layer1_outputs[3838]);
    assign layer2_outputs[1710] = (layer1_outputs[1890]) & (layer1_outputs[3640]);
    assign layer2_outputs[1711] = ~(layer1_outputs[389]);
    assign layer2_outputs[1712] = ~(layer1_outputs[3572]) | (layer1_outputs[4721]);
    assign layer2_outputs[1713] = 1'b0;
    assign layer2_outputs[1714] = 1'b0;
    assign layer2_outputs[1715] = ~(layer1_outputs[173]);
    assign layer2_outputs[1716] = 1'b1;
    assign layer2_outputs[1717] = layer1_outputs[4375];
    assign layer2_outputs[1718] = ~(layer1_outputs[3680]);
    assign layer2_outputs[1719] = (layer1_outputs[496]) & ~(layer1_outputs[338]);
    assign layer2_outputs[1720] = (layer1_outputs[506]) | (layer1_outputs[4823]);
    assign layer2_outputs[1721] = ~(layer1_outputs[450]) | (layer1_outputs[116]);
    assign layer2_outputs[1722] = 1'b1;
    assign layer2_outputs[1723] = layer1_outputs[4212];
    assign layer2_outputs[1724] = 1'b1;
    assign layer2_outputs[1725] = (layer1_outputs[3518]) & (layer1_outputs[1978]);
    assign layer2_outputs[1726] = ~((layer1_outputs[3978]) | (layer1_outputs[1368]));
    assign layer2_outputs[1727] = ~(layer1_outputs[1430]);
    assign layer2_outputs[1728] = (layer1_outputs[1177]) & ~(layer1_outputs[1201]);
    assign layer2_outputs[1729] = ~(layer1_outputs[621]);
    assign layer2_outputs[1730] = (layer1_outputs[4366]) & ~(layer1_outputs[2984]);
    assign layer2_outputs[1731] = ~((layer1_outputs[3903]) | (layer1_outputs[1607]));
    assign layer2_outputs[1732] = (layer1_outputs[3843]) & ~(layer1_outputs[1524]);
    assign layer2_outputs[1733] = (layer1_outputs[2883]) | (layer1_outputs[3558]);
    assign layer2_outputs[1734] = 1'b1;
    assign layer2_outputs[1735] = (layer1_outputs[3331]) & ~(layer1_outputs[19]);
    assign layer2_outputs[1736] = ~((layer1_outputs[2037]) | (layer1_outputs[2233]));
    assign layer2_outputs[1737] = 1'b0;
    assign layer2_outputs[1738] = 1'b0;
    assign layer2_outputs[1739] = 1'b1;
    assign layer2_outputs[1740] = 1'b0;
    assign layer2_outputs[1741] = 1'b0;
    assign layer2_outputs[1742] = ~(layer1_outputs[4861]) | (layer1_outputs[4353]);
    assign layer2_outputs[1743] = ~(layer1_outputs[555]);
    assign layer2_outputs[1744] = layer1_outputs[1761];
    assign layer2_outputs[1745] = ~((layer1_outputs[3372]) ^ (layer1_outputs[52]));
    assign layer2_outputs[1746] = (layer1_outputs[1718]) & (layer1_outputs[4426]);
    assign layer2_outputs[1747] = layer1_outputs[2754];
    assign layer2_outputs[1748] = layer1_outputs[1621];
    assign layer2_outputs[1749] = (layer1_outputs[2460]) | (layer1_outputs[1961]);
    assign layer2_outputs[1750] = layer1_outputs[986];
    assign layer2_outputs[1751] = (layer1_outputs[4876]) & (layer1_outputs[3160]);
    assign layer2_outputs[1752] = ~(layer1_outputs[2063]);
    assign layer2_outputs[1753] = ~((layer1_outputs[310]) | (layer1_outputs[2157]));
    assign layer2_outputs[1754] = (layer1_outputs[198]) & ~(layer1_outputs[744]);
    assign layer2_outputs[1755] = ~((layer1_outputs[2694]) ^ (layer1_outputs[4953]));
    assign layer2_outputs[1756] = ~(layer1_outputs[2340]) | (layer1_outputs[3925]);
    assign layer2_outputs[1757] = ~(layer1_outputs[2561]) | (layer1_outputs[811]);
    assign layer2_outputs[1758] = ~((layer1_outputs[5065]) & (layer1_outputs[3378]));
    assign layer2_outputs[1759] = ~(layer1_outputs[2454]);
    assign layer2_outputs[1760] = (layer1_outputs[61]) & ~(layer1_outputs[4655]);
    assign layer2_outputs[1761] = layer1_outputs[3073];
    assign layer2_outputs[1762] = (layer1_outputs[4951]) & ~(layer1_outputs[4665]);
    assign layer2_outputs[1763] = ~(layer1_outputs[1568]) | (layer1_outputs[2278]);
    assign layer2_outputs[1764] = (layer1_outputs[2594]) & (layer1_outputs[125]);
    assign layer2_outputs[1765] = 1'b1;
    assign layer2_outputs[1766] = ~(layer1_outputs[2528]) | (layer1_outputs[303]);
    assign layer2_outputs[1767] = (layer1_outputs[1408]) & ~(layer1_outputs[3384]);
    assign layer2_outputs[1768] = ~(layer1_outputs[2556]) | (layer1_outputs[3132]);
    assign layer2_outputs[1769] = ~(layer1_outputs[1105]);
    assign layer2_outputs[1770] = 1'b0;
    assign layer2_outputs[1771] = ~(layer1_outputs[5001]) | (layer1_outputs[3999]);
    assign layer2_outputs[1772] = (layer1_outputs[4483]) & ~(layer1_outputs[518]);
    assign layer2_outputs[1773] = 1'b0;
    assign layer2_outputs[1774] = ~(layer1_outputs[5100]);
    assign layer2_outputs[1775] = (layer1_outputs[3918]) & ~(layer1_outputs[4930]);
    assign layer2_outputs[1776] = (layer1_outputs[1294]) & ~(layer1_outputs[2577]);
    assign layer2_outputs[1777] = layer1_outputs[1992];
    assign layer2_outputs[1778] = (layer1_outputs[2607]) & (layer1_outputs[4080]);
    assign layer2_outputs[1779] = (layer1_outputs[2467]) | (layer1_outputs[4412]);
    assign layer2_outputs[1780] = 1'b0;
    assign layer2_outputs[1781] = ~((layer1_outputs[3087]) | (layer1_outputs[2383]));
    assign layer2_outputs[1782] = (layer1_outputs[787]) ^ (layer1_outputs[2269]);
    assign layer2_outputs[1783] = (layer1_outputs[3109]) & ~(layer1_outputs[4772]);
    assign layer2_outputs[1784] = 1'b0;
    assign layer2_outputs[1785] = (layer1_outputs[3336]) & ~(layer1_outputs[1865]);
    assign layer2_outputs[1786] = (layer1_outputs[302]) | (layer1_outputs[4367]);
    assign layer2_outputs[1787] = (layer1_outputs[802]) | (layer1_outputs[1896]);
    assign layer2_outputs[1788] = (layer1_outputs[1798]) & (layer1_outputs[107]);
    assign layer2_outputs[1789] = (layer1_outputs[1729]) & ~(layer1_outputs[3802]);
    assign layer2_outputs[1790] = ~(layer1_outputs[3587]);
    assign layer2_outputs[1791] = ~(layer1_outputs[1357]);
    assign layer2_outputs[1792] = 1'b1;
    assign layer2_outputs[1793] = 1'b0;
    assign layer2_outputs[1794] = layer1_outputs[2192];
    assign layer2_outputs[1795] = (layer1_outputs[2012]) & ~(layer1_outputs[1776]);
    assign layer2_outputs[1796] = ~((layer1_outputs[2844]) | (layer1_outputs[5079]));
    assign layer2_outputs[1797] = ~((layer1_outputs[4331]) | (layer1_outputs[4161]));
    assign layer2_outputs[1798] = ~(layer1_outputs[1264]) | (layer1_outputs[4002]);
    assign layer2_outputs[1799] = (layer1_outputs[4698]) | (layer1_outputs[4176]);
    assign layer2_outputs[1800] = ~(layer1_outputs[1218]) | (layer1_outputs[3896]);
    assign layer2_outputs[1801] = 1'b0;
    assign layer2_outputs[1802] = ~(layer1_outputs[135]) | (layer1_outputs[3542]);
    assign layer2_outputs[1803] = 1'b1;
    assign layer2_outputs[1804] = layer1_outputs[989];
    assign layer2_outputs[1805] = ~(layer1_outputs[3738]) | (layer1_outputs[4637]);
    assign layer2_outputs[1806] = layer1_outputs[3856];
    assign layer2_outputs[1807] = ~(layer1_outputs[4858]);
    assign layer2_outputs[1808] = (layer1_outputs[2619]) & (layer1_outputs[137]);
    assign layer2_outputs[1809] = layer1_outputs[3151];
    assign layer2_outputs[1810] = layer1_outputs[3073];
    assign layer2_outputs[1811] = 1'b1;
    assign layer2_outputs[1812] = 1'b0;
    assign layer2_outputs[1813] = 1'b0;
    assign layer2_outputs[1814] = 1'b0;
    assign layer2_outputs[1815] = layer1_outputs[1835];
    assign layer2_outputs[1816] = (layer1_outputs[3767]) & (layer1_outputs[1822]);
    assign layer2_outputs[1817] = 1'b1;
    assign layer2_outputs[1818] = ~(layer1_outputs[2309]);
    assign layer2_outputs[1819] = ~((layer1_outputs[537]) | (layer1_outputs[774]));
    assign layer2_outputs[1820] = ~((layer1_outputs[1990]) | (layer1_outputs[4097]));
    assign layer2_outputs[1821] = layer1_outputs[3636];
    assign layer2_outputs[1822] = 1'b1;
    assign layer2_outputs[1823] = ~(layer1_outputs[1270]);
    assign layer2_outputs[1824] = (layer1_outputs[3942]) & (layer1_outputs[4899]);
    assign layer2_outputs[1825] = layer1_outputs[3419];
    assign layer2_outputs[1826] = 1'b0;
    assign layer2_outputs[1827] = ~((layer1_outputs[2303]) ^ (layer1_outputs[820]));
    assign layer2_outputs[1828] = ~(layer1_outputs[1761]);
    assign layer2_outputs[1829] = ~(layer1_outputs[1590]) | (layer1_outputs[2798]);
    assign layer2_outputs[1830] = layer1_outputs[324];
    assign layer2_outputs[1831] = (layer1_outputs[1764]) ^ (layer1_outputs[4516]);
    assign layer2_outputs[1832] = ~(layer1_outputs[1508]);
    assign layer2_outputs[1833] = ~(layer1_outputs[1887]) | (layer1_outputs[3410]);
    assign layer2_outputs[1834] = ~(layer1_outputs[1177]) | (layer1_outputs[3013]);
    assign layer2_outputs[1835] = (layer1_outputs[4343]) & (layer1_outputs[3119]);
    assign layer2_outputs[1836] = ~(layer1_outputs[168]) | (layer1_outputs[4283]);
    assign layer2_outputs[1837] = ~((layer1_outputs[4619]) | (layer1_outputs[4767]));
    assign layer2_outputs[1838] = (layer1_outputs[4226]) & (layer1_outputs[1891]);
    assign layer2_outputs[1839] = ~(layer1_outputs[4164]) | (layer1_outputs[2260]);
    assign layer2_outputs[1840] = layer1_outputs[1641];
    assign layer2_outputs[1841] = (layer1_outputs[5074]) | (layer1_outputs[3378]);
    assign layer2_outputs[1842] = ~(layer1_outputs[2422]);
    assign layer2_outputs[1843] = layer1_outputs[1417];
    assign layer2_outputs[1844] = layer1_outputs[1690];
    assign layer2_outputs[1845] = ~(layer1_outputs[5099]);
    assign layer2_outputs[1846] = 1'b0;
    assign layer2_outputs[1847] = ~(layer1_outputs[174]) | (layer1_outputs[2395]);
    assign layer2_outputs[1848] = ~(layer1_outputs[3028]);
    assign layer2_outputs[1849] = ~(layer1_outputs[2347]) | (layer1_outputs[4376]);
    assign layer2_outputs[1850] = layer1_outputs[1863];
    assign layer2_outputs[1851] = ~((layer1_outputs[1777]) | (layer1_outputs[4390]));
    assign layer2_outputs[1852] = (layer1_outputs[1256]) & (layer1_outputs[4860]);
    assign layer2_outputs[1853] = layer1_outputs[3994];
    assign layer2_outputs[1854] = layer1_outputs[4987];
    assign layer2_outputs[1855] = ~(layer1_outputs[1329]);
    assign layer2_outputs[1856] = ~(layer1_outputs[846]);
    assign layer2_outputs[1857] = (layer1_outputs[2718]) | (layer1_outputs[1699]);
    assign layer2_outputs[1858] = ~(layer1_outputs[2491]);
    assign layer2_outputs[1859] = (layer1_outputs[4819]) | (layer1_outputs[2397]);
    assign layer2_outputs[1860] = ~(layer1_outputs[4820]);
    assign layer2_outputs[1861] = (layer1_outputs[3478]) & ~(layer1_outputs[776]);
    assign layer2_outputs[1862] = ~(layer1_outputs[584]);
    assign layer2_outputs[1863] = ~(layer1_outputs[74]);
    assign layer2_outputs[1864] = ~(layer1_outputs[1298]) | (layer1_outputs[1184]);
    assign layer2_outputs[1865] = ~(layer1_outputs[2473]);
    assign layer2_outputs[1866] = (layer1_outputs[297]) | (layer1_outputs[2542]);
    assign layer2_outputs[1867] = ~(layer1_outputs[2142]) | (layer1_outputs[3433]);
    assign layer2_outputs[1868] = ~((layer1_outputs[227]) & (layer1_outputs[5023]));
    assign layer2_outputs[1869] = ~(layer1_outputs[3162]);
    assign layer2_outputs[1870] = (layer1_outputs[2768]) & ~(layer1_outputs[4357]);
    assign layer2_outputs[1871] = layer1_outputs[4647];
    assign layer2_outputs[1872] = 1'b1;
    assign layer2_outputs[1873] = layer1_outputs[175];
    assign layer2_outputs[1874] = ~((layer1_outputs[516]) ^ (layer1_outputs[2659]));
    assign layer2_outputs[1875] = ~(layer1_outputs[1531]);
    assign layer2_outputs[1876] = (layer1_outputs[4205]) & (layer1_outputs[2623]);
    assign layer2_outputs[1877] = (layer1_outputs[242]) & ~(layer1_outputs[964]);
    assign layer2_outputs[1878] = (layer1_outputs[3703]) | (layer1_outputs[374]);
    assign layer2_outputs[1879] = layer1_outputs[991];
    assign layer2_outputs[1880] = ~(layer1_outputs[822]) | (layer1_outputs[4502]);
    assign layer2_outputs[1881] = ~((layer1_outputs[956]) & (layer1_outputs[4296]));
    assign layer2_outputs[1882] = (layer1_outputs[1958]) & (layer1_outputs[32]);
    assign layer2_outputs[1883] = (layer1_outputs[4616]) & ~(layer1_outputs[2805]);
    assign layer2_outputs[1884] = layer1_outputs[4355];
    assign layer2_outputs[1885] = layer1_outputs[4648];
    assign layer2_outputs[1886] = layer1_outputs[1032];
    assign layer2_outputs[1887] = (layer1_outputs[1704]) & (layer1_outputs[265]);
    assign layer2_outputs[1888] = (layer1_outputs[2390]) | (layer1_outputs[1594]);
    assign layer2_outputs[1889] = (layer1_outputs[4786]) & (layer1_outputs[501]);
    assign layer2_outputs[1890] = ~(layer1_outputs[1880]);
    assign layer2_outputs[1891] = ~(layer1_outputs[4215]) | (layer1_outputs[3238]);
    assign layer2_outputs[1892] = ~((layer1_outputs[2399]) | (layer1_outputs[2609]));
    assign layer2_outputs[1893] = ~(layer1_outputs[2673]);
    assign layer2_outputs[1894] = 1'b1;
    assign layer2_outputs[1895] = ~(layer1_outputs[2523]);
    assign layer2_outputs[1896] = (layer1_outputs[350]) & ~(layer1_outputs[3650]);
    assign layer2_outputs[1897] = (layer1_outputs[1809]) & ~(layer1_outputs[28]);
    assign layer2_outputs[1898] = (layer1_outputs[2033]) & ~(layer1_outputs[2802]);
    assign layer2_outputs[1899] = ~(layer1_outputs[3465]) | (layer1_outputs[1687]);
    assign layer2_outputs[1900] = ~(layer1_outputs[2807]) | (layer1_outputs[2120]);
    assign layer2_outputs[1901] = (layer1_outputs[2479]) & ~(layer1_outputs[3005]);
    assign layer2_outputs[1902] = layer1_outputs[3972];
    assign layer2_outputs[1903] = (layer1_outputs[3331]) & ~(layer1_outputs[105]);
    assign layer2_outputs[1904] = 1'b0;
    assign layer2_outputs[1905] = 1'b0;
    assign layer2_outputs[1906] = ~(layer1_outputs[4160]) | (layer1_outputs[631]);
    assign layer2_outputs[1907] = 1'b1;
    assign layer2_outputs[1908] = 1'b0;
    assign layer2_outputs[1909] = layer1_outputs[2183];
    assign layer2_outputs[1910] = ~((layer1_outputs[3634]) | (layer1_outputs[3161]));
    assign layer2_outputs[1911] = (layer1_outputs[677]) | (layer1_outputs[4118]);
    assign layer2_outputs[1912] = (layer1_outputs[1889]) & ~(layer1_outputs[3462]);
    assign layer2_outputs[1913] = (layer1_outputs[3758]) | (layer1_outputs[1144]);
    assign layer2_outputs[1914] = (layer1_outputs[1697]) ^ (layer1_outputs[2599]);
    assign layer2_outputs[1915] = ~(layer1_outputs[2739]);
    assign layer2_outputs[1916] = (layer1_outputs[4715]) ^ (layer1_outputs[1161]);
    assign layer2_outputs[1917] = ~(layer1_outputs[704]);
    assign layer2_outputs[1918] = (layer1_outputs[703]) & ~(layer1_outputs[5079]);
    assign layer2_outputs[1919] = ~((layer1_outputs[511]) & (layer1_outputs[2374]));
    assign layer2_outputs[1920] = layer1_outputs[2600];
    assign layer2_outputs[1921] = (layer1_outputs[3677]) ^ (layer1_outputs[3117]);
    assign layer2_outputs[1922] = ~(layer1_outputs[4665]);
    assign layer2_outputs[1923] = ~(layer1_outputs[186]);
    assign layer2_outputs[1924] = layer1_outputs[274];
    assign layer2_outputs[1925] = ~(layer1_outputs[1246]);
    assign layer2_outputs[1926] = ~(layer1_outputs[1069]) | (layer1_outputs[1845]);
    assign layer2_outputs[1927] = ~((layer1_outputs[5116]) ^ (layer1_outputs[4638]));
    assign layer2_outputs[1928] = layer1_outputs[1096];
    assign layer2_outputs[1929] = (layer1_outputs[401]) | (layer1_outputs[2205]);
    assign layer2_outputs[1930] = (layer1_outputs[4395]) & ~(layer1_outputs[199]);
    assign layer2_outputs[1931] = (layer1_outputs[3008]) & ~(layer1_outputs[4347]);
    assign layer2_outputs[1932] = ~(layer1_outputs[1086]) | (layer1_outputs[2067]);
    assign layer2_outputs[1933] = ~((layer1_outputs[2362]) & (layer1_outputs[4015]));
    assign layer2_outputs[1934] = 1'b1;
    assign layer2_outputs[1935] = layer1_outputs[2226];
    assign layer2_outputs[1936] = 1'b1;
    assign layer2_outputs[1937] = (layer1_outputs[2945]) ^ (layer1_outputs[3540]);
    assign layer2_outputs[1938] = layer1_outputs[4587];
    assign layer2_outputs[1939] = layer1_outputs[1928];
    assign layer2_outputs[1940] = 1'b1;
    assign layer2_outputs[1941] = ~(layer1_outputs[3528]) | (layer1_outputs[5099]);
    assign layer2_outputs[1942] = 1'b1;
    assign layer2_outputs[1943] = layer1_outputs[20];
    assign layer2_outputs[1944] = 1'b1;
    assign layer2_outputs[1945] = ~(layer1_outputs[2058]);
    assign layer2_outputs[1946] = 1'b1;
    assign layer2_outputs[1947] = (layer1_outputs[289]) & (layer1_outputs[2214]);
    assign layer2_outputs[1948] = (layer1_outputs[184]) | (layer1_outputs[1886]);
    assign layer2_outputs[1949] = ~(layer1_outputs[873]) | (layer1_outputs[1953]);
    assign layer2_outputs[1950] = 1'b1;
    assign layer2_outputs[1951] = (layer1_outputs[4768]) & ~(layer1_outputs[3897]);
    assign layer2_outputs[1952] = 1'b0;
    assign layer2_outputs[1953] = 1'b1;
    assign layer2_outputs[1954] = ~((layer1_outputs[1491]) & (layer1_outputs[5067]));
    assign layer2_outputs[1955] = (layer1_outputs[2296]) | (layer1_outputs[3790]);
    assign layer2_outputs[1956] = ~(layer1_outputs[2793]);
    assign layer2_outputs[1957] = layer1_outputs[1682];
    assign layer2_outputs[1958] = (layer1_outputs[2184]) ^ (layer1_outputs[443]);
    assign layer2_outputs[1959] = (layer1_outputs[1561]) & ~(layer1_outputs[4489]);
    assign layer2_outputs[1960] = layer1_outputs[1839];
    assign layer2_outputs[1961] = ~(layer1_outputs[4735]);
    assign layer2_outputs[1962] = layer1_outputs[2610];
    assign layer2_outputs[1963] = 1'b1;
    assign layer2_outputs[1964] = ~((layer1_outputs[4763]) & (layer1_outputs[123]));
    assign layer2_outputs[1965] = ~(layer1_outputs[4472]) | (layer1_outputs[3864]);
    assign layer2_outputs[1966] = ~(layer1_outputs[2919]);
    assign layer2_outputs[1967] = (layer1_outputs[1709]) & (layer1_outputs[3503]);
    assign layer2_outputs[1968] = (layer1_outputs[4389]) & (layer1_outputs[4716]);
    assign layer2_outputs[1969] = layer1_outputs[1321];
    assign layer2_outputs[1970] = layer1_outputs[789];
    assign layer2_outputs[1971] = ~(layer1_outputs[1807]);
    assign layer2_outputs[1972] = ~(layer1_outputs[3639]) | (layer1_outputs[826]);
    assign layer2_outputs[1973] = ~(layer1_outputs[3460]);
    assign layer2_outputs[1974] = (layer1_outputs[2485]) & ~(layer1_outputs[2322]);
    assign layer2_outputs[1975] = ~((layer1_outputs[142]) & (layer1_outputs[3773]));
    assign layer2_outputs[1976] = (layer1_outputs[1912]) | (layer1_outputs[67]);
    assign layer2_outputs[1977] = 1'b0;
    assign layer2_outputs[1978] = 1'b0;
    assign layer2_outputs[1979] = ~(layer1_outputs[559]);
    assign layer2_outputs[1980] = layer1_outputs[3836];
    assign layer2_outputs[1981] = ~(layer1_outputs[3359]);
    assign layer2_outputs[1982] = 1'b0;
    assign layer2_outputs[1983] = ~((layer1_outputs[4704]) | (layer1_outputs[3408]));
    assign layer2_outputs[1984] = ~((layer1_outputs[2244]) | (layer1_outputs[407]));
    assign layer2_outputs[1985] = 1'b1;
    assign layer2_outputs[1986] = layer1_outputs[1356];
    assign layer2_outputs[1987] = (layer1_outputs[5002]) & ~(layer1_outputs[1824]);
    assign layer2_outputs[1988] = ~((layer1_outputs[3737]) | (layer1_outputs[4966]));
    assign layer2_outputs[1989] = ~(layer1_outputs[2918]);
    assign layer2_outputs[1990] = (layer1_outputs[3762]) | (layer1_outputs[1716]);
    assign layer2_outputs[1991] = ~(layer1_outputs[3666]) | (layer1_outputs[4253]);
    assign layer2_outputs[1992] = (layer1_outputs[4871]) | (layer1_outputs[2034]);
    assign layer2_outputs[1993] = layer1_outputs[2875];
    assign layer2_outputs[1994] = (layer1_outputs[3856]) & ~(layer1_outputs[2820]);
    assign layer2_outputs[1995] = ~(layer1_outputs[2603]) | (layer1_outputs[4504]);
    assign layer2_outputs[1996] = (layer1_outputs[257]) & ~(layer1_outputs[4432]);
    assign layer2_outputs[1997] = ~(layer1_outputs[2931]);
    assign layer2_outputs[1998] = layer1_outputs[4539];
    assign layer2_outputs[1999] = ~(layer1_outputs[314]);
    assign layer2_outputs[2000] = ~((layer1_outputs[977]) & (layer1_outputs[2433]));
    assign layer2_outputs[2001] = ~(layer1_outputs[4228]);
    assign layer2_outputs[2002] = layer1_outputs[3780];
    assign layer2_outputs[2003] = ~(layer1_outputs[1672]) | (layer1_outputs[757]);
    assign layer2_outputs[2004] = layer1_outputs[4386];
    assign layer2_outputs[2005] = (layer1_outputs[4777]) | (layer1_outputs[2009]);
    assign layer2_outputs[2006] = layer1_outputs[3945];
    assign layer2_outputs[2007] = (layer1_outputs[3971]) | (layer1_outputs[4835]);
    assign layer2_outputs[2008] = ~((layer1_outputs[1139]) | (layer1_outputs[2761]));
    assign layer2_outputs[2009] = 1'b1;
    assign layer2_outputs[2010] = (layer1_outputs[3948]) & (layer1_outputs[2237]);
    assign layer2_outputs[2011] = 1'b1;
    assign layer2_outputs[2012] = 1'b0;
    assign layer2_outputs[2013] = ~(layer1_outputs[3727]);
    assign layer2_outputs[2014] = (layer1_outputs[3739]) & (layer1_outputs[523]);
    assign layer2_outputs[2015] = (layer1_outputs[604]) ^ (layer1_outputs[1828]);
    assign layer2_outputs[2016] = (layer1_outputs[571]) | (layer1_outputs[4906]);
    assign layer2_outputs[2017] = (layer1_outputs[490]) & (layer1_outputs[4409]);
    assign layer2_outputs[2018] = (layer1_outputs[4773]) & ~(layer1_outputs[2753]);
    assign layer2_outputs[2019] = ~(layer1_outputs[2160]) | (layer1_outputs[4608]);
    assign layer2_outputs[2020] = 1'b0;
    assign layer2_outputs[2021] = layer1_outputs[3677];
    assign layer2_outputs[2022] = (layer1_outputs[4097]) & (layer1_outputs[1614]);
    assign layer2_outputs[2023] = (layer1_outputs[2039]) ^ (layer1_outputs[4161]);
    assign layer2_outputs[2024] = (layer1_outputs[4907]) & (layer1_outputs[595]);
    assign layer2_outputs[2025] = ~(layer1_outputs[2631]);
    assign layer2_outputs[2026] = ~((layer1_outputs[3919]) | (layer1_outputs[4324]));
    assign layer2_outputs[2027] = (layer1_outputs[562]) | (layer1_outputs[88]);
    assign layer2_outputs[2028] = ~(layer1_outputs[3661]);
    assign layer2_outputs[2029] = (layer1_outputs[1473]) | (layer1_outputs[2525]);
    assign layer2_outputs[2030] = ~(layer1_outputs[2527]) | (layer1_outputs[2824]);
    assign layer2_outputs[2031] = (layer1_outputs[4299]) & ~(layer1_outputs[4145]);
    assign layer2_outputs[2032] = (layer1_outputs[2842]) & (layer1_outputs[3072]);
    assign layer2_outputs[2033] = layer1_outputs[3032];
    assign layer2_outputs[2034] = ~(layer1_outputs[16]);
    assign layer2_outputs[2035] = (layer1_outputs[4483]) | (layer1_outputs[3819]);
    assign layer2_outputs[2036] = layer1_outputs[229];
    assign layer2_outputs[2037] = 1'b0;
    assign layer2_outputs[2038] = ~((layer1_outputs[2552]) | (layer1_outputs[3047]));
    assign layer2_outputs[2039] = ~(layer1_outputs[981]) | (layer1_outputs[2393]);
    assign layer2_outputs[2040] = ~(layer1_outputs[1301]);
    assign layer2_outputs[2041] = ~(layer1_outputs[4305]) | (layer1_outputs[3538]);
    assign layer2_outputs[2042] = (layer1_outputs[3554]) & ~(layer1_outputs[1480]);
    assign layer2_outputs[2043] = layer1_outputs[4978];
    assign layer2_outputs[2044] = ~(layer1_outputs[3694]);
    assign layer2_outputs[2045] = ~((layer1_outputs[2876]) & (layer1_outputs[2621]));
    assign layer2_outputs[2046] = (layer1_outputs[4675]) & (layer1_outputs[1962]);
    assign layer2_outputs[2047] = ~(layer1_outputs[3244]) | (layer1_outputs[3806]);
    assign layer2_outputs[2048] = ~(layer1_outputs[2850]);
    assign layer2_outputs[2049] = layer1_outputs[341];
    assign layer2_outputs[2050] = ~(layer1_outputs[3576]);
    assign layer2_outputs[2051] = (layer1_outputs[1575]) & (layer1_outputs[590]);
    assign layer2_outputs[2052] = (layer1_outputs[173]) | (layer1_outputs[2752]);
    assign layer2_outputs[2053] = layer1_outputs[461];
    assign layer2_outputs[2054] = ~((layer1_outputs[1959]) | (layer1_outputs[4513]));
    assign layer2_outputs[2055] = ~((layer1_outputs[4754]) | (layer1_outputs[4237]));
    assign layer2_outputs[2056] = ~(layer1_outputs[4508]);
    assign layer2_outputs[2057] = (layer1_outputs[3299]) & ~(layer1_outputs[216]);
    assign layer2_outputs[2058] = ~(layer1_outputs[3977]) | (layer1_outputs[3482]);
    assign layer2_outputs[2059] = (layer1_outputs[3862]) & ~(layer1_outputs[3204]);
    assign layer2_outputs[2060] = (layer1_outputs[4271]) & ~(layer1_outputs[2136]);
    assign layer2_outputs[2061] = 1'b1;
    assign layer2_outputs[2062] = ~(layer1_outputs[3725]) | (layer1_outputs[2859]);
    assign layer2_outputs[2063] = layer1_outputs[4912];
    assign layer2_outputs[2064] = layer1_outputs[4201];
    assign layer2_outputs[2065] = (layer1_outputs[3500]) & (layer1_outputs[2912]);
    assign layer2_outputs[2066] = (layer1_outputs[3002]) & ~(layer1_outputs[4605]);
    assign layer2_outputs[2067] = ~(layer1_outputs[3996]);
    assign layer2_outputs[2068] = ~(layer1_outputs[4101]);
    assign layer2_outputs[2069] = 1'b0;
    assign layer2_outputs[2070] = layer1_outputs[1523];
    assign layer2_outputs[2071] = ~(layer1_outputs[847]);
    assign layer2_outputs[2072] = 1'b0;
    assign layer2_outputs[2073] = ~(layer1_outputs[47]) | (layer1_outputs[2211]);
    assign layer2_outputs[2074] = layer1_outputs[2536];
    assign layer2_outputs[2075] = ~((layer1_outputs[1717]) | (layer1_outputs[338]));
    assign layer2_outputs[2076] = layer1_outputs[4048];
    assign layer2_outputs[2077] = ~(layer1_outputs[2472]) | (layer1_outputs[2386]);
    assign layer2_outputs[2078] = ~((layer1_outputs[2317]) & (layer1_outputs[543]));
    assign layer2_outputs[2079] = layer1_outputs[2344];
    assign layer2_outputs[2080] = ~(layer1_outputs[2602]);
    assign layer2_outputs[2081] = layer1_outputs[3993];
    assign layer2_outputs[2082] = ~(layer1_outputs[1403]) | (layer1_outputs[431]);
    assign layer2_outputs[2083] = 1'b0;
    assign layer2_outputs[2084] = ~(layer1_outputs[3936]) | (layer1_outputs[988]);
    assign layer2_outputs[2085] = (layer1_outputs[2261]) & ~(layer1_outputs[2643]);
    assign layer2_outputs[2086] = layer1_outputs[5035];
    assign layer2_outputs[2087] = ~(layer1_outputs[198]);
    assign layer2_outputs[2088] = ~(layer1_outputs[4456]);
    assign layer2_outputs[2089] = (layer1_outputs[891]) & (layer1_outputs[2020]);
    assign layer2_outputs[2090] = (layer1_outputs[4956]) & ~(layer1_outputs[4955]);
    assign layer2_outputs[2091] = (layer1_outputs[845]) & (layer1_outputs[4851]);
    assign layer2_outputs[2092] = (layer1_outputs[862]) | (layer1_outputs[880]);
    assign layer2_outputs[2093] = layer1_outputs[81];
    assign layer2_outputs[2094] = ~(layer1_outputs[4197]) | (layer1_outputs[3215]);
    assign layer2_outputs[2095] = ~((layer1_outputs[3346]) & (layer1_outputs[3992]));
    assign layer2_outputs[2096] = ~(layer1_outputs[4353]);
    assign layer2_outputs[2097] = 1'b1;
    assign layer2_outputs[2098] = (layer1_outputs[4813]) ^ (layer1_outputs[2486]);
    assign layer2_outputs[2099] = ~(layer1_outputs[5092]) | (layer1_outputs[5021]);
    assign layer2_outputs[2100] = (layer1_outputs[1463]) & ~(layer1_outputs[2201]);
    assign layer2_outputs[2101] = (layer1_outputs[327]) & (layer1_outputs[4312]);
    assign layer2_outputs[2102] = layer1_outputs[3912];
    assign layer2_outputs[2103] = (layer1_outputs[2684]) & ~(layer1_outputs[1009]);
    assign layer2_outputs[2104] = (layer1_outputs[352]) & ~(layer1_outputs[342]);
    assign layer2_outputs[2105] = layer1_outputs[1705];
    assign layer2_outputs[2106] = (layer1_outputs[2904]) & ~(layer1_outputs[2176]);
    assign layer2_outputs[2107] = ~(layer1_outputs[784]);
    assign layer2_outputs[2108] = (layer1_outputs[783]) & ~(layer1_outputs[4249]);
    assign layer2_outputs[2109] = (layer1_outputs[724]) ^ (layer1_outputs[347]);
    assign layer2_outputs[2110] = ~((layer1_outputs[2808]) | (layer1_outputs[3487]));
    assign layer2_outputs[2111] = ~((layer1_outputs[1018]) | (layer1_outputs[4536]));
    assign layer2_outputs[2112] = (layer1_outputs[438]) & ~(layer1_outputs[3057]);
    assign layer2_outputs[2113] = (layer1_outputs[4204]) ^ (layer1_outputs[2285]);
    assign layer2_outputs[2114] = ~(layer1_outputs[2256]);
    assign layer2_outputs[2115] = ~(layer1_outputs[2492]);
    assign layer2_outputs[2116] = ~(layer1_outputs[262]) | (layer1_outputs[2896]);
    assign layer2_outputs[2117] = ~((layer1_outputs[898]) & (layer1_outputs[2455]));
    assign layer2_outputs[2118] = 1'b1;
    assign layer2_outputs[2119] = (layer1_outputs[3200]) & (layer1_outputs[1627]);
    assign layer2_outputs[2120] = (layer1_outputs[674]) | (layer1_outputs[4223]);
    assign layer2_outputs[2121] = layer1_outputs[3755];
    assign layer2_outputs[2122] = layer1_outputs[3631];
    assign layer2_outputs[2123] = layer1_outputs[2914];
    assign layer2_outputs[2124] = (layer1_outputs[3041]) & ~(layer1_outputs[2207]);
    assign layer2_outputs[2125] = layer1_outputs[2424];
    assign layer2_outputs[2126] = (layer1_outputs[189]) | (layer1_outputs[3294]);
    assign layer2_outputs[2127] = (layer1_outputs[1840]) & ~(layer1_outputs[983]);
    assign layer2_outputs[2128] = ~((layer1_outputs[4727]) & (layer1_outputs[4816]));
    assign layer2_outputs[2129] = layer1_outputs[2731];
    assign layer2_outputs[2130] = ~(layer1_outputs[512]);
    assign layer2_outputs[2131] = ~(layer1_outputs[2711]) | (layer1_outputs[3125]);
    assign layer2_outputs[2132] = ~(layer1_outputs[2557]) | (layer1_outputs[3220]);
    assign layer2_outputs[2133] = (layer1_outputs[2070]) & (layer1_outputs[2552]);
    assign layer2_outputs[2134] = (layer1_outputs[574]) & ~(layer1_outputs[1438]);
    assign layer2_outputs[2135] = ~((layer1_outputs[508]) ^ (layer1_outputs[400]));
    assign layer2_outputs[2136] = 1'b1;
    assign layer2_outputs[2137] = (layer1_outputs[1487]) & ~(layer1_outputs[418]);
    assign layer2_outputs[2138] = ~(layer1_outputs[2190]) | (layer1_outputs[2279]);
    assign layer2_outputs[2139] = (layer1_outputs[3011]) & ~(layer1_outputs[810]);
    assign layer2_outputs[2140] = (layer1_outputs[4406]) & ~(layer1_outputs[3911]);
    assign layer2_outputs[2141] = (layer1_outputs[1219]) | (layer1_outputs[2282]);
    assign layer2_outputs[2142] = (layer1_outputs[2463]) | (layer1_outputs[371]);
    assign layer2_outputs[2143] = 1'b1;
    assign layer2_outputs[2144] = ~((layer1_outputs[456]) | (layer1_outputs[453]));
    assign layer2_outputs[2145] = ~(layer1_outputs[893]) | (layer1_outputs[3400]);
    assign layer2_outputs[2146] = layer1_outputs[348];
    assign layer2_outputs[2147] = ~(layer1_outputs[3619]);
    assign layer2_outputs[2148] = ~(layer1_outputs[344]) | (layer1_outputs[773]);
    assign layer2_outputs[2149] = (layer1_outputs[3050]) | (layer1_outputs[3257]);
    assign layer2_outputs[2150] = ~(layer1_outputs[1451]) | (layer1_outputs[4848]);
    assign layer2_outputs[2151] = ~(layer1_outputs[4217]) | (layer1_outputs[2027]);
    assign layer2_outputs[2152] = (layer1_outputs[2181]) & (layer1_outputs[4425]);
    assign layer2_outputs[2153] = (layer1_outputs[5016]) & ~(layer1_outputs[3453]);
    assign layer2_outputs[2154] = layer1_outputs[5004];
    assign layer2_outputs[2155] = ~((layer1_outputs[3753]) | (layer1_outputs[1688]));
    assign layer2_outputs[2156] = (layer1_outputs[4030]) & (layer1_outputs[3966]);
    assign layer2_outputs[2157] = layer1_outputs[999];
    assign layer2_outputs[2158] = (layer1_outputs[1427]) & ~(layer1_outputs[1067]);
    assign layer2_outputs[2159] = (layer1_outputs[2638]) | (layer1_outputs[2773]);
    assign layer2_outputs[2160] = ~((layer1_outputs[1282]) & (layer1_outputs[3708]));
    assign layer2_outputs[2161] = 1'b0;
    assign layer2_outputs[2162] = layer1_outputs[3547];
    assign layer2_outputs[2163] = layer1_outputs[4671];
    assign layer2_outputs[2164] = (layer1_outputs[3603]) | (layer1_outputs[3178]);
    assign layer2_outputs[2165] = 1'b1;
    assign layer2_outputs[2166] = layer1_outputs[3077];
    assign layer2_outputs[2167] = (layer1_outputs[4673]) & (layer1_outputs[2067]);
    assign layer2_outputs[2168] = (layer1_outputs[3192]) & ~(layer1_outputs[4372]);
    assign layer2_outputs[2169] = layer1_outputs[2650];
    assign layer2_outputs[2170] = layer1_outputs[2881];
    assign layer2_outputs[2171] = layer1_outputs[5055];
    assign layer2_outputs[2172] = (layer1_outputs[4577]) & ~(layer1_outputs[4895]);
    assign layer2_outputs[2173] = ~(layer1_outputs[1241]);
    assign layer2_outputs[2174] = (layer1_outputs[1119]) & ~(layer1_outputs[3888]);
    assign layer2_outputs[2175] = (layer1_outputs[2133]) & ~(layer1_outputs[1186]);
    assign layer2_outputs[2176] = ~((layer1_outputs[5046]) & (layer1_outputs[2046]));
    assign layer2_outputs[2177] = ~(layer1_outputs[3239]) | (layer1_outputs[3000]);
    assign layer2_outputs[2178] = (layer1_outputs[1360]) & (layer1_outputs[2349]);
    assign layer2_outputs[2179] = layer1_outputs[2464];
    assign layer2_outputs[2180] = (layer1_outputs[3869]) & (layer1_outputs[4132]);
    assign layer2_outputs[2181] = (layer1_outputs[1173]) & ~(layer1_outputs[1466]);
    assign layer2_outputs[2182] = ~(layer1_outputs[3032]);
    assign layer2_outputs[2183] = ~(layer1_outputs[667]);
    assign layer2_outputs[2184] = ~((layer1_outputs[1380]) | (layer1_outputs[3948]));
    assign layer2_outputs[2185] = layer1_outputs[3641];
    assign layer2_outputs[2186] = (layer1_outputs[257]) & ~(layer1_outputs[3480]);
    assign layer2_outputs[2187] = (layer1_outputs[2485]) & (layer1_outputs[655]);
    assign layer2_outputs[2188] = (layer1_outputs[1993]) & ~(layer1_outputs[589]);
    assign layer2_outputs[2189] = (layer1_outputs[1877]) & ~(layer1_outputs[619]);
    assign layer2_outputs[2190] = ~(layer1_outputs[4790]);
    assign layer2_outputs[2191] = (layer1_outputs[1729]) & ~(layer1_outputs[2056]);
    assign layer2_outputs[2192] = ~((layer1_outputs[3488]) | (layer1_outputs[4609]));
    assign layer2_outputs[2193] = 1'b0;
    assign layer2_outputs[2194] = ~(layer1_outputs[4663]) | (layer1_outputs[1766]);
    assign layer2_outputs[2195] = ~(layer1_outputs[1081]) | (layer1_outputs[870]);
    assign layer2_outputs[2196] = 1'b1;
    assign layer2_outputs[2197] = 1'b1;
    assign layer2_outputs[2198] = ~((layer1_outputs[2961]) & (layer1_outputs[4558]));
    assign layer2_outputs[2199] = ~((layer1_outputs[1530]) & (layer1_outputs[4672]));
    assign layer2_outputs[2200] = 1'b0;
    assign layer2_outputs[2201] = ~(layer1_outputs[4434]);
    assign layer2_outputs[2202] = (layer1_outputs[1056]) & ~(layer1_outputs[1278]);
    assign layer2_outputs[2203] = ~(layer1_outputs[1630]) | (layer1_outputs[2405]);
    assign layer2_outputs[2204] = ~(layer1_outputs[1504]);
    assign layer2_outputs[2205] = (layer1_outputs[1908]) & (layer1_outputs[1762]);
    assign layer2_outputs[2206] = layer1_outputs[4329];
    assign layer2_outputs[2207] = 1'b0;
    assign layer2_outputs[2208] = ~(layer1_outputs[458]);
    assign layer2_outputs[2209] = (layer1_outputs[2350]) & (layer1_outputs[2708]);
    assign layer2_outputs[2210] = (layer1_outputs[4341]) | (layer1_outputs[1849]);
    assign layer2_outputs[2211] = 1'b1;
    assign layer2_outputs[2212] = ~((layer1_outputs[4983]) | (layer1_outputs[3849]));
    assign layer2_outputs[2213] = (layer1_outputs[719]) | (layer1_outputs[1681]);
    assign layer2_outputs[2214] = layer1_outputs[2608];
    assign layer2_outputs[2215] = (layer1_outputs[3218]) & ~(layer1_outputs[2756]);
    assign layer2_outputs[2216] = 1'b0;
    assign layer2_outputs[2217] = 1'b1;
    assign layer2_outputs[2218] = ~(layer1_outputs[2097]);
    assign layer2_outputs[2219] = ~(layer1_outputs[3205]);
    assign layer2_outputs[2220] = ~(layer1_outputs[4037]) | (layer1_outputs[3030]);
    assign layer2_outputs[2221] = ~((layer1_outputs[1453]) | (layer1_outputs[955]));
    assign layer2_outputs[2222] = (layer1_outputs[3017]) & ~(layer1_outputs[3937]);
    assign layer2_outputs[2223] = ~(layer1_outputs[2175]);
    assign layer2_outputs[2224] = ~(layer1_outputs[1636]);
    assign layer2_outputs[2225] = (layer1_outputs[2720]) & (layer1_outputs[686]);
    assign layer2_outputs[2226] = ~(layer1_outputs[5024]) | (layer1_outputs[4635]);
    assign layer2_outputs[2227] = ~(layer1_outputs[4553]);
    assign layer2_outputs[2228] = (layer1_outputs[5096]) & ~(layer1_outputs[876]);
    assign layer2_outputs[2229] = ~(layer1_outputs[2072]) | (layer1_outputs[5061]);
    assign layer2_outputs[2230] = (layer1_outputs[720]) & ~(layer1_outputs[182]);
    assign layer2_outputs[2231] = 1'b0;
    assign layer2_outputs[2232] = ~((layer1_outputs[1290]) & (layer1_outputs[3093]));
    assign layer2_outputs[2233] = layer1_outputs[89];
    assign layer2_outputs[2234] = layer1_outputs[3720];
    assign layer2_outputs[2235] = ~((layer1_outputs[3644]) & (layer1_outputs[1942]));
    assign layer2_outputs[2236] = layer1_outputs[3522];
    assign layer2_outputs[2237] = ~((layer1_outputs[133]) & (layer1_outputs[1150]));
    assign layer2_outputs[2238] = layer1_outputs[4227];
    assign layer2_outputs[2239] = ~(layer1_outputs[3625]);
    assign layer2_outputs[2240] = 1'b1;
    assign layer2_outputs[2241] = ~(layer1_outputs[1792]);
    assign layer2_outputs[2242] = (layer1_outputs[148]) & ~(layer1_outputs[3780]);
    assign layer2_outputs[2243] = (layer1_outputs[4584]) | (layer1_outputs[2275]);
    assign layer2_outputs[2244] = (layer1_outputs[3957]) & ~(layer1_outputs[3090]);
    assign layer2_outputs[2245] = layer1_outputs[753];
    assign layer2_outputs[2246] = ~((layer1_outputs[2745]) & (layer1_outputs[1058]));
    assign layer2_outputs[2247] = ~(layer1_outputs[3286]);
    assign layer2_outputs[2248] = (layer1_outputs[228]) & ~(layer1_outputs[4484]);
    assign layer2_outputs[2249] = 1'b0;
    assign layer2_outputs[2250] = 1'b0;
    assign layer2_outputs[2251] = ~(layer1_outputs[3308]);
    assign layer2_outputs[2252] = ~(layer1_outputs[4918]);
    assign layer2_outputs[2253] = ~((layer1_outputs[1410]) & (layer1_outputs[5022]));
    assign layer2_outputs[2254] = ~(layer1_outputs[4713]) | (layer1_outputs[4548]);
    assign layer2_outputs[2255] = 1'b0;
    assign layer2_outputs[2256] = layer1_outputs[1073];
    assign layer2_outputs[2257] = ~(layer1_outputs[199]);
    assign layer2_outputs[2258] = ~(layer1_outputs[3347]);
    assign layer2_outputs[2259] = ~(layer1_outputs[4987]) | (layer1_outputs[2231]);
    assign layer2_outputs[2260] = ~((layer1_outputs[616]) & (layer1_outputs[1132]));
    assign layer2_outputs[2261] = ~(layer1_outputs[1500]);
    assign layer2_outputs[2262] = ~((layer1_outputs[2243]) & (layer1_outputs[2348]));
    assign layer2_outputs[2263] = ~((layer1_outputs[2350]) | (layer1_outputs[4990]));
    assign layer2_outputs[2264] = ~(layer1_outputs[2224]) | (layer1_outputs[4807]);
    assign layer2_outputs[2265] = (layer1_outputs[4061]) & (layer1_outputs[4776]);
    assign layer2_outputs[2266] = layer1_outputs[2416];
    assign layer2_outputs[2267] = (layer1_outputs[1013]) & (layer1_outputs[2206]);
    assign layer2_outputs[2268] = layer1_outputs[1814];
    assign layer2_outputs[2269] = (layer1_outputs[4159]) & ~(layer1_outputs[1168]);
    assign layer2_outputs[2270] = ~(layer1_outputs[408]) | (layer1_outputs[4689]);
    assign layer2_outputs[2271] = (layer1_outputs[4971]) & ~(layer1_outputs[1971]);
    assign layer2_outputs[2272] = 1'b1;
    assign layer2_outputs[2273] = ~(layer1_outputs[4054]);
    assign layer2_outputs[2274] = 1'b0;
    assign layer2_outputs[2275] = ~((layer1_outputs[2494]) & (layer1_outputs[2917]));
    assign layer2_outputs[2276] = (layer1_outputs[3938]) & ~(layer1_outputs[3555]);
    assign layer2_outputs[2277] = ~(layer1_outputs[2853]);
    assign layer2_outputs[2278] = layer1_outputs[1181];
    assign layer2_outputs[2279] = ~(layer1_outputs[3423]) | (layer1_outputs[4020]);
    assign layer2_outputs[2280] = ~((layer1_outputs[1588]) | (layer1_outputs[4629]));
    assign layer2_outputs[2281] = layer1_outputs[1309];
    assign layer2_outputs[2282] = ~((layer1_outputs[316]) ^ (layer1_outputs[2317]));
    assign layer2_outputs[2283] = ~((layer1_outputs[4121]) | (layer1_outputs[297]));
    assign layer2_outputs[2284] = ~(layer1_outputs[1618]) | (layer1_outputs[1510]);
    assign layer2_outputs[2285] = layer1_outputs[2112];
    assign layer2_outputs[2286] = ~(layer1_outputs[2247]) | (layer1_outputs[3781]);
    assign layer2_outputs[2287] = ~((layer1_outputs[557]) | (layer1_outputs[1249]));
    assign layer2_outputs[2288] = (layer1_outputs[3079]) & ~(layer1_outputs[2742]);
    assign layer2_outputs[2289] = layer1_outputs[4265];
    assign layer2_outputs[2290] = ~(layer1_outputs[2747]);
    assign layer2_outputs[2291] = 1'b1;
    assign layer2_outputs[2292] = (layer1_outputs[2631]) & (layer1_outputs[4797]);
    assign layer2_outputs[2293] = ~(layer1_outputs[1874]) | (layer1_outputs[503]);
    assign layer2_outputs[2294] = layer1_outputs[1916];
    assign layer2_outputs[2295] = layer1_outputs[2416];
    assign layer2_outputs[2296] = layer1_outputs[3920];
    assign layer2_outputs[2297] = (layer1_outputs[4459]) & ~(layer1_outputs[3061]);
    assign layer2_outputs[2298] = layer1_outputs[3719];
    assign layer2_outputs[2299] = layer1_outputs[2675];
    assign layer2_outputs[2300] = ~((layer1_outputs[439]) & (layer1_outputs[5041]));
    assign layer2_outputs[2301] = (layer1_outputs[4288]) & ~(layer1_outputs[4471]);
    assign layer2_outputs[2302] = layer1_outputs[2407];
    assign layer2_outputs[2303] = ~(layer1_outputs[3818]) | (layer1_outputs[1029]);
    assign layer2_outputs[2304] = 1'b1;
    assign layer2_outputs[2305] = ~(layer1_outputs[3126]);
    assign layer2_outputs[2306] = (layer1_outputs[3116]) & (layer1_outputs[4788]);
    assign layer2_outputs[2307] = ~(layer1_outputs[4418]);
    assign layer2_outputs[2308] = ~(layer1_outputs[851]) | (layer1_outputs[2210]);
    assign layer2_outputs[2309] = ~(layer1_outputs[114]) | (layer1_outputs[1679]);
    assign layer2_outputs[2310] = ~(layer1_outputs[2806]);
    assign layer2_outputs[2311] = (layer1_outputs[1235]) | (layer1_outputs[378]);
    assign layer2_outputs[2312] = (layer1_outputs[3479]) & ~(layer1_outputs[1755]);
    assign layer2_outputs[2313] = layer1_outputs[4265];
    assign layer2_outputs[2314] = layer1_outputs[4685];
    assign layer2_outputs[2315] = ~((layer1_outputs[4198]) ^ (layer1_outputs[4631]));
    assign layer2_outputs[2316] = (layer1_outputs[3899]) | (layer1_outputs[4321]);
    assign layer2_outputs[2317] = layer1_outputs[2223];
    assign layer2_outputs[2318] = (layer1_outputs[4332]) & ~(layer1_outputs[1554]);
    assign layer2_outputs[2319] = layer1_outputs[1268];
    assign layer2_outputs[2320] = layer1_outputs[1838];
    assign layer2_outputs[2321] = layer1_outputs[2963];
    assign layer2_outputs[2322] = layer1_outputs[1713];
    assign layer2_outputs[2323] = ~(layer1_outputs[3942]) | (layer1_outputs[2503]);
    assign layer2_outputs[2324] = ~(layer1_outputs[3456]) | (layer1_outputs[2014]);
    assign layer2_outputs[2325] = ~(layer1_outputs[1687]);
    assign layer2_outputs[2326] = ~(layer1_outputs[2533]);
    assign layer2_outputs[2327] = (layer1_outputs[1376]) & (layer1_outputs[896]);
    assign layer2_outputs[2328] = layer1_outputs[3273];
    assign layer2_outputs[2329] = ~(layer1_outputs[2160]) | (layer1_outputs[2143]);
    assign layer2_outputs[2330] = (layer1_outputs[4859]) & ~(layer1_outputs[3134]);
    assign layer2_outputs[2331] = 1'b1;
    assign layer2_outputs[2332] = 1'b0;
    assign layer2_outputs[2333] = ~(layer1_outputs[1711]) | (layer1_outputs[4135]);
    assign layer2_outputs[2334] = ~(layer1_outputs[1191]);
    assign layer2_outputs[2335] = (layer1_outputs[3880]) ^ (layer1_outputs[2000]);
    assign layer2_outputs[2336] = ~(layer1_outputs[4793]);
    assign layer2_outputs[2337] = ~(layer1_outputs[153]) | (layer1_outputs[1947]);
    assign layer2_outputs[2338] = ~((layer1_outputs[641]) | (layer1_outputs[466]));
    assign layer2_outputs[2339] = ~((layer1_outputs[5012]) | (layer1_outputs[3536]));
    assign layer2_outputs[2340] = ~(layer1_outputs[1275]);
    assign layer2_outputs[2341] = ~((layer1_outputs[859]) | (layer1_outputs[277]));
    assign layer2_outputs[2342] = ~(layer1_outputs[4001]) | (layer1_outputs[1014]);
    assign layer2_outputs[2343] = (layer1_outputs[4047]) & (layer1_outputs[5083]);
    assign layer2_outputs[2344] = ~(layer1_outputs[2712]) | (layer1_outputs[5084]);
    assign layer2_outputs[2345] = 1'b1;
    assign layer2_outputs[2346] = 1'b0;
    assign layer2_outputs[2347] = (layer1_outputs[2746]) & ~(layer1_outputs[149]);
    assign layer2_outputs[2348] = (layer1_outputs[2983]) & (layer1_outputs[1541]);
    assign layer2_outputs[2349] = layer1_outputs[4527];
    assign layer2_outputs[2350] = ~((layer1_outputs[1807]) | (layer1_outputs[2754]));
    assign layer2_outputs[2351] = ~(layer1_outputs[2486]);
    assign layer2_outputs[2352] = ~(layer1_outputs[1074]) | (layer1_outputs[3786]);
    assign layer2_outputs[2353] = (layer1_outputs[2581]) | (layer1_outputs[4225]);
    assign layer2_outputs[2354] = ~(layer1_outputs[3972]);
    assign layer2_outputs[2355] = ~((layer1_outputs[920]) | (layer1_outputs[3507]));
    assign layer2_outputs[2356] = layer1_outputs[313];
    assign layer2_outputs[2357] = layer1_outputs[1622];
    assign layer2_outputs[2358] = (layer1_outputs[1627]) | (layer1_outputs[1505]);
    assign layer2_outputs[2359] = (layer1_outputs[452]) & ~(layer1_outputs[2335]);
    assign layer2_outputs[2360] = layer1_outputs[2656];
    assign layer2_outputs[2361] = layer1_outputs[2074];
    assign layer2_outputs[2362] = (layer1_outputs[4132]) | (layer1_outputs[17]);
    assign layer2_outputs[2363] = 1'b0;
    assign layer2_outputs[2364] = ~(layer1_outputs[3334]);
    assign layer2_outputs[2365] = layer1_outputs[3700];
    assign layer2_outputs[2366] = (layer1_outputs[3352]) & ~(layer1_outputs[3908]);
    assign layer2_outputs[2367] = ~((layer1_outputs[259]) | (layer1_outputs[1635]));
    assign layer2_outputs[2368] = layer1_outputs[943];
    assign layer2_outputs[2369] = layer1_outputs[4223];
    assign layer2_outputs[2370] = (layer1_outputs[424]) & ~(layer1_outputs[2672]);
    assign layer2_outputs[2371] = ~(layer1_outputs[2661]);
    assign layer2_outputs[2372] = (layer1_outputs[3486]) & ~(layer1_outputs[1472]);
    assign layer2_outputs[2373] = (layer1_outputs[1465]) & (layer1_outputs[4710]);
    assign layer2_outputs[2374] = ~((layer1_outputs[3880]) | (layer1_outputs[3627]));
    assign layer2_outputs[2375] = (layer1_outputs[2170]) & ~(layer1_outputs[4394]);
    assign layer2_outputs[2376] = layer1_outputs[1367];
    assign layer2_outputs[2377] = layer1_outputs[4422];
    assign layer2_outputs[2378] = ~(layer1_outputs[823]);
    assign layer2_outputs[2379] = (layer1_outputs[544]) | (layer1_outputs[1616]);
    assign layer2_outputs[2380] = layer1_outputs[4863];
    assign layer2_outputs[2381] = ~(layer1_outputs[2970]);
    assign layer2_outputs[2382] = ~(layer1_outputs[724]) | (layer1_outputs[856]);
    assign layer2_outputs[2383] = layer1_outputs[130];
    assign layer2_outputs[2384] = ~(layer1_outputs[989]) | (layer1_outputs[2450]);
    assign layer2_outputs[2385] = ~(layer1_outputs[1068]);
    assign layer2_outputs[2386] = ~((layer1_outputs[4880]) & (layer1_outputs[2865]));
    assign layer2_outputs[2387] = ~(layer1_outputs[483]) | (layer1_outputs[312]);
    assign layer2_outputs[2388] = (layer1_outputs[245]) & (layer1_outputs[1322]);
    assign layer2_outputs[2389] = ~((layer1_outputs[3283]) & (layer1_outputs[167]));
    assign layer2_outputs[2390] = (layer1_outputs[1785]) & ~(layer1_outputs[2262]);
    assign layer2_outputs[2391] = (layer1_outputs[1841]) | (layer1_outputs[4619]);
    assign layer2_outputs[2392] = 1'b0;
    assign layer2_outputs[2393] = 1'b1;
    assign layer2_outputs[2394] = layer1_outputs[4735];
    assign layer2_outputs[2395] = ~((layer1_outputs[2801]) ^ (layer1_outputs[3389]));
    assign layer2_outputs[2396] = (layer1_outputs[2852]) | (layer1_outputs[2717]);
    assign layer2_outputs[2397] = 1'b0;
    assign layer2_outputs[2398] = ~(layer1_outputs[5075]) | (layer1_outputs[17]);
    assign layer2_outputs[2399] = 1'b1;
    assign layer2_outputs[2400] = layer1_outputs[4361];
    assign layer2_outputs[2401] = ~(layer1_outputs[2354]) | (layer1_outputs[4294]);
    assign layer2_outputs[2402] = 1'b0;
    assign layer2_outputs[2403] = layer1_outputs[2961];
    assign layer2_outputs[2404] = layer1_outputs[3227];
    assign layer2_outputs[2405] = ~(layer1_outputs[1026]) | (layer1_outputs[3851]);
    assign layer2_outputs[2406] = ~((layer1_outputs[2803]) & (layer1_outputs[4118]));
    assign layer2_outputs[2407] = 1'b1;
    assign layer2_outputs[2408] = ~(layer1_outputs[2928]) | (layer1_outputs[1021]);
    assign layer2_outputs[2409] = layer1_outputs[3600];
    assign layer2_outputs[2410] = layer1_outputs[4717];
    assign layer2_outputs[2411] = ~(layer1_outputs[2894]);
    assign layer2_outputs[2412] = layer1_outputs[3076];
    assign layer2_outputs[2413] = ~(layer1_outputs[2825]) | (layer1_outputs[1141]);
    assign layer2_outputs[2414] = ~(layer1_outputs[2088]);
    assign layer2_outputs[2415] = (layer1_outputs[4122]) & ~(layer1_outputs[578]);
    assign layer2_outputs[2416] = ~((layer1_outputs[2334]) & (layer1_outputs[1189]));
    assign layer2_outputs[2417] = ~(layer1_outputs[1468]) | (layer1_outputs[2634]);
    assign layer2_outputs[2418] = ~(layer1_outputs[1917]);
    assign layer2_outputs[2419] = ~(layer1_outputs[3370]);
    assign layer2_outputs[2420] = ~((layer1_outputs[247]) | (layer1_outputs[546]));
    assign layer2_outputs[2421] = layer1_outputs[1608];
    assign layer2_outputs[2422] = ~(layer1_outputs[2429]) | (layer1_outputs[2022]);
    assign layer2_outputs[2423] = layer1_outputs[1715];
    assign layer2_outputs[2424] = (layer1_outputs[3997]) | (layer1_outputs[4385]);
    assign layer2_outputs[2425] = ~(layer1_outputs[1303]);
    assign layer2_outputs[2426] = ~(layer1_outputs[1993]) | (layer1_outputs[740]);
    assign layer2_outputs[2427] = ~(layer1_outputs[4033]);
    assign layer2_outputs[2428] = layer1_outputs[2540];
    assign layer2_outputs[2429] = ~(layer1_outputs[3830]) | (layer1_outputs[2234]);
    assign layer2_outputs[2430] = 1'b0;
    assign layer2_outputs[2431] = (layer1_outputs[2800]) & (layer1_outputs[4503]);
    assign layer2_outputs[2432] = ~((layer1_outputs[2596]) & (layer1_outputs[90]));
    assign layer2_outputs[2433] = (layer1_outputs[4623]) & (layer1_outputs[4729]);
    assign layer2_outputs[2434] = ~(layer1_outputs[4626]);
    assign layer2_outputs[2435] = layer1_outputs[346];
    assign layer2_outputs[2436] = (layer1_outputs[1331]) & ~(layer1_outputs[1518]);
    assign layer2_outputs[2437] = ~(layer1_outputs[2295]);
    assign layer2_outputs[2438] = (layer1_outputs[1224]) & (layer1_outputs[4031]);
    assign layer2_outputs[2439] = ~(layer1_outputs[4074]);
    assign layer2_outputs[2440] = ~((layer1_outputs[2216]) | (layer1_outputs[207]));
    assign layer2_outputs[2441] = ~(layer1_outputs[1858]);
    assign layer2_outputs[2442] = 1'b1;
    assign layer2_outputs[2443] = ~((layer1_outputs[3683]) & (layer1_outputs[1756]));
    assign layer2_outputs[2444] = ~(layer1_outputs[1662]) | (layer1_outputs[4720]);
    assign layer2_outputs[2445] = (layer1_outputs[291]) & ~(layer1_outputs[1667]);
    assign layer2_outputs[2446] = (layer1_outputs[2677]) | (layer1_outputs[3305]);
    assign layer2_outputs[2447] = layer1_outputs[5006];
    assign layer2_outputs[2448] = 1'b1;
    assign layer2_outputs[2449] = (layer1_outputs[4782]) & (layer1_outputs[4225]);
    assign layer2_outputs[2450] = ~(layer1_outputs[3704]) | (layer1_outputs[537]);
    assign layer2_outputs[2451] = ~(layer1_outputs[4532]) | (layer1_outputs[4217]);
    assign layer2_outputs[2452] = (layer1_outputs[4910]) & (layer1_outputs[1314]);
    assign layer2_outputs[2453] = (layer1_outputs[1083]) & (layer1_outputs[4997]);
    assign layer2_outputs[2454] = ~(layer1_outputs[2647]) | (layer1_outputs[156]);
    assign layer2_outputs[2455] = ~((layer1_outputs[5030]) & (layer1_outputs[2361]));
    assign layer2_outputs[2456] = ~(layer1_outputs[2548]) | (layer1_outputs[2238]);
    assign layer2_outputs[2457] = ~(layer1_outputs[1001]);
    assign layer2_outputs[2458] = ~(layer1_outputs[3801]) | (layer1_outputs[1610]);
    assign layer2_outputs[2459] = (layer1_outputs[2803]) & ~(layer1_outputs[4605]);
    assign layer2_outputs[2460] = ~(layer1_outputs[4674]) | (layer1_outputs[4428]);
    assign layer2_outputs[2461] = layer1_outputs[2011];
    assign layer2_outputs[2462] = layer1_outputs[926];
    assign layer2_outputs[2463] = (layer1_outputs[2624]) & ~(layer1_outputs[5008]);
    assign layer2_outputs[2464] = ~(layer1_outputs[2369]);
    assign layer2_outputs[2465] = ~(layer1_outputs[3217]) | (layer1_outputs[3401]);
    assign layer2_outputs[2466] = layer1_outputs[1233];
    assign layer2_outputs[2467] = ~((layer1_outputs[3108]) & (layer1_outputs[2291]));
    assign layer2_outputs[2468] = 1'b1;
    assign layer2_outputs[2469] = layer1_outputs[810];
    assign layer2_outputs[2470] = (layer1_outputs[222]) & ~(layer1_outputs[1911]);
    assign layer2_outputs[2471] = layer1_outputs[54];
    assign layer2_outputs[2472] = (layer1_outputs[96]) | (layer1_outputs[3265]);
    assign layer2_outputs[2473] = ~((layer1_outputs[4289]) & (layer1_outputs[1151]));
    assign layer2_outputs[2474] = 1'b1;
    assign layer2_outputs[2475] = layer1_outputs[2495];
    assign layer2_outputs[2476] = layer1_outputs[4834];
    assign layer2_outputs[2477] = ~((layer1_outputs[3425]) | (layer1_outputs[1398]));
    assign layer2_outputs[2478] = 1'b1;
    assign layer2_outputs[2479] = ~(layer1_outputs[4603]) | (layer1_outputs[3272]);
    assign layer2_outputs[2480] = layer1_outputs[2637];
    assign layer2_outputs[2481] = layer1_outputs[4231];
    assign layer2_outputs[2482] = 1'b0;
    assign layer2_outputs[2483] = (layer1_outputs[4927]) & ~(layer1_outputs[70]);
    assign layer2_outputs[2484] = ~(layer1_outputs[3848]);
    assign layer2_outputs[2485] = ~(layer1_outputs[4373]);
    assign layer2_outputs[2486] = (layer1_outputs[4604]) & ~(layer1_outputs[2043]);
    assign layer2_outputs[2487] = ~((layer1_outputs[169]) | (layer1_outputs[2671]));
    assign layer2_outputs[2488] = (layer1_outputs[2951]) & (layer1_outputs[437]);
    assign layer2_outputs[2489] = layer1_outputs[30];
    assign layer2_outputs[2490] = ~((layer1_outputs[1101]) | (layer1_outputs[185]));
    assign layer2_outputs[2491] = ~(layer1_outputs[3083]) | (layer1_outputs[4519]);
    assign layer2_outputs[2492] = (layer1_outputs[169]) | (layer1_outputs[1712]);
    assign layer2_outputs[2493] = (layer1_outputs[1085]) & ~(layer1_outputs[282]);
    assign layer2_outputs[2494] = ~(layer1_outputs[1831]);
    assign layer2_outputs[2495] = ~(layer1_outputs[1133]);
    assign layer2_outputs[2496] = ~((layer1_outputs[2811]) & (layer1_outputs[3697]));
    assign layer2_outputs[2497] = ~((layer1_outputs[548]) | (layer1_outputs[3251]));
    assign layer2_outputs[2498] = ~(layer1_outputs[1378]) | (layer1_outputs[4255]);
    assign layer2_outputs[2499] = (layer1_outputs[1344]) & ~(layer1_outputs[2560]);
    assign layer2_outputs[2500] = ~((layer1_outputs[2646]) ^ (layer1_outputs[3689]));
    assign layer2_outputs[2501] = ~((layer1_outputs[2413]) ^ (layer1_outputs[1090]));
    assign layer2_outputs[2502] = 1'b0;
    assign layer2_outputs[2503] = (layer1_outputs[2597]) & ~(layer1_outputs[3086]);
    assign layer2_outputs[2504] = ~((layer1_outputs[1024]) | (layer1_outputs[3468]));
    assign layer2_outputs[2505] = ~(layer1_outputs[3913]) | (layer1_outputs[529]);
    assign layer2_outputs[2506] = (layer1_outputs[5018]) & ~(layer1_outputs[783]);
    assign layer2_outputs[2507] = 1'b1;
    assign layer2_outputs[2508] = layer1_outputs[3742];
    assign layer2_outputs[2509] = (layer1_outputs[2871]) & ~(layer1_outputs[365]);
    assign layer2_outputs[2510] = ~((layer1_outputs[1077]) | (layer1_outputs[3571]));
    assign layer2_outputs[2511] = (layer1_outputs[469]) & ~(layer1_outputs[236]);
    assign layer2_outputs[2512] = ~(layer1_outputs[4391]);
    assign layer2_outputs[2513] = layer1_outputs[214];
    assign layer2_outputs[2514] = (layer1_outputs[3364]) | (layer1_outputs[3693]);
    assign layer2_outputs[2515] = 1'b0;
    assign layer2_outputs[2516] = ~(layer1_outputs[268]);
    assign layer2_outputs[2517] = (layer1_outputs[1824]) & ~(layer1_outputs[478]);
    assign layer2_outputs[2518] = ~(layer1_outputs[4872]) | (layer1_outputs[372]);
    assign layer2_outputs[2519] = layer1_outputs[3129];
    assign layer2_outputs[2520] = ~((layer1_outputs[734]) & (layer1_outputs[3422]));
    assign layer2_outputs[2521] = ~(layer1_outputs[5076]) | (layer1_outputs[3184]);
    assign layer2_outputs[2522] = layer1_outputs[3955];
    assign layer2_outputs[2523] = 1'b0;
    assign layer2_outputs[2524] = 1'b0;
    assign layer2_outputs[2525] = ~(layer1_outputs[239]) | (layer1_outputs[1293]);
    assign layer2_outputs[2526] = ~(layer1_outputs[2377]) | (layer1_outputs[2641]);
    assign layer2_outputs[2527] = ~(layer1_outputs[4271]) | (layer1_outputs[2499]);
    assign layer2_outputs[2528] = ~((layer1_outputs[1335]) & (layer1_outputs[897]));
    assign layer2_outputs[2529] = ~(layer1_outputs[227]);
    assign layer2_outputs[2530] = ~((layer1_outputs[3695]) | (layer1_outputs[1686]));
    assign layer2_outputs[2531] = ~(layer1_outputs[3287]);
    assign layer2_outputs[2532] = layer1_outputs[280];
    assign layer2_outputs[2533] = ~(layer1_outputs[3612]);
    assign layer2_outputs[2534] = ~((layer1_outputs[4659]) | (layer1_outputs[1157]));
    assign layer2_outputs[2535] = ~(layer1_outputs[3330]) | (layer1_outputs[45]);
    assign layer2_outputs[2536] = ~(layer1_outputs[2364]);
    assign layer2_outputs[2537] = (layer1_outputs[3792]) | (layer1_outputs[1429]);
    assign layer2_outputs[2538] = ~(layer1_outputs[3804]) | (layer1_outputs[2781]);
    assign layer2_outputs[2539] = (layer1_outputs[3914]) | (layer1_outputs[4757]);
    assign layer2_outputs[2540] = (layer1_outputs[4338]) & ~(layer1_outputs[4706]);
    assign layer2_outputs[2541] = layer1_outputs[3459];
    assign layer2_outputs[2542] = (layer1_outputs[1345]) | (layer1_outputs[3898]);
    assign layer2_outputs[2543] = 1'b0;
    assign layer2_outputs[2544] = (layer1_outputs[1879]) ^ (layer1_outputs[613]);
    assign layer2_outputs[2545] = ~(layer1_outputs[3320]) | (layer1_outputs[1359]);
    assign layer2_outputs[2546] = (layer1_outputs[3049]) & (layer1_outputs[213]);
    assign layer2_outputs[2547] = (layer1_outputs[4985]) ^ (layer1_outputs[4005]);
    assign layer2_outputs[2548] = ~(layer1_outputs[2938]) | (layer1_outputs[2748]);
    assign layer2_outputs[2549] = ~(layer1_outputs[1670]);
    assign layer2_outputs[2550] = (layer1_outputs[4554]) & (layer1_outputs[3924]);
    assign layer2_outputs[2551] = (layer1_outputs[1512]) & ~(layer1_outputs[3668]);
    assign layer2_outputs[2552] = (layer1_outputs[917]) & (layer1_outputs[4190]);
    assign layer2_outputs[2553] = 1'b1;
    assign layer2_outputs[2554] = ~(layer1_outputs[402]);
    assign layer2_outputs[2555] = ~((layer1_outputs[515]) & (layer1_outputs[4446]));
    assign layer2_outputs[2556] = (layer1_outputs[3427]) & (layer1_outputs[3849]);
    assign layer2_outputs[2557] = ~(layer1_outputs[1399]) | (layer1_outputs[4967]);
    assign layer2_outputs[2558] = layer1_outputs[4671];
    assign layer2_outputs[2559] = layer1_outputs[3288];
    assign layer2_outputs[2560] = ~((layer1_outputs[511]) ^ (layer1_outputs[1811]));
    assign layer2_outputs[2561] = 1'b1;
    assign layer2_outputs[2562] = (layer1_outputs[2706]) & ~(layer1_outputs[4293]);
    assign layer2_outputs[2563] = (layer1_outputs[2752]) ^ (layer1_outputs[2483]);
    assign layer2_outputs[2564] = layer1_outputs[5034];
    assign layer2_outputs[2565] = ~((layer1_outputs[4887]) ^ (layer1_outputs[403]));
    assign layer2_outputs[2566] = (layer1_outputs[4471]) ^ (layer1_outputs[4757]);
    assign layer2_outputs[2567] = 1'b1;
    assign layer2_outputs[2568] = (layer1_outputs[1084]) & (layer1_outputs[72]);
    assign layer2_outputs[2569] = 1'b1;
    assign layer2_outputs[2570] = ~((layer1_outputs[544]) | (layer1_outputs[2899]));
    assign layer2_outputs[2571] = layer1_outputs[4559];
    assign layer2_outputs[2572] = ~(layer1_outputs[4854]) | (layer1_outputs[4818]);
    assign layer2_outputs[2573] = (layer1_outputs[982]) | (layer1_outputs[965]);
    assign layer2_outputs[2574] = ~((layer1_outputs[170]) | (layer1_outputs[3220]));
    assign layer2_outputs[2575] = ~((layer1_outputs[4273]) & (layer1_outputs[2206]));
    assign layer2_outputs[2576] = (layer1_outputs[3797]) & (layer1_outputs[2403]);
    assign layer2_outputs[2577] = ~((layer1_outputs[965]) & (layer1_outputs[2132]));
    assign layer2_outputs[2578] = ~(layer1_outputs[2057]);
    assign layer2_outputs[2579] = ~((layer1_outputs[4281]) | (layer1_outputs[903]));
    assign layer2_outputs[2580] = (layer1_outputs[3611]) & ~(layer1_outputs[3407]);
    assign layer2_outputs[2581] = ~(layer1_outputs[29]) | (layer1_outputs[313]);
    assign layer2_outputs[2582] = ~((layer1_outputs[2529]) & (layer1_outputs[2069]));
    assign layer2_outputs[2583] = (layer1_outputs[2110]) & ~(layer1_outputs[545]);
    assign layer2_outputs[2584] = (layer1_outputs[2373]) & ~(layer1_outputs[3290]);
    assign layer2_outputs[2585] = ~(layer1_outputs[3827]);
    assign layer2_outputs[2586] = (layer1_outputs[3340]) & ~(layer1_outputs[1137]);
    assign layer2_outputs[2587] = 1'b0;
    assign layer2_outputs[2588] = ~(layer1_outputs[558]);
    assign layer2_outputs[2589] = 1'b0;
    assign layer2_outputs[2590] = (layer1_outputs[3834]) | (layer1_outputs[2759]);
    assign layer2_outputs[2591] = (layer1_outputs[963]) & (layer1_outputs[863]);
    assign layer2_outputs[2592] = ~(layer1_outputs[1823]);
    assign layer2_outputs[2593] = ~(layer1_outputs[3182]) | (layer1_outputs[3648]);
    assign layer2_outputs[2594] = 1'b0;
    assign layer2_outputs[2595] = layer1_outputs[5036];
    assign layer2_outputs[2596] = layer1_outputs[2525];
    assign layer2_outputs[2597] = (layer1_outputs[2177]) | (layer1_outputs[2574]);
    assign layer2_outputs[2598] = ~(layer1_outputs[3441]) | (layer1_outputs[4195]);
    assign layer2_outputs[2599] = ~(layer1_outputs[10]) | (layer1_outputs[860]);
    assign layer2_outputs[2600] = ~((layer1_outputs[1806]) & (layer1_outputs[1047]));
    assign layer2_outputs[2601] = ~((layer1_outputs[1079]) | (layer1_outputs[3727]));
    assign layer2_outputs[2602] = (layer1_outputs[3592]) & ~(layer1_outputs[4477]);
    assign layer2_outputs[2603] = (layer1_outputs[869]) & ~(layer1_outputs[2205]);
    assign layer2_outputs[2604] = layer1_outputs[4295];
    assign layer2_outputs[2605] = (layer1_outputs[1009]) & ~(layer1_outputs[2045]);
    assign layer2_outputs[2606] = (layer1_outputs[2922]) & ~(layer1_outputs[1492]);
    assign layer2_outputs[2607] = ~((layer1_outputs[2624]) | (layer1_outputs[2288]));
    assign layer2_outputs[2608] = ~(layer1_outputs[1629]);
    assign layer2_outputs[2609] = (layer1_outputs[3532]) | (layer1_outputs[2055]);
    assign layer2_outputs[2610] = ~(layer1_outputs[4134]) | (layer1_outputs[1520]);
    assign layer2_outputs[2611] = layer1_outputs[1533];
    assign layer2_outputs[2612] = (layer1_outputs[390]) & ~(layer1_outputs[830]);
    assign layer2_outputs[2613] = (layer1_outputs[1558]) & ~(layer1_outputs[3759]);
    assign layer2_outputs[2614] = ~(layer1_outputs[906]) | (layer1_outputs[3267]);
    assign layer2_outputs[2615] = layer1_outputs[2971];
    assign layer2_outputs[2616] = (layer1_outputs[3788]) & ~(layer1_outputs[392]);
    assign layer2_outputs[2617] = ~(layer1_outputs[2188]);
    assign layer2_outputs[2618] = ~((layer1_outputs[5013]) & (layer1_outputs[88]));
    assign layer2_outputs[2619] = ~((layer1_outputs[3266]) & (layer1_outputs[1609]));
    assign layer2_outputs[2620] = layer1_outputs[4688];
    assign layer2_outputs[2621] = (layer1_outputs[3835]) | (layer1_outputs[3989]);
    assign layer2_outputs[2622] = 1'b0;
    assign layer2_outputs[2623] = (layer1_outputs[3133]) & ~(layer1_outputs[1098]);
    assign layer2_outputs[2624] = ~(layer1_outputs[698]);
    assign layer2_outputs[2625] = 1'b0;
    assign layer2_outputs[2626] = 1'b1;
    assign layer2_outputs[2627] = ~(layer1_outputs[1441]);
    assign layer2_outputs[2628] = ~(layer1_outputs[4480]);
    assign layer2_outputs[2629] = ~(layer1_outputs[1999]);
    assign layer2_outputs[2630] = ~((layer1_outputs[4354]) | (layer1_outputs[4529]));
    assign layer2_outputs[2631] = (layer1_outputs[2565]) & ~(layer1_outputs[2642]);
    assign layer2_outputs[2632] = ~(layer1_outputs[975]) | (layer1_outputs[3869]);
    assign layer2_outputs[2633] = layer1_outputs[1465];
    assign layer2_outputs[2634] = ~(layer1_outputs[3307]);
    assign layer2_outputs[2635] = ~((layer1_outputs[3389]) | (layer1_outputs[2544]));
    assign layer2_outputs[2636] = (layer1_outputs[3083]) & (layer1_outputs[1134]);
    assign layer2_outputs[2637] = ~((layer1_outputs[530]) | (layer1_outputs[5028]));
    assign layer2_outputs[2638] = ~((layer1_outputs[2944]) | (layer1_outputs[2885]));
    assign layer2_outputs[2639] = (layer1_outputs[2103]) & ~(layer1_outputs[3506]);
    assign layer2_outputs[2640] = layer1_outputs[2877];
    assign layer2_outputs[2641] = ~((layer1_outputs[1207]) | (layer1_outputs[4668]));
    assign layer2_outputs[2642] = (layer1_outputs[3710]) & ~(layer1_outputs[4016]);
    assign layer2_outputs[2643] = layer1_outputs[3325];
    assign layer2_outputs[2644] = layer1_outputs[876];
    assign layer2_outputs[2645] = (layer1_outputs[1793]) ^ (layer1_outputs[362]);
    assign layer2_outputs[2646] = (layer1_outputs[1446]) & (layer1_outputs[2103]);
    assign layer2_outputs[2647] = layer1_outputs[793];
    assign layer2_outputs[2648] = ~(layer1_outputs[2690]);
    assign layer2_outputs[2649] = layer1_outputs[792];
    assign layer2_outputs[2650] = (layer1_outputs[4311]) | (layer1_outputs[1448]);
    assign layer2_outputs[2651] = ~((layer1_outputs[3471]) | (layer1_outputs[4521]));
    assign layer2_outputs[2652] = layer1_outputs[4091];
    assign layer2_outputs[2653] = (layer1_outputs[4661]) | (layer1_outputs[1608]);
    assign layer2_outputs[2654] = ~(layer1_outputs[2052]) | (layer1_outputs[3512]);
    assign layer2_outputs[2655] = ~(layer1_outputs[4496]);
    assign layer2_outputs[2656] = ~(layer1_outputs[2689]);
    assign layer2_outputs[2657] = (layer1_outputs[672]) & (layer1_outputs[3475]);
    assign layer2_outputs[2658] = (layer1_outputs[2434]) & (layer1_outputs[1872]);
    assign layer2_outputs[2659] = (layer1_outputs[4124]) & ~(layer1_outputs[284]);
    assign layer2_outputs[2660] = ~(layer1_outputs[2414]) | (layer1_outputs[4286]);
    assign layer2_outputs[2661] = (layer1_outputs[2997]) & ~(layer1_outputs[1060]);
    assign layer2_outputs[2662] = layer1_outputs[1961];
    assign layer2_outputs[2663] = (layer1_outputs[1117]) | (layer1_outputs[771]);
    assign layer2_outputs[2664] = ~(layer1_outputs[3222]) | (layer1_outputs[4138]);
    assign layer2_outputs[2665] = (layer1_outputs[3850]) & ~(layer1_outputs[1699]);
    assign layer2_outputs[2666] = 1'b0;
    assign layer2_outputs[2667] = layer1_outputs[2036];
    assign layer2_outputs[2668] = (layer1_outputs[4950]) ^ (layer1_outputs[4734]);
    assign layer2_outputs[2669] = ~(layer1_outputs[3421]);
    assign layer2_outputs[2670] = layer1_outputs[451];
    assign layer2_outputs[2671] = (layer1_outputs[1410]) & ~(layer1_outputs[4751]);
    assign layer2_outputs[2672] = ~(layer1_outputs[1914]);
    assign layer2_outputs[2673] = layer1_outputs[606];
    assign layer2_outputs[2674] = ~((layer1_outputs[3324]) | (layer1_outputs[2901]));
    assign layer2_outputs[2675] = ~(layer1_outputs[605]);
    assign layer2_outputs[2676] = (layer1_outputs[270]) & (layer1_outputs[2302]);
    assign layer2_outputs[2677] = (layer1_outputs[231]) & ~(layer1_outputs[1129]);
    assign layer2_outputs[2678] = layer1_outputs[4515];
    assign layer2_outputs[2679] = ~(layer1_outputs[1302]);
    assign layer2_outputs[2680] = (layer1_outputs[3262]) & (layer1_outputs[4625]);
    assign layer2_outputs[2681] = 1'b0;
    assign layer2_outputs[2682] = (layer1_outputs[3336]) ^ (layer1_outputs[4419]);
    assign layer2_outputs[2683] = ~((layer1_outputs[321]) & (layer1_outputs[406]));
    assign layer2_outputs[2684] = ~(layer1_outputs[4098]);
    assign layer2_outputs[2685] = ~(layer1_outputs[4633]) | (layer1_outputs[4731]);
    assign layer2_outputs[2686] = ~((layer1_outputs[314]) | (layer1_outputs[3726]));
    assign layer2_outputs[2687] = (layer1_outputs[3053]) | (layer1_outputs[1859]);
    assign layer2_outputs[2688] = (layer1_outputs[3575]) | (layer1_outputs[2887]);
    assign layer2_outputs[2689] = layer1_outputs[542];
    assign layer2_outputs[2690] = (layer1_outputs[4573]) & ~(layer1_outputs[2915]);
    assign layer2_outputs[2691] = layer1_outputs[1503];
    assign layer2_outputs[2692] = ~(layer1_outputs[5009]);
    assign layer2_outputs[2693] = ~((layer1_outputs[1931]) & (layer1_outputs[3847]));
    assign layer2_outputs[2694] = ~(layer1_outputs[4522]);
    assign layer2_outputs[2695] = ~(layer1_outputs[3361]);
    assign layer2_outputs[2696] = ~((layer1_outputs[3306]) & (layer1_outputs[3776]));
    assign layer2_outputs[2697] = ~((layer1_outputs[141]) ^ (layer1_outputs[680]));
    assign layer2_outputs[2698] = (layer1_outputs[3185]) & ~(layer1_outputs[2445]);
    assign layer2_outputs[2699] = ~(layer1_outputs[3680]);
    assign layer2_outputs[2700] = ~(layer1_outputs[4799]);
    assign layer2_outputs[2701] = (layer1_outputs[3577]) & (layer1_outputs[3062]);
    assign layer2_outputs[2702] = (layer1_outputs[4117]) & ~(layer1_outputs[4219]);
    assign layer2_outputs[2703] = ~(layer1_outputs[3639]);
    assign layer2_outputs[2704] = ~(layer1_outputs[1108]);
    assign layer2_outputs[2705] = ~(layer1_outputs[2996]);
    assign layer2_outputs[2706] = (layer1_outputs[2094]) | (layer1_outputs[4440]);
    assign layer2_outputs[2707] = 1'b0;
    assign layer2_outputs[2708] = ~(layer1_outputs[790]);
    assign layer2_outputs[2709] = ~(layer1_outputs[54]);
    assign layer2_outputs[2710] = layer1_outputs[3591];
    assign layer2_outputs[2711] = layer1_outputs[2747];
    assign layer2_outputs[2712] = ~(layer1_outputs[303]);
    assign layer2_outputs[2713] = (layer1_outputs[215]) & (layer1_outputs[4889]);
    assign layer2_outputs[2714] = layer1_outputs[3218];
    assign layer2_outputs[2715] = (layer1_outputs[533]) & ~(layer1_outputs[3589]);
    assign layer2_outputs[2716] = (layer1_outputs[4551]) & ~(layer1_outputs[308]);
    assign layer2_outputs[2717] = ~(layer1_outputs[2438]);
    assign layer2_outputs[2718] = (layer1_outputs[3244]) & ~(layer1_outputs[1327]);
    assign layer2_outputs[2719] = (layer1_outputs[2427]) | (layer1_outputs[281]);
    assign layer2_outputs[2720] = layer1_outputs[1453];
    assign layer2_outputs[2721] = ~((layer1_outputs[2502]) | (layer1_outputs[3122]));
    assign layer2_outputs[2722] = ~((layer1_outputs[3520]) | (layer1_outputs[4319]));
    assign layer2_outputs[2723] = 1'b0;
    assign layer2_outputs[2724] = ~(layer1_outputs[569]) | (layer1_outputs[1967]);
    assign layer2_outputs[2725] = ~((layer1_outputs[2355]) & (layer1_outputs[4151]));
    assign layer2_outputs[2726] = ~(layer1_outputs[2371]) | (layer1_outputs[3620]);
    assign layer2_outputs[2727] = (layer1_outputs[4440]) & ~(layer1_outputs[4737]);
    assign layer2_outputs[2728] = ~((layer1_outputs[1633]) | (layer1_outputs[3396]));
    assign layer2_outputs[2729] = layer1_outputs[4268];
    assign layer2_outputs[2730] = (layer1_outputs[2241]) | (layer1_outputs[109]);
    assign layer2_outputs[2731] = ~((layer1_outputs[1862]) & (layer1_outputs[1887]));
    assign layer2_outputs[2732] = ~(layer1_outputs[5047]);
    assign layer2_outputs[2733] = ~((layer1_outputs[1628]) | (layer1_outputs[3822]));
    assign layer2_outputs[2734] = ~(layer1_outputs[1106]);
    assign layer2_outputs[2735] = (layer1_outputs[754]) | (layer1_outputs[4431]);
    assign layer2_outputs[2736] = layer1_outputs[2118];
    assign layer2_outputs[2737] = ~(layer1_outputs[894]) | (layer1_outputs[5098]);
    assign layer2_outputs[2738] = ~(layer1_outputs[1348]);
    assign layer2_outputs[2739] = (layer1_outputs[1143]) ^ (layer1_outputs[2972]);
    assign layer2_outputs[2740] = ~(layer1_outputs[1621]) | (layer1_outputs[4867]);
    assign layer2_outputs[2741] = layer1_outputs[617];
    assign layer2_outputs[2742] = ~((layer1_outputs[930]) & (layer1_outputs[3145]));
    assign layer2_outputs[2743] = ~((layer1_outputs[2193]) & (layer1_outputs[2413]));
    assign layer2_outputs[2744] = 1'b0;
    assign layer2_outputs[2745] = layer1_outputs[2497];
    assign layer2_outputs[2746] = ~((layer1_outputs[2280]) & (layer1_outputs[4676]));
    assign layer2_outputs[2747] = layer1_outputs[308];
    assign layer2_outputs[2748] = ~(layer1_outputs[1419]) | (layer1_outputs[1763]);
    assign layer2_outputs[2749] = ~((layer1_outputs[1629]) & (layer1_outputs[2719]));
    assign layer2_outputs[2750] = (layer1_outputs[3823]) & ~(layer1_outputs[3852]);
    assign layer2_outputs[2751] = (layer1_outputs[3295]) | (layer1_outputs[2135]);
    assign layer2_outputs[2752] = ~((layer1_outputs[3569]) | (layer1_outputs[668]));
    assign layer2_outputs[2753] = 1'b1;
    assign layer2_outputs[2754] = ~(layer1_outputs[2641]);
    assign layer2_outputs[2755] = layer1_outputs[4194];
    assign layer2_outputs[2756] = (layer1_outputs[2277]) & ~(layer1_outputs[1634]);
    assign layer2_outputs[2757] = layer1_outputs[710];
    assign layer2_outputs[2758] = (layer1_outputs[1039]) & (layer1_outputs[2863]);
    assign layer2_outputs[2759] = layer1_outputs[1741];
    assign layer2_outputs[2760] = (layer1_outputs[3796]) ^ (layer1_outputs[3698]);
    assign layer2_outputs[2761] = ~(layer1_outputs[510]);
    assign layer2_outputs[2762] = (layer1_outputs[2305]) & ~(layer1_outputs[1555]);
    assign layer2_outputs[2763] = layer1_outputs[579];
    assign layer2_outputs[2764] = layer1_outputs[3254];
    assign layer2_outputs[2765] = layer1_outputs[3777];
    assign layer2_outputs[2766] = (layer1_outputs[1223]) & (layer1_outputs[2054]);
    assign layer2_outputs[2767] = 1'b0;
    assign layer2_outputs[2768] = 1'b0;
    assign layer2_outputs[2769] = 1'b0;
    assign layer2_outputs[2770] = ~((layer1_outputs[1927]) & (layer1_outputs[2721]));
    assign layer2_outputs[2771] = 1'b1;
    assign layer2_outputs[2772] = (layer1_outputs[3467]) & ~(layer1_outputs[2137]);
    assign layer2_outputs[2773] = (layer1_outputs[3838]) & ~(layer1_outputs[3402]);
    assign layer2_outputs[2774] = layer1_outputs[778];
    assign layer2_outputs[2775] = 1'b1;
    assign layer2_outputs[2776] = ~(layer1_outputs[1667]);
    assign layer2_outputs[2777] = (layer1_outputs[4843]) & (layer1_outputs[3762]);
    assign layer2_outputs[2778] = ~(layer1_outputs[625]);
    assign layer2_outputs[2779] = ~((layer1_outputs[2771]) | (layer1_outputs[2130]));
    assign layer2_outputs[2780] = ~((layer1_outputs[1578]) | (layer1_outputs[1092]));
    assign layer2_outputs[2781] = ~(layer1_outputs[3810]);
    assign layer2_outputs[2782] = layer1_outputs[4664];
    assign layer2_outputs[2783] = (layer1_outputs[60]) | (layer1_outputs[1902]);
    assign layer2_outputs[2784] = (layer1_outputs[4380]) & ~(layer1_outputs[1015]);
    assign layer2_outputs[2785] = (layer1_outputs[952]) & (layer1_outputs[1142]);
    assign layer2_outputs[2786] = ~((layer1_outputs[1650]) & (layer1_outputs[1225]));
    assign layer2_outputs[2787] = (layer1_outputs[5104]) & (layer1_outputs[4505]);
    assign layer2_outputs[2788] = 1'b1;
    assign layer2_outputs[2789] = ~(layer1_outputs[1653]);
    assign layer2_outputs[2790] = (layer1_outputs[2230]) & ~(layer1_outputs[856]);
    assign layer2_outputs[2791] = 1'b0;
    assign layer2_outputs[2792] = 1'b0;
    assign layer2_outputs[2793] = ~((layer1_outputs[3479]) | (layer1_outputs[3293]));
    assign layer2_outputs[2794] = layer1_outputs[2259];
    assign layer2_outputs[2795] = layer1_outputs[3841];
    assign layer2_outputs[2796] = (layer1_outputs[4426]) & ~(layer1_outputs[3823]);
    assign layer2_outputs[2797] = (layer1_outputs[2905]) & ~(layer1_outputs[918]);
    assign layer2_outputs[2798] = 1'b1;
    assign layer2_outputs[2799] = ~((layer1_outputs[463]) | (layer1_outputs[4242]));
    assign layer2_outputs[2800] = 1'b0;
    assign layer2_outputs[2801] = (layer1_outputs[4005]) & (layer1_outputs[4999]);
    assign layer2_outputs[2802] = ~(layer1_outputs[4998]) | (layer1_outputs[1327]);
    assign layer2_outputs[2803] = ~(layer1_outputs[4485]);
    assign layer2_outputs[2804] = (layer1_outputs[4556]) & ~(layer1_outputs[1619]);
    assign layer2_outputs[2805] = 1'b0;
    assign layer2_outputs[2806] = (layer1_outputs[2530]) | (layer1_outputs[3203]);
    assign layer2_outputs[2807] = ~((layer1_outputs[2488]) | (layer1_outputs[4490]));
    assign layer2_outputs[2808] = (layer1_outputs[5115]) & ~(layer1_outputs[4992]);
    assign layer2_outputs[2809] = layer1_outputs[4902];
    assign layer2_outputs[2810] = (layer1_outputs[225]) | (layer1_outputs[5056]);
    assign layer2_outputs[2811] = ~((layer1_outputs[3789]) & (layer1_outputs[3776]));
    assign layer2_outputs[2812] = (layer1_outputs[1781]) & ~(layer1_outputs[928]);
    assign layer2_outputs[2813] = ~((layer1_outputs[5031]) & (layer1_outputs[441]));
    assign layer2_outputs[2814] = 1'b0;
    assign layer2_outputs[2815] = ~((layer1_outputs[4586]) | (layer1_outputs[1889]));
    assign layer2_outputs[2816] = 1'b1;
    assign layer2_outputs[2817] = ~(layer1_outputs[3333]) | (layer1_outputs[3168]);
    assign layer2_outputs[2818] = (layer1_outputs[987]) & ~(layer1_outputs[4943]);
    assign layer2_outputs[2819] = ~(layer1_outputs[3580]) | (layer1_outputs[3932]);
    assign layer2_outputs[2820] = ~((layer1_outputs[2252]) & (layer1_outputs[743]));
    assign layer2_outputs[2821] = (layer1_outputs[716]) & ~(layer1_outputs[86]);
    assign layer2_outputs[2822] = ~(layer1_outputs[4277]);
    assign layer2_outputs[2823] = 1'b0;
    assign layer2_outputs[2824] = ~(layer1_outputs[3605]) | (layer1_outputs[415]);
    assign layer2_outputs[2825] = 1'b1;
    assign layer2_outputs[2826] = layer1_outputs[1831];
    assign layer2_outputs[2827] = (layer1_outputs[3068]) & ~(layer1_outputs[2073]);
    assign layer2_outputs[2828] = ~((layer1_outputs[2858]) | (layer1_outputs[1982]));
    assign layer2_outputs[2829] = ~(layer1_outputs[2456]);
    assign layer2_outputs[2830] = ~((layer1_outputs[5029]) | (layer1_outputs[2855]));
    assign layer2_outputs[2831] = 1'b1;
    assign layer2_outputs[2832] = layer1_outputs[3170];
    assign layer2_outputs[2833] = (layer1_outputs[1199]) | (layer1_outputs[256]);
    assign layer2_outputs[2834] = (layer1_outputs[1516]) & ~(layer1_outputs[1591]);
    assign layer2_outputs[2835] = 1'b0;
    assign layer2_outputs[2836] = layer1_outputs[592];
    assign layer2_outputs[2837] = ~(layer1_outputs[1826]);
    assign layer2_outputs[2838] = 1'b1;
    assign layer2_outputs[2839] = (layer1_outputs[1037]) & ~(layer1_outputs[4746]);
    assign layer2_outputs[2840] = ~(layer1_outputs[2006]);
    assign layer2_outputs[2841] = ~((layer1_outputs[1976]) & (layer1_outputs[874]));
    assign layer2_outputs[2842] = ~(layer1_outputs[3554]) | (layer1_outputs[1912]);
    assign layer2_outputs[2843] = ~(layer1_outputs[2670]) | (layer1_outputs[5014]);
    assign layer2_outputs[2844] = layer1_outputs[494];
    assign layer2_outputs[2845] = 1'b0;
    assign layer2_outputs[2846] = ~(layer1_outputs[3282]);
    assign layer2_outputs[2847] = 1'b1;
    assign layer2_outputs[2848] = layer1_outputs[1113];
    assign layer2_outputs[2849] = layer1_outputs[1915];
    assign layer2_outputs[2850] = layer1_outputs[2775];
    assign layer2_outputs[2851] = (layer1_outputs[391]) | (layer1_outputs[1436]);
    assign layer2_outputs[2852] = 1'b0;
    assign layer2_outputs[2853] = layer1_outputs[3660];
    assign layer2_outputs[2854] = 1'b0;
    assign layer2_outputs[2855] = ~((layer1_outputs[3470]) & (layer1_outputs[4565]));
    assign layer2_outputs[2856] = (layer1_outputs[1775]) & ~(layer1_outputs[2730]);
    assign layer2_outputs[2857] = ~((layer1_outputs[1972]) | (layer1_outputs[2008]));
    assign layer2_outputs[2858] = ~(layer1_outputs[5071]);
    assign layer2_outputs[2859] = layer1_outputs[3247];
    assign layer2_outputs[2860] = layer1_outputs[2779];
    assign layer2_outputs[2861] = layer1_outputs[2864];
    assign layer2_outputs[2862] = 1'b0;
    assign layer2_outputs[2863] = ~(layer1_outputs[574]) | (layer1_outputs[2729]);
    assign layer2_outputs[2864] = ~((layer1_outputs[4815]) | (layer1_outputs[2081]));
    assign layer2_outputs[2865] = 1'b0;
    assign layer2_outputs[2866] = ~((layer1_outputs[3537]) & (layer1_outputs[4636]));
    assign layer2_outputs[2867] = ~(layer1_outputs[2030]);
    assign layer2_outputs[2868] = ~((layer1_outputs[1320]) | (layer1_outputs[3187]));
    assign layer2_outputs[2869] = ~(layer1_outputs[1507]);
    assign layer2_outputs[2870] = layer1_outputs[5025];
    assign layer2_outputs[2871] = (layer1_outputs[546]) & ~(layer1_outputs[4608]);
    assign layer2_outputs[2872] = layer1_outputs[2981];
    assign layer2_outputs[2873] = ~(layer1_outputs[1696]);
    assign layer2_outputs[2874] = ~((layer1_outputs[4847]) & (layer1_outputs[1065]));
    assign layer2_outputs[2875] = ~(layer1_outputs[4110]) | (layer1_outputs[3968]);
    assign layer2_outputs[2876] = layer1_outputs[4163];
    assign layer2_outputs[2877] = 1'b0;
    assign layer2_outputs[2878] = 1'b1;
    assign layer2_outputs[2879] = layer1_outputs[3744];
    assign layer2_outputs[2880] = ~(layer1_outputs[3989]) | (layer1_outputs[913]);
    assign layer2_outputs[2881] = ~((layer1_outputs[2714]) ^ (layer1_outputs[4881]));
    assign layer2_outputs[2882] = (layer1_outputs[1152]) & ~(layer1_outputs[2123]);
    assign layer2_outputs[2883] = (layer1_outputs[224]) | (layer1_outputs[5097]);
    assign layer2_outputs[2884] = ~((layer1_outputs[2078]) | (layer1_outputs[2290]));
    assign layer2_outputs[2885] = 1'b0;
    assign layer2_outputs[2886] = 1'b1;
    assign layer2_outputs[2887] = ~((layer1_outputs[4641]) | (layer1_outputs[4449]));
    assign layer2_outputs[2888] = ~((layer1_outputs[4221]) | (layer1_outputs[2524]));
    assign layer2_outputs[2889] = layer1_outputs[4077];
    assign layer2_outputs[2890] = ~(layer1_outputs[708]);
    assign layer2_outputs[2891] = (layer1_outputs[1689]) | (layer1_outputs[3490]);
    assign layer2_outputs[2892] = 1'b0;
    assign layer2_outputs[2893] = ~((layer1_outputs[271]) | (layer1_outputs[4655]));
    assign layer2_outputs[2894] = ~(layer1_outputs[4186]) | (layer1_outputs[837]);
    assign layer2_outputs[2895] = ~(layer1_outputs[357]);
    assign layer2_outputs[2896] = (layer1_outputs[4162]) & ~(layer1_outputs[2853]);
    assign layer2_outputs[2897] = (layer1_outputs[1045]) | (layer1_outputs[1794]);
    assign layer2_outputs[2898] = (layer1_outputs[1915]) & ~(layer1_outputs[1950]);
    assign layer2_outputs[2899] = layer1_outputs[4640];
    assign layer2_outputs[2900] = (layer1_outputs[1041]) & ~(layer1_outputs[4479]);
    assign layer2_outputs[2901] = ~(layer1_outputs[256]) | (layer1_outputs[2151]);
    assign layer2_outputs[2902] = ~(layer1_outputs[3321]) | (layer1_outputs[5093]);
    assign layer2_outputs[2903] = layer1_outputs[2673];
    assign layer2_outputs[2904] = (layer1_outputs[3433]) | (layer1_outputs[402]);
    assign layer2_outputs[2905] = layer1_outputs[915];
    assign layer2_outputs[2906] = ~(layer1_outputs[4934]) | (layer1_outputs[2870]);
    assign layer2_outputs[2907] = ~(layer1_outputs[3859]);
    assign layer2_outputs[2908] = (layer1_outputs[2882]) & ~(layer1_outputs[3652]);
    assign layer2_outputs[2909] = 1'b1;
    assign layer2_outputs[2910] = (layer1_outputs[4762]) | (layer1_outputs[3553]);
    assign layer2_outputs[2911] = ~((layer1_outputs[971]) & (layer1_outputs[1804]));
    assign layer2_outputs[2912] = ~((layer1_outputs[1950]) ^ (layer1_outputs[1726]));
    assign layer2_outputs[2913] = ~((layer1_outputs[4266]) & (layer1_outputs[2976]));
    assign layer2_outputs[2914] = (layer1_outputs[3197]) & (layer1_outputs[1588]);
    assign layer2_outputs[2915] = ~(layer1_outputs[3041]) | (layer1_outputs[3124]);
    assign layer2_outputs[2916] = ~(layer1_outputs[19]);
    assign layer2_outputs[2917] = ~(layer1_outputs[4306]);
    assign layer2_outputs[2918] = ~(layer1_outputs[1693]) | (layer1_outputs[3964]);
    assign layer2_outputs[2919] = layer1_outputs[155];
    assign layer2_outputs[2920] = 1'b0;
    assign layer2_outputs[2921] = layer1_outputs[1537];
    assign layer2_outputs[2922] = layer1_outputs[4662];
    assign layer2_outputs[2923] = (layer1_outputs[1227]) | (layer1_outputs[3871]);
    assign layer2_outputs[2924] = (layer1_outputs[2770]) & ~(layer1_outputs[4018]);
    assign layer2_outputs[2925] = ~((layer1_outputs[498]) ^ (layer1_outputs[4387]));
    assign layer2_outputs[2926] = ~(layer1_outputs[3733]);
    assign layer2_outputs[2927] = layer1_outputs[4292];
    assign layer2_outputs[2928] = ~((layer1_outputs[1458]) | (layer1_outputs[1071]));
    assign layer2_outputs[2929] = layer1_outputs[4521];
    assign layer2_outputs[2930] = ~(layer1_outputs[740]) | (layer1_outputs[3706]);
    assign layer2_outputs[2931] = (layer1_outputs[230]) | (layer1_outputs[2809]);
    assign layer2_outputs[2932] = layer1_outputs[5054];
    assign layer2_outputs[2933] = 1'b1;
    assign layer2_outputs[2934] = layer1_outputs[4252];
    assign layer2_outputs[2935] = layer1_outputs[3841];
    assign layer2_outputs[2936] = 1'b1;
    assign layer2_outputs[2937] = ~(layer1_outputs[3613]) | (layer1_outputs[1085]);
    assign layer2_outputs[2938] = ~((layer1_outputs[3620]) | (layer1_outputs[3654]));
    assign layer2_outputs[2939] = (layer1_outputs[193]) | (layer1_outputs[409]);
    assign layer2_outputs[2940] = ~((layer1_outputs[2783]) & (layer1_outputs[332]));
    assign layer2_outputs[2941] = ~((layer1_outputs[4688]) | (layer1_outputs[2296]));
    assign layer2_outputs[2942] = ~((layer1_outputs[3379]) & (layer1_outputs[487]));
    assign layer2_outputs[2943] = layer1_outputs[4478];
    assign layer2_outputs[2944] = (layer1_outputs[960]) & (layer1_outputs[2927]);
    assign layer2_outputs[2945] = 1'b1;
    assign layer2_outputs[2946] = ~((layer1_outputs[3998]) | (layer1_outputs[4835]));
    assign layer2_outputs[2947] = (layer1_outputs[162]) & ~(layer1_outputs[1249]);
    assign layer2_outputs[2948] = layer1_outputs[4467];
    assign layer2_outputs[2949] = ~(layer1_outputs[288]);
    assign layer2_outputs[2950] = layer1_outputs[2575];
    assign layer2_outputs[2951] = ~(layer1_outputs[4546]);
    assign layer2_outputs[2952] = ~((layer1_outputs[245]) ^ (layer1_outputs[2050]));
    assign layer2_outputs[2953] = ~(layer1_outputs[3468]);
    assign layer2_outputs[2954] = ~((layer1_outputs[1214]) ^ (layer1_outputs[4643]));
    assign layer2_outputs[2955] = (layer1_outputs[736]) & ~(layer1_outputs[777]);
    assign layer2_outputs[2956] = ~((layer1_outputs[1702]) | (layer1_outputs[2273]));
    assign layer2_outputs[2957] = ~(layer1_outputs[2622]);
    assign layer2_outputs[2958] = layer1_outputs[4315];
    assign layer2_outputs[2959] = (layer1_outputs[2306]) | (layer1_outputs[938]);
    assign layer2_outputs[2960] = ~((layer1_outputs[1029]) | (layer1_outputs[643]));
    assign layer2_outputs[2961] = layer1_outputs[4455];
    assign layer2_outputs[2962] = 1'b1;
    assign layer2_outputs[2963] = ~((layer1_outputs[3376]) | (layer1_outputs[1205]));
    assign layer2_outputs[2964] = layer1_outputs[1224];
    assign layer2_outputs[2965] = 1'b0;
    assign layer2_outputs[2966] = (layer1_outputs[1076]) | (layer1_outputs[4369]);
    assign layer2_outputs[2967] = 1'b0;
    assign layer2_outputs[2968] = ~(layer1_outputs[2797]) | (layer1_outputs[2404]);
    assign layer2_outputs[2969] = layer1_outputs[2617];
    assign layer2_outputs[2970] = (layer1_outputs[1042]) & ~(layer1_outputs[2634]);
    assign layer2_outputs[2971] = ~(layer1_outputs[4363]);
    assign layer2_outputs[2972] = ~((layer1_outputs[1330]) & (layer1_outputs[4020]));
    assign layer2_outputs[2973] = layer1_outputs[501];
    assign layer2_outputs[2974] = 1'b0;
    assign layer2_outputs[2975] = ~(layer1_outputs[4239]) | (layer1_outputs[4544]);
    assign layer2_outputs[2976] = layer1_outputs[821];
    assign layer2_outputs[2977] = ~(layer1_outputs[53]) | (layer1_outputs[2691]);
    assign layer2_outputs[2978] = ~(layer1_outputs[2854]) | (layer1_outputs[4295]);
    assign layer2_outputs[2979] = (layer1_outputs[3622]) & ~(layer1_outputs[3413]);
    assign layer2_outputs[2980] = ~((layer1_outputs[261]) | (layer1_outputs[76]));
    assign layer2_outputs[2981] = layer1_outputs[808];
    assign layer2_outputs[2982] = ~((layer1_outputs[4701]) & (layer1_outputs[367]));
    assign layer2_outputs[2983] = layer1_outputs[554];
    assign layer2_outputs[2984] = layer1_outputs[1664];
    assign layer2_outputs[2985] = (layer1_outputs[517]) & ~(layer1_outputs[4849]);
    assign layer2_outputs[2986] = (layer1_outputs[4942]) & ~(layer1_outputs[1247]);
    assign layer2_outputs[2987] = ~((layer1_outputs[1046]) | (layer1_outputs[1602]));
    assign layer2_outputs[2988] = (layer1_outputs[1724]) & (layer1_outputs[1978]);
    assign layer2_outputs[2989] = 1'b1;
    assign layer2_outputs[2990] = ~(layer1_outputs[2663]) | (layer1_outputs[4300]);
    assign layer2_outputs[2991] = layer1_outputs[747];
    assign layer2_outputs[2992] = ~((layer1_outputs[353]) & (layer1_outputs[3458]));
    assign layer2_outputs[2993] = (layer1_outputs[383]) & ~(layer1_outputs[3916]);
    assign layer2_outputs[2994] = ~(layer1_outputs[563]);
    assign layer2_outputs[2995] = ~(layer1_outputs[1451]);
    assign layer2_outputs[2996] = (layer1_outputs[3832]) & ~(layer1_outputs[3311]);
    assign layer2_outputs[2997] = ~(layer1_outputs[3457]) | (layer1_outputs[82]);
    assign layer2_outputs[2998] = ~(layer1_outputs[3892]) | (layer1_outputs[2636]);
    assign layer2_outputs[2999] = ~(layer1_outputs[3544]);
    assign layer2_outputs[3000] = ~(layer1_outputs[4805]) | (layer1_outputs[352]);
    assign layer2_outputs[3001] = (layer1_outputs[185]) & ~(layer1_outputs[3503]);
    assign layer2_outputs[3002] = ~(layer1_outputs[2143]) | (layer1_outputs[3113]);
    assign layer2_outputs[3003] = layer1_outputs[5108];
    assign layer2_outputs[3004] = ~(layer1_outputs[3653]);
    assign layer2_outputs[3005] = 1'b0;
    assign layer2_outputs[3006] = layer1_outputs[3469];
    assign layer2_outputs[3007] = 1'b0;
    assign layer2_outputs[3008] = ~(layer1_outputs[1638]);
    assign layer2_outputs[3009] = ~((layer1_outputs[4396]) & (layer1_outputs[2338]));
    assign layer2_outputs[3010] = (layer1_outputs[2709]) ^ (layer1_outputs[2768]);
    assign layer2_outputs[3011] = ~((layer1_outputs[3100]) | (layer1_outputs[1]));
    assign layer2_outputs[3012] = ~(layer1_outputs[4896]);
    assign layer2_outputs[3013] = ~((layer1_outputs[1582]) & (layer1_outputs[2083]));
    assign layer2_outputs[3014] = (layer1_outputs[824]) & (layer1_outputs[4806]);
    assign layer2_outputs[3015] = 1'b1;
    assign layer2_outputs[3016] = ~((layer1_outputs[3429]) & (layer1_outputs[211]));
    assign layer2_outputs[3017] = ~(layer1_outputs[5033]) | (layer1_outputs[3995]);
    assign layer2_outputs[3018] = ~((layer1_outputs[2841]) & (layer1_outputs[753]));
    assign layer2_outputs[3019] = (layer1_outputs[3276]) & (layer1_outputs[2511]);
    assign layer2_outputs[3020] = ~(layer1_outputs[4699]);
    assign layer2_outputs[3021] = layer1_outputs[2655];
    assign layer2_outputs[3022] = ~(layer1_outputs[4361]) | (layer1_outputs[3485]);
    assign layer2_outputs[3023] = (layer1_outputs[253]) & ~(layer1_outputs[2045]);
    assign layer2_outputs[3024] = ~((layer1_outputs[433]) | (layer1_outputs[3304]));
    assign layer2_outputs[3025] = (layer1_outputs[4120]) & ~(layer1_outputs[5095]);
    assign layer2_outputs[3026] = (layer1_outputs[4202]) & ~(layer1_outputs[924]);
    assign layer2_outputs[3027] = ~((layer1_outputs[4105]) & (layer1_outputs[3340]));
    assign layer2_outputs[3028] = ~(layer1_outputs[3443]);
    assign layer2_outputs[3029] = (layer1_outputs[3461]) & (layer1_outputs[3158]);
    assign layer2_outputs[3030] = ~(layer1_outputs[2896]);
    assign layer2_outputs[3031] = ~(layer1_outputs[5051]);
    assign layer2_outputs[3032] = ~(layer1_outputs[2592]);
    assign layer2_outputs[3033] = ~((layer1_outputs[4889]) & (layer1_outputs[3348]));
    assign layer2_outputs[3034] = ~(layer1_outputs[2378]);
    assign layer2_outputs[3035] = 1'b0;
    assign layer2_outputs[3036] = (layer1_outputs[5103]) | (layer1_outputs[774]);
    assign layer2_outputs[3037] = 1'b0;
    assign layer2_outputs[3038] = ~(layer1_outputs[1295]);
    assign layer2_outputs[3039] = (layer1_outputs[2366]) & ~(layer1_outputs[568]);
    assign layer2_outputs[3040] = (layer1_outputs[1300]) & ~(layer1_outputs[3359]);
    assign layer2_outputs[3041] = ~(layer1_outputs[2041]) | (layer1_outputs[853]);
    assign layer2_outputs[3042] = (layer1_outputs[831]) & (layer1_outputs[4574]);
    assign layer2_outputs[3043] = ~(layer1_outputs[3464]) | (layer1_outputs[1194]);
    assign layer2_outputs[3044] = ~(layer1_outputs[4855]);
    assign layer2_outputs[3045] = ~((layer1_outputs[1925]) & (layer1_outputs[1943]));
    assign layer2_outputs[3046] = (layer1_outputs[2369]) & ~(layer1_outputs[1176]);
    assign layer2_outputs[3047] = layer1_outputs[648];
    assign layer2_outputs[3048] = ~(layer1_outputs[1773]);
    assign layer2_outputs[3049] = ~(layer1_outputs[645]) | (layer1_outputs[2394]);
    assign layer2_outputs[3050] = (layer1_outputs[3401]) | (layer1_outputs[3304]);
    assign layer2_outputs[3051] = ~(layer1_outputs[3911]);
    assign layer2_outputs[3052] = (layer1_outputs[1149]) & (layer1_outputs[3342]);
    assign layer2_outputs[3053] = layer1_outputs[1115];
    assign layer2_outputs[3054] = layer1_outputs[4627];
    assign layer2_outputs[3055] = ~((layer1_outputs[4492]) & (layer1_outputs[2728]));
    assign layer2_outputs[3056] = (layer1_outputs[4056]) & (layer1_outputs[1905]);
    assign layer2_outputs[3057] = (layer1_outputs[4692]) & ~(layer1_outputs[799]);
    assign layer2_outputs[3058] = ~(layer1_outputs[4852]);
    assign layer2_outputs[3059] = ~(layer1_outputs[1368]) | (layer1_outputs[2445]);
    assign layer2_outputs[3060] = layer1_outputs[1148];
    assign layer2_outputs[3061] = layer1_outputs[2582];
    assign layer2_outputs[3062] = ~(layer1_outputs[5088]) | (layer1_outputs[1966]);
    assign layer2_outputs[3063] = layer1_outputs[3115];
    assign layer2_outputs[3064] = layer1_outputs[1694];
    assign layer2_outputs[3065] = ~(layer1_outputs[3952]) | (layer1_outputs[982]);
    assign layer2_outputs[3066] = 1'b0;
    assign layer2_outputs[3067] = layer1_outputs[1949];
    assign layer2_outputs[3068] = layer1_outputs[4402];
    assign layer2_outputs[3069] = 1'b1;
    assign layer2_outputs[3070] = ~((layer1_outputs[2200]) ^ (layer1_outputs[1820]));
    assign layer2_outputs[3071] = (layer1_outputs[1769]) & ~(layer1_outputs[2686]);
    assign layer2_outputs[3072] = (layer1_outputs[5052]) | (layer1_outputs[3110]);
    assign layer2_outputs[3073] = layer1_outputs[226];
    assign layer2_outputs[3074] = ~((layer1_outputs[3456]) | (layer1_outputs[2625]));
    assign layer2_outputs[3075] = (layer1_outputs[504]) | (layer1_outputs[4450]);
    assign layer2_outputs[3076] = ~(layer1_outputs[4021]);
    assign layer2_outputs[3077] = layer1_outputs[166];
    assign layer2_outputs[3078] = 1'b0;
    assign layer2_outputs[3079] = ~(layer1_outputs[4133]) | (layer1_outputs[837]);
    assign layer2_outputs[3080] = ~(layer1_outputs[777]);
    assign layer2_outputs[3081] = 1'b0;
    assign layer2_outputs[3082] = ~(layer1_outputs[221]);
    assign layer2_outputs[3083] = ~((layer1_outputs[4653]) | (layer1_outputs[1514]));
    assign layer2_outputs[3084] = (layer1_outputs[2837]) & ~(layer1_outputs[4989]);
    assign layer2_outputs[3085] = 1'b0;
    assign layer2_outputs[3086] = ~((layer1_outputs[2149]) & (layer1_outputs[2452]));
    assign layer2_outputs[3087] = 1'b0;
    assign layer2_outputs[3088] = (layer1_outputs[81]) & ~(layer1_outputs[1723]);
    assign layer2_outputs[3089] = ~(layer1_outputs[2563]) | (layer1_outputs[4192]);
    assign layer2_outputs[3090] = (layer1_outputs[2242]) ^ (layer1_outputs[3232]);
    assign layer2_outputs[3091] = ~((layer1_outputs[4952]) & (layer1_outputs[2814]));
    assign layer2_outputs[3092] = (layer1_outputs[3444]) | (layer1_outputs[1057]);
    assign layer2_outputs[3093] = 1'b0;
    assign layer2_outputs[3094] = ~((layer1_outputs[1476]) & (layer1_outputs[2012]));
    assign layer2_outputs[3095] = (layer1_outputs[1818]) & ~(layer1_outputs[1427]);
    assign layer2_outputs[3096] = ~(layer1_outputs[2920]) | (layer1_outputs[95]);
    assign layer2_outputs[3097] = ~((layer1_outputs[4813]) ^ (layer1_outputs[2980]));
    assign layer2_outputs[3098] = (layer1_outputs[1728]) | (layer1_outputs[3186]);
    assign layer2_outputs[3099] = 1'b1;
    assign layer2_outputs[3100] = ~((layer1_outputs[2184]) | (layer1_outputs[1118]));
    assign layer2_outputs[3101] = ~((layer1_outputs[4258]) | (layer1_outputs[1380]));
    assign layer2_outputs[3102] = ~((layer1_outputs[2756]) | (layer1_outputs[3450]));
    assign layer2_outputs[3103] = 1'b1;
    assign layer2_outputs[3104] = layer1_outputs[3596];
    assign layer2_outputs[3105] = 1'b1;
    assign layer2_outputs[3106] = layer1_outputs[2018];
    assign layer2_outputs[3107] = (layer1_outputs[2233]) & ~(layer1_outputs[4828]);
    assign layer2_outputs[3108] = ~(layer1_outputs[765]);
    assign layer2_outputs[3109] = ~(layer1_outputs[835]) | (layer1_outputs[186]);
    assign layer2_outputs[3110] = ~(layer1_outputs[350]);
    assign layer2_outputs[3111] = ~(layer1_outputs[3745]);
    assign layer2_outputs[3112] = layer1_outputs[3565];
    assign layer2_outputs[3113] = (layer1_outputs[4789]) | (layer1_outputs[4058]);
    assign layer2_outputs[3114] = ~(layer1_outputs[2600]);
    assign layer2_outputs[3115] = ~((layer1_outputs[2240]) & (layer1_outputs[3969]));
    assign layer2_outputs[3116] = layer1_outputs[260];
    assign layer2_outputs[3117] = layer1_outputs[307];
    assign layer2_outputs[3118] = (layer1_outputs[5062]) | (layer1_outputs[611]);
    assign layer2_outputs[3119] = ~(layer1_outputs[4786]) | (layer1_outputs[3264]);
    assign layer2_outputs[3120] = ~(layer1_outputs[2588]);
    assign layer2_outputs[3121] = layer1_outputs[3470];
    assign layer2_outputs[3122] = ~((layer1_outputs[1422]) | (layer1_outputs[1390]));
    assign layer2_outputs[3123] = layer1_outputs[13];
    assign layer2_outputs[3124] = (layer1_outputs[2434]) & (layer1_outputs[3409]);
    assign layer2_outputs[3125] = ~(layer1_outputs[1869]);
    assign layer2_outputs[3126] = layer1_outputs[1139];
    assign layer2_outputs[3127] = 1'b0;
    assign layer2_outputs[3128] = ~(layer1_outputs[3883]) | (layer1_outputs[5039]);
    assign layer2_outputs[3129] = ~(layer1_outputs[3419]) | (layer1_outputs[2466]);
    assign layer2_outputs[3130] = ~(layer1_outputs[901]);
    assign layer2_outputs[3131] = ~(layer1_outputs[4937]) | (layer1_outputs[4155]);
    assign layer2_outputs[3132] = layer1_outputs[1233];
    assign layer2_outputs[3133] = 1'b1;
    assign layer2_outputs[3134] = (layer1_outputs[3575]) | (layer1_outputs[50]);
    assign layer2_outputs[3135] = layer1_outputs[761];
    assign layer2_outputs[3136] = ~((layer1_outputs[3728]) & (layer1_outputs[3568]));
    assign layer2_outputs[3137] = layer1_outputs[4634];
    assign layer2_outputs[3138] = layer1_outputs[1784];
    assign layer2_outputs[3139] = ~(layer1_outputs[464]);
    assign layer2_outputs[3140] = (layer1_outputs[2581]) & (layer1_outputs[3839]);
    assign layer2_outputs[3141] = (layer1_outputs[2509]) & ~(layer1_outputs[3630]);
    assign layer2_outputs[3142] = ~(layer1_outputs[4507]);
    assign layer2_outputs[3143] = (layer1_outputs[99]) & ~(layer1_outputs[31]);
    assign layer2_outputs[3144] = ~(layer1_outputs[1719]);
    assign layer2_outputs[3145] = ~((layer1_outputs[4302]) | (layer1_outputs[3276]));
    assign layer2_outputs[3146] = ~((layer1_outputs[204]) & (layer1_outputs[3847]));
    assign layer2_outputs[3147] = ~(layer1_outputs[2338]) | (layer1_outputs[2890]);
    assign layer2_outputs[3148] = ~(layer1_outputs[2558]);
    assign layer2_outputs[3149] = ~(layer1_outputs[355]);
    assign layer2_outputs[3150] = (layer1_outputs[2663]) | (layer1_outputs[3812]);
    assign layer2_outputs[3151] = ~(layer1_outputs[4904]) | (layer1_outputs[2906]);
    assign layer2_outputs[3152] = (layer1_outputs[4758]) | (layer1_outputs[2236]);
    assign layer2_outputs[3153] = 1'b0;
    assign layer2_outputs[3154] = ~(layer1_outputs[125]);
    assign layer2_outputs[3155] = (layer1_outputs[2773]) | (layer1_outputs[3850]);
    assign layer2_outputs[3156] = ~((layer1_outputs[371]) | (layer1_outputs[5049]));
    assign layer2_outputs[3157] = ~(layer1_outputs[786]);
    assign layer2_outputs[3158] = ~(layer1_outputs[1494]) | (layer1_outputs[4779]);
    assign layer2_outputs[3159] = ~(layer1_outputs[5057]);
    assign layer2_outputs[3160] = ~((layer1_outputs[330]) ^ (layer1_outputs[3807]));
    assign layer2_outputs[3161] = (layer1_outputs[3026]) & ~(layer1_outputs[1873]);
    assign layer2_outputs[3162] = layer1_outputs[101];
    assign layer2_outputs[3163] = layer1_outputs[3785];
    assign layer2_outputs[3164] = (layer1_outputs[3888]) & ~(layer1_outputs[2948]);
    assign layer2_outputs[3165] = (layer1_outputs[2846]) & ~(layer1_outputs[2698]);
    assign layer2_outputs[3166] = layer1_outputs[1665];
    assign layer2_outputs[3167] = layer1_outputs[3394];
    assign layer2_outputs[3168] = layer1_outputs[1461];
    assign layer2_outputs[3169] = ~((layer1_outputs[403]) | (layer1_outputs[597]));
    assign layer2_outputs[3170] = 1'b0;
    assign layer2_outputs[3171] = (layer1_outputs[2262]) & ~(layer1_outputs[692]);
    assign layer2_outputs[3172] = ~((layer1_outputs[1028]) ^ (layer1_outputs[43]));
    assign layer2_outputs[3173] = 1'b1;
    assign layer2_outputs[3174] = ~(layer1_outputs[2526]);
    assign layer2_outputs[3175] = (layer1_outputs[666]) ^ (layer1_outputs[2800]);
    assign layer2_outputs[3176] = (layer1_outputs[3973]) & ~(layer1_outputs[2359]);
    assign layer2_outputs[3177] = (layer1_outputs[117]) | (layer1_outputs[509]);
    assign layer2_outputs[3178] = ~((layer1_outputs[3893]) | (layer1_outputs[3271]));
    assign layer2_outputs[3179] = ~(layer1_outputs[1971]);
    assign layer2_outputs[3180] = ~((layer1_outputs[3579]) & (layer1_outputs[2425]));
    assign layer2_outputs[3181] = ~((layer1_outputs[4850]) | (layer1_outputs[294]));
    assign layer2_outputs[3182] = 1'b0;
    assign layer2_outputs[3183] = layer1_outputs[5090];
    assign layer2_outputs[3184] = 1'b1;
    assign layer2_outputs[3185] = (layer1_outputs[2328]) | (layer1_outputs[377]);
    assign layer2_outputs[3186] = layer1_outputs[1565];
    assign layer2_outputs[3187] = (layer1_outputs[1732]) ^ (layer1_outputs[2071]);
    assign layer2_outputs[3188] = (layer1_outputs[1137]) & ~(layer1_outputs[2291]);
    assign layer2_outputs[3189] = (layer1_outputs[1740]) & ~(layer1_outputs[3897]);
    assign layer2_outputs[3190] = ~((layer1_outputs[2484]) & (layer1_outputs[2089]));
    assign layer2_outputs[3191] = ~(layer1_outputs[444]);
    assign layer2_outputs[3192] = layer1_outputs[4951];
    assign layer2_outputs[3193] = (layer1_outputs[4994]) & (layer1_outputs[4106]);
    assign layer2_outputs[3194] = (layer1_outputs[2429]) | (layer1_outputs[966]);
    assign layer2_outputs[3195] = ~((layer1_outputs[2715]) ^ (layer1_outputs[2267]));
    assign layer2_outputs[3196] = ~(layer1_outputs[3067]);
    assign layer2_outputs[3197] = 1'b1;
    assign layer2_outputs[3198] = ~(layer1_outputs[3011]) | (layer1_outputs[921]);
    assign layer2_outputs[3199] = 1'b1;
    assign layer2_outputs[3200] = ~((layer1_outputs[4533]) & (layer1_outputs[2633]));
    assign layer2_outputs[3201] = ~((layer1_outputs[1870]) | (layer1_outputs[4024]));
    assign layer2_outputs[3202] = ~((layer1_outputs[819]) | (layer1_outputs[1053]));
    assign layer2_outputs[3203] = 1'b0;
    assign layer2_outputs[3204] = ~(layer1_outputs[2386]);
    assign layer2_outputs[3205] = ~((layer1_outputs[2036]) & (layer1_outputs[4961]));
    assign layer2_outputs[3206] = layer1_outputs[1805];
    assign layer2_outputs[3207] = (layer1_outputs[305]) & (layer1_outputs[3685]);
    assign layer2_outputs[3208] = (layer1_outputs[372]) & ~(layer1_outputs[2090]);
    assign layer2_outputs[3209] = ~(layer1_outputs[3291]);
    assign layer2_outputs[3210] = ~(layer1_outputs[1263]);
    assign layer2_outputs[3211] = layer1_outputs[4711];
    assign layer2_outputs[3212] = ~(layer1_outputs[298]) | (layer1_outputs[5064]);
    assign layer2_outputs[3213] = layer1_outputs[4169];
    assign layer2_outputs[3214] = (layer1_outputs[1339]) & ~(layer1_outputs[1665]);
    assign layer2_outputs[3215] = layer1_outputs[2670];
    assign layer2_outputs[3216] = ~(layer1_outputs[2515]);
    assign layer2_outputs[3217] = (layer1_outputs[1456]) & ~(layer1_outputs[1477]);
    assign layer2_outputs[3218] = (layer1_outputs[4569]) | (layer1_outputs[3711]);
    assign layer2_outputs[3219] = layer1_outputs[264];
    assign layer2_outputs[3220] = (layer1_outputs[2652]) | (layer1_outputs[1916]);
    assign layer2_outputs[3221] = (layer1_outputs[1506]) & ~(layer1_outputs[2707]);
    assign layer2_outputs[3222] = ~((layer1_outputs[4609]) & (layer1_outputs[1382]));
    assign layer2_outputs[3223] = (layer1_outputs[4487]) & (layer1_outputs[3681]);
    assign layer2_outputs[3224] = ~(layer1_outputs[929]) | (layer1_outputs[4173]);
    assign layer2_outputs[3225] = (layer1_outputs[4421]) ^ (layer1_outputs[1167]);
    assign layer2_outputs[3226] = (layer1_outputs[4723]) & ~(layer1_outputs[615]);
    assign layer2_outputs[3227] = ~(layer1_outputs[1612]) | (layer1_outputs[2863]);
    assign layer2_outputs[3228] = (layer1_outputs[3252]) & ~(layer1_outputs[146]);
    assign layer2_outputs[3229] = (layer1_outputs[3229]) & (layer1_outputs[4629]);
    assign layer2_outputs[3230] = ~(layer1_outputs[3891]);
    assign layer2_outputs[3231] = layer1_outputs[2432];
    assign layer2_outputs[3232] = ~((layer1_outputs[3539]) | (layer1_outputs[2500]));
    assign layer2_outputs[3233] = ~((layer1_outputs[2968]) & (layer1_outputs[4494]));
    assign layer2_outputs[3234] = ~(layer1_outputs[1182]);
    assign layer2_outputs[3235] = 1'b1;
    assign layer2_outputs[3236] = layer1_outputs[524];
    assign layer2_outputs[3237] = layer1_outputs[229];
    assign layer2_outputs[3238] = ~(layer1_outputs[656]);
    assign layer2_outputs[3239] = layer1_outputs[976];
    assign layer2_outputs[3240] = ~(layer1_outputs[3434]) | (layer1_outputs[5080]);
    assign layer2_outputs[3241] = layer1_outputs[1981];
    assign layer2_outputs[3242] = layer1_outputs[609];
    assign layer2_outputs[3243] = 1'b1;
    assign layer2_outputs[3244] = (layer1_outputs[129]) & (layer1_outputs[8]);
    assign layer2_outputs[3245] = (layer1_outputs[3391]) & (layer1_outputs[2454]);
    assign layer2_outputs[3246] = (layer1_outputs[717]) & ~(layer1_outputs[1079]);
    assign layer2_outputs[3247] = ~(layer1_outputs[3250]);
    assign layer2_outputs[3248] = (layer1_outputs[1867]) & ~(layer1_outputs[3655]);
    assign layer2_outputs[3249] = layer1_outputs[4797];
    assign layer2_outputs[3250] = ~((layer1_outputs[605]) & (layer1_outputs[319]));
    assign layer2_outputs[3251] = (layer1_outputs[4579]) ^ (layer1_outputs[4208]);
    assign layer2_outputs[3252] = ~(layer1_outputs[4633]);
    assign layer2_outputs[3253] = ~((layer1_outputs[2953]) | (layer1_outputs[284]));
    assign layer2_outputs[3254] = ~(layer1_outputs[2289]);
    assign layer2_outputs[3255] = (layer1_outputs[1658]) & ~(layer1_outputs[4844]);
    assign layer2_outputs[3256] = ~((layer1_outputs[27]) | (layer1_outputs[4631]));
    assign layer2_outputs[3257] = (layer1_outputs[1373]) ^ (layer1_outputs[1678]);
    assign layer2_outputs[3258] = ~(layer1_outputs[4461]) | (layer1_outputs[2457]);
    assign layer2_outputs[3259] = layer1_outputs[2134];
    assign layer2_outputs[3260] = 1'b1;
    assign layer2_outputs[3261] = ~((layer1_outputs[3826]) & (layer1_outputs[2384]));
    assign layer2_outputs[3262] = ~(layer1_outputs[1363]) | (layer1_outputs[2702]);
    assign layer2_outputs[3263] = (layer1_outputs[3045]) & ~(layer1_outputs[485]);
    assign layer2_outputs[3264] = ~((layer1_outputs[1180]) ^ (layer1_outputs[2164]));
    assign layer2_outputs[3265] = ~(layer1_outputs[4759]);
    assign layer2_outputs[3266] = ~(layer1_outputs[1159]) | (layer1_outputs[488]);
    assign layer2_outputs[3267] = (layer1_outputs[3509]) | (layer1_outputs[1277]);
    assign layer2_outputs[3268] = ~(layer1_outputs[2706]);
    assign layer2_outputs[3269] = ~((layer1_outputs[4809]) & (layer1_outputs[4436]));
    assign layer2_outputs[3270] = (layer1_outputs[4319]) & (layer1_outputs[1389]);
    assign layer2_outputs[3271] = 1'b0;
    assign layer2_outputs[3272] = layer1_outputs[4925];
    assign layer2_outputs[3273] = ~(layer1_outputs[361]) | (layer1_outputs[3514]);
    assign layer2_outputs[3274] = 1'b0;
    assign layer2_outputs[3275] = ~(layer1_outputs[1926]);
    assign layer2_outputs[3276] = (layer1_outputs[2549]) & (layer1_outputs[997]);
    assign layer2_outputs[3277] = 1'b1;
    assign layer2_outputs[3278] = (layer1_outputs[2428]) & ~(layer1_outputs[1168]);
    assign layer2_outputs[3279] = ~((layer1_outputs[3452]) & (layer1_outputs[4045]));
    assign layer2_outputs[3280] = ~(layer1_outputs[4027]);
    assign layer2_outputs[3281] = layer1_outputs[4872];
    assign layer2_outputs[3282] = ~(layer1_outputs[4630]);
    assign layer2_outputs[3283] = (layer1_outputs[2388]) & ~(layer1_outputs[3171]);
    assign layer2_outputs[3284] = ~(layer1_outputs[808]) | (layer1_outputs[495]);
    assign layer2_outputs[3285] = 1'b1;
    assign layer2_outputs[3286] = ~(layer1_outputs[3721]) | (layer1_outputs[962]);
    assign layer2_outputs[3287] = 1'b0;
    assign layer2_outputs[3288] = 1'b1;
    assign layer2_outputs[3289] = (layer1_outputs[2921]) & (layer1_outputs[4445]);
    assign layer2_outputs[3290] = (layer1_outputs[3187]) & ~(layer1_outputs[1790]);
    assign layer2_outputs[3291] = 1'b1;
    assign layer2_outputs[3292] = ~(layer1_outputs[738]);
    assign layer2_outputs[3293] = ~(layer1_outputs[843]) | (layer1_outputs[984]);
    assign layer2_outputs[3294] = ~(layer1_outputs[1337]);
    assign layer2_outputs[3295] = layer1_outputs[5088];
    assign layer2_outputs[3296] = (layer1_outputs[855]) & ~(layer1_outputs[1060]);
    assign layer2_outputs[3297] = ~(layer1_outputs[834]);
    assign layer2_outputs[3298] = ~(layer1_outputs[84]) | (layer1_outputs[4307]);
    assign layer2_outputs[3299] = (layer1_outputs[4395]) | (layer1_outputs[3621]);
    assign layer2_outputs[3300] = (layer1_outputs[2955]) & (layer1_outputs[3448]);
    assign layer2_outputs[3301] = (layer1_outputs[3043]) & (layer1_outputs[3258]);
    assign layer2_outputs[3302] = ~((layer1_outputs[2751]) & (layer1_outputs[2504]));
    assign layer2_outputs[3303] = ~(layer1_outputs[722]);
    assign layer2_outputs[3304] = ~(layer1_outputs[1940]) | (layer1_outputs[2100]);
    assign layer2_outputs[3305] = (layer1_outputs[1268]) & ~(layer1_outputs[121]);
    assign layer2_outputs[3306] = layer1_outputs[3533];
    assign layer2_outputs[3307] = ~(layer1_outputs[923]) | (layer1_outputs[3395]);
    assign layer2_outputs[3308] = 1'b0;
    assign layer2_outputs[3309] = layer1_outputs[434];
    assign layer2_outputs[3310] = ~(layer1_outputs[4557]);
    assign layer2_outputs[3311] = 1'b1;
    assign layer2_outputs[3312] = layer1_outputs[4453];
    assign layer2_outputs[3313] = layer1_outputs[126];
    assign layer2_outputs[3314] = ~(layer1_outputs[3610]) | (layer1_outputs[1219]);
    assign layer2_outputs[3315] = 1'b1;
    assign layer2_outputs[3316] = (layer1_outputs[3491]) | (layer1_outputs[1442]);
    assign layer2_outputs[3317] = ~(layer1_outputs[4326]) | (layer1_outputs[2209]);
    assign layer2_outputs[3318] = ~(layer1_outputs[4940]);
    assign layer2_outputs[3319] = ~(layer1_outputs[4095]) | (layer1_outputs[1550]);
    assign layer2_outputs[3320] = 1'b0;
    assign layer2_outputs[3321] = layer1_outputs[3143];
    assign layer2_outputs[3322] = ~((layer1_outputs[2104]) | (layer1_outputs[2913]));
    assign layer2_outputs[3323] = layer1_outputs[406];
    assign layer2_outputs[3324] = layer1_outputs[1598];
    assign layer2_outputs[3325] = 1'b0;
    assign layer2_outputs[3326] = layer1_outputs[2024];
    assign layer2_outputs[3327] = (layer1_outputs[1032]) & ~(layer1_outputs[2405]);
    assign layer2_outputs[3328] = ~(layer1_outputs[3959]) | (layer1_outputs[2555]);
    assign layer2_outputs[3329] = layer1_outputs[3582];
    assign layer2_outputs[3330] = ~(layer1_outputs[289]) | (layer1_outputs[1668]);
    assign layer2_outputs[3331] = (layer1_outputs[283]) ^ (layer1_outputs[240]);
    assign layer2_outputs[3332] = 1'b1;
    assign layer2_outputs[3333] = ~(layer1_outputs[1686]);
    assign layer2_outputs[3334] = (layer1_outputs[977]) & ~(layer1_outputs[4117]);
    assign layer2_outputs[3335] = layer1_outputs[3164];
    assign layer2_outputs[3336] = ~(layer1_outputs[519]);
    assign layer2_outputs[3337] = (layer1_outputs[2950]) & (layer1_outputs[3635]);
    assign layer2_outputs[3338] = ~(layer1_outputs[5118]) | (layer1_outputs[979]);
    assign layer2_outputs[3339] = layer1_outputs[1564];
    assign layer2_outputs[3340] = (layer1_outputs[2239]) ^ (layer1_outputs[539]);
    assign layer2_outputs[3341] = ~(layer1_outputs[1059]) | (layer1_outputs[3109]);
    assign layer2_outputs[3342] = (layer1_outputs[2813]) & ~(layer1_outputs[3403]);
    assign layer2_outputs[3343] = 1'b0;
    assign layer2_outputs[3344] = (layer1_outputs[1524]) & (layer1_outputs[851]);
    assign layer2_outputs[3345] = layer1_outputs[4260];
    assign layer2_outputs[3346] = (layer1_outputs[745]) & (layer1_outputs[2952]);
    assign layer2_outputs[3347] = (layer1_outputs[1951]) & ~(layer1_outputs[3138]);
    assign layer2_outputs[3348] = 1'b1;
    assign layer2_outputs[3349] = ~((layer1_outputs[1174]) | (layer1_outputs[2615]));
    assign layer2_outputs[3350] = (layer1_outputs[2767]) & (layer1_outputs[2902]);
    assign layer2_outputs[3351] = (layer1_outputs[1999]) ^ (layer1_outputs[1521]);
    assign layer2_outputs[3352] = layer1_outputs[1375];
    assign layer2_outputs[3353] = 1'b0;
    assign layer2_outputs[3354] = 1'b1;
    assign layer2_outputs[3355] = ~((layer1_outputs[3255]) | (layer1_outputs[2314]));
    assign layer2_outputs[3356] = (layer1_outputs[1334]) | (layer1_outputs[1632]);
    assign layer2_outputs[3357] = ~((layer1_outputs[3567]) | (layer1_outputs[1700]));
    assign layer2_outputs[3358] = (layer1_outputs[2267]) & (layer1_outputs[4038]);
    assign layer2_outputs[3359] = ~(layer1_outputs[2812]);
    assign layer2_outputs[3360] = ~((layer1_outputs[1655]) ^ (layer1_outputs[1845]));
    assign layer2_outputs[3361] = layer1_outputs[2916];
    assign layer2_outputs[3362] = (layer1_outputs[664]) & ~(layer1_outputs[2328]);
    assign layer2_outputs[3363] = (layer1_outputs[219]) | (layer1_outputs[3226]);
    assign layer2_outputs[3364] = layer1_outputs[2698];
    assign layer2_outputs[3365] = ~(layer1_outputs[2931]);
    assign layer2_outputs[3366] = ~(layer1_outputs[5051]) | (layer1_outputs[2166]);
    assign layer2_outputs[3367] = 1'b0;
    assign layer2_outputs[3368] = ~((layer1_outputs[2772]) ^ (layer1_outputs[5040]));
    assign layer2_outputs[3369] = ~((layer1_outputs[2936]) & (layer1_outputs[4601]));
    assign layer2_outputs[3370] = ~((layer1_outputs[277]) | (layer1_outputs[633]));
    assign layer2_outputs[3371] = ~((layer1_outputs[1956]) | (layer1_outputs[425]));
    assign layer2_outputs[3372] = (layer1_outputs[489]) & (layer1_outputs[5037]);
    assign layer2_outputs[3373] = layer1_outputs[2493];
    assign layer2_outputs[3374] = (layer1_outputs[4697]) & (layer1_outputs[2015]);
    assign layer2_outputs[3375] = ~((layer1_outputs[2677]) | (layer1_outputs[1592]));
    assign layer2_outputs[3376] = 1'b0;
    assign layer2_outputs[3377] = ~(layer1_outputs[11]);
    assign layer2_outputs[3378] = ~((layer1_outputs[2385]) & (layer1_outputs[64]));
    assign layer2_outputs[3379] = (layer1_outputs[2816]) & (layer1_outputs[4059]);
    assign layer2_outputs[3380] = 1'b1;
    assign layer2_outputs[3381] = ~(layer1_outputs[3348]) | (layer1_outputs[315]);
    assign layer2_outputs[3382] = (layer1_outputs[2298]) & (layer1_outputs[1882]);
    assign layer2_outputs[3383] = ~(layer1_outputs[890]) | (layer1_outputs[3862]);
    assign layer2_outputs[3384] = 1'b1;
    assign layer2_outputs[3385] = ~(layer1_outputs[1488]) | (layer1_outputs[4267]);
    assign layer2_outputs[3386] = layer1_outputs[2716];
    assign layer2_outputs[3387] = layer1_outputs[3248];
    assign layer2_outputs[3388] = (layer1_outputs[2066]) | (layer1_outputs[4324]);
    assign layer2_outputs[3389] = 1'b0;
    assign layer2_outputs[3390] = ~(layer1_outputs[4556]);
    assign layer2_outputs[3391] = (layer1_outputs[3525]) | (layer1_outputs[2935]);
    assign layer2_outputs[3392] = ~(layer1_outputs[1216]);
    assign layer2_outputs[3393] = ~(layer1_outputs[1450]) | (layer1_outputs[1435]);
    assign layer2_outputs[3394] = 1'b0;
    assign layer2_outputs[3395] = ~(layer1_outputs[2996]);
    assign layer2_outputs[3396] = ~(layer1_outputs[986]);
    assign layer2_outputs[3397] = ~(layer1_outputs[3345]);
    assign layer2_outputs[3398] = 1'b0;
    assign layer2_outputs[3399] = 1'b1;
    assign layer2_outputs[3400] = ~(layer1_outputs[4555]);
    assign layer2_outputs[3401] = (layer1_outputs[196]) & ~(layer1_outputs[4703]);
    assign layer2_outputs[3402] = (layer1_outputs[4774]) & (layer1_outputs[903]);
    assign layer2_outputs[3403] = 1'b0;
    assign layer2_outputs[3404] = (layer1_outputs[3590]) ^ (layer1_outputs[1666]);
    assign layer2_outputs[3405] = (layer1_outputs[1892]) & ~(layer1_outputs[4085]);
    assign layer2_outputs[3406] = (layer1_outputs[3741]) & ~(layer1_outputs[3715]);
    assign layer2_outputs[3407] = ~(layer1_outputs[1120]);
    assign layer2_outputs[3408] = (layer1_outputs[2236]) & ~(layer1_outputs[2319]);
    assign layer2_outputs[3409] = (layer1_outputs[3190]) & ~(layer1_outputs[993]);
    assign layer2_outputs[3410] = ~(layer1_outputs[398]) | (layer1_outputs[2914]);
    assign layer2_outputs[3411] = ~(layer1_outputs[3100]);
    assign layer2_outputs[3412] = ~(layer1_outputs[4566]) | (layer1_outputs[444]);
    assign layer2_outputs[3413] = layer1_outputs[3695];
    assign layer2_outputs[3414] = ~(layer1_outputs[3060]);
    assign layer2_outputs[3415] = ~(layer1_outputs[1337]) | (layer1_outputs[4742]);
    assign layer2_outputs[3416] = ~(layer1_outputs[1482]);
    assign layer2_outputs[3417] = ~(layer1_outputs[3199]);
    assign layer2_outputs[3418] = ~((layer1_outputs[3991]) | (layer1_outputs[4990]));
    assign layer2_outputs[3419] = (layer1_outputs[762]) | (layer1_outputs[368]);
    assign layer2_outputs[3420] = (layer1_outputs[1923]) & ~(layer1_outputs[1691]);
    assign layer2_outputs[3421] = ~(layer1_outputs[3821]);
    assign layer2_outputs[3422] = layer1_outputs[1940];
    assign layer2_outputs[3423] = ~(layer1_outputs[1116]) | (layer1_outputs[3669]);
    assign layer2_outputs[3424] = layer1_outputs[4996];
    assign layer2_outputs[3425] = (layer1_outputs[2795]) & ~(layer1_outputs[1326]);
    assign layer2_outputs[3426] = (layer1_outputs[4248]) | (layer1_outputs[1161]);
    assign layer2_outputs[3427] = ~(layer1_outputs[2794]);
    assign layer2_outputs[3428] = ~((layer1_outputs[1449]) | (layer1_outputs[1898]));
    assign layer2_outputs[3429] = ~(layer1_outputs[3501]) | (layer1_outputs[3152]);
    assign layer2_outputs[3430] = ~(layer1_outputs[512]);
    assign layer2_outputs[3431] = ~(layer1_outputs[2732]) | (layer1_outputs[4530]);
    assign layer2_outputs[3432] = (layer1_outputs[661]) & ~(layer1_outputs[1531]);
    assign layer2_outputs[3433] = layer1_outputs[4988];
    assign layer2_outputs[3434] = (layer1_outputs[4599]) & (layer1_outputs[4492]);
    assign layer2_outputs[3435] = ~((layer1_outputs[2334]) & (layer1_outputs[4831]));
    assign layer2_outputs[3436] = 1'b0;
    assign layer2_outputs[3437] = layer1_outputs[1792];
    assign layer2_outputs[3438] = layer1_outputs[4582];
    assign layer2_outputs[3439] = ~(layer1_outputs[4239]);
    assign layer2_outputs[3440] = ~((layer1_outputs[4083]) | (layer1_outputs[1391]));
    assign layer2_outputs[3441] = 1'b1;
    assign layer2_outputs[3442] = (layer1_outputs[2903]) & (layer1_outputs[1408]);
    assign layer2_outputs[3443] = layer1_outputs[3734];
    assign layer2_outputs[3444] = layer1_outputs[3915];
    assign layer2_outputs[3445] = ~((layer1_outputs[833]) & (layer1_outputs[746]));
    assign layer2_outputs[3446] = ~((layer1_outputs[3584]) | (layer1_outputs[295]));
    assign layer2_outputs[3447] = ~(layer1_outputs[4932]) | (layer1_outputs[2182]);
    assign layer2_outputs[3448] = ~(layer1_outputs[597]);
    assign layer2_outputs[3449] = ~(layer1_outputs[4348]);
    assign layer2_outputs[3450] = ~(layer1_outputs[2220]);
    assign layer2_outputs[3451] = ~((layer1_outputs[4788]) | (layer1_outputs[1585]));
    assign layer2_outputs[3452] = (layer1_outputs[802]) & (layer1_outputs[4096]);
    assign layer2_outputs[3453] = ~((layer1_outputs[4301]) & (layer1_outputs[3981]));
    assign layer2_outputs[3454] = layer1_outputs[616];
    assign layer2_outputs[3455] = (layer1_outputs[353]) | (layer1_outputs[821]);
    assign layer2_outputs[3456] = (layer1_outputs[1948]) & (layer1_outputs[4122]);
    assign layer2_outputs[3457] = 1'b0;
    assign layer2_outputs[3458] = 1'b0;
    assign layer2_outputs[3459] = 1'b0;
    assign layer2_outputs[3460] = ~(layer1_outputs[4833]);
    assign layer2_outputs[3461] = layer1_outputs[3957];
    assign layer2_outputs[3462] = layer1_outputs[1995];
    assign layer2_outputs[3463] = (layer1_outputs[1672]) & ~(layer1_outputs[4421]);
    assign layer2_outputs[3464] = (layer1_outputs[266]) & (layer1_outputs[1742]);
    assign layer2_outputs[3465] = ~((layer1_outputs[4091]) & (layer1_outputs[522]));
    assign layer2_outputs[3466] = (layer1_outputs[2332]) & ~(layer1_outputs[1044]);
    assign layer2_outputs[3467] = (layer1_outputs[4455]) ^ (layer1_outputs[1498]);
    assign layer2_outputs[3468] = ~(layer1_outputs[1251]) | (layer1_outputs[130]);
    assign layer2_outputs[3469] = ~((layer1_outputs[3983]) ^ (layer1_outputs[1763]));
    assign layer2_outputs[3470] = 1'b0;
    assign layer2_outputs[3471] = layer1_outputs[3980];
    assign layer2_outputs[3472] = ~(layer1_outputs[3814]) | (layer1_outputs[2867]);
    assign layer2_outputs[3473] = ~(layer1_outputs[2095]) | (layer1_outputs[4171]);
    assign layer2_outputs[3474] = 1'b1;
    assign layer2_outputs[3475] = (layer1_outputs[1479]) & (layer1_outputs[852]);
    assign layer2_outputs[3476] = 1'b0;
    assign layer2_outputs[3477] = layer1_outputs[3099];
    assign layer2_outputs[3478] = layer1_outputs[3538];
    assign layer2_outputs[3479] = ~((layer1_outputs[62]) & (layer1_outputs[3386]));
    assign layer2_outputs[3480] = ~((layer1_outputs[4821]) | (layer1_outputs[4092]));
    assign layer2_outputs[3481] = ~((layer1_outputs[1597]) ^ (layer1_outputs[384]));
    assign layer2_outputs[3482] = ~(layer1_outputs[1567]);
    assign layer2_outputs[3483] = (layer1_outputs[627]) & (layer1_outputs[2298]);
    assign layer2_outputs[3484] = ~(layer1_outputs[3471]);
    assign layer2_outputs[3485] = ~((layer1_outputs[1598]) | (layer1_outputs[481]));
    assign layer2_outputs[3486] = layer1_outputs[4224];
    assign layer2_outputs[3487] = layer1_outputs[4289];
    assign layer2_outputs[3488] = layer1_outputs[1611];
    assign layer2_outputs[3489] = 1'b1;
    assign layer2_outputs[3490] = ~(layer1_outputs[4885]);
    assign layer2_outputs[3491] = ~((layer1_outputs[3633]) ^ (layer1_outputs[2411]));
    assign layer2_outputs[3492] = (layer1_outputs[2544]) & (layer1_outputs[3763]);
    assign layer2_outputs[3493] = ~(layer1_outputs[3208]);
    assign layer2_outputs[3494] = (layer1_outputs[1642]) & (layer1_outputs[4905]);
    assign layer2_outputs[3495] = 1'b0;
    assign layer2_outputs[3496] = ~((layer1_outputs[2474]) & (layer1_outputs[4142]));
    assign layer2_outputs[3497] = 1'b1;
    assign layer2_outputs[3498] = (layer1_outputs[1652]) ^ (layer1_outputs[2306]);
    assign layer2_outputs[3499] = (layer1_outputs[3119]) & (layer1_outputs[4695]);
    assign layer2_outputs[3500] = 1'b0;
    assign layer2_outputs[3501] = ~(layer1_outputs[798]);
    assign layer2_outputs[3502] = 1'b0;
    assign layer2_outputs[3503] = ~((layer1_outputs[1214]) & (layer1_outputs[455]));
    assign layer2_outputs[3504] = layer1_outputs[565];
    assign layer2_outputs[3505] = layer1_outputs[2778];
    assign layer2_outputs[3506] = layer1_outputs[1884];
    assign layer2_outputs[3507] = (layer1_outputs[3201]) & (layer1_outputs[1674]);
    assign layer2_outputs[3508] = ~(layer1_outputs[1600]) | (layer1_outputs[3302]);
    assign layer2_outputs[3509] = ~(layer1_outputs[1764]);
    assign layer2_outputs[3510] = ~(layer1_outputs[703]) | (layer1_outputs[234]);
    assign layer2_outputs[3511] = ~(layer1_outputs[900]);
    assign layer2_outputs[3512] = ~(layer1_outputs[4193]);
    assign layer2_outputs[3513] = 1'b0;
    assign layer2_outputs[3514] = 1'b1;
    assign layer2_outputs[3515] = 1'b0;
    assign layer2_outputs[3516] = (layer1_outputs[888]) & ~(layer1_outputs[2797]);
    assign layer2_outputs[3517] = ~((layer1_outputs[4032]) & (layer1_outputs[3509]));
    assign layer2_outputs[3518] = ~((layer1_outputs[2591]) | (layer1_outputs[3436]));
    assign layer2_outputs[3519] = 1'b1;
    assign layer2_outputs[3520] = ~(layer1_outputs[3091]) | (layer1_outputs[2194]);
    assign layer2_outputs[3521] = ~(layer1_outputs[2278]);
    assign layer2_outputs[3522] = ~(layer1_outputs[111]);
    assign layer2_outputs[3523] = ~(layer1_outputs[414]) | (layer1_outputs[1232]);
    assign layer2_outputs[3524] = (layer1_outputs[3598]) ^ (layer1_outputs[4335]);
    assign layer2_outputs[3525] = layer1_outputs[216];
    assign layer2_outputs[3526] = layer1_outputs[933];
    assign layer2_outputs[3527] = (layer1_outputs[348]) & ~(layer1_outputs[1893]);
    assign layer2_outputs[3528] = 1'b1;
    assign layer2_outputs[3529] = ~((layer1_outputs[2255]) | (layer1_outputs[3523]));
    assign layer2_outputs[3530] = ~(layer1_outputs[3595]);
    assign layer2_outputs[3531] = ~(layer1_outputs[2152]);
    assign layer2_outputs[3532] = ~(layer1_outputs[3566]);
    assign layer2_outputs[3533] = ~(layer1_outputs[2847]);
    assign layer2_outputs[3534] = layer1_outputs[3932];
    assign layer2_outputs[3535] = ~(layer1_outputs[3739]);
    assign layer2_outputs[3536] = ~(layer1_outputs[2449]) | (layer1_outputs[2102]);
    assign layer2_outputs[3537] = 1'b1;
    assign layer2_outputs[3538] = (layer1_outputs[4228]) & ~(layer1_outputs[2235]);
    assign layer2_outputs[3539] = ~((layer1_outputs[1907]) | (layer1_outputs[4661]));
    assign layer2_outputs[3540] = 1'b1;
    assign layer2_outputs[3541] = ~(layer1_outputs[4365]);
    assign layer2_outputs[3542] = layer1_outputs[3607];
    assign layer2_outputs[3543] = ~((layer1_outputs[4346]) & (layer1_outputs[5061]));
    assign layer2_outputs[3544] = ~((layer1_outputs[3210]) | (layer1_outputs[4562]));
    assign layer2_outputs[3545] = (layer1_outputs[3063]) | (layer1_outputs[2120]);
    assign layer2_outputs[3546] = ~(layer1_outputs[3213]);
    assign layer2_outputs[3547] = ~(layer1_outputs[2943]) | (layer1_outputs[4401]);
    assign layer2_outputs[3548] = (layer1_outputs[1890]) & (layer1_outputs[4420]);
    assign layer2_outputs[3549] = ~(layer1_outputs[942]);
    assign layer2_outputs[3550] = (layer1_outputs[1455]) ^ (layer1_outputs[3290]);
    assign layer2_outputs[3551] = ~(layer1_outputs[4422]);
    assign layer2_outputs[3552] = ~((layer1_outputs[2697]) | (layer1_outputs[598]));
    assign layer2_outputs[3553] = 1'b0;
    assign layer2_outputs[3554] = ~(layer1_outputs[3736]) | (layer1_outputs[2358]);
    assign layer2_outputs[3555] = ~(layer1_outputs[4306]) | (layer1_outputs[3949]);
    assign layer2_outputs[3556] = ~((layer1_outputs[4437]) & (layer1_outputs[2125]));
    assign layer2_outputs[3557] = ~((layer1_outputs[5111]) | (layer1_outputs[4689]));
    assign layer2_outputs[3558] = (layer1_outputs[1336]) | (layer1_outputs[2804]);
    assign layer2_outputs[3559] = 1'b1;
    assign layer2_outputs[3560] = layer1_outputs[994];
    assign layer2_outputs[3561] = layer1_outputs[4920];
    assign layer2_outputs[3562] = 1'b0;
    assign layer2_outputs[3563] = ~(layer1_outputs[945]);
    assign layer2_outputs[3564] = ~(layer1_outputs[52]) | (layer1_outputs[1289]);
    assign layer2_outputs[3565] = ~(layer1_outputs[1815]);
    assign layer2_outputs[3566] = (layer1_outputs[5027]) & (layer1_outputs[2621]);
    assign layer2_outputs[3567] = ~((layer1_outputs[405]) | (layer1_outputs[4258]));
    assign layer2_outputs[3568] = (layer1_outputs[128]) & ~(layer1_outputs[2293]);
    assign layer2_outputs[3569] = 1'b0;
    assign layer2_outputs[3570] = ~(layer1_outputs[1174]);
    assign layer2_outputs[3571] = ~((layer1_outputs[5038]) ^ (layer1_outputs[380]));
    assign layer2_outputs[3572] = ~((layer1_outputs[3018]) | (layer1_outputs[4869]));
    assign layer2_outputs[3573] = (layer1_outputs[2282]) & ~(layer1_outputs[261]);
    assign layer2_outputs[3574] = (layer1_outputs[613]) ^ (layer1_outputs[4268]);
    assign layer2_outputs[3575] = ~(layer1_outputs[4112]) | (layer1_outputs[860]);
    assign layer2_outputs[3576] = 1'b1;
    assign layer2_outputs[3577] = 1'b0;
    assign layer2_outputs[3578] = layer1_outputs[567];
    assign layer2_outputs[3579] = ~((layer1_outputs[2257]) & (layer1_outputs[2645]));
    assign layer2_outputs[3580] = (layer1_outputs[2676]) & ~(layer1_outputs[3403]);
    assign layer2_outputs[3581] = (layer1_outputs[178]) & ~(layer1_outputs[3357]);
    assign layer2_outputs[3582] = 1'b0;
    assign layer2_outputs[3583] = (layer1_outputs[3277]) & ~(layer1_outputs[93]);
    assign layer2_outputs[3584] = 1'b0;
    assign layer2_outputs[3585] = (layer1_outputs[3167]) & (layer1_outputs[4297]);
    assign layer2_outputs[3586] = (layer1_outputs[4787]) & ~(layer1_outputs[2320]);
    assign layer2_outputs[3587] = layer1_outputs[3505];
    assign layer2_outputs[3588] = ~(layer1_outputs[1210]);
    assign layer2_outputs[3589] = layer1_outputs[2665];
    assign layer2_outputs[3590] = ~((layer1_outputs[4281]) & (layer1_outputs[3679]));
    assign layer2_outputs[3591] = layer1_outputs[4109];
    assign layer2_outputs[3592] = (layer1_outputs[2651]) & ~(layer1_outputs[3689]);
    assign layer2_outputs[3593] = 1'b1;
    assign layer2_outputs[3594] = ~(layer1_outputs[1160]);
    assign layer2_outputs[3595] = ~((layer1_outputs[3922]) & (layer1_outputs[3928]));
    assign layer2_outputs[3596] = layer1_outputs[1799];
    assign layer2_outputs[3597] = (layer1_outputs[1779]) ^ (layer1_outputs[1273]);
    assign layer2_outputs[3598] = layer1_outputs[2305];
    assign layer2_outputs[3599] = layer1_outputs[2522];
    assign layer2_outputs[3600] = ~((layer1_outputs[4250]) | (layer1_outputs[3516]));
    assign layer2_outputs[3601] = ~(layer1_outputs[1310]);
    assign layer2_outputs[3602] = (layer1_outputs[721]) | (layer1_outputs[5105]);
    assign layer2_outputs[3603] = (layer1_outputs[3592]) | (layer1_outputs[3072]);
    assign layer2_outputs[3604] = ~(layer1_outputs[1056]);
    assign layer2_outputs[3605] = (layer1_outputs[1815]) & (layer1_outputs[2541]);
    assign layer2_outputs[3606] = ~(layer1_outputs[2153]) | (layer1_outputs[228]);
    assign layer2_outputs[3607] = 1'b1;
    assign layer2_outputs[3608] = ~(layer1_outputs[3559]) | (layer1_outputs[935]);
    assign layer2_outputs[3609] = 1'b1;
    assign layer2_outputs[3610] = (layer1_outputs[3445]) & ~(layer1_outputs[4015]);
    assign layer2_outputs[3611] = 1'b1;
    assign layer2_outputs[3612] = 1'b1;
    assign layer2_outputs[3613] = layer1_outputs[2843];
    assign layer2_outputs[3614] = layer1_outputs[1963];
    assign layer2_outputs[3615] = layer1_outputs[499];
    assign layer2_outputs[3616] = (layer1_outputs[2126]) & ~(layer1_outputs[1909]);
    assign layer2_outputs[3617] = 1'b0;
    assign layer2_outputs[3618] = ~(layer1_outputs[1171]) | (layer1_outputs[5058]);
    assign layer2_outputs[3619] = (layer1_outputs[2422]) & (layer1_outputs[1153]);
    assign layer2_outputs[3620] = (layer1_outputs[4743]) & ~(layer1_outputs[2728]);
    assign layer2_outputs[3621] = 1'b0;
    assign layer2_outputs[3622] = layer1_outputs[4720];
    assign layer2_outputs[3623] = ~(layer1_outputs[4980]) | (layer1_outputs[1338]);
    assign layer2_outputs[3624] = (layer1_outputs[260]) | (layer1_outputs[4473]);
    assign layer2_outputs[3625] = (layer1_outputs[750]) & ~(layer1_outputs[630]);
    assign layer2_outputs[3626] = layer1_outputs[767];
    assign layer2_outputs[3627] = ~(layer1_outputs[2109]);
    assign layer2_outputs[3628] = (layer1_outputs[2867]) & ~(layer1_outputs[1366]);
    assign layer2_outputs[3629] = (layer1_outputs[286]) & ~(layer1_outputs[1568]);
    assign layer2_outputs[3630] = ~(layer1_outputs[4488]) | (layer1_outputs[1560]);
    assign layer2_outputs[3631] = layer1_outputs[1067];
    assign layer2_outputs[3632] = ~(layer1_outputs[2587]) | (layer1_outputs[2147]);
    assign layer2_outputs[3633] = ~(layer1_outputs[1778]) | (layer1_outputs[3483]);
    assign layer2_outputs[3634] = ~(layer1_outputs[1964]);
    assign layer2_outputs[3635] = ~(layer1_outputs[340]) | (layer1_outputs[2455]);
    assign layer2_outputs[3636] = ~(layer1_outputs[1928]) | (layer1_outputs[4867]);
    assign layer2_outputs[3637] = ~((layer1_outputs[3560]) | (layer1_outputs[3716]));
    assign layer2_outputs[3638] = layer1_outputs[2058];
    assign layer2_outputs[3639] = ~(layer1_outputs[4022]);
    assign layer2_outputs[3640] = 1'b1;
    assign layer2_outputs[3641] = ~((layer1_outputs[3551]) & (layer1_outputs[711]));
    assign layer2_outputs[3642] = (layer1_outputs[987]) & ~(layer1_outputs[3200]);
    assign layer2_outputs[3643] = (layer1_outputs[3873]) & ~(layer1_outputs[4589]);
    assign layer2_outputs[3644] = (layer1_outputs[1274]) & ~(layer1_outputs[3172]);
    assign layer2_outputs[3645] = ~(layer1_outputs[2535]);
    assign layer2_outputs[3646] = ~(layer1_outputs[2021]);
    assign layer2_outputs[3647] = ~(layer1_outputs[2053]) | (layer1_outputs[1696]);
    assign layer2_outputs[3648] = ~((layer1_outputs[3268]) & (layer1_outputs[2428]));
    assign layer2_outputs[3649] = 1'b1;
    assign layer2_outputs[3650] = (layer1_outputs[2959]) ^ (layer1_outputs[2595]);
    assign layer2_outputs[3651] = 1'b1;
    assign layer2_outputs[3652] = 1'b1;
    assign layer2_outputs[3653] = 1'b1;
    assign layer2_outputs[3654] = (layer1_outputs[97]) & (layer1_outputs[452]);
    assign layer2_outputs[3655] = ~((layer1_outputs[4814]) | (layer1_outputs[1744]));
    assign layer2_outputs[3656] = ~((layer1_outputs[1103]) | (layer1_outputs[1402]));
    assign layer2_outputs[3657] = ~(layer1_outputs[4610]) | (layer1_outputs[2259]);
    assign layer2_outputs[3658] = layer1_outputs[3915];
    assign layer2_outputs[3659] = ~(layer1_outputs[1083]) | (layer1_outputs[5109]);
    assign layer2_outputs[3660] = layer1_outputs[2419];
    assign layer2_outputs[3661] = layer1_outputs[2027];
    assign layer2_outputs[3662] = (layer1_outputs[3285]) & ~(layer1_outputs[2769]);
    assign layer2_outputs[3663] = ~(layer1_outputs[4241]);
    assign layer2_outputs[3664] = ~(layer1_outputs[2246]) | (layer1_outputs[1979]);
    assign layer2_outputs[3665] = 1'b0;
    assign layer2_outputs[3666] = layer1_outputs[4632];
    assign layer2_outputs[3667] = 1'b1;
    assign layer2_outputs[3668] = ~(layer1_outputs[3545]) | (layer1_outputs[1513]);
    assign layer2_outputs[3669] = (layer1_outputs[1692]) & ~(layer1_outputs[3979]);
    assign layer2_outputs[3670] = 1'b0;
    assign layer2_outputs[3671] = layer1_outputs[3573];
    assign layer2_outputs[3672] = ~(layer1_outputs[3534]) | (layer1_outputs[2122]);
    assign layer2_outputs[3673] = ~((layer1_outputs[2603]) ^ (layer1_outputs[878]));
    assign layer2_outputs[3674] = (layer1_outputs[1676]) | (layer1_outputs[939]);
    assign layer2_outputs[3675] = (layer1_outputs[711]) & ~(layer1_outputs[66]);
    assign layer2_outputs[3676] = layer1_outputs[4475];
    assign layer2_outputs[3677] = ~(layer1_outputs[3396]);
    assign layer2_outputs[3678] = ~(layer1_outputs[1812]) | (layer1_outputs[3941]);
    assign layer2_outputs[3679] = layer1_outputs[3645];
    assign layer2_outputs[3680] = layer1_outputs[1420];
    assign layer2_outputs[3681] = ~(layer1_outputs[4714]);
    assign layer2_outputs[3682] = (layer1_outputs[4891]) | (layer1_outputs[2115]);
    assign layer2_outputs[3683] = 1'b0;
    assign layer2_outputs[3684] = ~(layer1_outputs[3489]) | (layer1_outputs[1880]);
    assign layer2_outputs[3685] = ~(layer1_outputs[884]) | (layer1_outputs[2750]);
    assign layer2_outputs[3686] = ~((layer1_outputs[2313]) & (layer1_outputs[4667]));
    assign layer2_outputs[3687] = layer1_outputs[2478];
    assign layer2_outputs[3688] = ~(layer1_outputs[1781]);
    assign layer2_outputs[3689] = (layer1_outputs[3482]) | (layer1_outputs[93]);
    assign layer2_outputs[3690] = layer1_outputs[2765];
    assign layer2_outputs[3691] = 1'b0;
    assign layer2_outputs[3692] = (layer1_outputs[3105]) & ~(layer1_outputs[4152]);
    assign layer2_outputs[3693] = (layer1_outputs[4403]) & (layer1_outputs[3667]);
    assign layer2_outputs[3694] = layer1_outputs[901];
    assign layer2_outputs[3695] = layer1_outputs[918];
    assign layer2_outputs[3696] = ~(layer1_outputs[4444]);
    assign layer2_outputs[3697] = ~((layer1_outputs[3235]) & (layer1_outputs[2873]));
    assign layer2_outputs[3698] = (layer1_outputs[4333]) & ~(layer1_outputs[3730]);
    assign layer2_outputs[3699] = layer1_outputs[3492];
    assign layer2_outputs[3700] = layer1_outputs[4126];
    assign layer2_outputs[3701] = ~(layer1_outputs[2865]);
    assign layer2_outputs[3702] = ~(layer1_outputs[2214]);
    assign layer2_outputs[3703] = ~((layer1_outputs[2437]) | (layer1_outputs[360]));
    assign layer2_outputs[3704] = layer1_outputs[3397];
    assign layer2_outputs[3705] = (layer1_outputs[3585]) & (layer1_outputs[409]);
    assign layer2_outputs[3706] = 1'b0;
    assign layer2_outputs[3707] = ~(layer1_outputs[326]) | (layer1_outputs[3549]);
    assign layer2_outputs[3708] = ~(layer1_outputs[2649]);
    assign layer2_outputs[3709] = layer1_outputs[773];
    assign layer2_outputs[3710] = ~((layer1_outputs[523]) & (layer1_outputs[4219]));
    assign layer2_outputs[3711] = 1'b1;
    assign layer2_outputs[3712] = layer1_outputs[2922];
    assign layer2_outputs[3713] = layer1_outputs[3296];
    assign layer2_outputs[3714] = 1'b1;
    assign layer2_outputs[3715] = layer1_outputs[2108];
    assign layer2_outputs[3716] = ~((layer1_outputs[1797]) & (layer1_outputs[3412]));
    assign layer2_outputs[3717] = layer1_outputs[2019];
    assign layer2_outputs[3718] = 1'b1;
    assign layer2_outputs[3719] = ~(layer1_outputs[1038]);
    assign layer2_outputs[3720] = ~(layer1_outputs[1303]) | (layer1_outputs[2749]);
    assign layer2_outputs[3721] = ~(layer1_outputs[3622]) | (layer1_outputs[999]);
    assign layer2_outputs[3722] = (layer1_outputs[708]) | (layer1_outputs[871]);
    assign layer2_outputs[3723] = layer1_outputs[895];
    assign layer2_outputs[3724] = ~(layer1_outputs[4139]) | (layer1_outputs[2759]);
    assign layer2_outputs[3725] = layer1_outputs[2789];
    assign layer2_outputs[3726] = (layer1_outputs[4681]) | (layer1_outputs[3309]);
    assign layer2_outputs[3727] = ~(layer1_outputs[3582]);
    assign layer2_outputs[3728] = (layer1_outputs[3194]) | (layer1_outputs[527]);
    assign layer2_outputs[3729] = (layer1_outputs[1183]) & ~(layer1_outputs[2129]);
    assign layer2_outputs[3730] = 1'b0;
    assign layer2_outputs[3731] = (layer1_outputs[4342]) | (layer1_outputs[1932]);
    assign layer2_outputs[3732] = 1'b1;
    assign layer2_outputs[3733] = ~(layer1_outputs[2449]);
    assign layer2_outputs[3734] = (layer1_outputs[1684]) & (layer1_outputs[3211]);
    assign layer2_outputs[3735] = layer1_outputs[1924];
    assign layer2_outputs[3736] = layer1_outputs[1648];
    assign layer2_outputs[3737] = (layer1_outputs[90]) & (layer1_outputs[3673]);
    assign layer2_outputs[3738] = ~((layer1_outputs[4668]) | (layer1_outputs[4983]));
    assign layer2_outputs[3739] = ~(layer1_outputs[4253]) | (layer1_outputs[2007]);
    assign layer2_outputs[3740] = 1'b0;
    assign layer2_outputs[3741] = ~(layer1_outputs[651]) | (layer1_outputs[767]);
    assign layer2_outputs[3742] = ~(layer1_outputs[3350]);
    assign layer2_outputs[3743] = 1'b0;
    assign layer2_outputs[3744] = (layer1_outputs[140]) & ~(layer1_outputs[2144]);
    assign layer2_outputs[3745] = (layer1_outputs[1770]) & ~(layer1_outputs[2967]);
    assign layer2_outputs[3746] = (layer1_outputs[961]) ^ (layer1_outputs[2502]);
    assign layer2_outputs[3747] = ~((layer1_outputs[500]) | (layer1_outputs[1018]));
    assign layer2_outputs[3748] = (layer1_outputs[2392]) & (layer1_outputs[2002]);
    assign layer2_outputs[3749] = ~((layer1_outputs[4824]) | (layer1_outputs[4626]));
    assign layer2_outputs[3750] = (layer1_outputs[4062]) & (layer1_outputs[581]);
    assign layer2_outputs[3751] = 1'b1;
    assign layer2_outputs[3752] = ~(layer1_outputs[3380]) | (layer1_outputs[4158]);
    assign layer2_outputs[3753] = (layer1_outputs[1261]) & ~(layer1_outputs[4645]);
    assign layer2_outputs[3754] = ~(layer1_outputs[224]) | (layer1_outputs[4950]);
    assign layer2_outputs[3755] = ~(layer1_outputs[5018]) | (layer1_outputs[479]);
    assign layer2_outputs[3756] = (layer1_outputs[2570]) | (layer1_outputs[2148]);
    assign layer2_outputs[3757] = ~((layer1_outputs[1936]) | (layer1_outputs[3145]));
    assign layer2_outputs[3758] = ~((layer1_outputs[2480]) | (layer1_outputs[383]));
    assign layer2_outputs[3759] = ~(layer1_outputs[543]);
    assign layer2_outputs[3760] = (layer1_outputs[190]) | (layer1_outputs[2394]);
    assign layer2_outputs[3761] = ~(layer1_outputs[4340]);
    assign layer2_outputs[3762] = layer1_outputs[4501];
    assign layer2_outputs[3763] = ~(layer1_outputs[1883]);
    assign layer2_outputs[3764] = ~(layer1_outputs[4761]);
    assign layer2_outputs[3765] = ~(layer1_outputs[1394]);
    assign layer2_outputs[3766] = (layer1_outputs[4635]) & ~(layer1_outputs[447]);
    assign layer2_outputs[3767] = layer1_outputs[4657];
    assign layer2_outputs[3768] = (layer1_outputs[1513]) & (layer1_outputs[273]);
    assign layer2_outputs[3769] = ~(layer1_outputs[4843]) | (layer1_outputs[2849]);
    assign layer2_outputs[3770] = ~(layer1_outputs[5059]);
    assign layer2_outputs[3771] = ~((layer1_outputs[3381]) | (layer1_outputs[1491]));
    assign layer2_outputs[3772] = ~(layer1_outputs[3955]);
    assign layer2_outputs[3773] = (layer1_outputs[2415]) & (layer1_outputs[4368]);
    assign layer2_outputs[3774] = ~((layer1_outputs[3867]) | (layer1_outputs[1483]));
    assign layer2_outputs[3775] = 1'b1;
    assign layer2_outputs[3776] = 1'b0;
    assign layer2_outputs[3777] = ~((layer1_outputs[4033]) & (layer1_outputs[279]));
    assign layer2_outputs[3778] = 1'b0;
    assign layer2_outputs[3779] = (layer1_outputs[1519]) | (layer1_outputs[4790]);
    assign layer2_outputs[3780] = layer1_outputs[3339];
    assign layer2_outputs[3781] = 1'b0;
    assign layer2_outputs[3782] = ~((layer1_outputs[5035]) | (layer1_outputs[3131]));
    assign layer2_outputs[3783] = (layer1_outputs[4300]) & (layer1_outputs[1559]);
    assign layer2_outputs[3784] = ~(layer1_outputs[2701]);
    assign layer2_outputs[3785] = (layer1_outputs[3698]) & ~(layer1_outputs[2629]);
    assign layer2_outputs[3786] = 1'b0;
    assign layer2_outputs[3787] = (layer1_outputs[3012]) & (layer1_outputs[3889]);
    assign layer2_outputs[3788] = 1'b0;
    assign layer2_outputs[3789] = ~(layer1_outputs[2506]);
    assign layer2_outputs[3790] = ~((layer1_outputs[2330]) & (layer1_outputs[3564]));
    assign layer2_outputs[3791] = ~((layer1_outputs[1996]) | (layer1_outputs[760]));
    assign layer2_outputs[3792] = ~((layer1_outputs[4839]) | (layer1_outputs[3104]));
    assign layer2_outputs[3793] = ~(layer1_outputs[477]);
    assign layer2_outputs[3794] = (layer1_outputs[1637]) & ~(layer1_outputs[759]);
    assign layer2_outputs[3795] = (layer1_outputs[4660]) ^ (layer1_outputs[5118]);
    assign layer2_outputs[3796] = (layer1_outputs[3615]) & ~(layer1_outputs[2662]);
    assign layer2_outputs[3797] = layer1_outputs[3741];
    assign layer2_outputs[3798] = ~(layer1_outputs[1381]);
    assign layer2_outputs[3799] = layer1_outputs[3993];
    assign layer2_outputs[3800] = ~((layer1_outputs[3987]) & (layer1_outputs[1490]));
    assign layer2_outputs[3801] = (layer1_outputs[2034]) ^ (layer1_outputs[1897]);
    assign layer2_outputs[3802] = ~((layer1_outputs[4590]) | (layer1_outputs[1613]));
    assign layer2_outputs[3803] = ~(layer1_outputs[2159]);
    assign layer2_outputs[3804] = layer1_outputs[2778];
    assign layer2_outputs[3805] = 1'b1;
    assign layer2_outputs[3806] = ~((layer1_outputs[3742]) | (layer1_outputs[3599]));
    assign layer2_outputs[3807] = ~(layer1_outputs[4678]);
    assign layer2_outputs[3808] = ~(layer1_outputs[3526]) | (layer1_outputs[1772]);
    assign layer2_outputs[3809] = ~(layer1_outputs[2753]);
    assign layer2_outputs[3810] = ~(layer1_outputs[3126]);
    assign layer2_outputs[3811] = ~((layer1_outputs[1726]) & (layer1_outputs[2193]));
    assign layer2_outputs[3812] = 1'b0;
    assign layer2_outputs[3813] = ~(layer1_outputs[972]) | (layer1_outputs[3887]);
    assign layer2_outputs[3814] = ~(layer1_outputs[3519]);
    assign layer2_outputs[3815] = ~(layer1_outputs[180]);
    assign layer2_outputs[3816] = (layer1_outputs[4275]) | (layer1_outputs[974]);
    assign layer2_outputs[3817] = (layer1_outputs[4808]) & ~(layer1_outputs[3900]);
    assign layer2_outputs[3818] = (layer1_outputs[3084]) & (layer1_outputs[968]);
    assign layer2_outputs[3819] = layer1_outputs[68];
    assign layer2_outputs[3820] = (layer1_outputs[1201]) & (layer1_outputs[143]);
    assign layer2_outputs[3821] = (layer1_outputs[1757]) & (layer1_outputs[3866]);
    assign layer2_outputs[3822] = 1'b1;
    assign layer2_outputs[3823] = 1'b0;
    assign layer2_outputs[3824] = layer1_outputs[4216];
    assign layer2_outputs[3825] = ~((layer1_outputs[1645]) | (layer1_outputs[984]));
    assign layer2_outputs[3826] = (layer1_outputs[4168]) & ~(layer1_outputs[4393]);
    assign layer2_outputs[3827] = ~(layer1_outputs[748]);
    assign layer2_outputs[3828] = 1'b1;
    assign layer2_outputs[3829] = ~(layer1_outputs[908]);
    assign layer2_outputs[3830] = layer1_outputs[4543];
    assign layer2_outputs[3831] = ~((layer1_outputs[2087]) & (layer1_outputs[2823]));
    assign layer2_outputs[3832] = ~(layer1_outputs[4567]);
    assign layer2_outputs[3833] = layer1_outputs[2769];
    assign layer2_outputs[3834] = layer1_outputs[2215];
    assign layer2_outputs[3835] = (layer1_outputs[2746]) & (layer1_outputs[5086]);
    assign layer2_outputs[3836] = (layer1_outputs[3845]) & (layer1_outputs[640]);
    assign layer2_outputs[3837] = (layer1_outputs[3255]) & ~(layer1_outputs[1222]);
    assign layer2_outputs[3838] = (layer1_outputs[208]) | (layer1_outputs[4014]);
    assign layer2_outputs[3839] = layer1_outputs[3111];
    assign layer2_outputs[3840] = ~(layer1_outputs[191]) | (layer1_outputs[4846]);
    assign layer2_outputs[3841] = ~(layer1_outputs[5030]);
    assign layer2_outputs[3842] = (layer1_outputs[4062]) ^ (layer1_outputs[3953]);
    assign layer2_outputs[3843] = ~(layer1_outputs[3421]);
    assign layer2_outputs[3844] = ~((layer1_outputs[364]) & (layer1_outputs[1127]));
    assign layer2_outputs[3845] = ~((layer1_outputs[3096]) & (layer1_outputs[3699]));
    assign layer2_outputs[3846] = (layer1_outputs[1625]) ^ (layer1_outputs[735]);
    assign layer2_outputs[3847] = (layer1_outputs[549]) & ~(layer1_outputs[4322]);
    assign layer2_outputs[3848] = 1'b0;
    assign layer2_outputs[3849] = layer1_outputs[2832];
    assign layer2_outputs[3850] = (layer1_outputs[79]) & (layer1_outputs[2827]);
    assign layer2_outputs[3851] = ~((layer1_outputs[2796]) | (layer1_outputs[423]));
    assign layer2_outputs[3852] = layer1_outputs[789];
    assign layer2_outputs[3853] = layer1_outputs[4686];
    assign layer2_outputs[3854] = ~(layer1_outputs[2287]) | (layer1_outputs[2606]);
    assign layer2_outputs[3855] = (layer1_outputs[4247]) & ~(layer1_outputs[3522]);
    assign layer2_outputs[3856] = ~((layer1_outputs[2964]) & (layer1_outputs[3866]));
    assign layer2_outputs[3857] = ~(layer1_outputs[4819]);
    assign layer2_outputs[3858] = ~((layer1_outputs[4427]) ^ (layer1_outputs[775]));
    assign layer2_outputs[3859] = layer1_outputs[772];
    assign layer2_outputs[3860] = (layer1_outputs[4531]) & ~(layer1_outputs[2382]);
    assign layer2_outputs[3861] = (layer1_outputs[1446]) & ~(layer1_outputs[1404]);
    assign layer2_outputs[3862] = ~((layer1_outputs[243]) & (layer1_outputs[2363]));
    assign layer2_outputs[3863] = ~((layer1_outputs[1038]) ^ (layer1_outputs[1133]));
    assign layer2_outputs[3864] = ~(layer1_outputs[1352]);
    assign layer2_outputs[3865] = 1'b1;
    assign layer2_outputs[3866] = (layer1_outputs[1]) & ~(layer1_outputs[4982]);
    assign layer2_outputs[3867] = ~((layer1_outputs[3019]) | (layer1_outputs[3313]));
    assign layer2_outputs[3868] = ~(layer1_outputs[3390]);
    assign layer2_outputs[3869] = (layer1_outputs[1172]) | (layer1_outputs[3667]);
    assign layer2_outputs[3870] = layer1_outputs[3945];
    assign layer2_outputs[3871] = ~(layer1_outputs[2110]) | (layer1_outputs[381]);
    assign layer2_outputs[3872] = (layer1_outputs[828]) & (layer1_outputs[2749]);
    assign layer2_outputs[3873] = layer1_outputs[3107];
    assign layer2_outputs[3874] = 1'b1;
    assign layer2_outputs[3875] = ~((layer1_outputs[3700]) | (layer1_outputs[4728]));
    assign layer2_outputs[3876] = (layer1_outputs[3588]) | (layer1_outputs[4682]);
    assign layer2_outputs[3877] = (layer1_outputs[3449]) & ~(layer1_outputs[3182]);
    assign layer2_outputs[3878] = layer1_outputs[3328];
    assign layer2_outputs[3879] = ~(layer1_outputs[4564]);
    assign layer2_outputs[3880] = layer1_outputs[4396];
    assign layer2_outputs[3881] = (layer1_outputs[4071]) & (layer1_outputs[1470]);
    assign layer2_outputs[3882] = ~(layer1_outputs[967]) | (layer1_outputs[73]);
    assign layer2_outputs[3883] = ~((layer1_outputs[804]) | (layer1_outputs[4613]));
    assign layer2_outputs[3884] = 1'b0;
    assign layer2_outputs[3885] = (layer1_outputs[4769]) & (layer1_outputs[4549]);
    assign layer2_outputs[3886] = layer1_outputs[2286];
    assign layer2_outputs[3887] = ~(layer1_outputs[1544]);
    assign layer2_outputs[3888] = ~(layer1_outputs[764]) | (layer1_outputs[2065]);
    assign layer2_outputs[3889] = layer1_outputs[614];
    assign layer2_outputs[3890] = (layer1_outputs[4955]) & (layer1_outputs[3905]);
    assign layer2_outputs[3891] = 1'b0;
    assign layer2_outputs[3892] = ~((layer1_outputs[3807]) ^ (layer1_outputs[4525]));
    assign layer2_outputs[3893] = ~((layer1_outputs[3077]) | (layer1_outputs[1571]));
    assign layer2_outputs[3894] = ~(layer1_outputs[2897]);
    assign layer2_outputs[3895] = ~((layer1_outputs[4329]) ^ (layer1_outputs[1388]));
    assign layer2_outputs[3896] = layer1_outputs[653];
    assign layer2_outputs[3897] = ~(layer1_outputs[1007]) | (layer1_outputs[4202]);
    assign layer2_outputs[3898] = ~(layer1_outputs[4836]);
    assign layer2_outputs[3899] = 1'b0;
    assign layer2_outputs[3900] = 1'b1;
    assign layer2_outputs[3901] = ~((layer1_outputs[4339]) | (layer1_outputs[3280]));
    assign layer2_outputs[3902] = (layer1_outputs[5019]) & (layer1_outputs[5092]);
    assign layer2_outputs[3903] = layer1_outputs[4167];
    assign layer2_outputs[3904] = ~(layer1_outputs[1710]);
    assign layer2_outputs[3905] = (layer1_outputs[4658]) & ~(layer1_outputs[1200]);
    assign layer2_outputs[3906] = ~(layer1_outputs[4130]) | (layer1_outputs[1359]);
    assign layer2_outputs[3907] = (layer1_outputs[2726]) ^ (layer1_outputs[1734]);
    assign layer2_outputs[3908] = ~(layer1_outputs[4082]) | (layer1_outputs[3616]);
    assign layer2_outputs[3909] = layer1_outputs[3624];
    assign layer2_outputs[3910] = ~(layer1_outputs[3969]) | (layer1_outputs[4560]);
    assign layer2_outputs[3911] = layer1_outputs[3358];
    assign layer2_outputs[3912] = (layer1_outputs[3292]) & (layer1_outputs[1795]);
    assign layer2_outputs[3913] = (layer1_outputs[3819]) & ~(layer1_outputs[713]);
    assign layer2_outputs[3914] = (layer1_outputs[252]) & ~(layer1_outputs[1669]);
    assign layer2_outputs[3915] = ~(layer1_outputs[2976]);
    assign layer2_outputs[3916] = ~(layer1_outputs[3568]);
    assign layer2_outputs[3917] = 1'b1;
    assign layer2_outputs[3918] = layer1_outputs[4481];
    assign layer2_outputs[3919] = (layer1_outputs[3177]) & ~(layer1_outputs[4308]);
    assign layer2_outputs[3920] = ~(layer1_outputs[3694]) | (layer1_outputs[3723]);
    assign layer2_outputs[3921] = layer1_outputs[106];
    assign layer2_outputs[3922] = (layer1_outputs[2475]) & ~(layer1_outputs[1579]);
    assign layer2_outputs[3923] = ~(layer1_outputs[3269]) | (layer1_outputs[3222]);
    assign layer2_outputs[3924] = 1'b0;
    assign layer2_outputs[3925] = ~((layer1_outputs[2941]) | (layer1_outputs[2699]));
    assign layer2_outputs[3926] = ~(layer1_outputs[4186]) | (layer1_outputs[4144]);
    assign layer2_outputs[3927] = ~(layer1_outputs[2066]);
    assign layer2_outputs[3928] = ~(layer1_outputs[1301]);
    assign layer2_outputs[3929] = ~(layer1_outputs[4157]);
    assign layer2_outputs[3930] = ~(layer1_outputs[2134]);
    assign layer2_outputs[3931] = ~(layer1_outputs[1107]);
    assign layer2_outputs[3932] = (layer1_outputs[3458]) & ~(layer1_outputs[661]);
    assign layer2_outputs[3933] = ~((layer1_outputs[3393]) & (layer1_outputs[1671]));
    assign layer2_outputs[3934] = (layer1_outputs[4597]) & (layer1_outputs[569]);
    assign layer2_outputs[3935] = ~((layer1_outputs[707]) & (layer1_outputs[3489]));
    assign layer2_outputs[3936] = 1'b0;
    assign layer2_outputs[3937] = layer1_outputs[38];
    assign layer2_outputs[3938] = 1'b0;
    assign layer2_outputs[3939] = ~(layer1_outputs[4278]) | (layer1_outputs[2489]);
    assign layer2_outputs[3940] = ~((layer1_outputs[731]) & (layer1_outputs[391]));
    assign layer2_outputs[3941] = ~((layer1_outputs[2990]) & (layer1_outputs[1590]));
    assign layer2_outputs[3942] = ~(layer1_outputs[25]) | (layer1_outputs[2590]);
    assign layer2_outputs[3943] = ~((layer1_outputs[2171]) & (layer1_outputs[3487]));
    assign layer2_outputs[3944] = layer1_outputs[2030];
    assign layer2_outputs[3945] = ~((layer1_outputs[4476]) & (layer1_outputs[1322]));
    assign layer2_outputs[3946] = ~(layer1_outputs[2519]);
    assign layer2_outputs[3947] = layer1_outputs[2346];
    assign layer2_outputs[3948] = layer1_outputs[2930];
    assign layer2_outputs[3949] = layer1_outputs[3811];
    assign layer2_outputs[3950] = layer1_outputs[5];
    assign layer2_outputs[3951] = ~(layer1_outputs[2321]) | (layer1_outputs[950]);
    assign layer2_outputs[3952] = layer1_outputs[475];
    assign layer2_outputs[3953] = (layer1_outputs[1714]) & (layer1_outputs[4547]);
    assign layer2_outputs[3954] = (layer1_outputs[2816]) & (layer1_outputs[2246]);
    assign layer2_outputs[3955] = (layer1_outputs[3399]) & ~(layer1_outputs[3905]);
    assign layer2_outputs[3956] = 1'b0;
    assign layer2_outputs[3957] = layer1_outputs[3662];
    assign layer2_outputs[3958] = (layer1_outputs[997]) & ~(layer1_outputs[4517]);
    assign layer2_outputs[3959] = (layer1_outputs[1617]) | (layer1_outputs[4820]);
    assign layer2_outputs[3960] = ~((layer1_outputs[3541]) & (layer1_outputs[1954]));
    assign layer2_outputs[3961] = ~((layer1_outputs[3332]) ^ (layer1_outputs[3513]));
    assign layer2_outputs[3962] = ~(layer1_outputs[3889]) | (layer1_outputs[763]);
    assign layer2_outputs[3963] = ~((layer1_outputs[716]) | (layer1_outputs[2774]));
    assign layer2_outputs[3964] = ~(layer1_outputs[3065]);
    assign layer2_outputs[3965] = layer1_outputs[2793];
    assign layer2_outputs[3966] = ~(layer1_outputs[2649]);
    assign layer2_outputs[3967] = ~(layer1_outputs[2693]);
    assign layer2_outputs[3968] = (layer1_outputs[1158]) & ~(layer1_outputs[3965]);
    assign layer2_outputs[3969] = 1'b0;
    assign layer2_outputs[3970] = 1'b0;
    assign layer2_outputs[3971] = layer1_outputs[3601];
    assign layer2_outputs[3972] = 1'b0;
    assign layer2_outputs[3973] = ~((layer1_outputs[58]) | (layer1_outputs[3338]));
    assign layer2_outputs[3974] = (layer1_outputs[2335]) & ~(layer1_outputs[1642]);
    assign layer2_outputs[3975] = (layer1_outputs[5048]) & ~(layer1_outputs[1264]);
    assign layer2_outputs[3976] = (layer1_outputs[628]) & (layer1_outputs[3319]);
    assign layer2_outputs[3977] = ~((layer1_outputs[4369]) | (layer1_outputs[1064]));
    assign layer2_outputs[3978] = (layer1_outputs[3351]) & ~(layer1_outputs[3671]);
    assign layer2_outputs[3979] = ~((layer1_outputs[3418]) & (layer1_outputs[3524]));
    assign layer2_outputs[3980] = ~((layer1_outputs[3341]) | (layer1_outputs[2499]));
    assign layer2_outputs[3981] = ~((layer1_outputs[4330]) | (layer1_outputs[2420]));
    assign layer2_outputs[3982] = ~(layer1_outputs[1844]);
    assign layer2_outputs[3983] = (layer1_outputs[1692]) & ~(layer1_outputs[4868]);
    assign layer2_outputs[3984] = ~(layer1_outputs[1979]);
    assign layer2_outputs[3985] = layer1_outputs[4345];
    assign layer2_outputs[3986] = ~(layer1_outputs[29]);
    assign layer2_outputs[3987] = 1'b0;
    assign layer2_outputs[3988] = ~(layer1_outputs[3511]) | (layer1_outputs[1443]);
    assign layer2_outputs[3989] = 1'b1;
    assign layer2_outputs[3990] = 1'b0;
    assign layer2_outputs[3991] = ~(layer1_outputs[3820]);
    assign layer2_outputs[3992] = 1'b1;
    assign layer2_outputs[3993] = ~((layer1_outputs[1497]) | (layer1_outputs[3247]));
    assign layer2_outputs[3994] = ~((layer1_outputs[464]) | (layer1_outputs[3366]));
    assign layer2_outputs[3995] = (layer1_outputs[3383]) & (layer1_outputs[2956]);
    assign layer2_outputs[3996] = (layer1_outputs[2133]) & ~(layer1_outputs[725]);
    assign layer2_outputs[3997] = 1'b0;
    assign layer2_outputs[3998] = 1'b0;
    assign layer2_outputs[3999] = ~(layer1_outputs[1399]);
    assign layer2_outputs[4000] = (layer1_outputs[4508]) & ~(layer1_outputs[601]);
    assign layer2_outputs[4001] = ~(layer1_outputs[100]);
    assign layer2_outputs[4002] = 1'b0;
    assign layer2_outputs[4003] = (layer1_outputs[3420]) & ~(layer1_outputs[2696]);
    assign layer2_outputs[4004] = layer1_outputs[1165];
    assign layer2_outputs[4005] = (layer1_outputs[4287]) & ~(layer1_outputs[1897]);
    assign layer2_outputs[4006] = (layer1_outputs[1311]) | (layer1_outputs[91]);
    assign layer2_outputs[4007] = ~(layer1_outputs[682]);
    assign layer2_outputs[4008] = ~(layer1_outputs[2380]);
    assign layer2_outputs[4009] = (layer1_outputs[2315]) & ~(layer1_outputs[4725]);
    assign layer2_outputs[4010] = 1'b0;
    assign layer2_outputs[4011] = ~(layer1_outputs[1305]) | (layer1_outputs[741]);
    assign layer2_outputs[4012] = ~(layer1_outputs[739]) | (layer1_outputs[2596]);
    assign layer2_outputs[4013] = (layer1_outputs[69]) | (layer1_outputs[3926]);
    assign layer2_outputs[4014] = (layer1_outputs[1109]) & (layer1_outputs[4466]);
    assign layer2_outputs[4015] = 1'b1;
    assign layer2_outputs[4016] = (layer1_outputs[1748]) & (layer1_outputs[2999]);
    assign layer2_outputs[4017] = ~(layer1_outputs[1898]);
    assign layer2_outputs[4018] = layer1_outputs[980];
    assign layer2_outputs[4019] = ~(layer1_outputs[1095]);
    assign layer2_outputs[4020] = layer1_outputs[2908];
    assign layer2_outputs[4021] = layer1_outputs[2351];
    assign layer2_outputs[4022] = (layer1_outputs[5100]) | (layer1_outputs[508]);
    assign layer2_outputs[4023] = (layer1_outputs[4375]) | (layer1_outputs[4417]);
    assign layer2_outputs[4024] = layer1_outputs[4355];
    assign layer2_outputs[4025] = ~(layer1_outputs[765]);
    assign layer2_outputs[4026] = ~(layer1_outputs[1064]) | (layer1_outputs[2437]);
    assign layer2_outputs[4027] = ~(layer1_outputs[768]) | (layer1_outputs[4855]);
    assign layer2_outputs[4028] = ~(layer1_outputs[2294]);
    assign layer2_outputs[4029] = ~((layer1_outputs[3081]) | (layer1_outputs[4730]));
    assign layer2_outputs[4030] = ~(layer1_outputs[4758]);
    assign layer2_outputs[4031] = ~((layer1_outputs[644]) | (layer1_outputs[660]));
    assign layer2_outputs[4032] = (layer1_outputs[2559]) & ~(layer1_outputs[4435]);
    assign layer2_outputs[4033] = 1'b1;
    assign layer2_outputs[4034] = ~(layer1_outputs[2704]) | (layer1_outputs[1277]);
    assign layer2_outputs[4035] = (layer1_outputs[1791]) | (layer1_outputs[1150]);
    assign layer2_outputs[4036] = ~(layer1_outputs[1960]) | (layer1_outputs[231]);
    assign layer2_outputs[4037] = (layer1_outputs[4038]) ^ (layer1_outputs[2079]);
    assign layer2_outputs[4038] = (layer1_outputs[2658]) & (layer1_outputs[5082]);
    assign layer2_outputs[4039] = (layer1_outputs[4636]) & ~(layer1_outputs[916]);
    assign layer2_outputs[4040] = ~((layer1_outputs[2613]) & (layer1_outputs[343]));
    assign layer2_outputs[4041] = (layer1_outputs[2084]) | (layer1_outputs[4350]);
    assign layer2_outputs[4042] = ~((layer1_outputs[1423]) | (layer1_outputs[2426]));
    assign layer2_outputs[4043] = layer1_outputs[2163];
    assign layer2_outputs[4044] = 1'b1;
    assign layer2_outputs[4045] = layer1_outputs[3825];
    assign layer2_outputs[4046] = layer1_outputs[3061];
    assign layer2_outputs[4047] = ~((layer1_outputs[2618]) & (layer1_outputs[102]));
    assign layer2_outputs[4048] = (layer1_outputs[1031]) & ~(layer1_outputs[4588]);
    assign layer2_outputs[4049] = 1'b0;
    assign layer2_outputs[4050] = ~(layer1_outputs[2712]);
    assign layer2_outputs[4051] = ~(layer1_outputs[5091]) | (layer1_outputs[3163]);
    assign layer2_outputs[4052] = layer1_outputs[3399];
    assign layer2_outputs[4053] = 1'b0;
    assign layer2_outputs[4054] = 1'b1;
    assign layer2_outputs[4055] = 1'b0;
    assign layer2_outputs[4056] = 1'b0;
    assign layer2_outputs[4057] = (layer1_outputs[2355]) | (layer1_outputs[2593]);
    assign layer2_outputs[4058] = ~((layer1_outputs[1002]) & (layer1_outputs[3562]));
    assign layer2_outputs[4059] = ~((layer1_outputs[4462]) | (layer1_outputs[3789]));
    assign layer2_outputs[4060] = ~((layer1_outputs[3863]) & (layer1_outputs[4514]));
    assign layer2_outputs[4061] = ~(layer1_outputs[142]) | (layer1_outputs[2300]);
    assign layer2_outputs[4062] = ~(layer1_outputs[1666]) | (layer1_outputs[4084]);
    assign layer2_outputs[4063] = ~((layer1_outputs[4845]) | (layer1_outputs[122]));
    assign layer2_outputs[4064] = (layer1_outputs[2179]) & ~(layer1_outputs[2818]);
    assign layer2_outputs[4065] = layer1_outputs[1914];
    assign layer2_outputs[4066] = layer1_outputs[1814];
    assign layer2_outputs[4067] = (layer1_outputs[1463]) & ~(layer1_outputs[1340]);
    assign layer2_outputs[4068] = (layer1_outputs[5022]) & ~(layer1_outputs[4766]);
    assign layer2_outputs[4069] = ~((layer1_outputs[298]) & (layer1_outputs[3020]));
    assign layer2_outputs[4070] = 1'b0;
    assign layer2_outputs[4071] = ~(layer1_outputs[3753]) | (layer1_outputs[1206]);
    assign layer2_outputs[4072] = (layer1_outputs[2063]) & (layer1_outputs[791]);
    assign layer2_outputs[4073] = ~(layer1_outputs[4141]);
    assign layer2_outputs[4074] = ~(layer1_outputs[34]);
    assign layer2_outputs[4075] = ~(layer1_outputs[2051]) | (layer1_outputs[5105]);
    assign layer2_outputs[4076] = (layer1_outputs[4900]) & ~(layer1_outputs[235]);
    assign layer2_outputs[4077] = layer1_outputs[1649];
    assign layer2_outputs[4078] = layer1_outputs[3353];
    assign layer2_outputs[4079] = (layer1_outputs[1019]) & (layer1_outputs[4873]);
    assign layer2_outputs[4080] = ~(layer1_outputs[3294]) | (layer1_outputs[4151]);
    assign layer2_outputs[4081] = layer1_outputs[1634];
    assign layer2_outputs[4082] = layer1_outputs[3943];
    assign layer2_outputs[4083] = 1'b0;
    assign layer2_outputs[4084] = ~((layer1_outputs[3857]) & (layer1_outputs[1030]));
    assign layer2_outputs[4085] = 1'b1;
    assign layer2_outputs[4086] = (layer1_outputs[3904]) & ~(layer1_outputs[2681]);
    assign layer2_outputs[4087] = ~((layer1_outputs[4175]) | (layer1_outputs[3242]));
    assign layer2_outputs[4088] = ~(layer1_outputs[1180]) | (layer1_outputs[3193]);
    assign layer2_outputs[4089] = ~((layer1_outputs[688]) & (layer1_outputs[2167]));
    assign layer2_outputs[4090] = (layer1_outputs[2501]) & ~(layer1_outputs[4926]);
    assign layer2_outputs[4091] = ~((layer1_outputs[2000]) | (layer1_outputs[2483]));
    assign layer2_outputs[4092] = ~(layer1_outputs[4680]) | (layer1_outputs[3461]);
    assign layer2_outputs[4093] = ~((layer1_outputs[902]) & (layer1_outputs[3874]));
    assign layer2_outputs[4094] = ~((layer1_outputs[4960]) & (layer1_outputs[5007]));
    assign layer2_outputs[4095] = layer1_outputs[3881];
    assign layer2_outputs[4096] = 1'b1;
    assign layer2_outputs[4097] = ~(layer1_outputs[519]);
    assign layer2_outputs[4098] = 1'b1;
    assign layer2_outputs[4099] = ~(layer1_outputs[3137]) | (layer1_outputs[3135]);
    assign layer2_outputs[4100] = ~(layer1_outputs[2412]);
    assign layer2_outputs[4101] = (layer1_outputs[3273]) & (layer1_outputs[3587]);
    assign layer2_outputs[4102] = layer1_outputs[250];
    assign layer2_outputs[4103] = ~((layer1_outputs[179]) | (layer1_outputs[1226]));
    assign layer2_outputs[4104] = ~((layer1_outputs[3217]) | (layer1_outputs[3679]));
    assign layer2_outputs[4105] = ~(layer1_outputs[3325]);
    assign layer2_outputs[4106] = (layer1_outputs[3670]) | (layer1_outputs[3292]);
    assign layer2_outputs[4107] = (layer1_outputs[1737]) | (layer1_outputs[1062]);
    assign layer2_outputs[4108] = ~((layer1_outputs[684]) | (layer1_outputs[4468]));
    assign layer2_outputs[4109] = layer1_outputs[200];
    assign layer2_outputs[4110] = 1'b0;
    assign layer2_outputs[4111] = (layer1_outputs[492]) & (layer1_outputs[1960]);
    assign layer2_outputs[4112] = ~((layer1_outputs[4553]) & (layer1_outputs[2212]));
    assign layer2_outputs[4113] = ~(layer1_outputs[1572]) | (layer1_outputs[3686]);
    assign layer2_outputs[4114] = ~(layer1_outputs[2744]);
    assign layer2_outputs[4115] = (layer1_outputs[1426]) & ~(layer1_outputs[2477]);
    assign layer2_outputs[4116] = 1'b1;
    assign layer2_outputs[4117] = ~(layer1_outputs[1393]);
    assign layer2_outputs[4118] = 1'b1;
    assign layer2_outputs[4119] = layer1_outputs[5068];
    assign layer2_outputs[4120] = ~((layer1_outputs[3446]) | (layer1_outputs[3155]));
    assign layer2_outputs[4121] = (layer1_outputs[3537]) & ~(layer1_outputs[1179]);
    assign layer2_outputs[4122] = ~(layer1_outputs[2190]) | (layer1_outputs[1097]);
    assign layer2_outputs[4123] = ~(layer1_outputs[975]) | (layer1_outputs[3519]);
    assign layer2_outputs[4124] = 1'b1;
    assign layer2_outputs[4125] = 1'b0;
    assign layer2_outputs[4126] = (layer1_outputs[4611]) & ~(layer1_outputs[3402]);
    assign layer2_outputs[4127] = ~(layer1_outputs[2510]);
    assign layer2_outputs[4128] = (layer1_outputs[2210]) | (layer1_outputs[2142]);
    assign layer2_outputs[4129] = 1'b1;
    assign layer2_outputs[4130] = layer1_outputs[2357];
    assign layer2_outputs[4131] = (layer1_outputs[2623]) ^ (layer1_outputs[3397]);
    assign layer2_outputs[4132] = 1'b0;
    assign layer2_outputs[4133] = ~((layer1_outputs[4599]) | (layer1_outputs[539]));
    assign layer2_outputs[4134] = ~((layer1_outputs[4899]) | (layer1_outputs[2269]));
    assign layer2_outputs[4135] = 1'b1;
    assign layer2_outputs[4136] = 1'b1;
    assign layer2_outputs[4137] = ~((layer1_outputs[2925]) | (layer1_outputs[4917]));
    assign layer2_outputs[4138] = ~((layer1_outputs[2542]) | (layer1_outputs[1377]));
    assign layer2_outputs[4139] = ~(layer1_outputs[2936]);
    assign layer2_outputs[4140] = layer1_outputs[160];
    assign layer2_outputs[4141] = 1'b0;
    assign layer2_outputs[4142] = (layer1_outputs[1581]) & ~(layer1_outputs[184]);
    assign layer2_outputs[4143] = ~(layer1_outputs[2771]);
    assign layer2_outputs[4144] = (layer1_outputs[1445]) & (layer1_outputs[3930]);
    assign layer2_outputs[4145] = (layer1_outputs[2092]) & ~(layer1_outputs[4344]);
    assign layer2_outputs[4146] = ~((layer1_outputs[360]) & (layer1_outputs[278]));
    assign layer2_outputs[4147] = ~(layer1_outputs[3647]);
    assign layer2_outputs[4148] = (layer1_outputs[1698]) & (layer1_outputs[318]);
    assign layer2_outputs[4149] = (layer1_outputs[2550]) & (layer1_outputs[2226]);
    assign layer2_outputs[4150] = ~((layer1_outputs[570]) | (layer1_outputs[124]));
    assign layer2_outputs[4151] = (layer1_outputs[1741]) & ~(layer1_outputs[4227]);
    assign layer2_outputs[4152] = ~((layer1_outputs[1051]) ^ (layer1_outputs[4943]));
    assign layer2_outputs[4153] = (layer1_outputs[15]) | (layer1_outputs[1785]);
    assign layer2_outputs[4154] = (layer1_outputs[162]) & ~(layer1_outputs[717]);
    assign layer2_outputs[4155] = layer1_outputs[4376];
    assign layer2_outputs[4156] = (layer1_outputs[1366]) | (layer1_outputs[4969]);
    assign layer2_outputs[4157] = (layer1_outputs[4070]) | (layer1_outputs[1938]);
    assign layer2_outputs[4158] = 1'b1;
    assign layer2_outputs[4159] = 1'b1;
    assign layer2_outputs[4160] = (layer1_outputs[3799]) & (layer1_outputs[1722]);
    assign layer2_outputs[4161] = ~(layer1_outputs[4806]);
    assign layer2_outputs[4162] = 1'b0;
    assign layer2_outputs[4163] = (layer1_outputs[2734]) & (layer1_outputs[752]);
    assign layer2_outputs[4164] = (layer1_outputs[143]) | (layer1_outputs[2527]);
    assign layer2_outputs[4165] = (layer1_outputs[736]) & ~(layer1_outputs[4260]);
    assign layer2_outputs[4166] = ~(layer1_outputs[4060]);
    assign layer2_outputs[4167] = ~(layer1_outputs[4972]);
    assign layer2_outputs[4168] = ~(layer1_outputs[1420]);
    assign layer2_outputs[4169] = 1'b0;
    assign layer2_outputs[4170] = ~(layer1_outputs[1935]) | (layer1_outputs[2513]);
    assign layer2_outputs[4171] = 1'b0;
    assign layer2_outputs[4172] = (layer1_outputs[2556]) & (layer1_outputs[1400]);
    assign layer2_outputs[4173] = ~(layer1_outputs[4911]) | (layer1_outputs[3047]);
    assign layer2_outputs[4174] = (layer1_outputs[507]) & ~(layer1_outputs[3483]);
    assign layer2_outputs[4175] = ~(layer1_outputs[3816]);
    assign layer2_outputs[4176] = (layer1_outputs[33]) | (layer1_outputs[2189]);
    assign layer2_outputs[4177] = (layer1_outputs[3121]) & ~(layer1_outputs[2227]);
    assign layer2_outputs[4178] = layer1_outputs[1871];
    assign layer2_outputs[4179] = (layer1_outputs[3813]) & ~(layer1_outputs[2026]);
    assign layer2_outputs[4180] = ~((layer1_outputs[1562]) & (layer1_outputs[4156]));
    assign layer2_outputs[4181] = 1'b1;
    assign layer2_outputs[4182] = ~(layer1_outputs[3191]);
    assign layer2_outputs[4183] = 1'b1;
    assign layer2_outputs[4184] = layer1_outputs[3040];
    assign layer2_outputs[4185] = (layer1_outputs[1989]) & ~(layer1_outputs[3297]);
    assign layer2_outputs[4186] = ~(layer1_outputs[112]);
    assign layer2_outputs[4187] = (layer1_outputs[705]) & ~(layer1_outputs[4607]);
    assign layer2_outputs[4188] = 1'b0;
    assign layer2_outputs[4189] = (layer1_outputs[9]) & ~(layer1_outputs[276]);
    assign layer2_outputs[4190] = ~(layer1_outputs[154]) | (layer1_outputs[4256]);
    assign layer2_outputs[4191] = ~(layer1_outputs[995]);
    assign layer2_outputs[4192] = (layer1_outputs[1636]) & ~(layer1_outputs[4584]);
    assign layer2_outputs[4193] = ~(layer1_outputs[3094]);
    assign layer2_outputs[4194] = 1'b1;
    assign layer2_outputs[4195] = (layer1_outputs[4113]) & (layer1_outputs[4383]);
    assign layer2_outputs[4196] = (layer1_outputs[3216]) & ~(layer1_outputs[2580]);
    assign layer2_outputs[4197] = (layer1_outputs[3317]) & (layer1_outputs[164]);
    assign layer2_outputs[4198] = 1'b0;
    assign layer2_outputs[4199] = ~(layer1_outputs[2512]);
    assign layer2_outputs[4200] = (layer1_outputs[2002]) & (layer1_outputs[4035]);
    assign layer2_outputs[4201] = ~(layer1_outputs[709]) | (layer1_outputs[3207]);
    assign layer2_outputs[4202] = (layer1_outputs[2653]) & ~(layer1_outputs[3345]);
    assign layer2_outputs[4203] = 1'b1;
    assign layer2_outputs[4204] = ~(layer1_outputs[2280]);
    assign layer2_outputs[4205] = ~(layer1_outputs[448]);
    assign layer2_outputs[4206] = ~(layer1_outputs[3834]) | (layer1_outputs[2526]);
    assign layer2_outputs[4207] = 1'b0;
    assign layer2_outputs[4208] = (layer1_outputs[1563]) | (layer1_outputs[2270]);
    assign layer2_outputs[4209] = ~((layer1_outputs[3249]) & (layer1_outputs[4170]));
    assign layer2_outputs[4210] = (layer1_outputs[4771]) & ~(layer1_outputs[1444]);
    assign layer2_outputs[4211] = layer1_outputs[2620];
    assign layer2_outputs[4212] = ~((layer1_outputs[4945]) & (layer1_outputs[4614]));
    assign layer2_outputs[4213] = ~(layer1_outputs[912]);
    assign layer2_outputs[4214] = (layer1_outputs[3970]) & ~(layer1_outputs[2245]);
    assign layer2_outputs[4215] = (layer1_outputs[1365]) & ~(layer1_outputs[4034]);
    assign layer2_outputs[4216] = ~(layer1_outputs[1458]);
    assign layer2_outputs[4217] = ~(layer1_outputs[861]);
    assign layer2_outputs[4218] = 1'b1;
    assign layer2_outputs[4219] = 1'b1;
    assign layer2_outputs[4220] = ~((layer1_outputs[1431]) & (layer1_outputs[3886]));
    assign layer2_outputs[4221] = (layer1_outputs[2975]) | (layer1_outputs[2163]);
    assign layer2_outputs[4222] = layer1_outputs[3411];
    assign layer2_outputs[4223] = (layer1_outputs[3635]) ^ (layer1_outputs[688]);
    assign layer2_outputs[4224] = (layer1_outputs[4042]) & ~(layer1_outputs[1787]);
    assign layer2_outputs[4225] = 1'b0;
    assign layer2_outputs[4226] = (layer1_outputs[4035]) | (layer1_outputs[4013]);
    assign layer2_outputs[4227] = ~(layer1_outputs[700]);
    assign layer2_outputs[4228] = layer1_outputs[2201];
    assign layer2_outputs[4229] = layer1_outputs[4545];
    assign layer2_outputs[4230] = 1'b0;
    assign layer2_outputs[4231] = layer1_outputs[4328];
    assign layer2_outputs[4232] = 1'b1;
    assign layer2_outputs[4233] = 1'b0;
    assign layer2_outputs[4234] = (layer1_outputs[735]) & (layer1_outputs[4559]);
    assign layer2_outputs[4235] = (layer1_outputs[2396]) & (layer1_outputs[5094]);
    assign layer2_outputs[4236] = ~(layer1_outputs[3750]);
    assign layer2_outputs[4237] = 1'b0;
    assign layer2_outputs[4238] = ~((layer1_outputs[3423]) & (layer1_outputs[1846]));
    assign layer2_outputs[4239] = 1'b1;
    assign layer2_outputs[4240] = layer1_outputs[4760];
    assign layer2_outputs[4241] = layer1_outputs[1830];
    assign layer2_outputs[4242] = ~(layer1_outputs[1599]);
    assign layer2_outputs[4243] = ~((layer1_outputs[3436]) | (layer1_outputs[2926]));
    assign layer2_outputs[4244] = ~((layer1_outputs[4567]) & (layer1_outputs[2741]));
    assign layer2_outputs[4245] = 1'b0;
    assign layer2_outputs[4246] = layer1_outputs[4504];
    assign layer2_outputs[4247] = (layer1_outputs[1395]) & ~(layer1_outputs[2866]);
    assign layer2_outputs[4248] = (layer1_outputs[4388]) | (layer1_outputs[664]);
    assign layer2_outputs[4249] = (layer1_outputs[1859]) | (layer1_outputs[4176]);
    assign layer2_outputs[4250] = (layer1_outputs[2733]) & ~(layer1_outputs[131]);
    assign layer2_outputs[4251] = (layer1_outputs[561]) & ~(layer1_outputs[7]);
    assign layer2_outputs[4252] = (layer1_outputs[4840]) & ~(layer1_outputs[1983]);
    assign layer2_outputs[4253] = ~((layer1_outputs[2987]) | (layer1_outputs[3475]));
    assign layer2_outputs[4254] = (layer1_outputs[4378]) | (layer1_outputs[3612]);
    assign layer2_outputs[4255] = ~(layer1_outputs[2985]);
    assign layer2_outputs[4256] = ~((layer1_outputs[534]) ^ (layer1_outputs[580]));
    assign layer2_outputs[4257] = 1'b0;
    assign layer2_outputs[4258] = (layer1_outputs[4203]) & ~(layer1_outputs[4753]);
    assign layer2_outputs[4259] = (layer1_outputs[1425]) & ~(layer1_outputs[4505]);
    assign layer2_outputs[4260] = 1'b0;
    assign layer2_outputs[4261] = layer1_outputs[336];
    assign layer2_outputs[4262] = layer1_outputs[1737];
    assign layer2_outputs[4263] = (layer1_outputs[1654]) | (layer1_outputs[1075]);
    assign layer2_outputs[4264] = 1'b1;
    assign layer2_outputs[4265] = layer1_outputs[2498];
    assign layer2_outputs[4266] = 1'b1;
    assign layer2_outputs[4267] = ~(layer1_outputs[3813]);
    assign layer2_outputs[4268] = ~(layer1_outputs[2068]) | (layer1_outputs[577]);
    assign layer2_outputs[4269] = 1'b0;
    assign layer2_outputs[4270] = layer1_outputs[2564];
    assign layer2_outputs[4271] = layer1_outputs[2080];
    assign layer2_outputs[4272] = layer1_outputs[3976];
    assign layer2_outputs[4273] = ~((layer1_outputs[341]) ^ (layer1_outputs[299]));
    assign layer2_outputs[4274] = ~(layer1_outputs[4029]);
    assign layer2_outputs[4275] = ~(layer1_outputs[323]);
    assign layer2_outputs[4276] = ~(layer1_outputs[1108]);
    assign layer2_outputs[4277] = (layer1_outputs[1724]) & ~(layer1_outputs[2049]);
    assign layer2_outputs[4278] = 1'b0;
    assign layer2_outputs[4279] = ~((layer1_outputs[3843]) | (layer1_outputs[1434]));
    assign layer2_outputs[4280] = layer1_outputs[1813];
    assign layer2_outputs[4281] = ~(layer1_outputs[1052]);
    assign layer2_outputs[4282] = (layer1_outputs[1624]) | (layer1_outputs[4803]);
    assign layer2_outputs[4283] = ~(layer1_outputs[4518]);
    assign layer2_outputs[4284] = (layer1_outputs[2691]) | (layer1_outputs[5116]);
    assign layer2_outputs[4285] = (layer1_outputs[2953]) & ~(layer1_outputs[4087]);
    assign layer2_outputs[4286] = (layer1_outputs[3685]) & ~(layer1_outputs[4719]);
    assign layer2_outputs[4287] = ~(layer1_outputs[472]) | (layer1_outputs[2687]);
    assign layer2_outputs[4288] = 1'b1;
    assign layer2_outputs[4289] = (layer1_outputs[3684]) & ~(layer1_outputs[1834]);
    assign layer2_outputs[4290] = ~(layer1_outputs[136]) | (layer1_outputs[4041]);
    assign layer2_outputs[4291] = layer1_outputs[3407];
    assign layer2_outputs[4292] = ~((layer1_outputs[2168]) & (layer1_outputs[925]));
    assign layer2_outputs[4293] = ~(layer1_outputs[3046]);
    assign layer2_outputs[4294] = (layer1_outputs[3510]) ^ (layer1_outputs[3245]);
    assign layer2_outputs[4295] = ~(layer1_outputs[4528]) | (layer1_outputs[2890]);
    assign layer2_outputs[4296] = layer1_outputs[4285];
    assign layer2_outputs[4297] = ~((layer1_outputs[2548]) & (layer1_outputs[2949]));
    assign layer2_outputs[4298] = 1'b1;
    assign layer2_outputs[4299] = ~((layer1_outputs[561]) & (layer1_outputs[5023]));
    assign layer2_outputs[4300] = (layer1_outputs[3263]) & ~(layer1_outputs[4125]);
    assign layer2_outputs[4301] = ~(layer1_outputs[1965]) | (layer1_outputs[2888]);
    assign layer2_outputs[4302] = 1'b1;
    assign layer2_outputs[4303] = 1'b1;
    assign layer2_outputs[4304] = layer1_outputs[806];
    assign layer2_outputs[4305] = (layer1_outputs[1918]) & ~(layer1_outputs[2127]);
    assign layer2_outputs[4306] = (layer1_outputs[4169]) & ~(layer1_outputs[3950]);
    assign layer2_outputs[4307] = layer1_outputs[1466];
    assign layer2_outputs[4308] = (layer1_outputs[4624]) & ~(layer1_outputs[3827]);
    assign layer2_outputs[4309] = layer1_outputs[1582];
    assign layer2_outputs[4310] = layer1_outputs[2607];
    assign layer2_outputs[4311] = ~(layer1_outputs[2817]);
    assign layer2_outputs[4312] = (layer1_outputs[5024]) | (layer1_outputs[567]);
    assign layer2_outputs[4313] = layer1_outputs[1061];
    assign layer2_outputs[4314] = ~((layer1_outputs[3427]) ^ (layer1_outputs[4506]));
    assign layer2_outputs[4315] = 1'b0;
    assign layer2_outputs[4316] = (layer1_outputs[2232]) ^ (layer1_outputs[4330]);
    assign layer2_outputs[4317] = ~((layer1_outputs[179]) | (layer1_outputs[2932]));
    assign layer2_outputs[4318] = layer1_outputs[2146];
    assign layer2_outputs[4319] = ~((layer1_outputs[3132]) & (layer1_outputs[4558]));
    assign layer2_outputs[4320] = (layer1_outputs[1635]) & (layer1_outputs[493]);
    assign layer2_outputs[4321] = (layer1_outputs[4140]) & (layer1_outputs[2844]);
    assign layer2_outputs[4322] = (layer1_outputs[1703]) & ~(layer1_outputs[4207]);
    assign layer2_outputs[4323] = 1'b0;
    assign layer2_outputs[4324] = 1'b0;
    assign layer2_outputs[4325] = ~((layer1_outputs[293]) ^ (layer1_outputs[4009]));
    assign layer2_outputs[4326] = (layer1_outputs[2516]) ^ (layer1_outputs[3954]);
    assign layer2_outputs[4327] = layer1_outputs[3082];
    assign layer2_outputs[4328] = (layer1_outputs[2281]) | (layer1_outputs[3314]);
    assign layer2_outputs[4329] = ~(layer1_outputs[471]);
    assign layer2_outputs[4330] = ~((layer1_outputs[3714]) | (layer1_outputs[2381]));
    assign layer2_outputs[4331] = (layer1_outputs[2256]) | (layer1_outputs[3675]);
    assign layer2_outputs[4332] = layer1_outputs[635];
    assign layer2_outputs[4333] = ~((layer1_outputs[446]) & (layer1_outputs[2165]));
    assign layer2_outputs[4334] = layer1_outputs[2221];
    assign layer2_outputs[4335] = (layer1_outputs[4812]) & ~(layer1_outputs[3692]);
    assign layer2_outputs[4336] = ~(layer1_outputs[412]);
    assign layer2_outputs[4337] = (layer1_outputs[3480]) & ~(layer1_outputs[2010]);
    assign layer2_outputs[4338] = 1'b0;
    assign layer2_outputs[4339] = 1'b1;
    assign layer2_outputs[4340] = ~(layer1_outputs[272]) | (layer1_outputs[4166]);
    assign layer2_outputs[4341] = ~((layer1_outputs[3858]) | (layer1_outputs[1768]));
    assign layer2_outputs[4342] = 1'b1;
    assign layer2_outputs[4343] = layer1_outputs[4387];
    assign layer2_outputs[4344] = ~(layer1_outputs[552]) | (layer1_outputs[2819]);
    assign layer2_outputs[4345] = (layer1_outputs[809]) & (layer1_outputs[2490]);
    assign layer2_outputs[4346] = 1'b0;
    assign layer2_outputs[4347] = 1'b0;
    assign layer2_outputs[4348] = layer1_outputs[87];
    assign layer2_outputs[4349] = 1'b0;
    assign layer2_outputs[4350] = ~(layer1_outputs[4887]);
    assign layer2_outputs[4351] = ~(layer1_outputs[1810]);
    assign layer2_outputs[4352] = (layer1_outputs[2568]) | (layer1_outputs[4871]);
    assign layer2_outputs[4353] = (layer1_outputs[1929]) | (layer1_outputs[4910]);
    assign layer2_outputs[4354] = (layer1_outputs[3785]) & ~(layer1_outputs[3951]);
    assign layer2_outputs[4355] = (layer1_outputs[3298]) & ~(layer1_outputs[4420]);
    assign layer2_outputs[4356] = layer1_outputs[4646];
    assign layer2_outputs[4357] = ~(layer1_outputs[3381]);
    assign layer2_outputs[4358] = layer1_outputs[2158];
    assign layer2_outputs[4359] = ~(layer1_outputs[2891]);
    assign layer2_outputs[4360] = ~(layer1_outputs[1660]);
    assign layer2_outputs[4361] = layer1_outputs[759];
    assign layer2_outputs[4362] = 1'b0;
    assign layer2_outputs[4363] = 1'b0;
    assign layer2_outputs[4364] = ~(layer1_outputs[3724]) | (layer1_outputs[3388]);
    assign layer2_outputs[4365] = ~(layer1_outputs[3654]);
    assign layer2_outputs[4366] = 1'b0;
    assign layer2_outputs[4367] = layer1_outputs[201];
    assign layer2_outputs[4368] = layer1_outputs[4000];
    assign layer2_outputs[4369] = ~(layer1_outputs[733]);
    assign layer2_outputs[4370] = 1'b1;
    assign layer2_outputs[4371] = layer1_outputs[787];
    assign layer2_outputs[4372] = (layer1_outputs[2530]) & ~(layer1_outputs[4999]);
    assign layer2_outputs[4373] = ~(layer1_outputs[2032]) | (layer1_outputs[2293]);
    assign layer2_outputs[4374] = ~(layer1_outputs[94]) | (layer1_outputs[3066]);
    assign layer2_outputs[4375] = layer1_outputs[637];
    assign layer2_outputs[4376] = layer1_outputs[1122];
    assign layer2_outputs[4377] = ~(layer1_outputs[1540]);
    assign layer2_outputs[4378] = (layer1_outputs[819]) | (layer1_outputs[1650]);
    assign layer2_outputs[4379] = (layer1_outputs[3873]) | (layer1_outputs[1343]);
    assign layer2_outputs[4380] = (layer1_outputs[1454]) | (layer1_outputs[4547]);
    assign layer2_outputs[4381] = ~((layer1_outputs[2327]) | (layer1_outputs[3071]));
    assign layer2_outputs[4382] = layer1_outputs[4848];
    assign layer2_outputs[4383] = layer1_outputs[1949];
    assign layer2_outputs[4384] = ~((layer1_outputs[3826]) | (layer1_outputs[658]));
    assign layer2_outputs[4385] = ~((layer1_outputs[1870]) & (layer1_outputs[2955]));
    assign layer2_outputs[4386] = 1'b1;
    assign layer2_outputs[4387] = 1'b0;
    assign layer2_outputs[4388] = ~((layer1_outputs[4601]) & (layer1_outputs[3608]));
    assign layer2_outputs[4389] = ~(layer1_outputs[3919]) | (layer1_outputs[2585]);
    assign layer2_outputs[4390] = ~(layer1_outputs[3570]);
    assign layer2_outputs[4391] = ~((layer1_outputs[2662]) | (layer1_outputs[4311]));
    assign layer2_outputs[4392] = ~(layer1_outputs[1556]) | (layer1_outputs[4212]);
    assign layer2_outputs[4393] = 1'b1;
    assign layer2_outputs[4394] = ~((layer1_outputs[2337]) | (layer1_outputs[2516]));
    assign layer2_outputs[4395] = 1'b1;
    assign layer2_outputs[4396] = 1'b1;
    assign layer2_outputs[4397] = ~((layer1_outputs[3958]) | (layer1_outputs[4449]));
    assign layer2_outputs[4398] = ~((layer1_outputs[3691]) & (layer1_outputs[1965]));
    assign layer2_outputs[4399] = ~(layer1_outputs[971]);
    assign layer2_outputs[4400] = (layer1_outputs[3327]) | (layer1_outputs[1362]);
    assign layer2_outputs[4401] = layer1_outputs[1008];
    assign layer2_outputs[4402] = (layer1_outputs[1354]) & ~(layer1_outputs[3036]);
    assign layer2_outputs[4403] = 1'b1;
    assign layer2_outputs[4404] = layer1_outputs[2567];
    assign layer2_outputs[4405] = ~((layer1_outputs[292]) | (layer1_outputs[4537]));
    assign layer2_outputs[4406] = 1'b0;
    assign layer2_outputs[4407] = (layer1_outputs[2686]) | (layer1_outputs[3237]);
    assign layer2_outputs[4408] = (layer1_outputs[1991]) & ~(layer1_outputs[892]);
    assign layer2_outputs[4409] = layer1_outputs[746];
    assign layer2_outputs[4410] = layer1_outputs[1822];
    assign layer2_outputs[4411] = layer1_outputs[5019];
    assign layer2_outputs[4412] = (layer1_outputs[2992]) & (layer1_outputs[4124]);
    assign layer2_outputs[4413] = 1'b0;
    assign layer2_outputs[4414] = ~((layer1_outputs[1173]) | (layer1_outputs[131]));
    assign layer2_outputs[4415] = ~((layer1_outputs[2532]) | (layer1_outputs[4598]));
    assign layer2_outputs[4416] = 1'b1;
    assign layer2_outputs[4417] = ~((layer1_outputs[1780]) | (layer1_outputs[3561]));
    assign layer2_outputs[4418] = ~((layer1_outputs[1375]) ^ (layer1_outputs[2196]));
    assign layer2_outputs[4419] = ~(layer1_outputs[710]);
    assign layer2_outputs[4420] = 1'b0;
    assign layer2_outputs[4421] = 1'b0;
    assign layer2_outputs[4422] = ~(layer1_outputs[387]);
    assign layer2_outputs[4423] = ~(layer1_outputs[1154]);
    assign layer2_outputs[4424] = 1'b1;
    assign layer2_outputs[4425] = layer1_outputs[3062];
    assign layer2_outputs[4426] = layer1_outputs[2761];
    assign layer2_outputs[4427] = ~(layer1_outputs[1361]) | (layer1_outputs[2632]);
    assign layer2_outputs[4428] = (layer1_outputs[4670]) | (layer1_outputs[4863]);
    assign layer2_outputs[4429] = (layer1_outputs[1862]) | (layer1_outputs[834]);
    assign layer2_outputs[4430] = (layer1_outputs[3380]) & (layer1_outputs[1401]);
    assign layer2_outputs[4431] = layer1_outputs[1989];
    assign layer2_outputs[4432] = (layer1_outputs[587]) & ~(layer1_outputs[2705]);
    assign layer2_outputs[4433] = ~((layer1_outputs[4382]) | (layer1_outputs[5090]));
    assign layer2_outputs[4434] = ~((layer1_outputs[4146]) ^ (layer1_outputs[3783]));
    assign layer2_outputs[4435] = (layer1_outputs[1280]) & ~(layer1_outputs[3967]);
    assign layer2_outputs[4436] = (layer1_outputs[2358]) & (layer1_outputs[5029]);
    assign layer2_outputs[4437] = layer1_outputs[3203];
    assign layer2_outputs[4438] = ~(layer1_outputs[4500]);
    assign layer2_outputs[4439] = ~(layer1_outputs[4439]);
    assign layer2_outputs[4440] = 1'b0;
    assign layer2_outputs[4441] = (layer1_outputs[4771]) & ~(layer1_outputs[97]);
    assign layer2_outputs[4442] = ~(layer1_outputs[2085]) | (layer1_outputs[336]);
    assign layer2_outputs[4443] = layer1_outputs[887];
    assign layer2_outputs[4444] = 1'b0;
    assign layer2_outputs[4445] = ~((layer1_outputs[3828]) & (layer1_outputs[3176]));
    assign layer2_outputs[4446] = ~(layer1_outputs[63]) | (layer1_outputs[2666]);
    assign layer2_outputs[4447] = ~(layer1_outputs[4693]);
    assign layer2_outputs[4448] = layer1_outputs[2783];
    assign layer2_outputs[4449] = 1'b1;
    assign layer2_outputs[4450] = (layer1_outputs[4163]) & (layer1_outputs[642]);
    assign layer2_outputs[4451] = (layer1_outputs[3322]) | (layer1_outputs[3991]);
    assign layer2_outputs[4452] = (layer1_outputs[265]) & ~(layer1_outputs[3912]);
    assign layer2_outputs[4453] = ~(layer1_outputs[3148]);
    assign layer2_outputs[4454] = ~((layer1_outputs[2460]) | (layer1_outputs[1141]));
    assign layer2_outputs[4455] = (layer1_outputs[1829]) & ~(layer1_outputs[1659]);
    assign layer2_outputs[4456] = ~(layer1_outputs[4149]);
    assign layer2_outputs[4457] = ~(layer1_outputs[1217]);
    assign layer2_outputs[4458] = (layer1_outputs[2763]) & ~(layer1_outputs[790]);
    assign layer2_outputs[4459] = layer1_outputs[2977];
    assign layer2_outputs[4460] = (layer1_outputs[5063]) | (layer1_outputs[868]);
    assign layer2_outputs[4461] = (layer1_outputs[3768]) ^ (layer1_outputs[3844]);
    assign layer2_outputs[4462] = (layer1_outputs[1986]) & ~(layer1_outputs[175]);
    assign layer2_outputs[4463] = ~(layer1_outputs[2185]);
    assign layer2_outputs[4464] = ~((layer1_outputs[2807]) | (layer1_outputs[109]));
    assign layer2_outputs[4465] = ~((layer1_outputs[2165]) & (layer1_outputs[147]));
    assign layer2_outputs[4466] = layer1_outputs[1900];
    assign layer2_outputs[4467] = (layer1_outputs[392]) & ~(layer1_outputs[1987]);
    assign layer2_outputs[4468] = layer1_outputs[3669];
    assign layer2_outputs[4469] = ~(layer1_outputs[321]);
    assign layer2_outputs[4470] = 1'b0;
    assign layer2_outputs[4471] = ~(layer1_outputs[1439]) | (layer1_outputs[3102]);
    assign layer2_outputs[4472] = ~(layer1_outputs[1682]);
    assign layer2_outputs[4473] = ~(layer1_outputs[4147]);
    assign layer2_outputs[4474] = ~(layer1_outputs[2668]) | (layer1_outputs[3339]);
    assign layer2_outputs[4475] = ~((layer1_outputs[1025]) & (layer1_outputs[3148]));
    assign layer2_outputs[4476] = layer1_outputs[3301];
    assign layer2_outputs[4477] = (layer1_outputs[4259]) & ~(layer1_outputs[4457]);
    assign layer2_outputs[4478] = (layer1_outputs[3215]) & ~(layer1_outputs[1358]);
    assign layer2_outputs[4479] = layer1_outputs[1517];
    assign layer2_outputs[4480] = layer1_outputs[646];
    assign layer2_outputs[4481] = ~(layer1_outputs[844]);
    assign layer2_outputs[4482] = ~(layer1_outputs[1443]);
    assign layer2_outputs[4483] = ~((layer1_outputs[2379]) | (layer1_outputs[3674]));
    assign layer2_outputs[4484] = (layer1_outputs[484]) | (layer1_outputs[5102]);
    assign layer2_outputs[4485] = 1'b0;
    assign layer2_outputs[4486] = layer1_outputs[4310];
    assign layer2_outputs[4487] = 1'b0;
    assign layer2_outputs[4488] = layer1_outputs[4666];
    assign layer2_outputs[4489] = 1'b0;
    assign layer2_outputs[4490] = ~(layer1_outputs[2018]);
    assign layer2_outputs[4491] = layer1_outputs[428];
    assign layer2_outputs[4492] = ~((layer1_outputs[2367]) & (layer1_outputs[1439]));
    assign layer2_outputs[4493] = (layer1_outputs[1280]) ^ (layer1_outputs[3237]);
    assign layer2_outputs[4494] = (layer1_outputs[2518]) & ~(layer1_outputs[1407]);
    assign layer2_outputs[4495] = layer1_outputs[36];
    assign layer2_outputs[4496] = (layer1_outputs[1055]) & ~(layer1_outputs[4224]);
    assign layer2_outputs[4497] = ~((layer1_outputs[2994]) & (layer1_outputs[3597]));
    assign layer2_outputs[4498] = (layer1_outputs[2606]) & ~(layer1_outputs[2995]);
    assign layer2_outputs[4499] = layer1_outputs[2092];
    assign layer2_outputs[4500] = 1'b0;
    assign layer2_outputs[4501] = 1'b0;
    assign layer2_outputs[4502] = layer1_outputs[3548];
    assign layer2_outputs[4503] = ~((layer1_outputs[3870]) & (layer1_outputs[1567]));
    assign layer2_outputs[4504] = 1'b0;
    assign layer2_outputs[4505] = (layer1_outputs[4613]) & ~(layer1_outputs[22]);
    assign layer2_outputs[4506] = ~((layer1_outputs[326]) & (layer1_outputs[879]));
    assign layer2_outputs[4507] = 1'b1;
    assign layer2_outputs[4508] = ~(layer1_outputs[1595]);
    assign layer2_outputs[4509] = layer1_outputs[2537];
    assign layer2_outputs[4510] = ~((layer1_outputs[1921]) ^ (layer1_outputs[1875]));
    assign layer2_outputs[4511] = ~((layer1_outputs[3812]) | (layer1_outputs[2777]));
    assign layer2_outputs[4512] = (layer1_outputs[106]) & (layer1_outputs[784]);
    assign layer2_outputs[4513] = (layer1_outputs[3417]) | (layer1_outputs[2891]);
    assign layer2_outputs[4514] = layer1_outputs[2303];
    assign layer2_outputs[4515] = layer1_outputs[1400];
    assign layer2_outputs[4516] = ~(layer1_outputs[3196]) | (layer1_outputs[2589]);
    assign layer2_outputs[4517] = ~((layer1_outputs[3967]) | (layer1_outputs[2229]));
    assign layer2_outputs[4518] = ~(layer1_outputs[4385]) | (layer1_outputs[2237]);
    assign layer2_outputs[4519] = 1'b0;
    assign layer2_outputs[4520] = ~((layer1_outputs[2023]) | (layer1_outputs[883]));
    assign layer2_outputs[4521] = 1'b1;
    assign layer2_outputs[4522] = (layer1_outputs[1457]) | (layer1_outputs[4296]);
    assign layer2_outputs[4523] = (layer1_outputs[255]) & (layer1_outputs[4093]);
    assign layer2_outputs[4524] = ~(layer1_outputs[3924]);
    assign layer2_outputs[4525] = (layer1_outputs[1099]) & ~(layer1_outputs[4154]);
    assign layer2_outputs[4526] = layer1_outputs[1767];
    assign layer2_outputs[4527] = 1'b1;
    assign layer2_outputs[4528] = (layer1_outputs[1828]) & ~(layer1_outputs[1551]);
    assign layer2_outputs[4529] = ~(layer1_outputs[4945]) | (layer1_outputs[4965]);
    assign layer2_outputs[4530] = layer1_outputs[4048];
    assign layer2_outputs[4531] = (layer1_outputs[4578]) & (layer1_outputs[123]);
    assign layer2_outputs[4532] = ~((layer1_outputs[985]) & (layer1_outputs[1572]));
    assign layer2_outputs[4533] = 1'b1;
    assign layer2_outputs[4534] = layer1_outputs[2368];
    assign layer2_outputs[4535] = ~((layer1_outputs[319]) | (layer1_outputs[1484]));
    assign layer2_outputs[4536] = ~((layer1_outputs[5072]) & (layer1_outputs[317]));
    assign layer2_outputs[4537] = ~(layer1_outputs[731]);
    assign layer2_outputs[4538] = ~(layer1_outputs[2324]);
    assign layer2_outputs[4539] = ~(layer1_outputs[604]);
    assign layer2_outputs[4540] = ~(layer1_outputs[3440]);
    assign layer2_outputs[4541] = ~((layer1_outputs[1922]) | (layer1_outputs[4653]));
    assign layer2_outputs[4542] = (layer1_outputs[3003]) & ~(layer1_outputs[741]);
    assign layer2_outputs[4543] = 1'b0;
    assign layer2_outputs[4544] = layer1_outputs[3269];
    assign layer2_outputs[4545] = (layer1_outputs[3310]) & ~(layer1_outputs[3477]);
    assign layer2_outputs[4546] = (layer1_outputs[2812]) & (layer1_outputs[2513]);
    assign layer2_outputs[4547] = (layer1_outputs[1342]) & ~(layer1_outputs[4652]);
    assign layer2_outputs[4548] = layer1_outputs[2682];
    assign layer2_outputs[4549] = (layer1_outputs[1218]) | (layer1_outputs[1930]);
    assign layer2_outputs[4550] = 1'b1;
    assign layer2_outputs[4551] = 1'b0;
    assign layer2_outputs[4552] = ~((layer1_outputs[4542]) | (layer1_outputs[3925]));
    assign layer2_outputs[4553] = ~(layer1_outputs[2439]) | (layer1_outputs[3256]);
    assign layer2_outputs[4554] = ~(layer1_outputs[1126]) | (layer1_outputs[4750]);
    assign layer2_outputs[4555] = ~(layer1_outputs[1607]) | (layer1_outputs[3080]);
    assign layer2_outputs[4556] = ~(layer1_outputs[1122]) | (layer1_outputs[1188]);
    assign layer2_outputs[4557] = ~((layer1_outputs[4040]) & (layer1_outputs[2441]));
    assign layer2_outputs[4558] = ~((layer1_outputs[339]) & (layer1_outputs[1372]));
    assign layer2_outputs[4559] = ~(layer1_outputs[1371]) | (layer1_outputs[3163]);
    assign layer2_outputs[4560] = layer1_outputs[4320];
    assign layer2_outputs[4561] = layer1_outputs[2894];
    assign layer2_outputs[4562] = (layer1_outputs[4750]) & (layer1_outputs[2911]);
    assign layer2_outputs[4563] = 1'b0;
    assign layer2_outputs[4564] = (layer1_outputs[3515]) & ~(layer1_outputs[3089]);
    assign layer2_outputs[4565] = ~(layer1_outputs[410]);
    assign layer2_outputs[4566] = 1'b1;
    assign layer2_outputs[4567] = (layer1_outputs[1573]) & ~(layer1_outputs[2620]);
    assign layer2_outputs[4568] = ~(layer1_outputs[4775]) | (layer1_outputs[4882]);
    assign layer2_outputs[4569] = (layer1_outputs[947]) & ~(layer1_outputs[4252]);
    assign layer2_outputs[4570] = (layer1_outputs[573]) & ~(layer1_outputs[2810]);
    assign layer2_outputs[4571] = (layer1_outputs[3916]) ^ (layer1_outputs[1048]);
    assign layer2_outputs[4572] = layer1_outputs[212];
    assign layer2_outputs[4573] = ~((layer1_outputs[3726]) | (layer1_outputs[2105]));
    assign layer2_outputs[4574] = layer1_outputs[1183];
    assign layer2_outputs[4575] = ~(layer1_outputs[3875]);
    assign layer2_outputs[4576] = 1'b0;
    assign layer2_outputs[4577] = 1'b1;
    assign layer2_outputs[4578] = ~(layer1_outputs[2310]) | (layer1_outputs[1013]);
    assign layer2_outputs[4579] = layer1_outputs[3943];
    assign layer2_outputs[4580] = ~((layer1_outputs[2819]) | (layer1_outputs[449]));
    assign layer2_outputs[4581] = (layer1_outputs[3594]) | (layer1_outputs[240]);
    assign layer2_outputs[4582] = ~(layer1_outputs[69]) | (layer1_outputs[3367]);
    assign layer2_outputs[4583] = (layer1_outputs[3985]) ^ (layer1_outputs[2669]);
    assign layer2_outputs[4584] = (layer1_outputs[3637]) | (layer1_outputs[334]);
    assign layer2_outputs[4585] = ~(layer1_outputs[269]);
    assign layer2_outputs[4586] = ~(layer1_outputs[1997]) | (layer1_outputs[1860]);
    assign layer2_outputs[4587] = 1'b1;
    assign layer2_outputs[4588] = 1'b1;
    assign layer2_outputs[4589] = (layer1_outputs[2187]) ^ (layer1_outputs[4196]);
    assign layer2_outputs[4590] = ~(layer1_outputs[1138]) | (layer1_outputs[3085]);
    assign layer2_outputs[4591] = ~(layer1_outputs[1089]) | (layer1_outputs[2060]);
    assign layer2_outputs[4592] = 1'b0;
    assign layer2_outputs[4593] = layer1_outputs[2360];
    assign layer2_outputs[4594] = ~((layer1_outputs[3672]) | (layer1_outputs[2366]));
    assign layer2_outputs[4595] = ~(layer1_outputs[467]);
    assign layer2_outputs[4596] = layer1_outputs[5058];
    assign layer2_outputs[4597] = ~((layer1_outputs[1469]) & (layer1_outputs[4832]));
    assign layer2_outputs[4598] = layer1_outputs[536];
    assign layer2_outputs[4599] = ~(layer1_outputs[2683]) | (layer1_outputs[1081]);
    assign layer2_outputs[4600] = layer1_outputs[3564];
    assign layer2_outputs[4601] = ~((layer1_outputs[3775]) | (layer1_outputs[699]));
    assign layer2_outputs[4602] = 1'b1;
    assign layer2_outputs[4603] = ~((layer1_outputs[1428]) | (layer1_outputs[12]));
    assign layer2_outputs[4604] = (layer1_outputs[582]) | (layer1_outputs[182]);
    assign layer2_outputs[4605] = ~(layer1_outputs[1758]) | (layer1_outputs[3149]);
    assign layer2_outputs[4606] = (layer1_outputs[1709]) | (layer1_outputs[525]);
    assign layer2_outputs[4607] = ~(layer1_outputs[2605]) | (layer1_outputs[5055]);
    assign layer2_outputs[4608] = ~(layer1_outputs[1295]);
    assign layer2_outputs[4609] = 1'b1;
    assign layer2_outputs[4610] = (layer1_outputs[4574]) & ~(layer1_outputs[1244]);
    assign layer2_outputs[4611] = ~(layer1_outputs[547]);
    assign layer2_outputs[4612] = layer1_outputs[1647];
    assign layer2_outputs[4613] = ~(layer1_outputs[831]);
    assign layer2_outputs[4614] = (layer1_outputs[1330]) & ~(layer1_outputs[2026]);
    assign layer2_outputs[4615] = ~(layer1_outputs[4443]) | (layer1_outputs[601]);
    assign layer2_outputs[4616] = ~(layer1_outputs[4320]);
    assign layer2_outputs[4617] = ~((layer1_outputs[775]) ^ (layer1_outputs[5066]));
    assign layer2_outputs[4618] = (layer1_outputs[2360]) & (layer1_outputs[2734]);
    assign layer2_outputs[4619] = ~((layer1_outputs[2091]) ^ (layer1_outputs[4942]));
    assign layer2_outputs[4620] = (layer1_outputs[3678]) & (layer1_outputs[493]);
    assign layer2_outputs[4621] = 1'b1;
    assign layer2_outputs[4622] = layer1_outputs[2099];
    assign layer2_outputs[4623] = (layer1_outputs[3085]) & (layer1_outputs[3508]);
    assign layer2_outputs[4624] = (layer1_outputs[4187]) ^ (layer1_outputs[3439]);
    assign layer2_outputs[4625] = ~(layer1_outputs[4888]) | (layer1_outputs[4715]);
    assign layer2_outputs[4626] = ~((layer1_outputs[4273]) | (layer1_outputs[4780]));
    assign layer2_outputs[4627] = ~(layer1_outputs[4432]);
    assign layer2_outputs[4628] = (layer1_outputs[1733]) & (layer1_outputs[121]);
    assign layer2_outputs[4629] = (layer1_outputs[981]) & (layer1_outputs[852]);
    assign layer2_outputs[4630] = ~(layer1_outputs[177]) | (layer1_outputs[920]);
    assign layer2_outputs[4631] = (layer1_outputs[798]) & ~(layer1_outputs[3796]);
    assign layer2_outputs[4632] = ~((layer1_outputs[3415]) ^ (layer1_outputs[1747]));
    assign layer2_outputs[4633] = layer1_outputs[4263];
    assign layer2_outputs[4634] = ~(layer1_outputs[4964]);
    assign layer2_outputs[4635] = ~((layer1_outputs[2791]) & (layer1_outputs[888]));
    assign layer2_outputs[4636] = ~(layer1_outputs[95]) | (layer1_outputs[302]);
    assign layer2_outputs[4637] = ~((layer1_outputs[2479]) | (layer1_outputs[2858]));
    assign layer2_outputs[4638] = (layer1_outputs[3535]) & ~(layer1_outputs[1733]);
    assign layer2_outputs[4639] = ~(layer1_outputs[4099]) | (layer1_outputs[2181]);
    assign layer2_outputs[4640] = ~(layer1_outputs[2461]) | (layer1_outputs[3344]);
    assign layer2_outputs[4641] = ~(layer1_outputs[4088]);
    assign layer2_outputs[4642] = layer1_outputs[1475];
    assign layer2_outputs[4643] = (layer1_outputs[3098]) & (layer1_outputs[2549]);
    assign layer2_outputs[4644] = ~((layer1_outputs[3681]) | (layer1_outputs[1044]));
    assign layer2_outputs[4645] = ~((layer1_outputs[4182]) & (layer1_outputs[5034]));
    assign layer2_outputs[4646] = layer1_outputs[3980];
    assign layer2_outputs[4647] = ~((layer1_outputs[2406]) & (layer1_outputs[136]));
    assign layer2_outputs[4648] = ~(layer1_outputs[2408]) | (layer1_outputs[2126]);
    assign layer2_outputs[4649] = ~(layer1_outputs[521]) | (layer1_outputs[1633]);
    assign layer2_outputs[4650] = (layer1_outputs[2885]) & (layer1_outputs[2007]);
    assign layer2_outputs[4651] = 1'b1;
    assign layer2_outputs[4652] = ~(layer1_outputs[3486]);
    assign layer2_outputs[4653] = ~((layer1_outputs[4767]) ^ (layer1_outputs[1450]));
    assign layer2_outputs[4654] = ~((layer1_outputs[118]) & (layer1_outputs[3059]));
    assign layer2_outputs[4655] = ~(layer1_outputs[3962]);
    assign layer2_outputs[4656] = layer1_outputs[911];
    assign layer2_outputs[4657] = layer1_outputs[4007];
    assign layer2_outputs[4658] = 1'b0;
    assign layer2_outputs[4659] = layer1_outputs[1104];
    assign layer2_outputs[4660] = 1'b1;
    assign layer2_outputs[4661] = 1'b1;
    assign layer2_outputs[4662] = 1'b1;
    assign layer2_outputs[4663] = 1'b1;
    assign layer2_outputs[4664] = (layer1_outputs[1262]) | (layer1_outputs[4946]);
    assign layer2_outputs[4665] = layer1_outputs[3150];
    assign layer2_outputs[4666] = layer1_outputs[4423];
    assign layer2_outputs[4667] = (layer1_outputs[3095]) & (layer1_outputs[607]);
    assign layer2_outputs[4668] = ~(layer1_outputs[2474]);
    assign layer2_outputs[4669] = ~((layer1_outputs[4130]) & (layer1_outputs[4583]));
    assign layer2_outputs[4670] = 1'b1;
    assign layer2_outputs[4671] = ~((layer1_outputs[4934]) & (layer1_outputs[4732]));
    assign layer2_outputs[4672] = (layer1_outputs[2838]) ^ (layer1_outputs[4146]);
    assign layer2_outputs[4673] = layer1_outputs[766];
    assign layer2_outputs[4674] = (layer1_outputs[846]) & (layer1_outputs[4]);
    assign layer2_outputs[4675] = ~(layer1_outputs[4089]) | (layer1_outputs[91]);
    assign layer2_outputs[4676] = (layer1_outputs[1771]) & ~(layer1_outputs[4541]);
    assign layer2_outputs[4677] = 1'b1;
    assign layer2_outputs[4678] = ~(layer1_outputs[4749]);
    assign layer2_outputs[4679] = layer1_outputs[1255];
    assign layer2_outputs[4680] = 1'b0;
    assign layer2_outputs[4681] = layer1_outputs[3769];
    assign layer2_outputs[4682] = ~(layer1_outputs[4792]) | (layer1_outputs[1775]);
    assign layer2_outputs[4683] = layer1_outputs[3548];
    assign layer2_outputs[4684] = layer1_outputs[2420];
    assign layer2_outputs[4685] = (layer1_outputs[2265]) ^ (layer1_outputs[2028]);
    assign layer2_outputs[4686] = ~(layer1_outputs[1528]);
    assign layer2_outputs[4687] = ~((layer1_outputs[4008]) | (layer1_outputs[3293]));
    assign layer2_outputs[4688] = (layer1_outputs[4200]) & ~(layer1_outputs[1527]);
    assign layer2_outputs[4689] = ~(layer1_outputs[3907]) | (layer1_outputs[1409]);
    assign layer2_outputs[4690] = (layer1_outputs[457]) & ~(layer1_outputs[3555]);
    assign layer2_outputs[4691] = 1'b0;
    assign layer2_outputs[4692] = (layer1_outputs[3234]) ^ (layer1_outputs[780]);
    assign layer2_outputs[4693] = ~(layer1_outputs[4960]);
    assign layer2_outputs[4694] = ~((layer1_outputs[2560]) | (layer1_outputs[4729]));
    assign layer2_outputs[4695] = 1'b1;
    assign layer2_outputs[4696] = (layer1_outputs[1735]) & (layer1_outputs[968]);
    assign layer2_outputs[4697] = ~(layer1_outputs[1860]);
    assign layer2_outputs[4698] = ~(layer1_outputs[4812]) | (layer1_outputs[3196]);
    assign layer2_outputs[4699] = (layer1_outputs[3368]) | (layer1_outputs[3404]);
    assign layer2_outputs[4700] = ~(layer1_outputs[1364]);
    assign layer2_outputs[4701] = ~((layer1_outputs[910]) & (layer1_outputs[2841]));
    assign layer2_outputs[4702] = ~(layer1_outputs[818]) | (layer1_outputs[781]);
    assign layer2_outputs[4703] = ~((layer1_outputs[4993]) | (layer1_outputs[4765]));
    assign layer2_outputs[4704] = ~(layer1_outputs[475]);
    assign layer2_outputs[4705] = ~((layer1_outputs[4615]) & (layer1_outputs[3435]));
    assign layer2_outputs[4706] = layer1_outputs[3877];
    assign layer2_outputs[4707] = ~(layer1_outputs[1378]);
    assign layer2_outputs[4708] = (layer1_outputs[1926]) & ~(layer1_outputs[4107]);
    assign layer2_outputs[4709] = 1'b0;
    assign layer2_outputs[4710] = layer1_outputs[931];
    assign layer2_outputs[4711] = 1'b1;
    assign layer2_outputs[4712] = (layer1_outputs[4833]) & (layer1_outputs[2001]);
    assign layer2_outputs[4713] = (layer1_outputs[4182]) & ~(layer1_outputs[1346]);
    assign layer2_outputs[4714] = layer1_outputs[1852];
    assign layer2_outputs[4715] = (layer1_outputs[4654]) & ~(layer1_outputs[4751]);
    assign layer2_outputs[4716] = 1'b0;
    assign layer2_outputs[4717] = (layer1_outputs[507]) | (layer1_outputs[3794]);
    assign layer2_outputs[4718] = ~(layer1_outputs[3629]) | (layer1_outputs[15]);
    assign layer2_outputs[4719] = ~(layer1_outputs[1752]) | (layer1_outputs[2573]);
    assign layer2_outputs[4720] = ~(layer1_outputs[629]) | (layer1_outputs[980]);
    assign layer2_outputs[4721] = layer1_outputs[1683];
    assign layer2_outputs[4722] = ~((layer1_outputs[622]) & (layer1_outputs[3505]));
    assign layer2_outputs[4723] = ~(layer1_outputs[4238]);
    assign layer2_outputs[4724] = ~((layer1_outputs[146]) & (layer1_outputs[4444]));
    assign layer2_outputs[4725] = (layer1_outputs[5005]) | (layer1_outputs[5048]);
    assign layer2_outputs[4726] = (layer1_outputs[4639]) & (layer1_outputs[5050]);
    assign layer2_outputs[4727] = layer1_outputs[3395];
    assign layer2_outputs[4728] = ~((layer1_outputs[2613]) & (layer1_outputs[4342]));
    assign layer2_outputs[4729] = (layer1_outputs[4684]) | (layer1_outputs[4303]);
    assign layer2_outputs[4730] = layer1_outputs[4856];
    assign layer2_outputs[4731] = 1'b0;
    assign layer2_outputs[4732] = ~(layer1_outputs[3890]) | (layer1_outputs[3274]);
    assign layer2_outputs[4733] = (layer1_outputs[1329]) & (layer1_outputs[310]);
    assign layer2_outputs[4734] = (layer1_outputs[440]) & ~(layer1_outputs[2451]);
    assign layer2_outputs[4735] = ~(layer1_outputs[4974]);
    assign layer2_outputs[4736] = ~(layer1_outputs[4775]);
    assign layer2_outputs[4737] = ~(layer1_outputs[1405]) | (layer1_outputs[4980]);
    assign layer2_outputs[4738] = (layer1_outputs[1316]) & ~(layer1_outputs[4847]);
    assign layer2_outputs[4739] = ~(layer1_outputs[4360]);
    assign layer2_outputs[4740] = layer1_outputs[3941];
    assign layer2_outputs[4741] = ~((layer1_outputs[230]) & (layer1_outputs[3917]));
    assign layer2_outputs[4742] = ~((layer1_outputs[5001]) | (layer1_outputs[900]));
    assign layer2_outputs[4743] = ~(layer1_outputs[246]);
    assign layer2_outputs[4744] = ~(layer1_outputs[2855]);
    assign layer2_outputs[4745] = ~(layer1_outputs[4262]) | (layer1_outputs[5040]);
    assign layer2_outputs[4746] = 1'b1;
    assign layer2_outputs[4747] = ~((layer1_outputs[4970]) ^ (layer1_outputs[3296]));
    assign layer2_outputs[4748] = ~(layer1_outputs[356]);
    assign layer2_outputs[4749] = ~(layer1_outputs[4656]);
    assign layer2_outputs[4750] = 1'b1;
    assign layer2_outputs[4751] = (layer1_outputs[2263]) & ~(layer1_outputs[2861]);
    assign layer2_outputs[4752] = layer1_outputs[312];
    assign layer2_outputs[4753] = (layer1_outputs[3451]) & (layer1_outputs[4036]);
    assign layer2_outputs[4754] = 1'b0;
    assign layer2_outputs[4755] = ~(layer1_outputs[912]);
    assign layer2_outputs[4756] = 1'b1;
    assign layer2_outputs[4757] = (layer1_outputs[4817]) & (layer1_outputs[2514]);
    assign layer2_outputs[4758] = (layer1_outputs[2496]) | (layer1_outputs[699]);
    assign layer2_outputs[4759] = layer1_outputs[640];
    assign layer2_outputs[4760] = (layer1_outputs[2540]) & ~(layer1_outputs[1968]);
    assign layer2_outputs[4761] = 1'b0;
    assign layer2_outputs[4762] = ~(layer1_outputs[3909]) | (layer1_outputs[4801]);
    assign layer2_outputs[4763] = ~((layer1_outputs[1759]) & (layer1_outputs[462]));
    assign layer2_outputs[4764] = layer1_outputs[2697];
    assign layer2_outputs[4765] = layer1_outputs[4206];
    assign layer2_outputs[4766] = ~(layer1_outputs[3524]) | (layer1_outputs[1864]);
    assign layer2_outputs[4767] = (layer1_outputs[3250]) & ~(layer1_outputs[3192]);
    assign layer2_outputs[4768] = (layer1_outputs[2235]) & ~(layer1_outputs[2924]);
    assign layer2_outputs[4769] = (layer1_outputs[4628]) & ~(layer1_outputs[2814]);
    assign layer2_outputs[4770] = ~((layer1_outputs[2016]) | (layer1_outputs[1643]));
    assign layer2_outputs[4771] = layer1_outputs[1919];
    assign layer2_outputs[4772] = ~(layer1_outputs[2151]) | (layer1_outputs[70]);
    assign layer2_outputs[4773] = (layer1_outputs[3846]) & ~(layer1_outputs[3431]);
    assign layer2_outputs[4774] = (layer1_outputs[1766]) & (layer1_outputs[2710]);
    assign layer2_outputs[4775] = ~(layer1_outputs[2569]) | (layer1_outputs[3500]);
    assign layer2_outputs[4776] = layer1_outputs[4677];
    assign layer2_outputs[4777] = layer1_outputs[1078];
    assign layer2_outputs[4778] = 1'b0;
    assign layer2_outputs[4779] = ~(layer1_outputs[3546]) | (layer1_outputs[1977]);
    assign layer2_outputs[4780] = 1'b0;
    assign layer2_outputs[4781] = (layer1_outputs[47]) | (layer1_outputs[4578]);
    assign layer2_outputs[4782] = (layer1_outputs[2903]) | (layer1_outputs[1236]);
    assign layer2_outputs[4783] = 1'b1;
    assign layer2_outputs[4784] = layer1_outputs[305];
    assign layer2_outputs[4785] = layer1_outputs[3014];
    assign layer2_outputs[4786] = ~(layer1_outputs[4099]);
    assign layer2_outputs[4787] = 1'b0;
    assign layer2_outputs[4788] = layer1_outputs[1885];
    assign layer2_outputs[4789] = ~(layer1_outputs[3825]);
    assign layer2_outputs[4790] = ~(layer1_outputs[4981]);
    assign layer2_outputs[4791] = layer1_outputs[31];
    assign layer2_outputs[4792] = layer1_outputs[4717];
    assign layer2_outputs[4793] = 1'b0;
    assign layer2_outputs[4794] = ~(layer1_outputs[1770]) | (layer1_outputs[5003]);
    assign layer2_outputs[4795] = ~(layer1_outputs[1471]);
    assign layer2_outputs[4796] = 1'b0;
    assign layer2_outputs[4797] = ~(layer1_outputs[1470]);
    assign layer2_outputs[4798] = layer1_outputs[2923];
    assign layer2_outputs[4799] = (layer1_outputs[2575]) & ~(layer1_outputs[932]);
    assign layer2_outputs[4800] = (layer1_outputs[2468]) | (layer1_outputs[3354]);
    assign layer2_outputs[4801] = ~(layer1_outputs[5114]);
    assign layer2_outputs[4802] = (layer1_outputs[1782]) | (layer1_outputs[397]);
    assign layer2_outputs[4803] = ~((layer1_outputs[992]) ^ (layer1_outputs[1623]));
    assign layer2_outputs[4804] = layer1_outputs[1182];
    assign layer2_outputs[4805] = layer1_outputs[487];
    assign layer2_outputs[4806] = (layer1_outputs[1012]) & ~(layer1_outputs[4486]);
    assign layer2_outputs[4807] = layer1_outputs[1904];
    assign layer2_outputs[4808] = (layer1_outputs[3165]) & (layer1_outputs[671]);
    assign layer2_outputs[4809] = (layer1_outputs[3617]) | (layer1_outputs[334]);
    assign layer2_outputs[4810] = layer1_outputs[612];
    assign layer2_outputs[4811] = ~(layer1_outputs[2762]) | (layer1_outputs[497]);
    assign layer2_outputs[4812] = layer1_outputs[850];
    assign layer2_outputs[4813] = layer1_outputs[1116];
    assign layer2_outputs[4814] = ~(layer1_outputs[3166]);
    assign layer2_outputs[4815] = 1'b1;
    assign layer2_outputs[4816] = ~(layer1_outputs[3782]);
    assign layer2_outputs[4817] = 1'b1;
    assign layer2_outputs[4818] = layer1_outputs[3183];
    assign layer2_outputs[4819] = 1'b1;
    assign layer2_outputs[4820] = layer1_outputs[3457];
    assign layer2_outputs[4821] = 1'b1;
    assign layer2_outputs[4822] = ~(layer1_outputs[1557]) | (layer1_outputs[1187]);
    assign layer2_outputs[4823] = layer1_outputs[1973];
    assign layer2_outputs[4824] = ~((layer1_outputs[3658]) | (layer1_outputs[3114]));
    assign layer2_outputs[4825] = 1'b0;
    assign layer2_outputs[4826] = ~(layer1_outputs[5057]) | (layer1_outputs[4649]);
    assign layer2_outputs[4827] = ~((layer1_outputs[4849]) & (layer1_outputs[49]));
    assign layer2_outputs[4828] = ~(layer1_outputs[2878]);
    assign layer2_outputs[4829] = ~(layer1_outputs[4642]);
    assign layer2_outputs[4830] = ~((layer1_outputs[3628]) & (layer1_outputs[1736]));
    assign layer2_outputs[4831] = (layer1_outputs[1925]) & (layer1_outputs[2059]);
    assign layer2_outputs[4832] = ~((layer1_outputs[4092]) & (layer1_outputs[1516]));
    assign layer2_outputs[4833] = ~((layer1_outputs[4106]) & (layer1_outputs[2471]));
    assign layer2_outputs[4834] = layer1_outputs[1591];
    assign layer2_outputs[4835] = layer1_outputs[56];
    assign layer2_outputs[4836] = (layer1_outputs[21]) ^ (layer1_outputs[2567]);
    assign layer2_outputs[4837] = ~(layer1_outputs[1336]);
    assign layer2_outputs[4838] = (layer1_outputs[4208]) & (layer1_outputs[1486]);
    assign layer2_outputs[4839] = layer1_outputs[1671];
    assign layer2_outputs[4840] = ~((layer1_outputs[413]) & (layer1_outputs[188]));
    assign layer2_outputs[4841] = (layer1_outputs[3253]) ^ (layer1_outputs[531]);
    assign layer2_outputs[4842] = ~(layer1_outputs[1240]);
    assign layer2_outputs[4843] = layer1_outputs[4732];
    assign layer2_outputs[4844] = ~(layer1_outputs[3623]);
    assign layer2_outputs[4845] = ~(layer1_outputs[590]);
    assign layer2_outputs[4846] = ~(layer1_outputs[1415]) | (layer1_outputs[2130]);
    assign layer2_outputs[4847] = layer1_outputs[4072];
    assign layer2_outputs[4848] = ~(layer1_outputs[2974]) | (layer1_outputs[108]);
    assign layer2_outputs[4849] = (layer1_outputs[1544]) & (layer1_outputs[3351]);
    assign layer2_outputs[4850] = 1'b0;
    assign layer2_outputs[4851] = 1'b0;
    assign layer2_outputs[4852] = ~((layer1_outputs[1170]) & (layer1_outputs[3002]));
    assign layer2_outputs[4853] = ~(layer1_outputs[1023]);
    assign layer2_outputs[4854] = (layer1_outputs[700]) & ~(layer1_outputs[1244]);
    assign layer2_outputs[4855] = layer1_outputs[1788];
    assign layer2_outputs[4856] = ~(layer1_outputs[108]) | (layer1_outputs[3091]);
    assign layer2_outputs[4857] = ~(layer1_outputs[4318]);
    assign layer2_outputs[4858] = (layer1_outputs[2576]) & ~(layer1_outputs[2250]);
    assign layer2_outputs[4859] = (layer1_outputs[3467]) & (layer1_outputs[2696]);
    assign layer2_outputs[4860] = ~(layer1_outputs[1903]) | (layer1_outputs[4963]);
    assign layer2_outputs[4861] = ~(layer1_outputs[2988]);
    assign layer2_outputs[4862] = (layer1_outputs[137]) & (layer1_outputs[1134]);
    assign layer2_outputs[4863] = ~(layer1_outputs[3284]);
    assign layer2_outputs[4864] = (layer1_outputs[3605]) & ~(layer1_outputs[991]);
    assign layer2_outputs[4865] = ~((layer1_outputs[3065]) & (layer1_outputs[3490]));
    assign layer2_outputs[4866] = ~(layer1_outputs[3438]);
    assign layer2_outputs[4867] = ~((layer1_outputs[2902]) & (layer1_outputs[3750]));
    assign layer2_outputs[4868] = (layer1_outputs[4988]) | (layer1_outputs[2833]);
    assign layer2_outputs[4869] = ~(layer1_outputs[650]) | (layer1_outputs[595]);
    assign layer2_outputs[4870] = (layer1_outputs[4627]) & (layer1_outputs[5098]);
    assign layer2_outputs[4871] = ~((layer1_outputs[3048]) & (layer1_outputs[4234]));
    assign layer2_outputs[4872] = ~((layer1_outputs[657]) ^ (layer1_outputs[2121]));
    assign layer2_outputs[4873] = ~((layer1_outputs[4313]) | (layer1_outputs[3390]));
    assign layer2_outputs[4874] = ~(layer1_outputs[2392]) | (layer1_outputs[651]);
    assign layer2_outputs[4875] = ~(layer1_outputs[3169]);
    assign layer2_outputs[4876] = 1'b1;
    assign layer2_outputs[4877] = 1'b0;
    assign layer2_outputs[4878] = ~((layer1_outputs[3930]) & (layer1_outputs[3439]));
    assign layer2_outputs[4879] = (layer1_outputs[2337]) & (layer1_outputs[4209]);
    assign layer2_outputs[4880] = (layer1_outputs[2912]) & ~(layer1_outputs[1981]);
    assign layer2_outputs[4881] = 1'b1;
    assign layer2_outputs[4882] = ~(layer1_outputs[1202]);
    assign layer2_outputs[4883] = layer1_outputs[4677];
    assign layer2_outputs[4884] = ~(layer1_outputs[3743]);
    assign layer2_outputs[4885] = ~(layer1_outputs[809]);
    assign layer2_outputs[4886] = layer1_outputs[3928];
    assign layer2_outputs[4887] = (layer1_outputs[3270]) & ~(layer1_outputs[159]);
    assign layer2_outputs[4888] = ~(layer1_outputs[4651]);
    assign layer2_outputs[4889] = layer1_outputs[1020];
    assign layer2_outputs[4890] = ~((layer1_outputs[3146]) | (layer1_outputs[1481]));
    assign layer2_outputs[4891] = (layer1_outputs[1909]) & ~(layer1_outputs[998]);
    assign layer2_outputs[4892] = ~(layer1_outputs[3128]) | (layer1_outputs[2654]);
    assign layer2_outputs[4893] = (layer1_outputs[771]) & ~(layer1_outputs[623]);
    assign layer2_outputs[4894] = 1'b0;
    assign layer2_outputs[4895] = ~((layer1_outputs[3120]) | (layer1_outputs[4971]));
    assign layer2_outputs[4896] = layer1_outputs[3791];
    assign layer2_outputs[4897] = layer1_outputs[1209];
    assign layer2_outputs[4898] = 1'b1;
    assign layer2_outputs[4899] = ~(layer1_outputs[4431]);
    assign layer2_outputs[4900] = ~((layer1_outputs[3746]) | (layer1_outputs[4975]));
    assign layer2_outputs[4901] = ~(layer1_outputs[4392]);
    assign layer2_outputs[4902] = (layer1_outputs[4198]) & ~(layer1_outputs[3886]);
    assign layer2_outputs[4903] = (layer1_outputs[1162]) | (layer1_outputs[1415]);
    assign layer2_outputs[4904] = layer1_outputs[552];
    assign layer2_outputs[4905] = layer1_outputs[945];
    assign layer2_outputs[4906] = ~(layer1_outputs[1740]) | (layer1_outputs[4442]);
    assign layer2_outputs[4907] = ~(layer1_outputs[857]);
    assign layer2_outputs[4908] = ~((layer1_outputs[3707]) & (layer1_outputs[419]));
    assign layer2_outputs[4909] = 1'b1;
    assign layer2_outputs[4910] = (layer1_outputs[4192]) & ~(layer1_outputs[940]);
    assign layer2_outputs[4911] = 1'b1;
    assign layer2_outputs[4912] = ~((layer1_outputs[780]) | (layer1_outputs[3129]));
    assign layer2_outputs[4913] = ~((layer1_outputs[3156]) & (layer1_outputs[4543]));
    assign layer2_outputs[4914] = ~((layer1_outputs[5016]) | (layer1_outputs[4550]));
    assign layer2_outputs[4915] = (layer1_outputs[2740]) | (layer1_outputs[3983]);
    assign layer2_outputs[4916] = ~(layer1_outputs[135]);
    assign layer2_outputs[4917] = (layer1_outputs[3583]) ^ (layer1_outputs[1933]);
    assign layer2_outputs[4918] = ~(layer1_outputs[1033]);
    assign layer2_outputs[4919] = (layer1_outputs[826]) & ~(layer1_outputs[2189]);
    assign layer2_outputs[4920] = (layer1_outputs[5007]) & ~(layer1_outputs[683]);
    assign layer2_outputs[4921] = (layer1_outputs[4817]) & ~(layer1_outputs[1163]);
    assign layer2_outputs[4922] = layer1_outputs[5039];
    assign layer2_outputs[4923] = (layer1_outputs[2068]) | (layer1_outputs[4211]);
    assign layer2_outputs[4924] = (layer1_outputs[2015]) & ~(layer1_outputs[4890]);
    assign layer2_outputs[4925] = ~((layer1_outputs[4388]) & (layer1_outputs[3410]));
    assign layer2_outputs[4926] = (layer1_outputs[482]) | (layer1_outputs[3446]);
    assign layer2_outputs[4927] = ~((layer1_outputs[1228]) & (layer1_outputs[80]));
    assign layer2_outputs[4928] = layer1_outputs[3556];
    assign layer2_outputs[4929] = 1'b1;
    assign layer2_outputs[4930] = ~((layer1_outputs[2860]) & (layer1_outputs[2646]));
    assign layer2_outputs[4931] = (layer1_outputs[3644]) & ~(layer1_outputs[3226]);
    assign layer2_outputs[4932] = (layer1_outputs[1679]) ^ (layer1_outputs[1752]);
    assign layer2_outputs[4933] = ~((layer1_outputs[4482]) ^ (layer1_outputs[3573]));
    assign layer2_outputs[4934] = 1'b1;
    assign layer2_outputs[4935] = ~(layer1_outputs[1259]);
    assign layer2_outputs[4936] = 1'b0;
    assign layer2_outputs[4937] = (layer1_outputs[1397]) & ~(layer1_outputs[4948]);
    assign layer2_outputs[4938] = layer1_outputs[2248];
    assign layer2_outputs[4939] = 1'b1;
    assign layer2_outputs[4940] = ~(layer1_outputs[2934]);
    assign layer2_outputs[4941] = ~(layer1_outputs[4588]);
    assign layer2_outputs[4942] = ~(layer1_outputs[3857]);
    assign layer2_outputs[4943] = ~((layer1_outputs[4866]) ^ (layer1_outputs[3504]));
    assign layer2_outputs[4944] = (layer1_outputs[4919]) & (layer1_outputs[4368]);
    assign layer2_outputs[4945] = layer1_outputs[102];
    assign layer2_outputs[4946] = layer1_outputs[1350];
    assign layer2_outputs[4947] = ~(layer1_outputs[4381]) | (layer1_outputs[841]);
    assign layer2_outputs[4948] = 1'b1;
    assign layer2_outputs[4949] = ~((layer1_outputs[3953]) | (layer1_outputs[2047]));
    assign layer2_outputs[4950] = ~(layer1_outputs[2283]);
    assign layer2_outputs[4951] = ~(layer1_outputs[591]);
    assign layer2_outputs[4952] = ~((layer1_outputs[643]) ^ (layer1_outputs[966]));
    assign layer2_outputs[4953] = ~(layer1_outputs[4612]);
    assign layer2_outputs[4954] = ~((layer1_outputs[1823]) | (layer1_outputs[5070]));
    assign layer2_outputs[4955] = ~(layer1_outputs[1997]);
    assign layer2_outputs[4956] = 1'b1;
    assign layer2_outputs[4957] = (layer1_outputs[4153]) & ~(layer1_outputs[160]);
    assign layer2_outputs[4958] = ~((layer1_outputs[1545]) & (layer1_outputs[3879]));
    assign layer2_outputs[4959] = ~(layer1_outputs[4008]);
    assign layer2_outputs[4960] = layer1_outputs[3206];
    assign layer2_outputs[4961] = ~((layer1_outputs[4180]) & (layer1_outputs[1684]));
    assign layer2_outputs[4962] = ~(layer1_outputs[3093]);
    assign layer2_outputs[4963] = 1'b0;
    assign layer2_outputs[4964] = ~(layer1_outputs[1600]) | (layer1_outputs[4188]);
    assign layer2_outputs[4965] = (layer1_outputs[934]) & (layer1_outputs[12]);
    assign layer2_outputs[4966] = 1'b0;
    assign layer2_outputs[4967] = layer1_outputs[4059];
    assign layer2_outputs[4968] = (layer1_outputs[1046]) & ~(layer1_outputs[4346]);
    assign layer2_outputs[4969] = layer1_outputs[355];
    assign layer2_outputs[4970] = ~(layer1_outputs[768]) | (layer1_outputs[1760]);
    assign layer2_outputs[4971] = ~(layer1_outputs[1012]) | (layer1_outputs[3506]);
    assign layer2_outputs[4972] = ~(layer1_outputs[2822]);
    assign layer2_outputs[4973] = (layer1_outputs[3082]) & ~(layer1_outputs[275]);
    assign layer2_outputs[4974] = 1'b1;
    assign layer2_outputs[4975] = ~(layer1_outputs[3125]);
    assign layer2_outputs[4976] = ~(layer1_outputs[4141]);
    assign layer2_outputs[4977] = ~(layer1_outputs[3688]) | (layer1_outputs[1700]);
    assign layer2_outputs[4978] = 1'b1;
    assign layer2_outputs[4979] = ~(layer1_outputs[4114]);
    assign layer2_outputs[4980] = ~(layer1_outputs[3355]) | (layer1_outputs[5094]);
    assign layer2_outputs[4981] = 1'b1;
    assign layer2_outputs[4982] = (layer1_outputs[1796]) | (layer1_outputs[960]);
    assign layer2_outputs[4983] = ~(layer1_outputs[1369]);
    assign layer2_outputs[4984] = layer1_outputs[2173];
    assign layer2_outputs[4985] = ~(layer1_outputs[1194]);
    assign layer2_outputs[4986] = ~(layer1_outputs[2378]);
    assign layer2_outputs[4987] = 1'b0;
    assign layer2_outputs[4988] = ~(layer1_outputs[5044]) | (layer1_outputs[582]);
    assign layer2_outputs[4989] = (layer1_outputs[2319]) & ~(layer1_outputs[2755]);
    assign layer2_outputs[4990] = layer1_outputs[4783];
    assign layer2_outputs[4991] = ~((layer1_outputs[2774]) | (layer1_outputs[4975]));
    assign layer2_outputs[4992] = ~(layer1_outputs[212]) | (layer1_outputs[4206]);
    assign layer2_outputs[4993] = ~(layer1_outputs[1199]) | (layer1_outputs[510]);
    assign layer2_outputs[4994] = ~((layer1_outputs[181]) & (layer1_outputs[4231]));
    assign layer2_outputs[4995] = (layer1_outputs[811]) | (layer1_outputs[1962]);
    assign layer2_outputs[4996] = (layer1_outputs[1801]) & ~(layer1_outputs[2547]);
    assign layer2_outputs[4997] = layer1_outputs[3474];
    assign layer2_outputs[4998] = ~((layer1_outputs[2038]) | (layer1_outputs[4878]));
    assign layer2_outputs[4999] = ~((layer1_outputs[271]) & (layer1_outputs[2616]));
    assign layer2_outputs[5000] = 1'b1;
    assign layer2_outputs[5001] = ~((layer1_outputs[1952]) & (layer1_outputs[5080]));
    assign layer2_outputs[5002] = 1'b1;
    assign layer2_outputs[5003] = ~(layer1_outputs[2174]);
    assign layer2_outputs[5004] = ~(layer1_outputs[4784]);
    assign layer2_outputs[5005] = (layer1_outputs[3159]) & ~(layer1_outputs[4283]);
    assign layer2_outputs[5006] = ~(layer1_outputs[4173]);
    assign layer2_outputs[5007] = layer1_outputs[4288];
    assign layer2_outputs[5008] = 1'b0;
    assign layer2_outputs[5009] = (layer1_outputs[411]) & ~(layer1_outputs[2742]);
    assign layer2_outputs[5010] = (layer1_outputs[556]) | (layer1_outputs[1746]);
    assign layer2_outputs[5011] = (layer1_outputs[2907]) & (layer1_outputs[2271]);
    assign layer2_outputs[5012] = ~(layer1_outputs[3241]);
    assign layer2_outputs[5013] = (layer1_outputs[2287]) & ~(layer1_outputs[4914]);
    assign layer2_outputs[5014] = ~(layer1_outputs[2285]);
    assign layer2_outputs[5015] = ~(layer1_outputs[1270]);
    assign layer2_outputs[5016] = 1'b0;
    assign layer2_outputs[5017] = layer1_outputs[4933];
    assign layer2_outputs[5018] = ~((layer1_outputs[853]) & (layer1_outputs[2723]));
    assign layer2_outputs[5019] = (layer1_outputs[2780]) & ~(layer1_outputs[3009]);
    assign layer2_outputs[5020] = 1'b1;
    assign layer2_outputs[5021] = ~(layer1_outputs[1430]);
    assign layer2_outputs[5022] = (layer1_outputs[4743]) & ~(layer1_outputs[4598]);
    assign layer2_outputs[5023] = ~(layer1_outputs[4175]);
    assign layer2_outputs[5024] = ~(layer1_outputs[3005]) | (layer1_outputs[3287]);
    assign layer2_outputs[5025] = ~((layer1_outputs[1539]) & (layer1_outputs[1917]));
    assign layer2_outputs[5026] = ~(layer1_outputs[3184]);
    assign layer2_outputs[5027] = ~(layer1_outputs[905]);
    assign layer2_outputs[5028] = (layer1_outputs[2179]) & (layer1_outputs[2770]);
    assign layer2_outputs[5029] = ~((layer1_outputs[4351]) | (layer1_outputs[2098]));
    assign layer2_outputs[5030] = layer1_outputs[4528];
    assign layer2_outputs[5031] = ~((layer1_outputs[2158]) | (layer1_outputs[4452]));
    assign layer2_outputs[5032] = (layer1_outputs[4414]) & ~(layer1_outputs[4389]);
    assign layer2_outputs[5033] = ~((layer1_outputs[4542]) & (layer1_outputs[2932]));
    assign layer2_outputs[5034] = (layer1_outputs[3152]) & ~(layer1_outputs[4102]);
    assign layer2_outputs[5035] = ~(layer1_outputs[4174]);
    assign layer2_outputs[5036] = (layer1_outputs[578]) & (layer1_outputs[2626]);
    assign layer2_outputs[5037] = ~(layer1_outputs[1886]);
    assign layer2_outputs[5038] = (layer1_outputs[715]) & ~(layer1_outputs[3198]);
    assign layer2_outputs[5039] = ~(layer1_outputs[4218]);
    assign layer2_outputs[5040] = layer1_outputs[2683];
    assign layer2_outputs[5041] = ~(layer1_outputs[37]);
    assign layer2_outputs[5042] = 1'b0;
    assign layer2_outputs[5043] = ~(layer1_outputs[755]) | (layer1_outputs[120]);
    assign layer2_outputs[5044] = ~(layer1_outputs[98]);
    assign layer2_outputs[5045] = ~(layer1_outputs[3116]);
    assign layer2_outputs[5046] = ~(layer1_outputs[460]) | (layer1_outputs[970]);
    assign layer2_outputs[5047] = (layer1_outputs[1948]) & (layer1_outputs[3761]);
    assign layer2_outputs[5048] = layer1_outputs[4552];
    assign layer2_outputs[5049] = (layer1_outputs[4051]) & (layer1_outputs[2538]);
    assign layer2_outputs[5050] = (layer1_outputs[5010]) & ~(layer1_outputs[2506]);
    assign layer2_outputs[5051] = ~(layer1_outputs[927]);
    assign layer2_outputs[5052] = layer1_outputs[2610];
    assign layer2_outputs[5053] = (layer1_outputs[4043]) & (layer1_outputs[632]);
    assign layer2_outputs[5054] = (layer1_outputs[4095]) | (layer1_outputs[2578]);
    assign layer2_outputs[5055] = 1'b1;
    assign layer2_outputs[5056] = ~(layer1_outputs[1374]);
    assign layer2_outputs[5057] = ~(layer1_outputs[3049]);
    assign layer2_outputs[5058] = ~((layer1_outputs[408]) ^ (layer1_outputs[4776]));
    assign layer2_outputs[5059] = 1'b0;
    assign layer2_outputs[5060] = (layer1_outputs[2514]) & ~(layer1_outputs[4055]);
    assign layer2_outputs[5061] = ~(layer1_outputs[5087]);
    assign layer2_outputs[5062] = (layer1_outputs[953]) & (layer1_outputs[2612]);
    assign layer2_outputs[5063] = layer1_outputs[4928];
    assign layer2_outputs[5064] = ~(layer1_outputs[2791]);
    assign layer2_outputs[5065] = 1'b0;
    assign layer2_outputs[5066] = (layer1_outputs[2186]) & ~(layer1_outputs[1215]);
    assign layer2_outputs[5067] = (layer1_outputs[291]) & ~(layer1_outputs[2301]);
    assign layer2_outputs[5068] = layer1_outputs[1654];
    assign layer2_outputs[5069] = ~((layer1_outputs[749]) & (layer1_outputs[3388]));
    assign layer2_outputs[5070] = 1'b1;
    assign layer2_outputs[5071] = ~(layer1_outputs[1125]);
    assign layer2_outputs[5072] = 1'b0;
    assign layer2_outputs[5073] = ~(layer1_outputs[3042]);
    assign layer2_outputs[5074] = layer1_outputs[398];
    assign layer2_outputs[5075] = (layer1_outputs[1239]) & ~(layer1_outputs[4807]);
    assign layer2_outputs[5076] = ~(layer1_outputs[2893]);
    assign layer2_outputs[5077] = ~((layer1_outputs[2418]) & (layer1_outputs[803]));
    assign layer2_outputs[5078] = ~((layer1_outputs[3039]) & (layer1_outputs[1095]));
    assign layer2_outputs[5079] = layer1_outputs[3224];
    assign layer2_outputs[5080] = ~((layer1_outputs[253]) | (layer1_outputs[4895]));
    assign layer2_outputs[5081] = ~(layer1_outputs[4802]) | (layer1_outputs[3130]);
    assign layer2_outputs[5082] = layer1_outputs[4075];
    assign layer2_outputs[5083] = ~(layer1_outputs[2523]);
    assign layer2_outputs[5084] = ~(layer1_outputs[141]) | (layer1_outputs[1198]);
    assign layer2_outputs[5085] = ~((layer1_outputs[3092]) & (layer1_outputs[4804]));
    assign layer2_outputs[5086] = (layer1_outputs[2440]) & ~(layer1_outputs[2900]);
    assign layer2_outputs[5087] = ~((layer1_outputs[4721]) | (layer1_outputs[3606]));
    assign layer2_outputs[5088] = (layer1_outputs[3155]) | (layer1_outputs[954]);
    assign layer2_outputs[5089] = ~(layer1_outputs[1791]);
    assign layer2_outputs[5090] = ~((layer1_outputs[3453]) | (layer1_outputs[3171]));
    assign layer2_outputs[5091] = layer1_outputs[4428];
    assign layer2_outputs[5092] = (layer1_outputs[3844]) & ~(layer1_outputs[3275]);
    assign layer2_outputs[5093] = layer1_outputs[2630];
    assign layer2_outputs[5094] = layer1_outputs[422];
    assign layer2_outputs[5095] = layer1_outputs[542];
    assign layer2_outputs[5096] = (layer1_outputs[586]) & ~(layer1_outputs[196]);
    assign layer2_outputs[5097] = ~((layer1_outputs[2169]) | (layer1_outputs[4072]));
    assign layer2_outputs[5098] = (layer1_outputs[1913]) ^ (layer1_outputs[3863]);
    assign layer2_outputs[5099] = layer1_outputs[4774];
    assign layer2_outputs[5100] = (layer1_outputs[1812]) & ~(layer1_outputs[2292]);
    assign layer2_outputs[5101] = layer1_outputs[1873];
    assign layer2_outputs[5102] = ~(layer1_outputs[3169]);
    assign layer2_outputs[5103] = layer1_outputs[3075];
    assign layer2_outputs[5104] = ~(layer1_outputs[2561]) | (layer1_outputs[3075]);
    assign layer2_outputs[5105] = ~(layer1_outputs[2307]);
    assign layer2_outputs[5106] = layer1_outputs[1945];
    assign layer2_outputs[5107] = ~(layer1_outputs[2942]) | (layer1_outputs[1560]);
    assign layer2_outputs[5108] = (layer1_outputs[4052]) & ~(layer1_outputs[39]);
    assign layer2_outputs[5109] = layer1_outputs[3173];
    assign layer2_outputs[5110] = (layer1_outputs[4748]) & (layer1_outputs[4063]);
    assign layer2_outputs[5111] = ~(layer1_outputs[909]);
    assign layer2_outputs[5112] = layer1_outputs[1771];
    assign layer2_outputs[5113] = ~(layer1_outputs[3821]) | (layer1_outputs[5089]);
    assign layer2_outputs[5114] = 1'b0;
    assign layer2_outputs[5115] = ~((layer1_outputs[1004]) ^ (layer1_outputs[476]));
    assign layer2_outputs[5116] = 1'b1;
    assign layer2_outputs[5117] = (layer1_outputs[1937]) & ~(layer1_outputs[5117]);
    assign layer2_outputs[5118] = layer1_outputs[4810];
    assign layer2_outputs[5119] = layer1_outputs[4284];
    assign layer3_outputs[0] = 1'b0;
    assign layer3_outputs[1] = ~(layer2_outputs[2410]);
    assign layer3_outputs[2] = (layer2_outputs[1137]) & ~(layer2_outputs[3348]);
    assign layer3_outputs[3] = ~(layer2_outputs[1750]) | (layer2_outputs[131]);
    assign layer3_outputs[4] = layer2_outputs[535];
    assign layer3_outputs[5] = ~(layer2_outputs[646]);
    assign layer3_outputs[6] = 1'b1;
    assign layer3_outputs[7] = (layer2_outputs[3867]) & ~(layer2_outputs[5033]);
    assign layer3_outputs[8] = ~(layer2_outputs[4796]) | (layer2_outputs[4247]);
    assign layer3_outputs[9] = ~(layer2_outputs[462]);
    assign layer3_outputs[10] = (layer2_outputs[2044]) & ~(layer2_outputs[1686]);
    assign layer3_outputs[11] = 1'b0;
    assign layer3_outputs[12] = 1'b1;
    assign layer3_outputs[13] = (layer2_outputs[3280]) & ~(layer2_outputs[812]);
    assign layer3_outputs[14] = ~((layer2_outputs[3322]) & (layer2_outputs[4235]));
    assign layer3_outputs[15] = (layer2_outputs[4711]) | (layer2_outputs[2013]);
    assign layer3_outputs[16] = (layer2_outputs[1267]) & (layer2_outputs[3309]);
    assign layer3_outputs[17] = ~((layer2_outputs[3323]) & (layer2_outputs[3300]));
    assign layer3_outputs[18] = layer2_outputs[1306];
    assign layer3_outputs[19] = ~((layer2_outputs[2368]) & (layer2_outputs[1945]));
    assign layer3_outputs[20] = (layer2_outputs[2071]) | (layer2_outputs[468]);
    assign layer3_outputs[21] = ~((layer2_outputs[4024]) & (layer2_outputs[597]));
    assign layer3_outputs[22] = ~(layer2_outputs[4951]) | (layer2_outputs[4359]);
    assign layer3_outputs[23] = ~(layer2_outputs[3878]);
    assign layer3_outputs[24] = (layer2_outputs[1448]) & (layer2_outputs[4710]);
    assign layer3_outputs[25] = (layer2_outputs[1275]) & (layer2_outputs[406]);
    assign layer3_outputs[26] = ~(layer2_outputs[2281]);
    assign layer3_outputs[27] = ~(layer2_outputs[259]) | (layer2_outputs[2488]);
    assign layer3_outputs[28] = ~(layer2_outputs[2934]);
    assign layer3_outputs[29] = layer2_outputs[1653];
    assign layer3_outputs[30] = ~((layer2_outputs[1605]) | (layer2_outputs[3761]));
    assign layer3_outputs[31] = (layer2_outputs[2444]) | (layer2_outputs[1702]);
    assign layer3_outputs[32] = (layer2_outputs[3032]) & ~(layer2_outputs[4675]);
    assign layer3_outputs[33] = layer2_outputs[3991];
    assign layer3_outputs[34] = (layer2_outputs[3629]) & ~(layer2_outputs[2770]);
    assign layer3_outputs[35] = ~((layer2_outputs[5055]) ^ (layer2_outputs[3739]));
    assign layer3_outputs[36] = ~((layer2_outputs[966]) & (layer2_outputs[2810]));
    assign layer3_outputs[37] = layer2_outputs[4180];
    assign layer3_outputs[38] = ~((layer2_outputs[88]) ^ (layer2_outputs[2069]));
    assign layer3_outputs[39] = ~(layer2_outputs[1097]) | (layer2_outputs[1840]);
    assign layer3_outputs[40] = ~((layer2_outputs[2318]) | (layer2_outputs[414]));
    assign layer3_outputs[41] = ~(layer2_outputs[2530]);
    assign layer3_outputs[42] = ~(layer2_outputs[4823]);
    assign layer3_outputs[43] = ~((layer2_outputs[729]) | (layer2_outputs[2417]));
    assign layer3_outputs[44] = ~(layer2_outputs[4327]);
    assign layer3_outputs[45] = layer2_outputs[58];
    assign layer3_outputs[46] = (layer2_outputs[2719]) & (layer2_outputs[2694]);
    assign layer3_outputs[47] = (layer2_outputs[1028]) & ~(layer2_outputs[4830]);
    assign layer3_outputs[48] = layer2_outputs[4397];
    assign layer3_outputs[49] = 1'b0;
    assign layer3_outputs[50] = (layer2_outputs[3522]) | (layer2_outputs[4362]);
    assign layer3_outputs[51] = ~(layer2_outputs[195]) | (layer2_outputs[2145]);
    assign layer3_outputs[52] = layer2_outputs[2539];
    assign layer3_outputs[53] = ~((layer2_outputs[3134]) | (layer2_outputs[2779]));
    assign layer3_outputs[54] = ~(layer2_outputs[534]);
    assign layer3_outputs[55] = layer2_outputs[4972];
    assign layer3_outputs[56] = (layer2_outputs[5069]) | (layer2_outputs[512]);
    assign layer3_outputs[57] = ~(layer2_outputs[619]);
    assign layer3_outputs[58] = 1'b0;
    assign layer3_outputs[59] = (layer2_outputs[3458]) & (layer2_outputs[3560]);
    assign layer3_outputs[60] = ~(layer2_outputs[4854]) | (layer2_outputs[5062]);
    assign layer3_outputs[61] = layer2_outputs[3121];
    assign layer3_outputs[62] = layer2_outputs[4689];
    assign layer3_outputs[63] = (layer2_outputs[2945]) & (layer2_outputs[4572]);
    assign layer3_outputs[64] = ~(layer2_outputs[4432]);
    assign layer3_outputs[65] = layer2_outputs[1335];
    assign layer3_outputs[66] = ~(layer2_outputs[994]) | (layer2_outputs[3151]);
    assign layer3_outputs[67] = ~(layer2_outputs[77]);
    assign layer3_outputs[68] = 1'b1;
    assign layer3_outputs[69] = ~((layer2_outputs[414]) & (layer2_outputs[2265]));
    assign layer3_outputs[70] = ~((layer2_outputs[523]) & (layer2_outputs[2150]));
    assign layer3_outputs[71] = ~(layer2_outputs[1995]) | (layer2_outputs[2]);
    assign layer3_outputs[72] = ~(layer2_outputs[4944]) | (layer2_outputs[993]);
    assign layer3_outputs[73] = ~((layer2_outputs[1360]) & (layer2_outputs[3462]));
    assign layer3_outputs[74] = ~((layer2_outputs[3479]) & (layer2_outputs[4755]));
    assign layer3_outputs[75] = ~((layer2_outputs[4480]) & (layer2_outputs[2541]));
    assign layer3_outputs[76] = ~(layer2_outputs[1659]);
    assign layer3_outputs[77] = layer2_outputs[2635];
    assign layer3_outputs[78] = (layer2_outputs[19]) & ~(layer2_outputs[109]);
    assign layer3_outputs[79] = layer2_outputs[391];
    assign layer3_outputs[80] = ~(layer2_outputs[1883]) | (layer2_outputs[1420]);
    assign layer3_outputs[81] = ~(layer2_outputs[128]) | (layer2_outputs[2361]);
    assign layer3_outputs[82] = (layer2_outputs[1826]) | (layer2_outputs[3179]);
    assign layer3_outputs[83] = ~(layer2_outputs[1685]);
    assign layer3_outputs[84] = ~(layer2_outputs[3810]);
    assign layer3_outputs[85] = ~(layer2_outputs[533]);
    assign layer3_outputs[86] = 1'b1;
    assign layer3_outputs[87] = ~(layer2_outputs[3400]);
    assign layer3_outputs[88] = layer2_outputs[4376];
    assign layer3_outputs[89] = ~((layer2_outputs[360]) & (layer2_outputs[724]));
    assign layer3_outputs[90] = 1'b1;
    assign layer3_outputs[91] = ~((layer2_outputs[4686]) & (layer2_outputs[910]));
    assign layer3_outputs[92] = ~((layer2_outputs[4390]) & (layer2_outputs[3594]));
    assign layer3_outputs[93] = ~(layer2_outputs[2959]);
    assign layer3_outputs[94] = ~((layer2_outputs[2639]) | (layer2_outputs[3012]));
    assign layer3_outputs[95] = (layer2_outputs[4042]) & (layer2_outputs[1789]);
    assign layer3_outputs[96] = ~(layer2_outputs[229]);
    assign layer3_outputs[97] = ~(layer2_outputs[2564]) | (layer2_outputs[984]);
    assign layer3_outputs[98] = (layer2_outputs[1091]) | (layer2_outputs[2314]);
    assign layer3_outputs[99] = ~((layer2_outputs[4518]) ^ (layer2_outputs[1493]));
    assign layer3_outputs[100] = ~(layer2_outputs[3372]);
    assign layer3_outputs[101] = (layer2_outputs[2898]) & (layer2_outputs[1535]);
    assign layer3_outputs[102] = (layer2_outputs[3080]) | (layer2_outputs[3739]);
    assign layer3_outputs[103] = ~(layer2_outputs[4052]);
    assign layer3_outputs[104] = (layer2_outputs[4318]) & ~(layer2_outputs[4681]);
    assign layer3_outputs[105] = layer2_outputs[2929];
    assign layer3_outputs[106] = 1'b1;
    assign layer3_outputs[107] = ~(layer2_outputs[1159]) | (layer2_outputs[1933]);
    assign layer3_outputs[108] = ~(layer2_outputs[1568]);
    assign layer3_outputs[109] = 1'b0;
    assign layer3_outputs[110] = ~(layer2_outputs[3142]) | (layer2_outputs[2440]);
    assign layer3_outputs[111] = 1'b1;
    assign layer3_outputs[112] = ~((layer2_outputs[3795]) & (layer2_outputs[1269]));
    assign layer3_outputs[113] = ~(layer2_outputs[3265]);
    assign layer3_outputs[114] = ~(layer2_outputs[3989]) | (layer2_outputs[3777]);
    assign layer3_outputs[115] = layer2_outputs[2346];
    assign layer3_outputs[116] = 1'b0;
    assign layer3_outputs[117] = 1'b1;
    assign layer3_outputs[118] = ~(layer2_outputs[3554]) | (layer2_outputs[4507]);
    assign layer3_outputs[119] = ~((layer2_outputs[4680]) | (layer2_outputs[2951]));
    assign layer3_outputs[120] = 1'b0;
    assign layer3_outputs[121] = (layer2_outputs[2295]) ^ (layer2_outputs[4324]);
    assign layer3_outputs[122] = 1'b0;
    assign layer3_outputs[123] = ~((layer2_outputs[4569]) & (layer2_outputs[3646]));
    assign layer3_outputs[124] = layer2_outputs[2356];
    assign layer3_outputs[125] = ~(layer2_outputs[109]);
    assign layer3_outputs[126] = ~(layer2_outputs[4697]);
    assign layer3_outputs[127] = (layer2_outputs[3427]) & ~(layer2_outputs[2773]);
    assign layer3_outputs[128] = layer2_outputs[4182];
    assign layer3_outputs[129] = ~(layer2_outputs[4271]);
    assign layer3_outputs[130] = ~(layer2_outputs[896]);
    assign layer3_outputs[131] = layer2_outputs[574];
    assign layer3_outputs[132] = layer2_outputs[3385];
    assign layer3_outputs[133] = (layer2_outputs[2249]) & ~(layer2_outputs[1646]);
    assign layer3_outputs[134] = ~(layer2_outputs[1369]);
    assign layer3_outputs[135] = ~(layer2_outputs[4915]);
    assign layer3_outputs[136] = layer2_outputs[2296];
    assign layer3_outputs[137] = 1'b0;
    assign layer3_outputs[138] = layer2_outputs[5105];
    assign layer3_outputs[139] = ~(layer2_outputs[952]) | (layer2_outputs[4386]);
    assign layer3_outputs[140] = (layer2_outputs[484]) & ~(layer2_outputs[1913]);
    assign layer3_outputs[141] = ~(layer2_outputs[3668]) | (layer2_outputs[5003]);
    assign layer3_outputs[142] = (layer2_outputs[224]) & ~(layer2_outputs[1424]);
    assign layer3_outputs[143] = layer2_outputs[4249];
    assign layer3_outputs[144] = ~((layer2_outputs[4749]) & (layer2_outputs[2937]));
    assign layer3_outputs[145] = ~(layer2_outputs[469]) | (layer2_outputs[948]);
    assign layer3_outputs[146] = ~(layer2_outputs[558]);
    assign layer3_outputs[147] = (layer2_outputs[4576]) & ~(layer2_outputs[3387]);
    assign layer3_outputs[148] = ~((layer2_outputs[2235]) ^ (layer2_outputs[573]));
    assign layer3_outputs[149] = layer2_outputs[2781];
    assign layer3_outputs[150] = ~((layer2_outputs[1080]) & (layer2_outputs[1151]));
    assign layer3_outputs[151] = ~(layer2_outputs[4165]) | (layer2_outputs[3393]);
    assign layer3_outputs[152] = ~(layer2_outputs[4431]);
    assign layer3_outputs[153] = 1'b0;
    assign layer3_outputs[154] = (layer2_outputs[1074]) & (layer2_outputs[2921]);
    assign layer3_outputs[155] = ~(layer2_outputs[3721]);
    assign layer3_outputs[156] = ~(layer2_outputs[1068]);
    assign layer3_outputs[157] = ~(layer2_outputs[2419]) | (layer2_outputs[4982]);
    assign layer3_outputs[158] = (layer2_outputs[3791]) & ~(layer2_outputs[1266]);
    assign layer3_outputs[159] = (layer2_outputs[1084]) & ~(layer2_outputs[4575]);
    assign layer3_outputs[160] = (layer2_outputs[4031]) ^ (layer2_outputs[2182]);
    assign layer3_outputs[161] = (layer2_outputs[2362]) & (layer2_outputs[1190]);
    assign layer3_outputs[162] = 1'b0;
    assign layer3_outputs[163] = ~(layer2_outputs[1378]) | (layer2_outputs[1524]);
    assign layer3_outputs[164] = 1'b1;
    assign layer3_outputs[165] = (layer2_outputs[5040]) & ~(layer2_outputs[4348]);
    assign layer3_outputs[166] = ~(layer2_outputs[1547]);
    assign layer3_outputs[167] = 1'b0;
    assign layer3_outputs[168] = ~(layer2_outputs[3316]);
    assign layer3_outputs[169] = ~(layer2_outputs[3376]) | (layer2_outputs[2078]);
    assign layer3_outputs[170] = (layer2_outputs[1829]) | (layer2_outputs[2724]);
    assign layer3_outputs[171] = ~(layer2_outputs[3934]) | (layer2_outputs[1151]);
    assign layer3_outputs[172] = ~(layer2_outputs[1865]) | (layer2_outputs[2376]);
    assign layer3_outputs[173] = ~(layer2_outputs[303]);
    assign layer3_outputs[174] = 1'b1;
    assign layer3_outputs[175] = ~(layer2_outputs[2480]);
    assign layer3_outputs[176] = ~(layer2_outputs[1243]);
    assign layer3_outputs[177] = ~((layer2_outputs[1990]) | (layer2_outputs[4967]));
    assign layer3_outputs[178] = (layer2_outputs[1355]) | (layer2_outputs[4398]);
    assign layer3_outputs[179] = (layer2_outputs[1974]) & ~(layer2_outputs[3632]);
    assign layer3_outputs[180] = 1'b0;
    assign layer3_outputs[181] = ~((layer2_outputs[1805]) ^ (layer2_outputs[1109]));
    assign layer3_outputs[182] = ~((layer2_outputs[394]) | (layer2_outputs[1923]));
    assign layer3_outputs[183] = layer2_outputs[508];
    assign layer3_outputs[184] = layer2_outputs[4047];
    assign layer3_outputs[185] = 1'b1;
    assign layer3_outputs[186] = layer2_outputs[2297];
    assign layer3_outputs[187] = ~(layer2_outputs[291]) | (layer2_outputs[645]);
    assign layer3_outputs[188] = (layer2_outputs[1697]) & ~(layer2_outputs[933]);
    assign layer3_outputs[189] = ~(layer2_outputs[3472]);
    assign layer3_outputs[190] = 1'b0;
    assign layer3_outputs[191] = (layer2_outputs[630]) | (layer2_outputs[2340]);
    assign layer3_outputs[192] = (layer2_outputs[2694]) & ~(layer2_outputs[4612]);
    assign layer3_outputs[193] = ~((layer2_outputs[270]) | (layer2_outputs[3951]));
    assign layer3_outputs[194] = layer2_outputs[1764];
    assign layer3_outputs[195] = (layer2_outputs[3143]) & ~(layer2_outputs[2311]);
    assign layer3_outputs[196] = ~(layer2_outputs[4405]) | (layer2_outputs[4739]);
    assign layer3_outputs[197] = ~(layer2_outputs[4211]) | (layer2_outputs[4262]);
    assign layer3_outputs[198] = ~(layer2_outputs[1391]) | (layer2_outputs[3408]);
    assign layer3_outputs[199] = 1'b1;
    assign layer3_outputs[200] = 1'b0;
    assign layer3_outputs[201] = ~(layer2_outputs[3597]) | (layer2_outputs[3944]);
    assign layer3_outputs[202] = layer2_outputs[3497];
    assign layer3_outputs[203] = ~(layer2_outputs[3091]);
    assign layer3_outputs[204] = ~(layer2_outputs[622]) | (layer2_outputs[3851]);
    assign layer3_outputs[205] = ~(layer2_outputs[3952]);
    assign layer3_outputs[206] = ~(layer2_outputs[1441]);
    assign layer3_outputs[207] = ~(layer2_outputs[5089]) | (layer2_outputs[4320]);
    assign layer3_outputs[208] = (layer2_outputs[2942]) & ~(layer2_outputs[1919]);
    assign layer3_outputs[209] = ~((layer2_outputs[529]) & (layer2_outputs[4644]));
    assign layer3_outputs[210] = 1'b1;
    assign layer3_outputs[211] = ~((layer2_outputs[17]) | (layer2_outputs[4538]));
    assign layer3_outputs[212] = 1'b1;
    assign layer3_outputs[213] = 1'b1;
    assign layer3_outputs[214] = ~(layer2_outputs[4287]);
    assign layer3_outputs[215] = ~(layer2_outputs[3772]);
    assign layer3_outputs[216] = 1'b1;
    assign layer3_outputs[217] = ~((layer2_outputs[1202]) & (layer2_outputs[110]));
    assign layer3_outputs[218] = ~((layer2_outputs[2514]) & (layer2_outputs[983]));
    assign layer3_outputs[219] = ~(layer2_outputs[3252]) | (layer2_outputs[4669]);
    assign layer3_outputs[220] = layer2_outputs[2163];
    assign layer3_outputs[221] = ~(layer2_outputs[2519]);
    assign layer3_outputs[222] = ~((layer2_outputs[2608]) & (layer2_outputs[1783]));
    assign layer3_outputs[223] = layer2_outputs[2712];
    assign layer3_outputs[224] = ~(layer2_outputs[4953]);
    assign layer3_outputs[225] = 1'b1;
    assign layer3_outputs[226] = ~(layer2_outputs[514]) | (layer2_outputs[1148]);
    assign layer3_outputs[227] = ~(layer2_outputs[3708]) | (layer2_outputs[217]);
    assign layer3_outputs[228] = ~((layer2_outputs[1409]) ^ (layer2_outputs[3850]));
    assign layer3_outputs[229] = ~(layer2_outputs[2022]) | (layer2_outputs[1462]);
    assign layer3_outputs[230] = layer2_outputs[475];
    assign layer3_outputs[231] = (layer2_outputs[1682]) & ~(layer2_outputs[2161]);
    assign layer3_outputs[232] = (layer2_outputs[2811]) & ~(layer2_outputs[934]);
    assign layer3_outputs[233] = (layer2_outputs[2348]) | (layer2_outputs[5050]);
    assign layer3_outputs[234] = ~(layer2_outputs[223]) | (layer2_outputs[5036]);
    assign layer3_outputs[235] = ~(layer2_outputs[2307]);
    assign layer3_outputs[236] = ~((layer2_outputs[2575]) | (layer2_outputs[2469]));
    assign layer3_outputs[237] = layer2_outputs[4283];
    assign layer3_outputs[238] = layer2_outputs[3419];
    assign layer3_outputs[239] = ~(layer2_outputs[1861]) | (layer2_outputs[3190]);
    assign layer3_outputs[240] = ~((layer2_outputs[1081]) | (layer2_outputs[3288]));
    assign layer3_outputs[241] = ~((layer2_outputs[3710]) | (layer2_outputs[292]));
    assign layer3_outputs[242] = (layer2_outputs[776]) ^ (layer2_outputs[3055]);
    assign layer3_outputs[243] = (layer2_outputs[1437]) | (layer2_outputs[4752]);
    assign layer3_outputs[244] = layer2_outputs[2967];
    assign layer3_outputs[245] = ~(layer2_outputs[147]);
    assign layer3_outputs[246] = ~(layer2_outputs[4708]);
    assign layer3_outputs[247] = ~((layer2_outputs[2889]) & (layer2_outputs[2116]));
    assign layer3_outputs[248] = ~(layer2_outputs[66]);
    assign layer3_outputs[249] = layer2_outputs[3522];
    assign layer3_outputs[250] = ~((layer2_outputs[3094]) & (layer2_outputs[3657]));
    assign layer3_outputs[251] = (layer2_outputs[464]) ^ (layer2_outputs[1045]);
    assign layer3_outputs[252] = layer2_outputs[775];
    assign layer3_outputs[253] = ~(layer2_outputs[4369]) | (layer2_outputs[399]);
    assign layer3_outputs[254] = (layer2_outputs[1684]) ^ (layer2_outputs[3204]);
    assign layer3_outputs[255] = (layer2_outputs[1796]) ^ (layer2_outputs[745]);
    assign layer3_outputs[256] = ~((layer2_outputs[3543]) & (layer2_outputs[3213]));
    assign layer3_outputs[257] = 1'b0;
    assign layer3_outputs[258] = ~(layer2_outputs[5008]) | (layer2_outputs[4460]);
    assign layer3_outputs[259] = 1'b1;
    assign layer3_outputs[260] = ~(layer2_outputs[4924]) | (layer2_outputs[4157]);
    assign layer3_outputs[261] = (layer2_outputs[3365]) & ~(layer2_outputs[4321]);
    assign layer3_outputs[262] = (layer2_outputs[1184]) | (layer2_outputs[2894]);
    assign layer3_outputs[263] = layer2_outputs[2202];
    assign layer3_outputs[264] = ~((layer2_outputs[924]) | (layer2_outputs[97]));
    assign layer3_outputs[265] = layer2_outputs[4149];
    assign layer3_outputs[266] = (layer2_outputs[235]) | (layer2_outputs[1159]);
    assign layer3_outputs[267] = ~(layer2_outputs[783]);
    assign layer3_outputs[268] = ~(layer2_outputs[4345]) | (layer2_outputs[1851]);
    assign layer3_outputs[269] = (layer2_outputs[3801]) | (layer2_outputs[56]);
    assign layer3_outputs[270] = layer2_outputs[1719];
    assign layer3_outputs[271] = (layer2_outputs[2995]) & ~(layer2_outputs[5009]);
    assign layer3_outputs[272] = layer2_outputs[2442];
    assign layer3_outputs[273] = ~(layer2_outputs[838]);
    assign layer3_outputs[274] = ~(layer2_outputs[3743]) | (layer2_outputs[31]);
    assign layer3_outputs[275] = ~((layer2_outputs[3249]) & (layer2_outputs[3954]));
    assign layer3_outputs[276] = ~(layer2_outputs[4107]);
    assign layer3_outputs[277] = (layer2_outputs[3728]) & ~(layer2_outputs[254]);
    assign layer3_outputs[278] = ~(layer2_outputs[1030]);
    assign layer3_outputs[279] = ~((layer2_outputs[1304]) & (layer2_outputs[3649]));
    assign layer3_outputs[280] = layer2_outputs[506];
    assign layer3_outputs[281] = ~((layer2_outputs[4876]) ^ (layer2_outputs[4395]));
    assign layer3_outputs[282] = (layer2_outputs[3759]) & (layer2_outputs[2717]);
    assign layer3_outputs[283] = ~((layer2_outputs[379]) & (layer2_outputs[1712]));
    assign layer3_outputs[284] = 1'b1;
    assign layer3_outputs[285] = ~((layer2_outputs[2203]) ^ (layer2_outputs[2327]));
    assign layer3_outputs[286] = 1'b1;
    assign layer3_outputs[287] = layer2_outputs[1440];
    assign layer3_outputs[288] = ~((layer2_outputs[1226]) & (layer2_outputs[261]));
    assign layer3_outputs[289] = layer2_outputs[2425];
    assign layer3_outputs[290] = 1'b0;
    assign layer3_outputs[291] = 1'b1;
    assign layer3_outputs[292] = (layer2_outputs[715]) & ~(layer2_outputs[5058]);
    assign layer3_outputs[293] = ~(layer2_outputs[1414]);
    assign layer3_outputs[294] = (layer2_outputs[461]) & ~(layer2_outputs[2204]);
    assign layer3_outputs[295] = (layer2_outputs[2643]) | (layer2_outputs[2414]);
    assign layer3_outputs[296] = ~((layer2_outputs[1497]) & (layer2_outputs[328]));
    assign layer3_outputs[297] = (layer2_outputs[2559]) & ~(layer2_outputs[2214]);
    assign layer3_outputs[298] = layer2_outputs[2866];
    assign layer3_outputs[299] = 1'b1;
    assign layer3_outputs[300] = ~(layer2_outputs[4973]) | (layer2_outputs[2820]);
    assign layer3_outputs[301] = ~(layer2_outputs[4610]) | (layer2_outputs[1628]);
    assign layer3_outputs[302] = 1'b1;
    assign layer3_outputs[303] = (layer2_outputs[1736]) | (layer2_outputs[3730]);
    assign layer3_outputs[304] = (layer2_outputs[4812]) | (layer2_outputs[4593]);
    assign layer3_outputs[305] = (layer2_outputs[1557]) & (layer2_outputs[3440]);
    assign layer3_outputs[306] = layer2_outputs[4698];
    assign layer3_outputs[307] = ~(layer2_outputs[5079]);
    assign layer3_outputs[308] = (layer2_outputs[2036]) & (layer2_outputs[4581]);
    assign layer3_outputs[309] = ~((layer2_outputs[611]) & (layer2_outputs[2224]));
    assign layer3_outputs[310] = (layer2_outputs[5074]) & ~(layer2_outputs[3940]);
    assign layer3_outputs[311] = 1'b0;
    assign layer3_outputs[312] = ~(layer2_outputs[4838]);
    assign layer3_outputs[313] = ~(layer2_outputs[3849]);
    assign layer3_outputs[314] = ~(layer2_outputs[2106]);
    assign layer3_outputs[315] = ~((layer2_outputs[2074]) & (layer2_outputs[897]));
    assign layer3_outputs[316] = (layer2_outputs[3862]) ^ (layer2_outputs[1586]);
    assign layer3_outputs[317] = layer2_outputs[2152];
    assign layer3_outputs[318] = (layer2_outputs[1730]) | (layer2_outputs[460]);
    assign layer3_outputs[319] = ~((layer2_outputs[1192]) ^ (layer2_outputs[3275]));
    assign layer3_outputs[320] = (layer2_outputs[1153]) | (layer2_outputs[5003]);
    assign layer3_outputs[321] = (layer2_outputs[3355]) & (layer2_outputs[1368]);
    assign layer3_outputs[322] = (layer2_outputs[2579]) & ~(layer2_outputs[460]);
    assign layer3_outputs[323] = layer2_outputs[181];
    assign layer3_outputs[324] = ~(layer2_outputs[2703]);
    assign layer3_outputs[325] = (layer2_outputs[1326]) & ~(layer2_outputs[4036]);
    assign layer3_outputs[326] = 1'b1;
    assign layer3_outputs[327] = layer2_outputs[1163];
    assign layer3_outputs[328] = layer2_outputs[4405];
    assign layer3_outputs[329] = 1'b1;
    assign layer3_outputs[330] = ~(layer2_outputs[949]);
    assign layer3_outputs[331] = ~(layer2_outputs[2837]) | (layer2_outputs[159]);
    assign layer3_outputs[332] = layer2_outputs[2966];
    assign layer3_outputs[333] = (layer2_outputs[4522]) | (layer2_outputs[726]);
    assign layer3_outputs[334] = ~(layer2_outputs[150]);
    assign layer3_outputs[335] = ~(layer2_outputs[4122]) | (layer2_outputs[4980]);
    assign layer3_outputs[336] = ~(layer2_outputs[4437]) | (layer2_outputs[2749]);
    assign layer3_outputs[337] = ~((layer2_outputs[3905]) & (layer2_outputs[2502]));
    assign layer3_outputs[338] = ~(layer2_outputs[1743]);
    assign layer3_outputs[339] = ~(layer2_outputs[4076]);
    assign layer3_outputs[340] = ~(layer2_outputs[1112]);
    assign layer3_outputs[341] = 1'b0;
    assign layer3_outputs[342] = (layer2_outputs[551]) & ~(layer2_outputs[3352]);
    assign layer3_outputs[343] = ~(layer2_outputs[1680]);
    assign layer3_outputs[344] = (layer2_outputs[3399]) & ~(layer2_outputs[3262]);
    assign layer3_outputs[345] = ~(layer2_outputs[3208]) | (layer2_outputs[2743]);
    assign layer3_outputs[346] = ~(layer2_outputs[2547]);
    assign layer3_outputs[347] = 1'b0;
    assign layer3_outputs[348] = 1'b0;
    assign layer3_outputs[349] = (layer2_outputs[2228]) & ~(layer2_outputs[4864]);
    assign layer3_outputs[350] = layer2_outputs[1082];
    assign layer3_outputs[351] = (layer2_outputs[403]) & ~(layer2_outputs[1636]);
    assign layer3_outputs[352] = ~(layer2_outputs[3003]) | (layer2_outputs[956]);
    assign layer3_outputs[353] = ~((layer2_outputs[360]) & (layer2_outputs[3398]));
    assign layer3_outputs[354] = ~(layer2_outputs[1075]) | (layer2_outputs[3007]);
    assign layer3_outputs[355] = ~(layer2_outputs[475]);
    assign layer3_outputs[356] = (layer2_outputs[2739]) & ~(layer2_outputs[2965]);
    assign layer3_outputs[357] = ~(layer2_outputs[647]);
    assign layer3_outputs[358] = 1'b1;
    assign layer3_outputs[359] = ~(layer2_outputs[648]);
    assign layer3_outputs[360] = 1'b0;
    assign layer3_outputs[361] = ~(layer2_outputs[819]);
    assign layer3_outputs[362] = layer2_outputs[2463];
    assign layer3_outputs[363] = ~(layer2_outputs[4054]) | (layer2_outputs[4228]);
    assign layer3_outputs[364] = layer2_outputs[2124];
    assign layer3_outputs[365] = ~((layer2_outputs[4168]) | (layer2_outputs[4952]));
    assign layer3_outputs[366] = 1'b0;
    assign layer3_outputs[367] = ~(layer2_outputs[1384]) | (layer2_outputs[1673]);
    assign layer3_outputs[368] = ~(layer2_outputs[4940]);
    assign layer3_outputs[369] = 1'b0;
    assign layer3_outputs[370] = 1'b1;
    assign layer3_outputs[371] = (layer2_outputs[1872]) | (layer2_outputs[2915]);
    assign layer3_outputs[372] = ~(layer2_outputs[735]) | (layer2_outputs[696]);
    assign layer3_outputs[373] = (layer2_outputs[2778]) & ~(layer2_outputs[2894]);
    assign layer3_outputs[374] = ~(layer2_outputs[1528]);
    assign layer3_outputs[375] = (layer2_outputs[1925]) | (layer2_outputs[2861]);
    assign layer3_outputs[376] = 1'b0;
    assign layer3_outputs[377] = ~((layer2_outputs[3458]) & (layer2_outputs[415]));
    assign layer3_outputs[378] = (layer2_outputs[3794]) & (layer2_outputs[2508]);
    assign layer3_outputs[379] = ~(layer2_outputs[1385]);
    assign layer3_outputs[380] = 1'b0;
    assign layer3_outputs[381] = layer2_outputs[143];
    assign layer3_outputs[382] = layer2_outputs[955];
    assign layer3_outputs[383] = ~((layer2_outputs[1672]) | (layer2_outputs[669]));
    assign layer3_outputs[384] = (layer2_outputs[605]) & (layer2_outputs[1253]);
    assign layer3_outputs[385] = layer2_outputs[2156];
    assign layer3_outputs[386] = ~((layer2_outputs[1138]) | (layer2_outputs[1418]));
    assign layer3_outputs[387] = ~((layer2_outputs[3552]) & (layer2_outputs[2766]));
    assign layer3_outputs[388] = ~(layer2_outputs[1747]) | (layer2_outputs[3799]);
    assign layer3_outputs[389] = (layer2_outputs[4095]) | (layer2_outputs[1403]);
    assign layer3_outputs[390] = ~(layer2_outputs[2172]);
    assign layer3_outputs[391] = ~(layer2_outputs[1173]);
    assign layer3_outputs[392] = ~(layer2_outputs[1253]) | (layer2_outputs[3871]);
    assign layer3_outputs[393] = (layer2_outputs[1633]) | (layer2_outputs[995]);
    assign layer3_outputs[394] = ~((layer2_outputs[3718]) | (layer2_outputs[1017]));
    assign layer3_outputs[395] = ~(layer2_outputs[1657]) | (layer2_outputs[1344]);
    assign layer3_outputs[396] = (layer2_outputs[4213]) & (layer2_outputs[3722]);
    assign layer3_outputs[397] = (layer2_outputs[3432]) & ~(layer2_outputs[3251]);
    assign layer3_outputs[398] = layer2_outputs[1740];
    assign layer3_outputs[399] = ~(layer2_outputs[2241]);
    assign layer3_outputs[400] = 1'b1;
    assign layer3_outputs[401] = 1'b0;
    assign layer3_outputs[402] = (layer2_outputs[715]) & ~(layer2_outputs[1284]);
    assign layer3_outputs[403] = layer2_outputs[2799];
    assign layer3_outputs[404] = (layer2_outputs[1522]) & (layer2_outputs[3443]);
    assign layer3_outputs[405] = ~(layer2_outputs[2891]);
    assign layer3_outputs[406] = (layer2_outputs[4274]) ^ (layer2_outputs[4489]);
    assign layer3_outputs[407] = ~(layer2_outputs[1583]);
    assign layer3_outputs[408] = layer2_outputs[2284];
    assign layer3_outputs[409] = 1'b0;
    assign layer3_outputs[410] = layer2_outputs[2494];
    assign layer3_outputs[411] = layer2_outputs[3402];
    assign layer3_outputs[412] = ~((layer2_outputs[918]) | (layer2_outputs[2603]));
    assign layer3_outputs[413] = (layer2_outputs[2231]) & ~(layer2_outputs[2496]);
    assign layer3_outputs[414] = ~(layer2_outputs[4329]);
    assign layer3_outputs[415] = ~((layer2_outputs[1630]) & (layer2_outputs[2515]));
    assign layer3_outputs[416] = layer2_outputs[3137];
    assign layer3_outputs[417] = (layer2_outputs[1501]) & ~(layer2_outputs[1136]);
    assign layer3_outputs[418] = (layer2_outputs[3912]) & ~(layer2_outputs[2665]);
    assign layer3_outputs[419] = layer2_outputs[3152];
    assign layer3_outputs[420] = ~(layer2_outputs[4950]);
    assign layer3_outputs[421] = (layer2_outputs[2590]) & ~(layer2_outputs[2562]);
    assign layer3_outputs[422] = (layer2_outputs[80]) & ~(layer2_outputs[942]);
    assign layer3_outputs[423] = layer2_outputs[3450];
    assign layer3_outputs[424] = (layer2_outputs[474]) | (layer2_outputs[3387]);
    assign layer3_outputs[425] = ~(layer2_outputs[233]);
    assign layer3_outputs[426] = (layer2_outputs[4711]) ^ (layer2_outputs[3054]);
    assign layer3_outputs[427] = ~(layer2_outputs[4830]);
    assign layer3_outputs[428] = ~(layer2_outputs[442]);
    assign layer3_outputs[429] = ~((layer2_outputs[2696]) ^ (layer2_outputs[1938]));
    assign layer3_outputs[430] = ~(layer2_outputs[4216]);
    assign layer3_outputs[431] = (layer2_outputs[4843]) & ~(layer2_outputs[2401]);
    assign layer3_outputs[432] = (layer2_outputs[1322]) | (layer2_outputs[561]);
    assign layer3_outputs[433] = ~(layer2_outputs[2938]);
    assign layer3_outputs[434] = (layer2_outputs[4206]) | (layer2_outputs[1010]);
    assign layer3_outputs[435] = 1'b1;
    assign layer3_outputs[436] = (layer2_outputs[1242]) | (layer2_outputs[1271]);
    assign layer3_outputs[437] = layer2_outputs[3704];
    assign layer3_outputs[438] = ~((layer2_outputs[2926]) | (layer2_outputs[3690]));
    assign layer3_outputs[439] = layer2_outputs[1319];
    assign layer3_outputs[440] = 1'b0;
    assign layer3_outputs[441] = (layer2_outputs[327]) & ~(layer2_outputs[1434]);
    assign layer3_outputs[442] = layer2_outputs[4748];
    assign layer3_outputs[443] = (layer2_outputs[927]) | (layer2_outputs[3731]);
    assign layer3_outputs[444] = layer2_outputs[3633];
    assign layer3_outputs[445] = 1'b1;
    assign layer3_outputs[446] = layer2_outputs[2674];
    assign layer3_outputs[447] = layer2_outputs[347];
    assign layer3_outputs[448] = (layer2_outputs[504]) | (layer2_outputs[4369]);
    assign layer3_outputs[449] = (layer2_outputs[4719]) & (layer2_outputs[2542]);
    assign layer3_outputs[450] = ~(layer2_outputs[333]);
    assign layer3_outputs[451] = ~((layer2_outputs[40]) | (layer2_outputs[2702]));
    assign layer3_outputs[452] = (layer2_outputs[2974]) & ~(layer2_outputs[5107]);
    assign layer3_outputs[453] = (layer2_outputs[4756]) | (layer2_outputs[2749]);
    assign layer3_outputs[454] = ~(layer2_outputs[2247]) | (layer2_outputs[1394]);
    assign layer3_outputs[455] = (layer2_outputs[1321]) & (layer2_outputs[4887]);
    assign layer3_outputs[456] = layer2_outputs[3524];
    assign layer3_outputs[457] = 1'b1;
    assign layer3_outputs[458] = layer2_outputs[3047];
    assign layer3_outputs[459] = 1'b1;
    assign layer3_outputs[460] = (layer2_outputs[3621]) & ~(layer2_outputs[3703]);
    assign layer3_outputs[461] = ~(layer2_outputs[932]);
    assign layer3_outputs[462] = 1'b0;
    assign layer3_outputs[463] = ~((layer2_outputs[2447]) | (layer2_outputs[3135]));
    assign layer3_outputs[464] = (layer2_outputs[388]) & ~(layer2_outputs[2454]);
    assign layer3_outputs[465] = (layer2_outputs[37]) & ~(layer2_outputs[2336]);
    assign layer3_outputs[466] = layer2_outputs[1131];
    assign layer3_outputs[467] = ~((layer2_outputs[4004]) & (layer2_outputs[4845]));
    assign layer3_outputs[468] = ~(layer2_outputs[4001]);
    assign layer3_outputs[469] = 1'b1;
    assign layer3_outputs[470] = ~(layer2_outputs[3290]);
    assign layer3_outputs[471] = (layer2_outputs[29]) | (layer2_outputs[568]);
    assign layer3_outputs[472] = (layer2_outputs[837]) ^ (layer2_outputs[856]);
    assign layer3_outputs[473] = layer2_outputs[5111];
    assign layer3_outputs[474] = (layer2_outputs[1290]) & ~(layer2_outputs[516]);
    assign layer3_outputs[475] = ~(layer2_outputs[180]) | (layer2_outputs[3109]);
    assign layer3_outputs[476] = ~(layer2_outputs[909]);
    assign layer3_outputs[477] = 1'b0;
    assign layer3_outputs[478] = ~(layer2_outputs[4930]);
    assign layer3_outputs[479] = ~(layer2_outputs[1011]);
    assign layer3_outputs[480] = ~(layer2_outputs[3657]) | (layer2_outputs[1849]);
    assign layer3_outputs[481] = 1'b1;
    assign layer3_outputs[482] = layer2_outputs[1753];
    assign layer3_outputs[483] = 1'b0;
    assign layer3_outputs[484] = ~(layer2_outputs[1692]);
    assign layer3_outputs[485] = layer2_outputs[4767];
    assign layer3_outputs[486] = ~(layer2_outputs[463]) | (layer2_outputs[3755]);
    assign layer3_outputs[487] = (layer2_outputs[4918]) & ~(layer2_outputs[4640]);
    assign layer3_outputs[488] = 1'b0;
    assign layer3_outputs[489] = ~((layer2_outputs[4197]) & (layer2_outputs[324]));
    assign layer3_outputs[490] = ~((layer2_outputs[2520]) | (layer2_outputs[796]));
    assign layer3_outputs[491] = (layer2_outputs[434]) & (layer2_outputs[3092]);
    assign layer3_outputs[492] = 1'b1;
    assign layer3_outputs[493] = (layer2_outputs[3176]) & (layer2_outputs[3552]);
    assign layer3_outputs[494] = layer2_outputs[2987];
    assign layer3_outputs[495] = ~((layer2_outputs[12]) | (layer2_outputs[3917]));
    assign layer3_outputs[496] = layer2_outputs[2677];
    assign layer3_outputs[497] = (layer2_outputs[1302]) & (layer2_outputs[2167]);
    assign layer3_outputs[498] = layer2_outputs[1656];
    assign layer3_outputs[499] = ~(layer2_outputs[4965]);
    assign layer3_outputs[500] = 1'b1;
    assign layer3_outputs[501] = 1'b0;
    assign layer3_outputs[502] = ~((layer2_outputs[1903]) | (layer2_outputs[3294]));
    assign layer3_outputs[503] = (layer2_outputs[4654]) ^ (layer2_outputs[1346]);
    assign layer3_outputs[504] = layer2_outputs[1655];
    assign layer3_outputs[505] = layer2_outputs[873];
    assign layer3_outputs[506] = ~((layer2_outputs[2500]) | (layer2_outputs[682]));
    assign layer3_outputs[507] = ~(layer2_outputs[2181]);
    assign layer3_outputs[508] = ~(layer2_outputs[3141]);
    assign layer3_outputs[509] = layer2_outputs[4890];
    assign layer3_outputs[510] = ~((layer2_outputs[3226]) & (layer2_outputs[661]));
    assign layer3_outputs[511] = ~((layer2_outputs[2789]) | (layer2_outputs[3423]));
    assign layer3_outputs[512] = layer2_outputs[4167];
    assign layer3_outputs[513] = layer2_outputs[4463];
    assign layer3_outputs[514] = 1'b0;
    assign layer3_outputs[515] = (layer2_outputs[4855]) & ~(layer2_outputs[4718]);
    assign layer3_outputs[516] = layer2_outputs[3681];
    assign layer3_outputs[517] = layer2_outputs[3661];
    assign layer3_outputs[518] = (layer2_outputs[1163]) & ~(layer2_outputs[2731]);
    assign layer3_outputs[519] = (layer2_outputs[2103]) & (layer2_outputs[3145]);
    assign layer3_outputs[520] = ~(layer2_outputs[1117]) | (layer2_outputs[3891]);
    assign layer3_outputs[521] = layer2_outputs[5010];
    assign layer3_outputs[522] = ~(layer2_outputs[3342]) | (layer2_outputs[4199]);
    assign layer3_outputs[523] = 1'b0;
    assign layer3_outputs[524] = (layer2_outputs[676]) | (layer2_outputs[4079]);
    assign layer3_outputs[525] = layer2_outputs[4905];
    assign layer3_outputs[526] = 1'b1;
    assign layer3_outputs[527] = ~((layer2_outputs[672]) & (layer2_outputs[4526]));
    assign layer3_outputs[528] = (layer2_outputs[2939]) ^ (layer2_outputs[4845]);
    assign layer3_outputs[529] = ~((layer2_outputs[3332]) | (layer2_outputs[976]));
    assign layer3_outputs[530] = layer2_outputs[4404];
    assign layer3_outputs[531] = (layer2_outputs[4341]) & ~(layer2_outputs[2638]);
    assign layer3_outputs[532] = ~((layer2_outputs[3197]) | (layer2_outputs[329]));
    assign layer3_outputs[533] = ~(layer2_outputs[2275]) | (layer2_outputs[2890]);
    assign layer3_outputs[534] = (layer2_outputs[2611]) & ~(layer2_outputs[1758]);
    assign layer3_outputs[535] = layer2_outputs[4895];
    assign layer3_outputs[536] = layer2_outputs[4249];
    assign layer3_outputs[537] = ~(layer2_outputs[3525]) | (layer2_outputs[129]);
    assign layer3_outputs[538] = layer2_outputs[1119];
    assign layer3_outputs[539] = layer2_outputs[4357];
    assign layer3_outputs[540] = 1'b0;
    assign layer3_outputs[541] = ~((layer2_outputs[1691]) | (layer2_outputs[922]));
    assign layer3_outputs[542] = ~(layer2_outputs[4477]) | (layer2_outputs[707]);
    assign layer3_outputs[543] = (layer2_outputs[2343]) & (layer2_outputs[741]);
    assign layer3_outputs[544] = layer2_outputs[4497];
    assign layer3_outputs[545] = ~((layer2_outputs[1853]) | (layer2_outputs[1446]));
    assign layer3_outputs[546] = (layer2_outputs[3133]) | (layer2_outputs[4974]);
    assign layer3_outputs[547] = ~((layer2_outputs[930]) & (layer2_outputs[859]));
    assign layer3_outputs[548] = layer2_outputs[4927];
    assign layer3_outputs[549] = ~(layer2_outputs[1353]) | (layer2_outputs[5047]);
    assign layer3_outputs[550] = 1'b0;
    assign layer3_outputs[551] = ~(layer2_outputs[1316]) | (layer2_outputs[1537]);
    assign layer3_outputs[552] = ~((layer2_outputs[502]) | (layer2_outputs[3110]));
    assign layer3_outputs[553] = layer2_outputs[4086];
    assign layer3_outputs[554] = (layer2_outputs[2754]) & ~(layer2_outputs[1615]);
    assign layer3_outputs[555] = ~((layer2_outputs[2254]) | (layer2_outputs[955]));
    assign layer3_outputs[556] = (layer2_outputs[30]) & ~(layer2_outputs[677]);
    assign layer3_outputs[557] = layer2_outputs[3507];
    assign layer3_outputs[558] = ~(layer2_outputs[3293]) | (layer2_outputs[1899]);
    assign layer3_outputs[559] = ~(layer2_outputs[4319]);
    assign layer3_outputs[560] = ~(layer2_outputs[4787]) | (layer2_outputs[1272]);
    assign layer3_outputs[561] = 1'b0;
    assign layer3_outputs[562] = ~((layer2_outputs[1254]) & (layer2_outputs[3754]));
    assign layer3_outputs[563] = 1'b0;
    assign layer3_outputs[564] = (layer2_outputs[4328]) & ~(layer2_outputs[1404]);
    assign layer3_outputs[565] = (layer2_outputs[1827]) & (layer2_outputs[3336]);
    assign layer3_outputs[566] = ~((layer2_outputs[4585]) ^ (layer2_outputs[2079]));
    assign layer3_outputs[567] = (layer2_outputs[5057]) & ~(layer2_outputs[2265]);
    assign layer3_outputs[568] = layer2_outputs[2208];
    assign layer3_outputs[569] = 1'b1;
    assign layer3_outputs[570] = ~(layer2_outputs[1614]);
    assign layer3_outputs[571] = 1'b0;
    assign layer3_outputs[572] = (layer2_outputs[4294]) ^ (layer2_outputs[1084]);
    assign layer3_outputs[573] = layer2_outputs[2716];
    assign layer3_outputs[574] = (layer2_outputs[4559]) & (layer2_outputs[42]);
    assign layer3_outputs[575] = ~(layer2_outputs[3638]);
    assign layer3_outputs[576] = 1'b0;
    assign layer3_outputs[577] = ~(layer2_outputs[181]);
    assign layer3_outputs[578] = ~(layer2_outputs[3433]);
    assign layer3_outputs[579] = (layer2_outputs[1205]) & (layer2_outputs[2420]);
    assign layer3_outputs[580] = layer2_outputs[1332];
    assign layer3_outputs[581] = (layer2_outputs[2525]) & ~(layer2_outputs[763]);
    assign layer3_outputs[582] = (layer2_outputs[2505]) & ~(layer2_outputs[3437]);
    assign layer3_outputs[583] = ~(layer2_outputs[620]);
    assign layer3_outputs[584] = ~((layer2_outputs[1926]) & (layer2_outputs[2138]));
    assign layer3_outputs[585] = ~((layer2_outputs[3764]) ^ (layer2_outputs[4390]));
    assign layer3_outputs[586] = layer2_outputs[1969];
    assign layer3_outputs[587] = ~(layer2_outputs[4045]);
    assign layer3_outputs[588] = ~(layer2_outputs[1224]);
    assign layer3_outputs[589] = 1'b0;
    assign layer3_outputs[590] = ~((layer2_outputs[448]) | (layer2_outputs[3537]));
    assign layer3_outputs[591] = (layer2_outputs[1897]) & ~(layer2_outputs[1170]);
    assign layer3_outputs[592] = (layer2_outputs[28]) | (layer2_outputs[760]);
    assign layer3_outputs[593] = (layer2_outputs[437]) & ~(layer2_outputs[351]);
    assign layer3_outputs[594] = (layer2_outputs[1352]) & ~(layer2_outputs[3395]);
    assign layer3_outputs[595] = ~((layer2_outputs[5017]) & (layer2_outputs[3511]));
    assign layer3_outputs[596] = ~(layer2_outputs[3999]) | (layer2_outputs[2558]);
    assign layer3_outputs[597] = (layer2_outputs[4439]) | (layer2_outputs[3738]);
    assign layer3_outputs[598] = ~((layer2_outputs[1398]) ^ (layer2_outputs[998]));
    assign layer3_outputs[599] = (layer2_outputs[3766]) | (layer2_outputs[4154]);
    assign layer3_outputs[600] = 1'b1;
    assign layer3_outputs[601] = ~((layer2_outputs[878]) | (layer2_outputs[974]));
    assign layer3_outputs[602] = ~(layer2_outputs[2755]);
    assign layer3_outputs[603] = ~((layer2_outputs[1161]) & (layer2_outputs[367]));
    assign layer3_outputs[604] = layer2_outputs[4594];
    assign layer3_outputs[605] = ~(layer2_outputs[4346]) | (layer2_outputs[1864]);
    assign layer3_outputs[606] = layer2_outputs[4148];
    assign layer3_outputs[607] = ~(layer2_outputs[2737]);
    assign layer3_outputs[608] = layer2_outputs[5006];
    assign layer3_outputs[609] = (layer2_outputs[5040]) | (layer2_outputs[1799]);
    assign layer3_outputs[610] = (layer2_outputs[3826]) & ~(layer2_outputs[4416]);
    assign layer3_outputs[611] = 1'b1;
    assign layer3_outputs[612] = ~(layer2_outputs[790]) | (layer2_outputs[1929]);
    assign layer3_outputs[613] = layer2_outputs[2693];
    assign layer3_outputs[614] = (layer2_outputs[4976]) & (layer2_outputs[824]);
    assign layer3_outputs[615] = ~(layer2_outputs[698]) | (layer2_outputs[3592]);
    assign layer3_outputs[616] = layer2_outputs[2153];
    assign layer3_outputs[617] = ~((layer2_outputs[2402]) & (layer2_outputs[1387]));
    assign layer3_outputs[618] = ~((layer2_outputs[4266]) ^ (layer2_outputs[1073]));
    assign layer3_outputs[619] = (layer2_outputs[2769]) & ~(layer2_outputs[395]);
    assign layer3_outputs[620] = ~((layer2_outputs[4190]) | (layer2_outputs[1295]));
    assign layer3_outputs[621] = (layer2_outputs[536]) & (layer2_outputs[2299]);
    assign layer3_outputs[622] = (layer2_outputs[5029]) ^ (layer2_outputs[1285]);
    assign layer3_outputs[623] = ~((layer2_outputs[2128]) & (layer2_outputs[2864]));
    assign layer3_outputs[624] = ~(layer2_outputs[1495]) | (layer2_outputs[4012]);
    assign layer3_outputs[625] = ~(layer2_outputs[5048]);
    assign layer3_outputs[626] = ~((layer2_outputs[2855]) & (layer2_outputs[2787]));
    assign layer3_outputs[627] = ~(layer2_outputs[4288]);
    assign layer3_outputs[628] = ~((layer2_outputs[4374]) & (layer2_outputs[4354]));
    assign layer3_outputs[629] = ~(layer2_outputs[5084]);
    assign layer3_outputs[630] = ~((layer2_outputs[65]) | (layer2_outputs[630]));
    assign layer3_outputs[631] = ~(layer2_outputs[3947]) | (layer2_outputs[991]);
    assign layer3_outputs[632] = layer2_outputs[1449];
    assign layer3_outputs[633] = (layer2_outputs[3840]) & ~(layer2_outputs[2654]);
    assign layer3_outputs[634] = (layer2_outputs[1642]) | (layer2_outputs[4304]);
    assign layer3_outputs[635] = 1'b0;
    assign layer3_outputs[636] = ~(layer2_outputs[1823]);
    assign layer3_outputs[637] = ~(layer2_outputs[2471]);
    assign layer3_outputs[638] = (layer2_outputs[1913]) & (layer2_outputs[797]);
    assign layer3_outputs[639] = (layer2_outputs[4285]) & (layer2_outputs[1729]);
    assign layer3_outputs[640] = (layer2_outputs[180]) & ~(layer2_outputs[332]);
    assign layer3_outputs[641] = (layer2_outputs[1700]) | (layer2_outputs[2856]);
    assign layer3_outputs[642] = ~((layer2_outputs[3732]) | (layer2_outputs[1208]));
    assign layer3_outputs[643] = layer2_outputs[3947];
    assign layer3_outputs[644] = layer2_outputs[5027];
    assign layer3_outputs[645] = 1'b0;
    assign layer3_outputs[646] = ~((layer2_outputs[4030]) & (layer2_outputs[844]));
    assign layer3_outputs[647] = (layer2_outputs[3256]) & ~(layer2_outputs[2956]);
    assign layer3_outputs[648] = 1'b1;
    assign layer3_outputs[649] = (layer2_outputs[1203]) & (layer2_outputs[967]);
    assign layer3_outputs[650] = (layer2_outputs[664]) & (layer2_outputs[3301]);
    assign layer3_outputs[651] = ~((layer2_outputs[4699]) | (layer2_outputs[3918]));
    assign layer3_outputs[652] = ~(layer2_outputs[4826]);
    assign layer3_outputs[653] = layer2_outputs[2979];
    assign layer3_outputs[654] = (layer2_outputs[1349]) & (layer2_outputs[3848]);
    assign layer3_outputs[655] = (layer2_outputs[3625]) & ~(layer2_outputs[748]);
    assign layer3_outputs[656] = ~((layer2_outputs[2950]) & (layer2_outputs[2422]));
    assign layer3_outputs[657] = layer2_outputs[2935];
    assign layer3_outputs[658] = ~((layer2_outputs[5117]) | (layer2_outputs[395]));
    assign layer3_outputs[659] = ~(layer2_outputs[98]);
    assign layer3_outputs[660] = layer2_outputs[1744];
    assign layer3_outputs[661] = layer2_outputs[3832];
    assign layer3_outputs[662] = ~((layer2_outputs[3641]) ^ (layer2_outputs[2985]));
    assign layer3_outputs[663] = ~((layer2_outputs[3388]) ^ (layer2_outputs[3233]));
    assign layer3_outputs[664] = layer2_outputs[3363];
    assign layer3_outputs[665] = 1'b0;
    assign layer3_outputs[666] = ~(layer2_outputs[4049]) | (layer2_outputs[245]);
    assign layer3_outputs[667] = ~((layer2_outputs[3238]) & (layer2_outputs[2506]));
    assign layer3_outputs[668] = ~(layer2_outputs[2436]);
    assign layer3_outputs[669] = (layer2_outputs[342]) & (layer2_outputs[2341]);
    assign layer3_outputs[670] = (layer2_outputs[1234]) & ~(layer2_outputs[3248]);
    assign layer3_outputs[671] = ~((layer2_outputs[555]) | (layer2_outputs[2129]));
    assign layer3_outputs[672] = ~(layer2_outputs[3688]);
    assign layer3_outputs[673] = ~(layer2_outputs[3083]);
    assign layer3_outputs[674] = 1'b0;
    assign layer3_outputs[675] = ~(layer2_outputs[3298]);
    assign layer3_outputs[676] = 1'b0;
    assign layer3_outputs[677] = layer2_outputs[4407];
    assign layer3_outputs[678] = ~(layer2_outputs[1300]);
    assign layer3_outputs[679] = layer2_outputs[3784];
    assign layer3_outputs[680] = (layer2_outputs[4130]) & (layer2_outputs[4217]);
    assign layer3_outputs[681] = ~((layer2_outputs[5065]) & (layer2_outputs[975]));
    assign layer3_outputs[682] = ~(layer2_outputs[3191]);
    assign layer3_outputs[683] = ~(layer2_outputs[5095]);
    assign layer3_outputs[684] = ~(layer2_outputs[310]) | (layer2_outputs[4324]);
    assign layer3_outputs[685] = layer2_outputs[2306];
    assign layer3_outputs[686] = layer2_outputs[2084];
    assign layer3_outputs[687] = layer2_outputs[3824];
    assign layer3_outputs[688] = ~(layer2_outputs[759]);
    assign layer3_outputs[689] = ~(layer2_outputs[623]);
    assign layer3_outputs[690] = layer2_outputs[1611];
    assign layer3_outputs[691] = (layer2_outputs[3827]) & ~(layer2_outputs[3931]);
    assign layer3_outputs[692] = 1'b1;
    assign layer3_outputs[693] = ~((layer2_outputs[3941]) & (layer2_outputs[2377]));
    assign layer3_outputs[694] = ~(layer2_outputs[1464]);
    assign layer3_outputs[695] = ~(layer2_outputs[338]) | (layer2_outputs[2261]);
    assign layer3_outputs[696] = ~((layer2_outputs[888]) | (layer2_outputs[2592]));
    assign layer3_outputs[697] = ~(layer2_outputs[2895]);
    assign layer3_outputs[698] = (layer2_outputs[2243]) ^ (layer2_outputs[131]);
    assign layer3_outputs[699] = layer2_outputs[3836];
    assign layer3_outputs[700] = 1'b1;
    assign layer3_outputs[701] = ~(layer2_outputs[212]);
    assign layer3_outputs[702] = ~(layer2_outputs[3298]) | (layer2_outputs[3591]);
    assign layer3_outputs[703] = ~((layer2_outputs[2063]) & (layer2_outputs[4339]));
    assign layer3_outputs[704] = (layer2_outputs[3404]) & ~(layer2_outputs[513]);
    assign layer3_outputs[705] = (layer2_outputs[628]) | (layer2_outputs[420]);
    assign layer3_outputs[706] = (layer2_outputs[2376]) & ~(layer2_outputs[3169]);
    assign layer3_outputs[707] = (layer2_outputs[3861]) & (layer2_outputs[1967]);
    assign layer3_outputs[708] = layer2_outputs[2682];
    assign layer3_outputs[709] = 1'b1;
    assign layer3_outputs[710] = ~(layer2_outputs[30]);
    assign layer3_outputs[711] = ~((layer2_outputs[2301]) & (layer2_outputs[2406]));
    assign layer3_outputs[712] = ~((layer2_outputs[2835]) ^ (layer2_outputs[1859]));
    assign layer3_outputs[713] = 1'b1;
    assign layer3_outputs[714] = ~((layer2_outputs[4447]) | (layer2_outputs[210]));
    assign layer3_outputs[715] = (layer2_outputs[761]) & (layer2_outputs[5041]);
    assign layer3_outputs[716] = ~(layer2_outputs[4082]) | (layer2_outputs[1058]);
    assign layer3_outputs[717] = layer2_outputs[842];
    assign layer3_outputs[718] = ~(layer2_outputs[2824]) | (layer2_outputs[330]);
    assign layer3_outputs[719] = (layer2_outputs[1568]) & (layer2_outputs[2456]);
    assign layer3_outputs[720] = 1'b1;
    assign layer3_outputs[721] = layer2_outputs[4583];
    assign layer3_outputs[722] = ~(layer2_outputs[4998]) | (layer2_outputs[1781]);
    assign layer3_outputs[723] = 1'b0;
    assign layer3_outputs[724] = (layer2_outputs[3925]) & (layer2_outputs[2239]);
    assign layer3_outputs[725] = (layer2_outputs[485]) & ~(layer2_outputs[2989]);
    assign layer3_outputs[726] = 1'b1;
    assign layer3_outputs[727] = (layer2_outputs[2507]) & ~(layer2_outputs[894]);
    assign layer3_outputs[728] = (layer2_outputs[804]) | (layer2_outputs[2928]);
    assign layer3_outputs[729] = layer2_outputs[1908];
    assign layer3_outputs[730] = ~(layer2_outputs[3155]) | (layer2_outputs[4963]);
    assign layer3_outputs[731] = 1'b1;
    assign layer3_outputs[732] = layer2_outputs[4708];
    assign layer3_outputs[733] = ~(layer2_outputs[1293]);
    assign layer3_outputs[734] = ~(layer2_outputs[3328]);
    assign layer3_outputs[735] = 1'b1;
    assign layer3_outputs[736] = 1'b1;
    assign layer3_outputs[737] = layer2_outputs[2381];
    assign layer3_outputs[738] = 1'b0;
    assign layer3_outputs[739] = (layer2_outputs[4216]) & ~(layer2_outputs[1034]);
    assign layer3_outputs[740] = ~(layer2_outputs[4425]);
    assign layer3_outputs[741] = layer2_outputs[4706];
    assign layer3_outputs[742] = (layer2_outputs[1818]) & (layer2_outputs[4859]);
    assign layer3_outputs[743] = layer2_outputs[432];
    assign layer3_outputs[744] = (layer2_outputs[3793]) & (layer2_outputs[1848]);
    assign layer3_outputs[745] = ~(layer2_outputs[2825]);
    assign layer3_outputs[746] = 1'b0;
    assign layer3_outputs[747] = 1'b0;
    assign layer3_outputs[748] = ~(layer2_outputs[3211]) | (layer2_outputs[104]);
    assign layer3_outputs[749] = ~(layer2_outputs[3255]) | (layer2_outputs[4299]);
    assign layer3_outputs[750] = (layer2_outputs[1129]) & ~(layer2_outputs[4069]);
    assign layer3_outputs[751] = ~(layer2_outputs[754]);
    assign layer3_outputs[752] = (layer2_outputs[5096]) & ~(layer2_outputs[882]);
    assign layer3_outputs[753] = ~((layer2_outputs[1532]) ^ (layer2_outputs[2076]));
    assign layer3_outputs[754] = (layer2_outputs[2648]) & ~(layer2_outputs[2900]);
    assign layer3_outputs[755] = ~(layer2_outputs[2703]);
    assign layer3_outputs[756] = layer2_outputs[753];
    assign layer3_outputs[757] = layer2_outputs[713];
    assign layer3_outputs[758] = layer2_outputs[4771];
    assign layer3_outputs[759] = ~(layer2_outputs[1380]) | (layer2_outputs[1475]);
    assign layer3_outputs[760] = (layer2_outputs[3476]) | (layer2_outputs[560]);
    assign layer3_outputs[761] = (layer2_outputs[2593]) & ~(layer2_outputs[1641]);
    assign layer3_outputs[762] = ~((layer2_outputs[4977]) | (layer2_outputs[3961]));
    assign layer3_outputs[763] = ~((layer2_outputs[937]) | (layer2_outputs[3018]));
    assign layer3_outputs[764] = layer2_outputs[686];
    assign layer3_outputs[765] = (layer2_outputs[2463]) & ~(layer2_outputs[761]);
    assign layer3_outputs[766] = (layer2_outputs[198]) | (layer2_outputs[204]);
    assign layer3_outputs[767] = ~(layer2_outputs[5107]) | (layer2_outputs[839]);
    assign layer3_outputs[768] = (layer2_outputs[4929]) | (layer2_outputs[1404]);
    assign layer3_outputs[769] = (layer2_outputs[2007]) & ~(layer2_outputs[3196]);
    assign layer3_outputs[770] = layer2_outputs[3849];
    assign layer3_outputs[771] = (layer2_outputs[1265]) & ~(layer2_outputs[3478]);
    assign layer3_outputs[772] = ~((layer2_outputs[1177]) ^ (layer2_outputs[3475]));
    assign layer3_outputs[773] = 1'b0;
    assign layer3_outputs[774] = ~(layer2_outputs[3008]);
    assign layer3_outputs[775] = (layer2_outputs[1539]) | (layer2_outputs[4979]);
    assign layer3_outputs[776] = ~(layer2_outputs[100]);
    assign layer3_outputs[777] = ~(layer2_outputs[1046]);
    assign layer3_outputs[778] = ~((layer2_outputs[3498]) | (layer2_outputs[3397]));
    assign layer3_outputs[779] = 1'b1;
    assign layer3_outputs[780] = (layer2_outputs[3057]) ^ (layer2_outputs[1340]);
    assign layer3_outputs[781] = ~(layer2_outputs[3266]) | (layer2_outputs[4255]);
    assign layer3_outputs[782] = (layer2_outputs[622]) & ~(layer2_outputs[2136]);
    assign layer3_outputs[783] = ~(layer2_outputs[3456]) | (layer2_outputs[2273]);
    assign layer3_outputs[784] = ~(layer2_outputs[632]) | (layer2_outputs[792]);
    assign layer3_outputs[785] = ~(layer2_outputs[3899]);
    assign layer3_outputs[786] = (layer2_outputs[1058]) & (layer2_outputs[1969]);
    assign layer3_outputs[787] = ~(layer2_outputs[3124]) | (layer2_outputs[1082]);
    assign layer3_outputs[788] = ~(layer2_outputs[814]);
    assign layer3_outputs[789] = 1'b1;
    assign layer3_outputs[790] = ~(layer2_outputs[2808]) | (layer2_outputs[2413]);
    assign layer3_outputs[791] = ~((layer2_outputs[3970]) | (layer2_outputs[1986]));
    assign layer3_outputs[792] = layer2_outputs[4935];
    assign layer3_outputs[793] = ~(layer2_outputs[869]);
    assign layer3_outputs[794] = ~(layer2_outputs[1447]) | (layer2_outputs[857]);
    assign layer3_outputs[795] = (layer2_outputs[3564]) | (layer2_outputs[4060]);
    assign layer3_outputs[796] = ~(layer2_outputs[4004]) | (layer2_outputs[983]);
    assign layer3_outputs[797] = (layer2_outputs[3846]) | (layer2_outputs[2994]);
    assign layer3_outputs[798] = 1'b1;
    assign layer3_outputs[799] = ~((layer2_outputs[3638]) | (layer2_outputs[2337]));
    assign layer3_outputs[800] = ~(layer2_outputs[2656]) | (layer2_outputs[4974]);
    assign layer3_outputs[801] = ~((layer2_outputs[4813]) | (layer2_outputs[4612]));
    assign layer3_outputs[802] = ~((layer2_outputs[2943]) & (layer2_outputs[820]));
    assign layer3_outputs[803] = ~(layer2_outputs[3568]);
    assign layer3_outputs[804] = 1'b1;
    assign layer3_outputs[805] = ~(layer2_outputs[1960]) | (layer2_outputs[4823]);
    assign layer3_outputs[806] = ~(layer2_outputs[476]);
    assign layer3_outputs[807] = (layer2_outputs[932]) | (layer2_outputs[63]);
    assign layer3_outputs[808] = 1'b1;
    assign layer3_outputs[809] = ~(layer2_outputs[3302]);
    assign layer3_outputs[810] = ~(layer2_outputs[4236]);
    assign layer3_outputs[811] = (layer2_outputs[2546]) | (layer2_outputs[1067]);
    assign layer3_outputs[812] = layer2_outputs[1542];
    assign layer3_outputs[813] = 1'b0;
    assign layer3_outputs[814] = 1'b0;
    assign layer3_outputs[815] = ~(layer2_outputs[1005]) | (layer2_outputs[2107]);
    assign layer3_outputs[816] = ~(layer2_outputs[1612]);
    assign layer3_outputs[817] = ~((layer2_outputs[2319]) & (layer2_outputs[4262]));
    assign layer3_outputs[818] = 1'b0;
    assign layer3_outputs[819] = 1'b0;
    assign layer3_outputs[820] = ~((layer2_outputs[2973]) & (layer2_outputs[3063]));
    assign layer3_outputs[821] = ~(layer2_outputs[2521]);
    assign layer3_outputs[822] = ~(layer2_outputs[2843]) | (layer2_outputs[4300]);
    assign layer3_outputs[823] = ~(layer2_outputs[15]);
    assign layer3_outputs[824] = layer2_outputs[2644];
    assign layer3_outputs[825] = ~(layer2_outputs[4436]);
    assign layer3_outputs[826] = ~(layer2_outputs[2944]) | (layer2_outputs[702]);
    assign layer3_outputs[827] = (layer2_outputs[3405]) & (layer2_outputs[2355]);
    assign layer3_outputs[828] = (layer2_outputs[102]) | (layer2_outputs[4870]);
    assign layer3_outputs[829] = (layer2_outputs[4825]) ^ (layer2_outputs[1172]);
    assign layer3_outputs[830] = 1'b1;
    assign layer3_outputs[831] = layer2_outputs[4098];
    assign layer3_outputs[832] = layer2_outputs[3943];
    assign layer3_outputs[833] = ~((layer2_outputs[947]) & (layer2_outputs[4661]));
    assign layer3_outputs[834] = layer2_outputs[2068];
    assign layer3_outputs[835] = 1'b1;
    assign layer3_outputs[836] = (layer2_outputs[719]) & ~(layer2_outputs[2277]);
    assign layer3_outputs[837] = (layer2_outputs[1341]) & ~(layer2_outputs[1888]);
    assign layer3_outputs[838] = ~(layer2_outputs[1703]);
    assign layer3_outputs[839] = 1'b1;
    assign layer3_outputs[840] = 1'b1;
    assign layer3_outputs[841] = (layer2_outputs[727]) & ~(layer2_outputs[1979]);
    assign layer3_outputs[842] = ~(layer2_outputs[2670]);
    assign layer3_outputs[843] = layer2_outputs[4467];
    assign layer3_outputs[844] = ~((layer2_outputs[2136]) | (layer2_outputs[937]));
    assign layer3_outputs[845] = (layer2_outputs[2804]) | (layer2_outputs[2817]);
    assign layer3_outputs[846] = 1'b0;
    assign layer3_outputs[847] = 1'b1;
    assign layer3_outputs[848] = (layer2_outputs[4482]) & ~(layer2_outputs[1581]);
    assign layer3_outputs[849] = ~(layer2_outputs[2305]);
    assign layer3_outputs[850] = ~((layer2_outputs[2812]) | (layer2_outputs[4879]));
    assign layer3_outputs[851] = layer2_outputs[3547];
    assign layer3_outputs[852] = layer2_outputs[2669];
    assign layer3_outputs[853] = (layer2_outputs[4149]) & ~(layer2_outputs[171]);
    assign layer3_outputs[854] = (layer2_outputs[931]) | (layer2_outputs[3126]);
    assign layer3_outputs[855] = 1'b0;
    assign layer3_outputs[856] = layer2_outputs[2042];
    assign layer3_outputs[857] = (layer2_outputs[2108]) | (layer2_outputs[4839]);
    assign layer3_outputs[858] = (layer2_outputs[111]) ^ (layer2_outputs[3763]);
    assign layer3_outputs[859] = 1'b1;
    assign layer3_outputs[860] = layer2_outputs[1710];
    assign layer3_outputs[861] = (layer2_outputs[1201]) & ~(layer2_outputs[3526]);
    assign layer3_outputs[862] = 1'b0;
    assign layer3_outputs[863] = layer2_outputs[2647];
    assign layer3_outputs[864] = 1'b1;
    assign layer3_outputs[865] = (layer2_outputs[2569]) & (layer2_outputs[1486]);
    assign layer3_outputs[866] = ~(layer2_outputs[3577]);
    assign layer3_outputs[867] = 1'b1;
    assign layer3_outputs[868] = (layer2_outputs[4891]) & (layer2_outputs[2148]);
    assign layer3_outputs[869] = (layer2_outputs[2983]) & (layer2_outputs[3711]);
    assign layer3_outputs[870] = ~((layer2_outputs[3856]) & (layer2_outputs[2241]));
    assign layer3_outputs[871] = layer2_outputs[3715];
    assign layer3_outputs[872] = ~(layer2_outputs[603]) | (layer2_outputs[5038]);
    assign layer3_outputs[873] = layer2_outputs[2938];
    assign layer3_outputs[874] = (layer2_outputs[3787]) & (layer2_outputs[1577]);
    assign layer3_outputs[875] = 1'b0;
    assign layer3_outputs[876] = ~(layer2_outputs[2415]) | (layer2_outputs[3728]);
    assign layer3_outputs[877] = layer2_outputs[4428];
    assign layer3_outputs[878] = ~((layer2_outputs[2034]) ^ (layer2_outputs[2797]));
    assign layer3_outputs[879] = ~(layer2_outputs[250]);
    assign layer3_outputs[880] = ~((layer2_outputs[5111]) & (layer2_outputs[1803]));
    assign layer3_outputs[881] = ~(layer2_outputs[1472]);
    assign layer3_outputs[882] = ~(layer2_outputs[2980]) | (layer2_outputs[696]);
    assign layer3_outputs[883] = ~((layer2_outputs[4386]) | (layer2_outputs[3514]));
    assign layer3_outputs[884] = (layer2_outputs[4204]) & ~(layer2_outputs[2267]);
    assign layer3_outputs[885] = ~(layer2_outputs[4509]);
    assign layer3_outputs[886] = ~((layer2_outputs[3881]) ^ (layer2_outputs[3468]));
    assign layer3_outputs[887] = (layer2_outputs[2902]) | (layer2_outputs[3273]);
    assign layer3_outputs[888] = ~(layer2_outputs[1054]);
    assign layer3_outputs[889] = 1'b1;
    assign layer3_outputs[890] = (layer2_outputs[1796]) | (layer2_outputs[4103]);
    assign layer3_outputs[891] = layer2_outputs[2843];
    assign layer3_outputs[892] = layer2_outputs[1893];
    assign layer3_outputs[893] = ~((layer2_outputs[2510]) | (layer2_outputs[1343]));
    assign layer3_outputs[894] = 1'b0;
    assign layer3_outputs[895] = 1'b1;
    assign layer3_outputs[896] = ~(layer2_outputs[2935]) | (layer2_outputs[1586]);
    assign layer3_outputs[897] = ~(layer2_outputs[1932]);
    assign layer3_outputs[898] = ~(layer2_outputs[1987]) | (layer2_outputs[2782]);
    assign layer3_outputs[899] = ~((layer2_outputs[1759]) & (layer2_outputs[352]));
    assign layer3_outputs[900] = 1'b0;
    assign layer3_outputs[901] = ~(layer2_outputs[1407]) | (layer2_outputs[3939]);
    assign layer3_outputs[902] = (layer2_outputs[2227]) & ~(layer2_outputs[4453]);
    assign layer3_outputs[903] = (layer2_outputs[3281]) | (layer2_outputs[3368]);
    assign layer3_outputs[904] = ~(layer2_outputs[4630]);
    assign layer3_outputs[905] = ~(layer2_outputs[588]);
    assign layer3_outputs[906] = ~(layer2_outputs[3944]) | (layer2_outputs[3727]);
    assign layer3_outputs[907] = ~(layer2_outputs[973]);
    assign layer3_outputs[908] = ~(layer2_outputs[3994]);
    assign layer3_outputs[909] = ~(layer2_outputs[5023]);
    assign layer3_outputs[910] = ~(layer2_outputs[962]) | (layer2_outputs[4255]);
    assign layer3_outputs[911] = 1'b0;
    assign layer3_outputs[912] = ~(layer2_outputs[4778]);
    assign layer3_outputs[913] = layer2_outputs[3990];
    assign layer3_outputs[914] = ~(layer2_outputs[1814]);
    assign layer3_outputs[915] = ~((layer2_outputs[118]) ^ (layer2_outputs[3932]));
    assign layer3_outputs[916] = layer2_outputs[3901];
    assign layer3_outputs[917] = 1'b1;
    assign layer3_outputs[918] = ~((layer2_outputs[1399]) ^ (layer2_outputs[4551]));
    assign layer3_outputs[919] = ~((layer2_outputs[3351]) ^ (layer2_outputs[2312]));
    assign layer3_outputs[920] = (layer2_outputs[189]) | (layer2_outputs[639]);
    assign layer3_outputs[921] = ~(layer2_outputs[2519]);
    assign layer3_outputs[922] = 1'b0;
    assign layer3_outputs[923] = ~(layer2_outputs[2903]);
    assign layer3_outputs[924] = 1'b1;
    assign layer3_outputs[925] = layer2_outputs[1980];
    assign layer3_outputs[926] = ~((layer2_outputs[4051]) | (layer2_outputs[667]));
    assign layer3_outputs[927] = ~((layer2_outputs[1725]) | (layer2_outputs[4674]));
    assign layer3_outputs[928] = (layer2_outputs[5007]) & ~(layer2_outputs[3199]);
    assign layer3_outputs[929] = ~((layer2_outputs[3560]) | (layer2_outputs[1805]));
    assign layer3_outputs[930] = ~(layer2_outputs[3403]);
    assign layer3_outputs[931] = (layer2_outputs[2412]) ^ (layer2_outputs[164]);
    assign layer3_outputs[932] = ~(layer2_outputs[4127]);
    assign layer3_outputs[933] = ~(layer2_outputs[4684]) | (layer2_outputs[2812]);
    assign layer3_outputs[934] = ~(layer2_outputs[904]) | (layer2_outputs[4335]);
    assign layer3_outputs[935] = ~(layer2_outputs[1653]);
    assign layer3_outputs[936] = ~(layer2_outputs[3236]) | (layer2_outputs[1885]);
    assign layer3_outputs[937] = ~(layer2_outputs[520]);
    assign layer3_outputs[938] = (layer2_outputs[243]) & ~(layer2_outputs[1354]);
    assign layer3_outputs[939] = ~((layer2_outputs[3311]) ^ (layer2_outputs[905]));
    assign layer3_outputs[940] = 1'b0;
    assign layer3_outputs[941] = ~(layer2_outputs[2481]);
    assign layer3_outputs[942] = (layer2_outputs[1502]) & (layer2_outputs[1260]);
    assign layer3_outputs[943] = (layer2_outputs[1561]) | (layer2_outputs[3594]);
    assign layer3_outputs[944] = ~(layer2_outputs[4025]);
    assign layer3_outputs[945] = (layer2_outputs[2083]) & (layer2_outputs[4351]);
    assign layer3_outputs[946] = ~(layer2_outputs[2166]) | (layer2_outputs[2177]);
    assign layer3_outputs[947] = ~((layer2_outputs[3368]) | (layer2_outputs[4988]));
    assign layer3_outputs[948] = (layer2_outputs[5101]) & (layer2_outputs[756]);
    assign layer3_outputs[949] = layer2_outputs[2278];
    assign layer3_outputs[950] = layer2_outputs[1868];
    assign layer3_outputs[951] = (layer2_outputs[3564]) | (layer2_outputs[4036]);
    assign layer3_outputs[952] = (layer2_outputs[4455]) & ~(layer2_outputs[4961]);
    assign layer3_outputs[953] = layer2_outputs[1365];
    assign layer3_outputs[954] = (layer2_outputs[1732]) & ~(layer2_outputs[743]);
    assign layer3_outputs[955] = layer2_outputs[3429];
    assign layer3_outputs[956] = (layer2_outputs[2286]) & (layer2_outputs[1508]);
    assign layer3_outputs[957] = (layer2_outputs[4289]) & (layer2_outputs[2972]);
    assign layer3_outputs[958] = (layer2_outputs[1779]) & (layer2_outputs[54]);
    assign layer3_outputs[959] = 1'b0;
    assign layer3_outputs[960] = ~(layer2_outputs[3889]) | (layer2_outputs[412]);
    assign layer3_outputs[961] = layer2_outputs[3492];
    assign layer3_outputs[962] = (layer2_outputs[2917]) ^ (layer2_outputs[2531]);
    assign layer3_outputs[963] = ~(layer2_outputs[1939]) | (layer2_outputs[2618]);
    assign layer3_outputs[964] = ~((layer2_outputs[4018]) ^ (layer2_outputs[3929]));
    assign layer3_outputs[965] = layer2_outputs[3383];
    assign layer3_outputs[966] = (layer2_outputs[1784]) & ~(layer2_outputs[2448]);
    assign layer3_outputs[967] = (layer2_outputs[3208]) ^ (layer2_outputs[4855]);
    assign layer3_outputs[968] = layer2_outputs[1949];
    assign layer3_outputs[969] = (layer2_outputs[2959]) & (layer2_outputs[552]);
    assign layer3_outputs[970] = (layer2_outputs[3181]) | (layer2_outputs[4038]);
    assign layer3_outputs[971] = 1'b1;
    assign layer3_outputs[972] = ~(layer2_outputs[3166]);
    assign layer3_outputs[973] = ~(layer2_outputs[370]);
    assign layer3_outputs[974] = (layer2_outputs[2090]) & ~(layer2_outputs[3343]);
    assign layer3_outputs[975] = ~(layer2_outputs[3885]) | (layer2_outputs[3953]);
    assign layer3_outputs[976] = layer2_outputs[2435];
    assign layer3_outputs[977] = (layer2_outputs[3400]) & ~(layer2_outputs[3903]);
    assign layer3_outputs[978] = ~((layer2_outputs[3224]) & (layer2_outputs[2879]));
    assign layer3_outputs[979] = (layer2_outputs[190]) & ~(layer2_outputs[2687]);
    assign layer3_outputs[980] = ~(layer2_outputs[4005]) | (layer2_outputs[3950]);
    assign layer3_outputs[981] = layer2_outputs[2229];
    assign layer3_outputs[982] = ~((layer2_outputs[2952]) | (layer2_outputs[2341]));
    assign layer3_outputs[983] = ~(layer2_outputs[372]) | (layer2_outputs[253]);
    assign layer3_outputs[984] = ~((layer2_outputs[3339]) & (layer2_outputs[362]));
    assign layer3_outputs[985] = ~(layer2_outputs[193]) | (layer2_outputs[3935]);
    assign layer3_outputs[986] = ~((layer2_outputs[418]) & (layer2_outputs[350]));
    assign layer3_outputs[987] = layer2_outputs[2302];
    assign layer3_outputs[988] = ~(layer2_outputs[3280]);
    assign layer3_outputs[989] = ~(layer2_outputs[3021]);
    assign layer3_outputs[990] = ~(layer2_outputs[3289]) | (layer2_outputs[1521]);
    assign layer3_outputs[991] = ~((layer2_outputs[4861]) ^ (layer2_outputs[4422]));
    assign layer3_outputs[992] = (layer2_outputs[4257]) & ~(layer2_outputs[655]);
    assign layer3_outputs[993] = ~((layer2_outputs[2333]) | (layer2_outputs[1360]));
    assign layer3_outputs[994] = layer2_outputs[2366];
    assign layer3_outputs[995] = 1'b0;
    assign layer3_outputs[996] = layer2_outputs[1075];
    assign layer3_outputs[997] = (layer2_outputs[3331]) & ~(layer2_outputs[4994]);
    assign layer3_outputs[998] = ~((layer2_outputs[3664]) | (layer2_outputs[1576]));
    assign layer3_outputs[999] = ~(layer2_outputs[1013]) | (layer2_outputs[1622]);
    assign layer3_outputs[1000] = layer2_outputs[2526];
    assign layer3_outputs[1001] = (layer2_outputs[1996]) | (layer2_outputs[1818]);
    assign layer3_outputs[1002] = ~(layer2_outputs[3928]) | (layer2_outputs[2876]);
    assign layer3_outputs[1003] = ~((layer2_outputs[2097]) & (layer2_outputs[2815]));
    assign layer3_outputs[1004] = ~(layer2_outputs[2359]) | (layer2_outputs[3222]);
    assign layer3_outputs[1005] = layer2_outputs[4884];
    assign layer3_outputs[1006] = ~(layer2_outputs[4452]);
    assign layer3_outputs[1007] = ~(layer2_outputs[426]);
    assign layer3_outputs[1008] = ~(layer2_outputs[3234]) | (layer2_outputs[1507]);
    assign layer3_outputs[1009] = (layer2_outputs[3183]) | (layer2_outputs[4636]);
    assign layer3_outputs[1010] = (layer2_outputs[1377]) & (layer2_outputs[3394]);
    assign layer3_outputs[1011] = layer2_outputs[1196];
    assign layer3_outputs[1012] = ~(layer2_outputs[2988]);
    assign layer3_outputs[1013] = ~((layer2_outputs[808]) | (layer2_outputs[356]));
    assign layer3_outputs[1014] = (layer2_outputs[3101]) | (layer2_outputs[455]);
    assign layer3_outputs[1015] = ~((layer2_outputs[100]) & (layer2_outputs[4347]));
    assign layer3_outputs[1016] = ~((layer2_outputs[3065]) & (layer2_outputs[985]));
    assign layer3_outputs[1017] = ~(layer2_outputs[2990]) | (layer2_outputs[3471]);
    assign layer3_outputs[1018] = (layer2_outputs[1132]) & (layer2_outputs[688]);
    assign layer3_outputs[1019] = (layer2_outputs[1640]) & ~(layer2_outputs[2718]);
    assign layer3_outputs[1020] = ~(layer2_outputs[2018]);
    assign layer3_outputs[1021] = ~(layer2_outputs[5098]) | (layer2_outputs[4011]);
    assign layer3_outputs[1022] = ~((layer2_outputs[4183]) | (layer2_outputs[509]));
    assign layer3_outputs[1023] = ~(layer2_outputs[1226]);
    assign layer3_outputs[1024] = (layer2_outputs[730]) | (layer2_outputs[1716]);
    assign layer3_outputs[1025] = ~(layer2_outputs[1387]);
    assign layer3_outputs[1026] = layer2_outputs[294];
    assign layer3_outputs[1027] = ~(layer2_outputs[4273]);
    assign layer3_outputs[1028] = ~(layer2_outputs[605]);
    assign layer3_outputs[1029] = ~(layer2_outputs[4875]) | (layer2_outputs[2668]);
    assign layer3_outputs[1030] = ~(layer2_outputs[4141]);
    assign layer3_outputs[1031] = 1'b1;
    assign layer3_outputs[1032] = layer2_outputs[2492];
    assign layer3_outputs[1033] = ~((layer2_outputs[226]) & (layer2_outputs[4212]));
    assign layer3_outputs[1034] = layer2_outputs[3843];
    assign layer3_outputs[1035] = ~(layer2_outputs[4350]);
    assign layer3_outputs[1036] = 1'b0;
    assign layer3_outputs[1037] = ~(layer2_outputs[4566]);
    assign layer3_outputs[1038] = ~((layer2_outputs[3533]) & (layer2_outputs[3782]));
    assign layer3_outputs[1039] = ~((layer2_outputs[936]) | (layer2_outputs[4620]));
    assign layer3_outputs[1040] = 1'b0;
    assign layer3_outputs[1041] = ~(layer2_outputs[3808]);
    assign layer3_outputs[1042] = (layer2_outputs[4309]) & ~(layer2_outputs[976]);
    assign layer3_outputs[1043] = ~(layer2_outputs[2677]) | (layer2_outputs[921]);
    assign layer3_outputs[1044] = (layer2_outputs[2257]) & (layer2_outputs[3295]);
    assign layer3_outputs[1045] = layer2_outputs[3468];
    assign layer3_outputs[1046] = (layer2_outputs[2347]) | (layer2_outputs[1476]);
    assign layer3_outputs[1047] = ~(layer2_outputs[3169]);
    assign layer3_outputs[1048] = layer2_outputs[489];
    assign layer3_outputs[1049] = 1'b1;
    assign layer3_outputs[1050] = ~(layer2_outputs[518]) | (layer2_outputs[212]);
    assign layer3_outputs[1051] = ~(layer2_outputs[1509]);
    assign layer3_outputs[1052] = layer2_outputs[4938];
    assign layer3_outputs[1053] = layer2_outputs[662];
    assign layer3_outputs[1054] = ~((layer2_outputs[1776]) & (layer2_outputs[2922]));
    assign layer3_outputs[1055] = ~((layer2_outputs[1323]) | (layer2_outputs[2561]));
    assign layer3_outputs[1056] = layer2_outputs[431];
    assign layer3_outputs[1057] = layer2_outputs[4383];
    assign layer3_outputs[1058] = layer2_outputs[4841];
    assign layer3_outputs[1059] = (layer2_outputs[3062]) & ~(layer2_outputs[4906]);
    assign layer3_outputs[1060] = 1'b0;
    assign layer3_outputs[1061] = 1'b1;
    assign layer3_outputs[1062] = layer2_outputs[4744];
    assign layer3_outputs[1063] = 1'b1;
    assign layer3_outputs[1064] = ~(layer2_outputs[2013]);
    assign layer3_outputs[1065] = layer2_outputs[1087];
    assign layer3_outputs[1066] = ~(layer2_outputs[1896]) | (layer2_outputs[644]);
    assign layer3_outputs[1067] = (layer2_outputs[2432]) ^ (layer2_outputs[1690]);
    assign layer3_outputs[1068] = (layer2_outputs[4491]) | (layer2_outputs[4619]);
    assign layer3_outputs[1069] = (layer2_outputs[2851]) | (layer2_outputs[3178]);
    assign layer3_outputs[1070] = (layer2_outputs[164]) & ~(layer2_outputs[2813]);
    assign layer3_outputs[1071] = ~(layer2_outputs[1201]) | (layer2_outputs[3920]);
    assign layer3_outputs[1072] = 1'b1;
    assign layer3_outputs[1073] = (layer2_outputs[3441]) & (layer2_outputs[602]);
    assign layer3_outputs[1074] = 1'b1;
    assign layer3_outputs[1075] = ~(layer2_outputs[1233]);
    assign layer3_outputs[1076] = 1'b0;
    assign layer3_outputs[1077] = 1'b0;
    assign layer3_outputs[1078] = layer2_outputs[1570];
    assign layer3_outputs[1079] = (layer2_outputs[3865]) & ~(layer2_outputs[894]);
    assign layer3_outputs[1080] = layer2_outputs[4780];
    assign layer3_outputs[1081] = ~((layer2_outputs[961]) & (layer2_outputs[3035]));
    assign layer3_outputs[1082] = ~(layer2_outputs[3853]);
    assign layer3_outputs[1083] = ~(layer2_outputs[2230]);
    assign layer3_outputs[1084] = ~(layer2_outputs[2941]) | (layer2_outputs[3508]);
    assign layer3_outputs[1085] = 1'b0;
    assign layer3_outputs[1086] = layer2_outputs[244];
    assign layer3_outputs[1087] = layer2_outputs[1057];
    assign layer3_outputs[1088] = 1'b1;
    assign layer3_outputs[1089] = ~(layer2_outputs[768]);
    assign layer3_outputs[1090] = ~((layer2_outputs[4523]) & (layer2_outputs[85]));
    assign layer3_outputs[1091] = layer2_outputs[1556];
    assign layer3_outputs[1092] = ~((layer2_outputs[2561]) & (layer2_outputs[4967]));
    assign layer3_outputs[1093] = (layer2_outputs[2200]) & (layer2_outputs[3193]);
    assign layer3_outputs[1094] = (layer2_outputs[537]) & (layer2_outputs[4695]);
    assign layer3_outputs[1095] = ~((layer2_outputs[3874]) ^ (layer2_outputs[60]));
    assign layer3_outputs[1096] = (layer2_outputs[700]) & ~(layer2_outputs[4228]);
    assign layer3_outputs[1097] = layer2_outputs[4046];
    assign layer3_outputs[1098] = layer2_outputs[384];
    assign layer3_outputs[1099] = layer2_outputs[4242];
    assign layer3_outputs[1100] = (layer2_outputs[1658]) & ~(layer2_outputs[2167]);
    assign layer3_outputs[1101] = (layer2_outputs[2113]) & ~(layer2_outputs[3501]);
    assign layer3_outputs[1102] = ~(layer2_outputs[3943]);
    assign layer3_outputs[1103] = (layer2_outputs[2418]) & ~(layer2_outputs[817]);
    assign layer3_outputs[1104] = ~(layer2_outputs[657]) | (layer2_outputs[1006]);
    assign layer3_outputs[1105] = (layer2_outputs[4058]) & (layer2_outputs[4411]);
    assign layer3_outputs[1106] = ~(layer2_outputs[3518]);
    assign layer3_outputs[1107] = (layer2_outputs[2453]) & ~(layer2_outputs[2003]);
    assign layer3_outputs[1108] = 1'b1;
    assign layer3_outputs[1109] = (layer2_outputs[2681]) & ~(layer2_outputs[1216]);
    assign layer3_outputs[1110] = 1'b1;
    assign layer3_outputs[1111] = (layer2_outputs[3587]) & (layer2_outputs[1438]);
    assign layer3_outputs[1112] = ~((layer2_outputs[454]) | (layer2_outputs[3675]));
    assign layer3_outputs[1113] = (layer2_outputs[3516]) & ~(layer2_outputs[4671]);
    assign layer3_outputs[1114] = (layer2_outputs[103]) | (layer2_outputs[3612]);
    assign layer3_outputs[1115] = ~(layer2_outputs[1438]) | (layer2_outputs[4631]);
    assign layer3_outputs[1116] = layer2_outputs[4593];
    assign layer3_outputs[1117] = ~((layer2_outputs[3708]) ^ (layer2_outputs[4656]));
    assign layer3_outputs[1118] = layer2_outputs[4585];
    assign layer3_outputs[1119] = ~(layer2_outputs[57]) | (layer2_outputs[2170]);
    assign layer3_outputs[1120] = 1'b1;
    assign layer3_outputs[1121] = ~(layer2_outputs[594]);
    assign layer3_outputs[1122] = layer2_outputs[4999];
    assign layer3_outputs[1123] = ~(layer2_outputs[3092]);
    assign layer3_outputs[1124] = ~(layer2_outputs[2714]) | (layer2_outputs[3677]);
    assign layer3_outputs[1125] = (layer2_outputs[5066]) ^ (layer2_outputs[3333]);
    assign layer3_outputs[1126] = 1'b0;
    assign layer3_outputs[1127] = layer2_outputs[3361];
    assign layer3_outputs[1128] = (layer2_outputs[795]) | (layer2_outputs[1559]);
    assign layer3_outputs[1129] = 1'b1;
    assign layer3_outputs[1130] = (layer2_outputs[3655]) & (layer2_outputs[1439]);
    assign layer3_outputs[1131] = layer2_outputs[4720];
    assign layer3_outputs[1132] = ~(layer2_outputs[3748]) | (layer2_outputs[2011]);
    assign layer3_outputs[1133] = 1'b0;
    assign layer3_outputs[1134] = 1'b1;
    assign layer3_outputs[1135] = 1'b0;
    assign layer3_outputs[1136] = ~(layer2_outputs[1767]);
    assign layer3_outputs[1137] = ~(layer2_outputs[4659]) | (layer2_outputs[1581]);
    assign layer3_outputs[1138] = ~(layer2_outputs[1682]) | (layer2_outputs[5017]);
    assign layer3_outputs[1139] = 1'b1;
    assign layer3_outputs[1140] = ~(layer2_outputs[3382]) | (layer2_outputs[3343]);
    assign layer3_outputs[1141] = (layer2_outputs[1027]) & ~(layer2_outputs[441]);
    assign layer3_outputs[1142] = 1'b1;
    assign layer3_outputs[1143] = ~(layer2_outputs[4103]);
    assign layer3_outputs[1144] = ~((layer2_outputs[4111]) & (layer2_outputs[890]));
    assign layer3_outputs[1145] = ~(layer2_outputs[5108]) | (layer2_outputs[4532]);
    assign layer3_outputs[1146] = 1'b0;
    assign layer3_outputs[1147] = 1'b1;
    assign layer3_outputs[1148] = layer2_outputs[2351];
    assign layer3_outputs[1149] = (layer2_outputs[320]) & (layer2_outputs[1415]);
    assign layer3_outputs[1150] = layer2_outputs[3801];
    assign layer3_outputs[1151] = ~((layer2_outputs[499]) | (layer2_outputs[221]));
    assign layer3_outputs[1152] = (layer2_outputs[3355]) & ~(layer2_outputs[53]);
    assign layer3_outputs[1153] = ~(layer2_outputs[4564]) | (layer2_outputs[194]);
    assign layer3_outputs[1154] = (layer2_outputs[3413]) | (layer2_outputs[2674]);
    assign layer3_outputs[1155] = ~(layer2_outputs[3644]);
    assign layer3_outputs[1156] = ~(layer2_outputs[2878]);
    assign layer3_outputs[1157] = ~((layer2_outputs[353]) & (layer2_outputs[2142]));
    assign layer3_outputs[1158] = ~(layer2_outputs[3059]);
    assign layer3_outputs[1159] = ~(layer2_outputs[2915]);
    assign layer3_outputs[1160] = ~(layer2_outputs[2898]) | (layer2_outputs[3291]);
    assign layer3_outputs[1161] = ~((layer2_outputs[1246]) ^ (layer2_outputs[4221]));
    assign layer3_outputs[1162] = 1'b0;
    assign layer3_outputs[1163] = ~(layer2_outputs[2890]) | (layer2_outputs[2474]);
    assign layer3_outputs[1164] = layer2_outputs[744];
    assign layer3_outputs[1165] = 1'b1;
    assign layer3_outputs[1166] = ~(layer2_outputs[2093]) | (layer2_outputs[4925]);
    assign layer3_outputs[1167] = (layer2_outputs[2887]) & (layer2_outputs[3625]);
    assign layer3_outputs[1168] = layer2_outputs[4007];
    assign layer3_outputs[1169] = (layer2_outputs[2867]) & (layer2_outputs[2321]);
    assign layer3_outputs[1170] = layer2_outputs[3034];
    assign layer3_outputs[1171] = ~((layer2_outputs[51]) & (layer2_outputs[1425]));
    assign layer3_outputs[1172] = ~(layer2_outputs[3354]) | (layer2_outputs[2631]);
    assign layer3_outputs[1173] = ~(layer2_outputs[4001]);
    assign layer3_outputs[1174] = (layer2_outputs[4193]) & (layer2_outputs[403]);
    assign layer3_outputs[1175] = (layer2_outputs[28]) & (layer2_outputs[787]);
    assign layer3_outputs[1176] = ~(layer2_outputs[2072]);
    assign layer3_outputs[1177] = layer2_outputs[81];
    assign layer3_outputs[1178] = ~((layer2_outputs[2018]) & (layer2_outputs[2839]));
    assign layer3_outputs[1179] = (layer2_outputs[968]) & ~(layer2_outputs[5021]);
    assign layer3_outputs[1180] = ~(layer2_outputs[3272]);
    assign layer3_outputs[1181] = ~((layer2_outputs[997]) & (layer2_outputs[4284]));
    assign layer3_outputs[1182] = (layer2_outputs[3870]) | (layer2_outputs[4303]);
    assign layer3_outputs[1183] = layer2_outputs[2726];
    assign layer3_outputs[1184] = ~(layer2_outputs[4083]) | (layer2_outputs[586]);
    assign layer3_outputs[1185] = ~(layer2_outputs[1356]);
    assign layer3_outputs[1186] = 1'b0;
    assign layer3_outputs[1187] = ~((layer2_outputs[3284]) | (layer2_outputs[2477]));
    assign layer3_outputs[1188] = layer2_outputs[4380];
    assign layer3_outputs[1189] = ~(layer2_outputs[3264]) | (layer2_outputs[296]);
    assign layer3_outputs[1190] = ~(layer2_outputs[2457]);
    assign layer3_outputs[1191] = ~((layer2_outputs[4980]) & (layer2_outputs[4097]));
    assign layer3_outputs[1192] = ~(layer2_outputs[3270]) | (layer2_outputs[2393]);
    assign layer3_outputs[1193] = ~(layer2_outputs[3756]);
    assign layer3_outputs[1194] = ~(layer2_outputs[2314]) | (layer2_outputs[119]);
    assign layer3_outputs[1195] = layer2_outputs[4285];
    assign layer3_outputs[1196] = ~((layer2_outputs[2170]) & (layer2_outputs[1177]));
    assign layer3_outputs[1197] = (layer2_outputs[4763]) | (layer2_outputs[2466]);
    assign layer3_outputs[1198] = ~(layer2_outputs[3516]);
    assign layer3_outputs[1199] = ~(layer2_outputs[3191]);
    assign layer3_outputs[1200] = layer2_outputs[1174];
    assign layer3_outputs[1201] = ~((layer2_outputs[2252]) | (layer2_outputs[1637]));
    assign layer3_outputs[1202] = layer2_outputs[4513];
    assign layer3_outputs[1203] = (layer2_outputs[4100]) | (layer2_outputs[1410]);
    assign layer3_outputs[1204] = (layer2_outputs[2641]) ^ (layer2_outputs[4070]);
    assign layer3_outputs[1205] = ~((layer2_outputs[3906]) | (layer2_outputs[1338]));
    assign layer3_outputs[1206] = (layer2_outputs[511]) & (layer2_outputs[954]);
    assign layer3_outputs[1207] = ~(layer2_outputs[144]);
    assign layer3_outputs[1208] = ~((layer2_outputs[1648]) & (layer2_outputs[4463]));
    assign layer3_outputs[1209] = layer2_outputs[2662];
    assign layer3_outputs[1210] = ~(layer2_outputs[850]);
    assign layer3_outputs[1211] = ~(layer2_outputs[2570]);
    assign layer3_outputs[1212] = (layer2_outputs[2193]) & ~(layer2_outputs[652]);
    assign layer3_outputs[1213] = ~((layer2_outputs[4077]) & (layer2_outputs[2342]));
    assign layer3_outputs[1214] = (layer2_outputs[532]) & ~(layer2_outputs[1613]);
    assign layer3_outputs[1215] = ~(layer2_outputs[1238]);
    assign layer3_outputs[1216] = layer2_outputs[3144];
    assign layer3_outputs[1217] = 1'b0;
    assign layer3_outputs[1218] = ~((layer2_outputs[3377]) ^ (layer2_outputs[2221]));
    assign layer3_outputs[1219] = ~((layer2_outputs[3716]) | (layer2_outputs[3061]));
    assign layer3_outputs[1220] = (layer2_outputs[3118]) & ~(layer2_outputs[1855]);
    assign layer3_outputs[1221] = 1'b1;
    assign layer3_outputs[1222] = 1'b0;
    assign layer3_outputs[1223] = 1'b0;
    assign layer3_outputs[1224] = (layer2_outputs[3349]) & (layer2_outputs[1145]);
    assign layer3_outputs[1225] = ~((layer2_outputs[4626]) & (layer2_outputs[3349]));
    assign layer3_outputs[1226] = layer2_outputs[4064];
    assign layer3_outputs[1227] = ~((layer2_outputs[1893]) | (layer2_outputs[1490]));
    assign layer3_outputs[1228] = 1'b0;
    assign layer3_outputs[1229] = ~((layer2_outputs[2783]) ^ (layer2_outputs[767]));
    assign layer3_outputs[1230] = layer2_outputs[383];
    assign layer3_outputs[1231] = ~((layer2_outputs[4984]) & (layer2_outputs[2451]));
    assign layer3_outputs[1232] = layer2_outputs[859];
    assign layer3_outputs[1233] = layer2_outputs[1335];
    assign layer3_outputs[1234] = ~((layer2_outputs[192]) & (layer2_outputs[1825]));
    assign layer3_outputs[1235] = layer2_outputs[2795];
    assign layer3_outputs[1236] = (layer2_outputs[4358]) ^ (layer2_outputs[853]);
    assign layer3_outputs[1237] = ~((layer2_outputs[1252]) | (layer2_outputs[2979]));
    assign layer3_outputs[1238] = ~(layer2_outputs[2698]) | (layer2_outputs[4580]);
    assign layer3_outputs[1239] = 1'b1;
    assign layer3_outputs[1240] = ~((layer2_outputs[1]) & (layer2_outputs[2831]));
    assign layer3_outputs[1241] = ~(layer2_outputs[260]);
    assign layer3_outputs[1242] = ~((layer2_outputs[3698]) & (layer2_outputs[4785]));
    assign layer3_outputs[1243] = ~(layer2_outputs[4672]);
    assign layer3_outputs[1244] = layer2_outputs[1198];
    assign layer3_outputs[1245] = ~(layer2_outputs[2552]) | (layer2_outputs[4491]);
    assign layer3_outputs[1246] = ~(layer2_outputs[253]);
    assign layer3_outputs[1247] = (layer2_outputs[2429]) | (layer2_outputs[4586]);
    assign layer3_outputs[1248] = ~(layer2_outputs[4989]);
    assign layer3_outputs[1249] = layer2_outputs[991];
    assign layer3_outputs[1250] = (layer2_outputs[1717]) | (layer2_outputs[862]);
    assign layer3_outputs[1251] = 1'b0;
    assign layer3_outputs[1252] = (layer2_outputs[3229]) & ~(layer2_outputs[95]);
    assign layer3_outputs[1253] = ~((layer2_outputs[4229]) | (layer2_outputs[718]));
    assign layer3_outputs[1254] = 1'b1;
    assign layer3_outputs[1255] = 1'b0;
    assign layer3_outputs[1256] = ~(layer2_outputs[1985]);
    assign layer3_outputs[1257] = layer2_outputs[4816];
    assign layer3_outputs[1258] = ~((layer2_outputs[3536]) | (layer2_outputs[568]));
    assign layer3_outputs[1259] = ~(layer2_outputs[421]);
    assign layer3_outputs[1260] = ~((layer2_outputs[307]) | (layer2_outputs[2455]));
    assign layer3_outputs[1261] = ~(layer2_outputs[2076]);
    assign layer3_outputs[1262] = ~(layer2_outputs[4467]) | (layer2_outputs[1023]);
    assign layer3_outputs[1263] = ~((layer2_outputs[4673]) & (layer2_outputs[187]));
    assign layer3_outputs[1264] = ~((layer2_outputs[1087]) & (layer2_outputs[934]));
    assign layer3_outputs[1265] = 1'b0;
    assign layer3_outputs[1266] = layer2_outputs[2560];
    assign layer3_outputs[1267] = layer2_outputs[3142];
    assign layer3_outputs[1268] = ~(layer2_outputs[520]);
    assign layer3_outputs[1269] = ~((layer2_outputs[2284]) | (layer2_outputs[149]));
    assign layer3_outputs[1270] = (layer2_outputs[241]) & (layer2_outputs[3617]);
    assign layer3_outputs[1271] = ~(layer2_outputs[4665]);
    assign layer3_outputs[1272] = ~(layer2_outputs[3161]);
    assign layer3_outputs[1273] = (layer2_outputs[1003]) & ~(layer2_outputs[928]);
    assign layer3_outputs[1274] = layer2_outputs[1412];
    assign layer3_outputs[1275] = (layer2_outputs[2029]) & ~(layer2_outputs[1317]);
    assign layer3_outputs[1276] = layer2_outputs[4837];
    assign layer3_outputs[1277] = (layer2_outputs[5028]) | (layer2_outputs[3398]);
    assign layer3_outputs[1278] = (layer2_outputs[953]) & (layer2_outputs[2484]);
    assign layer3_outputs[1279] = (layer2_outputs[3286]) & ~(layer2_outputs[3679]);
    assign layer3_outputs[1280] = layer2_outputs[1859];
    assign layer3_outputs[1281] = (layer2_outputs[2602]) & ~(layer2_outputs[821]);
    assign layer3_outputs[1282] = ~((layer2_outputs[1606]) & (layer2_outputs[2001]));
    assign layer3_outputs[1283] = ~(layer2_outputs[3663]);
    assign layer3_outputs[1284] = ~(layer2_outputs[2981]);
    assign layer3_outputs[1285] = (layer2_outputs[4519]) & (layer2_outputs[1741]);
    assign layer3_outputs[1286] = ~(layer2_outputs[4088]);
    assign layer3_outputs[1287] = (layer2_outputs[2806]) & (layer2_outputs[4722]);
    assign layer3_outputs[1288] = 1'b1;
    assign layer3_outputs[1289] = ~((layer2_outputs[4318]) | (layer2_outputs[2924]));
    assign layer3_outputs[1290] = ~((layer2_outputs[102]) | (layer2_outputs[2966]));
    assign layer3_outputs[1291] = 1'b0;
    assign layer3_outputs[1292] = ~(layer2_outputs[2310]);
    assign layer3_outputs[1293] = 1'b1;
    assign layer3_outputs[1294] = 1'b1;
    assign layer3_outputs[1295] = layer2_outputs[4850];
    assign layer3_outputs[1296] = layer2_outputs[1829];
    assign layer3_outputs[1297] = (layer2_outputs[152]) & (layer2_outputs[1965]);
    assign layer3_outputs[1298] = (layer2_outputs[1408]) & ~(layer2_outputs[2406]);
    assign layer3_outputs[1299] = ~(layer2_outputs[2676]) | (layer2_outputs[1487]);
    assign layer3_outputs[1300] = (layer2_outputs[2877]) & ~(layer2_outputs[2872]);
    assign layer3_outputs[1301] = ~(layer2_outputs[798]);
    assign layer3_outputs[1302] = (layer2_outputs[2056]) & (layer2_outputs[1083]);
    assign layer3_outputs[1303] = ~(layer2_outputs[3549]) | (layer2_outputs[2357]);
    assign layer3_outputs[1304] = (layer2_outputs[113]) | (layer2_outputs[2199]);
    assign layer3_outputs[1305] = ~((layer2_outputs[635]) & (layer2_outputs[2785]));
    assign layer3_outputs[1306] = ~(layer2_outputs[172]);
    assign layer3_outputs[1307] = ~(layer2_outputs[2395]);
    assign layer3_outputs[1308] = layer2_outputs[2088];
    assign layer3_outputs[1309] = layer2_outputs[1250];
    assign layer3_outputs[1310] = ~(layer2_outputs[138]) | (layer2_outputs[804]);
    assign layer3_outputs[1311] = ~((layer2_outputs[3499]) & (layer2_outputs[3263]));
    assign layer3_outputs[1312] = ~(layer2_outputs[3282]);
    assign layer3_outputs[1313] = layer2_outputs[272];
    assign layer3_outputs[1314] = layer2_outputs[956];
    assign layer3_outputs[1315] = ~((layer2_outputs[1985]) | (layer2_outputs[1251]));
    assign layer3_outputs[1316] = layer2_outputs[2722];
    assign layer3_outputs[1317] = 1'b0;
    assign layer3_outputs[1318] = ~((layer2_outputs[524]) | (layer2_outputs[4298]));
    assign layer3_outputs[1319] = (layer2_outputs[2026]) & ~(layer2_outputs[4971]);
    assign layer3_outputs[1320] = (layer2_outputs[1915]) | (layer2_outputs[193]);
    assign layer3_outputs[1321] = ~(layer2_outputs[1445]) | (layer2_outputs[1188]);
    assign layer3_outputs[1322] = ~(layer2_outputs[231]) | (layer2_outputs[38]);
    assign layer3_outputs[1323] = (layer2_outputs[1414]) & (layer2_outputs[3086]);
    assign layer3_outputs[1324] = ~(layer2_outputs[3630]);
    assign layer3_outputs[1325] = (layer2_outputs[1833]) & ~(layer2_outputs[3709]);
    assign layer3_outputs[1326] = ~(layer2_outputs[3850]);
    assign layer3_outputs[1327] = (layer2_outputs[283]) & ~(layer2_outputs[2911]);
    assign layer3_outputs[1328] = ~(layer2_outputs[3799]);
    assign layer3_outputs[1329] = layer2_outputs[4436];
    assign layer3_outputs[1330] = ~((layer2_outputs[306]) | (layer2_outputs[1432]));
    assign layer3_outputs[1331] = (layer2_outputs[472]) | (layer2_outputs[16]);
    assign layer3_outputs[1332] = ~(layer2_outputs[5053]);
    assign layer3_outputs[1333] = ~(layer2_outputs[3500]);
    assign layer3_outputs[1334] = ~(layer2_outputs[3665]) | (layer2_outputs[4624]);
    assign layer3_outputs[1335] = (layer2_outputs[4294]) & ~(layer2_outputs[356]);
    assign layer3_outputs[1336] = ~(layer2_outputs[4448]);
    assign layer3_outputs[1337] = ~(layer2_outputs[1782]);
    assign layer3_outputs[1338] = ~(layer2_outputs[2024]);
    assign layer3_outputs[1339] = 1'b0;
    assign layer3_outputs[1340] = layer2_outputs[1966];
    assign layer3_outputs[1341] = ~(layer2_outputs[1552]);
    assign layer3_outputs[1342] = layer2_outputs[895];
    assign layer3_outputs[1343] = ~((layer2_outputs[3319]) & (layer2_outputs[3241]));
    assign layer3_outputs[1344] = layer2_outputs[5046];
    assign layer3_outputs[1345] = layer2_outputs[513];
    assign layer3_outputs[1346] = (layer2_outputs[1374]) & ~(layer2_outputs[3452]);
    assign layer3_outputs[1347] = ~(layer2_outputs[788]) | (layer2_outputs[846]);
    assign layer3_outputs[1348] = (layer2_outputs[566]) & (layer2_outputs[1086]);
    assign layer3_outputs[1349] = ~(layer2_outputs[1806]);
    assign layer3_outputs[1350] = layer2_outputs[940];
    assign layer3_outputs[1351] = ~(layer2_outputs[3081]);
    assign layer3_outputs[1352] = layer2_outputs[4616];
    assign layer3_outputs[1353] = 1'b1;
    assign layer3_outputs[1354] = 1'b0;
    assign layer3_outputs[1355] = layer2_outputs[2596];
    assign layer3_outputs[1356] = 1'b0;
    assign layer3_outputs[1357] = (layer2_outputs[2963]) & ~(layer2_outputs[2162]);
    assign layer3_outputs[1358] = ~(layer2_outputs[2754]);
    assign layer3_outputs[1359] = (layer2_outputs[2460]) & ~(layer2_outputs[1325]);
    assign layer3_outputs[1360] = layer2_outputs[3605];
    assign layer3_outputs[1361] = ~(layer2_outputs[466]);
    assign layer3_outputs[1362] = (layer2_outputs[2583]) & ~(layer2_outputs[2471]);
    assign layer3_outputs[1363] = ~(layer2_outputs[14]);
    assign layer3_outputs[1364] = ~(layer2_outputs[1114]);
    assign layer3_outputs[1365] = 1'b0;
    assign layer3_outputs[1366] = ~((layer2_outputs[3443]) & (layer2_outputs[3]));
    assign layer3_outputs[1367] = 1'b0;
    assign layer3_outputs[1368] = ~(layer2_outputs[3701]);
    assign layer3_outputs[1369] = ~(layer2_outputs[3663]);
    assign layer3_outputs[1370] = (layer2_outputs[2254]) | (layer2_outputs[2220]);
    assign layer3_outputs[1371] = 1'b0;
    assign layer3_outputs[1372] = layer2_outputs[3356];
    assign layer3_outputs[1373] = (layer2_outputs[2418]) & ~(layer2_outputs[2759]);
    assign layer3_outputs[1374] = 1'b0;
    assign layer3_outputs[1375] = 1'b0;
    assign layer3_outputs[1376] = 1'b1;
    assign layer3_outputs[1377] = (layer2_outputs[933]) & (layer2_outputs[3816]);
    assign layer3_outputs[1378] = 1'b0;
    assign layer3_outputs[1379] = layer2_outputs[722];
    assign layer3_outputs[1380] = ~((layer2_outputs[3180]) | (layer2_outputs[4444]));
    assign layer3_outputs[1381] = (layer2_outputs[2649]) ^ (layer2_outputs[2658]);
    assign layer3_outputs[1382] = ~((layer2_outputs[3103]) | (layer2_outputs[2178]));
    assign layer3_outputs[1383] = ~(layer2_outputs[2093]);
    assign layer3_outputs[1384] = 1'b1;
    assign layer3_outputs[1385] = 1'b1;
    assign layer3_outputs[1386] = layer2_outputs[996];
    assign layer3_outputs[1387] = ~(layer2_outputs[5106]);
    assign layer3_outputs[1388] = layer2_outputs[3424];
    assign layer3_outputs[1389] = 1'b0;
    assign layer3_outputs[1390] = ~((layer2_outputs[1957]) ^ (layer2_outputs[4932]));
    assign layer3_outputs[1391] = ~(layer2_outputs[1688]) | (layer2_outputs[1079]);
    assign layer3_outputs[1392] = layer2_outputs[5026];
    assign layer3_outputs[1393] = ~(layer2_outputs[3377]);
    assign layer3_outputs[1394] = ~(layer2_outputs[2708]) | (layer2_outputs[2333]);
    assign layer3_outputs[1395] = layer2_outputs[4081];
    assign layer3_outputs[1396] = ~(layer2_outputs[263]);
    assign layer3_outputs[1397] = 1'b0;
    assign layer3_outputs[1398] = (layer2_outputs[3431]) & (layer2_outputs[2652]);
    assign layer3_outputs[1399] = 1'b1;
    assign layer3_outputs[1400] = (layer2_outputs[4673]) & ~(layer2_outputs[3543]);
    assign layer3_outputs[1401] = 1'b1;
    assign layer3_outputs[1402] = layer2_outputs[3068];
    assign layer3_outputs[1403] = 1'b0;
    assign layer3_outputs[1404] = 1'b0;
    assign layer3_outputs[1405] = ~((layer2_outputs[3968]) & (layer2_outputs[4148]));
    assign layer3_outputs[1406] = ~(layer2_outputs[546]) | (layer2_outputs[1709]);
    assign layer3_outputs[1407] = ~(layer2_outputs[1721]);
    assign layer3_outputs[1408] = ~((layer2_outputs[2042]) & (layer2_outputs[1761]));
    assign layer3_outputs[1409] = (layer2_outputs[651]) & ~(layer2_outputs[4799]);
    assign layer3_outputs[1410] = 1'b1;
    assign layer3_outputs[1411] = layer2_outputs[756];
    assign layer3_outputs[1412] = ~((layer2_outputs[2367]) & (layer2_outputs[2880]));
    assign layer3_outputs[1413] = layer2_outputs[3141];
    assign layer3_outputs[1414] = ~((layer2_outputs[614]) ^ (layer2_outputs[3608]));
    assign layer3_outputs[1415] = ~((layer2_outputs[2617]) ^ (layer2_outputs[564]));
    assign layer3_outputs[1416] = 1'b1;
    assign layer3_outputs[1417] = layer2_outputs[2922];
    assign layer3_outputs[1418] = ~(layer2_outputs[4215]);
    assign layer3_outputs[1419] = ~(layer2_outputs[1165]) | (layer2_outputs[4005]);
    assign layer3_outputs[1420] = (layer2_outputs[2949]) & ~(layer2_outputs[343]);
    assign layer3_outputs[1421] = (layer2_outputs[2128]) & (layer2_outputs[4508]);
    assign layer3_outputs[1422] = (layer2_outputs[194]) & ~(layer2_outputs[1949]);
    assign layer3_outputs[1423] = ~((layer2_outputs[4295]) & (layer2_outputs[3544]));
    assign layer3_outputs[1424] = 1'b1;
    assign layer3_outputs[1425] = ~(layer2_outputs[2565]) | (layer2_outputs[517]);
    assign layer3_outputs[1426] = ~((layer2_outputs[3448]) | (layer2_outputs[1274]));
    assign layer3_outputs[1427] = (layer2_outputs[4106]) & ~(layer2_outputs[3529]);
    assign layer3_outputs[1428] = ~(layer2_outputs[2629]) | (layer2_outputs[3892]);
    assign layer3_outputs[1429] = ~(layer2_outputs[1554]);
    assign layer3_outputs[1430] = layer2_outputs[4186];
    assign layer3_outputs[1431] = ~((layer2_outputs[5031]) & (layer2_outputs[3061]));
    assign layer3_outputs[1432] = (layer2_outputs[2661]) & ~(layer2_outputs[273]);
    assign layer3_outputs[1433] = ~((layer2_outputs[2372]) & (layer2_outputs[4305]));
    assign layer3_outputs[1434] = ~(layer2_outputs[2809]);
    assign layer3_outputs[1435] = ~((layer2_outputs[3470]) ^ (layer2_outputs[1911]));
    assign layer3_outputs[1436] = ~(layer2_outputs[2619]);
    assign layer3_outputs[1437] = ~(layer2_outputs[3139]) | (layer2_outputs[3372]);
    assign layer3_outputs[1438] = ~(layer2_outputs[3090]);
    assign layer3_outputs[1439] = layer2_outputs[4047];
    assign layer3_outputs[1440] = ~(layer2_outputs[463]) | (layer2_outputs[2109]);
    assign layer3_outputs[1441] = ~(layer2_outputs[2741]);
    assign layer3_outputs[1442] = ~(layer2_outputs[119]);
    assign layer3_outputs[1443] = layer2_outputs[4360];
    assign layer3_outputs[1444] = 1'b1;
    assign layer3_outputs[1445] = ~((layer2_outputs[858]) & (layer2_outputs[1937]));
    assign layer3_outputs[1446] = ~((layer2_outputs[4435]) ^ (layer2_outputs[2275]));
    assign layer3_outputs[1447] = 1'b1;
    assign layer3_outputs[1448] = layer2_outputs[3449];
    assign layer3_outputs[1449] = layer2_outputs[1725];
    assign layer3_outputs[1450] = ~((layer2_outputs[4877]) & (layer2_outputs[5114]));
    assign layer3_outputs[1451] = ~(layer2_outputs[1114]);
    assign layer3_outputs[1452] = ~((layer2_outputs[3174]) | (layer2_outputs[2923]));
    assign layer3_outputs[1453] = layer2_outputs[2305];
    assign layer3_outputs[1454] = (layer2_outputs[1599]) | (layer2_outputs[4824]);
    assign layer3_outputs[1455] = (layer2_outputs[4609]) ^ (layer2_outputs[1777]);
    assign layer3_outputs[1456] = (layer2_outputs[3725]) | (layer2_outputs[438]);
    assign layer3_outputs[1457] = ~(layer2_outputs[2639]) | (layer2_outputs[1511]);
    assign layer3_outputs[1458] = 1'b1;
    assign layer3_outputs[1459] = ~(layer2_outputs[3888]) | (layer2_outputs[3300]);
    assign layer3_outputs[1460] = ~(layer2_outputs[3318]);
    assign layer3_outputs[1461] = ~(layer2_outputs[1902]) | (layer2_outputs[3242]);
    assign layer3_outputs[1462] = ~((layer2_outputs[3433]) & (layer2_outputs[2582]));
    assign layer3_outputs[1463] = ~(layer2_outputs[1915]);
    assign layer3_outputs[1464] = (layer2_outputs[3847]) & ~(layer2_outputs[234]);
    assign layer3_outputs[1465] = 1'b1;
    assign layer3_outputs[1466] = layer2_outputs[4952];
    assign layer3_outputs[1467] = (layer2_outputs[2977]) & ~(layer2_outputs[3912]);
    assign layer3_outputs[1468] = ~(layer2_outputs[1569]);
    assign layer3_outputs[1469] = layer2_outputs[228];
    assign layer3_outputs[1470] = (layer2_outputs[1377]) & ~(layer2_outputs[3871]);
    assign layer3_outputs[1471] = ~(layer2_outputs[1737]) | (layer2_outputs[1624]);
    assign layer3_outputs[1472] = (layer2_outputs[3621]) & ~(layer2_outputs[1179]);
    assign layer3_outputs[1473] = ~(layer2_outputs[1124]);
    assign layer3_outputs[1474] = (layer2_outputs[2086]) & ~(layer2_outputs[527]);
    assign layer3_outputs[1475] = (layer2_outputs[3610]) & (layer2_outputs[3972]);
    assign layer3_outputs[1476] = layer2_outputs[887];
    assign layer3_outputs[1477] = ~(layer2_outputs[4000]);
    assign layer3_outputs[1478] = layer2_outputs[3157];
    assign layer3_outputs[1479] = ~(layer2_outputs[3618]) | (layer2_outputs[1838]);
    assign layer3_outputs[1480] = ~(layer2_outputs[3212]) | (layer2_outputs[129]);
    assign layer3_outputs[1481] = ~(layer2_outputs[4368]);
    assign layer3_outputs[1482] = layer2_outputs[2080];
    assign layer3_outputs[1483] = (layer2_outputs[2925]) & (layer2_outputs[3938]);
    assign layer3_outputs[1484] = ~(layer2_outputs[2441]) | (layer2_outputs[4919]);
    assign layer3_outputs[1485] = ~((layer2_outputs[3084]) & (layer2_outputs[1085]));
    assign layer3_outputs[1486] = 1'b1;
    assign layer3_outputs[1487] = 1'b0;
    assign layer3_outputs[1488] = (layer2_outputs[186]) & ~(layer2_outputs[1451]);
    assign layer3_outputs[1489] = ~(layer2_outputs[2755]) | (layer2_outputs[4625]);
    assign layer3_outputs[1490] = ~(layer2_outputs[169]);
    assign layer3_outputs[1491] = ~((layer2_outputs[1622]) & (layer2_outputs[1479]));
    assign layer3_outputs[1492] = (layer2_outputs[3461]) & ~(layer2_outputs[1697]);
    assign layer3_outputs[1493] = (layer2_outputs[3896]) & ~(layer2_outputs[4323]);
    assign layer3_outputs[1494] = (layer2_outputs[3463]) & (layer2_outputs[3956]);
    assign layer3_outputs[1495] = 1'b0;
    assign layer3_outputs[1496] = layer2_outputs[724];
    assign layer3_outputs[1497] = layer2_outputs[432];
    assign layer3_outputs[1498] = layer2_outputs[2452];
    assign layer3_outputs[1499] = layer2_outputs[3186];
    assign layer3_outputs[1500] = ~(layer2_outputs[466]) | (layer2_outputs[3052]);
    assign layer3_outputs[1501] = layer2_outputs[399];
    assign layer3_outputs[1502] = (layer2_outputs[5098]) & ~(layer2_outputs[4552]);
    assign layer3_outputs[1503] = (layer2_outputs[13]) & ~(layer2_outputs[4445]);
    assign layer3_outputs[1504] = (layer2_outputs[2239]) & ~(layer2_outputs[3575]);
    assign layer3_outputs[1505] = 1'b0;
    assign layer3_outputs[1506] = layer2_outputs[3770];
    assign layer3_outputs[1507] = layer2_outputs[1408];
    assign layer3_outputs[1508] = (layer2_outputs[3168]) & ~(layer2_outputs[2089]);
    assign layer3_outputs[1509] = (layer2_outputs[1486]) & (layer2_outputs[3189]);
    assign layer3_outputs[1510] = ~(layer2_outputs[4127]) | (layer2_outputs[4145]);
    assign layer3_outputs[1511] = layer2_outputs[1569];
    assign layer3_outputs[1512] = ~((layer2_outputs[2802]) & (layer2_outputs[2771]));
    assign layer3_outputs[1513] = ~((layer2_outputs[4382]) & (layer2_outputs[1567]));
    assign layer3_outputs[1514] = (layer2_outputs[973]) & ~(layer2_outputs[3244]);
    assign layer3_outputs[1515] = (layer2_outputs[2381]) & ~(layer2_outputs[429]);
    assign layer3_outputs[1516] = ~(layer2_outputs[3709]);
    assign layer3_outputs[1517] = (layer2_outputs[3607]) | (layer2_outputs[5000]);
    assign layer3_outputs[1518] = ~(layer2_outputs[3477]);
    assign layer3_outputs[1519] = layer2_outputs[1238];
    assign layer3_outputs[1520] = ~(layer2_outputs[2472]);
    assign layer3_outputs[1521] = (layer2_outputs[3271]) & ~(layer2_outputs[3553]);
    assign layer3_outputs[1522] = (layer2_outputs[1388]) & ~(layer2_outputs[4454]);
    assign layer3_outputs[1523] = 1'b1;
    assign layer3_outputs[1524] = layer2_outputs[945];
    assign layer3_outputs[1525] = ~(layer2_outputs[319]);
    assign layer3_outputs[1526] = 1'b1;
    assign layer3_outputs[1527] = layer2_outputs[459];
    assign layer3_outputs[1528] = layer2_outputs[388];
    assign layer3_outputs[1529] = (layer2_outputs[3592]) & ~(layer2_outputs[3317]);
    assign layer3_outputs[1530] = ~(layer2_outputs[229]);
    assign layer3_outputs[1531] = layer2_outputs[5113];
    assign layer3_outputs[1532] = ~((layer2_outputs[1588]) ^ (layer2_outputs[1083]));
    assign layer3_outputs[1533] = layer2_outputs[3770];
    assign layer3_outputs[1534] = ~((layer2_outputs[218]) & (layer2_outputs[3379]));
    assign layer3_outputs[1535] = ~(layer2_outputs[3653]);
    assign layer3_outputs[1536] = (layer2_outputs[2795]) & ~(layer2_outputs[1768]);
    assign layer3_outputs[1537] = ~((layer2_outputs[2334]) & (layer2_outputs[4301]));
    assign layer3_outputs[1538] = (layer2_outputs[3817]) & (layer2_outputs[663]);
    assign layer3_outputs[1539] = (layer2_outputs[4541]) & (layer2_outputs[861]);
    assign layer3_outputs[1540] = ~(layer2_outputs[4172]);
    assign layer3_outputs[1541] = ~((layer2_outputs[3487]) | (layer2_outputs[1572]));
    assign layer3_outputs[1542] = (layer2_outputs[401]) & ~(layer2_outputs[4484]);
    assign layer3_outputs[1543] = layer2_outputs[1976];
    assign layer3_outputs[1544] = 1'b0;
    assign layer3_outputs[1545] = 1'b0;
    assign layer3_outputs[1546] = (layer2_outputs[3167]) & ~(layer2_outputs[2537]);
    assign layer3_outputs[1547] = layer2_outputs[3622];
    assign layer3_outputs[1548] = ~((layer2_outputs[3955]) | (layer2_outputs[471]));
    assign layer3_outputs[1549] = ~((layer2_outputs[2252]) ^ (layer2_outputs[4962]));
    assign layer3_outputs[1550] = layer2_outputs[829];
    assign layer3_outputs[1551] = ~(layer2_outputs[3547]) | (layer2_outputs[2213]);
    assign layer3_outputs[1552] = ~(layer2_outputs[18]);
    assign layer3_outputs[1553] = ~(layer2_outputs[4499]);
    assign layer3_outputs[1554] = layer2_outputs[1089];
    assign layer3_outputs[1555] = (layer2_outputs[3967]) | (layer2_outputs[4138]);
    assign layer3_outputs[1556] = 1'b0;
    assign layer3_outputs[1557] = (layer2_outputs[3297]) & (layer2_outputs[2230]);
    assign layer3_outputs[1558] = (layer2_outputs[5043]) & ~(layer2_outputs[1520]);
    assign layer3_outputs[1559] = (layer2_outputs[3192]) & ~(layer2_outputs[3335]);
    assign layer3_outputs[1560] = (layer2_outputs[2313]) & ~(layer2_outputs[2849]);
    assign layer3_outputs[1561] = ~(layer2_outputs[4096]) | (layer2_outputs[2002]);
    assign layer3_outputs[1562] = ~((layer2_outputs[1263]) ^ (layer2_outputs[1378]));
    assign layer3_outputs[1563] = (layer2_outputs[4323]) & ~(layer2_outputs[453]);
    assign layer3_outputs[1564] = ~(layer2_outputs[4355]) | (layer2_outputs[1685]);
    assign layer3_outputs[1565] = ~(layer2_outputs[2450]);
    assign layer3_outputs[1566] = ~((layer2_outputs[3456]) | (layer2_outputs[3807]));
    assign layer3_outputs[1567] = ~((layer2_outputs[3145]) | (layer2_outputs[417]));
    assign layer3_outputs[1568] = (layer2_outputs[4432]) & ~(layer2_outputs[1277]);
    assign layer3_outputs[1569] = ~(layer2_outputs[1484]) | (layer2_outputs[4313]);
    assign layer3_outputs[1570] = ~((layer2_outputs[3684]) | (layer2_outputs[450]));
    assign layer3_outputs[1571] = (layer2_outputs[4638]) | (layer2_outputs[1689]);
    assign layer3_outputs[1572] = layer2_outputs[1843];
    assign layer3_outputs[1573] = 1'b0;
    assign layer3_outputs[1574] = layer2_outputs[153];
    assign layer3_outputs[1575] = (layer2_outputs[2785]) & ~(layer2_outputs[1997]);
    assign layer3_outputs[1576] = layer2_outputs[199];
    assign layer3_outputs[1577] = layer2_outputs[308];
    assign layer3_outputs[1578] = 1'b1;
    assign layer3_outputs[1579] = ~(layer2_outputs[2410]);
    assign layer3_outputs[1580] = layer2_outputs[353];
    assign layer3_outputs[1581] = (layer2_outputs[4095]) | (layer2_outputs[4209]);
    assign layer3_outputs[1582] = ~((layer2_outputs[674]) | (layer2_outputs[1943]));
    assign layer3_outputs[1583] = ~(layer2_outputs[1711]);
    assign layer3_outputs[1584] = (layer2_outputs[1380]) & (layer2_outputs[2404]);
    assign layer3_outputs[1585] = (layer2_outputs[481]) & ~(layer2_outputs[3322]);
    assign layer3_outputs[1586] = ~(layer2_outputs[1751]) | (layer2_outputs[2982]);
    assign layer3_outputs[1587] = layer2_outputs[4997];
    assign layer3_outputs[1588] = ~((layer2_outputs[2082]) | (layer2_outputs[634]));
    assign layer3_outputs[1589] = ~(layer2_outputs[1563]);
    assign layer3_outputs[1590] = layer2_outputs[2075];
    assign layer3_outputs[1591] = layer2_outputs[2651];
    assign layer3_outputs[1592] = ~((layer2_outputs[1835]) & (layer2_outputs[530]));
    assign layer3_outputs[1593] = 1'b1;
    assign layer3_outputs[1594] = layer2_outputs[4626];
    assign layer3_outputs[1595] = layer2_outputs[1150];
    assign layer3_outputs[1596] = ~(layer2_outputs[1402]) | (layer2_outputs[4881]);
    assign layer3_outputs[1597] = (layer2_outputs[4939]) ^ (layer2_outputs[854]);
    assign layer3_outputs[1598] = ~(layer2_outputs[869]) | (layer2_outputs[2687]);
    assign layer3_outputs[1599] = ~(layer2_outputs[1667]) | (layer2_outputs[3414]);
    assign layer3_outputs[1600] = (layer2_outputs[3348]) | (layer2_outputs[4117]);
    assign layer3_outputs[1601] = (layer2_outputs[3269]) | (layer2_outputs[1204]);
    assign layer3_outputs[1602] = ~((layer2_outputs[4225]) ^ (layer2_outputs[2763]));
    assign layer3_outputs[1603] = ~(layer2_outputs[2006]);
    assign layer3_outputs[1604] = ~(layer2_outputs[2126]);
    assign layer3_outputs[1605] = (layer2_outputs[3789]) & ~(layer2_outputs[4351]);
    assign layer3_outputs[1606] = ~(layer2_outputs[4709]) | (layer2_outputs[3672]);
    assign layer3_outputs[1607] = ~(layer2_outputs[4982]);
    assign layer3_outputs[1608] = layer2_outputs[2513];
    assign layer3_outputs[1609] = (layer2_outputs[4352]) | (layer2_outputs[3146]);
    assign layer3_outputs[1610] = ~(layer2_outputs[2067]);
    assign layer3_outputs[1611] = ~(layer2_outputs[2107]);
    assign layer3_outputs[1612] = layer2_outputs[2735];
    assign layer3_outputs[1613] = (layer2_outputs[2273]) | (layer2_outputs[3220]);
    assign layer3_outputs[1614] = (layer2_outputs[2000]) & (layer2_outputs[4666]);
    assign layer3_outputs[1615] = (layer2_outputs[1118]) ^ (layer2_outputs[3031]);
    assign layer3_outputs[1616] = ~(layer2_outputs[3038]);
    assign layer3_outputs[1617] = ~(layer2_outputs[809]);
    assign layer3_outputs[1618] = (layer2_outputs[61]) & (layer2_outputs[412]);
    assign layer3_outputs[1619] = (layer2_outputs[1978]) & (layer2_outputs[4200]);
    assign layer3_outputs[1620] = ~(layer2_outputs[1141]);
    assign layer3_outputs[1621] = layer2_outputs[175];
    assign layer3_outputs[1622] = ~(layer2_outputs[2053]) | (layer2_outputs[4807]);
    assign layer3_outputs[1623] = ~((layer2_outputs[3230]) | (layer2_outputs[2633]));
    assign layer3_outputs[1624] = (layer2_outputs[2204]) & ~(layer2_outputs[2512]);
    assign layer3_outputs[1625] = ~((layer2_outputs[2163]) & (layer2_outputs[3337]));
    assign layer3_outputs[1626] = ~((layer2_outputs[4152]) | (layer2_outputs[2802]));
    assign layer3_outputs[1627] = (layer2_outputs[4849]) & (layer2_outputs[3103]);
    assign layer3_outputs[1628] = (layer2_outputs[4838]) | (layer2_outputs[413]);
    assign layer3_outputs[1629] = 1'b0;
    assign layer3_outputs[1630] = layer2_outputs[855];
    assign layer3_outputs[1631] = ~(layer2_outputs[2829]) | (layer2_outputs[1996]);
    assign layer3_outputs[1632] = ~(layer2_outputs[2099]);
    assign layer3_outputs[1633] = ~(layer2_outputs[1188]);
    assign layer3_outputs[1634] = 1'b1;
    assign layer3_outputs[1635] = layer2_outputs[512];
    assign layer3_outputs[1636] = layer2_outputs[2905];
    assign layer3_outputs[1637] = ~(layer2_outputs[626]);
    assign layer3_outputs[1638] = ~(layer2_outputs[3283]);
    assign layer3_outputs[1639] = 1'b1;
    assign layer3_outputs[1640] = (layer2_outputs[214]) | (layer2_outputs[668]);
    assign layer3_outputs[1641] = ~(layer2_outputs[3693]) | (layer2_outputs[3879]);
    assign layer3_outputs[1642] = ~((layer2_outputs[3410]) | (layer2_outputs[1517]));
    assign layer3_outputs[1643] = (layer2_outputs[1037]) | (layer2_outputs[2303]);
    assign layer3_outputs[1644] = (layer2_outputs[4856]) & ~(layer2_outputs[1098]);
    assign layer3_outputs[1645] = 1'b0;
    assign layer3_outputs[1646] = (layer2_outputs[2509]) | (layer2_outputs[3908]);
    assign layer3_outputs[1647] = ~(layer2_outputs[3478]) | (layer2_outputs[2255]);
    assign layer3_outputs[1648] = (layer2_outputs[177]) ^ (layer2_outputs[3527]);
    assign layer3_outputs[1649] = ~(layer2_outputs[4691]);
    assign layer3_outputs[1650] = layer2_outputs[3795];
    assign layer3_outputs[1651] = ~(layer2_outputs[616]) | (layer2_outputs[1120]);
    assign layer3_outputs[1652] = ~(layer2_outputs[777]);
    assign layer3_outputs[1653] = ~(layer2_outputs[3135]) | (layer2_outputs[1698]);
    assign layer3_outputs[1654] = ~((layer2_outputs[963]) ^ (layer2_outputs[4131]));
    assign layer3_outputs[1655] = 1'b0;
    assign layer3_outputs[1656] = ~((layer2_outputs[25]) & (layer2_outputs[1077]));
    assign layer3_outputs[1657] = (layer2_outputs[2805]) & ~(layer2_outputs[4958]);
    assign layer3_outputs[1658] = layer2_outputs[3102];
    assign layer3_outputs[1659] = 1'b1;
    assign layer3_outputs[1660] = ~((layer2_outputs[2300]) & (layer2_outputs[4899]));
    assign layer3_outputs[1661] = ~(layer2_outputs[1795]);
    assign layer3_outputs[1662] = (layer2_outputs[2223]) & ~(layer2_outputs[1761]);
    assign layer3_outputs[1663] = ~(layer2_outputs[2155]) | (layer2_outputs[3640]);
    assign layer3_outputs[1664] = ~(layer2_outputs[446]) | (layer2_outputs[320]);
    assign layer3_outputs[1665] = 1'b1;
    assign layer3_outputs[1666] = 1'b1;
    assign layer3_outputs[1667] = (layer2_outputs[740]) & ~(layer2_outputs[4757]);
    assign layer3_outputs[1668] = ~(layer2_outputs[655]);
    assign layer3_outputs[1669] = ~(layer2_outputs[2134]);
    assign layer3_outputs[1670] = ~(layer2_outputs[117]);
    assign layer3_outputs[1671] = ~((layer2_outputs[1787]) ^ (layer2_outputs[247]));
    assign layer3_outputs[1672] = (layer2_outputs[430]) & (layer2_outputs[473]);
    assign layer3_outputs[1673] = ~(layer2_outputs[2005]);
    assign layer3_outputs[1674] = ~(layer2_outputs[1476]) | (layer2_outputs[4139]);
    assign layer3_outputs[1675] = (layer2_outputs[4766]) | (layer2_outputs[3240]);
    assign layer3_outputs[1676] = ~(layer2_outputs[3412]);
    assign layer3_outputs[1677] = layer2_outputs[1089];
    assign layer3_outputs[1678] = ~((layer2_outputs[4413]) ^ (layer2_outputs[841]));
    assign layer3_outputs[1679] = (layer2_outputs[3520]) & (layer2_outputs[1513]);
    assign layer3_outputs[1680] = ~(layer2_outputs[106]);
    assign layer3_outputs[1681] = ~(layer2_outputs[351]);
    assign layer3_outputs[1682] = layer2_outputs[999];
    assign layer3_outputs[1683] = ~(layer2_outputs[4832]) | (layer2_outputs[1673]);
    assign layer3_outputs[1684] = layer2_outputs[3246];
    assign layer3_outputs[1685] = (layer2_outputs[492]) & ~(layer2_outputs[4728]);
    assign layer3_outputs[1686] = (layer2_outputs[1508]) & ~(layer2_outputs[1957]);
    assign layer3_outputs[1687] = layer2_outputs[686];
    assign layer3_outputs[1688] = ~(layer2_outputs[4226]);
    assign layer3_outputs[1689] = ~(layer2_outputs[739]);
    assign layer3_outputs[1690] = (layer2_outputs[2132]) & ~(layer2_outputs[3822]);
    assign layer3_outputs[1691] = (layer2_outputs[596]) | (layer2_outputs[2794]);
    assign layer3_outputs[1692] = ~(layer2_outputs[2964]) | (layer2_outputs[810]);
    assign layer3_outputs[1693] = ~(layer2_outputs[2875]) | (layer2_outputs[2640]);
    assign layer3_outputs[1694] = ~((layer2_outputs[2553]) | (layer2_outputs[4073]));
    assign layer3_outputs[1695] = ~((layer2_outputs[690]) | (layer2_outputs[2529]));
    assign layer3_outputs[1696] = ~(layer2_outputs[4158]) | (layer2_outputs[4833]);
    assign layer3_outputs[1697] = layer2_outputs[3643];
    assign layer3_outputs[1698] = ~(layer2_outputs[3122]);
    assign layer3_outputs[1699] = layer2_outputs[772];
    assign layer3_outputs[1700] = ~(layer2_outputs[428]) | (layer2_outputs[4916]);
    assign layer3_outputs[1701] = ~(layer2_outputs[3404]) | (layer2_outputs[3671]);
    assign layer3_outputs[1702] = (layer2_outputs[1620]) & (layer2_outputs[2048]);
    assign layer3_outputs[1703] = layer2_outputs[134];
    assign layer3_outputs[1704] = (layer2_outputs[5018]) & ~(layer2_outputs[1503]);
    assign layer3_outputs[1705] = ~(layer2_outputs[3904]);
    assign layer3_outputs[1706] = layer2_outputs[3043];
    assign layer3_outputs[1707] = ~(layer2_outputs[3660]);
    assign layer3_outputs[1708] = layer2_outputs[2766];
    assign layer3_outputs[1709] = layer2_outputs[1446];
    assign layer3_outputs[1710] = ~(layer2_outputs[3589]);
    assign layer3_outputs[1711] = ~(layer2_outputs[3097]) | (layer2_outputs[592]);
    assign layer3_outputs[1712] = ~(layer2_outputs[2710]);
    assign layer3_outputs[1713] = ~(layer2_outputs[300]);
    assign layer3_outputs[1714] = (layer2_outputs[1999]) & ~(layer2_outputs[4199]);
    assign layer3_outputs[1715] = layer2_outputs[3773];
    assign layer3_outputs[1716] = 1'b1;
    assign layer3_outputs[1717] = (layer2_outputs[4193]) & ~(layer2_outputs[161]);
    assign layer3_outputs[1718] = ~(layer2_outputs[3841]) | (layer2_outputs[5080]);
    assign layer3_outputs[1719] = (layer2_outputs[4159]) | (layer2_outputs[1926]);
    assign layer3_outputs[1720] = ~(layer2_outputs[4860]);
    assign layer3_outputs[1721] = ~(layer2_outputs[3307]) | (layer2_outputs[4426]);
    assign layer3_outputs[1722] = 1'b0;
    assign layer3_outputs[1723] = ~(layer2_outputs[4101]) | (layer2_outputs[3389]);
    assign layer3_outputs[1724] = ~((layer2_outputs[4223]) | (layer2_outputs[781]));
    assign layer3_outputs[1725] = ~(layer2_outputs[3875]);
    assign layer3_outputs[1726] = (layer2_outputs[1048]) & ~(layer2_outputs[4914]);
    assign layer3_outputs[1727] = ~(layer2_outputs[1607]);
    assign layer3_outputs[1728] = ~(layer2_outputs[3417]);
    assign layer3_outputs[1729] = (layer2_outputs[4759]) ^ (layer2_outputs[1870]);
    assign layer3_outputs[1730] = (layer2_outputs[4579]) ^ (layer2_outputs[170]);
    assign layer3_outputs[1731] = (layer2_outputs[169]) & ~(layer2_outputs[2009]);
    assign layer3_outputs[1732] = ~(layer2_outputs[2761]) | (layer2_outputs[1675]);
    assign layer3_outputs[1733] = 1'b1;
    assign layer3_outputs[1734] = (layer2_outputs[3888]) & ~(layer2_outputs[905]);
    assign layer3_outputs[1735] = (layer2_outputs[2616]) & ~(layer2_outputs[2154]);
    assign layer3_outputs[1736] = layer2_outputs[4853];
    assign layer3_outputs[1737] = (layer2_outputs[242]) & ~(layer2_outputs[1580]);
    assign layer3_outputs[1738] = layer2_outputs[4633];
    assign layer3_outputs[1739] = (layer2_outputs[3513]) & (layer2_outputs[1483]);
    assign layer3_outputs[1740] = ~(layer2_outputs[2543]) | (layer2_outputs[1206]);
    assign layer3_outputs[1741] = 1'b0;
    assign layer3_outputs[1742] = 1'b0;
    assign layer3_outputs[1743] = (layer2_outputs[4660]) ^ (layer2_outputs[3634]);
    assign layer3_outputs[1744] = (layer2_outputs[1989]) & ~(layer2_outputs[4511]);
    assign layer3_outputs[1745] = 1'b0;
    assign layer3_outputs[1746] = ~((layer2_outputs[882]) & (layer2_outputs[4514]));
    assign layer3_outputs[1747] = ~(layer2_outputs[1873]) | (layer2_outputs[2165]);
    assign layer3_outputs[1748] = 1'b1;
    assign layer3_outputs[1749] = layer2_outputs[2492];
    assign layer3_outputs[1750] = (layer2_outputs[5056]) & (layer2_outputs[3521]);
    assign layer3_outputs[1751] = ~(layer2_outputs[3292]);
    assign layer3_outputs[1752] = ~(layer2_outputs[2506]) | (layer2_outputs[5070]);
    assign layer3_outputs[1753] = 1'b0;
    assign layer3_outputs[1754] = (layer2_outputs[4935]) & ~(layer2_outputs[1473]);
    assign layer3_outputs[1755] = layer2_outputs[2926];
    assign layer3_outputs[1756] = ~(layer2_outputs[3680]);
    assign layer3_outputs[1757] = layer2_outputs[2701];
    assign layer3_outputs[1758] = ~(layer2_outputs[1535]);
    assign layer3_outputs[1759] = 1'b1;
    assign layer3_outputs[1760] = ~(layer2_outputs[1071]);
    assign layer3_outputs[1761] = layer2_outputs[3897];
    assign layer3_outputs[1762] = ~((layer2_outputs[3403]) & (layer2_outputs[4037]));
    assign layer3_outputs[1763] = ~((layer2_outputs[3033]) | (layer2_outputs[4170]));
    assign layer3_outputs[1764] = 1'b0;
    assign layer3_outputs[1765] = (layer2_outputs[1187]) & (layer2_outputs[3687]);
    assign layer3_outputs[1766] = 1'b0;
    assign layer3_outputs[1767] = layer2_outputs[4059];
    assign layer3_outputs[1768] = (layer2_outputs[1593]) & ~(layer2_outputs[3321]);
    assign layer3_outputs[1769] = (layer2_outputs[814]) & ~(layer2_outputs[4528]);
    assign layer3_outputs[1770] = ~(layer2_outputs[1639]);
    assign layer3_outputs[1771] = layer2_outputs[2616];
    assign layer3_outputs[1772] = layer2_outputs[1225];
    assign layer3_outputs[1773] = layer2_outputs[4248];
    assign layer3_outputs[1774] = (layer2_outputs[1066]) & ~(layer2_outputs[5066]);
    assign layer3_outputs[1775] = (layer2_outputs[292]) | (layer2_outputs[1760]);
    assign layer3_outputs[1776] = 1'b1;
    assign layer3_outputs[1777] = ~(layer2_outputs[427]);
    assign layer3_outputs[1778] = (layer2_outputs[683]) ^ (layer2_outputs[1747]);
    assign layer3_outputs[1779] = ~((layer2_outputs[3546]) | (layer2_outputs[1946]));
    assign layer3_outputs[1780] = ~(layer2_outputs[571]);
    assign layer3_outputs[1781] = layer2_outputs[4495];
    assign layer3_outputs[1782] = ~(layer2_outputs[1004]);
    assign layer3_outputs[1783] = ~((layer2_outputs[2189]) ^ (layer2_outputs[1974]));
    assign layer3_outputs[1784] = (layer2_outputs[3699]) | (layer2_outputs[4903]);
    assign layer3_outputs[1785] = (layer2_outputs[1713]) & ~(layer2_outputs[4283]);
    assign layer3_outputs[1786] = ~(layer2_outputs[218]);
    assign layer3_outputs[1787] = ~(layer2_outputs[586]) | (layer2_outputs[1846]);
    assign layer3_outputs[1788] = ~((layer2_outputs[5102]) & (layer2_outputs[3385]));
    assign layer3_outputs[1789] = (layer2_outputs[3193]) & (layer2_outputs[101]);
    assign layer3_outputs[1790] = ~((layer2_outputs[2148]) ^ (layer2_outputs[3636]));
    assign layer3_outputs[1791] = ~(layer2_outputs[4891]) | (layer2_outputs[3007]);
    assign layer3_outputs[1792] = ~(layer2_outputs[450]);
    assign layer3_outputs[1793] = layer2_outputs[2179];
    assign layer3_outputs[1794] = ~(layer2_outputs[889]);
    assign layer3_outputs[1795] = (layer2_outputs[3457]) & (layer2_outputs[2787]);
    assign layer3_outputs[1796] = layer2_outputs[3725];
    assign layer3_outputs[1797] = (layer2_outputs[2455]) & (layer2_outputs[4222]);
    assign layer3_outputs[1798] = layer2_outputs[1773];
    assign layer3_outputs[1799] = ~(layer2_outputs[3173]) | (layer2_outputs[4603]);
    assign layer3_outputs[1800] = ~(layer2_outputs[3452]) | (layer2_outputs[4957]);
    assign layer3_outputs[1801] = ~(layer2_outputs[2636]);
    assign layer3_outputs[1802] = layer2_outputs[3565];
    assign layer3_outputs[1803] = (layer2_outputs[4141]) & ~(layer2_outputs[4222]);
    assign layer3_outputs[1804] = 1'b0;
    assign layer3_outputs[1805] = ~(layer2_outputs[1452]) | (layer2_outputs[4955]);
    assign layer3_outputs[1806] = layer2_outputs[587];
    assign layer3_outputs[1807] = layer2_outputs[1516];
    assign layer3_outputs[1808] = ~((layer2_outputs[1062]) & (layer2_outputs[4589]));
    assign layer3_outputs[1809] = ~(layer2_outputs[2770]) | (layer2_outputs[4740]);
    assign layer3_outputs[1810] = layer2_outputs[1107];
    assign layer3_outputs[1811] = ~((layer2_outputs[4775]) | (layer2_outputs[2817]));
    assign layer3_outputs[1812] = (layer2_outputs[2100]) | (layer2_outputs[3992]);
    assign layer3_outputs[1813] = (layer2_outputs[2390]) & ~(layer2_outputs[4976]);
    assign layer3_outputs[1814] = (layer2_outputs[114]) & ~(layer2_outputs[3957]);
    assign layer3_outputs[1815] = 1'b0;
    assign layer3_outputs[1816] = ~(layer2_outputs[486]);
    assign layer3_outputs[1817] = (layer2_outputs[3324]) & ~(layer2_outputs[15]);
    assign layer3_outputs[1818] = (layer2_outputs[3068]) & (layer2_outputs[202]);
    assign layer3_outputs[1819] = 1'b1;
    assign layer3_outputs[1820] = ~(layer2_outputs[4785]) | (layer2_outputs[3879]);
    assign layer3_outputs[1821] = (layer2_outputs[3774]) ^ (layer2_outputs[4546]);
    assign layer3_outputs[1822] = ~((layer2_outputs[329]) ^ (layer2_outputs[2841]));
    assign layer3_outputs[1823] = ~(layer2_outputs[3206]);
    assign layer3_outputs[1824] = (layer2_outputs[4860]) & ~(layer2_outputs[1192]);
    assign layer3_outputs[1825] = ~(layer2_outputs[942]) | (layer2_outputs[4232]);
    assign layer3_outputs[1826] = ~(layer2_outputs[4810]);
    assign layer3_outputs[1827] = 1'b0;
    assign layer3_outputs[1828] = (layer2_outputs[3373]) | (layer2_outputs[4330]);
    assign layer3_outputs[1829] = ~(layer2_outputs[764]);
    assign layer3_outputs[1830] = 1'b0;
    assign layer3_outputs[1831] = ~((layer2_outputs[1526]) & (layer2_outputs[2512]));
    assign layer3_outputs[1832] = (layer2_outputs[511]) & ~(layer2_outputs[4099]);
    assign layer3_outputs[1833] = (layer2_outputs[4965]) & ~(layer2_outputs[3704]);
    assign layer3_outputs[1834] = layer2_outputs[877];
    assign layer3_outputs[1835] = (layer2_outputs[4039]) & ~(layer2_outputs[3380]);
    assign layer3_outputs[1836] = ~(layer2_outputs[3940]);
    assign layer3_outputs[1837] = ~(layer2_outputs[3747]);
    assign layer3_outputs[1838] = (layer2_outputs[2700]) | (layer2_outputs[886]);
    assign layer3_outputs[1839] = 1'b1;
    assign layer3_outputs[1840] = ~(layer2_outputs[3721]);
    assign layer3_outputs[1841] = layer2_outputs[4159];
    assign layer3_outputs[1842] = (layer2_outputs[4738]) ^ (layer2_outputs[5063]);
    assign layer3_outputs[1843] = ~((layer2_outputs[3444]) & (layer2_outputs[4780]));
    assign layer3_outputs[1844] = ~(layer2_outputs[610]);
    assign layer3_outputs[1845] = (layer2_outputs[2293]) | (layer2_outputs[3396]);
    assign layer3_outputs[1846] = (layer2_outputs[175]) & ~(layer2_outputs[273]);
    assign layer3_outputs[1847] = (layer2_outputs[1298]) | (layer2_outputs[1319]);
    assign layer3_outputs[1848] = ~((layer2_outputs[2309]) | (layer2_outputs[3445]));
    assign layer3_outputs[1849] = layer2_outputs[2467];
    assign layer3_outputs[1850] = ~((layer2_outputs[4796]) ^ (layer2_outputs[1325]));
    assign layer3_outputs[1851] = ~((layer2_outputs[2449]) & (layer2_outputs[67]));
    assign layer3_outputs[1852] = layer2_outputs[2901];
    assign layer3_outputs[1853] = ~(layer2_outputs[1333]) | (layer2_outputs[4160]);
    assign layer3_outputs[1854] = ~((layer2_outputs[629]) | (layer2_outputs[4811]));
    assign layer3_outputs[1855] = ~(layer2_outputs[1871]);
    assign layer3_outputs[1856] = ~(layer2_outputs[2423]);
    assign layer3_outputs[1857] = ~((layer2_outputs[3384]) | (layer2_outputs[970]));
    assign layer3_outputs[1858] = ~(layer2_outputs[4410]) | (layer2_outputs[2130]);
    assign layer3_outputs[1859] = 1'b0;
    assign layer3_outputs[1860] = ~(layer2_outputs[4637]) | (layer2_outputs[3334]);
    assign layer3_outputs[1861] = (layer2_outputs[4873]) & ~(layer2_outputs[179]);
    assign layer3_outputs[1862] = (layer2_outputs[4373]) | (layer2_outputs[1679]);
    assign layer3_outputs[1863] = (layer2_outputs[563]) ^ (layer2_outputs[3149]);
    assign layer3_outputs[1864] = ~((layer2_outputs[4418]) & (layer2_outputs[1351]));
    assign layer3_outputs[1865] = ~(layer2_outputs[713]);
    assign layer3_outputs[1866] = layer2_outputs[2524];
    assign layer3_outputs[1867] = ~(layer2_outputs[470]) | (layer2_outputs[1424]);
    assign layer3_outputs[1868] = ~((layer2_outputs[4263]) & (layer2_outputs[4753]));
    assign layer3_outputs[1869] = layer2_outputs[3426];
    assign layer3_outputs[1870] = ~((layer2_outputs[3369]) | (layer2_outputs[2359]));
    assign layer3_outputs[1871] = (layer2_outputs[1154]) & ~(layer2_outputs[975]);
    assign layer3_outputs[1872] = ~(layer2_outputs[1369]);
    assign layer3_outputs[1873] = ~(layer2_outputs[1241]);
    assign layer3_outputs[1874] = (layer2_outputs[4603]) & (layer2_outputs[3417]);
    assign layer3_outputs[1875] = 1'b0;
    assign layer3_outputs[1876] = ~(layer2_outputs[2390]) | (layer2_outputs[2465]);
    assign layer3_outputs[1877] = ~(layer2_outputs[1123]);
    assign layer3_outputs[1878] = layer2_outputs[1024];
    assign layer3_outputs[1879] = ~((layer2_outputs[1420]) | (layer2_outputs[4231]));
    assign layer3_outputs[1880] = (layer2_outputs[4104]) & (layer2_outputs[314]);
    assign layer3_outputs[1881] = layer2_outputs[2860];
    assign layer3_outputs[1882] = 1'b1;
    assign layer3_outputs[1883] = (layer2_outputs[2405]) | (layer2_outputs[1382]);
    assign layer3_outputs[1884] = ~(layer2_outputs[790]);
    assign layer3_outputs[1885] = (layer2_outputs[1401]) & ~(layer2_outputs[902]);
    assign layer3_outputs[1886] = (layer2_outputs[89]) | (layer2_outputs[930]);
    assign layer3_outputs[1887] = ~(layer2_outputs[749]);
    assign layer3_outputs[1888] = ~(layer2_outputs[3063]);
    assign layer3_outputs[1889] = 1'b0;
    assign layer3_outputs[1890] = (layer2_outputs[3716]) ^ (layer2_outputs[1247]);
    assign layer3_outputs[1891] = ~((layer2_outputs[1708]) | (layer2_outputs[1097]));
    assign layer3_outputs[1892] = ~(layer2_outputs[1971]) | (layer2_outputs[34]);
    assign layer3_outputs[1893] = (layer2_outputs[3615]) | (layer2_outputs[2515]);
    assign layer3_outputs[1894] = ~((layer2_outputs[3883]) | (layer2_outputs[2529]));
    assign layer3_outputs[1895] = ~(layer2_outputs[2408]);
    assign layer3_outputs[1896] = (layer2_outputs[1342]) & ~(layer2_outputs[2077]);
    assign layer3_outputs[1897] = layer2_outputs[3652];
    assign layer3_outputs[1898] = 1'b1;
    assign layer3_outputs[1899] = ~(layer2_outputs[547]);
    assign layer3_outputs[1900] = (layer2_outputs[3114]) & ~(layer2_outputs[2832]);
    assign layer3_outputs[1901] = ~((layer2_outputs[2765]) ^ (layer2_outputs[3]));
    assign layer3_outputs[1902] = (layer2_outputs[1046]) & ~(layer2_outputs[4597]);
    assign layer3_outputs[1903] = (layer2_outputs[2122]) & (layer2_outputs[4886]);
    assign layer3_outputs[1904] = ~(layer2_outputs[650]);
    assign layer3_outputs[1905] = (layer2_outputs[631]) & ~(layer2_outputs[4703]);
    assign layer3_outputs[1906] = layer2_outputs[326];
    assign layer3_outputs[1907] = ~(layer2_outputs[3907]) | (layer2_outputs[4653]);
    assign layer3_outputs[1908] = ~(layer2_outputs[4487]) | (layer2_outputs[1318]);
    assign layer3_outputs[1909] = ~(layer2_outputs[4412]);
    assign layer3_outputs[1910] = ~((layer2_outputs[893]) & (layer2_outputs[537]));
    assign layer3_outputs[1911] = (layer2_outputs[1293]) | (layer2_outputs[712]);
    assign layer3_outputs[1912] = ~(layer2_outputs[1608]) | (layer2_outputs[4719]);
    assign layer3_outputs[1913] = layer2_outputs[3254];
    assign layer3_outputs[1914] = (layer2_outputs[3779]) & ~(layer2_outputs[4078]);
    assign layer3_outputs[1915] = layer2_outputs[3635];
    assign layer3_outputs[1916] = ~((layer2_outputs[5031]) | (layer2_outputs[1922]));
    assign layer3_outputs[1917] = ~(layer2_outputs[2554]);
    assign layer3_outputs[1918] = ~((layer2_outputs[1264]) | (layer2_outputs[1676]));
    assign layer3_outputs[1919] = (layer2_outputs[4678]) & ~(layer2_outputs[4981]);
    assign layer3_outputs[1920] = (layer2_outputs[524]) & ~(layer2_outputs[3261]);
    assign layer3_outputs[1921] = 1'b1;
    assign layer3_outputs[1922] = ~(layer2_outputs[3760]);
    assign layer3_outputs[1923] = ~((layer2_outputs[2874]) & (layer2_outputs[3518]));
    assign layer3_outputs[1924] = ~(layer2_outputs[2573]);
    assign layer3_outputs[1925] = layer2_outputs[3845];
    assign layer3_outputs[1926] = ~((layer2_outputs[3604]) & (layer2_outputs[3824]));
    assign layer3_outputs[1927] = ~((layer2_outputs[2475]) & (layer2_outputs[1323]));
    assign layer3_outputs[1928] = ~(layer2_outputs[580]);
    assign layer3_outputs[1929] = ~(layer2_outputs[2601]) | (layer2_outputs[782]);
    assign layer3_outputs[1930] = layer2_outputs[113];
    assign layer3_outputs[1931] = 1'b1;
    assign layer3_outputs[1932] = (layer2_outputs[143]) & ~(layer2_outputs[401]);
    assign layer3_outputs[1933] = 1'b0;
    assign layer3_outputs[1934] = ~(layer2_outputs[4084]) | (layer2_outputs[916]);
    assign layer3_outputs[1935] = ~(layer2_outputs[828]) | (layer2_outputs[2165]);
    assign layer3_outputs[1936] = layer2_outputs[620];
    assign layer3_outputs[1937] = ~((layer2_outputs[4006]) & (layer2_outputs[3258]));
    assign layer3_outputs[1938] = layer2_outputs[2957];
    assign layer3_outputs[1939] = (layer2_outputs[3251]) & (layer2_outputs[1941]);
    assign layer3_outputs[1940] = (layer2_outputs[2062]) & (layer2_outputs[1958]);
    assign layer3_outputs[1941] = (layer2_outputs[1411]) ^ (layer2_outputs[3381]);
    assign layer3_outputs[1942] = ~((layer2_outputs[4577]) | (layer2_outputs[2159]));
    assign layer3_outputs[1943] = ~(layer2_outputs[2936]);
    assign layer3_outputs[1944] = 1'b1;
    assign layer3_outputs[1945] = ~((layer2_outputs[831]) | (layer2_outputs[2780]));
    assign layer3_outputs[1946] = ~(layer2_outputs[1370]);
    assign layer3_outputs[1947] = 1'b0;
    assign layer3_outputs[1948] = layer2_outputs[311];
    assign layer3_outputs[1949] = ~((layer2_outputs[1641]) ^ (layer2_outputs[1749]));
    assign layer3_outputs[1950] = ~(layer2_outputs[2215]);
    assign layer3_outputs[1951] = ~((layer2_outputs[4911]) & (layer2_outputs[1509]));
    assign layer3_outputs[1952] = (layer2_outputs[2046]) ^ (layer2_outputs[2245]);
    assign layer3_outputs[1953] = layer2_outputs[4417];
    assign layer3_outputs[1954] = (layer2_outputs[424]) & (layer2_outputs[3250]);
    assign layer3_outputs[1955] = ~((layer2_outputs[2806]) ^ (layer2_outputs[215]));
    assign layer3_outputs[1956] = ~((layer2_outputs[1916]) | (layer2_outputs[1531]));
    assign layer3_outputs[1957] = ~(layer2_outputs[4140]);
    assign layer3_outputs[1958] = ~(layer2_outputs[2031]);
    assign layer3_outputs[1959] = layer2_outputs[1947];
    assign layer3_outputs[1960] = 1'b0;
    assign layer3_outputs[1961] = 1'b1;
    assign layer3_outputs[1962] = layer2_outputs[4900];
    assign layer3_outputs[1963] = ~(layer2_outputs[3467]) | (layer2_outputs[1333]);
    assign layer3_outputs[1964] = (layer2_outputs[1873]) & (layer2_outputs[548]);
    assign layer3_outputs[1965] = layer2_outputs[844];
    assign layer3_outputs[1966] = layer2_outputs[2068];
    assign layer3_outputs[1967] = layer2_outputs[2765];
    assign layer3_outputs[1968] = ~((layer2_outputs[199]) & (layer2_outputs[2896]));
    assign layer3_outputs[1969] = 1'b1;
    assign layer3_outputs[1970] = ~((layer2_outputs[4989]) | (layer2_outputs[646]));
    assign layer3_outputs[1971] = ~(layer2_outputs[2644]) | (layer2_outputs[1249]);
    assign layer3_outputs[1972] = 1'b0;
    assign layer3_outputs[1973] = (layer2_outputs[2054]) & ~(layer2_outputs[1640]);
    assign layer3_outputs[1974] = ~(layer2_outputs[2536]) | (layer2_outputs[4504]);
    assign layer3_outputs[1975] = (layer2_outputs[2710]) & ~(layer2_outputs[880]);
    assign layer3_outputs[1976] = ~(layer2_outputs[4560]);
    assign layer3_outputs[1977] = (layer2_outputs[3153]) & ~(layer2_outputs[4552]);
    assign layer3_outputs[1978] = layer2_outputs[1901];
    assign layer3_outputs[1979] = layer2_outputs[2907];
    assign layer3_outputs[1980] = ~(layer2_outputs[39]);
    assign layer3_outputs[1981] = layer2_outputs[235];
    assign layer3_outputs[1982] = ~(layer2_outputs[4909]);
    assign layer3_outputs[1983] = layer2_outputs[732];
    assign layer3_outputs[1984] = (layer2_outputs[2978]) | (layer2_outputs[1660]);
    assign layer3_outputs[1985] = (layer2_outputs[4299]) & (layer2_outputs[4143]);
    assign layer3_outputs[1986] = (layer2_outputs[176]) | (layer2_outputs[3299]);
    assign layer3_outputs[1987] = ~(layer2_outputs[500]);
    assign layer3_outputs[1988] = ~(layer2_outputs[1549]);
    assign layer3_outputs[1989] = layer2_outputs[3634];
    assign layer3_outputs[1990] = ~(layer2_outputs[2059]);
    assign layer3_outputs[1991] = ~(layer2_outputs[3095]);
    assign layer3_outputs[1992] = ~(layer2_outputs[2446]);
    assign layer3_outputs[1993] = ~(layer2_outputs[2591]);
    assign layer3_outputs[1994] = layer2_outputs[4798];
    assign layer3_outputs[1995] = ~((layer2_outputs[1493]) | (layer2_outputs[1008]));
    assign layer3_outputs[1996] = 1'b0;
    assign layer3_outputs[1997] = ~(layer2_outputs[922]);
    assign layer3_outputs[1998] = ~((layer2_outputs[3462]) & (layer2_outputs[1892]));
    assign layer3_outputs[1999] = ~(layer2_outputs[3984]) | (layer2_outputs[4101]);
    assign layer3_outputs[2000] = ~((layer2_outputs[2962]) | (layer2_outputs[13]));
    assign layer3_outputs[2001] = ~(layer2_outputs[1158]);
    assign layer3_outputs[2002] = ~(layer2_outputs[2656]) | (layer2_outputs[748]);
    assign layer3_outputs[2003] = (layer2_outputs[4253]) & ~(layer2_outputs[1106]);
    assign layer3_outputs[2004] = (layer2_outputs[3461]) | (layer2_outputs[2826]);
    assign layer3_outputs[2005] = ~(layer2_outputs[1174]);
    assign layer3_outputs[2006] = (layer2_outputs[2980]) & (layer2_outputs[1099]);
    assign layer3_outputs[2007] = 1'b1;
    assign layer3_outputs[2008] = ~((layer2_outputs[1710]) | (layer2_outputs[3724]));
    assign layer3_outputs[2009] = 1'b0;
    assign layer3_outputs[2010] = ~(layer2_outputs[4502]) | (layer2_outputs[3740]);
    assign layer3_outputs[2011] = ~((layer2_outputs[3395]) & (layer2_outputs[2022]));
    assign layer3_outputs[2012] = 1'b0;
    assign layer3_outputs[2013] = layer2_outputs[623];
    assign layer3_outputs[2014] = ~(layer2_outputs[5014]);
    assign layer3_outputs[2015] = (layer2_outputs[4616]) & (layer2_outputs[1644]);
    assign layer3_outputs[2016] = (layer2_outputs[4641]) & ~(layer2_outputs[912]);
    assign layer3_outputs[2017] = (layer2_outputs[4158]) | (layer2_outputs[4181]);
    assign layer3_outputs[2018] = ~(layer2_outputs[4991]) | (layer2_outputs[137]);
    assign layer3_outputs[2019] = ~(layer2_outputs[1951]);
    assign layer3_outputs[2020] = (layer2_outputs[1051]) | (layer2_outputs[3852]);
    assign layer3_outputs[2021] = ~(layer2_outputs[1497]) | (layer2_outputs[1136]);
    assign layer3_outputs[2022] = ~(layer2_outputs[4658]) | (layer2_outputs[4803]);
    assign layer3_outputs[2023] = ~(layer2_outputs[3839]);
    assign layer3_outputs[2024] = ~((layer2_outputs[1322]) & (layer2_outputs[2041]));
    assign layer3_outputs[2025] = ~(layer2_outputs[286]) | (layer2_outputs[2517]);
    assign layer3_outputs[2026] = ~((layer2_outputs[2640]) | (layer2_outputs[246]));
    assign layer3_outputs[2027] = (layer2_outputs[4548]) | (layer2_outputs[3070]);
    assign layer3_outputs[2028] = (layer2_outputs[1543]) | (layer2_outputs[4784]);
    assign layer3_outputs[2029] = ~(layer2_outputs[2973]) | (layer2_outputs[2758]);
    assign layer3_outputs[2030] = ~((layer2_outputs[677]) ^ (layer2_outputs[1925]));
    assign layer3_outputs[2031] = ~(layer2_outputs[4483]) | (layer2_outputs[1276]);
    assign layer3_outputs[2032] = ~(layer2_outputs[1707]);
    assign layer3_outputs[2033] = layer2_outputs[1288];
    assign layer3_outputs[2034] = ~((layer2_outputs[2668]) ^ (layer2_outputs[3572]));
    assign layer3_outputs[2035] = 1'b1;
    assign layer3_outputs[2036] = layer2_outputs[4450];
    assign layer3_outputs[2037] = ~(layer2_outputs[1782]) | (layer2_outputs[4926]);
    assign layer3_outputs[2038] = (layer2_outputs[3381]) | (layer2_outputs[2527]);
    assign layer3_outputs[2039] = layer2_outputs[4892];
    assign layer3_outputs[2040] = ~(layer2_outputs[3194]);
    assign layer3_outputs[2041] = ~((layer2_outputs[580]) | (layer2_outputs[4586]));
    assign layer3_outputs[2042] = ~(layer2_outputs[3283]) | (layer2_outputs[4508]);
    assign layer3_outputs[2043] = layer2_outputs[3609];
    assign layer3_outputs[2044] = (layer2_outputs[2385]) & ~(layer2_outputs[4582]);
    assign layer3_outputs[2045] = ~(layer2_outputs[1488]) | (layer2_outputs[4124]);
    assign layer3_outputs[2046] = layer2_outputs[2125];
    assign layer3_outputs[2047] = (layer2_outputs[694]) & ~(layer2_outputs[4461]);
    assign layer3_outputs[2048] = 1'b1;
    assign layer3_outputs[2049] = 1'b0;
    assign layer3_outputs[2050] = ~((layer2_outputs[3992]) | (layer2_outputs[721]));
    assign layer3_outputs[2051] = (layer2_outputs[1152]) & (layer2_outputs[673]);
    assign layer3_outputs[2052] = ~(layer2_outputs[2288]);
    assign layer3_outputs[2053] = ~((layer2_outputs[2548]) | (layer2_outputs[1739]));
    assign layer3_outputs[2054] = layer2_outputs[4473];
    assign layer3_outputs[2055] = (layer2_outputs[3515]) & ~(layer2_outputs[2262]);
    assign layer3_outputs[2056] = ~((layer2_outputs[5059]) & (layer2_outputs[2004]));
    assign layer3_outputs[2057] = ~((layer2_outputs[3363]) & (layer2_outputs[4468]));
    assign layer3_outputs[2058] = ~(layer2_outputs[3830]);
    assign layer3_outputs[2059] = 1'b0;
    assign layer3_outputs[2060] = ~(layer2_outputs[1881]);
    assign layer3_outputs[2061] = ~(layer2_outputs[4331]) | (layer2_outputs[636]);
    assign layer3_outputs[2062] = ~((layer2_outputs[547]) ^ (layer2_outputs[2828]));
    assign layer3_outputs[2063] = layer2_outputs[4571];
    assign layer3_outputs[2064] = layer2_outputs[4615];
    assign layer3_outputs[2065] = 1'b0;
    assign layer3_outputs[2066] = layer2_outputs[1336];
    assign layer3_outputs[2067] = layer2_outputs[3916];
    assign layer3_outputs[2068] = (layer2_outputs[392]) & (layer2_outputs[184]);
    assign layer3_outputs[2069] = ~(layer2_outputs[4198]) | (layer2_outputs[1639]);
    assign layer3_outputs[2070] = (layer2_outputs[1626]) & (layer2_outputs[4956]);
    assign layer3_outputs[2071] = (layer2_outputs[1545]) | (layer2_outputs[3027]);
    assign layer3_outputs[2072] = ~(layer2_outputs[1165]) | (layer2_outputs[17]);
    assign layer3_outputs[2073] = layer2_outputs[1224];
    assign layer3_outputs[2074] = (layer2_outputs[1002]) & ~(layer2_outputs[875]);
    assign layer3_outputs[2075] = layer2_outputs[784];
    assign layer3_outputs[2076] = ~(layer2_outputs[839]);
    assign layer3_outputs[2077] = ~(layer2_outputs[2339]);
    assign layer3_outputs[2078] = layer2_outputs[3425];
    assign layer3_outputs[2079] = ~(layer2_outputs[542]);
    assign layer3_outputs[2080] = ~(layer2_outputs[660]) | (layer2_outputs[1766]);
    assign layer3_outputs[2081] = ~(layer2_outputs[2206]);
    assign layer3_outputs[2082] = ~(layer2_outputs[416]) | (layer2_outputs[575]);
    assign layer3_outputs[2083] = ~(layer2_outputs[2848]);
    assign layer3_outputs[2084] = ~(layer2_outputs[4751]);
    assign layer3_outputs[2085] = ~(layer2_outputs[4760]) | (layer2_outputs[2316]);
    assign layer3_outputs[2086] = ~(layer2_outputs[704]) | (layer2_outputs[4632]);
    assign layer3_outputs[2087] = (layer2_outputs[2398]) | (layer2_outputs[3991]);
    assign layer3_outputs[2088] = (layer2_outputs[1745]) ^ (layer2_outputs[73]);
    assign layer3_outputs[2089] = 1'b1;
    assign layer3_outputs[2090] = 1'b1;
    assign layer3_outputs[2091] = (layer2_outputs[456]) & ~(layer2_outputs[4883]);
    assign layer3_outputs[2092] = ~((layer2_outputs[2499]) ^ (layer2_outputs[2139]));
    assign layer3_outputs[2093] = (layer2_outputs[4287]) & ~(layer2_outputs[5001]);
    assign layer3_outputs[2094] = ~(layer2_outputs[4367]);
    assign layer3_outputs[2095] = ~((layer2_outputs[2937]) & (layer2_outputs[3030]));
    assign layer3_outputs[2096] = 1'b0;
    assign layer3_outputs[2097] = ~(layer2_outputs[3702]);
    assign layer3_outputs[2098] = (layer2_outputs[3585]) & (layer2_outputs[2949]);
    assign layer3_outputs[2099] = 1'b1;
    assign layer3_outputs[2100] = ~(layer2_outputs[3883]);
    assign layer3_outputs[2101] = 1'b1;
    assign layer3_outputs[2102] = layer2_outputs[1049];
    assign layer3_outputs[2103] = (layer2_outputs[2709]) & ~(layer2_outputs[4643]);
    assign layer3_outputs[2104] = ~(layer2_outputs[3868]) | (layer2_outputs[4019]);
    assign layer3_outputs[2105] = ~(layer2_outputs[3750]);
    assign layer3_outputs[2106] = (layer2_outputs[927]) | (layer2_outputs[4366]);
    assign layer3_outputs[2107] = (layer2_outputs[2904]) | (layer2_outputs[2253]);
    assign layer3_outputs[2108] = ~(layer2_outputs[2585]);
    assign layer3_outputs[2109] = layer2_outputs[2099];
    assign layer3_outputs[2110] = ~(layer2_outputs[4481]) | (layer2_outputs[261]);
    assign layer3_outputs[2111] = (layer2_outputs[1943]) | (layer2_outputs[788]);
    assign layer3_outputs[2112] = ~(layer2_outputs[2188]) | (layer2_outputs[1193]);
    assign layer3_outputs[2113] = (layer2_outputs[3330]) | (layer2_outputs[3466]);
    assign layer3_outputs[2114] = 1'b1;
    assign layer3_outputs[2115] = (layer2_outputs[4437]) & (layer2_outputs[225]);
    assign layer3_outputs[2116] = (layer2_outputs[4565]) | (layer2_outputs[142]);
    assign layer3_outputs[2117] = layer2_outputs[4954];
    assign layer3_outputs[2118] = ~((layer2_outputs[3150]) | (layer2_outputs[1657]));
    assign layer3_outputs[2119] = 1'b1;
    assign layer3_outputs[2120] = (layer2_outputs[3313]) & ~(layer2_outputs[3358]);
    assign layer3_outputs[2121] = (layer2_outputs[805]) | (layer2_outputs[2634]);
    assign layer3_outputs[2122] = (layer2_outputs[2403]) & ~(layer2_outputs[2925]);
    assign layer3_outputs[2123] = layer2_outputs[4789];
    assign layer3_outputs[2124] = ~(layer2_outputs[1445]) | (layer2_outputs[4909]);
    assign layer3_outputs[2125] = (layer2_outputs[1627]) ^ (layer2_outputs[4259]);
    assign layer3_outputs[2126] = ~(layer2_outputs[3837]);
    assign layer3_outputs[2127] = 1'b1;
    assign layer3_outputs[2128] = ~(layer2_outputs[4110]) | (layer2_outputs[1466]);
    assign layer3_outputs[2129] = (layer2_outputs[2117]) & ~(layer2_outputs[3252]);
    assign layer3_outputs[2130] = 1'b0;
    assign layer3_outputs[2131] = layer2_outputs[3843];
    assign layer3_outputs[2132] = ~((layer2_outputs[3258]) | (layer2_outputs[1001]));
    assign layer3_outputs[2133] = 1'b0;
    assign layer3_outputs[2134] = layer2_outputs[25];
    assign layer3_outputs[2135] = (layer2_outputs[1531]) & ~(layer2_outputs[2363]);
    assign layer3_outputs[2136] = ~(layer2_outputs[1313]);
    assign layer3_outputs[2137] = ~(layer2_outputs[3963]) | (layer2_outputs[574]);
    assign layer3_outputs[2138] = ~(layer2_outputs[1013]);
    assign layer3_outputs[2139] = ~((layer2_outputs[4943]) & (layer2_outputs[155]));
    assign layer3_outputs[2140] = 1'b1;
    assign layer3_outputs[2141] = 1'b0;
    assign layer3_outputs[2142] = layer2_outputs[536];
    assign layer3_outputs[2143] = 1'b1;
    assign layer3_outputs[2144] = ~(layer2_outputs[4642]) | (layer2_outputs[2799]);
    assign layer3_outputs[2145] = 1'b1;
    assign layer3_outputs[2146] = (layer2_outputs[1258]) & ~(layer2_outputs[1124]);
    assign layer3_outputs[2147] = 1'b1;
    assign layer3_outputs[2148] = layer2_outputs[735];
    assign layer3_outputs[2149] = ~(layer2_outputs[2424]) | (layer2_outputs[3675]);
    assign layer3_outputs[2150] = ~(layer2_outputs[1884]);
    assign layer3_outputs[2151] = ~(layer2_outputs[904]);
    assign layer3_outputs[2152] = (layer2_outputs[3742]) ^ (layer2_outputs[4850]);
    assign layer3_outputs[2153] = ~(layer2_outputs[1006]) | (layer2_outputs[4672]);
    assign layer3_outputs[2154] = (layer2_outputs[708]) & ~(layer2_outputs[4582]);
    assign layer3_outputs[2155] = 1'b1;
    assign layer3_outputs[2156] = layer2_outputs[262];
    assign layer3_outputs[2157] = ~(layer2_outputs[1918]) | (layer2_outputs[1603]);
    assign layer3_outputs[2158] = ~((layer2_outputs[1350]) & (layer2_outputs[1406]));
    assign layer3_outputs[2159] = layer2_outputs[2721];
    assign layer3_outputs[2160] = 1'b0;
    assign layer3_outputs[2161] = layer2_outputs[4635];
    assign layer3_outputs[2162] = (layer2_outputs[4045]) | (layer2_outputs[252]);
    assign layer3_outputs[2163] = (layer2_outputs[1801]) & ~(layer2_outputs[4312]);
    assign layer3_outputs[2164] = 1'b0;
    assign layer3_outputs[2165] = ~((layer2_outputs[4484]) & (layer2_outputs[4897]));
    assign layer3_outputs[2166] = layer2_outputs[4710];
    assign layer3_outputs[2167] = ~(layer2_outputs[4173]);
    assign layer3_outputs[2168] = (layer2_outputs[2491]) | (layer2_outputs[3064]);
    assign layer3_outputs[2169] = (layer2_outputs[2871]) & ~(layer2_outputs[4041]);
    assign layer3_outputs[2170] = 1'b0;
    assign layer3_outputs[2171] = (layer2_outputs[3593]) & ~(layer2_outputs[3270]);
    assign layer3_outputs[2172] = (layer2_outputs[173]) & ~(layer2_outputs[746]);
    assign layer3_outputs[2173] = ~(layer2_outputs[3361]);
    assign layer3_outputs[2174] = (layer2_outputs[279]) & ~(layer2_outputs[5023]);
    assign layer3_outputs[2175] = ~((layer2_outputs[3281]) & (layer2_outputs[691]));
    assign layer3_outputs[2176] = ~(layer2_outputs[5039]);
    assign layer3_outputs[2177] = (layer2_outputs[2055]) & ~(layer2_outputs[117]);
    assign layer3_outputs[2178] = 1'b1;
    assign layer3_outputs[2179] = ~(layer2_outputs[1200]);
    assign layer3_outputs[2180] = ~(layer2_outputs[1274]);
    assign layer3_outputs[2181] = ~(layer2_outputs[4604]);
    assign layer3_outputs[2182] = (layer2_outputs[5016]) & ~(layer2_outputs[3733]);
    assign layer3_outputs[2183] = ~(layer2_outputs[4772]);
    assign layer3_outputs[2184] = ~(layer2_outputs[3137]);
    assign layer3_outputs[2185] = (layer2_outputs[2360]) & (layer2_outputs[762]);
    assign layer3_outputs[2186] = (layer2_outputs[1477]) & (layer2_outputs[2094]);
    assign layer3_outputs[2187] = (layer2_outputs[2335]) & ~(layer2_outputs[665]);
    assign layer3_outputs[2188] = ~((layer2_outputs[1749]) | (layer2_outputs[319]));
    assign layer3_outputs[2189] = ~(layer2_outputs[4185]);
    assign layer3_outputs[2190] = (layer2_outputs[656]) | (layer2_outputs[2910]);
    assign layer3_outputs[2191] = ~(layer2_outputs[2764]);
    assign layer3_outputs[2192] = ~(layer2_outputs[2723]);
    assign layer3_outputs[2193] = layer2_outputs[151];
    assign layer3_outputs[2194] = ~((layer2_outputs[2144]) & (layer2_outputs[3911]));
    assign layer3_outputs[2195] = 1'b1;
    assign layer3_outputs[2196] = ~((layer2_outputs[1560]) & (layer2_outputs[3446]));
    assign layer3_outputs[2197] = ~(layer2_outputs[2289]) | (layer2_outputs[281]);
    assign layer3_outputs[2198] = (layer2_outputs[683]) & ~(layer2_outputs[3792]);
    assign layer3_outputs[2199] = ~(layer2_outputs[4151]);
    assign layer3_outputs[2200] = 1'b1;
    assign layer3_outputs[2201] = 1'b1;
    assign layer3_outputs[2202] = layer2_outputs[1258];
    assign layer3_outputs[2203] = ~(layer2_outputs[531]);
    assign layer3_outputs[2204] = ~(layer2_outputs[2501]);
    assign layer3_outputs[2205] = ~(layer2_outputs[4751]);
    assign layer3_outputs[2206] = ~((layer2_outputs[2888]) | (layer2_outputs[1794]));
    assign layer3_outputs[2207] = ~((layer2_outputs[1837]) ^ (layer2_outputs[3814]));
    assign layer3_outputs[2208] = (layer2_outputs[5029]) & ~(layer2_outputs[940]);
    assign layer3_outputs[2209] = ~((layer2_outputs[2858]) & (layer2_outputs[4012]));
    assign layer3_outputs[2210] = 1'b1;
    assign layer3_outputs[2211] = 1'b1;
    assign layer3_outputs[2212] = layer2_outputs[2918];
    assign layer3_outputs[2213] = (layer2_outputs[4242]) & ~(layer2_outputs[4275]);
    assign layer3_outputs[2214] = ~((layer2_outputs[4352]) ^ (layer2_outputs[2081]));
    assign layer3_outputs[2215] = (layer2_outputs[642]) | (layer2_outputs[4902]);
    assign layer3_outputs[2216] = ~(layer2_outputs[2374]) | (layer2_outputs[4400]);
    assign layer3_outputs[2217] = layer2_outputs[3282];
    assign layer3_outputs[2218] = (layer2_outputs[1677]) | (layer2_outputs[42]);
    assign layer3_outputs[2219] = ~(layer2_outputs[3783]);
    assign layer3_outputs[2220] = ~((layer2_outputs[583]) | (layer2_outputs[3185]));
    assign layer3_outputs[2221] = ~(layer2_outputs[3484]) | (layer2_outputs[4393]);
    assign layer3_outputs[2222] = (layer2_outputs[3112]) & (layer2_outputs[567]);
    assign layer3_outputs[2223] = ~(layer2_outputs[4014]);
    assign layer3_outputs[2224] = (layer2_outputs[4296]) & ~(layer2_outputs[2244]);
    assign layer3_outputs[2225] = ~(layer2_outputs[998]);
    assign layer3_outputs[2226] = (layer2_outputs[1636]) & ~(layer2_outputs[1125]);
    assign layer3_outputs[2227] = ~(layer2_outputs[1021]) | (layer2_outputs[4724]);
    assign layer3_outputs[2228] = layer2_outputs[4502];
    assign layer3_outputs[2229] = 1'b1;
    assign layer3_outputs[2230] = ~((layer2_outputs[2044]) ^ (layer2_outputs[3865]));
    assign layer3_outputs[2231] = layer2_outputs[3623];
    assign layer3_outputs[2232] = (layer2_outputs[1602]) & ~(layer2_outputs[1032]);
    assign layer3_outputs[2233] = ~((layer2_outputs[54]) & (layer2_outputs[3119]));
    assign layer3_outputs[2234] = ~(layer2_outputs[211]);
    assign layer3_outputs[2235] = ~(layer2_outputs[731]);
    assign layer3_outputs[2236] = (layer2_outputs[2246]) & ~(layer2_outputs[2943]);
    assign layer3_outputs[2237] = ~(layer2_outputs[3974]) | (layer2_outputs[4167]);
    assign layer3_outputs[2238] = (layer2_outputs[3232]) | (layer2_outputs[1096]);
    assign layer3_outputs[2239] = (layer2_outputs[368]) ^ (layer2_outputs[4520]);
    assign layer3_outputs[2240] = (layer2_outputs[4574]) & ~(layer2_outputs[923]);
    assign layer3_outputs[2241] = layer2_outputs[993];
    assign layer3_outputs[2242] = ~((layer2_outputs[2782]) | (layer2_outputs[157]));
    assign layer3_outputs[2243] = (layer2_outputs[4383]) | (layer2_outputs[4503]);
    assign layer3_outputs[2244] = ~(layer2_outputs[5110]);
    assign layer3_outputs[2245] = ~((layer2_outputs[2905]) ^ (layer2_outputs[4954]));
    assign layer3_outputs[2246] = ~(layer2_outputs[3008]);
    assign layer3_outputs[2247] = layer2_outputs[2655];
    assign layer3_outputs[2248] = ~(layer2_outputs[4617]) | (layer2_outputs[1042]);
    assign layer3_outputs[2249] = ~((layer2_outputs[652]) ^ (layer2_outputs[3981]));
    assign layer3_outputs[2250] = (layer2_outputs[56]) & ~(layer2_outputs[2003]);
    assign layer3_outputs[2251] = ~(layer2_outputs[3895]);
    assign layer3_outputs[2252] = (layer2_outputs[4741]) & (layer2_outputs[3696]);
    assign layer3_outputs[2253] = (layer2_outputs[2385]) | (layer2_outputs[4277]);
    assign layer3_outputs[2254] = (layer2_outputs[2157]) | (layer2_outputs[3162]);
    assign layer3_outputs[2255] = layer2_outputs[3604];
    assign layer3_outputs[2256] = ~(layer2_outputs[4842]) | (layer2_outputs[1755]);
    assign layer3_outputs[2257] = 1'b0;
    assign layer3_outputs[2258] = layer2_outputs[1031];
    assign layer3_outputs[2259] = layer2_outputs[1435];
    assign layer3_outputs[2260] = ~((layer2_outputs[3183]) | (layer2_outputs[2236]));
    assign layer3_outputs[2261] = ~((layer2_outputs[794]) | (layer2_outputs[2001]));
    assign layer3_outputs[2262] = 1'b1;
    assign layer3_outputs[2263] = ~((layer2_outputs[4385]) | (layer2_outputs[3891]));
    assign layer3_outputs[2264] = layer2_outputs[2329];
    assign layer3_outputs[2265] = layer2_outputs[1069];
    assign layer3_outputs[2266] = (layer2_outputs[1842]) | (layer2_outputs[4779]);
    assign layer3_outputs[2267] = layer2_outputs[3297];
    assign layer3_outputs[2268] = (layer2_outputs[105]) & ~(layer2_outputs[127]);
    assign layer3_outputs[2269] = (layer2_outputs[3373]) & ~(layer2_outputs[4016]);
    assign layer3_outputs[2270] = ~(layer2_outputs[3477]) | (layer2_outputs[3515]);
    assign layer3_outputs[2271] = ~((layer2_outputs[2844]) | (layer2_outputs[3506]));
    assign layer3_outputs[2272] = ~((layer2_outputs[560]) | (layer2_outputs[497]));
    assign layer3_outputs[2273] = ~(layer2_outputs[2533]);
    assign layer3_outputs[2274] = ~(layer2_outputs[4567]) | (layer2_outputs[3501]);
    assign layer3_outputs[2275] = (layer2_outputs[4651]) & ~(layer2_outputs[705]);
    assign layer3_outputs[2276] = ~(layer2_outputs[2228]);
    assign layer3_outputs[2277] = layer2_outputs[126];
    assign layer3_outputs[2278] = ~(layer2_outputs[878]);
    assign layer3_outputs[2279] = ~(layer2_outputs[1854]);
    assign layer3_outputs[2280] = layer2_outputs[2187];
    assign layer3_outputs[2281] = 1'b0;
    assign layer3_outputs[2282] = 1'b0;
    assign layer3_outputs[2283] = (layer2_outputs[1858]) & ~(layer2_outputs[2608]);
    assign layer3_outputs[2284] = (layer2_outputs[4739]) | (layer2_outputs[1259]);
    assign layer3_outputs[2285] = 1'b0;
    assign layer3_outputs[2286] = ~(layer2_outputs[1789]);
    assign layer3_outputs[2287] = layer2_outputs[4628];
    assign layer3_outputs[2288] = (layer2_outputs[2632]) & (layer2_outputs[2029]);
    assign layer3_outputs[2289] = ~(layer2_outputs[4572]);
    assign layer3_outputs[2290] = (layer2_outputs[2913]) & ~(layer2_outputs[925]);
    assign layer3_outputs[2291] = ~(layer2_outputs[1816]);
    assign layer3_outputs[2292] = 1'b0;
    assign layer3_outputs[2293] = (layer2_outputs[4485]) & (layer2_outputs[3806]);
    assign layer3_outputs[2294] = ~((layer2_outputs[4622]) | (layer2_outputs[4397]));
    assign layer3_outputs[2295] = (layer2_outputs[1530]) & ~(layer2_outputs[4327]);
    assign layer3_outputs[2296] = 1'b0;
    assign layer3_outputs[2297] = ~(layer2_outputs[4289]);
    assign layer3_outputs[2298] = ~((layer2_outputs[1233]) | (layer2_outputs[2464]));
    assign layer3_outputs[2299] = ~(layer2_outputs[3914]);
    assign layer3_outputs[2300] = ~((layer2_outputs[214]) | (layer2_outputs[3378]));
    assign layer3_outputs[2301] = (layer2_outputs[4662]) ^ (layer2_outputs[3107]);
    assign layer3_outputs[2302] = (layer2_outputs[1465]) & (layer2_outputs[203]);
    assign layer3_outputs[2303] = ~((layer2_outputs[2092]) ^ (layer2_outputs[2298]));
    assign layer3_outputs[2304] = ~(layer2_outputs[1334]) | (layer2_outputs[1187]);
    assign layer3_outputs[2305] = ~(layer2_outputs[1003]);
    assign layer3_outputs[2306] = ~((layer2_outputs[3671]) & (layer2_outputs[59]));
    assign layer3_outputs[2307] = layer2_outputs[2119];
    assign layer3_outputs[2308] = (layer2_outputs[803]) & ~(layer2_outputs[64]);
    assign layer3_outputs[2309] = layer2_outputs[2800];
    assign layer3_outputs[2310] = ~((layer2_outputs[368]) | (layer2_outputs[1122]));
    assign layer3_outputs[2311] = 1'b1;
    assign layer3_outputs[2312] = layer2_outputs[20];
    assign layer3_outputs[2313] = ~(layer2_outputs[1197]);
    assign layer3_outputs[2314] = ~(layer2_outputs[3374]);
    assign layer3_outputs[2315] = layer2_outputs[4131];
    assign layer3_outputs[2316] = ~(layer2_outputs[2111]);
    assign layer3_outputs[2317] = layer2_outputs[2695];
    assign layer3_outputs[2318] = ~(layer2_outputs[2386]);
    assign layer3_outputs[2319] = ~(layer2_outputs[4625]) | (layer2_outputs[1924]);
    assign layer3_outputs[2320] = ~(layer2_outputs[1127]) | (layer2_outputs[1014]);
    assign layer3_outputs[2321] = ~(layer2_outputs[4479]);
    assign layer3_outputs[2322] = (layer2_outputs[2589]) & ~(layer2_outputs[3099]);
    assign layer3_outputs[2323] = ~(layer2_outputs[4498]);
    assign layer3_outputs[2324] = ~(layer2_outputs[4030]);
    assign layer3_outputs[2325] = (layer2_outputs[1112]) ^ (layer2_outputs[1383]);
    assign layer3_outputs[2326] = (layer2_outputs[1842]) | (layer2_outputs[4091]);
    assign layer3_outputs[2327] = 1'b1;
    assign layer3_outputs[2328] = ~(layer2_outputs[4473]);
    assign layer3_outputs[2329] = layer2_outputs[2741];
    assign layer3_outputs[2330] = 1'b0;
    assign layer3_outputs[2331] = (layer2_outputs[1422]) & ~(layer2_outputs[380]);
    assign layer3_outputs[2332] = ~((layer2_outputs[1207]) & (layer2_outputs[478]));
    assign layer3_outputs[2333] = 1'b0;
    assign layer3_outputs[2334] = 1'b1;
    assign layer3_outputs[2335] = ~(layer2_outputs[907]) | (layer2_outputs[2714]);
    assign layer3_outputs[2336] = (layer2_outputs[213]) & (layer2_outputs[4465]);
    assign layer3_outputs[2337] = ~(layer2_outputs[3203]) | (layer2_outputs[90]);
    assign layer3_outputs[2338] = ~(layer2_outputs[2309]) | (layer2_outputs[2667]);
    assign layer3_outputs[2339] = (layer2_outputs[2280]) & (layer2_outputs[4650]);
    assign layer3_outputs[2340] = (layer2_outputs[469]) | (layer2_outputs[2240]);
    assign layer3_outputs[2341] = (layer2_outputs[4575]) | (layer2_outputs[4529]);
    assign layer3_outputs[2342] = (layer2_outputs[832]) | (layer2_outputs[4852]);
    assign layer3_outputs[2343] = 1'b1;
    assign layer3_outputs[2344] = (layer2_outputs[4510]) & ~(layer2_outputs[2853]);
    assign layer3_outputs[2345] = 1'b0;
    assign layer3_outputs[2346] = layer2_outputs[3748];
    assign layer3_outputs[2347] = ~(layer2_outputs[2263]);
    assign layer3_outputs[2348] = ~(layer2_outputs[2063]);
    assign layer3_outputs[2349] = ~(layer2_outputs[2666]) | (layer2_outputs[3701]);
    assign layer3_outputs[2350] = ~((layer2_outputs[1591]) | (layer2_outputs[2369]));
    assign layer3_outputs[2351] = (layer2_outputs[1499]) & ~(layer2_outputs[2884]);
    assign layer3_outputs[2352] = ~((layer2_outputs[3859]) ^ (layer2_outputs[2388]));
    assign layer3_outputs[2353] = (layer2_outputs[3436]) & (layer2_outputs[680]);
    assign layer3_outputs[2354] = ~(layer2_outputs[4713]) | (layer2_outputs[2303]);
    assign layer3_outputs[2355] = ~(layer2_outputs[5110]) | (layer2_outputs[598]);
    assign layer3_outputs[2356] = ~((layer2_outputs[1922]) | (layer2_outputs[2885]));
    assign layer3_outputs[2357] = (layer2_outputs[4438]) ^ (layer2_outputs[2267]);
    assign layer3_outputs[2358] = ~(layer2_outputs[386]);
    assign layer3_outputs[2359] = ~((layer2_outputs[610]) ^ (layer2_outputs[2489]));
    assign layer3_outputs[2360] = layer2_outputs[2549];
    assign layer3_outputs[2361] = (layer2_outputs[4003]) ^ (layer2_outputs[1421]);
    assign layer3_outputs[2362] = ~(layer2_outputs[4791]);
    assign layer3_outputs[2363] = (layer2_outputs[1466]) ^ (layer2_outputs[4462]);
    assign layer3_outputs[2364] = ~(layer2_outputs[386]);
    assign layer3_outputs[2365] = ~((layer2_outputs[1762]) | (layer2_outputs[1810]));
    assign layer3_outputs[2366] = (layer2_outputs[48]) & (layer2_outputs[3406]);
    assign layer3_outputs[2367] = ~(layer2_outputs[1832]);
    assign layer3_outputs[2368] = ~((layer2_outputs[5051]) ^ (layer2_outputs[2073]));
    assign layer3_outputs[2369] = layer2_outputs[679];
    assign layer3_outputs[2370] = ~(layer2_outputs[16]);
    assign layer3_outputs[2371] = (layer2_outputs[4053]) ^ (layer2_outputs[1857]);
    assign layer3_outputs[2372] = 1'b1;
    assign layer3_outputs[2373] = (layer2_outputs[2944]) ^ (layer2_outputs[1952]);
    assign layer3_outputs[2374] = ~((layer2_outputs[4608]) & (layer2_outputs[5018]));
    assign layer3_outputs[2375] = layer2_outputs[3369];
    assign layer3_outputs[2376] = layer2_outputs[4758];
    assign layer3_outputs[2377] = layer2_outputs[1548];
    assign layer3_outputs[2378] = ~((layer2_outputs[4431]) | (layer2_outputs[3389]));
    assign layer3_outputs[2379] = (layer2_outputs[2470]) & (layer2_outputs[3567]);
    assign layer3_outputs[2380] = (layer2_outputs[4937]) & (layer2_outputs[3217]);
    assign layer3_outputs[2381] = 1'b0;
    assign layer3_outputs[2382] = 1'b0;
    assign layer3_outputs[2383] = 1'b0;
    assign layer3_outputs[2384] = ~(layer2_outputs[1733]) | (layer2_outputs[2033]);
    assign layer3_outputs[2385] = ~(layer2_outputs[4944]);
    assign layer3_outputs[2386] = layer2_outputs[2372];
    assign layer3_outputs[2387] = layer2_outputs[2706];
    assign layer3_outputs[2388] = layer2_outputs[126];
    assign layer3_outputs[2389] = (layer2_outputs[2032]) ^ (layer2_outputs[464]);
    assign layer3_outputs[2390] = ~((layer2_outputs[2216]) & (layer2_outputs[3584]));
    assign layer3_outputs[2391] = layer2_outputs[3538];
    assign layer3_outputs[2392] = ~(layer2_outputs[1115]) | (layer2_outputs[3435]);
    assign layer3_outputs[2393] = layer2_outputs[1800];
    assign layer3_outputs[2394] = ~(layer2_outputs[4945]);
    assign layer3_outputs[2395] = (layer2_outputs[137]) | (layer2_outputs[3399]);
    assign layer3_outputs[2396] = ~(layer2_outputs[372]) | (layer2_outputs[4640]);
    assign layer3_outputs[2397] = (layer2_outputs[1816]) | (layer2_outputs[222]);
    assign layer3_outputs[2398] = ~(layer2_outputs[2511]);
    assign layer3_outputs[2399] = layer2_outputs[3892];
    assign layer3_outputs[2400] = 1'b0;
    assign layer3_outputs[2401] = (layer2_outputs[1139]) & ~(layer2_outputs[3430]);
    assign layer3_outputs[2402] = ~((layer2_outputs[540]) | (layer2_outputs[2185]));
    assign layer3_outputs[2403] = (layer2_outputs[470]) & (layer2_outputs[82]);
    assign layer3_outputs[2404] = (layer2_outputs[2539]) & ~(layer2_outputs[298]);
    assign layer3_outputs[2405] = layer2_outputs[1699];
    assign layer3_outputs[2406] = (layer2_outputs[1836]) & ~(layer2_outputs[4234]);
    assign layer3_outputs[2407] = ~(layer2_outputs[4108]);
    assign layer3_outputs[2408] = layer2_outputs[5079];
    assign layer3_outputs[2409] = ~(layer2_outputs[3044]);
    assign layer3_outputs[2410] = (layer2_outputs[1249]) & (layer2_outputs[3301]);
    assign layer3_outputs[2411] = ~((layer2_outputs[1403]) ^ (layer2_outputs[3807]));
    assign layer3_outputs[2412] = ~(layer2_outputs[2913]);
    assign layer3_outputs[2413] = (layer2_outputs[4196]) | (layer2_outputs[4331]);
    assign layer3_outputs[2414] = layer2_outputs[777];
    assign layer3_outputs[2415] = layer2_outputs[2992];
    assign layer3_outputs[2416] = (layer2_outputs[5062]) | (layer2_outputs[2464]);
    assign layer3_outputs[2417] = 1'b1;
    assign layer3_outputs[2418] = ~(layer2_outputs[3726]);
    assign layer3_outputs[2419] = (layer2_outputs[1078]) | (layer2_outputs[519]);
    assign layer3_outputs[2420] = (layer2_outputs[1791]) | (layer2_outputs[4]);
    assign layer3_outputs[2421] = ~((layer2_outputs[2438]) | (layer2_outputs[3536]));
    assign layer3_outputs[2422] = layer2_outputs[4786];
    assign layer3_outputs[2423] = 1'b0;
    assign layer3_outputs[2424] = layer2_outputs[1164];
    assign layer3_outputs[2425] = ~(layer2_outputs[4784]) | (layer2_outputs[2826]);
    assign layer3_outputs[2426] = ~((layer2_outputs[4055]) | (layer2_outputs[2564]));
    assign layer3_outputs[2427] = 1'b1;
    assign layer3_outputs[2428] = layer2_outputs[4334];
    assign layer3_outputs[2429] = (layer2_outputs[4812]) & ~(layer2_outputs[1524]);
    assign layer3_outputs[2430] = ~(layer2_outputs[1412]);
    assign layer3_outputs[2431] = (layer2_outputs[4774]) & (layer2_outputs[1908]);
    assign layer3_outputs[2432] = (layer2_outputs[3422]) & (layer2_outputs[1752]);
    assign layer3_outputs[2433] = ~((layer2_outputs[4829]) & (layer2_outputs[1294]));
    assign layer3_outputs[2434] = (layer2_outputs[2174]) & ~(layer2_outputs[2030]);
    assign layer3_outputs[2435] = 1'b0;
    assign layer3_outputs[2436] = layer2_outputs[4702];
    assign layer3_outputs[2437] = layer2_outputs[79];
    assign layer3_outputs[2438] = ~(layer2_outputs[1426]);
    assign layer3_outputs[2439] = ~(layer2_outputs[3965]) | (layer2_outputs[681]);
    assign layer3_outputs[2440] = (layer2_outputs[3803]) & ~(layer2_outputs[4968]);
    assign layer3_outputs[2441] = (layer2_outputs[2699]) & ~(layer2_outputs[3447]);
    assign layer3_outputs[2442] = (layer2_outputs[1905]) & (layer2_outputs[63]);
    assign layer3_outputs[2443] = layer2_outputs[3712];
    assign layer3_outputs[2444] = layer2_outputs[613];
    assign layer3_outputs[2445] = layer2_outputs[3261];
    assign layer3_outputs[2446] = ~(layer2_outputs[3175]);
    assign layer3_outputs[2447] = (layer2_outputs[309]) & ~(layer2_outputs[1386]);
    assign layer3_outputs[2448] = (layer2_outputs[2070]) & ~(layer2_outputs[3334]);
    assign layer3_outputs[2449] = ~((layer2_outputs[3495]) & (layer2_outputs[1478]));
    assign layer3_outputs[2450] = (layer2_outputs[1905]) & (layer2_outputs[110]);
    assign layer3_outputs[2451] = 1'b0;
    assign layer3_outputs[2452] = layer2_outputs[2751];
    assign layer3_outputs[2453] = ~(layer2_outputs[4975]) | (layer2_outputs[90]);
    assign layer3_outputs[2454] = ~(layer2_outputs[969]);
    assign layer3_outputs[2455] = ~((layer2_outputs[1754]) & (layer2_outputs[3877]));
    assign layer3_outputs[2456] = ~(layer2_outputs[3994]);
    assign layer3_outputs[2457] = ~(layer2_outputs[4433]) | (layer2_outputs[41]);
    assign layer3_outputs[2458] = ~((layer2_outputs[1551]) ^ (layer2_outputs[1232]));
    assign layer3_outputs[2459] = layer2_outputs[4017];
    assign layer3_outputs[2460] = (layer2_outputs[1808]) ^ (layer2_outputs[2400]);
    assign layer3_outputs[2461] = layer2_outputs[1590];
    assign layer3_outputs[2462] = ~((layer2_outputs[599]) | (layer2_outputs[1199]));
    assign layer3_outputs[2463] = layer2_outputs[2764];
    assign layer3_outputs[2464] = ~(layer2_outputs[4081]);
    assign layer3_outputs[2465] = ~(layer2_outputs[359]);
    assign layer3_outputs[2466] = ~((layer2_outputs[1467]) & (layer2_outputs[1381]));
    assign layer3_outputs[2467] = ~((layer2_outputs[660]) | (layer2_outputs[2487]));
    assign layer3_outputs[2468] = layer2_outputs[2373];
    assign layer3_outputs[2469] = ~((layer2_outputs[640]) ^ (layer2_outputs[239]));
    assign layer3_outputs[2470] = ~(layer2_outputs[3846]);
    assign layer3_outputs[2471] = (layer2_outputs[3148]) & ~(layer2_outputs[1968]);
    assign layer3_outputs[2472] = layer2_outputs[570];
    assign layer3_outputs[2473] = layer2_outputs[2027];
    assign layer3_outputs[2474] = ~(layer2_outputs[2691]);
    assign layer3_outputs[2475] = (layer2_outputs[2550]) & (layer2_outputs[2061]);
    assign layer3_outputs[2476] = ~((layer2_outputs[1945]) & (layer2_outputs[2760]));
    assign layer3_outputs[2477] = ~((layer2_outputs[1463]) | (layer2_outputs[3512]));
    assign layer3_outputs[2478] = (layer2_outputs[1183]) | (layer2_outputs[3809]);
    assign layer3_outputs[2479] = ~(layer2_outputs[1741]) | (layer2_outputs[2746]);
    assign layer3_outputs[2480] = ~(layer2_outputs[4668]);
    assign layer3_outputs[2481] = (layer2_outputs[1667]) | (layer2_outputs[2650]);
    assign layer3_outputs[2482] = ~(layer2_outputs[2884]);
    assign layer3_outputs[2483] = ~(layer2_outputs[3411]);
    assign layer3_outputs[2484] = layer2_outputs[4788];
    assign layer3_outputs[2485] = ~(layer2_outputs[3051]);
    assign layer3_outputs[2486] = layer2_outputs[3874];
    assign layer3_outputs[2487] = layer2_outputs[1939];
    assign layer3_outputs[2488] = ~(layer2_outputs[293]);
    assign layer3_outputs[2489] = (layer2_outputs[2052]) | (layer2_outputs[3447]);
    assign layer3_outputs[2490] = ~((layer2_outputs[2260]) ^ (layer2_outputs[3570]));
    assign layer3_outputs[2491] = 1'b0;
    assign layer3_outputs[2492] = ~(layer2_outputs[374]);
    assign layer3_outputs[2493] = (layer2_outputs[3672]) | (layer2_outputs[1935]);
    assign layer3_outputs[2494] = ~((layer2_outputs[2098]) | (layer2_outputs[3561]));
    assign layer3_outputs[2495] = (layer2_outputs[2854]) & ~(layer2_outputs[4769]);
    assign layer3_outputs[2496] = layer2_outputs[4946];
    assign layer3_outputs[2497] = ~((layer2_outputs[3486]) | (layer2_outputs[3111]));
    assign layer3_outputs[2498] = ~((layer2_outputs[5061]) & (layer2_outputs[847]));
    assign layer3_outputs[2499] = ~(layer2_outputs[2689]) | (layer2_outputs[806]);
    assign layer3_outputs[2500] = layer2_outputs[3976];
    assign layer3_outputs[2501] = layer2_outputs[4140];
    assign layer3_outputs[2502] = (layer2_outputs[1510]) & ~(layer2_outputs[3260]);
    assign layer3_outputs[2503] = (layer2_outputs[4414]) & ~(layer2_outputs[945]);
    assign layer3_outputs[2504] = ~(layer2_outputs[1886]);
    assign layer3_outputs[2505] = (layer2_outputs[274]) | (layer2_outputs[4601]);
    assign layer3_outputs[2506] = ~(layer2_outputs[4842]);
    assign layer3_outputs[2507] = ~(layer2_outputs[2320]) | (layer2_outputs[4754]);
    assign layer3_outputs[2508] = 1'b1;
    assign layer3_outputs[2509] = ~(layer2_outputs[4265]);
    assign layer3_outputs[2510] = layer2_outputs[929];
    assign layer3_outputs[2511] = (layer2_outputs[1376]) & (layer2_outputs[600]);
    assign layer3_outputs[2512] = ~(layer2_outputs[2478]) | (layer2_outputs[4475]);
    assign layer3_outputs[2513] = (layer2_outputs[2501]) | (layer2_outputs[3198]);
    assign layer3_outputs[2514] = layer2_outputs[925];
    assign layer3_outputs[2515] = ~(layer2_outputs[1347]);
    assign layer3_outputs[2516] = ~(layer2_outputs[240]);
    assign layer3_outputs[2517] = ~((layer2_outputs[1681]) | (layer2_outputs[4818]));
    assign layer3_outputs[2518] = ~(layer2_outputs[695]) | (layer2_outputs[1726]);
    assign layer3_outputs[2519] = 1'b1;
    assign layer3_outputs[2520] = ~((layer2_outputs[5115]) | (layer2_outputs[2104]));
    assign layer3_outputs[2521] = ~(layer2_outputs[1372]);
    assign layer3_outputs[2522] = (layer2_outputs[3096]) | (layer2_outputs[5004]);
    assign layer3_outputs[2523] = ~(layer2_outputs[599]) | (layer2_outputs[501]);
    assign layer3_outputs[2524] = 1'b1;
    assign layer3_outputs[2525] = layer2_outputs[958];
    assign layer3_outputs[2526] = ~(layer2_outputs[4555]);
    assign layer3_outputs[2527] = (layer2_outputs[3895]) & ~(layer2_outputs[3530]);
    assign layer3_outputs[2528] = ~((layer2_outputs[3337]) & (layer2_outputs[3980]));
    assign layer3_outputs[2529] = layer2_outputs[828];
    assign layer3_outputs[2530] = (layer2_outputs[3745]) & ~(layer2_outputs[4192]);
    assign layer3_outputs[2531] = layer2_outputs[2738];
    assign layer3_outputs[2532] = ~(layer2_outputs[564]);
    assign layer3_outputs[2533] = layer2_outputs[2369];
    assign layer3_outputs[2534] = 1'b1;
    assign layer3_outputs[2535] = ~((layer2_outputs[267]) | (layer2_outputs[4943]));
    assign layer3_outputs[2536] = layer2_outputs[1632];
    assign layer3_outputs[2537] = (layer2_outputs[845]) ^ (layer2_outputs[1301]);
    assign layer3_outputs[2538] = ~(layer2_outputs[1736]);
    assign layer3_outputs[2539] = (layer2_outputs[257]) & ~(layer2_outputs[1519]);
    assign layer3_outputs[2540] = layer2_outputs[3439];
    assign layer3_outputs[2541] = ~(layer2_outputs[2421]) | (layer2_outputs[2734]);
    assign layer3_outputs[2542] = layer2_outputs[4092];
    assign layer3_outputs[2543] = 1'b0;
    assign layer3_outputs[2544] = 1'b1;
    assign layer3_outputs[2545] = (layer2_outputs[4406]) & ~(layer2_outputs[3129]);
    assign layer3_outputs[2546] = ~(layer2_outputs[4567]) | (layer2_outputs[3209]);
    assign layer3_outputs[2547] = (layer2_outputs[2699]) ^ (layer2_outputs[49]);
    assign layer3_outputs[2548] = ~((layer2_outputs[4303]) & (layer2_outputs[4737]));
    assign layer3_outputs[2549] = ~(layer2_outputs[2461]);
    assign layer3_outputs[2550] = (layer2_outputs[3955]) & (layer2_outputs[2634]);
    assign layer3_outputs[2551] = ~(layer2_outputs[2054]) | (layer2_outputs[2646]);
    assign layer3_outputs[2552] = ~(layer2_outputs[390]);
    assign layer3_outputs[2553] = layer2_outputs[1683];
    assign layer3_outputs[2554] = 1'b1;
    assign layer3_outputs[2555] = ~(layer2_outputs[4024]);
    assign layer3_outputs[2556] = (layer2_outputs[1770]) | (layer2_outputs[1528]);
    assign layer3_outputs[2557] = ~(layer2_outputs[4333]) | (layer2_outputs[2030]);
    assign layer3_outputs[2558] = (layer2_outputs[2630]) & (layer2_outputs[2100]);
    assign layer3_outputs[2559] = layer2_outputs[865];
    assign layer3_outputs[2560] = ~(layer2_outputs[2965]) | (layer2_outputs[1992]);
    assign layer3_outputs[2561] = ~(layer2_outputs[4755]);
    assign layer3_outputs[2562] = 1'b0;
    assign layer3_outputs[2563] = 1'b1;
    assign layer3_outputs[2564] = layer2_outputs[3569];
    assign layer3_outputs[2565] = (layer2_outputs[4918]) ^ (layer2_outputs[5013]);
    assign layer3_outputs[2566] = 1'b1;
    assign layer3_outputs[2567] = layer2_outputs[3076];
    assign layer3_outputs[2568] = (layer2_outputs[2508]) | (layer2_outputs[2609]);
    assign layer3_outputs[2569] = (layer2_outputs[3226]) ^ (layer2_outputs[1063]);
    assign layer3_outputs[2570] = ~(layer2_outputs[1817]) | (layer2_outputs[4715]);
    assign layer3_outputs[2571] = layer2_outputs[4930];
    assign layer3_outputs[2572] = 1'b0;
    assign layer3_outputs[2573] = ~(layer2_outputs[1554]) | (layer2_outputs[1663]);
    assign layer3_outputs[2574] = layer2_outputs[974];
    assign layer3_outputs[2575] = 1'b0;
    assign layer3_outputs[2576] = 1'b1;
    assign layer3_outputs[2577] = layer2_outputs[4008];
    assign layer3_outputs[2578] = ~((layer2_outputs[1638]) & (layer2_outputs[1617]));
    assign layer3_outputs[2579] = layer2_outputs[2518];
    assign layer3_outputs[2580] = ~(layer2_outputs[3152]);
    assign layer3_outputs[2581] = layer2_outputs[185];
    assign layer3_outputs[2582] = (layer2_outputs[3815]) | (layer2_outputs[4853]);
    assign layer3_outputs[2583] = (layer2_outputs[4652]) & ~(layer2_outputs[675]);
    assign layer3_outputs[2584] = 1'b0;
    assign layer3_outputs[2585] = ~(layer2_outputs[4479]);
    assign layer3_outputs[2586] = layer2_outputs[1208];
    assign layer3_outputs[2587] = (layer2_outputs[478]) & ~(layer2_outputs[876]);
    assign layer3_outputs[2588] = 1'b0;
    assign layer3_outputs[2589] = ~(layer2_outputs[2131]) | (layer2_outputs[1885]);
    assign layer3_outputs[2590] = ~((layer2_outputs[4137]) & (layer2_outputs[4496]));
    assign layer3_outputs[2591] = ~(layer2_outputs[3423]);
    assign layer3_outputs[2592] = (layer2_outputs[4403]) & ~(layer2_outputs[4434]);
    assign layer3_outputs[2593] = 1'b0;
    assign layer3_outputs[2594] = layer2_outputs[1714];
    assign layer3_outputs[2595] = 1'b0;
    assign layer3_outputs[2596] = ~((layer2_outputs[2784]) ^ (layer2_outputs[3170]));
    assign layer3_outputs[2597] = (layer2_outputs[1740]) | (layer2_outputs[4407]);
    assign layer3_outputs[2598] = ~((layer2_outputs[1718]) | (layer2_outputs[1645]));
    assign layer3_outputs[2599] = ~(layer2_outputs[2683]) | (layer2_outputs[1261]);
    assign layer3_outputs[2600] = layer2_outputs[1012];
    assign layer3_outputs[2601] = 1'b1;
    assign layer3_outputs[2602] = (layer2_outputs[515]) & ~(layer2_outputs[1255]);
    assign layer3_outputs[2603] = ~(layer2_outputs[4171]);
    assign layer3_outputs[2604] = 1'b1;
    assign layer3_outputs[2605] = ~((layer2_outputs[4378]) ^ (layer2_outputs[3459]));
    assign layer3_outputs[2606] = layer2_outputs[2546];
    assign layer3_outputs[2607] = (layer2_outputs[4394]) & (layer2_outputs[3562]);
    assign layer3_outputs[2608] = layer2_outputs[2614];
    assign layer3_outputs[2609] = ~(layer2_outputs[3098]);
    assign layer3_outputs[2610] = ~(layer2_outputs[108]);
    assign layer3_outputs[2611] = ~((layer2_outputs[3023]) | (layer2_outputs[507]));
    assign layer3_outputs[2612] = ~(layer2_outputs[3326]);
    assign layer3_outputs[2613] = (layer2_outputs[265]) & ~(layer2_outputs[3113]);
    assign layer3_outputs[2614] = ~((layer2_outputs[4319]) | (layer2_outputs[1984]));
    assign layer3_outputs[2615] = layer2_outputs[338];
    assign layer3_outputs[2616] = layer2_outputs[627];
    assign layer3_outputs[2617] = ~(layer2_outputs[2207]) | (layer2_outputs[4084]);
    assign layer3_outputs[2618] = ~(layer2_outputs[3050]);
    assign layer3_outputs[2619] = (layer2_outputs[5024]) | (layer2_outputs[1181]);
    assign layer3_outputs[2620] = layer2_outputs[2295];
    assign layer3_outputs[2621] = ~((layer2_outputs[4204]) | (layer2_outputs[965]));
    assign layer3_outputs[2622] = ~(layer2_outputs[3907]) | (layer2_outputs[2955]);
    assign layer3_outputs[2623] = (layer2_outputs[3164]) & ~(layer2_outputs[1220]);
    assign layer3_outputs[2624] = (layer2_outputs[3049]) ^ (layer2_outputs[1123]);
    assign layer3_outputs[2625] = 1'b1;
    assign layer3_outputs[2626] = (layer2_outputs[208]) & ~(layer2_outputs[236]);
    assign layer3_outputs[2627] = 1'b1;
    assign layer3_outputs[2628] = (layer2_outputs[1394]) & (layer2_outputs[3783]);
    assign layer3_outputs[2629] = ~(layer2_outputs[4515]) | (layer2_outputs[1821]);
    assign layer3_outputs[2630] = 1'b0;
    assign layer3_outputs[2631] = ~((layer2_outputs[1742]) | (layer2_outputs[4876]));
    assign layer3_outputs[2632] = layer2_outputs[299];
    assign layer3_outputs[2633] = ~(layer2_outputs[4611]);
    assign layer3_outputs[2634] = 1'b0;
    assign layer3_outputs[2635] = ~((layer2_outputs[545]) | (layer2_outputs[1598]));
    assign layer3_outputs[2636] = ~(layer2_outputs[4703]);
    assign layer3_outputs[2637] = ~((layer2_outputs[566]) & (layer2_outputs[3797]));
    assign layer3_outputs[2638] = 1'b1;
    assign layer3_outputs[2639] = (layer2_outputs[781]) & (layer2_outputs[2043]);
    assign layer3_outputs[2640] = (layer2_outputs[747]) | (layer2_outputs[1765]);
    assign layer3_outputs[2641] = ~((layer2_outputs[980]) | (layer2_outputs[3893]));
    assign layer3_outputs[2642] = layer2_outputs[840];
    assign layer3_outputs[2643] = layer2_outputs[1854];
    assign layer3_outputs[2644] = ~(layer2_outputs[5067]) | (layer2_outputs[2822]);
    assign layer3_outputs[2645] = (layer2_outputs[1664]) & ~(layer2_outputs[1811]);
    assign layer3_outputs[2646] = ~(layer2_outputs[643]);
    assign layer3_outputs[2647] = (layer2_outputs[5109]) & ~(layer2_outputs[1287]);
    assign layer3_outputs[2648] = layer2_outputs[2017];
    assign layer3_outputs[2649] = ~(layer2_outputs[2301]);
    assign layer3_outputs[2650] = ~(layer2_outputs[2576]);
    assign layer3_outputs[2651] = layer2_outputs[3202];
    assign layer3_outputs[2652] = layer2_outputs[287];
    assign layer3_outputs[2653] = layer2_outputs[3673];
    assign layer3_outputs[2654] = ~(layer2_outputs[4218]) | (layer2_outputs[1614]);
    assign layer3_outputs[2655] = (layer2_outputs[269]) & ~(layer2_outputs[1756]);
    assign layer3_outputs[2656] = 1'b1;
    assign layer3_outputs[2657] = 1'b0;
    assign layer3_outputs[2658] = (layer2_outputs[480]) & ~(layer2_outputs[3591]);
    assign layer3_outputs[2659] = ~((layer2_outputs[3015]) | (layer2_outputs[4050]));
    assign layer3_outputs[2660] = layer2_outputs[559];
    assign layer3_outputs[2661] = layer2_outputs[4457];
    assign layer3_outputs[2662] = 1'b0;
    assign layer3_outputs[2663] = (layer2_outputs[2986]) & (layer2_outputs[4906]);
    assign layer3_outputs[2664] = (layer2_outputs[2531]) ^ (layer2_outputs[582]);
    assign layer3_outputs[2665] = (layer2_outputs[1364]) & (layer2_outputs[2428]);
    assign layer3_outputs[2666] = ~(layer2_outputs[4120]);
    assign layer3_outputs[2667] = (layer2_outputs[569]) & ~(layer2_outputs[2149]);
    assign layer3_outputs[2668] = ~(layer2_outputs[4896]);
    assign layer3_outputs[2669] = ~(layer2_outputs[350]) | (layer2_outputs[2727]);
    assign layer3_outputs[2670] = ~((layer2_outputs[2164]) & (layer2_outputs[4375]));
    assign layer3_outputs[2671] = ~(layer2_outputs[835]) | (layer2_outputs[4146]);
    assign layer3_outputs[2672] = layer2_outputs[2462];
    assign layer3_outputs[2673] = (layer2_outputs[339]) & (layer2_outputs[834]);
    assign layer3_outputs[2674] = 1'b0;
    assign layer3_outputs[2675] = ~((layer2_outputs[3056]) & (layer2_outputs[4928]));
    assign layer3_outputs[2676] = ~(layer2_outputs[5112]) | (layer2_outputs[2399]);
    assign layer3_outputs[2677] = (layer2_outputs[3455]) & ~(layer2_outputs[3430]);
    assign layer3_outputs[2678] = 1'b0;
    assign layer3_outputs[2679] = layer2_outputs[1059];
    assign layer3_outputs[2680] = ~((layer2_outputs[23]) ^ (layer2_outputs[4568]));
    assign layer3_outputs[2681] = ~((layer2_outputs[2195]) | (layer2_outputs[77]));
    assign layer3_outputs[2682] = layer2_outputs[2274];
    assign layer3_outputs[2683] = ~(layer2_outputs[2846]);
    assign layer3_outputs[2684] = layer2_outputs[770];
    assign layer3_outputs[2685] = ~((layer2_outputs[2179]) ^ (layer2_outputs[3130]));
    assign layer3_outputs[2686] = 1'b1;
    assign layer3_outputs[2687] = 1'b1;
    assign layer3_outputs[2688] = layer2_outputs[123];
    assign layer3_outputs[2689] = ~(layer2_outputs[174]);
    assign layer3_outputs[2690] = (layer2_outputs[2186]) & (layer2_outputs[504]);
    assign layer3_outputs[2691] = (layer2_outputs[4754]) & ~(layer2_outputs[282]);
    assign layer3_outputs[2692] = ~(layer2_outputs[2171]);
    assign layer3_outputs[2693] = ~(layer2_outputs[4245]) | (layer2_outputs[2416]);
    assign layer3_outputs[2694] = ~(layer2_outputs[831]) | (layer2_outputs[2833]);
    assign layer3_outputs[2695] = ~(layer2_outputs[1390]);
    assign layer3_outputs[2696] = ~(layer2_outputs[243]) | (layer2_outputs[1506]);
    assign layer3_outputs[2697] = ~((layer2_outputs[4212]) | (layer2_outputs[287]));
    assign layer3_outputs[2698] = (layer2_outputs[2675]) & ~(layer2_outputs[2986]);
    assign layer3_outputs[2699] = ~(layer2_outputs[509]) | (layer2_outputs[3838]);
    assign layer3_outputs[2700] = ~(layer2_outputs[2999]);
    assign layer3_outputs[2701] = (layer2_outputs[61]) ^ (layer2_outputs[2555]);
    assign layer3_outputs[2702] = ~((layer2_outputs[4198]) & (layer2_outputs[374]));
    assign layer3_outputs[2703] = ~((layer2_outputs[160]) & (layer2_outputs[2007]));
    assign layer3_outputs[2704] = ~(layer2_outputs[2577]);
    assign layer3_outputs[2705] = layer2_outputs[3009];
    assign layer3_outputs[2706] = ~((layer2_outputs[4459]) & (layer2_outputs[860]));
    assign layer3_outputs[2707] = (layer2_outputs[1797]) & ~(layer2_outputs[4460]);
    assign layer3_outputs[2708] = ~(layer2_outputs[1863]);
    assign layer3_outputs[2709] = ~(layer2_outputs[4057]) | (layer2_outputs[2294]);
    assign layer3_outputs[2710] = ~(layer2_outputs[2050]) | (layer2_outputs[4959]);
    assign layer3_outputs[2711] = (layer2_outputs[3204]) & ~(layer2_outputs[2920]);
    assign layer3_outputs[2712] = (layer2_outputs[3917]) & ~(layer2_outputs[108]);
    assign layer3_outputs[2713] = (layer2_outputs[532]) | (layer2_outputs[4990]);
    assign layer3_outputs[2714] = (layer2_outputs[4056]) & ~(layer2_outputs[3311]);
    assign layer3_outputs[2715] = 1'b1;
    assign layer3_outputs[2716] = (layer2_outputs[93]) | (layer2_outputs[3482]);
    assign layer3_outputs[2717] = ~((layer2_outputs[2299]) | (layer2_outputs[1126]));
    assign layer3_outputs[2718] = layer2_outputs[293];
    assign layer3_outputs[2719] = layer2_outputs[746];
    assign layer3_outputs[2720] = layer2_outputs[3958];
    assign layer3_outputs[2721] = ~(layer2_outputs[1025]);
    assign layer3_outputs[2722] = (layer2_outputs[4160]) & (layer2_outputs[624]);
    assign layer3_outputs[2723] = layer2_outputs[2235];
    assign layer3_outputs[2724] = 1'b1;
    assign layer3_outputs[2725] = ~(layer2_outputs[4789]);
    assign layer3_outputs[2726] = (layer2_outputs[3072]) | (layer2_outputs[2479]);
    assign layer3_outputs[2727] = layer2_outputs[1868];
    assign layer3_outputs[2728] = ~(layer2_outputs[4247]);
    assign layer3_outputs[2729] = ~(layer2_outputs[2919]) | (layer2_outputs[707]);
    assign layer3_outputs[2730] = ~(layer2_outputs[1061]);
    assign layer3_outputs[2731] = ~((layer2_outputs[381]) & (layer2_outputs[1373]));
    assign layer3_outputs[2732] = (layer2_outputs[1214]) & ~(layer2_outputs[4584]);
    assign layer3_outputs[2733] = ~(layer2_outputs[2010]) | (layer2_outputs[2578]);
    assign layer3_outputs[2734] = ~(layer2_outputs[2994]);
    assign layer3_outputs[2735] = layer2_outputs[4377];
    assign layer3_outputs[2736] = ~(layer2_outputs[4391]) | (layer2_outputs[2477]);
    assign layer3_outputs[2737] = 1'b1;
    assign layer3_outputs[2738] = ~(layer2_outputs[3032]) | (layer2_outputs[3104]);
    assign layer3_outputs[2739] = ~(layer2_outputs[720]) | (layer2_outputs[3800]);
    assign layer3_outputs[2740] = ~(layer2_outputs[2893]) | (layer2_outputs[1280]);
    assign layer3_outputs[2741] = 1'b1;
    assign layer3_outputs[2742] = (layer2_outputs[1744]) | (layer2_outputs[4419]);
    assign layer3_outputs[2743] = ~(layer2_outputs[1988]);
    assign layer3_outputs[2744] = ~(layer2_outputs[2272]) | (layer2_outputs[1372]);
    assign layer3_outputs[2745] = ~((layer2_outputs[3542]) ^ (layer2_outputs[4207]));
    assign layer3_outputs[2746] = 1'b1;
    assign layer3_outputs[2747] = ~(layer2_outputs[1962]);
    assign layer3_outputs[2748] = ~(layer2_outputs[1064]);
    assign layer3_outputs[2749] = ~(layer2_outputs[4556]) | (layer2_outputs[980]);
    assign layer3_outputs[2750] = (layer2_outputs[4563]) & ~(layer2_outputs[3291]);
    assign layer3_outputs[2751] = layer2_outputs[3223];
    assign layer3_outputs[2752] = ~(layer2_outputs[1955]);
    assign layer3_outputs[2753] = ~(layer2_outputs[2459]) | (layer2_outputs[2977]);
    assign layer3_outputs[2754] = (layer2_outputs[4442]) & ~(layer2_outputs[2848]);
    assign layer3_outputs[2755] = ~(layer2_outputs[5021]);
    assign layer3_outputs[2756] = ~((layer2_outputs[3608]) ^ (layer2_outputs[4201]));
    assign layer3_outputs[2757] = ~(layer2_outputs[3420]);
    assign layer3_outputs[2758] = (layer2_outputs[3401]) & ~(layer2_outputs[465]);
    assign layer3_outputs[2759] = 1'b1;
    assign layer3_outputs[2760] = (layer2_outputs[4203]) | (layer2_outputs[3069]);
    assign layer3_outputs[2761] = ~((layer2_outputs[4034]) | (layer2_outputs[4746]));
    assign layer3_outputs[2762] = (layer2_outputs[2057]) & ~(layer2_outputs[4297]);
    assign layer3_outputs[2763] = ~((layer2_outputs[2326]) & (layer2_outputs[1149]));
    assign layer3_outputs[2764] = (layer2_outputs[1934]) | (layer2_outputs[4583]);
    assign layer3_outputs[2765] = (layer2_outputs[3392]) & ~(layer2_outputs[4210]);
    assign layer3_outputs[2766] = (layer2_outputs[2602]) & ~(layer2_outputs[4657]);
    assign layer3_outputs[2767] = (layer2_outputs[3151]) & ~(layer2_outputs[2005]);
    assign layer3_outputs[2768] = layer2_outputs[1705];
    assign layer3_outputs[2769] = ~(layer2_outputs[2060]);
    assign layer3_outputs[2770] = layer2_outputs[4494];
    assign layer3_outputs[2771] = ~(layer2_outputs[385]) | (layer2_outputs[4985]);
    assign layer3_outputs[2772] = (layer2_outputs[1649]) & ~(layer2_outputs[3157]);
    assign layer3_outputs[2773] = ~(layer2_outputs[1215]);
    assign layer3_outputs[2774] = 1'b0;
    assign layer3_outputs[2775] = layer2_outputs[2422];
    assign layer3_outputs[2776] = ~((layer2_outputs[775]) & (layer2_outputs[4734]));
    assign layer3_outputs[2777] = ~((layer2_outputs[4521]) | (layer2_outputs[1027]));
    assign layer3_outputs[2778] = 1'b0;
    assign layer3_outputs[2779] = layer2_outputs[3993];
    assign layer3_outputs[2780] = layer2_outputs[1596];
    assign layer3_outputs[2781] = ~((layer2_outputs[2579]) | (layer2_outputs[4941]));
    assign layer3_outputs[2782] = layer2_outputs[2183];
    assign layer3_outputs[2783] = 1'b1;
    assign layer3_outputs[2784] = (layer2_outputs[2456]) | (layer2_outputs[1615]);
    assign layer3_outputs[2785] = ~(layer2_outputs[2289]) | (layer2_outputs[597]);
    assign layer3_outputs[2786] = ~(layer2_outputs[1533]);
    assign layer3_outputs[2787] = (layer2_outputs[2212]) & (layer2_outputs[4924]);
    assign layer3_outputs[2788] = layer2_outputs[4248];
    assign layer3_outputs[2789] = ~(layer2_outputs[4559]);
    assign layer3_outputs[2790] = (layer2_outputs[1917]) ^ (layer2_outputs[2156]);
    assign layer3_outputs[2791] = ~((layer2_outputs[3820]) ^ (layer2_outputs[5052]));
    assign layer3_outputs[2792] = ~(layer2_outputs[1856]);
    assign layer3_outputs[2793] = layer2_outputs[1869];
    assign layer3_outputs[2794] = ~((layer2_outputs[2319]) | (layer2_outputs[3782]));
    assign layer3_outputs[2795] = layer2_outputs[2792];
    assign layer3_outputs[2796] = layer2_outputs[1209];
    assign layer3_outputs[2797] = ~((layer2_outputs[4819]) & (layer2_outputs[2821]));
    assign layer3_outputs[2798] = ~(layer2_outputs[3558]) | (layer2_outputs[1711]);
    assign layer3_outputs[2799] = 1'b1;
    assign layer3_outputs[2800] = layer2_outputs[2190];
    assign layer3_outputs[2801] = ~((layer2_outputs[2851]) | (layer2_outputs[682]));
    assign layer3_outputs[2802] = layer2_outputs[5094];
    assign layer3_outputs[2803] = (layer2_outputs[2595]) & ~(layer2_outputs[1090]);
    assign layer3_outputs[2804] = layer2_outputs[992];
    assign layer3_outputs[2805] = ~(layer2_outputs[2034]);
    assign layer3_outputs[2806] = ~((layer2_outputs[2840]) | (layer2_outputs[4825]));
    assign layer3_outputs[2807] = 1'b0;
    assign layer3_outputs[2808] = 1'b1;
    assign layer3_outputs[2809] = (layer2_outputs[709]) & (layer2_outputs[2751]);
    assign layer3_outputs[2810] = (layer2_outputs[4372]) & ~(layer2_outputs[1456]);
    assign layer3_outputs[2811] = 1'b1;
    assign layer3_outputs[2812] = (layer2_outputs[3144]) & ~(layer2_outputs[4013]);
    assign layer3_outputs[2813] = 1'b1;
    assign layer3_outputs[2814] = layer2_outputs[1200];
    assign layer3_outputs[2815] = (layer2_outputs[723]) ^ (layer2_outputs[4434]);
    assign layer3_outputs[2816] = ~((layer2_outputs[2343]) & (layer2_outputs[3680]));
    assign layer3_outputs[2817] = ~(layer2_outputs[2859]) | (layer2_outputs[4524]);
    assign layer3_outputs[2818] = ~(layer2_outputs[2794]) | (layer2_outputs[2849]);
    assign layer3_outputs[2819] = ~(layer2_outputs[1520]) | (layer2_outputs[4903]);
    assign layer3_outputs[2820] = layer2_outputs[2624];
    assign layer3_outputs[2821] = ~(layer2_outputs[1971]);
    assign layer3_outputs[2822] = (layer2_outputs[166]) | (layer2_outputs[3260]);
    assign layer3_outputs[2823] = (layer2_outputs[4682]) | (layer2_outputs[1506]);
    assign layer3_outputs[2824] = ~((layer2_outputs[1289]) & (layer2_outputs[2844]));
    assign layer3_outputs[2825] = (layer2_outputs[4194]) ^ (layer2_outputs[559]);
    assign layer3_outputs[2826] = 1'b0;
    assign layer3_outputs[2827] = (layer2_outputs[2901]) & (layer2_outputs[4993]);
    assign layer3_outputs[2828] = 1'b1;
    assign layer3_outputs[2829] = (layer2_outputs[1327]) & ~(layer2_outputs[4189]);
    assign layer3_outputs[2830] = (layer2_outputs[4085]) & ~(layer2_outputs[4376]);
    assign layer3_outputs[2831] = ~((layer2_outputs[2194]) | (layer2_outputs[4244]));
    assign layer3_outputs[2832] = ~(layer2_outputs[4900]) | (layer2_outputs[3235]);
    assign layer3_outputs[2833] = ~(layer2_outputs[327]) | (layer2_outputs[827]);
    assign layer3_outputs[2834] = (layer2_outputs[4273]) | (layer2_outputs[2135]);
    assign layer3_outputs[2835] = (layer2_outputs[1144]) | (layer2_outputs[3487]);
    assign layer3_outputs[2836] = layer2_outputs[200];
    assign layer3_outputs[2837] = (layer2_outputs[2045]) & (layer2_outputs[2195]);
    assign layer3_outputs[2838] = ~(layer2_outputs[1544]);
    assign layer3_outputs[2839] = 1'b1;
    assign layer3_outputs[2840] = ~(layer2_outputs[2182]);
    assign layer3_outputs[2841] = ~((layer2_outputs[2929]) ^ (layer2_outputs[4265]));
    assign layer3_outputs[2842] = layer2_outputs[2606];
    assign layer3_outputs[2843] = ~(layer2_outputs[4844]) | (layer2_outputs[1894]);
    assign layer3_outputs[2844] = ~(layer2_outputs[3899]) | (layer2_outputs[4176]);
    assign layer3_outputs[2845] = ~(layer2_outputs[2584]);
    assign layer3_outputs[2846] = ~(layer2_outputs[4806]) | (layer2_outputs[3131]);
    assign layer3_outputs[2847] = ~(layer2_outputs[4257]);
    assign layer3_outputs[2848] = (layer2_outputs[624]) & ~(layer2_outputs[2740]);
    assign layer3_outputs[2849] = ~(layer2_outputs[3743]);
    assign layer3_outputs[2850] = layer2_outputs[877];
    assign layer3_outputs[2851] = 1'b1;
    assign layer3_outputs[2852] = ~(layer2_outputs[1603]);
    assign layer3_outputs[2853] = (layer2_outputs[1940]) | (layer2_outputs[2572]);
    assign layer3_outputs[2854] = layer2_outputs[4280];
    assign layer3_outputs[2855] = ~((layer2_outputs[1379]) | (layer2_outputs[1550]));
    assign layer3_outputs[2856] = ~(layer2_outputs[780]) | (layer2_outputs[1625]);
    assign layer3_outputs[2857] = ~(layer2_outputs[3622]) | (layer2_outputs[95]);
    assign layer3_outputs[2858] = 1'b1;
    assign layer3_outputs[2859] = ~((layer2_outputs[4642]) | (layer2_outputs[617]));
    assign layer3_outputs[2860] = layer2_outputs[5061];
    assign layer3_outputs[2861] = ~(layer2_outputs[2067]);
    assign layer3_outputs[2862] = ~((layer2_outputs[3102]) | (layer2_outputs[498]));
    assign layer3_outputs[2863] = ~(layer2_outputs[4291]);
    assign layer3_outputs[2864] = ~(layer2_outputs[5064]);
    assign layer3_outputs[2865] = 1'b1;
    assign layer3_outputs[2866] = ~(layer2_outputs[2830]) | (layer2_outputs[1004]);
    assign layer3_outputs[2867] = 1'b0;
    assign layer3_outputs[2868] = ~(layer2_outputs[1670]);
    assign layer3_outputs[2869] = ~(layer2_outputs[1020]);
    assign layer3_outputs[2870] = ~(layer2_outputs[220]) | (layer2_outputs[2551]);
    assign layer3_outputs[2871] = (layer2_outputs[4717]) & ~(layer2_outputs[2047]);
    assign layer3_outputs[2872] = (layer2_outputs[1196]) | (layer2_outputs[1065]);
    assign layer3_outputs[2873] = layer2_outputs[1597];
    assign layer3_outputs[2874] = ~(layer2_outputs[4252]) | (layer2_outputs[3510]);
    assign layer3_outputs[2875] = ~(layer2_outputs[4570]);
    assign layer3_outputs[2876] = (layer2_outputs[4517]) & ~(layer2_outputs[5102]);
    assign layer3_outputs[2877] = ~(layer2_outputs[4758]);
    assign layer3_outputs[2878] = ~(layer2_outputs[4516]) | (layer2_outputs[3639]);
    assign layer3_outputs[2879] = layer2_outputs[4088];
    assign layer3_outputs[2880] = ~(layer2_outputs[494]);
    assign layer3_outputs[2881] = 1'b1;
    assign layer3_outputs[2882] = layer2_outputs[3862];
    assign layer3_outputs[2883] = 1'b1;
    assign layer3_outputs[2884] = ~((layer2_outputs[2540]) | (layer2_outputs[2832]));
    assign layer3_outputs[2885] = ~((layer2_outputs[4750]) & (layer2_outputs[3921]));
    assign layer3_outputs[2886] = (layer2_outputs[3160]) & ~(layer2_outputs[1500]);
    assign layer3_outputs[2887] = 1'b0;
    assign layer3_outputs[2888] = ~((layer2_outputs[449]) & (layer2_outputs[1557]));
    assign layer3_outputs[2889] = 1'b0;
    assign layer3_outputs[2890] = ~(layer2_outputs[1296]) | (layer2_outputs[3432]);
    assign layer3_outputs[2891] = (layer2_outputs[2571]) | (layer2_outputs[1156]);
    assign layer3_outputs[2892] = layer2_outputs[1474];
    assign layer3_outputs[2893] = layer2_outputs[3383];
    assign layer3_outputs[2894] = layer2_outputs[1727];
    assign layer3_outputs[2895] = ~(layer2_outputs[1786]) | (layer2_outputs[4544]);
    assign layer3_outputs[2896] = (layer2_outputs[2173]) & (layer2_outputs[3088]);
    assign layer3_outputs[2897] = ~(layer2_outputs[4464]) | (layer2_outputs[162]);
    assign layer3_outputs[2898] = ~((layer2_outputs[4923]) | (layer2_outputs[4794]));
    assign layer3_outputs[2899] = (layer2_outputs[1951]) | (layer2_outputs[3923]);
    assign layer3_outputs[2900] = ~(layer2_outputs[2627]) | (layer2_outputs[4958]);
    assign layer3_outputs[2901] = ~(layer2_outputs[4898]) | (layer2_outputs[3603]);
    assign layer3_outputs[2902] = ~((layer2_outputs[3834]) ^ (layer2_outputs[526]));
    assign layer3_outputs[2903] = (layer2_outputs[812]) | (layer2_outputs[3324]);
    assign layer3_outputs[2904] = ~((layer2_outputs[3954]) & (layer2_outputs[4348]));
    assign layer3_outputs[2905] = layer2_outputs[1584];
    assign layer3_outputs[2906] = ~(layer2_outputs[447]);
    assign layer3_outputs[2907] = ~((layer2_outputs[2807]) & (layer2_outputs[1264]));
    assign layer3_outputs[2908] = ~(layer2_outputs[1045]);
    assign layer3_outputs[2909] = layer2_outputs[2917];
    assign layer3_outputs[2910] = ~(layer2_outputs[1872]) | (layer2_outputs[1954]);
    assign layer3_outputs[2911] = layer2_outputs[1059];
    assign layer3_outputs[2912] = (layer2_outputs[1300]) & ~(layer2_outputs[2888]);
    assign layer3_outputs[2913] = ~(layer2_outputs[1794]);
    assign layer3_outputs[2914] = ~(layer2_outputs[4288]);
    assign layer3_outputs[2915] = layer2_outputs[1979];
    assign layer3_outputs[2916] = layer2_outputs[429];
    assign layer3_outputs[2917] = (layer2_outputs[4509]) & ~(layer2_outputs[5070]);
    assign layer3_outputs[2918] = layer2_outputs[1564];
    assign layer3_outputs[2919] = ~(layer2_outputs[4439]);
    assign layer3_outputs[2920] = (layer2_outputs[4767]) & ~(layer2_outputs[3630]);
    assign layer3_outputs[2921] = (layer2_outputs[2049]) ^ (layer2_outputs[1193]);
    assign layer3_outputs[2922] = ~(layer2_outputs[4382]);
    assign layer3_outputs[2923] = ~(layer2_outputs[2368]) | (layer2_outputs[2057]);
    assign layer3_outputs[2924] = 1'b0;
    assign layer3_outputs[2925] = ~(layer2_outputs[4735]);
    assign layer3_outputs[2926] = (layer2_outputs[4685]) & (layer2_outputs[317]);
    assign layer3_outputs[2927] = layer2_outputs[3042];
    assign layer3_outputs[2928] = layer2_outputs[666];
    assign layer3_outputs[2929] = ~(layer2_outputs[445]) | (layer2_outputs[1429]);
    assign layer3_outputs[2930] = 1'b0;
    assign layer3_outputs[2931] = ~((layer2_outputs[4409]) & (layer2_outputs[1198]));
    assign layer3_outputs[2932] = 1'b0;
    assign layer3_outputs[2933] = ~(layer2_outputs[4481]);
    assign layer3_outputs[2934] = ~(layer2_outputs[20]) | (layer2_outputs[2370]);
    assign layer3_outputs[2935] = ~(layer2_outputs[2991]);
    assign layer3_outputs[2936] = ~(layer2_outputs[38]) | (layer2_outputs[405]);
    assign layer3_outputs[2937] = layer2_outputs[2745];
    assign layer3_outputs[2938] = ~(layer2_outputs[4600]);
    assign layer3_outputs[2939] = (layer2_outputs[716]) | (layer2_outputs[3588]);
    assign layer3_outputs[2940] = (layer2_outputs[1580]) & ~(layer2_outputs[4121]);
    assign layer3_outputs[2941] = layer2_outputs[2729];
    assign layer3_outputs[2942] = layer2_outputs[1733];
    assign layer3_outputs[2943] = layer2_outputs[209];
    assign layer3_outputs[2944] = ~((layer2_outputs[373]) ^ (layer2_outputs[4649]));
    assign layer3_outputs[2945] = ~(layer2_outputs[4568]);
    assign layer3_outputs[2946] = ~(layer2_outputs[3804]) | (layer2_outputs[5077]);
    assign layer3_outputs[2947] = ~(layer2_outputs[842]) | (layer2_outputs[4946]);
    assign layer3_outputs[2948] = layer2_outputs[2846];
    assign layer3_outputs[2949] = layer2_outputs[964];
    assign layer3_outputs[2950] = (layer2_outputs[3870]) | (layer2_outputs[619]);
    assign layer3_outputs[2951] = (layer2_outputs[3108]) & ~(layer2_outputs[965]);
    assign layer3_outputs[2952] = ~(layer2_outputs[2708]);
    assign layer3_outputs[2953] = layer2_outputs[2784];
    assign layer3_outputs[2954] = ~(layer2_outputs[3855]) | (layer2_outputs[3659]);
    assign layer3_outputs[2955] = ~((layer2_outputs[1251]) | (layer2_outputs[4555]));
    assign layer3_outputs[2956] = layer2_outputs[3789];
    assign layer3_outputs[2957] = ~((layer2_outputs[3451]) ^ (layer2_outputs[3678]));
    assign layer3_outputs[2958] = (layer2_outputs[2000]) & ~(layer2_outputs[3960]);
    assign layer3_outputs[2959] = ~((layer2_outputs[3511]) & (layer2_outputs[3935]));
    assign layer3_outputs[2960] = (layer2_outputs[3318]) & ~(layer2_outputs[4418]);
    assign layer3_outputs[2961] = ~(layer2_outputs[4175]);
    assign layer3_outputs[2962] = layer2_outputs[3093];
    assign layer3_outputs[2963] = ~((layer2_outputs[458]) & (layer2_outputs[1715]));
    assign layer3_outputs[2964] = layer2_outputs[5013];
    assign layer3_outputs[2965] = layer2_outputs[3424];
    assign layer3_outputs[2966] = ~(layer2_outputs[2360]);
    assign layer3_outputs[2967] = ~((layer2_outputs[3192]) & (layer2_outputs[4398]));
    assign layer3_outputs[2968] = layer2_outputs[3290];
    assign layer3_outputs[2969] = ~(layer2_outputs[2338]);
    assign layer3_outputs[2970] = layer2_outputs[1426];
    assign layer3_outputs[2971] = ~(layer2_outputs[2008]) | (layer2_outputs[2600]);
    assign layer3_outputs[2972] = layer2_outputs[1785];
    assign layer3_outputs[2973] = ~(layer2_outputs[2349]);
    assign layer3_outputs[2974] = layer2_outputs[601];
    assign layer3_outputs[2975] = (layer2_outputs[3407]) & ~(layer2_outputs[3010]);
    assign layer3_outputs[2976] = (layer2_outputs[4316]) & ~(layer2_outputs[4857]);
    assign layer3_outputs[2977] = 1'b0;
    assign layer3_outputs[2978] = layer2_outputs[2330];
    assign layer3_outputs[2979] = ~(layer2_outputs[2565]) | (layer2_outputs[2457]);
    assign layer3_outputs[2980] = ~(layer2_outputs[142]);
    assign layer3_outputs[2981] = ~(layer2_outputs[4759]);
    assign layer3_outputs[2982] = ~(layer2_outputs[6]) | (layer2_outputs[3225]);
    assign layer3_outputs[2983] = ~(layer2_outputs[836]) | (layer2_outputs[3946]);
    assign layer3_outputs[2984] = ~((layer2_outputs[2201]) & (layer2_outputs[3550]));
    assign layer3_outputs[2985] = ~((layer2_outputs[1953]) | (layer2_outputs[4913]));
    assign layer3_outputs[2986] = 1'b1;
    assign layer3_outputs[2987] = (layer2_outputs[2722]) & (layer2_outputs[1316]);
    assign layer3_outputs[2988] = layer2_outputs[1833];
    assign layer3_outputs[2989] = 1'b1;
    assign layer3_outputs[2990] = ~((layer2_outputs[3987]) & (layer2_outputs[2250]));
    assign layer3_outputs[2991] = ~(layer2_outputs[270]);
    assign layer3_outputs[2992] = layer2_outputs[4652];
    assign layer3_outputs[2993] = layer2_outputs[2721];
    assign layer3_outputs[2994] = (layer2_outputs[1795]) & ~(layer2_outputs[5012]);
    assign layer3_outputs[2995] = ~(layer2_outputs[873]);
    assign layer3_outputs[2996] = (layer2_outputs[3200]) & (layer2_outputs[1775]);
    assign layer3_outputs[2997] = ~(layer2_outputs[1128]) | (layer2_outputs[3338]);
    assign layer3_outputs[2998] = (layer2_outputs[3803]) & (layer2_outputs[1717]);
    assign layer3_outputs[2999] = (layer2_outputs[2732]) & ~(layer2_outputs[1235]);
    assign layer3_outputs[3000] = ~(layer2_outputs[2984]);
    assign layer3_outputs[3001] = (layer2_outputs[2632]) & ~(layer2_outputs[4009]);
    assign layer3_outputs[3002] = (layer2_outputs[3982]) & ~(layer2_outputs[1049]);
    assign layer3_outputs[3003] = ~(layer2_outputs[2248]);
    assign layer3_outputs[3004] = (layer2_outputs[1223]) & ~(layer2_outputs[3022]);
    assign layer3_outputs[3005] = ~((layer2_outputs[2993]) & (layer2_outputs[2635]));
    assign layer3_outputs[3006] = ~((layer2_outputs[3184]) & (layer2_outputs[2483]));
    assign layer3_outputs[3007] = 1'b1;
    assign layer3_outputs[3008] = 1'b0;
    assign layer3_outputs[3009] = ~(layer2_outputs[4769]);
    assign layer3_outputs[3010] = (layer2_outputs[4020]) | (layer2_outputs[3644]);
    assign layer3_outputs[3011] = 1'b0;
    assign layer3_outputs[3012] = (layer2_outputs[2683]) | (layer2_outputs[4782]);
    assign layer3_outputs[3013] = ~(layer2_outputs[362]) | (layer2_outputs[3913]);
    assign layer3_outputs[3014] = ~((layer2_outputs[3444]) | (layer2_outputs[931]));
    assign layer3_outputs[3015] = 1'b0;
    assign layer3_outputs[3016] = (layer2_outputs[120]) & (layer2_outputs[3081]);
    assign layer3_outputs[3017] = (layer2_outputs[3694]) | (layer2_outputs[4251]);
    assign layer3_outputs[3018] = ~((layer2_outputs[848]) | (layer2_outputs[2653]));
    assign layer3_outputs[3019] = (layer2_outputs[2358]) & ~(layer2_outputs[2663]);
    assign layer3_outputs[3020] = (layer2_outputs[2686]) & (layer2_outputs[768]);
    assign layer3_outputs[3021] = 1'b1;
    assign layer3_outputs[3022] = (layer2_outputs[4295]) | (layer2_outputs[3682]);
    assign layer3_outputs[3023] = ~(layer2_outputs[744]);
    assign layer3_outputs[3024] = (layer2_outputs[3948]) | (layer2_outputs[3442]);
    assign layer3_outputs[3025] = (layer2_outputs[1776]) | (layer2_outputs[4050]);
    assign layer3_outputs[3026] = layer2_outputs[1342];
    assign layer3_outputs[3027] = layer2_outputs[91];
    assign layer3_outputs[3028] = ~(layer2_outputs[1788]);
    assign layer3_outputs[3029] = 1'b0;
    assign layer3_outputs[3030] = ~(layer2_outputs[779]);
    assign layer3_outputs[3031] = layer2_outputs[2019];
    assign layer3_outputs[3032] = (layer2_outputs[1302]) & (layer2_outputs[4694]);
    assign layer3_outputs[3033] = 1'b1;
    assign layer3_outputs[3034] = (layer2_outputs[2692]) & ~(layer2_outputs[1910]);
    assign layer3_outputs[3035] = ~(layer2_outputs[3242]);
    assign layer3_outputs[3036] = (layer2_outputs[4614]) ^ (layer2_outputs[615]);
    assign layer3_outputs[3037] = ~((layer2_outputs[3823]) ^ (layer2_outputs[662]));
    assign layer3_outputs[3038] = layer2_outputs[4092];
    assign layer3_outputs[3039] = (layer2_outputs[1488]) | (layer2_outputs[3531]);
    assign layer3_outputs[3040] = layer2_outputs[4146];
    assign layer3_outputs[3041] = 1'b1;
    assign layer3_outputs[3042] = ~((layer2_outputs[1853]) | (layer2_outputs[1721]));
    assign layer3_outputs[3043] = layer2_outputs[3601];
    assign layer3_outputs[3044] = 1'b0;
    assign layer3_outputs[3045] = ~(layer2_outputs[1609]) | (layer2_outputs[771]);
    assign layer3_outputs[3046] = layer2_outputs[2549];
    assign layer3_outputs[3047] = 1'b0;
    assign layer3_outputs[3048] = layer2_outputs[5074];
    assign layer3_outputs[3049] = ~(layer2_outputs[4455]) | (layer2_outputs[1906]);
    assign layer3_outputs[3050] = (layer2_outputs[1748]) & ~(layer2_outputs[2811]);
    assign layer3_outputs[3051] = ~(layer2_outputs[5045]) | (layer2_outputs[950]);
    assign layer3_outputs[3052] = ~((layer2_outputs[1221]) | (layer2_outputs[423]));
    assign layer3_outputs[3053] = layer2_outputs[3603];
    assign layer3_outputs[3054] = ~(layer2_outputs[4322]);
    assign layer3_outputs[3055] = ~(layer2_outputs[555]) | (layer2_outputs[2678]);
    assign layer3_outputs[3056] = layer2_outputs[1086];
    assign layer3_outputs[3057] = 1'b0;
    assign layer3_outputs[3058] = layer2_outputs[2219];
    assign layer3_outputs[3059] = (layer2_outputs[3760]) ^ (layer2_outputs[725]);
    assign layer3_outputs[3060] = layer2_outputs[772];
    assign layer3_outputs[3061] = ~((layer2_outputs[2522]) | (layer2_outputs[2255]));
    assign layer3_outputs[3062] = ~((layer2_outputs[2121]) | (layer2_outputs[159]));
    assign layer3_outputs[3063] = ~(layer2_outputs[2327]) | (layer2_outputs[2394]);
    assign layer3_outputs[3064] = layer2_outputs[2563];
    assign layer3_outputs[3065] = ~(layer2_outputs[334]) | (layer2_outputs[709]);
    assign layer3_outputs[3066] = 1'b1;
    assign layer3_outputs[3067] = 1'b1;
    assign layer3_outputs[3068] = ~((layer2_outputs[1808]) & (layer2_outputs[3872]));
    assign layer3_outputs[3069] = (layer2_outputs[2845]) | (layer2_outputs[1503]);
    assign layer3_outputs[3070] = layer2_outputs[3753];
    assign layer3_outputs[3071] = ~((layer2_outputs[519]) & (layer2_outputs[2910]));
    assign layer3_outputs[3072] = ~((layer2_outputs[4773]) ^ (layer2_outputs[2384]));
    assign layer3_outputs[3073] = (layer2_outputs[3707]) & ~(layer2_outputs[4135]);
    assign layer3_outputs[3074] = layer2_outputs[3020];
    assign layer3_outputs[3075] = layer2_outputs[1001];
    assign layer3_outputs[3076] = (layer2_outputs[2690]) ^ (layer2_outputs[279]);
    assign layer3_outputs[3077] = (layer2_outputs[2665]) & ~(layer2_outputs[1079]);
    assign layer3_outputs[3078] = ~(layer2_outputs[2331]) | (layer2_outputs[3002]);
    assign layer3_outputs[3079] = ~(layer2_outputs[4270]);
    assign layer3_outputs[3080] = (layer2_outputs[1814]) & ~(layer2_outputs[2628]);
    assign layer3_outputs[3081] = (layer2_outputs[2709]) | (layer2_outputs[4344]);
    assign layer3_outputs[3082] = ~((layer2_outputs[1465]) | (layer2_outputs[1344]));
    assign layer3_outputs[3083] = (layer2_outputs[2134]) & ~(layer2_outputs[5090]);
    assign layer3_outputs[3084] = (layer2_outputs[4245]) & (layer2_outputs[3346]);
    assign layer3_outputs[3085] = ~(layer2_outputs[3496]);
    assign layer3_outputs[3086] = layer2_outputs[1494];
    assign layer3_outputs[3087] = (layer2_outputs[178]) & ~(layer2_outputs[3707]);
    assign layer3_outputs[3088] = ~(layer2_outputs[2095]) | (layer2_outputs[1245]);
    assign layer3_outputs[3089] = ~(layer2_outputs[2697]);
    assign layer3_outputs[3090] = (layer2_outputs[3662]) & ~(layer2_outputs[413]);
    assign layer3_outputs[3091] = (layer2_outputs[2736]) & ~(layer2_outputs[3579]);
    assign layer3_outputs[3092] = (layer2_outputs[4363]) & ~(layer2_outputs[3805]);
    assign layer3_outputs[3093] = 1'b1;
    assign layer3_outputs[3094] = ~(layer2_outputs[3683]);
    assign layer3_outputs[3095] = 1'b0;
    assign layer3_outputs[3096] = ~((layer2_outputs[1435]) | (layer2_outputs[275]));
    assign layer3_outputs[3097] = (layer2_outputs[4679]) & (layer2_outputs[921]);
    assign layer3_outputs[3098] = ~(layer2_outputs[553]);
    assign layer3_outputs[3099] = ~(layer2_outputs[280]);
    assign layer3_outputs[3100] = ~(layer2_outputs[4117]);
    assign layer3_outputs[3101] = 1'b0;
    assign layer3_outputs[3102] = (layer2_outputs[2258]) & (layer2_outputs[3450]);
    assign layer3_outputs[3103] = 1'b1;
    assign layer3_outputs[3104] = ~(layer2_outputs[2783]) | (layer2_outputs[2836]);
    assign layer3_outputs[3105] = (layer2_outputs[3005]) & (layer2_outputs[1229]);
    assign layer3_outputs[3106] = layer2_outputs[4046];
    assign layer3_outputs[3107] = 1'b1;
    assign layer3_outputs[3108] = layer2_outputs[428];
    assign layer3_outputs[3109] = ~((layer2_outputs[3569]) & (layer2_outputs[786]));
    assign layer3_outputs[3110] = ~(layer2_outputs[3833]);
    assign layer3_outputs[3111] = (layer2_outputs[4921]) & ~(layer2_outputs[1548]);
    assign layer3_outputs[3112] = (layer2_outputs[2996]) & (layer2_outputs[3713]);
    assign layer3_outputs[3113] = (layer2_outputs[4743]) & (layer2_outputs[4804]);
    assign layer3_outputs[3114] = layer2_outputs[2404];
    assign layer3_outputs[3115] = ~(layer2_outputs[4591]) | (layer2_outputs[1650]);
    assign layer3_outputs[3116] = ~(layer2_outputs[1347]);
    assign layer3_outputs[3117] = ~((layer2_outputs[4090]) & (layer2_outputs[1389]));
    assign layer3_outputs[3118] = 1'b1;
    assign layer3_outputs[3119] = 1'b0;
    assign layer3_outputs[3120] = (layer2_outputs[2541]) & ~(layer2_outputs[551]);
    assign layer3_outputs[3121] = (layer2_outputs[1186]) & ~(layer2_outputs[2127]);
    assign layer3_outputs[3122] = 1'b0;
    assign layer3_outputs[3123] = layer2_outputs[4788];
    assign layer3_outputs[3124] = ~(layer2_outputs[4844]);
    assign layer3_outputs[3125] = ~(layer2_outputs[2881]) | (layer2_outputs[2468]);
    assign layer3_outputs[3126] = 1'b1;
    assign layer3_outputs[3127] = (layer2_outputs[4246]) & (layer2_outputs[2443]);
    assign layer3_outputs[3128] = ~(layer2_outputs[1539]) | (layer2_outputs[2371]);
    assign layer3_outputs[3129] = ~(layer2_outputs[3902]);
    assign layer3_outputs[3130] = layer2_outputs[763];
    assign layer3_outputs[3131] = layer2_outputs[1582];
    assign layer3_outputs[3132] = (layer2_outputs[5096]) & ~(layer2_outputs[750]);
    assign layer3_outputs[3133] = (layer2_outputs[5091]) & ~(layer2_outputs[2606]);
    assign layer3_outputs[3134] = (layer2_outputs[3078]) ^ (layer2_outputs[4654]);
    assign layer3_outputs[3135] = layer2_outputs[124];
    assign layer3_outputs[3136] = (layer2_outputs[2623]) & ~(layer2_outputs[4848]);
    assign layer3_outputs[3137] = layer2_outputs[2070];
    assign layer3_outputs[3138] = ~(layer2_outputs[4109]);
    assign layer3_outputs[3139] = layer2_outputs[833];
    assign layer3_outputs[3140] = (layer2_outputs[717]) & ~(layer2_outputs[3435]);
    assign layer3_outputs[3141] = (layer2_outputs[3160]) & (layer2_outputs[3105]);
    assign layer3_outputs[3142] = (layer2_outputs[2671]) & ~(layer2_outputs[2595]);
    assign layer3_outputs[3143] = (layer2_outputs[1642]) & (layer2_outputs[2348]);
    assign layer3_outputs[3144] = 1'b0;
    assign layer3_outputs[3145] = layer2_outputs[671];
    assign layer3_outputs[3146] = ~(layer2_outputs[1507]);
    assign layer3_outputs[3147] = layer2_outputs[2533];
    assign layer3_outputs[3148] = layer2_outputs[3470];
    assign layer3_outputs[3149] = ~((layer2_outputs[2566]) | (layer2_outputs[1116]));
    assign layer3_outputs[3150] = layer2_outputs[2776];
    assign layer3_outputs[3151] = ~(layer2_outputs[3749]);
    assign layer3_outputs[3152] = 1'b0;
    assign layer3_outputs[3153] = ~((layer2_outputs[3159]) | (layer2_outputs[4203]));
    assign layer3_outputs[3154] = ~(layer2_outputs[3205]);
    assign layer3_outputs[3155] = ~((layer2_outputs[1052]) | (layer2_outputs[2883]));
    assign layer3_outputs[3156] = (layer2_outputs[146]) & ~(layer2_outputs[4174]);
    assign layer3_outputs[3157] = ~((layer2_outputs[1091]) & (layer2_outputs[4814]));
    assign layer3_outputs[3158] = 1'b1;
    assign layer3_outputs[3159] = ~(layer2_outputs[4655]);
    assign layer3_outputs[3160] = layer2_outputs[3656];
    assign layer3_outputs[3161] = (layer2_outputs[3977]) & ~(layer2_outputs[3125]);
    assign layer3_outputs[3162] = (layer2_outputs[604]) & (layer2_outputs[3268]);
    assign layer3_outputs[3163] = layer2_outputs[4770];
    assign layer3_outputs[3164] = ~(layer2_outputs[1558]) | (layer2_outputs[1527]);
    assign layer3_outputs[3165] = ~((layer2_outputs[4441]) & (layer2_outputs[1135]));
    assign layer3_outputs[3166] = (layer2_outputs[2711]) | (layer2_outputs[227]);
    assign layer3_outputs[3167] = ~(layer2_outputs[4608]);
    assign layer3_outputs[3168] = layer2_outputs[2119];
    assign layer3_outputs[3169] = ~((layer2_outputs[2873]) & (layer2_outputs[2651]));
    assign layer3_outputs[3170] = ~((layer2_outputs[75]) | (layer2_outputs[1048]));
    assign layer3_outputs[3171] = (layer2_outputs[3985]) | (layer2_outputs[3733]);
    assign layer3_outputs[3172] = ~(layer2_outputs[2911]) | (layer2_outputs[4392]);
    assign layer3_outputs[3173] = (layer2_outputs[422]) | (layer2_outputs[5078]);
    assign layer3_outputs[3174] = ~(layer2_outputs[4745]) | (layer2_outputs[1108]);
    assign layer3_outputs[3175] = 1'b0;
    assign layer3_outputs[3176] = 1'b1;
    assign layer3_outputs[3177] = ~((layer2_outputs[3465]) | (layer2_outputs[4542]));
    assign layer3_outputs[3178] = ~(layer2_outputs[1055]);
    assign layer3_outputs[3179] = (layer2_outputs[2325]) & ~(layer2_outputs[4189]);
    assign layer3_outputs[3180] = ~((layer2_outputs[4032]) & (layer2_outputs[4400]));
    assign layer3_outputs[3181] = ~(layer2_outputs[3868]);
    assign layer3_outputs[3182] = (layer2_outputs[856]) & ~(layer2_outputs[4653]);
    assign layer3_outputs[3183] = ~(layer2_outputs[2752]) | (layer2_outputs[751]);
    assign layer3_outputs[3184] = ~((layer2_outputs[188]) | (layer2_outputs[2120]));
    assign layer3_outputs[3185] = (layer2_outputs[3734]) & (layer2_outputs[2021]);
    assign layer3_outputs[3186] = layer2_outputs[295];
    assign layer3_outputs[3187] = (layer2_outputs[1900]) | (layer2_outputs[36]);
    assign layer3_outputs[3188] = (layer2_outputs[4864]) ^ (layer2_outputs[510]);
    assign layer3_outputs[3189] = (layer2_outputs[3237]) & (layer2_outputs[363]);
    assign layer3_outputs[3190] = (layer2_outputs[2657]) & ~(layer2_outputs[3367]);
    assign layer3_outputs[3191] = 1'b1;
    assign layer3_outputs[3192] = (layer2_outputs[1076]) & (layer2_outputs[1169]);
    assign layer3_outputs[3193] = layer2_outputs[3937];
    assign layer3_outputs[3194] = layer2_outputs[690];
    assign layer3_outputs[3195] = (layer2_outputs[836]) | (layer2_outputs[4162]);
    assign layer3_outputs[3196] = 1'b0;
    assign layer3_outputs[3197] = ~((layer2_outputs[2040]) & (layer2_outputs[5109]));
    assign layer3_outputs[3198] = ~(layer2_outputs[4310]);
    assign layer3_outputs[3199] = ~(layer2_outputs[4470]) | (layer2_outputs[4757]);
    assign layer3_outputs[3200] = 1'b1;
    assign layer3_outputs[3201] = ~((layer2_outputs[4002]) & (layer2_outputs[4920]));
    assign layer3_outputs[3202] = (layer2_outputs[1811]) ^ (layer2_outputs[1970]);
    assign layer3_outputs[3203] = 1'b0;
    assign layer3_outputs[3204] = (layer2_outputs[2047]) & ~(layer2_outputs[1555]);
    assign layer3_outputs[3205] = 1'b0;
    assign layer3_outputs[3206] = 1'b1;
    assign layer3_outputs[3207] = ~(layer2_outputs[3295]);
    assign layer3_outputs[3208] = ~(layer2_outputs[2258]) | (layer2_outputs[4874]);
    assign layer3_outputs[3209] = ~(layer2_outputs[1330]);
    assign layer3_outputs[3210] = ~((layer2_outputs[2407]) & (layer2_outputs[4085]));
    assign layer3_outputs[3211] = layer2_outputs[4365];
    assign layer3_outputs[3212] = layer2_outputs[1102];
    assign layer3_outputs[3213] = ~(layer2_outputs[4315]) | (layer2_outputs[205]);
    assign layer3_outputs[3214] = layer2_outputs[1882];
    assign layer3_outputs[3215] = ~((layer2_outputs[1607]) & (layer2_outputs[4786]));
    assign layer3_outputs[3216] = ~(layer2_outputs[4306]);
    assign layer3_outputs[3217] = (layer2_outputs[486]) & ~(layer2_outputs[1763]);
    assign layer3_outputs[3218] = (layer2_outputs[3540]) ^ (layer2_outputs[1840]);
    assign layer3_outputs[3219] = ~(layer2_outputs[247]) | (layer2_outputs[1746]);
    assign layer3_outputs[3220] = ~(layer2_outputs[3121]);
    assign layer3_outputs[3221] = layer2_outputs[2211];
    assign layer3_outputs[3222] = (layer2_outputs[1942]) & (layer2_outputs[156]);
    assign layer3_outputs[3223] = layer2_outputs[3830];
    assign layer3_outputs[3224] = ~(layer2_outputs[289]) | (layer2_outputs[98]);
    assign layer3_outputs[3225] = ~(layer2_outputs[4394]) | (layer2_outputs[4343]);
    assign layer3_outputs[3226] = layer2_outputs[3930];
    assign layer3_outputs[3227] = ~(layer2_outputs[4630]);
    assign layer3_outputs[3228] = 1'b0;
    assign layer3_outputs[3229] = (layer2_outputs[3039]) ^ (layer2_outputs[4520]);
    assign layer3_outputs[3230] = layer2_outputs[71];
    assign layer3_outputs[3231] = ~(layer2_outputs[70]);
    assign layer3_outputs[3232] = ~((layer2_outputs[1390]) & (layer2_outputs[4580]));
    assign layer3_outputs[3233] = layer2_outputs[1469];
    assign layer3_outputs[3234] = ~(layer2_outputs[2505]);
    assign layer3_outputs[3235] = ~(layer2_outputs[1931]);
    assign layer3_outputs[3236] = (layer2_outputs[1555]) & (layer2_outputs[490]);
    assign layer3_outputs[3237] = ~(layer2_outputs[4675]);
    assign layer3_outputs[3238] = (layer2_outputs[1008]) & ~(layer2_outputs[4868]);
    assign layer3_outputs[3239] = layer2_outputs[1895];
    assign layer3_outputs[3240] = ~(layer2_outputs[2320]);
    assign layer3_outputs[3241] = layer2_outputs[4281];
    assign layer3_outputs[3242] = ~(layer2_outputs[3555]);
    assign layer3_outputs[3243] = ~((layer2_outputs[3578]) & (layer2_outputs[308]));
    assign layer3_outputs[3244] = layer2_outputs[2588];
    assign layer3_outputs[3245] = layer2_outputs[3500];
    assign layer3_outputs[3246] = ~(layer2_outputs[2279]);
    assign layer3_outputs[3247] = layer2_outputs[1861];
    assign layer3_outputs[3248] = 1'b1;
    assign layer3_outputs[3249] = (layer2_outputs[3668]) & ~(layer2_outputs[249]);
    assign layer3_outputs[3250] = ~((layer2_outputs[1695]) | (layer2_outputs[1057]));
    assign layer3_outputs[3251] = layer2_outputs[4942];
    assign layer3_outputs[3252] = ~(layer2_outputs[1605]);
    assign layer3_outputs[3253] = ~(layer2_outputs[2643]);
    assign layer3_outputs[3254] = ~(layer2_outputs[4820]);
    assign layer3_outputs[3255] = ~((layer2_outputs[2175]) & (layer2_outputs[4121]));
    assign layer3_outputs[3256] = 1'b0;
    assign layer3_outputs[3257] = (layer2_outputs[4736]) & ~(layer2_outputs[971]);
    assign layer3_outputs[3258] = (layer2_outputs[2058]) & ~(layer2_outputs[4683]);
    assign layer3_outputs[3259] = layer2_outputs[919];
    assign layer3_outputs[3260] = ~(layer2_outputs[4893]);
    assign layer3_outputs[3261] = (layer2_outputs[265]) & ~(layer2_outputs[3123]);
    assign layer3_outputs[3262] = ~(layer2_outputs[400]);
    assign layer3_outputs[3263] = (layer2_outputs[1928]) | (layer2_outputs[2049]);
    assign layer3_outputs[3264] = ~(layer2_outputs[1489]) | (layer2_outputs[3553]);
    assign layer3_outputs[3265] = (layer2_outputs[3650]) ^ (layer2_outputs[4304]);
    assign layer3_outputs[3266] = ~(layer2_outputs[4733]);
    assign layer3_outputs[3267] = ~((layer2_outputs[1499]) & (layer2_outputs[40]));
    assign layer3_outputs[3268] = (layer2_outputs[3816]) & ~(layer2_outputs[4824]);
    assign layer3_outputs[3269] = (layer2_outputs[2960]) & (layer2_outputs[2240]);
    assign layer3_outputs[3270] = layer2_outputs[827];
    assign layer3_outputs[3271] = layer2_outputs[4882];
    assign layer3_outputs[3272] = ~(layer2_outputs[1270]) | (layer2_outputs[4006]);
    assign layer3_outputs[3273] = (layer2_outputs[3762]) & ~(layer2_outputs[987]);
    assign layer3_outputs[3274] = layer2_outputs[4488];
    assign layer3_outputs[3275] = 1'b0;
    assign layer3_outputs[3276] = layer2_outputs[1774];
    assign layer3_outputs[3277] = ~(layer2_outputs[1676]);
    assign layer3_outputs[3278] = ~(layer2_outputs[522]) | (layer2_outputs[2788]);
    assign layer3_outputs[3279] = (layer2_outputs[3884]) & ~(layer2_outputs[737]);
    assign layer3_outputs[3280] = layer2_outputs[2198];
    assign layer3_outputs[3281] = ~(layer2_outputs[3120]);
    assign layer3_outputs[3282] = layer2_outputs[3136];
    assign layer3_outputs[3283] = ~(layer2_outputs[2065]) | (layer2_outputs[411]);
    assign layer3_outputs[3284] = ~(layer2_outputs[1831]) | (layer2_outputs[133]);
    assign layer3_outputs[3285] = layer2_outputs[3360];
    assign layer3_outputs[3286] = ~(layer2_outputs[2015]);
    assign layer3_outputs[3287] = ~(layer2_outputs[2383]);
    assign layer3_outputs[3288] = ~((layer2_outputs[2728]) & (layer2_outputs[808]));
    assign layer3_outputs[3289] = ~(layer2_outputs[864]);
    assign layer3_outputs[3290] = (layer2_outputs[2395]) | (layer2_outputs[4368]);
    assign layer3_outputs[3291] = layer2_outputs[1110];
    assign layer3_outputs[3292] = 1'b0;
    assign layer3_outputs[3293] = layer2_outputs[4426];
    assign layer3_outputs[3294] = (layer2_outputs[3194]) | (layer2_outputs[1722]);
    assign layer3_outputs[3295] = 1'b1;
    assign layer3_outputs[3296] = (layer2_outputs[4986]) ^ (layer2_outputs[3713]);
    assign layer3_outputs[3297] = ~(layer2_outputs[1107]);
    assign layer3_outputs[3298] = (layer2_outputs[3831]) | (layer2_outputs[2628]);
    assign layer3_outputs[3299] = 1'b1;
    assign layer3_outputs[3300] = ~((layer2_outputs[1756]) & (layer2_outputs[774]));
    assign layer3_outputs[3301] = layer2_outputs[4537];
    assign layer3_outputs[3302] = ~(layer2_outputs[398]);
    assign layer3_outputs[3303] = layer2_outputs[2427];
    assign layer3_outputs[3304] = ~(layer2_outputs[2985]) | (layer2_outputs[1948]);
    assign layer3_outputs[3305] = ~(layer2_outputs[3214]);
    assign layer3_outputs[3306] = (layer2_outputs[387]) & ~(layer2_outputs[565]);
    assign layer3_outputs[3307] = layer2_outputs[2391];
    assign layer3_outputs[3308] = layer2_outputs[2050];
    assign layer3_outputs[3309] = 1'b0;
    assign layer3_outputs[3310] = ~(layer2_outputs[2035]);
    assign layer3_outputs[3311] = (layer2_outputs[3236]) & ~(layer2_outputs[134]);
    assign layer3_outputs[3312] = ~(layer2_outputs[2271]) | (layer2_outputs[393]);
    assign layer3_outputs[3313] = 1'b0;
    assign layer3_outputs[3314] = ~(layer2_outputs[1696]) | (layer2_outputs[743]);
    assign layer3_outputs[3315] = (layer2_outputs[3627]) & ~(layer2_outputs[3118]);
    assign layer3_outputs[3316] = ~(layer2_outputs[3315]);
    assign layer3_outputs[3317] = ~(layer2_outputs[2352]) | (layer2_outputs[2554]);
    assign layer3_outputs[3318] = 1'b1;
    assign layer3_outputs[3319] = (layer2_outputs[4293]) & ~(layer2_outputs[3275]);
    assign layer3_outputs[3320] = (layer2_outputs[911]) & ~(layer2_outputs[2266]);
    assign layer3_outputs[3321] = ~((layer2_outputs[4873]) ^ (layer2_outputs[127]));
    assign layer3_outputs[3322] = layer2_outputs[1393];
    assign layer3_outputs[3323] = (layer2_outputs[978]) & (layer2_outputs[2201]);
    assign layer3_outputs[3324] = (layer2_outputs[1847]) & (layer2_outputs[3167]);
    assign layer3_outputs[3325] = ~(layer2_outputs[3557]);
    assign layer3_outputs[3326] = ~((layer2_outputs[5060]) | (layer2_outputs[3541]));
    assign layer3_outputs[3327] = 1'b0;
    assign layer3_outputs[3328] = ~(layer2_outputs[337]) | (layer2_outputs[2867]);
    assign layer3_outputs[3329] = layer2_outputs[4707];
    assign layer3_outputs[3330] = ~(layer2_outputs[4044]) | (layer2_outputs[661]);
    assign layer3_outputs[3331] = ~((layer2_outputs[3259]) ^ (layer2_outputs[439]));
    assign layer3_outputs[3332] = (layer2_outputs[3937]) & (layer2_outputs[3987]);
    assign layer3_outputs[3333] = ~(layer2_outputs[826]);
    assign layer3_outputs[3334] = ~(layer2_outputs[1035]);
    assign layer3_outputs[3335] = ~(layer2_outputs[1306]);
    assign layer3_outputs[3336] = layer2_outputs[1727];
    assign layer3_outputs[3337] = layer2_outputs[1989];
    assign layer3_outputs[3338] = (layer2_outputs[3836]) & ~(layer2_outputs[3123]);
    assign layer3_outputs[3339] = (layer2_outputs[1324]) & (layer2_outputs[130]);
    assign layer3_outputs[3340] = layer2_outputs[835];
    assign layer3_outputs[3341] = layer2_outputs[251];
    assign layer3_outputs[3342] = ~((layer2_outputs[1329]) & (layer2_outputs[3740]));
    assign layer3_outputs[3343] = 1'b0;
    assign layer3_outputs[3344] = (layer2_outputs[3979]) | (layer2_outputs[2285]);
    assign layer3_outputs[3345] = ~(layer2_outputs[1995]);
    assign layer3_outputs[3346] = (layer2_outputs[3880]) & (layer2_outputs[2970]);
    assign layer3_outputs[3347] = ~(layer2_outputs[3576]);
    assign layer3_outputs[3348] = ~((layer2_outputs[3503]) | (layer2_outputs[809]));
    assign layer3_outputs[3349] = ~((layer2_outputs[4492]) | (layer2_outputs[4576]));
    assign layer3_outputs[3350] = ~(layer2_outputs[400]);
    assign layer3_outputs[3351] = 1'b1;
    assign layer3_outputs[3352] = (layer2_outputs[813]) & ~(layer2_outputs[4540]);
    assign layer3_outputs[3353] = layer2_outputs[2495];
    assign layer3_outputs[3354] = ~((layer2_outputs[5060]) & (layer2_outputs[340]));
    assign layer3_outputs[3355] = (layer2_outputs[4329]) & ~(layer2_outputs[2534]);
    assign layer3_outputs[3356] = ~((layer2_outputs[5099]) & (layer2_outputs[1162]));
    assign layer3_outputs[3357] = ~(layer2_outputs[2192]);
    assign layer3_outputs[3358] = ~(layer2_outputs[1256]) | (layer2_outputs[1786]);
    assign layer3_outputs[3359] = ~(layer2_outputs[2712]);
    assign layer3_outputs[3360] = ~(layer2_outputs[18]);
    assign layer3_outputs[3361] = layer2_outputs[3571];
    assign layer3_outputs[3362] = ~(layer2_outputs[2307]);
    assign layer3_outputs[3363] = ~(layer2_outputs[5087]);
    assign layer3_outputs[3364] = 1'b1;
    assign layer3_outputs[3365] = (layer2_outputs[1865]) & ~(layer2_outputs[5119]);
    assign layer3_outputs[3366] = 1'b1;
    assign layer3_outputs[3367] = ~(layer2_outputs[4714]);
    assign layer3_outputs[3368] = ~(layer2_outputs[5105]);
    assign layer3_outputs[3369] = (layer2_outputs[50]) & (layer2_outputs[1157]);
    assign layer3_outputs[3370] = layer2_outputs[3684];
    assign layer3_outputs[3371] = ~((layer2_outputs[1000]) | (layer2_outputs[4410]));
    assign layer3_outputs[3372] = layer2_outputs[1461];
    assign layer3_outputs[3373] = layer2_outputs[1769];
    assign layer3_outputs[3374] = (layer2_outputs[1309]) & (layer2_outputs[3676]);
    assign layer3_outputs[3375] = 1'b0;
    assign layer3_outputs[3376] = ~((layer2_outputs[999]) | (layer2_outputs[2349]));
    assign layer3_outputs[3377] = (layer2_outputs[810]) & ~(layer2_outputs[3028]);
    assign layer3_outputs[3378] = layer2_outputs[3838];
    assign layer3_outputs[3379] = ~(layer2_outputs[4904]);
    assign layer3_outputs[3380] = layer2_outputs[1900];
    assign layer3_outputs[3381] = ~((layer2_outputs[4595]) ^ (layer2_outputs[31]));
    assign layer3_outputs[3382] = 1'b1;
    assign layer3_outputs[3383] = (layer2_outputs[3670]) & ~(layer2_outputs[2798]);
    assign layer3_outputs[3384] = (layer2_outputs[3565]) | (layer2_outputs[4968]);
    assign layer3_outputs[3385] = ~(layer2_outputs[3305]);
    assign layer3_outputs[3386] = ~(layer2_outputs[4551]);
    assign layer3_outputs[3387] = (layer2_outputs[1374]) & (layer2_outputs[4747]);
    assign layer3_outputs[3388] = (layer2_outputs[408]) & ~(layer2_outputs[2132]);
    assign layer3_outputs[3389] = layer2_outputs[1470];
    assign layer3_outputs[3390] = ~(layer2_outputs[3268]) | (layer2_outputs[2767]);
    assign layer3_outputs[3391] = (layer2_outputs[2791]) | (layer2_outputs[1454]);
    assign layer3_outputs[3392] = layer2_outputs[4847];
    assign layer3_outputs[3393] = ~(layer2_outputs[4219]);
    assign layer3_outputs[3394] = ~(layer2_outputs[2852]) | (layer2_outputs[1866]);
    assign layer3_outputs[3395] = (layer2_outputs[1101]) | (layer2_outputs[4108]);
    assign layer3_outputs[3396] = layer2_outputs[1884];
    assign layer3_outputs[3397] = 1'b1;
    assign layer3_outputs[3398] = layer2_outputs[4301];
    assign layer3_outputs[3399] = ~(layer2_outputs[2409]);
    assign layer3_outputs[3400] = ~(layer2_outputs[4960]);
    assign layer3_outputs[3401] = (layer2_outputs[3923]) & ~(layer2_outputs[1331]);
    assign layer3_outputs[3402] = ~(layer2_outputs[4534]) | (layer2_outputs[959]);
    assign layer3_outputs[3403] = layer2_outputs[2928];
    assign layer3_outputs[3404] = (layer2_outputs[4641]) & ~(layer2_outputs[4668]);
    assign layer3_outputs[3405] = 1'b0;
    assign layer3_outputs[3406] = (layer2_outputs[2767]) & (layer2_outputs[3156]);
    assign layer3_outputs[3407] = ~(layer2_outputs[3829]) | (layer2_outputs[4742]);
    assign layer3_outputs[3408] = (layer2_outputs[4517]) & (layer2_outputs[902]);
    assign layer3_outputs[3409] = ~(layer2_outputs[4986]);
    assign layer3_outputs[3410] = 1'b1;
    assign layer3_outputs[3411] = (layer2_outputs[4856]) & ~(layer2_outputs[2346]);
    assign layer3_outputs[3412] = ~(layer2_outputs[3025]);
    assign layer3_outputs[3413] = 1'b1;
    assign layer3_outputs[3414] = (layer2_outputs[840]) & ~(layer2_outputs[1035]);
    assign layer3_outputs[3415] = ~(layer2_outputs[3116]);
    assign layer3_outputs[3416] = layer2_outputs[1329];
    assign layer3_outputs[3417] = (layer2_outputs[195]) & ~(layer2_outputs[2269]);
    assign layer3_outputs[3418] = ~(layer2_outputs[4880]) | (layer2_outputs[2138]);
    assign layer3_outputs[3419] = ~(layer2_outputs[1978]) | (layer2_outputs[3514]);
    assign layer3_outputs[3420] = ~((layer2_outputs[820]) ^ (layer2_outputs[602]));
    assign layer3_outputs[3421] = ~((layer2_outputs[4388]) & (layer2_outputs[2268]));
    assign layer3_outputs[3422] = ~(layer2_outputs[1807]);
    assign layer3_outputs[3423] = 1'b0;
    assign layer3_outputs[3424] = ~(layer2_outputs[238]);
    assign layer3_outputs[3425] = (layer2_outputs[2473]) & ~(layer2_outputs[2891]);
    assign layer3_outputs[3426] = (layer2_outputs[33]) | (layer2_outputs[4656]);
    assign layer3_outputs[3427] = ~((layer2_outputs[3187]) | (layer2_outputs[335]));
    assign layer3_outputs[3428] = (layer2_outputs[2629]) & ~(layer2_outputs[3128]);
    assign layer3_outputs[3429] = 1'b0;
    assign layer3_outputs[3430] = (layer2_outputs[4999]) | (layer2_outputs[2196]);
    assign layer3_outputs[3431] = ~((layer2_outputs[1981]) | (layer2_outputs[1016]));
    assign layer3_outputs[3432] = ~(layer2_outputs[3532]);
    assign layer3_outputs[3433] = layer2_outputs[1511];
    assign layer3_outputs[3434] = (layer2_outputs[4862]) ^ (layer2_outputs[494]);
    assign layer3_outputs[3435] = (layer2_outputs[2499]) & ~(layer2_outputs[147]);
    assign layer3_outputs[3436] = ~(layer2_outputs[3308]) | (layer2_outputs[4221]);
    assign layer3_outputs[3437] = ~(layer2_outputs[1147]);
    assign layer3_outputs[3438] = (layer2_outputs[4905]) & ~(layer2_outputs[1616]);
    assign layer3_outputs[3439] = ~(layer2_outputs[1870]);
    assign layer3_outputs[3440] = ~(layer2_outputs[3930]);
    assign layer3_outputs[3441] = (layer2_outputs[1318]) & ~(layer2_outputs[4992]);
    assign layer3_outputs[3442] = (layer2_outputs[89]) & ~(layer2_outputs[1204]);
    assign layer3_outputs[3443] = (layer2_outputs[3942]) | (layer2_outputs[4536]);
    assign layer3_outputs[3444] = (layer2_outputs[3405]) & ~(layer2_outputs[2011]);
    assign layer3_outputs[3445] = ~(layer2_outputs[4558]) | (layer2_outputs[628]);
    assign layer3_outputs[3446] = ~(layer2_outputs[3927]);
    assign layer3_outputs[3447] = 1'b1;
    assign layer3_outputs[3448] = ~(layer2_outputs[205]) | (layer2_outputs[1179]);
    assign layer3_outputs[3449] = ~(layer2_outputs[3112]);
    assign layer3_outputs[3450] = ~(layer2_outputs[5095]);
    assign layer3_outputs[3451] = ~(layer2_outputs[2648]) | (layer2_outputs[581]);
    assign layer3_outputs[3452] = (layer2_outputs[3498]) & (layer2_outputs[4721]);
    assign layer3_outputs[3453] = (layer2_outputs[3086]) & ~(layer2_outputs[3033]);
    assign layer3_outputs[3454] = ~(layer2_outputs[1628]);
    assign layer3_outputs[3455] = (layer2_outputs[741]) & (layer2_outputs[5019]);
    assign layer3_outputs[3456] = (layer2_outputs[4772]) & (layer2_outputs[2028]);
    assign layer3_outputs[3457] = ~((layer2_outputs[770]) | (layer2_outputs[2685]));
    assign layer3_outputs[3458] = (layer2_outputs[2331]) | (layer2_outputs[5026]);
    assign layer3_outputs[3459] = (layer2_outputs[2682]) | (layer2_outputs[675]);
    assign layer3_outputs[3460] = ~(layer2_outputs[4105]);
    assign layer3_outputs[3461] = ~(layer2_outputs[1878]) | (layer2_outputs[4888]);
    assign layer3_outputs[3462] = ~((layer2_outputs[2800]) & (layer2_outputs[309]));
    assign layer3_outputs[3463] = (layer2_outputs[1551]) ^ (layer2_outputs[238]);
    assign layer3_outputs[3464] = layer2_outputs[2497];
    assign layer3_outputs[3465] = ~(layer2_outputs[4997]);
    assign layer3_outputs[3466] = ~(layer2_outputs[3771]);
    assign layer3_outputs[3467] = (layer2_outputs[4238]) | (layer2_outputs[712]);
    assign layer3_outputs[3468] = ~(layer2_outputs[1348]);
    assign layer3_outputs[3469] = layer2_outputs[954];
    assign layer3_outputs[3470] = (layer2_outputs[4281]) & ~(layer2_outputs[1920]);
    assign layer3_outputs[3471] = (layer2_outputs[3490]) & ~(layer2_outputs[1442]);
    assign layer3_outputs[3472] = ~((layer2_outputs[216]) ^ (layer2_outputs[3555]));
    assign layer3_outputs[3473] = ~(layer2_outputs[4753]);
    assign layer3_outputs[3474] = (layer2_outputs[436]) & ~(layer2_outputs[4698]);
    assign layer3_outputs[3475] = (layer2_outputs[2981]) & ~(layer2_outputs[3934]);
    assign layer3_outputs[3476] = 1'b1;
    assign layer3_outputs[3477] = layer2_outputs[4959];
    assign layer3_outputs[3478] = ~(layer2_outputs[255]);
    assign layer3_outputs[3479] = layer2_outputs[3699];
    assign layer3_outputs[3480] = (layer2_outputs[1678]) & (layer2_outputs[2344]);
    assign layer3_outputs[3481] = (layer2_outputs[2919]) ^ (layer2_outputs[764]);
    assign layer3_outputs[3482] = 1'b1;
    assign layer3_outputs[3483] = ~(layer2_outputs[3734]) | (layer2_outputs[3810]);
    assign layer3_outputs[3484] = ~(layer2_outputs[482]);
    assign layer3_outputs[3485] = (layer2_outputs[4422]) & ~(layer2_outputs[5097]);
    assign layer3_outputs[3486] = 1'b1;
    assign layer3_outputs[3487] = 1'b0;
    assign layer3_outputs[3488] = ~((layer2_outputs[1095]) ^ (layer2_outputs[3787]));
    assign layer3_outputs[3489] = layer2_outputs[4516];
    assign layer3_outputs[3490] = (layer2_outputs[3959]) & (layer2_outputs[3797]);
    assign layer3_outputs[3491] = (layer2_outputs[2598]) | (layer2_outputs[2437]);
    assign layer3_outputs[3492] = (layer2_outputs[213]) & ~(layer2_outputs[4349]);
    assign layer3_outputs[3493] = ~(layer2_outputs[1906]);
    assign layer3_outputs[3494] = 1'b1;
    assign layer3_outputs[3495] = layer2_outputs[4598];
    assign layer3_outputs[3496] = 1'b1;
    assign layer3_outputs[3497] = 1'b0;
    assign layer3_outputs[3498] = ~(layer2_outputs[3697]);
    assign layer3_outputs[3499] = layer2_outputs[4639];
    assign layer3_outputs[3500] = ~(layer2_outputs[3048]);
    assign layer3_outputs[3501] = ~(layer2_outputs[1631]);
    assign layer3_outputs[3502] = ~(layer2_outputs[3598]);
    assign layer3_outputs[3503] = (layer2_outputs[917]) & ~(layer2_outputs[3130]);
    assign layer3_outputs[3504] = 1'b1;
    assign layer3_outputs[3505] = layer2_outputs[3494];
    assign layer3_outputs[3506] = layer2_outputs[1194];
    assign layer3_outputs[3507] = layer2_outputs[3889];
    assign layer3_outputs[3508] = ~(layer2_outputs[22]) | (layer2_outputs[3765]);
    assign layer3_outputs[3509] = (layer2_outputs[2094]) & (layer2_outputs[1310]);
    assign layer3_outputs[3510] = ~((layer2_outputs[4843]) ^ (layer2_outputs[2815]));
    assign layer3_outputs[3511] = ~((layer2_outputs[3764]) | (layer2_outputs[2304]));
    assign layer3_outputs[3512] = ~(layer2_outputs[1326]);
    assign layer3_outputs[3513] = ~(layer2_outputs[276]);
    assign layer3_outputs[3514] = (layer2_outputs[2411]) | (layer2_outputs[4450]);
    assign layer3_outputs[3515] = layer2_outputs[2362];
    assign layer3_outputs[3516] = (layer2_outputs[442]) & (layer2_outputs[510]);
    assign layer3_outputs[3517] = (layer2_outputs[1770]) & ~(layer2_outputs[1709]);
    assign layer3_outputs[3518] = ~(layer2_outputs[426]);
    assign layer3_outputs[3519] = (layer2_outputs[676]) & ~(layer2_outputs[4401]);
    assign layer3_outputs[3520] = (layer2_outputs[2400]) & ~(layer2_outputs[3401]);
    assign layer3_outputs[3521] = layer2_outputs[1482];
    assign layer3_outputs[3522] = (layer2_outputs[3471]) & ~(layer2_outputs[4342]);
    assign layer3_outputs[3523] = ~(layer2_outputs[2736]) | (layer2_outputs[2930]);
    assign layer3_outputs[3524] = 1'b0;
    assign layer3_outputs[3525] = ~((layer2_outputs[981]) | (layer2_outputs[1623]));
    assign layer3_outputs[3526] = 1'b0;
    assign layer3_outputs[3527] = (layer2_outputs[4142]) & (layer2_outputs[4498]);
    assign layer3_outputs[3528] = ~(layer2_outputs[434]);
    assign layer3_outputs[3529] = (layer2_outputs[3172]) | (layer2_outputs[3216]);
    assign layer3_outputs[3530] = ~((layer2_outputs[385]) & (layer2_outputs[4161]));
    assign layer3_outputs[3531] = ~(layer2_outputs[2571]);
    assign layer3_outputs[3532] = (layer2_outputs[2621]) | (layer2_outputs[2256]);
    assign layer3_outputs[3533] = 1'b0;
    assign layer3_outputs[3534] = layer2_outputs[104];
    assign layer3_outputs[3535] = ~(layer2_outputs[4805]);
    assign layer3_outputs[3536] = (layer2_outputs[453]) ^ (layer2_outputs[4019]);
    assign layer3_outputs[3537] = layer2_outputs[1113];
    assign layer3_outputs[3538] = ~((layer2_outputs[997]) | (layer2_outputs[1305]));
    assign layer3_outputs[3539] = (layer2_outputs[2557]) & (layer2_outputs[1018]);
    assign layer3_outputs[3540] = ~((layer2_outputs[3327]) & (layer2_outputs[1439]));
    assign layer3_outputs[3541] = ~(layer2_outputs[4991]);
    assign layer3_outputs[3542] = ~(layer2_outputs[2729]);
    assign layer3_outputs[3543] = ~(layer2_outputs[734]);
    assign layer3_outputs[3544] = (layer2_outputs[701]) & (layer2_outputs[3247]);
    assign layer3_outputs[3545] = (layer2_outputs[3963]) | (layer2_outputs[3727]);
    assign layer3_outputs[3546] = (layer2_outputs[2526]) ^ (layer2_outputs[837]);
    assign layer3_outputs[3547] = ~(layer2_outputs[1527]);
    assign layer3_outputs[3548] = (layer2_outputs[2108]) & ~(layer2_outputs[2952]);
    assign layer3_outputs[3549] = layer2_outputs[721];
    assign layer3_outputs[3550] = layer2_outputs[1146];
    assign layer3_outputs[3551] = (layer2_outputs[4602]) & (layer2_outputs[4279]);
    assign layer3_outputs[3552] = layer2_outputs[4486];
    assign layer3_outputs[3553] = ~(layer2_outputs[4293]);
    assign layer3_outputs[3554] = layer2_outputs[2256];
    assign layer3_outputs[3555] = layer2_outputs[4700];
    assign layer3_outputs[3556] = layer2_outputs[1748];
    assign layer3_outputs[3557] = ~(layer2_outputs[2310]);
    assign layer3_outputs[3558] = 1'b1;
    assign layer3_outputs[3559] = ~(layer2_outputs[1283]);
    assign layer3_outputs[3560] = ~(layer2_outputs[4804]);
    assign layer3_outputs[3561] = (layer2_outputs[2778]) & ~(layer2_outputs[491]);
    assign layer3_outputs[3562] = layer2_outputs[4200];
    assign layer3_outputs[3563] = (layer2_outputs[2760]) | (layer2_outputs[4872]);
    assign layer3_outputs[3564] = 1'b0;
    assign layer3_outputs[3565] = ~((layer2_outputs[830]) & (layer2_outputs[1237]));
    assign layer3_outputs[3566] = layer2_outputs[958];
    assign layer3_outputs[3567] = (layer2_outputs[3982]) & ~(layer2_outputs[654]);
    assign layer3_outputs[3568] = ~(layer2_outputs[4687]);
    assign layer3_outputs[3569] = ~(layer2_outputs[1575]);
    assign layer3_outputs[3570] = ~(layer2_outputs[3491]);
    assign layer3_outputs[3571] = layer2_outputs[3211];
    assign layer3_outputs[3572] = layer2_outputs[3624];
    assign layer3_outputs[3573] = ~((layer2_outputs[1731]) & (layer2_outputs[3279]));
    assign layer3_outputs[3574] = ~((layer2_outputs[249]) | (layer2_outputs[425]));
    assign layer3_outputs[3575] = ~((layer2_outputs[2520]) | (layer2_outputs[4055]));
    assign layer3_outputs[3576] = layer2_outputs[4511];
    assign layer3_outputs[3577] = 1'b1;
    assign layer3_outputs[3578] = (layer2_outputs[487]) | (layer2_outputs[2528]);
    assign layer3_outputs[3579] = ~(layer2_outputs[4627]);
    assign layer3_outputs[3580] = ~(layer2_outputs[3524]);
    assign layer3_outputs[3581] = layer2_outputs[2151];
    assign layer3_outputs[3582] = 1'b0;
    assign layer3_outputs[3583] = (layer2_outputs[649]) & (layer2_outputs[4720]);
    assign layer3_outputs[3584] = (layer2_outputs[1361]) & (layer2_outputs[4681]);
    assign layer3_outputs[3585] = 1'b1;
    assign layer3_outputs[3586] = (layer2_outputs[1422]) & ~(layer2_outputs[4590]);
    assign layer3_outputs[3587] = ~(layer2_outputs[3542]) | (layer2_outputs[726]);
    assign layer3_outputs[3588] = ~(layer2_outputs[750]);
    assign layer3_outputs[3589] = (layer2_outputs[4490]) & (layer2_outputs[4763]);
    assign layer3_outputs[3590] = (layer2_outputs[2603]) & (layer2_outputs[378]);
    assign layer3_outputs[3591] = layer2_outputs[5048];
    assign layer3_outputs[3592] = ~(layer2_outputs[4184]);
    assign layer3_outputs[3593] = 1'b0;
    assign layer3_outputs[3594] = layer2_outputs[4186];
    assign layer3_outputs[3595] = ~(layer2_outputs[2789]);
    assign layer3_outputs[3596] = ~((layer2_outputs[609]) | (layer2_outputs[461]));
    assign layer3_outputs[3597] = (layer2_outputs[1343]) & (layer2_outputs[3231]);
    assign layer3_outputs[3598] = ~((layer2_outputs[2451]) | (layer2_outputs[4093]));
    assign layer3_outputs[3599] = (layer2_outputs[3752]) & (layer2_outputs[2290]);
    assign layer3_outputs[3600] = ~(layer2_outputs[3971]);
    assign layer3_outputs[3601] = ~(layer2_outputs[666]);
    assign layer3_outputs[3602] = 1'b0;
    assign layer3_outputs[3603] = (layer2_outputs[1120]) ^ (layer2_outputs[4256]);
    assign layer3_outputs[3604] = (layer2_outputs[1877]) & (layer2_outputs[2646]);
    assign layer3_outputs[3605] = layer2_outputs[2856];
    assign layer3_outputs[3606] = ~(layer2_outputs[801]) | (layer2_outputs[2530]);
    assign layer3_outputs[3607] = layer2_outputs[46];
    assign layer3_outputs[3608] = ~(layer2_outputs[107]);
    assign layer3_outputs[3609] = (layer2_outputs[5053]) & ~(layer2_outputs[2984]);
    assign layer3_outputs[3610] = ~(layer2_outputs[3312]) | (layer2_outputs[1373]);
    assign layer3_outputs[3611] = ~(layer2_outputs[5112]) | (layer2_outputs[3224]);
    assign layer3_outputs[3612] = layer2_outputs[3806];
    assign layer3_outputs[3613] = ~(layer2_outputs[548]) | (layer2_outputs[816]);
    assign layer3_outputs[3614] = ~(layer2_outputs[41]);
    assign layer3_outputs[3615] = ~(layer2_outputs[2026]) | (layer2_outputs[2954]);
    assign layer3_outputs[3616] = (layer2_outputs[4561]) & (layer2_outputs[2394]);
    assign layer3_outputs[3617] = (layer2_outputs[1194]) & (layer2_outputs[1679]);
    assign layer3_outputs[3618] = ~(layer2_outputs[1621]);
    assign layer3_outputs[3619] = ~((layer2_outputs[2790]) | (layer2_outputs[2750]));
    assign layer3_outputs[3620] = layer2_outputs[2374];
    assign layer3_outputs[3621] = ~(layer2_outputs[2940]) | (layer2_outputs[99]);
    assign layer3_outputs[3622] = ~(layer2_outputs[3415]);
    assign layer3_outputs[3623] = layer2_outputs[76];
    assign layer3_outputs[3624] = layer2_outputs[3237];
    assign layer3_outputs[3625] = 1'b1;
    assign layer3_outputs[3626] = 1'b1;
    assign layer3_outputs[3627] = (layer2_outputs[4538]) & ~(layer2_outputs[1695]);
    assign layer3_outputs[3628] = ~(layer2_outputs[1320]) | (layer2_outputs[4349]);
    assign layer3_outputs[3629] = layer2_outputs[755];
    assign layer3_outputs[3630] = ~(layer2_outputs[3239]) | (layer2_outputs[798]);
    assign layer3_outputs[3631] = 1'b0;
    assign layer3_outputs[3632] = ~(layer2_outputs[3938]);
    assign layer3_outputs[3633] = ~(layer2_outputs[3411]) | (layer2_outputs[135]);
    assign layer3_outputs[3634] = ~(layer2_outputs[4530]);
    assign layer3_outputs[3635] = ~(layer2_outputs[2566]);
    assign layer3_outputs[3636] = ~(layer2_outputs[3975]) | (layer2_outputs[595]);
    assign layer3_outputs[3637] = layer2_outputs[1573];
    assign layer3_outputs[3638] = 1'b1;
    assign layer3_outputs[3639] = (layer2_outputs[138]) & ~(layer2_outputs[2036]);
    assign layer3_outputs[3640] = ~(layer2_outputs[4202]) | (layer2_outputs[4894]);
    assign layer3_outputs[3641] = (layer2_outputs[4806]) & ~(layer2_outputs[4442]);
    assign layer3_outputs[3642] = 1'b0;
    assign layer3_outputs[3643] = layer2_outputs[3517];
    assign layer3_outputs[3644] = ~((layer2_outputs[946]) & (layer2_outputs[1090]));
    assign layer3_outputs[3645] = ~((layer2_outputs[310]) ^ (layer2_outputs[2967]));
    assign layer3_outputs[3646] = (layer2_outputs[2168]) | (layer2_outputs[1366]);
    assign layer3_outputs[3647] = (layer2_outputs[3267]) & ~(layer2_outputs[962]);
    assign layer3_outputs[3648] = layer2_outputs[2306];
    assign layer3_outputs[3649] = ~((layer2_outputs[972]) & (layer2_outputs[3639]));
    assign layer3_outputs[3650] = ~(layer2_outputs[1891]);
    assign layer3_outputs[3651] = ~(layer2_outputs[1265]);
    assign layer3_outputs[3652] = 1'b0;
    assign layer3_outputs[3653] = ~(layer2_outputs[484]);
    assign layer3_outputs[3654] = ~((layer2_outputs[148]) ^ (layer2_outputs[3463]));
    assign layer3_outputs[3655] = ~(layer2_outputs[4579]);
    assign layer3_outputs[3656] = 1'b0;
    assign layer3_outputs[3657] = (layer2_outputs[4507]) ^ (layer2_outputs[2847]);
    assign layer3_outputs[3658] = layer2_outputs[1168];
    assign layer3_outputs[3659] = layer2_outputs[776];
    assign layer3_outputs[3660] = (layer2_outputs[1558]) ^ (layer2_outputs[1444]);
    assign layer3_outputs[3661] = ~(layer2_outputs[654]);
    assign layer3_outputs[3662] = ~((layer2_outputs[3454]) & (layer2_outputs[2392]));
    assign layer3_outputs[3663] = ~((layer2_outputs[1170]) | (layer2_outputs[4094]));
    assign layer3_outputs[3664] = 1'b0;
    assign layer3_outputs[3665] = ~(layer2_outputs[1956]);
    assign layer3_outputs[3666] = ~((layer2_outputs[1862]) | (layer2_outputs[4781]));
    assign layer3_outputs[3667] = ~((layer2_outputs[2126]) & (layer2_outputs[4296]));
    assign layer3_outputs[3668] = (layer2_outputs[4279]) & (layer2_outputs[4164]);
    assign layer3_outputs[3669] = 1'b0;
    assign layer3_outputs[3670] = (layer2_outputs[1501]) & ~(layer2_outputs[832]);
    assign layer3_outputs[3671] = ~((layer2_outputs[116]) | (layer2_outputs[2298]));
    assign layer3_outputs[3672] = (layer2_outputs[1357]) | (layer2_outputs[55]);
    assign layer3_outputs[3673] = layer2_outputs[1537];
    assign layer3_outputs[3674] = ~((layer2_outputs[1553]) & (layer2_outputs[2916]));
    assign layer3_outputs[3675] = (layer2_outputs[4730]) | (layer2_outputs[3809]);
    assign layer3_outputs[3676] = ~(layer2_outputs[968]);
    assign layer3_outputs[3677] = ~((layer2_outputs[992]) & (layer2_outputs[165]));
    assign layer3_outputs[3678] = layer2_outputs[4021];
    assign layer3_outputs[3679] = (layer2_outputs[4665]) | (layer2_outputs[656]);
    assign layer3_outputs[3680] = ~(layer2_outputs[2004]) | (layer2_outputs[3860]);
    assign layer3_outputs[3681] = layer2_outputs[4524];
    assign layer3_outputs[3682] = (layer2_outputs[2570]) & ~(layer2_outputs[718]);
    assign layer3_outputs[3683] = ~((layer2_outputs[1485]) | (layer2_outputs[4409]));
    assign layer3_outputs[3684] = (layer2_outputs[5118]) & ~(layer2_outputs[1690]);
    assign layer3_outputs[3685] = layer2_outputs[2160];
    assign layer3_outputs[3686] = ~((layer2_outputs[3174]) & (layer2_outputs[2932]));
    assign layer3_outputs[3687] = 1'b1;
    assign layer3_outputs[3688] = layer2_outputs[886];
    assign layer3_outputs[3689] = ~((layer2_outputs[4464]) & (layer2_outputs[1007]));
    assign layer3_outputs[3690] = ~(layer2_outputs[465]);
    assign layer3_outputs[3691] = (layer2_outputs[3370]) | (layer2_outputs[2062]);
    assign layer3_outputs[3692] = ~(layer2_outputs[3541]);
    assign layer3_outputs[3693] = 1'b0;
    assign layer3_outputs[3694] = ~(layer2_outputs[1972]);
    assign layer3_outputs[3695] = ~((layer2_outputs[1822]) | (layer2_outputs[4960]));
    assign layer3_outputs[3696] = ~(layer2_outputs[1998]) | (layer2_outputs[3187]);
    assign layer3_outputs[3697] = layer2_outputs[2855];
    assign layer3_outputs[3698] = ~(layer2_outputs[5030]);
    assign layer3_outputs[3699] = (layer2_outputs[2101]) & ~(layer2_outputs[1421]);
    assign layer3_outputs[3700] = layer2_outputs[920];
    assign layer3_outputs[3701] = (layer2_outputs[84]) & ~(layer2_outputs[1874]);
    assign layer3_outputs[3702] = layer2_outputs[913];
    assign layer3_outputs[3703] = ~(layer2_outputs[1994]);
    assign layer3_outputs[3704] = ~((layer2_outputs[3097]) & (layer2_outputs[3216]));
    assign layer3_outputs[3705] = (layer2_outputs[2659]) & ~(layer2_outputs[684]);
    assign layer3_outputs[3706] = (layer2_outputs[2934]) ^ (layer2_outputs[2324]);
    assign layer3_outputs[3707] = ~((layer2_outputs[1889]) & (layer2_outputs[1532]));
    assign layer3_outputs[3708] = 1'b1;
    assign layer3_outputs[3709] = ~(layer2_outputs[3011]) | (layer2_outputs[4093]);
    assign layer3_outputs[3710] = ~(layer2_outputs[4360]);
    assign layer3_outputs[3711] = (layer2_outputs[5044]) & (layer2_outputs[3062]);
    assign layer3_outputs[3712] = layer2_outputs[2439];
    assign layer3_outputs[3713] = ~(layer2_outputs[1514]);
    assign layer3_outputs[3714] = layer2_outputs[4969];
    assign layer3_outputs[3715] = layer2_outputs[5045];
    assign layer3_outputs[3716] = (layer2_outputs[4578]) | (layer2_outputs[4099]);
    assign layer3_outputs[3717] = ~((layer2_outputs[4660]) ^ (layer2_outputs[1283]));
    assign layer3_outputs[3718] = ~(layer2_outputs[1661]) | (layer2_outputs[2019]);
    assign layer3_outputs[3719] = ~((layer2_outputs[1839]) | (layer2_outputs[3597]));
    assign layer3_outputs[3720] = ~(layer2_outputs[2885]) | (layer2_outputs[2874]);
    assign layer3_outputs[3721] = (layer2_outputs[4933]) & ~(layer2_outputs[2058]);
    assign layer3_outputs[3722] = ~(layer2_outputs[211]) | (layer2_outputs[2761]);
    assign layer3_outputs[3723] = ~(layer2_outputs[1073]);
    assign layer3_outputs[3724] = ~(layer2_outputs[2183]) | (layer2_outputs[2137]);
    assign layer3_outputs[3725] = (layer2_outputs[838]) & ~(layer2_outputs[753]);
    assign layer3_outputs[3726] = ~((layer2_outputs[2859]) | (layer2_outputs[140]));
    assign layer3_outputs[3727] = ~(layer2_outputs[457]) | (layer2_outputs[2189]);
    assign layer3_outputs[3728] = ~(layer2_outputs[5037]);
    assign layer3_outputs[3729] = ~(layer2_outputs[277]);
    assign layer3_outputs[3730] = ~(layer2_outputs[1809]);
    assign layer3_outputs[3731] = ~(layer2_outputs[3578]);
    assign layer3_outputs[3732] = layer2_outputs[1547];
    assign layer3_outputs[3733] = ~(layer2_outputs[492]);
    assign layer3_outputs[3734] = ~(layer2_outputs[1386]) | (layer2_outputs[4732]);
    assign layer3_outputs[3735] = layer2_outputs[1225];
    assign layer3_outputs[3736] = (layer2_outputs[4828]) & ~(layer2_outputs[1888]);
    assign layer3_outputs[3737] = (layer2_outputs[1772]) & (layer2_outputs[2837]);
    assign layer3_outputs[3738] = (layer2_outputs[1757]) & (layer2_outputs[4707]);
    assign layer3_outputs[3739] = 1'b1;
    assign layer3_outputs[3740] = (layer2_outputs[2274]) & ~(layer2_outputs[906]);
    assign layer3_outputs[3741] = ~((layer2_outputs[2478]) | (layer2_outputs[3802]));
    assign layer3_outputs[3742] = (layer2_outputs[121]) & ~(layer2_outputs[3474]);
    assign layer3_outputs[3743] = ~((layer2_outputs[2238]) | (layer2_outputs[4076]));
    assign layer3_outputs[3744] = (layer2_outputs[3323]) & ~(layer2_outputs[3052]);
    assign layer3_outputs[3745] = ~(layer2_outputs[291]);
    assign layer3_outputs[3746] = ~(layer2_outputs[1052]) | (layer2_outputs[3857]);
    assign layer3_outputs[3747] = 1'b1;
    assign layer3_outputs[3748] = ~((layer2_outputs[3619]) | (layer2_outputs[2089]));
    assign layer3_outputs[3749] = (layer2_outputs[2941]) | (layer2_outputs[4745]);
    assign layer3_outputs[3750] = layer2_outputs[1415];
    assign layer3_outputs[3751] = ~(layer2_outputs[889]) | (layer2_outputs[80]);
    assign layer3_outputs[3752] = (layer2_outputs[773]) & (layer2_outputs[4232]);
    assign layer3_outputs[3753] = ~(layer2_outputs[2313]);
    assign layer3_outputs[3754] = layer2_outputs[4151];
    assign layer3_outputs[3755] = ~(layer2_outputs[1604]);
    assign layer3_outputs[3756] = ~(layer2_outputs[4477]) | (layer2_outputs[1726]);
    assign layer3_outputs[3757] = ~(layer2_outputs[4335]) | (layer2_outputs[2594]);
    assign layer3_outputs[3758] = ~((layer2_outputs[1595]) ^ (layer2_outputs[2055]));
    assign layer3_outputs[3759] = ~(layer2_outputs[888]) | (layer2_outputs[3956]);
    assign layer3_outputs[3760] = ~(layer2_outputs[1440]) | (layer2_outputs[1205]);
    assign layer3_outputs[3761] = (layer2_outputs[1777]) ^ (layer2_outputs[3757]);
    assign layer3_outputs[3762] = 1'b1;
    assign layer3_outputs[3763] = ~(layer2_outputs[3313]);
    assign layer3_outputs[3764] = (layer2_outputs[2087]) & (layer2_outputs[1728]);
    assign layer3_outputs[3765] = ~(layer2_outputs[3438]);
    assign layer3_outputs[3766] = (layer2_outputs[416]) & (layer2_outputs[2580]);
    assign layer3_outputs[3767] = ~(layer2_outputs[4276]);
    assign layer3_outputs[3768] = 1'b1;
    assign layer3_outputs[3769] = 1'b0;
    assign layer3_outputs[3770] = (layer2_outputs[2151]) & ~(layer2_outputs[2280]);
    assign layer3_outputs[3771] = ~((layer2_outputs[3969]) & (layer2_outputs[3768]));
    assign layer3_outputs[3772] = ~(layer2_outputs[1564]) | (layer2_outputs[527]);
    assign layer3_outputs[3773] = 1'b1;
    assign layer3_outputs[3774] = 1'b0;
    assign layer3_outputs[3775] = ~(layer2_outputs[5046]);
    assign layer3_outputs[3776] = 1'b1;
    assign layer3_outputs[3777] = layer2_outputs[4000];
    assign layer3_outputs[3778] = (layer2_outputs[4150]) & (layer2_outputs[2379]);
    assign layer3_outputs[3779] = (layer2_outputs[4483]) & ~(layer2_outputs[1541]);
    assign layer3_outputs[3780] = (layer2_outputs[590]) & ~(layer2_outputs[4401]);
    assign layer3_outputs[3781] = layer2_outputs[2257];
    assign layer3_outputs[3782] = ~((layer2_outputs[4933]) ^ (layer2_outputs[209]));
    assign layer3_outputs[3783] = ~((layer2_outputs[65]) | (layer2_outputs[885]));
    assign layer3_outputs[3784] = 1'b1;
    assign layer3_outputs[3785] = (layer2_outputs[4457]) & ~(layer2_outputs[1921]);
    assign layer3_outputs[3786] = ~(layer2_outputs[1514]) | (layer2_outputs[704]);
    assign layer3_outputs[3787] = (layer2_outputs[3302]) | (layer2_outputs[4022]);
    assign layer3_outputs[3788] = layer2_outputs[3688];
    assign layer3_outputs[3789] = ~((layer2_outputs[3375]) | (layer2_outputs[4374]));
    assign layer3_outputs[3790] = ~(layer2_outputs[1134]) | (layer2_outputs[1708]);
    assign layer3_outputs[3791] = layer2_outputs[2407];
    assign layer3_outputs[3792] = ~(layer2_outputs[2490]);
    assign layer3_outputs[3793] = ~((layer2_outputs[324]) & (layer2_outputs[4953]));
    assign layer3_outputs[3794] = 1'b1;
    assign layer3_outputs[3795] = ~((layer2_outputs[2198]) ^ (layer2_outputs[2365]));
    assign layer3_outputs[3796] = layer2_outputs[326];
    assign layer3_outputs[3797] = ~((layer2_outputs[2906]) | (layer2_outputs[3388]));
    assign layer3_outputs[3798] = layer2_outputs[3949];
    assign layer3_outputs[3799] = (layer2_outputs[3273]) | (layer2_outputs[1540]);
    assign layer3_outputs[3800] = ~(layer2_outputs[3294]) | (layer2_outputs[3922]);
    assign layer3_outputs[3801] = ~(layer2_outputs[2594]);
    assign layer3_outputs[3802] = ~((layer2_outputs[4589]) & (layer2_outputs[681]));
    assign layer3_outputs[3803] = 1'b0;
    assign layer3_outputs[3804] = layer2_outputs[3215];
    assign layer3_outputs[3805] = 1'b1;
    assign layer3_outputs[3806] = 1'b0;
    assign layer3_outputs[3807] = ~(layer2_outputs[219]) | (layer2_outputs[3376]);
    assign layer3_outputs[3808] = ~((layer2_outputs[4087]) | (layer2_outputs[139]));
    assign layer3_outputs[3809] = (layer2_outputs[122]) & (layer2_outputs[5056]);
    assign layer3_outputs[3810] = layer2_outputs[57];
    assign layer3_outputs[3811] = ~(layer2_outputs[1879]);
    assign layer3_outputs[3812] = 1'b0;
    assign layer3_outputs[3813] = 1'b1;
    assign layer3_outputs[3814] = ~(layer2_outputs[2192]);
    assign layer3_outputs[3815] = (layer2_outputs[4461]) & ~(layer2_outputs[2061]);
    assign layer3_outputs[3816] = 1'b0;
    assign layer3_outputs[3817] = layer2_outputs[1881];
    assign layer3_outputs[3818] = layer2_outputs[1239];
    assign layer3_outputs[3819] = layer2_outputs[3044];
    assign layer3_outputs[3820] = ~((layer2_outputs[3918]) | (layer2_outputs[2160]));
    assign layer3_outputs[3821] = ~((layer2_outputs[544]) & (layer2_outputs[201]));
    assign layer3_outputs[3822] = layer2_outputs[4643];
    assign layer3_outputs[3823] = layer2_outputs[2686];
    assign layer3_outputs[3824] = 1'b1;
    assign layer3_outputs[3825] = ~(layer2_outputs[4530]);
    assign layer3_outputs[3826] = ~(layer2_outputs[3574]);
    assign layer3_outputs[3827] = (layer2_outputs[1409]) & ~(layer2_outputs[4211]);
    assign layer3_outputs[3828] = (layer2_outputs[585]) | (layer2_outputs[549]);
    assign layer3_outputs[3829] = 1'b0;
    assign layer3_outputs[3830] = ~(layer2_outputs[2939]);
    assign layer3_outputs[3831] = (layer2_outputs[3315]) ^ (layer2_outputs[780]);
    assign layer3_outputs[3832] = (layer2_outputs[3023]) & ~(layer2_outputs[2300]);
    assign layer3_outputs[3833] = ~(layer2_outputs[5014]);
    assign layer3_outputs[3834] = layer2_outputs[2115];
    assign layer3_outputs[3835] = layer2_outputs[2344];
    assign layer3_outputs[3836] = (layer2_outputs[1324]) & ~(layer2_outputs[1869]);
    assign layer3_outputs[3837] = 1'b0;
    assign layer3_outputs[3838] = layer2_outputs[892];
    assign layer3_outputs[3839] = ~((layer2_outputs[1185]) | (layer2_outputs[2472]));
    assign layer3_outputs[3840] = ~((layer2_outputs[1178]) & (layer2_outputs[1311]));
    assign layer3_outputs[3841] = layer2_outputs[3758];
    assign layer3_outputs[3842] = layer2_outputs[3894];
    assign layer3_outputs[3843] = 1'b1;
    assign layer3_outputs[3844] = layer2_outputs[979];
    assign layer3_outputs[3845] = ~(layer2_outputs[2663]) | (layer2_outputs[4714]);
    assign layer3_outputs[3846] = ~(layer2_outputs[1345]);
    assign layer3_outputs[3847] = ~((layer2_outputs[2353]) | (layer2_outputs[3188]));
    assign layer3_outputs[3848] = 1'b1;
    assign layer3_outputs[3849] = (layer2_outputs[1991]) & ~(layer2_outputs[4205]);
    assign layer3_outputs[3850] = layer2_outputs[1604];
    assign layer3_outputs[3851] = layer2_outputs[4145];
    assign layer3_outputs[3852] = (layer2_outputs[3645]) ^ (layer2_outputs[2828]);
    assign layer3_outputs[3853] = ~((layer2_outputs[4466]) & (layer2_outputs[4599]));
    assign layer3_outputs[3854] = (layer2_outputs[4596]) | (layer2_outputs[4202]);
    assign layer3_outputs[3855] = 1'b0;
    assign layer3_outputs[3856] = ~(layer2_outputs[76]);
    assign layer3_outputs[3857] = ~(layer2_outputs[2251]) | (layer2_outputs[3179]);
    assign layer3_outputs[3858] = 1'b0;
    assign layer3_outputs[3859] = ~(layer2_outputs[4928]);
    assign layer3_outputs[3860] = ~(layer2_outputs[793]) | (layer2_outputs[299]);
    assign layer3_outputs[3861] = layer2_outputs[4130];
    assign layer3_outputs[3862] = (layer2_outputs[1376]) & ~(layer2_outputs[3360]);
    assign layer3_outputs[3863] = ~(layer2_outputs[4764]);
    assign layer3_outputs[3864] = ~(layer2_outputs[868]);
    assign layer3_outputs[3865] = layer2_outputs[3072];
    assign layer3_outputs[3866] = ~(layer2_outputs[420]);
    assign layer3_outputs[3867] = ~((layer2_outputs[2523]) & (layer2_outputs[3205]));
    assign layer3_outputs[3868] = 1'b0;
    assign layer3_outputs[3869] = ~(layer2_outputs[85]) | (layer2_outputs[2206]);
    assign layer3_outputs[3870] = 1'b0;
    assign layer3_outputs[3871] = (layer2_outputs[2575]) | (layer2_outputs[1305]);
    assign layer3_outputs[3872] = ~((layer2_outputs[2437]) | (layer2_outputs[3697]));
    assign layer3_outputs[3873] = (layer2_outputs[2642]) & (layer2_outputs[1180]);
    assign layer3_outputs[3874] = (layer2_outputs[3041]) | (layer2_outputs[2145]);
    assign layer3_outputs[3875] = (layer2_outputs[2023]) & ~(layer2_outputs[2225]);
    assign layer3_outputs[3876] = (layer2_outputs[3035]) & (layer2_outputs[4311]);
    assign layer3_outputs[3877] = (layer2_outputs[1683]) & ~(layer2_outputs[346]);
    assign layer3_outputs[3878] = ~(layer2_outputs[266]);
    assign layer3_outputs[3879] = (layer2_outputs[11]) & ~(layer2_outputs[1271]);
    assign layer3_outputs[3880] = ~(layer2_outputs[3545]) | (layer2_outputs[3004]);
    assign layer3_outputs[3881] = ~(layer2_outputs[284]);
    assign layer3_outputs[3882] = (layer2_outputs[2104]) & (layer2_outputs[2732]);
    assign layer3_outputs[3883] = ~((layer2_outputs[3919]) ^ (layer2_outputs[1454]));
    assign layer3_outputs[3884] = ~(layer2_outputs[2756]);
    assign layer3_outputs[3885] = ~((layer2_outputs[1053]) | (layer2_outputs[2009]));
    assign layer3_outputs[3886] = (layer2_outputs[2317]) & (layer2_outputs[312]);
    assign layer3_outputs[3887] = (layer2_outputs[826]) & ~(layer2_outputs[1055]);
    assign layer3_outputs[3888] = ~(layer2_outputs[2833]) | (layer2_outputs[1505]);
    assign layer3_outputs[3889] = ~(layer2_outputs[3378]);
    assign layer3_outputs[3890] = (layer2_outputs[228]) & (layer2_outputs[1291]);
    assign layer3_outputs[3891] = layer2_outputs[3771];
    assign layer3_outputs[3892] = layer2_outputs[2066];
    assign layer3_outputs[3893] = layer2_outputs[4655];
    assign layer3_outputs[3894] = layer2_outputs[778];
    assign layer3_outputs[3895] = layer2_outputs[435];
    assign layer3_outputs[3896] = (layer2_outputs[1494]) | (layer2_outputs[653]);
    assign layer3_outputs[3897] = ~((layer2_outputs[1834]) & (layer2_outputs[4790]));
    assign layer3_outputs[3898] = layer2_outputs[4868];
    assign layer3_outputs[3899] = layer2_outputs[2266];
    assign layer3_outputs[3900] = ~(layer2_outputs[4392]);
    assign layer3_outputs[3901] = ~(layer2_outputs[5083]);
    assign layer3_outputs[3902] = ~((layer2_outputs[5050]) & (layer2_outputs[3979]));
    assign layer3_outputs[3903] = ~(layer2_outputs[637]);
    assign layer3_outputs[3904] = layer2_outputs[456];
    assign layer3_outputs[3905] = ~((layer2_outputs[2244]) & (layer2_outputs[994]));
    assign layer3_outputs[3906] = ~(layer2_outputs[3347]) | (layer2_outputs[4116]);
    assign layer3_outputs[3907] = (layer2_outputs[1759]) & ~(layer2_outputs[4525]);
    assign layer3_outputs[3908] = (layer2_outputs[3185]) & (layer2_outputs[3983]);
    assign layer3_outputs[3909] = (layer2_outputs[7]) & ~(layer2_outputs[4902]);
    assign layer3_outputs[3910] = (layer2_outputs[3454]) | (layer2_outputs[2724]);
    assign layer3_outputs[3911] = ~((layer2_outputs[2403]) ^ (layer2_outputs[2296]));
    assign layer3_outputs[3912] = (layer2_outputs[2645]) & ~(layer2_outputs[3256]);
    assign layer3_outputs[3913] = ~(layer2_outputs[457]);
    assign layer3_outputs[3914] = ~(layer2_outputs[3537]);
    assign layer3_outputs[3915] = 1'b0;
    assign layer3_outputs[3916] = layer2_outputs[392];
    assign layer3_outputs[3917] = (layer2_outputs[2768]) & ~(layer2_outputs[3854]);
    assign layer3_outputs[3918] = 1'b0;
    assign layer3_outputs[3919] = ~(layer2_outputs[2538]) | (layer2_outputs[136]);
    assign layer3_outputs[3920] = ~(layer2_outputs[4350]) | (layer2_outputs[3485]);
    assign layer3_outputs[3921] = ~(layer2_outputs[3230]) | (layer2_outputs[1098]);
    assign layer3_outputs[3922] = ~((layer2_outputs[4421]) & (layer2_outputs[4506]));
    assign layer3_outputs[3923] = layer2_outputs[53];
    assign layer3_outputs[3924] = ~((layer2_outputs[4532]) | (layer2_outputs[2176]));
    assign layer3_outputs[3925] = (layer2_outputs[263]) & (layer2_outputs[70]);
    assign layer3_outputs[3926] = (layer2_outputs[4240]) | (layer2_outputs[1041]);
    assign layer3_outputs[3927] = 1'b0;
    assign layer3_outputs[3928] = layer2_outputs[2102];
    assign layer3_outputs[3929] = (layer2_outputs[2516]) & ~(layer2_outputs[3409]);
    assign layer3_outputs[3930] = (layer2_outputs[4936]) & ~(layer2_outputs[1312]);
    assign layer3_outputs[3931] = (layer2_outputs[3929]) & (layer2_outputs[1125]);
    assign layer3_outputs[3932] = layer2_outputs[182];
    assign layer3_outputs[3933] = layer2_outputs[2115];
    assign layer3_outputs[3934] = 1'b1;
    assign layer3_outputs[3935] = ~((layer2_outputs[4766]) & (layer2_outputs[3736]));
    assign layer3_outputs[3936] = (layer2_outputs[1363]) | (layer2_outputs[1443]);
    assign layer3_outputs[3937] = ~(layer2_outputs[1284]) | (layer2_outputs[769]);
    assign layer3_outputs[3938] = ~(layer2_outputs[887]);
    assign layer3_outputs[3939] = ~((layer2_outputs[3272]) ^ (layer2_outputs[4344]));
    assign layer3_outputs[3940] = (layer2_outputs[1462]) | (layer2_outputs[3959]);
    assign layer3_outputs[3941] = ~(layer2_outputs[4634]);
    assign layer3_outputs[3942] = (layer2_outputs[1634]) & ~(layer2_outputs[285]);
    assign layer3_outputs[3943] = 1'b0;
    assign layer3_outputs[3944] = ~(layer2_outputs[3460]);
    assign layer3_outputs[3945] = layer2_outputs[3866];
    assign layer3_outputs[3946] = ~(layer2_outputs[3493]) | (layer2_outputs[4829]);
    assign layer3_outputs[3947] = ~((layer2_outputs[4546]) | (layer2_outputs[1665]));
    assign layer3_outputs[3948] = ~(layer2_outputs[4638]) | (layer2_outputs[1011]);
    assign layer3_outputs[3949] = ~(layer2_outputs[3827]);
    assign layer3_outputs[3950] = 1'b1;
    assign layer3_outputs[3951] = (layer2_outputs[1785]) & ~(layer2_outputs[4501]);
    assign layer3_outputs[3952] = ~(layer2_outputs[4134]);
    assign layer3_outputs[3953] = ~(layer2_outputs[2352]) | (layer2_outputs[4527]);
    assign layer3_outputs[3954] = (layer2_outputs[4750]) & ~(layer2_outputs[1413]);
    assign layer3_outputs[3955] = ~(layer2_outputs[892]) | (layer2_outputs[2276]);
    assign layer3_outputs[3956] = ~(layer2_outputs[3860]);
    assign layer3_outputs[3957] = ~(layer2_outputs[4514]);
    assign layer3_outputs[3958] = (layer2_outputs[4175]) & (layer2_outputs[3263]);
    assign layer3_outputs[3959] = (layer2_outputs[4494]) & ~(layer2_outputs[1601]);
    assign layer3_outputs[3960] = ~((layer2_outputs[4114]) | (layer2_outputs[5099]));
    assign layer3_outputs[3961] = 1'b0;
    assign layer3_outputs[3962] = layer2_outputs[4837];
    assign layer3_outputs[3963] = 1'b1;
    assign layer3_outputs[3964] = ~(layer2_outputs[4163]) | (layer2_outputs[3090]);
    assign layer3_outputs[3965] = (layer2_outputs[2680]) | (layer2_outputs[3117]);
    assign layer3_outputs[3966] = ~(layer2_outputs[2742]);
    assign layer3_outputs[3967] = ~(layer2_outputs[2654]);
    assign layer3_outputs[3968] = 1'b1;
    assign layer3_outputs[3969] = ~((layer2_outputs[2854]) ^ (layer2_outputs[508]));
    assign layer3_outputs[3970] = ~(layer2_outputs[252]);
    assign layer3_outputs[3971] = ~(layer2_outputs[2152]) | (layer2_outputs[1017]);
    assign layer3_outputs[3972] = ~(layer2_outputs[5020]) | (layer2_outputs[2569]);
    assign layer3_outputs[3973] = (layer2_outputs[3659]) & (layer2_outputs[4679]);
    assign layer3_outputs[3974] = (layer2_outputs[4764]) & ~(layer2_outputs[4080]);
    assign layer3_outputs[3975] = (layer2_outputs[1778]) & (layer2_outputs[3875]);
    assign layer3_outputs[3976] = ~(layer2_outputs[4029]) | (layer2_outputs[1938]);
    assign layer3_outputs[3977] = layer2_outputs[1268];
    assign layer3_outputs[3978] = layer2_outputs[4345];
    assign layer3_outputs[3979] = layer2_outputs[2114];
    assign layer3_outputs[3980] = ~(layer2_outputs[3091]) | (layer2_outputs[3508]);
    assign layer3_outputs[3981] = (layer2_outputs[2078]) & ~(layer2_outputs[4522]);
    assign layer3_outputs[3982] = ~(layer2_outputs[3254]) | (layer2_outputs[3087]);
    assign layer3_outputs[3983] = (layer2_outputs[4705]) & ~(layer2_outputs[4880]);
    assign layer3_outputs[3984] = ~(layer2_outputs[3717]);
    assign layer3_outputs[3985] = (layer2_outputs[3867]) & ~(layer2_outputs[3253]);
    assign layer3_outputs[3986] = 1'b1;
    assign layer3_outputs[3987] = (layer2_outputs[151]) | (layer2_outputs[2220]);
    assign layer3_outputs[3988] = 1'b0;
    assign layer3_outputs[3989] = ~(layer2_outputs[4998]) | (layer2_outputs[2825]);
    assign layer3_outputs[3990] = 1'b1;
    assign layer3_outputs[3991] = ~(layer2_outputs[33]);
    assign layer3_outputs[3992] = (layer2_outputs[3788]) & ~(layer2_outputs[587]);
    assign layer3_outputs[3993] = ~(layer2_outputs[4133]);
    assign layer3_outputs[3994] = (layer2_outputs[1512]) & ~(layer2_outputs[2159]);
    assign layer3_outputs[3995] = 1'b0;
    assign layer3_outputs[3996] = ~(layer2_outputs[4600]);
    assign layer3_outputs[3997] = (layer2_outputs[2281]) & (layer2_outputs[2707]);
    assign layer3_outputs[3998] = ~(layer2_outputs[3757]);
    assign layer3_outputs[3999] = (layer2_outputs[4862]) & ~(layer2_outputs[2474]);
    assign layer3_outputs[4000] = ~(layer2_outputs[1135]) | (layer2_outputs[5091]);
    assign layer3_outputs[4001] = (layer2_outputs[957]) | (layer2_outputs[1935]);
    assign layer3_outputs[4002] = (layer2_outputs[723]) & ~(layer2_outputs[1154]);
    assign layer3_outputs[4003] = ~((layer2_outputs[2964]) | (layer2_outputs[3150]));
    assign layer3_outputs[4004] = (layer2_outputs[3017]) & ~(layer2_outputs[4073]);
    assign layer3_outputs[4005] = layer2_outputs[4807];
    assign layer3_outputs[4006] = 1'b0;
    assign layer3_outputs[4007] = layer2_outputs[1100];
    assign layer3_outputs[4008] = 1'b0;
    assign layer3_outputs[4009] = (layer2_outputs[3147]) | (layer2_outputs[313]);
    assign layer3_outputs[4010] = (layer2_outputs[237]) & ~(layer2_outputs[4680]);
    assign layer3_outputs[4011] = ~(layer2_outputs[900]);
    assign layer3_outputs[4012] = (layer2_outputs[911]) & ~(layer2_outputs[3529]);
    assign layer3_outputs[4013] = (layer2_outputs[4981]) | (layer2_outputs[3800]);
    assign layer3_outputs[4014] = layer2_outputs[3784];
    assign layer3_outputs[4015] = layer2_outputs[4695];
    assign layer3_outputs[4016] = ~((layer2_outputs[3580]) | (layer2_outputs[1396]));
    assign layer3_outputs[4017] = ~(layer2_outputs[917]) | (layer2_outputs[5117]);
    assign layer3_outputs[4018] = (layer2_outputs[4669]) & ~(layer2_outputs[4613]);
    assign layer3_outputs[4019] = (layer2_outputs[2772]) | (layer2_outputs[585]);
    assign layer3_outputs[4020] = 1'b0;
    assign layer3_outputs[4021] = (layer2_outputs[1774]) & (layer2_outputs[2072]);
    assign layer3_outputs[4022] = ~(layer2_outputs[3428]) | (layer2_outputs[1203]);
    assign layer3_outputs[4023] = ~(layer2_outputs[949]);
    assign layer3_outputs[4024] = ~(layer2_outputs[3693]) | (layer2_outputs[183]);
    assign layer3_outputs[4025] = ~(layer2_outputs[1155]);
    assign layer3_outputs[4026] = ~(layer2_outputs[1281]);
    assign layer3_outputs[4027] = ~((layer2_outputs[505]) | (layer2_outputs[4667]));
    assign layer3_outputs[4028] = layer2_outputs[4008];
    assign layer3_outputs[4029] = layer2_outputs[3636];
    assign layer3_outputs[4030] = (layer2_outputs[1023]) | (layer2_outputs[4449]);
    assign layer3_outputs[4031] = ~(layer2_outputs[3117]);
    assign layer3_outputs[4032] = ~(layer2_outputs[4443]);
    assign layer3_outputs[4033] = (layer2_outputs[4841]) & ~(layer2_outputs[1783]);
    assign layer3_outputs[4034] = ~((layer2_outputs[3386]) | (layer2_outputs[1178]));
    assign layer3_outputs[4035] = ~(layer2_outputs[304]);
    assign layer3_outputs[4036] = ~((layer2_outputs[4415]) & (layer2_outputs[2453]));
    assign layer3_outputs[4037] = ~(layer2_outputs[3416]);
    assign layer3_outputs[4038] = ~(layer2_outputs[4456]) | (layer2_outputs[4794]);
    assign layer3_outputs[4039] = 1'b1;
    assign layer3_outputs[4040] = (layer2_outputs[3566]) & ~(layer2_outputs[1312]);
    assign layer3_outputs[4041] = ~(layer2_outputs[1244]);
    assign layer3_outputs[4042] = (layer2_outputs[3495]) & ~(layer2_outputs[2425]);
    assign layer3_outputs[4043] = ~(layer2_outputs[39]) | (layer2_outputs[1563]);
    assign layer3_outputs[4044] = ~((layer2_outputs[823]) & (layer2_outputs[3043]));
    assign layer3_outputs[4045] = layer2_outputs[4553];
    assign layer3_outputs[4046] = (layer2_outputs[4889]) & ~(layer2_outputs[2718]);
    assign layer3_outputs[4047] = 1'b1;
    assign layer3_outputs[4048] = layer2_outputs[3587];
    assign layer3_outputs[4049] = (layer2_outputs[1431]) | (layer2_outputs[272]);
    assign layer3_outputs[4050] = layer2_outputs[2325];
    assign layer3_outputs[4051] = layer2_outputs[2238];
    assign layer3_outputs[4052] = ~(layer2_outputs[613]);
    assign layer3_outputs[4053] = (layer2_outputs[1874]) & ~(layer2_outputs[4267]);
    assign layer3_outputs[4054] = (layer2_outputs[3276]) | (layer2_outputs[3737]);
    assign layer3_outputs[4055] = layer2_outputs[1634];
    assign layer3_outputs[4056] = ~(layer2_outputs[4598]) | (layer2_outputs[4118]);
    assign layer3_outputs[4057] = ~(layer2_outputs[3833]);
    assign layer3_outputs[4058] = layer2_outputs[3788];
    assign layer3_outputs[4059] = (layer2_outputs[2436]) & ~(layer2_outputs[4337]);
    assign layer3_outputs[4060] = 1'b1;
    assign layer3_outputs[4061] = ~((layer2_outputs[783]) | (layer2_outputs[3180]));
    assign layer3_outputs[4062] = ~((layer2_outputs[4429]) | (layer2_outputs[2633]));
    assign layer3_outputs[4063] = 1'b0;
    assign layer3_outputs[4064] = ~(layer2_outputs[1804]) | (layer2_outputs[1618]);
    assign layer3_outputs[4065] = (layer2_outputs[4420]) & ~(layer2_outputs[433]);
    assign layer3_outputs[4066] = ~((layer2_outputs[5103]) | (layer2_outputs[47]));
    assign layer3_outputs[4067] = ~((layer2_outputs[3197]) | (layer2_outputs[5081]));
    assign layer3_outputs[4068] = layer2_outputs[3724];
    assign layer3_outputs[4069] = 1'b0;
    assign layer3_outputs[4070] = layer2_outputs[3431];
    assign layer3_outputs[4071] = layer2_outputs[2283];
    assign layer3_outputs[4072] = (layer2_outputs[3669]) & ~(layer2_outputs[1266]);
    assign layer3_outputs[4073] = ~(layer2_outputs[4922]) | (layer2_outputs[1074]);
    assign layer3_outputs[4074] = ~(layer2_outputs[3626]);
    assign layer3_outputs[4075] = (layer2_outputs[3416]) & ~(layer2_outputs[792]);
    assign layer3_outputs[4076] = (layer2_outputs[2568]) & (layer2_outputs[2185]);
    assign layer3_outputs[4077] = 1'b0;
    assign layer3_outputs[4078] = ~(layer2_outputs[2827]) | (layer2_outputs[1720]);
    assign layer3_outputs[4079] = ~(layer2_outputs[3877]);
    assign layer3_outputs[4080] = ~((layer2_outputs[3069]) | (layer2_outputs[331]));
    assign layer3_outputs[4081] = (layer2_outputs[2904]) & ~(layer2_outputs[1668]);
    assign layer3_outputs[4082] = (layer2_outputs[1033]) & ~(layer2_outputs[3995]);
    assign layer3_outputs[4083] = 1'b0;
    assign layer3_outputs[4084] = ~(layer2_outputs[1111]);
    assign layer3_outputs[4085] = ~((layer2_outputs[4415]) & (layer2_outputs[365]));
    assign layer3_outputs[4086] = 1'b1;
    assign layer3_outputs[4087] = (layer2_outputs[1692]) & ~(layer2_outputs[3140]);
    assign layer3_outputs[4088] = (layer2_outputs[4631]) & (layer2_outputs[1338]);
    assign layer3_outputs[4089] = 1'b0;
    assign layer3_outputs[4090] = layer2_outputs[2958];
    assign layer3_outputs[4091] = (layer2_outputs[439]) & ~(layer2_outputs[1236]);
    assign layer3_outputs[4092] = ~(layer2_outputs[2276]) | (layer2_outputs[4033]);
    assign layer3_outputs[4093] = ~(layer2_outputs[1932]) | (layer2_outputs[4079]);
    assign layer3_outputs[4094] = ~(layer2_outputs[1034]);
    assign layer3_outputs[4095] = ~(layer2_outputs[4762]);
    assign layer3_outputs[4096] = ~(layer2_outputs[3196]);
    assign layer3_outputs[4097] = ~((layer2_outputs[1757]) ^ (layer2_outputs[347]));
    assign layer3_outputs[4098] = ~(layer2_outputs[2085]);
    assign layer3_outputs[4099] = 1'b1;
    assign layer3_outputs[4100] = (layer2_outputs[3825]) & (layer2_outputs[3171]);
    assign layer3_outputs[4101] = ~((layer2_outputs[4590]) & (layer2_outputs[633]));
    assign layer3_outputs[4102] = ~(layer2_outputs[2912]);
    assign layer3_outputs[4103] = ~((layer2_outputs[376]) | (layer2_outputs[3848]));
    assign layer3_outputs[4104] = ~(layer2_outputs[2176]);
    assign layer3_outputs[4105] = layer2_outputs[4528];
    assign layer3_outputs[4106] = (layer2_outputs[3996]) & (layer2_outputs[2071]);
    assign layer3_outputs[4107] = layer2_outputs[1167];
    assign layer3_outputs[4108] = (layer2_outputs[5033]) & ~(layer2_outputs[514]);
    assign layer3_outputs[4109] = ~(layer2_outputs[5010]) | (layer2_outputs[4297]);
    assign layer3_outputs[4110] = (layer2_outputs[2804]) & ~(layer2_outputs[3951]);
    assign layer3_outputs[4111] = layer2_outputs[3244];
    assign layer3_outputs[4112] = 1'b0;
    assign layer3_outputs[4113] = ~((layer2_outputs[2282]) ^ (layer2_outputs[3288]));
    assign layer3_outputs[4114] = (layer2_outputs[680]) & ~(layer2_outputs[3449]);
    assign layer3_outputs[4115] = layer2_outputs[1291];
    assign layer3_outputs[4116] = (layer2_outputs[4306]) & ~(layer2_outputs[1461]);
    assign layer3_outputs[4117] = ~((layer2_outputs[2025]) & (layer2_outputs[2297]));
    assign layer3_outputs[4118] = (layer2_outputs[3983]) & ~(layer2_outputs[3133]);
    assign layer3_outputs[4119] = ~(layer2_outputs[884]) | (layer2_outputs[3384]);
    assign layer3_outputs[4120] = (layer2_outputs[3818]) & ~(layer2_outputs[4089]);
    assign layer3_outputs[4121] = ~(layer2_outputs[4223]) | (layer2_outputs[3583]);
    assign layer3_outputs[4122] = layer2_outputs[3752];
    assign layer3_outputs[4123] = ~(layer2_outputs[4052]);
    assign layer3_outputs[4124] = ~(layer2_outputs[914]);
    assign layer3_outputs[4125] = ~((layer2_outputs[2545]) & (layer2_outputs[2672]));
    assign layer3_outputs[4126] = ~((layer2_outputs[3602]) ^ (layer2_outputs[3549]));
    assign layer3_outputs[4127] = ~(layer2_outputs[2711]);
    assign layer3_outputs[4128] = 1'b1;
    assign layer3_outputs[4129] = ~(layer2_outputs[1296]) | (layer2_outputs[10]);
    assign layer3_outputs[4130] = ~(layer2_outputs[1257]);
    assign layer3_outputs[4131] = ~((layer2_outputs[1118]) | (layer2_outputs[2975]));
    assign layer3_outputs[4132] = ~(layer2_outputs[304]);
    assign layer3_outputs[4133] = ~(layer2_outputs[2620]);
    assign layer3_outputs[4134] = ~(layer2_outputs[2860]);
    assign layer3_outputs[4135] = layer2_outputs[4907];
    assign layer3_outputs[4136] = layer2_outputs[4646];
    assign layer3_outputs[4137] = (layer2_outputs[4371]) | (layer2_outputs[4545]);
    assign layer3_outputs[4138] = 1'b1;
    assign layer3_outputs[4139] = layer2_outputs[4123];
    assign layer3_outputs[4140] = 1'b1;
    assign layer3_outputs[4141] = layer2_outputs[1674];
    assign layer3_outputs[4142] = ~(layer2_outputs[1161]) | (layer2_outputs[4163]);
    assign layer3_outputs[4143] = ~(layer2_outputs[4857]);
    assign layer3_outputs[4144] = ~((layer2_outputs[1252]) ^ (layer2_outputs[914]));
    assign layer3_outputs[4145] = ~((layer2_outputs[2141]) | (layer2_outputs[4258]));
    assign layer3_outputs[4146] = (layer2_outputs[2112]) | (layer2_outputs[2738]);
    assign layer3_outputs[4147] = ~(layer2_outputs[531]);
    assign layer3_outputs[4148] = ~((layer2_outputs[4813]) ^ (layer2_outputs[3519]));
    assign layer3_outputs[4149] = ~((layer2_outputs[2290]) ^ (layer2_outputs[451]));
    assign layer3_outputs[4150] = ~((layer2_outputs[634]) | (layer2_outputs[3650]));
    assign layer3_outputs[4151] = (layer2_outputs[738]) & ~(layer2_outputs[4018]);
    assign layer3_outputs[4152] = ~(layer2_outputs[995]);
    assign layer3_outputs[4153] = ~((layer2_outputs[4741]) | (layer2_outputs[2813]));
    assign layer3_outputs[4154] = (layer2_outputs[984]) & (layer2_outputs[4256]);
    assign layer3_outputs[4155] = (layer2_outputs[4107]) & ~(layer2_outputs[3132]);
    assign layer3_outputs[4156] = (layer2_outputs[4250]) & (layer2_outputs[4043]);
    assign layer3_outputs[4157] = ~(layer2_outputs[4417]);
    assign layer3_outputs[4158] = (layer2_outputs[2131]) & ~(layer2_outputs[3312]);
    assign layer3_outputs[4159] = layer2_outputs[86];
    assign layer3_outputs[4160] = (layer2_outputs[4877]) | (layer2_outputs[4181]);
    assign layer3_outputs[4161] = ~(layer2_outputs[483]);
    assign layer3_outputs[4162] = ~(layer2_outputs[1070]);
    assign layer3_outputs[4163] = (layer2_outputs[1247]) & (layer2_outputs[4676]);
    assign layer3_outputs[4164] = layer2_outputs[335];
    assign layer3_outputs[4165] = (layer2_outputs[97]) | (layer2_outputs[3285]);
    assign layer3_outputs[4166] = ~(layer2_outputs[2958]);
    assign layer3_outputs[4167] = ~(layer2_outputs[4820]);
    assign layer3_outputs[4168] = (layer2_outputs[2158]) | (layer2_outputs[3039]);
    assign layer3_outputs[4169] = layer2_outputs[1820];
    assign layer3_outputs[4170] = ~(layer2_outputs[1197]) | (layer2_outputs[4154]);
    assign layer3_outputs[4171] = layer2_outputs[86];
    assign layer3_outputs[4172] = (layer2_outputs[459]) & (layer2_outputs[4178]);
    assign layer3_outputs[4173] = ~(layer2_outputs[2475]);
    assign layer3_outputs[4174] = ~(layer2_outputs[1941]);
    assign layer3_outputs[4175] = (layer2_outputs[1590]) | (layer2_outputs[2945]);
    assign layer3_outputs[4176] = ~((layer2_outputs[3690]) & (layer2_outputs[3464]));
    assign layer3_outputs[4177] = ~(layer2_outputs[3359]);
    assign layer3_outputs[4178] = layer2_outputs[3154];
    assign layer3_outputs[4179] = (layer2_outputs[4606]) & ~(layer2_outputs[2873]);
    assign layer3_outputs[4180] = layer2_outputs[1970];
    assign layer3_outputs[4181] = layer2_outputs[2096];
    assign layer3_outputs[4182] = (layer2_outputs[1626]) ^ (layer2_outputs[1619]);
    assign layer3_outputs[4183] = ~(layer2_outputs[284]) | (layer2_outputs[4468]);
    assign layer3_outputs[4184] = 1'b0;
    assign layer3_outputs[4185] = ~((layer2_outputs[979]) | (layer2_outputs[4894]));
    assign layer3_outputs[4186] = ~(layer2_outputs[3059]);
    assign layer3_outputs[4187] = ~(layer2_outputs[3873]);
    assign layer3_outputs[4188] = layer2_outputs[2171];
    assign layer3_outputs[4189] = ~(layer2_outputs[3225]);
    assign layer3_outputs[4190] = ~((layer2_outputs[1222]) | (layer2_outputs[1077]));
    assign layer3_outputs[4191] = ~((layer2_outputs[2862]) | (layer2_outputs[554]));
    assign layer3_outputs[4192] = ~((layer2_outputs[3004]) & (layer2_outputs[2662]));
    assign layer3_outputs[4193] = 1'b1;
    assign layer3_outputs[4194] = (layer2_outputs[1738]) & ~(layer2_outputs[2930]);
    assign layer3_outputs[4195] = (layer2_outputs[2664]) | (layer2_outputs[2153]);
    assign layer3_outputs[4196] = layer2_outputs[3905];
    assign layer3_outputs[4197] = (layer2_outputs[2277]) | (layer2_outputs[4337]);
    assign layer3_outputs[4198] = ~((layer2_outputs[1093]) | (layer2_outputs[2862]));
    assign layer3_outputs[4199] = layer2_outputs[3872];
    assign layer3_outputs[4200] = 1'b1;
    assign layer3_outputs[4201] = ~(layer2_outputs[758]) | (layer2_outputs[3336]);
    assign layer3_outputs[4202] = ~(layer2_outputs[1821]) | (layer2_outputs[1171]);
    assign layer3_outputs[4203] = layer2_outputs[4618];
    assign layer3_outputs[4204] = ~((layer2_outputs[1301]) & (layer2_outputs[3745]));
    assign layer3_outputs[4205] = layer2_outputs[3831];
    assign layer3_outputs[4206] = ~((layer2_outputs[3304]) | (layer2_outputs[961]));
    assign layer3_outputs[4207] = ~((layer2_outputs[1737]) & (layer2_outputs[1719]));
    assign layer3_outputs[4208] = ~((layer2_outputs[3631]) | (layer2_outputs[719]));
    assign layer3_outputs[4209] = ~(layer2_outputs[5059]) | (layer2_outputs[2396]);
    assign layer3_outputs[4210] = (layer2_outputs[4166]) | (layer2_outputs[4091]);
    assign layer3_outputs[4211] = layer2_outputs[1353];
    assign layer3_outputs[4212] = 1'b0;
    assign layer3_outputs[4213] = (layer2_outputs[4979]) & (layer2_outputs[2853]);
    assign layer3_outputs[4214] = (layer2_outputs[2942]) | (layer2_outputs[2278]);
    assign layer3_outputs[4215] = ~(layer2_outputs[2605]);
    assign layer3_outputs[4216] = (layer2_outputs[297]) & ~(layer2_outputs[5103]);
    assign layer3_outputs[4217] = ~(layer2_outputs[1631]) | (layer2_outputs[2335]);
    assign layer3_outputs[4218] = (layer2_outputs[546]) & (layer2_outputs[4486]);
    assign layer3_outputs[4219] = (layer2_outputs[1712]) & ~(layer2_outputs[3412]);
    assign layer3_outputs[4220] = ~((layer2_outputs[1724]) | (layer2_outputs[3880]));
    assign layer3_outputs[4221] = 1'b1;
    assign layer3_outputs[4222] = ~(layer2_outputs[2623]);
    assign layer3_outputs[4223] = ~(layer2_outputs[1633]);
    assign layer3_outputs[4224] = (layer2_outputs[2768]) & (layer2_outputs[2339]);
    assign layer3_outputs[4225] = ~(layer2_outputs[3166]) | (layer2_outputs[2584]);
    assign layer3_outputs[4226] = (layer2_outputs[3189]) & (layer2_outputs[1792]);
    assign layer3_outputs[4227] = ~((layer2_outputs[4027]) | (layer2_outputs[474]));
    assign layer3_outputs[4228] = 1'b1;
    assign layer3_outputs[4229] = layer2_outputs[4688];
    assign layer3_outputs[4230] = ~(layer2_outputs[3966]);
    assign layer3_outputs[4231] = layer2_outputs[1060];
    assign layer3_outputs[4232] = ~(layer2_outputs[584]);
    assign layer3_outputs[4233] = 1'b1;
    assign layer3_outputs[4234] = (layer2_outputs[4128]) & ~(layer2_outputs[3654]);
    assign layer3_outputs[4235] = ~(layer2_outputs[4028]) | (layer2_outputs[4408]);
    assign layer3_outputs[4236] = (layer2_outputs[161]) & ~(layer2_outputs[2731]);
    assign layer3_outputs[4237] = layer2_outputs[4162];
    assign layer3_outputs[4238] = (layer2_outputs[4701]) & ~(layer2_outputs[697]);
    assign layer3_outputs[4239] = layer2_outputs[3931];
    assign layer3_outputs[4240] = ~(layer2_outputs[2870]);
    assign layer3_outputs[4241] = (layer2_outputs[296]) & (layer2_outputs[4897]);
    assign layer3_outputs[4242] = ~(layer2_outputs[1092]);
    assign layer3_outputs[4243] = ~(layer2_outputs[2312]);
    assign layer3_outputs[4244] = layer2_outputs[4748];
    assign layer3_outputs[4245] = layer2_outputs[387];
    assign layer3_outputs[4246] = (layer2_outputs[5085]) & ~(layer2_outputs[2426]);
    assign layer3_outputs[4247] = (layer2_outputs[4613]) ^ (layer2_outputs[1765]);
    assign layer3_outputs[4248] = ~(layer2_outputs[2384]) | (layer2_outputs[2322]);
    assign layer3_outputs[4249] = ~((layer2_outputs[3720]) ^ (layer2_outputs[5104]));
    assign layer3_outputs[4250] = ~(layer2_outputs[1337]) | (layer2_outputs[3489]);
    assign layer3_outputs[4251] = ~(layer2_outputs[967]);
    assign layer3_outputs[4252] = 1'b1;
    assign layer3_outputs[4253] = layer2_outputs[23];
    assign layer3_outputs[4254] = (layer2_outputs[1307]) & ~(layer2_outputs[4803]);
    assign layer3_outputs[4255] = (layer2_outputs[3138]) & ~(layer2_outputs[4800]);
    assign layer3_outputs[4256] = (layer2_outputs[363]) & (layer2_outputs[2354]);
    assign layer3_outputs[4257] = (layer2_outputs[1799]) & (layer2_outputs[4765]);
    assign layer3_outputs[4258] = layer2_outputs[3505];
    assign layer3_outputs[4259] = (layer2_outputs[1016]) & ~(layer2_outputs[3479]);
    assign layer3_outputs[4260] = (layer2_outputs[1033]) & ~(layer2_outputs[897]);
    assign layer3_outputs[4261] = ~((layer2_outputs[3188]) | (layer2_outputs[1182]));
    assign layer3_outputs[4262] = (layer2_outputs[766]) & ~(layer2_outputs[3535]);
    assign layer3_outputs[4263] = (layer2_outputs[5038]) & (layer2_outputs[3832]);
    assign layer3_outputs[4264] = ~(layer2_outputs[936]) | (layer2_outputs[3660]);
    assign layer3_outputs[4265] = ~(layer2_outputs[1519]);
    assign layer3_outputs[4266] = (layer2_outputs[3296]) & (layer2_outputs[3950]);
    assign layer3_outputs[4267] = (layer2_outputs[4315]) & ~(layer2_outputs[1285]);
    assign layer3_outputs[4268] = ~(layer2_outputs[358]) | (layer2_outputs[46]);
    assign layer3_outputs[4269] = (layer2_outputs[3670]) & ~(layer2_outputs[2963]);
    assign layer3_outputs[4270] = ~(layer2_outputs[315]);
    assign layer3_outputs[4271] = 1'b0;
    assign layer3_outputs[4272] = layer2_outputs[3813];
    assign layer3_outputs[4273] = ~(layer2_outputs[1131]) | (layer2_outputs[361]);
    assign layer3_outputs[4274] = layer2_outputs[3003];
    assign layer3_outputs[4275] = (layer2_outputs[1321]) & ~(layer2_outputs[778]);
    assign layer3_outputs[4276] = ~((layer2_outputs[3710]) & (layer2_outputs[167]));
    assign layer3_outputs[4277] = ~(layer2_outputs[4863]);
    assign layer3_outputs[4278] = (layer2_outputs[2020]) & ~(layer2_outputs[364]);
    assign layer3_outputs[4279] = ~((layer2_outputs[2175]) & (layer2_outputs[2803]));
    assign layer3_outputs[4280] = layer2_outputs[1616];
    assign layer3_outputs[4281] = ~((layer2_outputs[240]) & (layer2_outputs[4913]));
    assign layer3_outputs[4282] = layer2_outputs[1973];
    assign layer3_outputs[4283] = ~(layer2_outputs[2412]);
    assign layer3_outputs[4284] = ~(layer2_outputs[4269]) | (layer2_outputs[2916]);
    assign layer3_outputs[4285] = 1'b1;
    assign layer3_outputs[4286] = layer2_outputs[3826];
    assign layer3_outputs[4287] = ~(layer2_outputs[4747]);
    assign layer3_outputs[4288] = (layer2_outputs[4596]) & ~(layer2_outputs[3901]);
    assign layer3_outputs[4289] = layer2_outputs[3249];
    assign layer3_outputs[4290] = ~((layer2_outputs[4888]) | (layer2_outputs[2191]));
    assign layer3_outputs[4291] = (layer2_outputs[4704]) | (layer2_outputs[3394]);
    assign layer3_outputs[4292] = layer2_outputs[2315];
    assign layer3_outputs[4293] = ~((layer2_outputs[2705]) | (layer2_outputs[1066]));
    assign layer3_outputs[4294] = 1'b0;
    assign layer3_outputs[4295] = layer2_outputs[1924];
    assign layer3_outputs[4296] = layer2_outputs[3407];
    assign layer3_outputs[4297] = ~((layer2_outputs[83]) & (layer2_outputs[3620]));
    assign layer3_outputs[4298] = layer2_outputs[4482];
    assign layer3_outputs[4299] = layer2_outputs[1297];
    assign layer3_outputs[4300] = 1'b1;
    assign layer3_outputs[4301] = ~(layer2_outputs[4190]);
    assign layer3_outputs[4302] = (layer2_outputs[2224]) & ~(layer2_outputs[525]);
    assign layer3_outputs[4303] = ~(layer2_outputs[4693]);
    assign layer3_outputs[4304] = 1'b1;
    assign layer3_outputs[4305] = ~((layer2_outputs[3737]) ^ (layer2_outputs[3338]));
    assign layer3_outputs[4306] = layer2_outputs[3504];
    assign layer3_outputs[4307] = layer2_outputs[155];
    assign layer3_outputs[4308] = (layer2_outputs[2248]) & ~(layer2_outputs[1257]);
    assign layer3_outputs[4309] = (layer2_outputs[4317]) & (layer2_outputs[2509]);
    assign layer3_outputs[4310] = ~((layer2_outputs[128]) ^ (layer2_outputs[2103]));
    assign layer3_outputs[4311] = ~(layer2_outputs[4402]);
    assign layer3_outputs[4312] = 1'b1;
    assign layer3_outputs[4313] = ~(layer2_outputs[2271]);
    assign layer3_outputs[4314] = (layer2_outputs[1202]) & (layer2_outputs[1182]);
    assign layer3_outputs[4315] = 1'b0;
    assign layer3_outputs[4316] = ~(layer2_outputs[2027]);
    assign layer3_outputs[4317] = (layer2_outputs[4346]) | (layer2_outputs[1530]);
    assign layer3_outputs[4318] = layer2_outputs[4229];
    assign layer3_outputs[4319] = 1'b0;
    assign layer3_outputs[4320] = 1'b0;
    assign layer3_outputs[4321] = ~(layer2_outputs[4241]);
    assign layer3_outputs[4322] = ~(layer2_outputs[4770]);
    assign layer3_outputs[4323] = ~(layer2_outputs[1750]) | (layer2_outputs[3589]);
    assign layer3_outputs[4324] = 1'b1;
    assign layer3_outputs[4325] = (layer2_outputs[4234]) | (layer2_outputs[1248]);
    assign layer3_outputs[4326] = ~(layer2_outputs[4260]) | (layer2_outputs[1282]);
    assign layer3_outputs[4327] = ~(layer2_outputs[384]);
    assign layer3_outputs[4328] = (layer2_outputs[5076]) & ~(layer2_outputs[3266]);
    assign layer3_outputs[4329] = ~(layer2_outputs[2659]) | (layer2_outputs[4961]);
    assign layer3_outputs[4330] = ~(layer2_outputs[132]);
    assign layer3_outputs[4331] = layer2_outputs[2604];
    assign layer3_outputs[4332] = layer2_outputs[2187];
    assign layer3_outputs[4333] = layer2_outputs[436];
    assign layer3_outputs[4334] = ~((layer2_outputs[3526]) ^ (layer2_outputs[4326]));
    assign layer3_outputs[4335] = ~(layer2_outputs[4761]);
    assign layer3_outputs[4336] = ~((layer2_outputs[5042]) | (layer2_outputs[742]));
    assign layer3_outputs[4337] = (layer2_outputs[2317]) ^ (layer2_outputs[2504]);
    assign layer3_outputs[4338] = (layer2_outputs[601]) & ~(layer2_outputs[1245]);
    assign layer3_outputs[4339] = ~((layer2_outputs[4715]) & (layer2_outputs[4866]));
    assign layer3_outputs[4340] = 1'b1;
    assign layer3_outputs[4341] = layer2_outputs[2169];
    assign layer3_outputs[4342] = 1'b0;
    assign layer3_outputs[4343] = 1'b1;
    assign layer3_outputs[4344] = layer2_outputs[3661];
    assign layer3_outputs[4345] = layer2_outputs[3027];
    assign layer3_outputs[4346] = ~((layer2_outputs[864]) | (layer2_outputs[2225]));
    assign layer3_outputs[4347] = ~((layer2_outputs[3559]) | (layer2_outputs[802]));
    assign layer3_outputs[4348] = layer2_outputs[1587];
    assign layer3_outputs[4349] = ~(layer2_outputs[530]) | (layer2_outputs[4554]);
    assign layer3_outputs[4350] = (layer2_outputs[2897]) & ~(layer2_outputs[1762]);
    assign layer3_outputs[4351] = layer2_outputs[2790];
    assign layer3_outputs[4352] = ~(layer2_outputs[2895]);
    assign layer3_outputs[4353] = ~((layer2_outputs[4010]) ^ (layer2_outputs[5093]));
    assign layer3_outputs[4354] = (layer2_outputs[717]) & (layer2_outputs[1156]);
    assign layer3_outputs[4355] = ~((layer2_outputs[3531]) & (layer2_outputs[850]));
    assign layer3_outputs[4356] = 1'b1;
    assign layer3_outputs[4357] = (layer2_outputs[2880]) ^ (layer2_outputs[5077]);
    assign layer3_outputs[4358] = ~(layer2_outputs[3599]) | (layer2_outputs[2105]);
    assign layer3_outputs[4359] = ~(layer2_outputs[2793]) | (layer2_outputs[526]);
    assign layer3_outputs[4360] = layer2_outputs[2700];
    assign layer3_outputs[4361] = ~(layer2_outputs[3024]);
    assign layer3_outputs[4362] = (layer2_outputs[2065]) | (layer2_outputs[332]);
    assign layer3_outputs[4363] = layer2_outputs[1348];
    assign layer3_outputs[4364] = layer2_outputs[1150];
    assign layer3_outputs[4365] = (layer2_outputs[1175]) | (layer2_outputs[3071]);
    assign layer3_outputs[4366] = (layer2_outputs[1702]) & ~(layer2_outputs[2356]);
    assign layer3_outputs[4367] = (layer2_outputs[1891]) & ~(layer2_outputs[3609]);
    assign layer3_outputs[4368] = (layer2_outputs[135]) | (layer2_outputs[4972]);
    assign layer3_outputs[4369] = (layer2_outputs[1852]) & (layer2_outputs[4307]);
    assign layer3_outputs[4370] = layer2_outputs[224];
    assign layer3_outputs[4371] = (layer2_outputs[2066]) & (layer2_outputs[4214]);
    assign layer3_outputs[4372] = 1'b0;
    assign layer3_outputs[4373] = (layer2_outputs[294]) & ~(layer2_outputs[4472]);
    assign layer3_outputs[4374] = 1'b1;
    assign layer3_outputs[4375] = layer2_outputs[3415];
    assign layer3_outputs[4376] = (layer2_outputs[166]) & ~(layer2_outputs[3029]);
    assign layer3_outputs[4377] = (layer2_outputs[2361]) & ~(layer2_outputs[66]);
    assign layer3_outputs[4378] = layer2_outputs[593];
    assign layer3_outputs[4379] = ~(layer2_outputs[1574]) | (layer2_outputs[4313]);
    assign layer3_outputs[4380] = ~(layer2_outputs[2345]) | (layer2_outputs[2006]);
    assign layer3_outputs[4381] = ~((layer2_outputs[4645]) | (layer2_outputs[2611]));
    assign layer3_outputs[4382] = ~(layer2_outputs[4136]) | (layer2_outputs[2035]);
    assign layer3_outputs[4383] = 1'b0;
    assign layer3_outputs[4384] = ~((layer2_outputs[4667]) & (layer2_outputs[3078]));
    assign layer3_outputs[4385] = (layer2_outputs[553]) & (layer2_outputs[2321]);
    assign layer3_outputs[4386] = (layer2_outputs[1706]) ^ (layer2_outputs[3186]);
    assign layer3_outputs[4387] = ~(layer2_outputs[266]);
    assign layer3_outputs[4388] = ~((layer2_outputs[5094]) & (layer2_outputs[1496]));
    assign layer3_outputs[4389] = ~(layer2_outputs[3317]) | (layer2_outputs[1427]);
    assign layer3_outputs[4390] = (layer2_outputs[2212]) ^ (layer2_outputs[163]);
    assign layer3_outputs[4391] = (layer2_outputs[1036]) ^ (layer2_outputs[819]);
    assign layer3_outputs[4392] = (layer2_outputs[5054]) & ~(layer2_outputs[3695]);
    assign layer3_outputs[4393] = ~(layer2_outputs[2388]) | (layer2_outputs[2109]);
    assign layer3_outputs[4394] = 1'b0;
    assign layer3_outputs[4395] = ~(layer2_outputs[3972]) | (layer2_outputs[1482]);
    assign layer3_outputs[4396] = (layer2_outputs[4768]) & ~(layer2_outputs[4209]);
    assign layer3_outputs[4397] = ~((layer2_outputs[1158]) | (layer2_outputs[3601]));
    assign layer3_outputs[4398] = ~((layer2_outputs[4547]) | (layer2_outputs[525]));
    assign layer3_outputs[4399] = ~(layer2_outputs[1804]);
    assign layer3_outputs[4400] = 1'b1;
    assign layer3_outputs[4401] = ~(layer2_outputs[2091]);
    assign layer3_outputs[4402] = ~(layer2_outputs[2355]) | (layer2_outputs[451]);
    assign layer3_outputs[4403] = (layer2_outputs[3714]) | (layer2_outputs[1963]);
    assign layer3_outputs[4404] = layer2_outputs[1180];
    assign layer3_outputs[4405] = layer2_outputs[1644];
    assign layer3_outputs[4406] = layer2_outputs[4727];
    assign layer3_outputs[4407] = layer2_outputs[1937];
    assign layer3_outputs[4408] = ~((layer2_outputs[821]) | (layer2_outputs[1389]));
    assign layer3_outputs[4409] = 1'b1;
    assign layer3_outputs[4410] = ~(layer2_outputs[3600]);
    assign layer3_outputs[4411] = 1'b0;
    assign layer3_outputs[4412] = ~(layer2_outputs[910]);
    assign layer3_outputs[4413] = layer2_outputs[1339];
    assign layer3_outputs[4414] = layer2_outputs[4356];
    assign layer3_outputs[4415] = layer2_outputs[3359];
    assign layer3_outputs[4416] = (layer2_outputs[5015]) & (layer2_outputs[381]);
    assign layer3_outputs[4417] = ~(layer2_outputs[2899]);
    assign layer3_outputs[4418] = layer2_outputs[96];
    assign layer3_outputs[4419] = ~(layer2_outputs[1886]) | (layer2_outputs[1222]);
    assign layer3_outputs[4420] = ~((layer2_outputs[217]) | (layer2_outputs[5016]));
    assign layer3_outputs[4421] = ~((layer2_outputs[177]) & (layer2_outputs[207]));
    assign layer3_outputs[4422] = (layer2_outputs[3278]) & ~(layer2_outputs[3882]);
    assign layer3_outputs[4423] = (layer2_outputs[1751]) & ~(layer2_outputs[4846]);
    assign layer3_outputs[4424] = ~(layer2_outputs[5022]) | (layer2_outputs[2373]);
    assign layer3_outputs[4425] = (layer2_outputs[2503]) & (layer2_outputs[4208]);
    assign layer3_outputs[4426] = ~((layer2_outputs[4177]) & (layer2_outputs[4391]));
    assign layer3_outputs[4427] = layer2_outputs[751];
    assign layer3_outputs[4428] = ~(layer2_outputs[1183]);
    assign layer3_outputs[4429] = ~(layer2_outputs[3245]);
    assign layer3_outputs[4430] = ~(layer2_outputs[4795]);
    assign layer3_outputs[4431] = ~(layer2_outputs[3753]);
    assign layer3_outputs[4432] = (layer2_outputs[699]) | (layer2_outputs[578]);
    assign layer3_outputs[4433] = (layer2_outputs[2598]) & ~(layer2_outputs[1080]);
    assign layer3_outputs[4434] = ~((layer2_outputs[3206]) & (layer2_outputs[4014]));
    assign layer3_outputs[4435] = layer2_outputs[3397];
    assign layer3_outputs[4436] = 1'b1;
    assign layer3_outputs[4437] = 1'b0;
    assign layer3_outputs[4438] = ~(layer2_outputs[248]) | (layer2_outputs[1850]);
    assign layer3_outputs[4439] = (layer2_outputs[4948]) & (layer2_outputs[4448]);
    assign layer3_outputs[4440] = 1'b0;
    assign layer3_outputs[4441] = ~((layer2_outputs[3894]) & (layer2_outputs[4908]));
    assign layer3_outputs[4442] = (layer2_outputs[5100]) | (layer2_outputs[1797]);
    assign layer3_outputs[4443] = ~(layer2_outputs[4381]);
    assign layer3_outputs[4444] = (layer2_outputs[2340]) & (layer2_outputs[2574]);
    assign layer3_outputs[4445] = (layer2_outputs[576]) & (layer2_outputs[2438]);
    assign layer3_outputs[4446] = (layer2_outputs[3067]) & ~(layer2_outputs[2950]);
    assign layer3_outputs[4447] = ~(layer2_outputs[1366]) | (layer2_outputs[4887]);
    assign layer3_outputs[4448] = (layer2_outputs[1847]) | (layer2_outputs[1128]);
    assign layer3_outputs[4449] = ~(layer2_outputs[1341]) | (layer2_outputs[4702]);
    assign layer3_outputs[4450] = layer2_outputs[4659];
    assign layer3_outputs[4451] = ~((layer2_outputs[1358]) & (layer2_outputs[3082]));
    assign layer3_outputs[4452] = layer2_outputs[1381];
    assign layer3_outputs[4453] = (layer2_outputs[3642]) & ~(layer2_outputs[1849]);
    assign layer3_outputs[4454] = layer2_outputs[2653];
    assign layer3_outputs[4455] = ~(layer2_outputs[49]) | (layer2_outputs[849]);
    assign layer3_outputs[4456] = layer2_outputs[4723];
    assign layer3_outputs[4457] = 1'b1;
    assign layer3_outputs[4458] = ~(layer2_outputs[3402]) | (layer2_outputs[685]);
    assign layer3_outputs[4459] = 1'b0;
    assign layer3_outputs[4460] = ~(layer2_outputs[1623]);
    assign layer3_outputs[4461] = layer2_outputs[3475];
    assign layer3_outputs[4462] = layer2_outputs[611];
    assign layer3_outputs[4463] = (layer2_outputs[1137]) & ~(layer2_outputs[5104]);
    assign layer3_outputs[4464] = (layer2_outputs[477]) | (layer2_outputs[875]);
    assign layer3_outputs[4465] = (layer2_outputs[2350]) & (layer2_outputs[2347]);
    assign layer3_outputs[4466] = ~((layer2_outputs[3723]) & (layer2_outputs[4201]));
    assign layer3_outputs[4467] = ~(layer2_outputs[4574]);
    assign layer3_outputs[4468] = ~((layer2_outputs[1848]) & (layer2_outputs[3706]));
    assign layer3_outputs[4469] = ~((layer2_outputs[495]) | (layer2_outputs[4996]));
    assign layer3_outputs[4470] = ~(layer2_outputs[4569]);
    assign layer3_outputs[4471] = ~((layer2_outputs[289]) & (layer2_outputs[2021]));
    assign layer3_outputs[4472] = 1'b1;
    assign layer3_outputs[4473] = ~(layer2_outputs[4251]) | (layer2_outputs[4378]);
    assign layer3_outputs[4474] = 1'b0;
    assign layer3_outputs[4475] = layer2_outputs[807];
    assign layer3_outputs[4476] = (layer2_outputs[4474]) | (layer2_outputs[349]);
    assign layer3_outputs[4477] = (layer2_outputs[4597]) | (layer2_outputs[2972]);
    assign layer3_outputs[4478] = ~(layer2_outputs[2791]);
    assign layer3_outputs[4479] = ~(layer2_outputs[4846]);
    assign layer3_outputs[4480] = ~((layer2_outputs[230]) | (layer2_outputs[78]));
    assign layer3_outputs[4481] = 1'b0;
    assign layer3_outputs[4482] = ~((layer2_outputs[3079]) | (layer2_outputs[4254]));
    assign layer3_outputs[4483] = ~((layer2_outputs[3623]) | (layer2_outputs[4605]));
    assign layer3_outputs[4484] = layer2_outputs[2535];
    assign layer3_outputs[4485] = (layer2_outputs[1594]) & ~(layer2_outputs[1498]);
    assign layer3_outputs[4486] = layer2_outputs[633];
    assign layer3_outputs[4487] = (layer2_outputs[2365]) ^ (layer2_outputs[2858]);
    assign layer3_outputs[4488] = 1'b0;
    assign layer3_outputs[4489] = (layer2_outputs[3120]) & ~(layer2_outputs[4795]);
    assign layer3_outputs[4490] = (layer2_outputs[4573]) & ~(layer2_outputs[800]);
    assign layer3_outputs[4491] = (layer2_outputs[1392]) & ~(layer2_outputs[4377]);
    assign layer3_outputs[4492] = ~(layer2_outputs[1944]);
    assign layer3_outputs[4493] = ~(layer2_outputs[528]);
    assign layer3_outputs[4494] = (layer2_outputs[2354]) & ~(layer2_outputs[2168]);
    assign layer3_outputs[4495] = (layer2_outputs[2641]) & ~(layer2_outputs[1262]);
    assign layer3_outputs[4496] = ~((layer2_outputs[1317]) & (layer2_outputs[1477]));
    assign layer3_outputs[4497] = (layer2_outputs[2218]) & ~(layer2_outputs[3978]);
    assign layer3_outputs[4498] = ~(layer2_outputs[1026]) | (layer2_outputs[1669]);
    assign layer3_outputs[4499] = ~(layer2_outputs[3813]);
    assign layer3_outputs[4500] = ~(layer2_outputs[2756]) | (layer2_outputs[695]);
    assign layer3_outputs[4501] = ~(layer2_outputs[3171]);
    assign layer3_outputs[4502] = (layer2_outputs[4357]) & ~(layer2_outputs[223]);
    assign layer3_outputs[4503] = ~(layer2_outputs[4938]);
    assign layer3_outputs[4504] = (layer2_outputs[3457]) & (layer2_outputs[1674]);
    assign layer3_outputs[4505] = 1'b1;
    assign layer3_outputs[4506] = 1'b1;
    assign layer3_outputs[4507] = 1'b1;
    assign layer3_outputs[4508] = ~(layer2_outputs[1275]) | (layer2_outputs[1314]);
    assign layer3_outputs[4509] = 1'b1;
    assign layer3_outputs[4510] = layer2_outputs[1367];
    assign layer3_outputs[4511] = layer2_outputs[4365];
    assign layer3_outputs[4512] = 1'b1;
    assign layer3_outputs[4513] = (layer2_outputs[3685]) | (layer2_outputs[2401]);
    assign layer3_outputs[4514] = (layer2_outputs[2364]) & ~(layer2_outputs[1468]);
    assign layer3_outputs[4515] = ~((layer2_outputs[3563]) | (layer2_outputs[10]));
    assign layer3_outputs[4516] = layer2_outputs[1780];
    assign layer3_outputs[4517] = (layer2_outputs[5008]) & ~(layer2_outputs[3822]);
    assign layer3_outputs[4518] = ~((layer2_outputs[941]) | (layer2_outputs[4926]));
    assign layer3_outputs[4519] = (layer2_outputs[4687]) & ~(layer2_outputs[3335]);
    assign layer3_outputs[4520] = layer2_outputs[150];
    assign layer3_outputs[4521] = layer2_outputs[3227];
    assign layer3_outputs[4522] = ~(layer2_outputs[754]);
    assign layer3_outputs[4523] = ~(layer2_outputs[4007]);
    assign layer3_outputs[4524] = (layer2_outputs[2046]) & ~(layer2_outputs[987]);
    assign layer3_outputs[4525] = ~(layer2_outputs[3952]);
    assign layer3_outputs[4526] = 1'b0;
    assign layer3_outputs[4527] = 1'b1;
    assign layer3_outputs[4528] = 1'b1;
    assign layer3_outputs[4529] = layer2_outputs[4692];
    assign layer3_outputs[4530] = ~(layer2_outputs[1843]);
    assign layer3_outputs[4531] = 1'b1;
    assign layer3_outputs[4532] = (layer2_outputs[1026]) & ~(layer2_outputs[4261]);
    assign layer3_outputs[4533] = layer2_outputs[3125];
    assign layer3_outputs[4534] = ~(layer2_outputs[1879]) | (layer2_outputs[692]);
    assign layer3_outputs[4535] = layer2_outputs[222];
    assign layer3_outputs[4536] = ~(layer2_outputs[3616]);
    assign layer3_outputs[4537] = 1'b1;
    assign layer3_outputs[4538] = (layer2_outputs[3434]) & ~(layer2_outputs[2233]);
    assign layer3_outputs[4539] = layer2_outputs[1896];
    assign layer3_outputs[4540] = layer2_outputs[2655];
    assign layer3_outputs[4541] = layer2_outputs[2850];
    assign layer3_outputs[4542] = layer2_outputs[5086];
    assign layer3_outputs[4543] = ~((layer2_outputs[1069]) & (layer2_outputs[1281]));
    assign layer3_outputs[4544] = layer2_outputs[4693];
    assign layer3_outputs[4545] = 1'b1;
    assign layer3_outputs[4546] = (layer2_outputs[26]) & (layer2_outputs[4810]);
    assign layer3_outputs[4547] = (layer2_outputs[2353]) & ~(layer2_outputs[139]);
    assign layer3_outputs[4548] = ~(layer2_outputs[1701]);
    assign layer3_outputs[4549] = layer2_outputs[1600];
    assign layer3_outputs[4550] = layer2_outputs[1947];
    assign layer3_outputs[4551] = 1'b1;
    assign layer3_outputs[4552] = ~(layer2_outputs[1585]) | (layer2_outputs[1450]);
    assign layer3_outputs[4553] = layer2_outputs[1384];
    assign layer3_outputs[4554] = ~(layer2_outputs[1579]);
    assign layer3_outputs[4555] = ~((layer2_outputs[858]) ^ (layer2_outputs[667]));
    assign layer3_outputs[4556] = 1'b1;
    assign layer3_outputs[4557] = ~((layer2_outputs[4564]) & (layer2_outputs[2389]));
    assign layer3_outputs[4558] = ~(layer2_outputs[1515]);
    assign layer3_outputs[4559] = ~((layer2_outputs[2866]) & (layer2_outputs[1898]));
    assign layer3_outputs[4560] = 1'b1;
    assign layer3_outputs[4561] = layer2_outputs[2940];
    assign layer3_outputs[4562] = layer2_outputs[1529];
    assign layer3_outputs[4563] = layer2_outputs[4678];
    assign layer3_outputs[4564] = layer2_outputs[4362];
    assign layer3_outputs[4565] = 1'b1;
    assign layer3_outputs[4566] = layer2_outputs[2383];
    assign layer3_outputs[4567] = ~((layer2_outputs[3047]) & (layer2_outputs[3548]));
    assign layer3_outputs[4568] = 1'b0;
    assign layer3_outputs[4569] = layer2_outputs[2733];
    assign layer3_outputs[4570] = ~(layer2_outputs[3181]) | (layer2_outputs[1056]);
    assign layer3_outputs[4571] = layer2_outputs[3614];
    assign layer3_outputs[4572] = (layer2_outputs[359]) & ~(layer2_outputs[1538]);
    assign layer3_outputs[4573] = 1'b1;
    assign layer3_outputs[4574] = layer2_outputs[4947];
    assign layer3_outputs[4575] = 1'b0;
    assign layer3_outputs[4576] = ~(layer2_outputs[657]) | (layer2_outputs[1254]);
    assign layer3_outputs[4577] = (layer2_outputs[1072]) & ~(layer2_outputs[4389]);
    assign layer3_outputs[4578] = layer2_outputs[4358];
    assign layer3_outputs[4579] = layer2_outputs[3890];
    assign layer3_outputs[4580] = ~(layer2_outputs[1962]) | (layer2_outputs[3534]);
    assign layer3_outputs[4581] = layer2_outputs[2169];
    assign layer3_outputs[4582] = ~(layer2_outputs[3364]);
    assign layer3_outputs[4583] = 1'b0;
    assign layer3_outputs[4584] = (layer2_outputs[3427]) & ~(layer2_outputs[36]);
    assign layer3_outputs[4585] = (layer2_outputs[3019]) & ~(layer2_outputs[538]);
    assign layer3_outputs[4586] = ~((layer2_outputs[3220]) | (layer2_outputs[4917]));
    assign layer3_outputs[4587] = (layer2_outputs[1474]) ^ (layer2_outputs[4635]);
    assign layer3_outputs[4588] = (layer2_outputs[3202]) & (layer2_outputs[3825]);
    assign layer3_outputs[4589] = layer2_outputs[447];
    assign layer3_outputs[4590] = 1'b1;
    assign layer3_outputs[4591] = layer2_outputs[3493];
    assign layer3_outputs[4592] = ~((layer2_outputs[866]) & (layer2_outputs[3933]));
    assign layer3_outputs[4593] = layer2_outputs[4388];
    assign layer3_outputs[4594] = (layer2_outputs[2831]) | (layer2_outputs[951]);
    assign layer3_outputs[4595] = (layer2_outputs[423]) & (layer2_outputs[4238]);
    assign layer3_outputs[4596] = (layer2_outputs[4733]) & ~(layer2_outputs[4859]);
    assign layer3_outputs[4597] = ~(layer2_outputs[3371]) | (layer2_outputs[3020]);
    assign layer3_outputs[4598] = ~(layer2_outputs[1845]);
    assign layer3_outputs[4599] = ~((layer2_outputs[4628]) & (layer2_outputs[2517]));
    assign layer3_outputs[4600] = ~(layer2_outputs[4765]);
    assign layer3_outputs[4601] = layer2_outputs[1658];
    assign layer3_outputs[4602] = ~(layer2_outputs[4543]) | (layer2_outputs[2194]);
    assign layer3_outputs[4603] = layer2_outputs[3738];
    assign layer3_outputs[4604] = layer2_outputs[4973];
    assign layer3_outputs[4605] = 1'b1;
    assign layer3_outputs[4606] = ~(layer2_outputs[1877]);
    assign layer3_outputs[4607] = 1'b0;
    assign layer3_outputs[4608] = 1'b1;
    assign layer3_outputs[4609] = ~(layer2_outputs[1061]);
    assign layer3_outputs[4610] = 1'b0;
    assign layer3_outputs[4611] = ~(layer2_outputs[4230]) | (layer2_outputs[2291]);
    assign layer3_outputs[4612] = (layer2_outputs[3425]) & ~(layer2_outputs[4075]);
    assign layer3_outputs[4613] = ~(layer2_outputs[1901]);
    assign layer3_outputs[4614] = ~(layer2_outputs[3658]);
    assign layer3_outputs[4615] = ~(layer2_outputs[1099]) | (layer2_outputs[4094]);
    assign layer3_outputs[4616] = (layer2_outputs[663]) & ~(layer2_outputs[4171]);
    assign layer3_outputs[4617] = layer2_outputs[1855];
    assign layer3_outputs[4618] = (layer2_outputs[4054]) & ~(layer2_outputs[4497]);
    assign layer3_outputs[4619] = (layer2_outputs[1315]) & ~(layer2_outputs[3329]);
    assign layer3_outputs[4620] = ~(layer2_outputs[2830]) | (layer2_outputs[2282]);
    assign layer3_outputs[4621] = ~(layer2_outputs[5101]);
    assign layer3_outputs[4622] = layer2_outputs[295];
    assign layer3_outputs[4623] = ~(layer2_outputs[5043]);
    assign layer3_outputs[4624] = layer2_outputs[27];
    assign layer3_outputs[4625] = ~((layer2_outputs[3504]) | (layer2_outputs[1427]));
    assign layer3_outputs[4626] = ~(layer2_outputs[3637]) | (layer2_outputs[4533]);
    assign layer3_outputs[4627] = ~(layer2_outputs[3662]);
    assign layer3_outputs[4628] = ~(layer2_outputs[562]);
    assign layer3_outputs[4629] = ~((layer2_outputs[1363]) & (layer2_outputs[345]));
    assign layer3_outputs[4630] = (layer2_outputs[658]) | (layer2_outputs[9]);
    assign layer3_outputs[4631] = ~(layer2_outputs[1593]);
    assign layer3_outputs[4632] = ~(layer2_outputs[1802]);
    assign layer3_outputs[4633] = (layer2_outputs[1618]) | (layer2_outputs[93]);
    assign layer3_outputs[4634] = ~((layer2_outputs[51]) & (layer2_outputs[3042]));
    assign layer3_outputs[4635] = ~(layer2_outputs[1365]);
    assign layer3_outputs[4636] = ~(layer2_outputs[2536]);
    assign layer3_outputs[4637] = ~(layer2_outputs[3563]);
    assign layer3_outputs[4638] = layer2_outputs[4233];
    assign layer3_outputs[4639] = (layer2_outputs[737]) & (layer2_outputs[3627]);
    assign layer3_outputs[4640] = ~(layer2_outputs[0]) | (layer2_outputs[4984]);
    assign layer3_outputs[4641] = layer2_outputs[3887];
    assign layer3_outputs[4642] = layer2_outputs[1469];
    assign layer3_outputs[4643] = ~(layer2_outputs[4375]) | (layer2_outputs[3390]);
    assign layer3_outputs[4644] = ~((layer2_outputs[4446]) | (layer2_outputs[2955]));
    assign layer3_outputs[4645] = ~(layer2_outputs[5055]);
    assign layer3_outputs[4646] = ~(layer2_outputs[271]) | (layer2_outputs[4429]);
    assign layer3_outputs[4647] = (layer2_outputs[2139]) & ~(layer2_outputs[1297]);
    assign layer3_outputs[4648] = (layer2_outputs[3246]) & ~(layer2_outputs[3986]);
    assign layer3_outputs[4649] = 1'b1;
    assign layer3_outputs[4650] = (layer2_outputs[2991]) & ~(layer2_outputs[2146]);
    assign layer3_outputs[4651] = ~(layer2_outputs[3781]) | (layer2_outputs[3703]);
    assign layer3_outputs[4652] = layer2_outputs[1138];
    assign layer3_outputs[4653] = layer2_outputs[2801];
    assign layer3_outputs[4654] = ~(layer2_outputs[157]);
    assign layer3_outputs[4655] = ~((layer2_outputs[1311]) | (layer2_outputs[1019]));
    assign layer3_outputs[4656] = (layer2_outputs[5069]) ^ (layer2_outputs[1456]);
    assign layer3_outputs[4657] = (layer2_outputs[258]) ^ (layer2_outputs[2745]);
    assign layer3_outputs[4658] = (layer2_outputs[3723]) & ~(layer2_outputs[4618]);
    assign layer3_outputs[4659] = layer2_outputs[2983];
    assign layer3_outputs[4660] = ~(layer2_outputs[43]);
    assign layer3_outputs[4661] = ~(layer2_outputs[94]);
    assign layer3_outputs[4662] = ~(layer2_outputs[895]) | (layer2_outputs[3115]);
    assign layer3_outputs[4663] = layer2_outputs[4196];
    assign layer3_outputs[4664] = layer2_outputs[3214];
    assign layer3_outputs[4665] = ~((layer2_outputs[2924]) & (layer2_outputs[557]));
    assign layer3_outputs[4666] = ~(layer2_outputs[1260]) | (layer2_outputs[1010]);
    assign layer3_outputs[4667] = layer2_outputs[4799];
    assign layer3_outputs[4668] = ~(layer2_outputs[2772]);
    assign layer3_outputs[4669] = layer2_outputs[2424];
    assign layer3_outputs[4670] = ~(layer2_outputs[3080]);
    assign layer3_outputs[4671] = layer2_outputs[1541];
    assign layer3_outputs[4672] = 1'b1;
    assign layer3_outputs[4673] = (layer2_outputs[4534]) & (layer2_outputs[4379]);
    assign layer3_outputs[4674] = layer2_outputs[4147];
    assign layer3_outputs[4675] = (layer2_outputs[2886]) | (layer2_outputs[3939]);
    assign layer3_outputs[4676] = ~(layer2_outputs[935]);
    assign layer3_outputs[4677] = ~(layer2_outputs[375]) | (layer2_outputs[626]);
    assign layer3_outputs[4678] = ~(layer2_outputs[4314]) | (layer2_outputs[3073]);
    assign layer3_outputs[4679] = (layer2_outputs[2592]) & (layer2_outputs[4610]);
    assign layer3_outputs[4680] = layer2_outputs[3566];
    assign layer3_outputs[4681] = ~(layer2_outputs[575]);
    assign layer3_outputs[4682] = ~(layer2_outputs[2430]) | (layer2_outputs[3053]);
    assign layer3_outputs[4683] = layer2_outputs[3034];
    assign layer3_outputs[4684] = (layer2_outputs[1540]) | (layer2_outputs[1562]);
    assign layer3_outputs[4685] = ~(layer2_outputs[1654]);
    assign layer3_outputs[4686] = ~((layer2_outputs[3481]) & (layer2_outputs[4087]));
    assign layer3_outputs[4687] = 1'b1;
    assign layer3_outputs[4688] = ~(layer2_outputs[3136]) | (layer2_outputs[2223]);
    assign layer3_outputs[4689] = layer2_outputs[471];
    assign layer3_outputs[4690] = ~((layer2_outputs[1672]) & (layer2_outputs[4696]));
    assign layer3_outputs[4691] = layer2_outputs[4950];
    assign layer3_outputs[4692] = 1'b1;
    assign layer3_outputs[4693] = ~(layer2_outputs[1860]) | (layer2_outputs[1763]);
    assign layer3_outputs[4694] = ~(layer2_outputs[4674]);
    assign layer3_outputs[4695] = 1'b0;
    assign layer3_outputs[4696] = layer2_outputs[4325];
    assign layer3_outputs[4697] = (layer2_outputs[3841]) | (layer2_outputs[1088]);
    assign layer3_outputs[4698] = (layer2_outputs[1585]) | (layer2_outputs[5072]);
    assign layer3_outputs[4699] = layer2_outputs[3808];
    assign layer3_outputs[4700] = ~(layer2_outputs[79]) | (layer2_outputs[3238]);
    assign layer3_outputs[4701] = ~(layer2_outputs[3100]) | (layer2_outputs[4834]);
    assign layer3_outputs[4702] = ~(layer2_outputs[2236]) | (layer2_outputs[2657]);
    assign layer3_outputs[4703] = (layer2_outputs[2226]) | (layer2_outputs[703]);
    assign layer3_outputs[4704] = 1'b1;
    assign layer3_outputs[4705] = ~(layer2_outputs[3599]);
    assign layer3_outputs[4706] = 1'b1;
    assign layer3_outputs[4707] = ~(layer2_outputs[4040]);
    assign layer3_outputs[4708] = (layer2_outputs[3786]) & ~(layer2_outputs[306]);
    assign layer3_outputs[4709] = layer2_outputs[2823];
    assign layer3_outputs[4710] = ~(layer2_outputs[1997]);
    assign layer3_outputs[4711] = ~((layer2_outputs[653]) | (layer2_outputs[2434]));
    assign layer3_outputs[4712] = layer2_outputs[1211];
    assign layer3_outputs[4713] = 1'b0;
    assign layer3_outputs[4714] = layer2_outputs[1798];
    assign layer3_outputs[4715] = 1'b0;
    assign layer3_outputs[4716] = (layer2_outputs[1921]) & ~(layer2_outputs[2788]);
    assign layer3_outputs[4717] = (layer2_outputs[4914]) & ~(layer2_outputs[2196]);
    assign layer3_outputs[4718] = layer2_outputs[4723];
    assign layer3_outputs[4719] = 1'b1;
    assign layer3_outputs[4720] = layer2_outputs[3975];
    assign layer3_outputs[4721] = layer2_outputs[3922];
    assign layer3_outputs[4722] = 1'b0;
    assign layer3_outputs[4723] = 1'b0;
    assign layer3_outputs[4724] = ~(layer2_outputs[1259]) | (layer2_outputs[1375]);
    assign layer3_outputs[4725] = ~(layer2_outputs[2219]);
    assign layer3_outputs[4726] = (layer2_outputs[225]) & (layer2_outputs[685]);
    assign layer3_outputs[4727] = ~(layer2_outputs[2110]) | (layer2_outputs[2666]);
    assign layer3_outputs[4728] = ~((layer2_outputs[818]) | (layer2_outputs[2440]));
    assign layer3_outputs[4729] = 1'b0;
    assign layer3_outputs[4730] = (layer2_outputs[2140]) & ~(layer2_outputs[3574]);
    assign layer3_outputs[4731] = ~(layer2_outputs[92]) | (layer2_outputs[1536]);
    assign layer3_outputs[4732] = (layer2_outputs[3557]) & ~(layer2_outputs[4371]);
    assign layer3_outputs[4733] = (layer2_outputs[3887]) | (layer2_outputs[627]);
    assign layer3_outputs[4734] = ~(layer2_outputs[1459]);
    assign layer3_outputs[4735] = ~(layer2_outputs[2445]);
    assign layer3_outputs[4736] = ~(layer2_outputs[2435]) | (layer2_outputs[4028]);
    assign layer3_outputs[4737] = ~(layer2_outputs[5035]);
    assign layer3_outputs[4738] = ~(layer2_outputs[3074]) | (layer2_outputs[4623]);
    assign layer3_outputs[4739] = ~(layer2_outputs[480]);
    assign layer3_outputs[4740] = layer2_outputs[1140];
    assign layer3_outputs[4741] = ~(layer2_outputs[1600]) | (layer2_outputs[3391]);
    assign layer3_outputs[4742] = (layer2_outputs[4272]) & ~(layer2_outputs[1696]);
    assign layer3_outputs[4743] = (layer2_outputs[4424]) & ~(layer2_outputs[3856]);
    assign layer3_outputs[4744] = layer2_outputs[488];
    assign layer3_outputs[4745] = ~((layer2_outputs[3060]) | (layer2_outputs[1145]));
    assign layer3_outputs[4746] = layer2_outputs[2744];
    assign layer3_outputs[4747] = 1'b1;
    assign layer3_outputs[4748] = layer2_outputs[1858];
    assign layer3_outputs[4749] = (layer2_outputs[2927]) | (layer2_outputs[688]);
    assign layer3_outputs[4750] = ~(layer2_outputs[3754]);
    assign layer3_outputs[4751] = ~(layer2_outputs[1707]);
    assign layer3_outputs[4752] = (layer2_outputs[1371]) & ~(layer2_outputs[1140]);
    assign layer3_outputs[4753] = ~(layer2_outputs[3946]);
    assign layer3_outputs[4754] = ~((layer2_outputs[3556]) | (layer2_outputs[4792]));
    assign layer3_outputs[4755] = ~(layer2_outputs[4977]);
    assign layer3_outputs[4756] = ~(layer2_outputs[2079]);
    assign layer3_outputs[4757] = ~(layer2_outputs[3958]) | (layer2_outputs[2074]);
    assign layer3_outputs[4758] = layer2_outputs[5044];
    assign layer3_outputs[4759] = layer2_outputs[3267];
    assign layer3_outputs[4760] = layer2_outputs[3058];
    assign layer3_outputs[4761] = ~(layer2_outputs[67]) | (layer2_outputs[3489]);
    assign layer3_outputs[4762] = 1'b1;
    assign layer3_outputs[4763] = ~(layer2_outputs[318]);
    assign layer3_outputs[4764] = ~(layer2_outputs[4065]);
    assign layer3_outputs[4765] = (layer2_outputs[2727]) & ~(layer2_outputs[3006]);
    assign layer3_outputs[4766] = (layer2_outputs[2971]) ^ (layer2_outputs[2544]);
    assign layer3_outputs[4767] = (layer2_outputs[2113]) & (layer2_outputs[2534]);
    assign layer3_outputs[4768] = 1'b0;
    assign layer3_outputs[4769] = ~((layer2_outputs[3775]) | (layer2_outputs[2447]));
    assign layer3_outputs[4770] = ~(layer2_outputs[941]);
    assign layer3_outputs[4771] = ~(layer2_outputs[4606]);
    assign layer3_outputs[4772] = ~((layer2_outputs[2684]) | (layer2_outputs[3227]));
    assign layer3_outputs[4773] = 1'b0;
    assign layer3_outputs[4774] = 1'b1;
    assign layer3_outputs[4775] = ~(layer2_outputs[3111]);
    assign layer3_outputs[4776] = ~(layer2_outputs[3509]);
    assign layer3_outputs[4777] = ~(layer2_outputs[5025]) | (layer2_outputs[900]);
    assign layer3_outputs[4778] = layer2_outputs[2585];
    assign layer3_outputs[4779] = ~(layer2_outputs[2080]);
    assign layer3_outputs[4780] = ~(layer2_outputs[4194]);
    assign layer3_outputs[4781] = (layer2_outputs[4165]) & ~(layer2_outputs[4062]);
    assign layer3_outputs[4782] = 1'b0;
    assign layer3_outputs[4783] = ~(layer2_outputs[2016]);
    assign layer3_outputs[4784] = (layer2_outputs[1072]) & (layer2_outputs[1764]);
    assign layer3_outputs[4785] = 1'b0;
    assign layer3_outputs[4786] = ~(layer2_outputs[3408]) | (layer2_outputs[670]);
    assign layer3_outputs[4787] = ~(layer2_outputs[1040]) | (layer2_outputs[4591]);
    assign layer3_outputs[4788] = (layer2_outputs[1820]) & (layer2_outputs[625]);
    assign layer3_outputs[4789] = ~((layer2_outputs[407]) | (layer2_outputs[2041]));
    assign layer3_outputs[4790] = ~(layer2_outputs[154]) | (layer2_outputs[3438]);
    assign layer3_outputs[4791] = (layer2_outputs[3075]) & ~(layer2_outputs[629]);
    assign layer3_outputs[4792] = (layer2_outputs[4276]) & ~(layer2_outputs[590]);
    assign layer3_outputs[4793] = ~(layer2_outputs[204]);
    assign layer3_outputs[4794] = ~((layer2_outputs[1402]) | (layer2_outputs[3962]));
    assign layer3_outputs[4795] = ~(layer2_outputs[1584]) | (layer2_outputs[3981]);
    assign layer3_outputs[4796] = layer2_outputs[1492];
    assign layer3_outputs[4797] = 1'b1;
    assign layer3_outputs[4798] = ~(layer2_outputs[977]);
    assign layer3_outputs[4799] = layer2_outputs[2260];
    assign layer3_outputs[4800] = 1'b0;
    assign layer3_outputs[4801] = ~((layer2_outputs[1213]) | (layer2_outputs[2251]));
    assign layer3_outputs[4802] = 1'b0;
    assign layer3_outputs[4803] = 1'b0;
    assign layer3_outputs[4804] = ~(layer2_outputs[4811]);
    assign layer3_outputs[4805] = (layer2_outputs[2838]) ^ (layer2_outputs[1788]);
    assign layer3_outputs[4806] = layer2_outputs[2563];
    assign layer3_outputs[4807] = 1'b0;
    assign layer3_outputs[4808] = layer2_outputs[419];
    assign layer3_outputs[4809] = ~((layer2_outputs[1428]) & (layer2_outputs[1767]));
    assign layer3_outputs[4810] = ~(layer2_outputs[3127]);
    assign layer3_outputs[4811] = (layer2_outputs[2869]) & ~(layer2_outputs[4957]);
    assign layer3_outputs[4812] = (layer2_outputs[2610]) & ~(layer2_outputs[2717]);
    assign layer3_outputs[4813] = ~((layer2_outputs[4292]) & (layer2_outputs[449]));
    assign layer3_outputs[4814] = (layer2_outputs[2056]) ^ (layer2_outputs[4684]);
    assign layer3_outputs[4815] = ~(layer2_outputs[1223]);
    assign layer3_outputs[4816] = (layer2_outputs[322]) & (layer2_outputs[4777]);
    assign layer3_outputs[4817] = ~(layer2_outputs[3613]);
    assign layer3_outputs[4818] = 1'b0;
    assign layer3_outputs[4819] = ~(layer2_outputs[1823]);
    assign layer3_outputs[4820] = 1'b1;
    assign layer3_outputs[4821] = layer2_outputs[2269];
    assign layer3_outputs[4822] = ~(layer2_outputs[4996]);
    assign layer3_outputs[4823] = layer2_outputs[4801];
    assign layer3_outputs[4824] = (layer2_outputs[4865]) ^ (layer2_outputs[2416]);
    assign layer3_outputs[4825] = (layer2_outputs[569]) ^ (layer2_outputs[1936]);
    assign layer3_outputs[4826] = ~(layer2_outputs[5052]);
    assign layer3_outputs[4827] = (layer2_outputs[354]) & (layer2_outputs[4692]);
    assign layer3_outputs[4828] = ~(layer2_outputs[1976]) | (layer2_outputs[3765]);
    assign layer3_outputs[4829] = 1'b0;
    assign layer3_outputs[4830] = ~(layer2_outputs[1129]);
    assign layer3_outputs[4831] = layer2_outputs[606];
    assign layer3_outputs[4832] = ~(layer2_outputs[4920]);
    assign layer3_outputs[4833] = ~((layer2_outputs[4408]) & (layer2_outputs[419]));
    assign layer3_outputs[4834] = ~(layer2_outputs[124]);
    assign layer3_outputs[4835] = layer2_outputs[4916];
    assign layer3_outputs[4836] = ~((layer2_outputs[1458]) | (layer2_outputs[2693]));
    assign layer3_outputs[4837] = layer2_outputs[4937];
    assign layer3_outputs[4838] = 1'b0;
    assign layer3_outputs[4839] = layer2_outputs[118];
    assign layer3_outputs[4840] = (layer2_outputs[2704]) | (layer2_outputs[4137]);
    assign layer3_outputs[4841] = layer2_outputs[614];
    assign layer3_outputs[4842] = layer2_outputs[2932];
    assign layer3_outputs[4843] = ~(layer2_outputs[784]);
    assign layer3_outputs[4844] = layer2_outputs[3523];
    assign layer3_outputs[4845] = layer2_outputs[2205];
    assign layer3_outputs[4846] = ~(layer2_outputs[2622]) | (layer2_outputs[1621]);
    assign layer3_outputs[4847] = layer2_outputs[762];
    assign layer3_outputs[4848] = layer2_outputs[3606];
    assign layer3_outputs[4849] = (layer2_outputs[1902]) | (layer2_outputs[2551]);
    assign layer3_outputs[4850] = ~((layer2_outputs[1071]) | (layer2_outputs[1769]));
    assign layer3_outputs[4851] = ~(layer2_outputs[647]);
    assign layer3_outputs[4852] = ~(layer2_outputs[1553]) | (layer2_outputs[1613]);
    assign layer3_outputs[4853] = (layer2_outputs[411]) ^ (layer2_outputs[1005]);
    assign layer3_outputs[4854] = (layer2_outputs[4983]) ^ (layer2_outputs[4536]);
    assign layer3_outputs[4855] = (layer2_outputs[4115]) ^ (layer2_outputs[35]);
    assign layer3_outputs[4856] = 1'b1;
    assign layer3_outputs[4857] = 1'b1;
    assign layer3_outputs[4858] = (layer2_outputs[609]) & ~(layer2_outputs[803]);
    assign layer3_outputs[4859] = (layer2_outputs[2017]) | (layer2_outputs[1189]);
    assign layer3_outputs[4860] = (layer2_outputs[2740]) | (layer2_outputs[2743]);
    assign layer3_outputs[4861] = ~(layer2_outputs[3921]) | (layer2_outputs[3655]);
    assign layer3_outputs[4862] = 1'b1;
    assign layer3_outputs[4863] = ~(layer2_outputs[3897]);
    assign layer3_outputs[4864] = ~(layer2_outputs[773]);
    assign layer3_outputs[4865] = ~(layer2_outputs[860]);
    assign layer3_outputs[4866] = ~(layer2_outputs[4443]);
    assign layer3_outputs[4867] = layer2_outputs[4632];
    assign layer3_outputs[4868] = (layer2_outputs[1638]) & ~(layer2_outputs[641]);
    assign layer3_outputs[4869] = layer2_outputs[3414];
    assign layer3_outputs[4870] = (layer2_outputs[2956]) & ~(layer2_outputs[4904]);
    assign layer3_outputs[4871] = ~(layer2_outputs[5072]);
    assign layer3_outputs[4872] = ~(layer2_outputs[767]);
    assign layer3_outputs[4873] = 1'b0;
    assign layer3_outputs[4874] = ~(layer2_outputs[2675]);
    assign layer3_outputs[4875] = (layer2_outputs[5063]) ^ (layer2_outputs[3030]);
    assign layer3_outputs[4876] = (layer2_outputs[3497]) | (layer2_outputs[1206]);
    assign layer3_outputs[4877] = ~(layer2_outputs[3058]) | (layer2_outputs[256]);
    assign layer3_outputs[4878] = (layer2_outputs[2796]) & (layer2_outputs[4063]);
    assign layer3_outputs[4879] = (layer2_outputs[4271]) | (layer2_outputs[2537]);
    assign layer3_outputs[4880] = layer2_outputs[1544];
    assign layer3_outputs[4881] = layer2_outputs[4808];
    assign layer3_outputs[4882] = ~(layer2_outputs[2673]) | (layer2_outputs[2713]);
    assign layer3_outputs[4883] = (layer2_outputs[1063]) | (layer2_outputs[479]);
    assign layer3_outputs[4884] = ~((layer2_outputs[4949]) | (layer2_outputs[824]));
    assign layer3_outputs[4885] = layer2_outputs[576];
    assign layer3_outputs[4886] = layer2_outputs[4666];
    assign layer3_outputs[4887] = ~(layer2_outputs[885]) | (layer2_outputs[4041]);
    assign layer3_outputs[4888] = 1'b1;
    assign layer3_outputs[4889] = (layer2_outputs[1020]) & (layer2_outputs[1972]);
    assign layer3_outputs[4890] = 1'b0;
    assign layer3_outputs[4891] = layer2_outputs[799];
    assign layer3_outputs[4892] = layer2_outputs[254];
    assign layer3_outputs[4893] = layer2_outputs[1502];
    assign layer3_outputs[4894] = layer2_outputs[2302];
    assign layer3_outputs[4895] = ~(layer2_outputs[533]);
    assign layer3_outputs[4896] = ~(layer2_outputs[1452]);
    assign layer3_outputs[4897] = ~(layer2_outputs[2082]) | (layer2_outputs[3873]);
    assign layer3_outputs[4898] = ~((layer2_outputs[4404]) ^ (layer2_outputs[959]));
    assign layer3_outputs[4899] = ~(layer2_outputs[2488]);
    assign layer3_outputs[4900] = 1'b1;
    assign layer3_outputs[4901] = layer2_outputs[4213];
    assign layer3_outputs[4902] = ~((layer2_outputs[2217]) | (layer2_outputs[4726]));
    assign layer3_outputs[4903] = ~(layer2_outputs[1610]) | (layer2_outputs[2692]);
    assign layer3_outputs[4904] = layer2_outputs[1635];
    assign layer3_outputs[4905] = layer2_outputs[165];
    assign layer3_outputs[4906] = ~(layer2_outputs[4447]);
    assign layer3_outputs[4907] = 1'b0;
    assign layer3_outputs[4908] = ~((layer2_outputs[4605]) & (layer2_outputs[220]));
    assign layer3_outputs[4909] = (layer2_outputs[3840]) & (layer2_outputs[3013]);
    assign layer3_outputs[4910] = layer2_outputs[4627];
    assign layer3_outputs[4911] = (layer2_outputs[4700]) & ~(layer2_outputs[3483]);
    assign layer3_outputs[4912] = ~(layer2_outputs[3596]);
    assign layer3_outputs[4913] = (layer2_outputs[794]) & (layer2_outputs[2114]);
    assign layer3_outputs[4914] = (layer2_outputs[1916]) & ~(layer2_outputs[711]);
    assign layer3_outputs[4915] = ~(layer2_outputs[156]);
    assign layer3_outputs[4916] = ~(layer2_outputs[1029]);
    assign layer3_outputs[4917] = ~((layer2_outputs[4921]) & (layer2_outputs[1171]));
    assign layer3_outputs[4918] = (layer2_outputs[59]) ^ (layer2_outputs[339]);
    assign layer3_outputs[4919] = ~(layer2_outputs[801]);
    assign layer3_outputs[4920] = ~(layer2_outputs[2408]);
    assign layer3_outputs[4921] = ~(layer2_outputs[3012]) | (layer2_outputs[3305]);
    assign layer3_outputs[4922] = ~((layer2_outputs[2933]) | (layer2_outputs[1104]));
    assign layer3_outputs[4923] = (layer2_outputs[1565]) & ~(layer2_outputs[3486]);
    assign layer3_outputs[4924] = (layer2_outputs[3864]) & ~(layer2_outputs[2141]);
    assign layer3_outputs[4925] = ~((layer2_outputs[1130]) & (layer2_outputs[4104]));
    assign layer3_outputs[4926] = layer2_outputs[2180];
    assign layer3_outputs[4927] = ~((layer2_outputs[2111]) & (layer2_outputs[267]));
    assign layer3_outputs[4928] = ~(layer2_outputs[1002]) | (layer2_outputs[1012]);
    assign layer3_outputs[4929] = (layer2_outputs[496]) & (layer2_outputs[1490]);
    assign layer3_outputs[4930] = ~(layer2_outputs[4594]) | (layer2_outputs[4396]);
    assign layer3_outputs[4931] = (layer2_outputs[1643]) | (layer2_outputs[4827]);
    assign layer3_outputs[4932] = ~(layer2_outputs[1237]) | (layer2_outputs[2613]);
    assign layer3_outputs[4933] = ~(layer2_outputs[3915]) | (layer2_outputs[635]);
    assign layer3_outputs[4934] = 1'b1;
    assign layer3_outputs[4935] = (layer2_outputs[2691]) & (layer2_outputs[4833]);
    assign layer3_outputs[4936] = 1'b0;
    assign layer3_outputs[4937] = ~((layer2_outputs[371]) | (layer2_outputs[4268]));
    assign layer3_outputs[4938] = ~((layer2_outputs[909]) & (layer2_outputs[2014]));
    assign layer3_outputs[4939] = (layer2_outputs[3448]) & (layer2_outputs[625]);
    assign layer3_outputs[4940] = 1'b1;
    assign layer3_outputs[4941] = layer2_outputs[2483];
    assign layer3_outputs[4942] = ~((layer2_outputs[2449]) | (layer2_outputs[490]));
    assign layer3_outputs[4943] = 1'b1;
    assign layer3_outputs[4944] = layer2_outputs[64];
    assign layer3_outputs[4945] = ~((layer2_outputs[2689]) & (layer2_outputs[3746]));
    assign layer3_outputs[4946] = layer2_outputs[2363];
    assign layer3_outputs[4947] = (layer2_outputs[1495]) & ~(layer2_outputs[2716]);
    assign layer3_outputs[4948] = layer2_outputs[2896];
    assign layer3_outputs[4949] = ~(layer2_outputs[1309]) | (layer2_outputs[4713]);
    assign layer3_outputs[4950] = 1'b1;
    assign layer3_outputs[4951] = 1'b1;
    assign layer3_outputs[4952] = ~(layer2_outputs[639]);
    assign layer3_outputs[4953] = 1'b0;
    assign layer3_outputs[4954] = ~((layer2_outputs[1489]) & (layer2_outputs[2933]));
    assign layer3_outputs[4955] = ~(layer2_outputs[4503]);
    assign layer3_outputs[4956] = layer2_outputs[787];
    assign layer3_outputs[4957] = (layer2_outputs[52]) & ~(layer2_outputs[9]);
    assign layer3_outputs[4958] = ~(layer2_outputs[1043]) | (layer2_outputs[2292]);
    assign layer3_outputs[4959] = ~(layer2_outputs[370]) | (layer2_outputs[4934]);
    assign layer3_outputs[4960] = (layer2_outputs[774]) & ~(layer2_outputs[1523]);
    assign layer3_outputs[4961] = ~(layer2_outputs[4080]);
    assign layer3_outputs[4962] = ~(layer2_outputs[3593]);
    assign layer3_outputs[4963] = ~((layer2_outputs[632]) ^ (layer2_outputs[2247]));
    assign layer3_outputs[4964] = (layer2_outputs[4939]) | (layer2_outputs[3751]);
    assign layer3_outputs[4965] = ~(layer2_outputs[2014]) | (layer2_outputs[2547]);
    assign layer3_outputs[4966] = (layer2_outputs[5092]) & ~(layer2_outputs[1451]);
    assign layer3_outputs[4967] = ~(layer2_outputs[260]) | (layer2_outputs[2073]);
    assign layer3_outputs[4968] = (layer2_outputs[4399]) | (layer2_outputs[1307]);
    assign layer3_outputs[4969] = ~((layer2_outputs[4885]) | (layer2_outputs[1270]));
    assign layer3_outputs[4970] = layer2_outputs[2154];
    assign layer3_outputs[4971] = (layer2_outputs[4320]) & (layer2_outputs[3476]);
    assign layer3_outputs[4972] = (layer2_outputs[1920]) | (layer2_outputs[422]);
    assign layer3_outputs[4973] = 1'b1;
    assign layer3_outputs[4974] = ~((layer2_outputs[578]) & (layer2_outputs[2818]));
    assign layer3_outputs[4975] = layer2_outputs[1142];
    assign layer3_outputs[4976] = (layer2_outputs[755]) | (layer2_outputs[1576]);
    assign layer3_outputs[4977] = layer2_outputs[4308];
    assign layer3_outputs[4978] = ~(layer2_outputs[5032]) | (layer2_outputs[4798]);
    assign layer3_outputs[4979] = (layer2_outputs[3857]) & ~(layer2_outputs[4241]);
    assign layer3_outputs[4980] = ~((layer2_outputs[4025]) & (layer2_outputs[2441]));
    assign layer3_outputs[4981] = (layer2_outputs[2865]) & ~(layer2_outputs[2931]);
    assign layer3_outputs[4982] = ~(layer2_outputs[2234]);
    assign layer3_outputs[4983] = ~(layer2_outputs[179]);
    assign layer3_outputs[4984] = ~(layer2_outputs[4648]);
    assign layer3_outputs[4985] = ~((layer2_outputs[668]) & (layer2_outputs[4931]));
    assign layer3_outputs[4986] = (layer2_outputs[928]) & ~(layer2_outputs[4987]);
    assign layer3_outputs[4987] = layer2_outputs[3581];
    assign layer3_outputs[4988] = ~(layer2_outputs[4015]) | (layer2_outputs[2763]);
    assign layer3_outputs[4989] = ~(layer2_outputs[2127]) | (layer2_outputs[4311]);
    assign layer3_outputs[4990] = 1'b1;
    assign layer3_outputs[4991] = layer2_outputs[4595];
    assign layer3_outputs[4992] = ~(layer2_outputs[2990]);
    assign layer3_outputs[4993] = ~(layer2_outputs[1601]);
    assign layer3_outputs[4994] = layer2_outputs[3635];
    assign layer3_outputs[4995] = (layer2_outputs[3550]) & ~(layer2_outputs[589]);
    assign layer3_outputs[4996] = ~((layer2_outputs[1250]) & (layer2_outputs[571]));
    assign layer3_outputs[4997] = 1'b0;
    assign layer3_outputs[4998] = (layer2_outputs[141]) | (layer2_outputs[868]);
    assign layer3_outputs[4999] = (layer2_outputs[1525]) | (layer2_outputs[1792]);
    assign layer3_outputs[5000] = ~(layer2_outputs[1102]) | (layer2_outputs[4280]);
    assign layer3_outputs[5001] = ~(layer2_outputs[3927]) | (layer2_outputs[4462]);
    assign layer3_outputs[5002] = layer2_outputs[4531];
    assign layer3_outputs[5003] = ~(layer2_outputs[3719]);
    assign layer3_outputs[5004] = 1'b1;
    assign layer3_outputs[5005] = ~(layer2_outputs[2379]);
    assign layer3_outputs[5006] = 1'b1;
    assign layer3_outputs[5007] = layer2_outputs[4834];
    assign layer3_outputs[5008] = ~(layer2_outputs[2075]) | (layer2_outputs[2432]);
    assign layer3_outputs[5009] = layer2_outputs[4185];
    assign layer3_outputs[5010] = (layer2_outputs[1723]) | (layer2_outputs[4725]);
    assign layer3_outputs[5011] = ~(layer2_outputs[3299]);
    assign layer3_outputs[5012] = ~((layer2_outputs[684]) | (layer2_outputs[4740]));
    assign layer3_outputs[5013] = ~((layer2_outputs[2997]) | (layer2_outputs[1041]));
    assign layer3_outputs[5014] = ~(layer2_outputs[1834]);
    assign layer3_outputs[5015] = ~(layer2_outputs[4312]);
    assign layer3_outputs[5016] = ~(layer2_outputs[3637]) | (layer2_outputs[4717]);
    assign layer3_outputs[5017] = (layer2_outputs[2304]) | (layer2_outputs[424]);
    assign layer3_outputs[5018] = (layer2_outputs[4071]) & (layer2_outputs[3046]);
    assign layer3_outputs[5019] = ~(layer2_outputs[4086]);
    assign layer3_outputs[5020] = ~((layer2_outputs[2597]) & (layer2_outputs[1286]));
    assign layer3_outputs[5021] = ~(layer2_outputs[4646]);
    assign layer3_outputs[5022] = ~(layer2_outputs[4570]) | (layer2_outputs[8]);
    assign layer3_outputs[5023] = layer2_outputs[268];
    assign layer3_outputs[5024] = 1'b0;
    assign layer3_outputs[5025] = ~(layer2_outputs[1295]) | (layer2_outputs[325]);
    assign layer3_outputs[5026] = layer2_outputs[4469];
    assign layer3_outputs[5027] = 1'b0;
    assign layer3_outputs[5028] = 1'b0;
    assign layer3_outputs[5029] = ~(layer2_outputs[268]);
    assign layer3_outputs[5030] = layer2_outputs[732];
    assign layer3_outputs[5031] = ~(layer2_outputs[2086]);
    assign layer3_outputs[5032] = ~((layer2_outputs[4063]) & (layer2_outputs[2914]));
    assign layer3_outputs[5033] = (layer2_outputs[427]) & ~(layer2_outputs[543]);
    assign layer3_outputs[5034] = (layer2_outputs[1448]) & (layer2_outputs[4808]);
    assign layer3_outputs[5035] = 1'b0;
    assign layer3_outputs[5036] = (layer2_outputs[863]) & ~(layer2_outputs[745]);
    assign layer3_outputs[5037] = layer2_outputs[926];
    assign layer3_outputs[5038] = layer2_outputs[1092];
    assign layer3_outputs[5039] = (layer2_outputs[4604]) | (layer2_outputs[4506]);
    assign layer3_outputs[5040] = ~(layer2_outputs[4736]);
    assign layer3_outputs[5041] = ~(layer2_outputs[408]) | (layer2_outputs[3576]);
    assign layer3_outputs[5042] = 1'b0;
    assign layer3_outputs[5043] = (layer2_outputs[1966]) | (layer2_outputs[312]);
    assign layer3_outputs[5044] = (layer2_outputs[149]) & ~(layer2_outputs[3834]);
    assign layer3_outputs[5045] = 1'b1;
    assign layer3_outputs[5046] = (layer2_outputs[2953]) & ~(layer2_outputs[445]);
    assign layer3_outputs[5047] = ~(layer2_outputs[4097]);
    assign layer3_outputs[5048] = ~((layer2_outputs[822]) ^ (layer2_outputs[3794]));
    assign layer3_outputs[5049] = layer2_outputs[1851];
    assign layer3_outputs[5050] = ~(layer2_outputs[323]);
    assign layer3_outputs[5051] = 1'b1;
    assign layer3_outputs[5052] = (layer2_outputs[5090]) & ~(layer2_outputs[4817]);
    assign layer3_outputs[5053] = layer2_outputs[3878];
    assign layer3_outputs[5054] = ~((layer2_outputs[4969]) ^ (layer2_outputs[2660]));
    assign layer3_outputs[5055] = (layer2_outputs[3502]) & (layer2_outputs[522]);
    assign layer3_outputs[5056] = (layer2_outputs[4244]) & ~(layer2_outputs[1706]);
    assign layer3_outputs[5057] = layer2_outputs[853];
    assign layer3_outputs[5058] = layer2_outputs[3964];
    assign layer3_outputs[5059] = 1'b1;
    assign layer3_outputs[5060] = (layer2_outputs[174]) & ~(layer2_outputs[3474]);
    assign layer3_outputs[5061] = (layer2_outputs[4124]) & (layer2_outputs[1589]);
    assign layer3_outputs[5062] = ~(layer2_outputs[354]);
    assign layer3_outputs[5063] = ~(layer2_outputs[1007]) | (layer2_outputs[1352]);
    assign layer3_outputs[5064] = layer2_outputs[404];
    assign layer3_outputs[5065] = ~(layer2_outputs[4705]) | (layer2_outputs[2583]);
    assign layer3_outputs[5066] = 1'b1;
    assign layer3_outputs[5067] = ~(layer2_outputs[32]);
    assign layer3_outputs[5068] = (layer2_outputs[172]) & ~(layer2_outputs[3241]);
    assign layer3_outputs[5069] = ~(layer2_outputs[2161]) | (layer2_outputs[4166]);
    assign layer3_outputs[5070] = (layer2_outputs[782]) & (layer2_outputs[607]);
    assign layer3_outputs[5071] = (layer2_outputs[4651]) & ~(layer2_outputs[926]);
    assign layer3_outputs[5072] = (layer2_outputs[3711]) & (layer2_outputs[1246]);
    assign layer3_outputs[5073] = ~((layer2_outputs[4250]) & (layer2_outputs[3685]));
    assign layer3_outputs[5074] = (layer2_outputs[497]) & ~(layer2_outputs[4290]);
    assign layer3_outputs[5075] = (layer2_outputs[3667]) | (layer2_outputs[3358]);
    assign layer3_outputs[5076] = ~(layer2_outputs[278]);
    assign layer3_outputs[5077] = 1'b0;
    assign layer3_outputs[5078] = layer2_outputs[4963];
    assign layer3_outputs[5079] = ~(layer2_outputs[1431]);
    assign layer3_outputs[5080] = (layer2_outputs[5087]) ^ (layer2_outputs[72]);
    assign layer3_outputs[5081] = (layer2_outputs[2818]) & ~(layer2_outputs[1880]);
    assign layer3_outputs[5082] = ~(layer2_outputs[4206]) | (layer2_outputs[1956]);
    assign layer3_outputs[5083] = (layer2_outputs[367]) | (layer2_outputs[2294]);
    assign layer3_outputs[5084] = (layer2_outputs[736]) | (layer2_outputs[341]);
    assign layer3_outputs[5085] = 1'b0;
    assign layer3_outputs[5086] = (layer2_outputs[644]) ^ (layer2_outputs[3805]);
    assign layer3_outputs[5087] = layer2_outputs[951];
    assign layer3_outputs[5088] = ~(layer2_outputs[3089]);
    assign layer3_outputs[5089] = ~(layer2_outputs[3278]);
    assign layer3_outputs[5090] = (layer2_outputs[4039]) & ~(layer2_outputs[4037]);
    assign layer3_outputs[5091] = layer2_outputs[4911];
    assign layer3_outputs[5092] = ~(layer2_outputs[1487]);
    assign layer3_outputs[5093] = layer2_outputs[2903];
    assign layer3_outputs[5094] = layer2_outputs[4537];
    assign layer3_outputs[5095] = (layer2_outputs[608]) & ~(layer2_outputs[1930]);
    assign layer3_outputs[5096] = ~(layer2_outputs[3519]);
    assign layer3_outputs[5097] = ~(layer2_outputs[3866]) | (layer2_outputs[290]);
    assign layer3_outputs[5098] = (layer2_outputs[2946]) ^ (layer2_outputs[1339]);
    assign layer3_outputs[5099] = (layer2_outputs[3679]) & ~(layer2_outputs[1401]);
    assign layer3_outputs[5100] = layer2_outputs[2706];
    assign layer3_outputs[5101] = ~(layer2_outputs[3692]) | (layer2_outputs[3647]);
    assign layer3_outputs[5102] = 1'b0;
    assign layer3_outputs[5103] = layer2_outputs[4729];
    assign layer3_outputs[5104] = ~((layer2_outputs[1108]) ^ (layer2_outputs[5106]));
    assign layer3_outputs[5105] = ~((layer2_outputs[2234]) | (layer2_outputs[2841]));
    assign layer3_outputs[5106] = ~(layer2_outputs[2377]) | (layer2_outputs[4884]);
    assign layer3_outputs[5107] = 1'b1;
    assign layer3_outputs[5108] = ~(layer2_outputs[3818]) | (layer2_outputs[183]);
    assign layer3_outputs[5109] = (layer2_outputs[2610]) | (layer2_outputs[3176]);
    assign layer3_outputs[5110] = (layer2_outputs[4210]) ^ (layer2_outputs[2821]);
    assign layer3_outputs[5111] = (layer2_outputs[1227]) | (layer2_outputs[3071]);
    assign layer3_outputs[5112] = (layer2_outputs[2613]) & ~(layer2_outputs[3250]);
    assign layer3_outputs[5113] = 1'b1;
    assign layer3_outputs[5114] = 1'b1;
    assign layer3_outputs[5115] = ~(layer2_outputs[2997]);
    assign layer3_outputs[5116] = 1'b0;
    assign layer3_outputs[5117] = (layer2_outputs[3823]) | (layer2_outputs[2726]);
    assign layer3_outputs[5118] = (layer2_outputs[2023]) & ~(layer2_outputs[2098]);
    assign layer3_outputs[5119] = (layer2_outputs[4290]) & ~(layer2_outputs[74]);
    assign layer4_outputs[0] = ~((layer3_outputs[5094]) ^ (layer3_outputs[1659]));
    assign layer4_outputs[1] = 1'b0;
    assign layer4_outputs[2] = layer3_outputs[5037];
    assign layer4_outputs[3] = ~(layer3_outputs[2894]) | (layer3_outputs[727]);
    assign layer4_outputs[4] = ~((layer3_outputs[898]) | (layer3_outputs[3178]));
    assign layer4_outputs[5] = layer3_outputs[218];
    assign layer4_outputs[6] = ~(layer3_outputs[4568]) | (layer3_outputs[2858]);
    assign layer4_outputs[7] = layer3_outputs[1474];
    assign layer4_outputs[8] = ~(layer3_outputs[4667]);
    assign layer4_outputs[9] = ~(layer3_outputs[1331]);
    assign layer4_outputs[10] = layer3_outputs[2279];
    assign layer4_outputs[11] = layer3_outputs[4341];
    assign layer4_outputs[12] = layer3_outputs[5057];
    assign layer4_outputs[13] = ~(layer3_outputs[1362]);
    assign layer4_outputs[14] = layer3_outputs[2386];
    assign layer4_outputs[15] = ~((layer3_outputs[1220]) | (layer3_outputs[3316]));
    assign layer4_outputs[16] = (layer3_outputs[3416]) & ~(layer3_outputs[4103]);
    assign layer4_outputs[17] = ~(layer3_outputs[2661]);
    assign layer4_outputs[18] = layer3_outputs[4678];
    assign layer4_outputs[19] = ~(layer3_outputs[2213]);
    assign layer4_outputs[20] = (layer3_outputs[2009]) | (layer3_outputs[410]);
    assign layer4_outputs[21] = layer3_outputs[4584];
    assign layer4_outputs[22] = layer3_outputs[3857];
    assign layer4_outputs[23] = layer3_outputs[2290];
    assign layer4_outputs[24] = 1'b1;
    assign layer4_outputs[25] = layer3_outputs[2438];
    assign layer4_outputs[26] = ~(layer3_outputs[4202]);
    assign layer4_outputs[27] = (layer3_outputs[366]) & ~(layer3_outputs[199]);
    assign layer4_outputs[28] = (layer3_outputs[4877]) ^ (layer3_outputs[575]);
    assign layer4_outputs[29] = ~(layer3_outputs[4181]);
    assign layer4_outputs[30] = layer3_outputs[3551];
    assign layer4_outputs[31] = ~(layer3_outputs[4444]);
    assign layer4_outputs[32] = ~(layer3_outputs[3735]);
    assign layer4_outputs[33] = ~(layer3_outputs[2903]) | (layer3_outputs[4658]);
    assign layer4_outputs[34] = ~(layer3_outputs[1582]) | (layer3_outputs[3447]);
    assign layer4_outputs[35] = 1'b0;
    assign layer4_outputs[36] = 1'b1;
    assign layer4_outputs[37] = 1'b1;
    assign layer4_outputs[38] = (layer3_outputs[4231]) & ~(layer3_outputs[4769]);
    assign layer4_outputs[39] = 1'b1;
    assign layer4_outputs[40] = layer3_outputs[1027];
    assign layer4_outputs[41] = (layer3_outputs[3907]) | (layer3_outputs[4321]);
    assign layer4_outputs[42] = ~(layer3_outputs[3306]);
    assign layer4_outputs[43] = ~(layer3_outputs[1862]);
    assign layer4_outputs[44] = (layer3_outputs[529]) & ~(layer3_outputs[1066]);
    assign layer4_outputs[45] = layer3_outputs[2126];
    assign layer4_outputs[46] = 1'b0;
    assign layer4_outputs[47] = ~((layer3_outputs[1260]) | (layer3_outputs[1709]));
    assign layer4_outputs[48] = layer3_outputs[4367];
    assign layer4_outputs[49] = 1'b1;
    assign layer4_outputs[50] = layer3_outputs[1560];
    assign layer4_outputs[51] = 1'b0;
    assign layer4_outputs[52] = (layer3_outputs[1861]) & (layer3_outputs[2143]);
    assign layer4_outputs[53] = layer3_outputs[2264];
    assign layer4_outputs[54] = (layer3_outputs[4705]) & (layer3_outputs[1250]);
    assign layer4_outputs[55] = layer3_outputs[4626];
    assign layer4_outputs[56] = 1'b1;
    assign layer4_outputs[57] = ~(layer3_outputs[2304]);
    assign layer4_outputs[58] = (layer3_outputs[1798]) & (layer3_outputs[5014]);
    assign layer4_outputs[59] = (layer3_outputs[4901]) | (layer3_outputs[3938]);
    assign layer4_outputs[60] = ~(layer3_outputs[309]);
    assign layer4_outputs[61] = ~(layer3_outputs[3508]);
    assign layer4_outputs[62] = (layer3_outputs[4203]) & ~(layer3_outputs[4998]);
    assign layer4_outputs[63] = ~(layer3_outputs[5017]) | (layer3_outputs[1793]);
    assign layer4_outputs[64] = 1'b1;
    assign layer4_outputs[65] = ~(layer3_outputs[3598]) | (layer3_outputs[2623]);
    assign layer4_outputs[66] = ~((layer3_outputs[4120]) | (layer3_outputs[3647]));
    assign layer4_outputs[67] = ~(layer3_outputs[937]) | (layer3_outputs[4218]);
    assign layer4_outputs[68] = 1'b1;
    assign layer4_outputs[69] = layer3_outputs[3676];
    assign layer4_outputs[70] = (layer3_outputs[2928]) & (layer3_outputs[1540]);
    assign layer4_outputs[71] = (layer3_outputs[1497]) & ~(layer3_outputs[2655]);
    assign layer4_outputs[72] = ~(layer3_outputs[3343]) | (layer3_outputs[4514]);
    assign layer4_outputs[73] = ~(layer3_outputs[4406]);
    assign layer4_outputs[74] = ~(layer3_outputs[3428]) | (layer3_outputs[2215]);
    assign layer4_outputs[75] = 1'b0;
    assign layer4_outputs[76] = (layer3_outputs[2704]) ^ (layer3_outputs[1286]);
    assign layer4_outputs[77] = (layer3_outputs[4058]) ^ (layer3_outputs[2266]);
    assign layer4_outputs[78] = (layer3_outputs[4671]) | (layer3_outputs[3334]);
    assign layer4_outputs[79] = 1'b0;
    assign layer4_outputs[80] = ~((layer3_outputs[4197]) | (layer3_outputs[3201]));
    assign layer4_outputs[81] = 1'b0;
    assign layer4_outputs[82] = ~((layer3_outputs[3471]) ^ (layer3_outputs[257]));
    assign layer4_outputs[83] = 1'b1;
    assign layer4_outputs[84] = (layer3_outputs[380]) ^ (layer3_outputs[1229]);
    assign layer4_outputs[85] = layer3_outputs[3415];
    assign layer4_outputs[86] = 1'b1;
    assign layer4_outputs[87] = (layer3_outputs[2693]) | (layer3_outputs[1642]);
    assign layer4_outputs[88] = ~(layer3_outputs[2525]);
    assign layer4_outputs[89] = 1'b1;
    assign layer4_outputs[90] = ~(layer3_outputs[1333]);
    assign layer4_outputs[91] = ~(layer3_outputs[820]);
    assign layer4_outputs[92] = ~(layer3_outputs[3911]);
    assign layer4_outputs[93] = layer3_outputs[3591];
    assign layer4_outputs[94] = (layer3_outputs[3369]) & (layer3_outputs[3995]);
    assign layer4_outputs[95] = ~(layer3_outputs[4694]);
    assign layer4_outputs[96] = layer3_outputs[4175];
    assign layer4_outputs[97] = (layer3_outputs[4927]) & ~(layer3_outputs[3188]);
    assign layer4_outputs[98] = layer3_outputs[4952];
    assign layer4_outputs[99] = layer3_outputs[1833];
    assign layer4_outputs[100] = (layer3_outputs[1846]) & ~(layer3_outputs[3417]);
    assign layer4_outputs[101] = layer3_outputs[1827];
    assign layer4_outputs[102] = layer3_outputs[4873];
    assign layer4_outputs[103] = (layer3_outputs[1689]) & ~(layer3_outputs[2151]);
    assign layer4_outputs[104] = layer3_outputs[3457];
    assign layer4_outputs[105] = (layer3_outputs[2589]) & ~(layer3_outputs[5042]);
    assign layer4_outputs[106] = ~(layer3_outputs[2920]) | (layer3_outputs[964]);
    assign layer4_outputs[107] = layer3_outputs[5001];
    assign layer4_outputs[108] = layer3_outputs[4346];
    assign layer4_outputs[109] = (layer3_outputs[1461]) & (layer3_outputs[3007]);
    assign layer4_outputs[110] = ~((layer3_outputs[934]) ^ (layer3_outputs[2176]));
    assign layer4_outputs[111] = layer3_outputs[1254];
    assign layer4_outputs[112] = layer3_outputs[2610];
    assign layer4_outputs[113] = ~(layer3_outputs[3139]);
    assign layer4_outputs[114] = 1'b0;
    assign layer4_outputs[115] = ~(layer3_outputs[4444]) | (layer3_outputs[4787]);
    assign layer4_outputs[116] = ~(layer3_outputs[432]) | (layer3_outputs[1651]);
    assign layer4_outputs[117] = ~(layer3_outputs[4658]);
    assign layer4_outputs[118] = layer3_outputs[2230];
    assign layer4_outputs[119] = ~((layer3_outputs[603]) ^ (layer3_outputs[3354]));
    assign layer4_outputs[120] = layer3_outputs[3727];
    assign layer4_outputs[121] = layer3_outputs[424];
    assign layer4_outputs[122] = (layer3_outputs[2300]) ^ (layer3_outputs[1452]);
    assign layer4_outputs[123] = 1'b1;
    assign layer4_outputs[124] = ~(layer3_outputs[4412]);
    assign layer4_outputs[125] = ~((layer3_outputs[2981]) | (layer3_outputs[4721]));
    assign layer4_outputs[126] = ~(layer3_outputs[195]) | (layer3_outputs[4689]);
    assign layer4_outputs[127] = ~((layer3_outputs[2436]) | (layer3_outputs[2160]));
    assign layer4_outputs[128] = (layer3_outputs[3213]) ^ (layer3_outputs[3207]);
    assign layer4_outputs[129] = ~(layer3_outputs[1420]) | (layer3_outputs[3307]);
    assign layer4_outputs[130] = ~(layer3_outputs[2735]);
    assign layer4_outputs[131] = layer3_outputs[884];
    assign layer4_outputs[132] = ~(layer3_outputs[4337]);
    assign layer4_outputs[133] = ~(layer3_outputs[1818]);
    assign layer4_outputs[134] = layer3_outputs[1767];
    assign layer4_outputs[135] = ~(layer3_outputs[79]);
    assign layer4_outputs[136] = 1'b0;
    assign layer4_outputs[137] = 1'b1;
    assign layer4_outputs[138] = ~((layer3_outputs[1305]) & (layer3_outputs[3854]));
    assign layer4_outputs[139] = ~(layer3_outputs[3670]) | (layer3_outputs[1061]);
    assign layer4_outputs[140] = ~(layer3_outputs[4596]) | (layer3_outputs[3506]);
    assign layer4_outputs[141] = ~(layer3_outputs[1836]);
    assign layer4_outputs[142] = (layer3_outputs[2071]) | (layer3_outputs[967]);
    assign layer4_outputs[143] = (layer3_outputs[4107]) & ~(layer3_outputs[2661]);
    assign layer4_outputs[144] = ~((layer3_outputs[3344]) | (layer3_outputs[4799]));
    assign layer4_outputs[145] = layer3_outputs[3892];
    assign layer4_outputs[146] = ~(layer3_outputs[2391]);
    assign layer4_outputs[147] = (layer3_outputs[2629]) ^ (layer3_outputs[1217]);
    assign layer4_outputs[148] = (layer3_outputs[3423]) & (layer3_outputs[4507]);
    assign layer4_outputs[149] = (layer3_outputs[4907]) & ~(layer3_outputs[766]);
    assign layer4_outputs[150] = layer3_outputs[237];
    assign layer4_outputs[151] = layer3_outputs[3025];
    assign layer4_outputs[152] = ~(layer3_outputs[4232]);
    assign layer4_outputs[153] = (layer3_outputs[4342]) & ~(layer3_outputs[3147]);
    assign layer4_outputs[154] = ~(layer3_outputs[2555]);
    assign layer4_outputs[155] = 1'b0;
    assign layer4_outputs[156] = (layer3_outputs[1199]) & ~(layer3_outputs[4802]);
    assign layer4_outputs[157] = ~((layer3_outputs[2613]) ^ (layer3_outputs[2265]));
    assign layer4_outputs[158] = layer3_outputs[215];
    assign layer4_outputs[159] = (layer3_outputs[3972]) & ~(layer3_outputs[234]);
    assign layer4_outputs[160] = ~(layer3_outputs[467]);
    assign layer4_outputs[161] = (layer3_outputs[4899]) | (layer3_outputs[1541]);
    assign layer4_outputs[162] = layer3_outputs[3537];
    assign layer4_outputs[163] = layer3_outputs[5111];
    assign layer4_outputs[164] = 1'b0;
    assign layer4_outputs[165] = layer3_outputs[3953];
    assign layer4_outputs[166] = layer3_outputs[4428];
    assign layer4_outputs[167] = ~(layer3_outputs[1693]) | (layer3_outputs[1738]);
    assign layer4_outputs[168] = ~(layer3_outputs[2878]) | (layer3_outputs[1151]);
    assign layer4_outputs[169] = ~((layer3_outputs[1963]) & (layer3_outputs[2730]));
    assign layer4_outputs[170] = ~(layer3_outputs[128]);
    assign layer4_outputs[171] = ~(layer3_outputs[4367]) | (layer3_outputs[3824]);
    assign layer4_outputs[172] = (layer3_outputs[3559]) & ~(layer3_outputs[2305]);
    assign layer4_outputs[173] = layer3_outputs[433];
    assign layer4_outputs[174] = ~((layer3_outputs[4662]) & (layer3_outputs[2446]));
    assign layer4_outputs[175] = (layer3_outputs[700]) | (layer3_outputs[1020]);
    assign layer4_outputs[176] = layer3_outputs[4177];
    assign layer4_outputs[177] = ~(layer3_outputs[3070]) | (layer3_outputs[1852]);
    assign layer4_outputs[178] = (layer3_outputs[2772]) & ~(layer3_outputs[252]);
    assign layer4_outputs[179] = ~(layer3_outputs[102]);
    assign layer4_outputs[180] = ~((layer3_outputs[3089]) & (layer3_outputs[3725]));
    assign layer4_outputs[181] = layer3_outputs[2750];
    assign layer4_outputs[182] = 1'b0;
    assign layer4_outputs[183] = 1'b1;
    assign layer4_outputs[184] = layer3_outputs[1801];
    assign layer4_outputs[185] = (layer3_outputs[3251]) & (layer3_outputs[79]);
    assign layer4_outputs[186] = ~(layer3_outputs[5003]);
    assign layer4_outputs[187] = ~(layer3_outputs[1209]);
    assign layer4_outputs[188] = ~((layer3_outputs[938]) & (layer3_outputs[2745]));
    assign layer4_outputs[189] = ~(layer3_outputs[2554]) | (layer3_outputs[2989]);
    assign layer4_outputs[190] = (layer3_outputs[2050]) ^ (layer3_outputs[2537]);
    assign layer4_outputs[191] = (layer3_outputs[1919]) & ~(layer3_outputs[484]);
    assign layer4_outputs[192] = ~(layer3_outputs[4357]) | (layer3_outputs[2100]);
    assign layer4_outputs[193] = ~(layer3_outputs[679]);
    assign layer4_outputs[194] = 1'b1;
    assign layer4_outputs[195] = (layer3_outputs[1720]) ^ (layer3_outputs[1530]);
    assign layer4_outputs[196] = (layer3_outputs[1893]) ^ (layer3_outputs[5098]);
    assign layer4_outputs[197] = ~(layer3_outputs[3574]);
    assign layer4_outputs[198] = (layer3_outputs[3574]) & (layer3_outputs[3971]);
    assign layer4_outputs[199] = ~(layer3_outputs[3878]);
    assign layer4_outputs[200] = 1'b1;
    assign layer4_outputs[201] = (layer3_outputs[2640]) ^ (layer3_outputs[1615]);
    assign layer4_outputs[202] = ~(layer3_outputs[4005]);
    assign layer4_outputs[203] = (layer3_outputs[4768]) & ~(layer3_outputs[4787]);
    assign layer4_outputs[204] = ~((layer3_outputs[3445]) | (layer3_outputs[3849]));
    assign layer4_outputs[205] = ~((layer3_outputs[2424]) | (layer3_outputs[673]));
    assign layer4_outputs[206] = ~(layer3_outputs[4914]);
    assign layer4_outputs[207] = layer3_outputs[3701];
    assign layer4_outputs[208] = (layer3_outputs[3202]) & ~(layer3_outputs[4840]);
    assign layer4_outputs[209] = 1'b1;
    assign layer4_outputs[210] = ~(layer3_outputs[3998]) | (layer3_outputs[648]);
    assign layer4_outputs[211] = ~(layer3_outputs[3941]);
    assign layer4_outputs[212] = ~((layer3_outputs[1851]) | (layer3_outputs[4432]));
    assign layer4_outputs[213] = ~(layer3_outputs[2542]);
    assign layer4_outputs[214] = ~(layer3_outputs[4384]);
    assign layer4_outputs[215] = (layer3_outputs[236]) & ~(layer3_outputs[5008]);
    assign layer4_outputs[216] = ~(layer3_outputs[1118]);
    assign layer4_outputs[217] = (layer3_outputs[4203]) | (layer3_outputs[1993]);
    assign layer4_outputs[218] = 1'b0;
    assign layer4_outputs[219] = ~((layer3_outputs[683]) & (layer3_outputs[2943]));
    assign layer4_outputs[220] = (layer3_outputs[1644]) & (layer3_outputs[4828]);
    assign layer4_outputs[221] = ~((layer3_outputs[3346]) & (layer3_outputs[750]));
    assign layer4_outputs[222] = ~(layer3_outputs[3355]);
    assign layer4_outputs[223] = ~(layer3_outputs[2808]);
    assign layer4_outputs[224] = (layer3_outputs[4566]) & (layer3_outputs[3516]);
    assign layer4_outputs[225] = (layer3_outputs[828]) & ~(layer3_outputs[444]);
    assign layer4_outputs[226] = layer3_outputs[2419];
    assign layer4_outputs[227] = ~((layer3_outputs[2807]) & (layer3_outputs[1487]));
    assign layer4_outputs[228] = ~(layer3_outputs[4505]);
    assign layer4_outputs[229] = ~(layer3_outputs[2620]);
    assign layer4_outputs[230] = ~((layer3_outputs[1061]) ^ (layer3_outputs[2448]));
    assign layer4_outputs[231] = layer3_outputs[1608];
    assign layer4_outputs[232] = (layer3_outputs[2461]) & (layer3_outputs[655]);
    assign layer4_outputs[233] = ~(layer3_outputs[186]);
    assign layer4_outputs[234] = ~(layer3_outputs[668]);
    assign layer4_outputs[235] = ~((layer3_outputs[3668]) | (layer3_outputs[972]));
    assign layer4_outputs[236] = layer3_outputs[3076];
    assign layer4_outputs[237] = ~(layer3_outputs[3249]);
    assign layer4_outputs[238] = layer3_outputs[180];
    assign layer4_outputs[239] = ~((layer3_outputs[470]) | (layer3_outputs[1528]));
    assign layer4_outputs[240] = (layer3_outputs[1988]) & ~(layer3_outputs[2488]);
    assign layer4_outputs[241] = ~(layer3_outputs[2777]) | (layer3_outputs[1390]);
    assign layer4_outputs[242] = ~(layer3_outputs[3472]);
    assign layer4_outputs[243] = ~(layer3_outputs[2612]);
    assign layer4_outputs[244] = ~(layer3_outputs[3506]);
    assign layer4_outputs[245] = ~(layer3_outputs[1614]);
    assign layer4_outputs[246] = (layer3_outputs[3501]) & (layer3_outputs[3441]);
    assign layer4_outputs[247] = ~(layer3_outputs[102]);
    assign layer4_outputs[248] = ~((layer3_outputs[4026]) & (layer3_outputs[1336]));
    assign layer4_outputs[249] = ~(layer3_outputs[4234]) | (layer3_outputs[2619]);
    assign layer4_outputs[250] = ~(layer3_outputs[1712]);
    assign layer4_outputs[251] = ~(layer3_outputs[496]);
    assign layer4_outputs[252] = ~(layer3_outputs[3192]);
    assign layer4_outputs[253] = (layer3_outputs[201]) ^ (layer3_outputs[3929]);
    assign layer4_outputs[254] = layer3_outputs[3319];
    assign layer4_outputs[255] = ~(layer3_outputs[1164]);
    assign layer4_outputs[256] = (layer3_outputs[4791]) & ~(layer3_outputs[2301]);
    assign layer4_outputs[257] = ~(layer3_outputs[3380]);
    assign layer4_outputs[258] = (layer3_outputs[1598]) | (layer3_outputs[1182]);
    assign layer4_outputs[259] = ~(layer3_outputs[3399]);
    assign layer4_outputs[260] = ~(layer3_outputs[3030]);
    assign layer4_outputs[261] = ~(layer3_outputs[4413]);
    assign layer4_outputs[262] = (layer3_outputs[2678]) | (layer3_outputs[54]);
    assign layer4_outputs[263] = (layer3_outputs[3898]) ^ (layer3_outputs[1617]);
    assign layer4_outputs[264] = ~(layer3_outputs[4369]);
    assign layer4_outputs[265] = ~((layer3_outputs[4372]) | (layer3_outputs[2306]));
    assign layer4_outputs[266] = (layer3_outputs[3507]) | (layer3_outputs[4844]);
    assign layer4_outputs[267] = ~(layer3_outputs[3244]);
    assign layer4_outputs[268] = (layer3_outputs[2517]) | (layer3_outputs[242]);
    assign layer4_outputs[269] = (layer3_outputs[2530]) & (layer3_outputs[341]);
    assign layer4_outputs[270] = layer3_outputs[3464];
    assign layer4_outputs[271] = layer3_outputs[2464];
    assign layer4_outputs[272] = (layer3_outputs[969]) & ~(layer3_outputs[661]);
    assign layer4_outputs[273] = (layer3_outputs[3888]) ^ (layer3_outputs[3897]);
    assign layer4_outputs[274] = ~(layer3_outputs[1011]) | (layer3_outputs[20]);
    assign layer4_outputs[275] = layer3_outputs[1934];
    assign layer4_outputs[276] = ~(layer3_outputs[3481]);
    assign layer4_outputs[277] = ~(layer3_outputs[561]);
    assign layer4_outputs[278] = (layer3_outputs[1531]) & (layer3_outputs[1858]);
    assign layer4_outputs[279] = (layer3_outputs[394]) | (layer3_outputs[3760]);
    assign layer4_outputs[280] = ~((layer3_outputs[4221]) ^ (layer3_outputs[58]));
    assign layer4_outputs[281] = layer3_outputs[5070];
    assign layer4_outputs[282] = (layer3_outputs[2479]) & ~(layer3_outputs[3341]);
    assign layer4_outputs[283] = layer3_outputs[5099];
    assign layer4_outputs[284] = (layer3_outputs[1496]) & ~(layer3_outputs[2813]);
    assign layer4_outputs[285] = ~(layer3_outputs[3181]);
    assign layer4_outputs[286] = layer3_outputs[4132];
    assign layer4_outputs[287] = ~((layer3_outputs[3368]) ^ (layer3_outputs[4594]));
    assign layer4_outputs[288] = ~(layer3_outputs[4850]) | (layer3_outputs[1321]);
    assign layer4_outputs[289] = layer3_outputs[801];
    assign layer4_outputs[290] = layer3_outputs[1590];
    assign layer4_outputs[291] = ~((layer3_outputs[2520]) | (layer3_outputs[761]));
    assign layer4_outputs[292] = (layer3_outputs[1071]) & ~(layer3_outputs[468]);
    assign layer4_outputs[293] = (layer3_outputs[2104]) ^ (layer3_outputs[4729]);
    assign layer4_outputs[294] = 1'b0;
    assign layer4_outputs[295] = (layer3_outputs[2494]) ^ (layer3_outputs[3988]);
    assign layer4_outputs[296] = (layer3_outputs[491]) ^ (layer3_outputs[4108]);
    assign layer4_outputs[297] = layer3_outputs[2925];
    assign layer4_outputs[298] = ~((layer3_outputs[1223]) | (layer3_outputs[3252]));
    assign layer4_outputs[299] = layer3_outputs[1386];
    assign layer4_outputs[300] = (layer3_outputs[1658]) & ~(layer3_outputs[5085]);
    assign layer4_outputs[301] = ~(layer3_outputs[1116]);
    assign layer4_outputs[302] = ~(layer3_outputs[3650]);
    assign layer4_outputs[303] = ~((layer3_outputs[2792]) & (layer3_outputs[2952]));
    assign layer4_outputs[304] = layer3_outputs[1889];
    assign layer4_outputs[305] = ~(layer3_outputs[2817]);
    assign layer4_outputs[306] = layer3_outputs[965];
    assign layer4_outputs[307] = (layer3_outputs[1147]) & (layer3_outputs[3338]);
    assign layer4_outputs[308] = layer3_outputs[1352];
    assign layer4_outputs[309] = ~(layer3_outputs[1861]);
    assign layer4_outputs[310] = (layer3_outputs[1170]) ^ (layer3_outputs[329]);
    assign layer4_outputs[311] = ~((layer3_outputs[3096]) | (layer3_outputs[2516]));
    assign layer4_outputs[312] = ~(layer3_outputs[1869]);
    assign layer4_outputs[313] = (layer3_outputs[556]) ^ (layer3_outputs[3190]);
    assign layer4_outputs[314] = (layer3_outputs[3546]) | (layer3_outputs[1264]);
    assign layer4_outputs[315] = (layer3_outputs[4263]) | (layer3_outputs[4206]);
    assign layer4_outputs[316] = (layer3_outputs[2596]) & ~(layer3_outputs[3267]);
    assign layer4_outputs[317] = ~(layer3_outputs[3355]);
    assign layer4_outputs[318] = (layer3_outputs[4240]) ^ (layer3_outputs[227]);
    assign layer4_outputs[319] = ~(layer3_outputs[4429]) | (layer3_outputs[4205]);
    assign layer4_outputs[320] = ~((layer3_outputs[3086]) ^ (layer3_outputs[3999]));
    assign layer4_outputs[321] = layer3_outputs[858];
    assign layer4_outputs[322] = (layer3_outputs[3751]) & (layer3_outputs[3450]);
    assign layer4_outputs[323] = ~(layer3_outputs[3542]) | (layer3_outputs[2927]);
    assign layer4_outputs[324] = 1'b1;
    assign layer4_outputs[325] = ~(layer3_outputs[2356]) | (layer3_outputs[320]);
    assign layer4_outputs[326] = ~(layer3_outputs[3716]);
    assign layer4_outputs[327] = ~(layer3_outputs[2795]) | (layer3_outputs[3434]);
    assign layer4_outputs[328] = ~(layer3_outputs[61]);
    assign layer4_outputs[329] = ~(layer3_outputs[3265]);
    assign layer4_outputs[330] = ~(layer3_outputs[4189]) | (layer3_outputs[1451]);
    assign layer4_outputs[331] = ~(layer3_outputs[2487]);
    assign layer4_outputs[332] = layer3_outputs[3460];
    assign layer4_outputs[333] = layer3_outputs[1262];
    assign layer4_outputs[334] = (layer3_outputs[1478]) & ~(layer3_outputs[3352]);
    assign layer4_outputs[335] = layer3_outputs[3469];
    assign layer4_outputs[336] = ~(layer3_outputs[327]);
    assign layer4_outputs[337] = layer3_outputs[752];
    assign layer4_outputs[338] = ~(layer3_outputs[1225]) | (layer3_outputs[4597]);
    assign layer4_outputs[339] = ~((layer3_outputs[2550]) & (layer3_outputs[877]));
    assign layer4_outputs[340] = layer3_outputs[5099];
    assign layer4_outputs[341] = ~(layer3_outputs[2246]) | (layer3_outputs[2674]);
    assign layer4_outputs[342] = (layer3_outputs[1735]) ^ (layer3_outputs[2074]);
    assign layer4_outputs[343] = ~((layer3_outputs[1270]) & (layer3_outputs[3914]));
    assign layer4_outputs[344] = (layer3_outputs[2977]) & (layer3_outputs[342]);
    assign layer4_outputs[345] = layer3_outputs[3230];
    assign layer4_outputs[346] = ~((layer3_outputs[407]) | (layer3_outputs[2157]));
    assign layer4_outputs[347] = ~((layer3_outputs[1071]) & (layer3_outputs[2988]));
    assign layer4_outputs[348] = (layer3_outputs[910]) | (layer3_outputs[4950]);
    assign layer4_outputs[349] = ~(layer3_outputs[1208]);
    assign layer4_outputs[350] = (layer3_outputs[4221]) | (layer3_outputs[1424]);
    assign layer4_outputs[351] = layer3_outputs[3923];
    assign layer4_outputs[352] = 1'b0;
    assign layer4_outputs[353] = (layer3_outputs[1878]) | (layer3_outputs[399]);
    assign layer4_outputs[354] = ~((layer3_outputs[3262]) | (layer3_outputs[4653]));
    assign layer4_outputs[355] = ~(layer3_outputs[433]) | (layer3_outputs[1478]);
    assign layer4_outputs[356] = (layer3_outputs[1772]) & (layer3_outputs[4856]);
    assign layer4_outputs[357] = 1'b0;
    assign layer4_outputs[358] = ~(layer3_outputs[919]);
    assign layer4_outputs[359] = layer3_outputs[3295];
    assign layer4_outputs[360] = ~(layer3_outputs[849]);
    assign layer4_outputs[361] = ~(layer3_outputs[423]) | (layer3_outputs[3135]);
    assign layer4_outputs[362] = ~(layer3_outputs[4540]);
    assign layer4_outputs[363] = ~(layer3_outputs[792]);
    assign layer4_outputs[364] = (layer3_outputs[1964]) & ~(layer3_outputs[3976]);
    assign layer4_outputs[365] = (layer3_outputs[5108]) | (layer3_outputs[1981]);
    assign layer4_outputs[366] = ~(layer3_outputs[919]) | (layer3_outputs[1840]);
    assign layer4_outputs[367] = ~(layer3_outputs[34]) | (layer3_outputs[3605]);
    assign layer4_outputs[368] = 1'b1;
    assign layer4_outputs[369] = layer3_outputs[1393];
    assign layer4_outputs[370] = ~(layer3_outputs[651]) | (layer3_outputs[2090]);
    assign layer4_outputs[371] = layer3_outputs[3850];
    assign layer4_outputs[372] = ~(layer3_outputs[1449]);
    assign layer4_outputs[373] = ~(layer3_outputs[4233]) | (layer3_outputs[1470]);
    assign layer4_outputs[374] = ~(layer3_outputs[5034]);
    assign layer4_outputs[375] = (layer3_outputs[2731]) & ~(layer3_outputs[2884]);
    assign layer4_outputs[376] = (layer3_outputs[312]) | (layer3_outputs[278]);
    assign layer4_outputs[377] = ~(layer3_outputs[3113]);
    assign layer4_outputs[378] = ~(layer3_outputs[1090]) | (layer3_outputs[2438]);
    assign layer4_outputs[379] = (layer3_outputs[2840]) ^ (layer3_outputs[1885]);
    assign layer4_outputs[380] = ~(layer3_outputs[2014]);
    assign layer4_outputs[381] = 1'b0;
    assign layer4_outputs[382] = layer3_outputs[4456];
    assign layer4_outputs[383] = 1'b1;
    assign layer4_outputs[384] = (layer3_outputs[2848]) & (layer3_outputs[2334]);
    assign layer4_outputs[385] = (layer3_outputs[1095]) ^ (layer3_outputs[3891]);
    assign layer4_outputs[386] = (layer3_outputs[2166]) & ~(layer3_outputs[1211]);
    assign layer4_outputs[387] = (layer3_outputs[2896]) & ~(layer3_outputs[5117]);
    assign layer4_outputs[388] = layer3_outputs[3016];
    assign layer4_outputs[389] = layer3_outputs[2373];
    assign layer4_outputs[390] = ~(layer3_outputs[3361]);
    assign layer4_outputs[391] = (layer3_outputs[1720]) & ~(layer3_outputs[4388]);
    assign layer4_outputs[392] = ~((layer3_outputs[4963]) & (layer3_outputs[4702]));
    assign layer4_outputs[393] = (layer3_outputs[4687]) & ~(layer3_outputs[3594]);
    assign layer4_outputs[394] = layer3_outputs[3207];
    assign layer4_outputs[395] = (layer3_outputs[520]) ^ (layer3_outputs[487]);
    assign layer4_outputs[396] = (layer3_outputs[425]) & (layer3_outputs[3595]);
    assign layer4_outputs[397] = ~(layer3_outputs[1376]);
    assign layer4_outputs[398] = ~(layer3_outputs[3010]) | (layer3_outputs[1250]);
    assign layer4_outputs[399] = ~(layer3_outputs[4886]) | (layer3_outputs[4236]);
    assign layer4_outputs[400] = ~((layer3_outputs[2505]) & (layer3_outputs[1500]));
    assign layer4_outputs[401] = 1'b0;
    assign layer4_outputs[402] = ~(layer3_outputs[108]) | (layer3_outputs[3554]);
    assign layer4_outputs[403] = (layer3_outputs[1068]) & ~(layer3_outputs[1507]);
    assign layer4_outputs[404] = ~(layer3_outputs[3703]);
    assign layer4_outputs[405] = ~((layer3_outputs[4390]) | (layer3_outputs[2215]));
    assign layer4_outputs[406] = (layer3_outputs[979]) | (layer3_outputs[1822]);
    assign layer4_outputs[407] = (layer3_outputs[396]) & (layer3_outputs[3430]);
    assign layer4_outputs[408] = 1'b0;
    assign layer4_outputs[409] = layer3_outputs[3853];
    assign layer4_outputs[410] = (layer3_outputs[2459]) & ~(layer3_outputs[4765]);
    assign layer4_outputs[411] = 1'b0;
    assign layer4_outputs[412] = layer3_outputs[47];
    assign layer4_outputs[413] = layer3_outputs[3088];
    assign layer4_outputs[414] = ~(layer3_outputs[754]);
    assign layer4_outputs[415] = ~(layer3_outputs[4065]) | (layer3_outputs[1646]);
    assign layer4_outputs[416] = ~((layer3_outputs[3824]) ^ (layer3_outputs[690]));
    assign layer4_outputs[417] = ~((layer3_outputs[4394]) | (layer3_outputs[1384]));
    assign layer4_outputs[418] = ~((layer3_outputs[699]) & (layer3_outputs[5087]));
    assign layer4_outputs[419] = (layer3_outputs[4761]) ^ (layer3_outputs[2007]);
    assign layer4_outputs[420] = ~(layer3_outputs[602]) | (layer3_outputs[1918]);
    assign layer4_outputs[421] = layer3_outputs[4151];
    assign layer4_outputs[422] = ~(layer3_outputs[632]);
    assign layer4_outputs[423] = 1'b0;
    assign layer4_outputs[424] = ~((layer3_outputs[4434]) | (layer3_outputs[2423]));
    assign layer4_outputs[425] = 1'b1;
    assign layer4_outputs[426] = (layer3_outputs[567]) ^ (layer3_outputs[807]);
    assign layer4_outputs[427] = (layer3_outputs[3791]) & (layer3_outputs[712]);
    assign layer4_outputs[428] = ~((layer3_outputs[1246]) | (layer3_outputs[4773]));
    assign layer4_outputs[429] = layer3_outputs[4463];
    assign layer4_outputs[430] = ~(layer3_outputs[2945]);
    assign layer4_outputs[431] = (layer3_outputs[3718]) & ~(layer3_outputs[4050]);
    assign layer4_outputs[432] = layer3_outputs[3690];
    assign layer4_outputs[433] = ~(layer3_outputs[3819]);
    assign layer4_outputs[434] = ~(layer3_outputs[2871]);
    assign layer4_outputs[435] = ~(layer3_outputs[868]) | (layer3_outputs[4439]);
    assign layer4_outputs[436] = (layer3_outputs[3765]) | (layer3_outputs[164]);
    assign layer4_outputs[437] = ~(layer3_outputs[304]);
    assign layer4_outputs[438] = layer3_outputs[4758];
    assign layer4_outputs[439] = (layer3_outputs[1856]) & ~(layer3_outputs[1952]);
    assign layer4_outputs[440] = layer3_outputs[1442];
    assign layer4_outputs[441] = layer3_outputs[3618];
    assign layer4_outputs[442] = ~(layer3_outputs[3534]);
    assign layer4_outputs[443] = layer3_outputs[4670];
    assign layer4_outputs[444] = (layer3_outputs[3430]) & ~(layer3_outputs[697]);
    assign layer4_outputs[445] = ~(layer3_outputs[3553]);
    assign layer4_outputs[446] = ~(layer3_outputs[2275]);
    assign layer4_outputs[447] = ~(layer3_outputs[2108]);
    assign layer4_outputs[448] = layer3_outputs[4737];
    assign layer4_outputs[449] = layer3_outputs[4355];
    assign layer4_outputs[450] = layer3_outputs[1344];
    assign layer4_outputs[451] = ~(layer3_outputs[4134]);
    assign layer4_outputs[452] = (layer3_outputs[3623]) ^ (layer3_outputs[1876]);
    assign layer4_outputs[453] = (layer3_outputs[37]) | (layer3_outputs[3733]);
    assign layer4_outputs[454] = layer3_outputs[338];
    assign layer4_outputs[455] = layer3_outputs[2736];
    assign layer4_outputs[456] = ~(layer3_outputs[3594]) | (layer3_outputs[365]);
    assign layer4_outputs[457] = (layer3_outputs[4196]) & (layer3_outputs[1098]);
    assign layer4_outputs[458] = layer3_outputs[4912];
    assign layer4_outputs[459] = ~(layer3_outputs[182]) | (layer3_outputs[163]);
    assign layer4_outputs[460] = ~(layer3_outputs[523]) | (layer3_outputs[1898]);
    assign layer4_outputs[461] = ~((layer3_outputs[3030]) | (layer3_outputs[2251]));
    assign layer4_outputs[462] = (layer3_outputs[4382]) ^ (layer3_outputs[2814]);
    assign layer4_outputs[463] = ~(layer3_outputs[199]);
    assign layer4_outputs[464] = ~(layer3_outputs[4135]) | (layer3_outputs[3167]);
    assign layer4_outputs[465] = layer3_outputs[194];
    assign layer4_outputs[466] = ~(layer3_outputs[2024]) | (layer3_outputs[881]);
    assign layer4_outputs[467] = ~(layer3_outputs[2966]) | (layer3_outputs[3389]);
    assign layer4_outputs[468] = 1'b1;
    assign layer4_outputs[469] = ~((layer3_outputs[3284]) | (layer3_outputs[546]));
    assign layer4_outputs[470] = 1'b1;
    assign layer4_outputs[471] = (layer3_outputs[782]) & (layer3_outputs[387]);
    assign layer4_outputs[472] = layer3_outputs[4847];
    assign layer4_outputs[473] = ~(layer3_outputs[1845]);
    assign layer4_outputs[474] = (layer3_outputs[4709]) ^ (layer3_outputs[2880]);
    assign layer4_outputs[475] = ~(layer3_outputs[1678]) | (layer3_outputs[4046]);
    assign layer4_outputs[476] = ~(layer3_outputs[4133]);
    assign layer4_outputs[477] = layer3_outputs[3895];
    assign layer4_outputs[478] = layer3_outputs[1400];
    assign layer4_outputs[479] = ~(layer3_outputs[3170]);
    assign layer4_outputs[480] = (layer3_outputs[2124]) | (layer3_outputs[1495]);
    assign layer4_outputs[481] = ~(layer3_outputs[2227]);
    assign layer4_outputs[482] = (layer3_outputs[2362]) & (layer3_outputs[377]);
    assign layer4_outputs[483] = ~(layer3_outputs[1849]) | (layer3_outputs[1524]);
    assign layer4_outputs[484] = ~(layer3_outputs[2084]) | (layer3_outputs[1175]);
    assign layer4_outputs[485] = ~(layer3_outputs[4450]);
    assign layer4_outputs[486] = 1'b1;
    assign layer4_outputs[487] = ~((layer3_outputs[2722]) ^ (layer3_outputs[3683]));
    assign layer4_outputs[488] = ~(layer3_outputs[4360]);
    assign layer4_outputs[489] = ~(layer3_outputs[4498]);
    assign layer4_outputs[490] = ~(layer3_outputs[4847]) | (layer3_outputs[3976]);
    assign layer4_outputs[491] = ~(layer3_outputs[4274]);
    assign layer4_outputs[492] = layer3_outputs[3463];
    assign layer4_outputs[493] = layer3_outputs[5031];
    assign layer4_outputs[494] = ~(layer3_outputs[1869]);
    assign layer4_outputs[495] = (layer3_outputs[555]) ^ (layer3_outputs[5009]);
    assign layer4_outputs[496] = ~((layer3_outputs[847]) ^ (layer3_outputs[929]));
    assign layer4_outputs[497] = layer3_outputs[430];
    assign layer4_outputs[498] = ~(layer3_outputs[513]);
    assign layer4_outputs[499] = layer3_outputs[1750];
    assign layer4_outputs[500] = ~(layer3_outputs[2150]);
    assign layer4_outputs[501] = ~(layer3_outputs[4531]);
    assign layer4_outputs[502] = ~(layer3_outputs[3112]) | (layer3_outputs[5057]);
    assign layer4_outputs[503] = (layer3_outputs[2257]) & (layer3_outputs[4464]);
    assign layer4_outputs[504] = layer3_outputs[4319];
    assign layer4_outputs[505] = layer3_outputs[4943];
    assign layer4_outputs[506] = layer3_outputs[4530];
    assign layer4_outputs[507] = (layer3_outputs[3580]) & ~(layer3_outputs[3960]);
    assign layer4_outputs[508] = layer3_outputs[2995];
    assign layer4_outputs[509] = (layer3_outputs[2388]) ^ (layer3_outputs[2991]);
    assign layer4_outputs[510] = (layer3_outputs[3287]) & ~(layer3_outputs[16]);
    assign layer4_outputs[511] = ~(layer3_outputs[4711]);
    assign layer4_outputs[512] = ~(layer3_outputs[942]) | (layer3_outputs[3451]);
    assign layer4_outputs[513] = 1'b0;
    assign layer4_outputs[514] = layer3_outputs[76];
    assign layer4_outputs[515] = ~(layer3_outputs[119]);
    assign layer4_outputs[516] = layer3_outputs[4228];
    assign layer4_outputs[517] = (layer3_outputs[1212]) & ~(layer3_outputs[48]);
    assign layer4_outputs[518] = (layer3_outputs[4042]) | (layer3_outputs[3480]);
    assign layer4_outputs[519] = ~(layer3_outputs[311]);
    assign layer4_outputs[520] = 1'b1;
    assign layer4_outputs[521] = ~(layer3_outputs[3780]) | (layer3_outputs[4223]);
    assign layer4_outputs[522] = (layer3_outputs[2363]) & ~(layer3_outputs[4357]);
    assign layer4_outputs[523] = ~((layer3_outputs[2263]) ^ (layer3_outputs[1438]));
    assign layer4_outputs[524] = layer3_outputs[4715];
    assign layer4_outputs[525] = ~((layer3_outputs[4708]) & (layer3_outputs[2690]));
    assign layer4_outputs[526] = ~(layer3_outputs[3966]);
    assign layer4_outputs[527] = (layer3_outputs[2908]) & ~(layer3_outputs[2870]);
    assign layer4_outputs[528] = ~((layer3_outputs[1763]) ^ (layer3_outputs[2834]));
    assign layer4_outputs[529] = layer3_outputs[615];
    assign layer4_outputs[530] = layer3_outputs[4008];
    assign layer4_outputs[531] = 1'b1;
    assign layer4_outputs[532] = (layer3_outputs[4139]) & ~(layer3_outputs[2606]);
    assign layer4_outputs[533] = ~(layer3_outputs[3372]);
    assign layer4_outputs[534] = (layer3_outputs[590]) | (layer3_outputs[343]);
    assign layer4_outputs[535] = ~((layer3_outputs[3014]) & (layer3_outputs[4345]));
    assign layer4_outputs[536] = ~((layer3_outputs[3128]) | (layer3_outputs[2333]));
    assign layer4_outputs[537] = 1'b1;
    assign layer4_outputs[538] = (layer3_outputs[778]) | (layer3_outputs[1901]);
    assign layer4_outputs[539] = (layer3_outputs[1280]) & ~(layer3_outputs[2508]);
    assign layer4_outputs[540] = ~(layer3_outputs[1106]);
    assign layer4_outputs[541] = ~((layer3_outputs[14]) | (layer3_outputs[4036]));
    assign layer4_outputs[542] = layer3_outputs[44];
    assign layer4_outputs[543] = ~(layer3_outputs[1308]);
    assign layer4_outputs[544] = ~(layer3_outputs[4294]) | (layer3_outputs[1231]);
    assign layer4_outputs[545] = 1'b1;
    assign layer4_outputs[546] = 1'b1;
    assign layer4_outputs[547] = 1'b0;
    assign layer4_outputs[548] = layer3_outputs[2111];
    assign layer4_outputs[549] = layer3_outputs[1028];
    assign layer4_outputs[550] = (layer3_outputs[1755]) | (layer3_outputs[3652]);
    assign layer4_outputs[551] = ~((layer3_outputs[1418]) | (layer3_outputs[1760]));
    assign layer4_outputs[552] = ~((layer3_outputs[333]) | (layer3_outputs[4528]));
    assign layer4_outputs[553] = (layer3_outputs[764]) | (layer3_outputs[4177]);
    assign layer4_outputs[554] = ~(layer3_outputs[2546]);
    assign layer4_outputs[555] = (layer3_outputs[4742]) & ~(layer3_outputs[4093]);
    assign layer4_outputs[556] = ~(layer3_outputs[4374]);
    assign layer4_outputs[557] = ~(layer3_outputs[1876]) | (layer3_outputs[223]);
    assign layer4_outputs[558] = ~((layer3_outputs[2559]) | (layer3_outputs[5008]));
    assign layer4_outputs[559] = ~(layer3_outputs[9]) | (layer3_outputs[1197]);
    assign layer4_outputs[560] = ~(layer3_outputs[428]);
    assign layer4_outputs[561] = (layer3_outputs[3508]) | (layer3_outputs[3407]);
    assign layer4_outputs[562] = ~(layer3_outputs[4341]);
    assign layer4_outputs[563] = ~(layer3_outputs[4755]) | (layer3_outputs[1353]);
    assign layer4_outputs[564] = (layer3_outputs[1489]) & (layer3_outputs[3466]);
    assign layer4_outputs[565] = (layer3_outputs[1524]) & ~(layer3_outputs[2129]);
    assign layer4_outputs[566] = ~(layer3_outputs[4142]);
    assign layer4_outputs[567] = 1'b1;
    assign layer4_outputs[568] = layer3_outputs[3834];
    assign layer4_outputs[569] = 1'b0;
    assign layer4_outputs[570] = layer3_outputs[1529];
    assign layer4_outputs[571] = ~(layer3_outputs[1529]);
    assign layer4_outputs[572] = (layer3_outputs[3400]) | (layer3_outputs[4853]);
    assign layer4_outputs[573] = layer3_outputs[624];
    assign layer4_outputs[574] = (layer3_outputs[4438]) | (layer3_outputs[698]);
    assign layer4_outputs[575] = layer3_outputs[4902];
    assign layer4_outputs[576] = ~((layer3_outputs[2765]) | (layer3_outputs[4410]));
    assign layer4_outputs[577] = ~(layer3_outputs[2793]);
    assign layer4_outputs[578] = (layer3_outputs[1448]) & ~(layer3_outputs[3799]);
    assign layer4_outputs[579] = (layer3_outputs[4515]) & (layer3_outputs[2331]);
    assign layer4_outputs[580] = layer3_outputs[2320];
    assign layer4_outputs[581] = ~((layer3_outputs[2899]) ^ (layer3_outputs[4706]));
    assign layer4_outputs[582] = layer3_outputs[5110];
    assign layer4_outputs[583] = ~((layer3_outputs[85]) ^ (layer3_outputs[3708]));
    assign layer4_outputs[584] = layer3_outputs[3312];
    assign layer4_outputs[585] = ~((layer3_outputs[3177]) ^ (layer3_outputs[4512]));
    assign layer4_outputs[586] = 1'b0;
    assign layer4_outputs[587] = (layer3_outputs[4017]) & ~(layer3_outputs[2389]);
    assign layer4_outputs[588] = ~(layer3_outputs[1510]);
    assign layer4_outputs[589] = 1'b1;
    assign layer4_outputs[590] = layer3_outputs[1873];
    assign layer4_outputs[591] = ~(layer3_outputs[4896]);
    assign layer4_outputs[592] = (layer3_outputs[3567]) & ~(layer3_outputs[3260]);
    assign layer4_outputs[593] = ~(layer3_outputs[473]) | (layer3_outputs[880]);
    assign layer4_outputs[594] = (layer3_outputs[5021]) ^ (layer3_outputs[1096]);
    assign layer4_outputs[595] = 1'b0;
    assign layer4_outputs[596] = ~((layer3_outputs[4620]) | (layer3_outputs[4560]));
    assign layer4_outputs[597] = layer3_outputs[4578];
    assign layer4_outputs[598] = ~(layer3_outputs[3069]) | (layer3_outputs[2507]);
    assign layer4_outputs[599] = ~(layer3_outputs[3779]) | (layer3_outputs[3866]);
    assign layer4_outputs[600] = ~(layer3_outputs[2196]);
    assign layer4_outputs[601] = ~(layer3_outputs[4542]) | (layer3_outputs[4349]);
    assign layer4_outputs[602] = (layer3_outputs[3008]) | (layer3_outputs[1190]);
    assign layer4_outputs[603] = ~(layer3_outputs[1911]) | (layer3_outputs[3522]);
    assign layer4_outputs[604] = ~(layer3_outputs[3763]);
    assign layer4_outputs[605] = (layer3_outputs[4408]) & ~(layer3_outputs[111]);
    assign layer4_outputs[606] = (layer3_outputs[2518]) & (layer3_outputs[3168]);
    assign layer4_outputs[607] = (layer3_outputs[2904]) & ~(layer3_outputs[2164]);
    assign layer4_outputs[608] = layer3_outputs[4887];
    assign layer4_outputs[609] = layer3_outputs[437];
    assign layer4_outputs[610] = (layer3_outputs[3095]) & ~(layer3_outputs[4418]);
    assign layer4_outputs[611] = ~((layer3_outputs[1701]) & (layer3_outputs[2062]));
    assign layer4_outputs[612] = layer3_outputs[3302];
    assign layer4_outputs[613] = ~(layer3_outputs[478]);
    assign layer4_outputs[614] = ~((layer3_outputs[2202]) | (layer3_outputs[2201]));
    assign layer4_outputs[615] = 1'b0;
    assign layer4_outputs[616] = (layer3_outputs[3540]) & (layer3_outputs[4288]);
    assign layer4_outputs[617] = layer3_outputs[4487];
    assign layer4_outputs[618] = layer3_outputs[324];
    assign layer4_outputs[619] = layer3_outputs[2827];
    assign layer4_outputs[620] = layer3_outputs[4007];
    assign layer4_outputs[621] = ~(layer3_outputs[364]);
    assign layer4_outputs[622] = ~(layer3_outputs[4269]) | (layer3_outputs[1157]);
    assign layer4_outputs[623] = ~(layer3_outputs[525]);
    assign layer4_outputs[624] = (layer3_outputs[353]) ^ (layer3_outputs[4622]);
    assign layer4_outputs[625] = ~(layer3_outputs[3117]);
    assign layer4_outputs[626] = layer3_outputs[425];
    assign layer4_outputs[627] = ~(layer3_outputs[4447]);
    assign layer4_outputs[628] = ~((layer3_outputs[2845]) | (layer3_outputs[3402]));
    assign layer4_outputs[629] = (layer3_outputs[3917]) & ~(layer3_outputs[3523]);
    assign layer4_outputs[630] = ~(layer3_outputs[2425]);
    assign layer4_outputs[631] = (layer3_outputs[1657]) | (layer3_outputs[3130]);
    assign layer4_outputs[632] = (layer3_outputs[965]) | (layer3_outputs[2337]);
    assign layer4_outputs[633] = ~(layer3_outputs[4201]);
    assign layer4_outputs[634] = layer3_outputs[694];
    assign layer4_outputs[635] = ~(layer3_outputs[740]) | (layer3_outputs[1568]);
    assign layer4_outputs[636] = layer3_outputs[2233];
    assign layer4_outputs[637] = layer3_outputs[3886];
    assign layer4_outputs[638] = (layer3_outputs[2620]) & ~(layer3_outputs[3928]);
    assign layer4_outputs[639] = layer3_outputs[3952];
    assign layer4_outputs[640] = (layer3_outputs[3737]) & (layer3_outputs[4879]);
    assign layer4_outputs[641] = 1'b1;
    assign layer4_outputs[642] = ~(layer3_outputs[4734]);
    assign layer4_outputs[643] = ~(layer3_outputs[2816]) | (layer3_outputs[2541]);
    assign layer4_outputs[644] = layer3_outputs[865];
    assign layer4_outputs[645] = (layer3_outputs[4823]) & ~(layer3_outputs[2758]);
    assign layer4_outputs[646] = (layer3_outputs[36]) & (layer3_outputs[1989]);
    assign layer4_outputs[647] = 1'b0;
    assign layer4_outputs[648] = layer3_outputs[4740];
    assign layer4_outputs[649] = ~(layer3_outputs[4431]);
    assign layer4_outputs[650] = (layer3_outputs[4947]) & ~(layer3_outputs[3309]);
    assign layer4_outputs[651] = layer3_outputs[2319];
    assign layer4_outputs[652] = ~(layer3_outputs[4920]) | (layer3_outputs[2891]);
    assign layer4_outputs[653] = layer3_outputs[3497];
    assign layer4_outputs[654] = layer3_outputs[177];
    assign layer4_outputs[655] = ~(layer3_outputs[5065]);
    assign layer4_outputs[656] = ~((layer3_outputs[2231]) & (layer3_outputs[492]));
    assign layer4_outputs[657] = ~(layer3_outputs[1338]);
    assign layer4_outputs[658] = 1'b1;
    assign layer4_outputs[659] = (layer3_outputs[3032]) | (layer3_outputs[3087]);
    assign layer4_outputs[660] = (layer3_outputs[1446]) & ~(layer3_outputs[1967]);
    assign layer4_outputs[661] = ~((layer3_outputs[1256]) ^ (layer3_outputs[4966]));
    assign layer4_outputs[662] = ~(layer3_outputs[2531]);
    assign layer4_outputs[663] = ~(layer3_outputs[3233]);
    assign layer4_outputs[664] = (layer3_outputs[3961]) & ~(layer3_outputs[1993]);
    assign layer4_outputs[665] = (layer3_outputs[754]) | (layer3_outputs[786]);
    assign layer4_outputs[666] = (layer3_outputs[4953]) ^ (layer3_outputs[1194]);
    assign layer4_outputs[667] = (layer3_outputs[4801]) & ~(layer3_outputs[2138]);
    assign layer4_outputs[668] = (layer3_outputs[3627]) & (layer3_outputs[4789]);
    assign layer4_outputs[669] = layer3_outputs[4098];
    assign layer4_outputs[670] = layer3_outputs[947];
    assign layer4_outputs[671] = layer3_outputs[3665];
    assign layer4_outputs[672] = ~(layer3_outputs[31]);
    assign layer4_outputs[673] = layer3_outputs[3255];
    assign layer4_outputs[674] = ~(layer3_outputs[2955]) | (layer3_outputs[914]);
    assign layer4_outputs[675] = (layer3_outputs[2950]) & ~(layer3_outputs[3753]);
    assign layer4_outputs[676] = (layer3_outputs[853]) & ~(layer3_outputs[26]);
    assign layer4_outputs[677] = ~(layer3_outputs[2484]);
    assign layer4_outputs[678] = ~(layer3_outputs[3186]);
    assign layer4_outputs[679] = ~((layer3_outputs[1394]) & (layer3_outputs[568]));
    assign layer4_outputs[680] = ~((layer3_outputs[2265]) & (layer3_outputs[4302]));
    assign layer4_outputs[681] = 1'b1;
    assign layer4_outputs[682] = ~(layer3_outputs[4245]);
    assign layer4_outputs[683] = ~(layer3_outputs[63]) | (layer3_outputs[3843]);
    assign layer4_outputs[684] = layer3_outputs[3243];
    assign layer4_outputs[685] = (layer3_outputs[4525]) & (layer3_outputs[1350]);
    assign layer4_outputs[686] = layer3_outputs[427];
    assign layer4_outputs[687] = (layer3_outputs[3456]) & ~(layer3_outputs[3533]);
    assign layer4_outputs[688] = (layer3_outputs[1554]) & (layer3_outputs[3736]);
    assign layer4_outputs[689] = ~(layer3_outputs[1918]);
    assign layer4_outputs[690] = ~(layer3_outputs[1062]) | (layer3_outputs[934]);
    assign layer4_outputs[691] = layer3_outputs[1358];
    assign layer4_outputs[692] = ~((layer3_outputs[1719]) & (layer3_outputs[873]));
    assign layer4_outputs[693] = (layer3_outputs[1647]) | (layer3_outputs[4385]);
    assign layer4_outputs[694] = ~(layer3_outputs[2360]);
    assign layer4_outputs[695] = ~(layer3_outputs[4246]);
    assign layer4_outputs[696] = ~(layer3_outputs[4158]);
    assign layer4_outputs[697] = ~((layer3_outputs[3560]) | (layer3_outputs[2660]));
    assign layer4_outputs[698] = layer3_outputs[2224];
    assign layer4_outputs[699] = layer3_outputs[3110];
    assign layer4_outputs[700] = layer3_outputs[1398];
    assign layer4_outputs[701] = ~(layer3_outputs[100]) | (layer3_outputs[3281]);
    assign layer4_outputs[702] = (layer3_outputs[2104]) | (layer3_outputs[3987]);
    assign layer4_outputs[703] = (layer3_outputs[282]) & ~(layer3_outputs[1963]);
    assign layer4_outputs[704] = layer3_outputs[4348];
    assign layer4_outputs[705] = layer3_outputs[3174];
    assign layer4_outputs[706] = layer3_outputs[1679];
    assign layer4_outputs[707] = layer3_outputs[2299];
    assign layer4_outputs[708] = ~((layer3_outputs[4672]) | (layer3_outputs[1008]));
    assign layer4_outputs[709] = ~(layer3_outputs[4603]);
    assign layer4_outputs[710] = layer3_outputs[134];
    assign layer4_outputs[711] = ~(layer3_outputs[2117]) | (layer3_outputs[3212]);
    assign layer4_outputs[712] = 1'b1;
    assign layer4_outputs[713] = ~(layer3_outputs[1676]);
    assign layer4_outputs[714] = ~(layer3_outputs[4813]) | (layer3_outputs[3419]);
    assign layer4_outputs[715] = layer3_outputs[40];
    assign layer4_outputs[716] = (layer3_outputs[1431]) | (layer3_outputs[3777]);
    assign layer4_outputs[717] = layer3_outputs[536];
    assign layer4_outputs[718] = ~(layer3_outputs[812]);
    assign layer4_outputs[719] = ~(layer3_outputs[1414]);
    assign layer4_outputs[720] = (layer3_outputs[1110]) | (layer3_outputs[1191]);
    assign layer4_outputs[721] = 1'b0;
    assign layer4_outputs[722] = layer3_outputs[1479];
    assign layer4_outputs[723] = (layer3_outputs[518]) | (layer3_outputs[1900]);
    assign layer4_outputs[724] = 1'b0;
    assign layer4_outputs[725] = (layer3_outputs[197]) & (layer3_outputs[128]);
    assign layer4_outputs[726] = layer3_outputs[3937];
    assign layer4_outputs[727] = ~((layer3_outputs[578]) | (layer3_outputs[633]));
    assign layer4_outputs[728] = (layer3_outputs[372]) & ~(layer3_outputs[4954]);
    assign layer4_outputs[729] = (layer3_outputs[3773]) | (layer3_outputs[4173]);
    assign layer4_outputs[730] = ~((layer3_outputs[203]) | (layer3_outputs[3568]));
    assign layer4_outputs[731] = ~(layer3_outputs[4539]);
    assign layer4_outputs[732] = ~((layer3_outputs[2029]) & (layer3_outputs[4604]));
    assign layer4_outputs[733] = ~((layer3_outputs[5104]) ^ (layer3_outputs[1359]));
    assign layer4_outputs[734] = ~(layer3_outputs[2974]);
    assign layer4_outputs[735] = layer3_outputs[990];
    assign layer4_outputs[736] = (layer3_outputs[4054]) | (layer3_outputs[4946]);
    assign layer4_outputs[737] = 1'b0;
    assign layer4_outputs[738] = ~(layer3_outputs[1215]);
    assign layer4_outputs[739] = ~(layer3_outputs[1995]) | (layer3_outputs[3581]);
    assign layer4_outputs[740] = ~(layer3_outputs[3542]);
    assign layer4_outputs[741] = layer3_outputs[1654];
    assign layer4_outputs[742] = ~((layer3_outputs[4859]) & (layer3_outputs[3089]));
    assign layer4_outputs[743] = ~(layer3_outputs[1378]);
    assign layer4_outputs[744] = (layer3_outputs[1161]) & ~(layer3_outputs[5032]);
    assign layer4_outputs[745] = ~(layer3_outputs[323]);
    assign layer4_outputs[746] = (layer3_outputs[2909]) ^ (layer3_outputs[1797]);
    assign layer4_outputs[747] = ~(layer3_outputs[2458]) | (layer3_outputs[2394]);
    assign layer4_outputs[748] = (layer3_outputs[4995]) & ~(layer3_outputs[2972]);
    assign layer4_outputs[749] = (layer3_outputs[3502]) & ~(layer3_outputs[2158]);
    assign layer4_outputs[750] = layer3_outputs[3616];
    assign layer4_outputs[751] = ~(layer3_outputs[1355]);
    assign layer4_outputs[752] = layer3_outputs[4642];
    assign layer4_outputs[753] = ~(layer3_outputs[4242]);
    assign layer4_outputs[754] = 1'b1;
    assign layer4_outputs[755] = layer3_outputs[4765];
    assign layer4_outputs[756] = (layer3_outputs[596]) & ~(layer3_outputs[2060]);
    assign layer4_outputs[757] = (layer3_outputs[2361]) | (layer3_outputs[1226]);
    assign layer4_outputs[758] = ~(layer3_outputs[1358]);
    assign layer4_outputs[759] = ~(layer3_outputs[3644]);
    assign layer4_outputs[760] = ~(layer3_outputs[1269]);
    assign layer4_outputs[761] = ~((layer3_outputs[5095]) & (layer3_outputs[1870]));
    assign layer4_outputs[762] = ~(layer3_outputs[832]) | (layer3_outputs[3092]);
    assign layer4_outputs[763] = ~(layer3_outputs[4863]);
    assign layer4_outputs[764] = ~(layer3_outputs[103]);
    assign layer4_outputs[765] = ~(layer3_outputs[4238]);
    assign layer4_outputs[766] = layer3_outputs[3137];
    assign layer4_outputs[767] = 1'b0;
    assign layer4_outputs[768] = ~((layer3_outputs[574]) & (layer3_outputs[2208]));
    assign layer4_outputs[769] = ~(layer3_outputs[3786]);
    assign layer4_outputs[770] = ~(layer3_outputs[2708]);
    assign layer4_outputs[771] = layer3_outputs[1904];
    assign layer4_outputs[772] = ~(layer3_outputs[3869]);
    assign layer4_outputs[773] = ~(layer3_outputs[3985]);
    assign layer4_outputs[774] = ~(layer3_outputs[3571]);
    assign layer4_outputs[775] = ~(layer3_outputs[1119]);
    assign layer4_outputs[776] = layer3_outputs[4268];
    assign layer4_outputs[777] = ~(layer3_outputs[3061]) | (layer3_outputs[4678]);
    assign layer4_outputs[778] = (layer3_outputs[1462]) ^ (layer3_outputs[4005]);
    assign layer4_outputs[779] = ~(layer3_outputs[4802]);
    assign layer4_outputs[780] = (layer3_outputs[2333]) & ~(layer3_outputs[4533]);
    assign layer4_outputs[781] = (layer3_outputs[4890]) & (layer3_outputs[4547]);
    assign layer4_outputs[782] = ~(layer3_outputs[587]);
    assign layer4_outputs[783] = layer3_outputs[3242];
    assign layer4_outputs[784] = layer3_outputs[4922];
    assign layer4_outputs[785] = (layer3_outputs[428]) & ~(layer3_outputs[3088]);
    assign layer4_outputs[786] = ~(layer3_outputs[5069]);
    assign layer4_outputs[787] = (layer3_outputs[569]) ^ (layer3_outputs[3975]);
    assign layer4_outputs[788] = ~(layer3_outputs[3432]);
    assign layer4_outputs[789] = ~(layer3_outputs[44]);
    assign layer4_outputs[790] = ~(layer3_outputs[1729]) | (layer3_outputs[2008]);
    assign layer4_outputs[791] = (layer3_outputs[4880]) & ~(layer3_outputs[2288]);
    assign layer4_outputs[792] = ~((layer3_outputs[1219]) & (layer3_outputs[4971]));
    assign layer4_outputs[793] = (layer3_outputs[3823]) & ~(layer3_outputs[1088]);
    assign layer4_outputs[794] = ~((layer3_outputs[2745]) ^ (layer3_outputs[4497]));
    assign layer4_outputs[795] = ~((layer3_outputs[5109]) | (layer3_outputs[3455]));
    assign layer4_outputs[796] = layer3_outputs[1089];
    assign layer4_outputs[797] = ~((layer3_outputs[2167]) | (layer3_outputs[2893]));
    assign layer4_outputs[798] = ~((layer3_outputs[4643]) ^ (layer3_outputs[4664]));
    assign layer4_outputs[799] = layer3_outputs[583];
    assign layer4_outputs[800] = (layer3_outputs[4120]) & ~(layer3_outputs[4753]);
    assign layer4_outputs[801] = (layer3_outputs[2033]) & ~(layer3_outputs[1522]);
    assign layer4_outputs[802] = 1'b1;
    assign layer4_outputs[803] = layer3_outputs[3297];
    assign layer4_outputs[804] = layer3_outputs[4003];
    assign layer4_outputs[805] = layer3_outputs[354];
    assign layer4_outputs[806] = (layer3_outputs[4099]) & (layer3_outputs[493]);
    assign layer4_outputs[807] = layer3_outputs[3580];
    assign layer4_outputs[808] = ~(layer3_outputs[1074]) | (layer3_outputs[3037]);
    assign layer4_outputs[809] = layer3_outputs[2049];
    assign layer4_outputs[810] = (layer3_outputs[623]) | (layer3_outputs[1127]);
    assign layer4_outputs[811] = (layer3_outputs[988]) | (layer3_outputs[4090]);
    assign layer4_outputs[812] = 1'b0;
    assign layer4_outputs[813] = layer3_outputs[525];
    assign layer4_outputs[814] = (layer3_outputs[1365]) ^ (layer3_outputs[3264]);
    assign layer4_outputs[815] = (layer3_outputs[2453]) ^ (layer3_outputs[4750]);
    assign layer4_outputs[816] = (layer3_outputs[2198]) & (layer3_outputs[724]);
    assign layer4_outputs[817] = layer3_outputs[2555];
    assign layer4_outputs[818] = ~(layer3_outputs[3653]);
    assign layer4_outputs[819] = ~(layer3_outputs[2195]);
    assign layer4_outputs[820] = layer3_outputs[1895];
    assign layer4_outputs[821] = ~(layer3_outputs[2082]);
    assign layer4_outputs[822] = (layer3_outputs[1129]) | (layer3_outputs[459]);
    assign layer4_outputs[823] = ~((layer3_outputs[4429]) & (layer3_outputs[2324]));
    assign layer4_outputs[824] = layer3_outputs[1867];
    assign layer4_outputs[825] = ~(layer3_outputs[1837]);
    assign layer4_outputs[826] = 1'b0;
    assign layer4_outputs[827] = (layer3_outputs[3822]) & ~(layer3_outputs[4634]);
    assign layer4_outputs[828] = ~(layer3_outputs[961]);
    assign layer4_outputs[829] = 1'b1;
    assign layer4_outputs[830] = ~(layer3_outputs[301]);
    assign layer4_outputs[831] = 1'b0;
    assign layer4_outputs[832] = ~(layer3_outputs[1591]);
    assign layer4_outputs[833] = ~(layer3_outputs[3757]);
    assign layer4_outputs[834] = 1'b1;
    assign layer4_outputs[835] = (layer3_outputs[2867]) & ~(layer3_outputs[4160]);
    assign layer4_outputs[836] = 1'b0;
    assign layer4_outputs[837] = ~(layer3_outputs[391]);
    assign layer4_outputs[838] = 1'b1;
    assign layer4_outputs[839] = ~((layer3_outputs[1238]) | (layer3_outputs[2686]));
    assign layer4_outputs[840] = 1'b0;
    assign layer4_outputs[841] = layer3_outputs[1091];
    assign layer4_outputs[842] = (layer3_outputs[573]) & ~(layer3_outputs[2371]);
    assign layer4_outputs[843] = ~((layer3_outputs[1273]) & (layer3_outputs[1346]));
    assign layer4_outputs[844] = ~((layer3_outputs[3655]) & (layer3_outputs[3408]));
    assign layer4_outputs[845] = ~(layer3_outputs[968]);
    assign layer4_outputs[846] = (layer3_outputs[4325]) | (layer3_outputs[1415]);
    assign layer4_outputs[847] = (layer3_outputs[704]) | (layer3_outputs[1275]);
    assign layer4_outputs[848] = 1'b0;
    assign layer4_outputs[849] = (layer3_outputs[3034]) & ~(layer3_outputs[38]);
    assign layer4_outputs[850] = layer3_outputs[2673];
    assign layer4_outputs[851] = (layer3_outputs[1549]) & ~(layer3_outputs[1517]);
    assign layer4_outputs[852] = layer3_outputs[1900];
    assign layer4_outputs[853] = layer3_outputs[1011];
    assign layer4_outputs[854] = (layer3_outputs[1771]) & (layer3_outputs[1190]);
    assign layer4_outputs[855] = ~(layer3_outputs[2171]) | (layer3_outputs[2477]);
    assign layer4_outputs[856] = ~((layer3_outputs[2140]) ^ (layer3_outputs[4405]));
    assign layer4_outputs[857] = layer3_outputs[2416];
    assign layer4_outputs[858] = (layer3_outputs[1789]) & (layer3_outputs[3558]);
    assign layer4_outputs[859] = (layer3_outputs[4908]) ^ (layer3_outputs[3973]);
    assign layer4_outputs[860] = 1'b0;
    assign layer4_outputs[861] = 1'b1;
    assign layer4_outputs[862] = ~(layer3_outputs[3448]);
    assign layer4_outputs[863] = ~((layer3_outputs[1195]) & (layer3_outputs[2083]));
    assign layer4_outputs[864] = layer3_outputs[252];
    assign layer4_outputs[865] = (layer3_outputs[1228]) | (layer3_outputs[2228]);
    assign layer4_outputs[866] = ~(layer3_outputs[1599]);
    assign layer4_outputs[867] = 1'b1;
    assign layer4_outputs[868] = ~(layer3_outputs[3612]) | (layer3_outputs[1406]);
    assign layer4_outputs[869] = (layer3_outputs[2272]) & ~(layer3_outputs[2207]);
    assign layer4_outputs[870] = ~((layer3_outputs[1966]) | (layer3_outputs[245]));
    assign layer4_outputs[871] = layer3_outputs[4519];
    assign layer4_outputs[872] = layer3_outputs[4494];
    assign layer4_outputs[873] = 1'b0;
    assign layer4_outputs[874] = (layer3_outputs[184]) | (layer3_outputs[3136]);
    assign layer4_outputs[875] = (layer3_outputs[1422]) & ~(layer3_outputs[4099]);
    assign layer4_outputs[876] = ~((layer3_outputs[863]) | (layer3_outputs[508]));
    assign layer4_outputs[877] = (layer3_outputs[4595]) | (layer3_outputs[3077]);
    assign layer4_outputs[878] = 1'b0;
    assign layer4_outputs[879] = 1'b1;
    assign layer4_outputs[880] = ~((layer3_outputs[3691]) & (layer3_outputs[3540]));
    assign layer4_outputs[881] = ~(layer3_outputs[3205]) | (layer3_outputs[1597]);
    assign layer4_outputs[882] = layer3_outputs[3646];
    assign layer4_outputs[883] = (layer3_outputs[4386]) & (layer3_outputs[4118]);
    assign layer4_outputs[884] = layer3_outputs[2913];
    assign layer4_outputs[885] = layer3_outputs[4722];
    assign layer4_outputs[886] = ~((layer3_outputs[663]) & (layer3_outputs[4883]));
    assign layer4_outputs[887] = layer3_outputs[687];
    assign layer4_outputs[888] = layer3_outputs[1171];
    assign layer4_outputs[889] = ~(layer3_outputs[4105]);
    assign layer4_outputs[890] = ~(layer3_outputs[1537]);
    assign layer4_outputs[891] = 1'b1;
    assign layer4_outputs[892] = ~(layer3_outputs[4164]);
    assign layer4_outputs[893] = (layer3_outputs[4662]) & ~(layer3_outputs[1280]);
    assign layer4_outputs[894] = (layer3_outputs[2717]) & ~(layer3_outputs[266]);
    assign layer4_outputs[895] = ~(layer3_outputs[2719]);
    assign layer4_outputs[896] = ~((layer3_outputs[115]) & (layer3_outputs[168]));
    assign layer4_outputs[897] = 1'b0;
    assign layer4_outputs[898] = (layer3_outputs[3950]) & ~(layer3_outputs[560]);
    assign layer4_outputs[899] = ~(layer3_outputs[267]) | (layer3_outputs[4091]);
    assign layer4_outputs[900] = ~((layer3_outputs[2311]) | (layer3_outputs[4854]));
    assign layer4_outputs[901] = ~(layer3_outputs[3164]) | (layer3_outputs[4918]);
    assign layer4_outputs[902] = ~(layer3_outputs[933]);
    assign layer4_outputs[903] = ~(layer3_outputs[1561]);
    assign layer4_outputs[904] = 1'b0;
    assign layer4_outputs[905] = ~(layer3_outputs[4265]);
    assign layer4_outputs[906] = layer3_outputs[4913];
    assign layer4_outputs[907] = ~(layer3_outputs[4686]);
    assign layer4_outputs[908] = ~(layer3_outputs[1364]);
    assign layer4_outputs[909] = (layer3_outputs[954]) & (layer3_outputs[2020]);
    assign layer4_outputs[910] = ~(layer3_outputs[3939]);
    assign layer4_outputs[911] = ~((layer3_outputs[678]) | (layer3_outputs[2584]));
    assign layer4_outputs[912] = layer3_outputs[3798];
    assign layer4_outputs[913] = 1'b0;
    assign layer4_outputs[914] = layer3_outputs[3634];
    assign layer4_outputs[915] = ~(layer3_outputs[2885]) | (layer3_outputs[4572]);
    assign layer4_outputs[916] = ~(layer3_outputs[4046]);
    assign layer4_outputs[917] = ~(layer3_outputs[81]) | (layer3_outputs[2704]);
    assign layer4_outputs[918] = ~(layer3_outputs[4579]) | (layer3_outputs[1319]);
    assign layer4_outputs[919] = ~((layer3_outputs[2085]) & (layer3_outputs[4144]));
    assign layer4_outputs[920] = 1'b1;
    assign layer4_outputs[921] = ~(layer3_outputs[4114]);
    assign layer4_outputs[922] = layer3_outputs[2583];
    assign layer4_outputs[923] = 1'b0;
    assign layer4_outputs[924] = layer3_outputs[1002];
    assign layer4_outputs[925] = ~((layer3_outputs[1735]) | (layer3_outputs[3348]));
    assign layer4_outputs[926] = ~(layer3_outputs[432]);
    assign layer4_outputs[927] = ~((layer3_outputs[3598]) & (layer3_outputs[1943]));
    assign layer4_outputs[928] = ~((layer3_outputs[368]) | (layer3_outputs[2990]));
    assign layer4_outputs[929] = ~(layer3_outputs[3916]);
    assign layer4_outputs[930] = (layer3_outputs[610]) & ~(layer3_outputs[4062]);
    assign layer4_outputs[931] = ~((layer3_outputs[417]) & (layer3_outputs[3028]));
    assign layer4_outputs[932] = ~((layer3_outputs[4293]) | (layer3_outputs[779]));
    assign layer4_outputs[933] = ~(layer3_outputs[5100]) | (layer3_outputs[253]);
    assign layer4_outputs[934] = ~((layer3_outputs[4754]) & (layer3_outputs[902]));
    assign layer4_outputs[935] = ~(layer3_outputs[3918]) | (layer3_outputs[4421]);
    assign layer4_outputs[936] = (layer3_outputs[2497]) & ~(layer3_outputs[3615]);
    assign layer4_outputs[937] = layer3_outputs[3590];
    assign layer4_outputs[938] = layer3_outputs[3933];
    assign layer4_outputs[939] = ~((layer3_outputs[4693]) ^ (layer3_outputs[332]));
    assign layer4_outputs[940] = ~(layer3_outputs[2255]);
    assign layer4_outputs[941] = (layer3_outputs[3614]) & (layer3_outputs[3889]);
    assign layer4_outputs[942] = ~((layer3_outputs[3396]) & (layer3_outputs[4070]));
    assign layer4_outputs[943] = (layer3_outputs[2077]) ^ (layer3_outputs[3122]);
    assign layer4_outputs[944] = ~(layer3_outputs[4518]);
    assign layer4_outputs[945] = (layer3_outputs[2445]) & ~(layer3_outputs[2667]);
    assign layer4_outputs[946] = ~(layer3_outputs[4475]) | (layer3_outputs[2448]);
    assign layer4_outputs[947] = ~(layer3_outputs[2948]);
    assign layer4_outputs[948] = (layer3_outputs[3412]) ^ (layer3_outputs[4243]);
    assign layer4_outputs[949] = ~(layer3_outputs[4123]);
    assign layer4_outputs[950] = (layer3_outputs[706]) & ~(layer3_outputs[4736]);
    assign layer4_outputs[951] = ~(layer3_outputs[3698]);
    assign layer4_outputs[952] = layer3_outputs[4911];
    assign layer4_outputs[953] = (layer3_outputs[1268]) & (layer3_outputs[5007]);
    assign layer4_outputs[954] = (layer3_outputs[3538]) & ~(layer3_outputs[3378]);
    assign layer4_outputs[955] = 1'b0;
    assign layer4_outputs[956] = ~((layer3_outputs[3516]) | (layer3_outputs[1297]));
    assign layer4_outputs[957] = layer3_outputs[3832];
    assign layer4_outputs[958] = ~(layer3_outputs[1847]) | (layer3_outputs[4184]);
    assign layer4_outputs[959] = ~((layer3_outputs[4582]) ^ (layer3_outputs[1798]));
    assign layer4_outputs[960] = 1'b1;
    assign layer4_outputs[961] = ~(layer3_outputs[697]);
    assign layer4_outputs[962] = ~(layer3_outputs[4041]);
    assign layer4_outputs[963] = ~((layer3_outputs[537]) | (layer3_outputs[2261]));
    assign layer4_outputs[964] = (layer3_outputs[4454]) & ~(layer3_outputs[3736]);
    assign layer4_outputs[965] = (layer3_outputs[4353]) & ~(layer3_outputs[3091]);
    assign layer4_outputs[966] = ~(layer3_outputs[5041]) | (layer3_outputs[303]);
    assign layer4_outputs[967] = ~(layer3_outputs[767]);
    assign layer4_outputs[968] = ~((layer3_outputs[710]) & (layer3_outputs[1322]));
    assign layer4_outputs[969] = (layer3_outputs[1112]) & ~(layer3_outputs[780]);
    assign layer4_outputs[970] = 1'b1;
    assign layer4_outputs[971] = layer3_outputs[4421];
    assign layer4_outputs[972] = ~(layer3_outputs[581]);
    assign layer4_outputs[973] = ~(layer3_outputs[5007]);
    assign layer4_outputs[974] = ~(layer3_outputs[4351]) | (layer3_outputs[4635]);
    assign layer4_outputs[975] = ~(layer3_outputs[3315]) | (layer3_outputs[1638]);
    assign layer4_outputs[976] = ~((layer3_outputs[2164]) & (layer3_outputs[4260]));
    assign layer4_outputs[977] = ~(layer3_outputs[4837]);
    assign layer4_outputs[978] = ~(layer3_outputs[305]) | (layer3_outputs[3299]);
    assign layer4_outputs[979] = ~((layer3_outputs[967]) ^ (layer3_outputs[2070]));
    assign layer4_outputs[980] = (layer3_outputs[2693]) | (layer3_outputs[1484]);
    assign layer4_outputs[981] = (layer3_outputs[810]) | (layer3_outputs[3031]);
    assign layer4_outputs[982] = 1'b0;
    assign layer4_outputs[983] = (layer3_outputs[3183]) | (layer3_outputs[2194]);
    assign layer4_outputs[984] = layer3_outputs[2487];
    assign layer4_outputs[985] = ~(layer3_outputs[1200]);
    assign layer4_outputs[986] = layer3_outputs[419];
    assign layer4_outputs[987] = ~(layer3_outputs[2431]) | (layer3_outputs[1003]);
    assign layer4_outputs[988] = layer3_outputs[2383];
    assign layer4_outputs[989] = layer3_outputs[4289];
    assign layer4_outputs[990] = ~(layer3_outputs[1398]);
    assign layer4_outputs[991] = 1'b1;
    assign layer4_outputs[992] = (layer3_outputs[4730]) & (layer3_outputs[1380]);
    assign layer4_outputs[993] = layer3_outputs[2326];
    assign layer4_outputs[994] = (layer3_outputs[3989]) & ~(layer3_outputs[1512]);
    assign layer4_outputs[995] = layer3_outputs[304];
    assign layer4_outputs[996] = ~(layer3_outputs[1628]) | (layer3_outputs[4305]);
    assign layer4_outputs[997] = (layer3_outputs[1880]) | (layer3_outputs[1893]);
    assign layer4_outputs[998] = ~(layer3_outputs[4435]);
    assign layer4_outputs[999] = layer3_outputs[3173];
    assign layer4_outputs[1000] = layer3_outputs[3286];
    assign layer4_outputs[1001] = layer3_outputs[3893];
    assign layer4_outputs[1002] = (layer3_outputs[1307]) & ~(layer3_outputs[2124]);
    assign layer4_outputs[1003] = (layer3_outputs[1427]) ^ (layer3_outputs[3722]);
    assign layer4_outputs[1004] = layer3_outputs[4106];
    assign layer4_outputs[1005] = layer3_outputs[4427];
    assign layer4_outputs[1006] = ~(layer3_outputs[178]) | (layer3_outputs[4125]);
    assign layer4_outputs[1007] = (layer3_outputs[1807]) & ~(layer3_outputs[73]);
    assign layer4_outputs[1008] = layer3_outputs[3168];
    assign layer4_outputs[1009] = (layer3_outputs[1626]) & ~(layer3_outputs[2963]);
    assign layer4_outputs[1010] = (layer3_outputs[999]) & ~(layer3_outputs[3894]);
    assign layer4_outputs[1011] = layer3_outputs[2355];
    assign layer4_outputs[1012] = layer3_outputs[5097];
    assign layer4_outputs[1013] = (layer3_outputs[3684]) ^ (layer3_outputs[4096]);
    assign layer4_outputs[1014] = layer3_outputs[3921];
    assign layer4_outputs[1015] = layer3_outputs[1976];
    assign layer4_outputs[1016] = layer3_outputs[3357];
    assign layer4_outputs[1017] = ~(layer3_outputs[94]);
    assign layer4_outputs[1018] = ~((layer3_outputs[2547]) | (layer3_outputs[3766]));
    assign layer4_outputs[1019] = ~(layer3_outputs[2913]);
    assign layer4_outputs[1020] = ~((layer3_outputs[1674]) ^ (layer3_outputs[3474]));
    assign layer4_outputs[1021] = ~(layer3_outputs[3239]);
    assign layer4_outputs[1022] = ~(layer3_outputs[3651]);
    assign layer4_outputs[1023] = layer3_outputs[160];
    assign layer4_outputs[1024] = ~(layer3_outputs[2523]);
    assign layer4_outputs[1025] = ~(layer3_outputs[230]);
    assign layer4_outputs[1026] = (layer3_outputs[4355]) & ~(layer3_outputs[1587]);
    assign layer4_outputs[1027] = layer3_outputs[1473];
    assign layer4_outputs[1028] = ~((layer3_outputs[2535]) & (layer3_outputs[257]));
    assign layer4_outputs[1029] = 1'b0;
    assign layer4_outputs[1030] = (layer3_outputs[5019]) & ~(layer3_outputs[1301]);
    assign layer4_outputs[1031] = ~((layer3_outputs[2760]) | (layer3_outputs[289]));
    assign layer4_outputs[1032] = (layer3_outputs[335]) & ~(layer3_outputs[3629]);
    assign layer4_outputs[1033] = (layer3_outputs[3908]) & ~(layer3_outputs[2742]);
    assign layer4_outputs[1034] = ~(layer3_outputs[1149]);
    assign layer4_outputs[1035] = ~(layer3_outputs[1631]);
    assign layer4_outputs[1036] = ~(layer3_outputs[660]) | (layer3_outputs[2488]);
    assign layer4_outputs[1037] = ~(layer3_outputs[4175]);
    assign layer4_outputs[1038] = ~(layer3_outputs[4655]) | (layer3_outputs[1669]);
    assign layer4_outputs[1039] = layer3_outputs[4896];
    assign layer4_outputs[1040] = ~((layer3_outputs[4848]) & (layer3_outputs[3082]));
    assign layer4_outputs[1041] = ~(layer3_outputs[3963]) | (layer3_outputs[4011]);
    assign layer4_outputs[1042] = layer3_outputs[2072];
    assign layer4_outputs[1043] = ~((layer3_outputs[2385]) | (layer3_outputs[1625]));
    assign layer4_outputs[1044] = ~((layer3_outputs[3948]) ^ (layer3_outputs[3293]));
    assign layer4_outputs[1045] = ~(layer3_outputs[4522]);
    assign layer4_outputs[1046] = (layer3_outputs[95]) ^ (layer3_outputs[2873]);
    assign layer4_outputs[1047] = ~(layer3_outputs[4465]) | (layer3_outputs[4786]);
    assign layer4_outputs[1048] = layer3_outputs[596];
    assign layer4_outputs[1049] = ~((layer3_outputs[317]) ^ (layer3_outputs[1846]));
    assign layer4_outputs[1050] = layer3_outputs[3671];
    assign layer4_outputs[1051] = layer3_outputs[4298];
    assign layer4_outputs[1052] = ~(layer3_outputs[149]);
    assign layer4_outputs[1053] = ~((layer3_outputs[2363]) | (layer3_outputs[666]));
    assign layer4_outputs[1054] = ~(layer3_outputs[3838]);
    assign layer4_outputs[1055] = layer3_outputs[1115];
    assign layer4_outputs[1056] = ~(layer3_outputs[4401]);
    assign layer4_outputs[1057] = ~(layer3_outputs[1075]);
    assign layer4_outputs[1058] = ~(layer3_outputs[4672]);
    assign layer4_outputs[1059] = (layer3_outputs[2517]) & ~(layer3_outputs[2029]);
    assign layer4_outputs[1060] = layer3_outputs[3645];
    assign layer4_outputs[1061] = (layer3_outputs[2407]) ^ (layer3_outputs[2600]);
    assign layer4_outputs[1062] = layer3_outputs[1906];
    assign layer4_outputs[1063] = ~(layer3_outputs[3426]) | (layer3_outputs[3622]);
    assign layer4_outputs[1064] = ~(layer3_outputs[1426]);
    assign layer4_outputs[1065] = (layer3_outputs[546]) & ~(layer3_outputs[3433]);
    assign layer4_outputs[1066] = ~(layer3_outputs[4519]);
    assign layer4_outputs[1067] = layer3_outputs[2938];
    assign layer4_outputs[1068] = (layer3_outputs[543]) & ~(layer3_outputs[800]);
    assign layer4_outputs[1069] = ~(layer3_outputs[2162]);
    assign layer4_outputs[1070] = ~(layer3_outputs[1152]);
    assign layer4_outputs[1071] = 1'b1;
    assign layer4_outputs[1072] = ~(layer3_outputs[1797]);
    assign layer4_outputs[1073] = ~(layer3_outputs[1325]);
    assign layer4_outputs[1074] = ~(layer3_outputs[4342]);
    assign layer4_outputs[1075] = ~(layer3_outputs[3586]);
    assign layer4_outputs[1076] = ~(layer3_outputs[1048]) | (layer3_outputs[2603]);
    assign layer4_outputs[1077] = layer3_outputs[1518];
    assign layer4_outputs[1078] = ~((layer3_outputs[1734]) ^ (layer3_outputs[26]));
    assign layer4_outputs[1079] = ~((layer3_outputs[89]) | (layer3_outputs[2902]));
    assign layer4_outputs[1080] = ~(layer3_outputs[1173]) | (layer3_outputs[1]);
    assign layer4_outputs[1081] = (layer3_outputs[351]) | (layer3_outputs[2048]);
    assign layer4_outputs[1082] = ~(layer3_outputs[16]) | (layer3_outputs[2636]);
    assign layer4_outputs[1083] = ~((layer3_outputs[1920]) | (layer3_outputs[2797]));
    assign layer4_outputs[1084] = (layer3_outputs[3068]) | (layer3_outputs[2372]);
    assign layer4_outputs[1085] = layer3_outputs[966];
    assign layer4_outputs[1086] = (layer3_outputs[2120]) & (layer3_outputs[657]);
    assign layer4_outputs[1087] = 1'b0;
    assign layer4_outputs[1088] = ~(layer3_outputs[4170]);
    assign layer4_outputs[1089] = (layer3_outputs[2115]) & ~(layer3_outputs[4960]);
    assign layer4_outputs[1090] = 1'b1;
    assign layer4_outputs[1091] = ~(layer3_outputs[2826]) | (layer3_outputs[2897]);
    assign layer4_outputs[1092] = 1'b0;
    assign layer4_outputs[1093] = 1'b0;
    assign layer4_outputs[1094] = (layer3_outputs[2465]) & ~(layer3_outputs[3818]);
    assign layer4_outputs[1095] = ~(layer3_outputs[643]);
    assign layer4_outputs[1096] = ~(layer3_outputs[929]);
    assign layer4_outputs[1097] = 1'b0;
    assign layer4_outputs[1098] = ~(layer3_outputs[175]);
    assign layer4_outputs[1099] = ~(layer3_outputs[4722]) | (layer3_outputs[3903]);
    assign layer4_outputs[1100] = 1'b1;
    assign layer4_outputs[1101] = layer3_outputs[4126];
    assign layer4_outputs[1102] = ~(layer3_outputs[2664]);
    assign layer4_outputs[1103] = layer3_outputs[823];
    assign layer4_outputs[1104] = ~(layer3_outputs[4152]);
    assign layer4_outputs[1105] = (layer3_outputs[3564]) & (layer3_outputs[1672]);
    assign layer4_outputs[1106] = ~(layer3_outputs[3187]);
    assign layer4_outputs[1107] = ~(layer3_outputs[334]);
    assign layer4_outputs[1108] = (layer3_outputs[1639]) & ~(layer3_outputs[4031]);
    assign layer4_outputs[1109] = layer3_outputs[3247];
    assign layer4_outputs[1110] = ~(layer3_outputs[143]);
    assign layer4_outputs[1111] = layer3_outputs[2297];
    assign layer4_outputs[1112] = (layer3_outputs[1776]) | (layer3_outputs[3687]);
    assign layer4_outputs[1113] = ~((layer3_outputs[3434]) ^ (layer3_outputs[171]));
    assign layer4_outputs[1114] = ~((layer3_outputs[204]) | (layer3_outputs[2752]));
    assign layer4_outputs[1115] = layer3_outputs[43];
    assign layer4_outputs[1116] = layer3_outputs[3900];
    assign layer4_outputs[1117] = 1'b1;
    assign layer4_outputs[1118] = (layer3_outputs[3063]) ^ (layer3_outputs[5052]);
    assign layer4_outputs[1119] = (layer3_outputs[211]) | (layer3_outputs[4350]);
    assign layer4_outputs[1120] = ~(layer3_outputs[3235]) | (layer3_outputs[3815]);
    assign layer4_outputs[1121] = (layer3_outputs[1616]) & ~(layer3_outputs[1067]);
    assign layer4_outputs[1122] = ~((layer3_outputs[65]) & (layer3_outputs[2806]));
    assign layer4_outputs[1123] = ~(layer3_outputs[3909]);
    assign layer4_outputs[1124] = (layer3_outputs[1132]) ^ (layer3_outputs[1554]);
    assign layer4_outputs[1125] = ~((layer3_outputs[3829]) ^ (layer3_outputs[962]));
    assign layer4_outputs[1126] = layer3_outputs[2369];
    assign layer4_outputs[1127] = (layer3_outputs[4048]) & ~(layer3_outputs[3658]);
    assign layer4_outputs[1128] = ~(layer3_outputs[1626]) | (layer3_outputs[1430]);
    assign layer4_outputs[1129] = ~(layer3_outputs[5111]);
    assign layer4_outputs[1130] = layer3_outputs[4251];
    assign layer4_outputs[1131] = layer3_outputs[4514];
    assign layer4_outputs[1132] = layer3_outputs[1080];
    assign layer4_outputs[1133] = ~((layer3_outputs[2727]) ^ (layer3_outputs[2366]));
    assign layer4_outputs[1134] = ~(layer3_outputs[2106]) | (layer3_outputs[3267]);
    assign layer4_outputs[1135] = (layer3_outputs[1128]) & (layer3_outputs[121]);
    assign layer4_outputs[1136] = ~((layer3_outputs[3172]) ^ (layer3_outputs[3813]));
    assign layer4_outputs[1137] = ~(layer3_outputs[1176]);
    assign layer4_outputs[1138] = (layer3_outputs[772]) & ~(layer3_outputs[1713]);
    assign layer4_outputs[1139] = layer3_outputs[4062];
    assign layer4_outputs[1140] = ~(layer3_outputs[152]);
    assign layer4_outputs[1141] = layer3_outputs[2500];
    assign layer4_outputs[1142] = 1'b1;
    assign layer4_outputs[1143] = (layer3_outputs[415]) & (layer3_outputs[802]);
    assign layer4_outputs[1144] = (layer3_outputs[2756]) & ~(layer3_outputs[1958]);
    assign layer4_outputs[1145] = ~(layer3_outputs[4225]);
    assign layer4_outputs[1146] = layer3_outputs[3403];
    assign layer4_outputs[1147] = layer3_outputs[64];
    assign layer4_outputs[1148] = ~((layer3_outputs[1289]) ^ (layer3_outputs[4983]));
    assign layer4_outputs[1149] = layer3_outputs[1001];
    assign layer4_outputs[1150] = ~(layer3_outputs[1155]);
    assign layer4_outputs[1151] = ~(layer3_outputs[3740]) | (layer3_outputs[519]);
    assign layer4_outputs[1152] = 1'b1;
    assign layer4_outputs[1153] = layer3_outputs[3626];
    assign layer4_outputs[1154] = ~(layer3_outputs[2189]);
    assign layer4_outputs[1155] = ~(layer3_outputs[3752]);
    assign layer4_outputs[1156] = ~((layer3_outputs[2820]) ^ (layer3_outputs[3648]));
    assign layer4_outputs[1157] = ~(layer3_outputs[421]);
    assign layer4_outputs[1158] = (layer3_outputs[3971]) & (layer3_outputs[3969]);
    assign layer4_outputs[1159] = ~(layer3_outputs[3487]) | (layer3_outputs[4513]);
    assign layer4_outputs[1160] = layer3_outputs[70];
    assign layer4_outputs[1161] = (layer3_outputs[2319]) & ~(layer3_outputs[3624]);
    assign layer4_outputs[1162] = ~(layer3_outputs[4808]);
    assign layer4_outputs[1163] = (layer3_outputs[2915]) & ~(layer3_outputs[162]);
    assign layer4_outputs[1164] = ~(layer3_outputs[1206]);
    assign layer4_outputs[1165] = layer3_outputs[3114];
    assign layer4_outputs[1166] = ~(layer3_outputs[2298]);
    assign layer4_outputs[1167] = layer3_outputs[3308];
    assign layer4_outputs[1168] = ~(layer3_outputs[2369]);
    assign layer4_outputs[1169] = ~(layer3_outputs[4173]);
    assign layer4_outputs[1170] = ~(layer3_outputs[4064]) | (layer3_outputs[4891]);
    assign layer4_outputs[1171] = layer3_outputs[2039];
    assign layer4_outputs[1172] = ~((layer3_outputs[4770]) ^ (layer3_outputs[1354]));
    assign layer4_outputs[1173] = (layer3_outputs[3200]) & ~(layer3_outputs[1180]);
    assign layer4_outputs[1174] = ~(layer3_outputs[3034]);
    assign layer4_outputs[1175] = (layer3_outputs[4024]) & ~(layer3_outputs[198]);
    assign layer4_outputs[1176] = (layer3_outputs[1431]) & (layer3_outputs[4365]);
    assign layer4_outputs[1177] = ~((layer3_outputs[872]) ^ (layer3_outputs[1877]));
    assign layer4_outputs[1178] = ~(layer3_outputs[3853]) | (layer3_outputs[2474]);
    assign layer4_outputs[1179] = (layer3_outputs[2663]) ^ (layer3_outputs[3536]);
    assign layer4_outputs[1180] = (layer3_outputs[2263]) | (layer3_outputs[3139]);
    assign layer4_outputs[1181] = (layer3_outputs[3062]) & ~(layer3_outputs[611]);
    assign layer4_outputs[1182] = ~(layer3_outputs[694]);
    assign layer4_outputs[1183] = (layer3_outputs[4794]) & ~(layer3_outputs[4949]);
    assign layer4_outputs[1184] = ~(layer3_outputs[3640]) | (layer3_outputs[5098]);
    assign layer4_outputs[1185] = layer3_outputs[3295];
    assign layer4_outputs[1186] = layer3_outputs[1493];
    assign layer4_outputs[1187] = ~(layer3_outputs[3904]);
    assign layer4_outputs[1188] = ~(layer3_outputs[1189]);
    assign layer4_outputs[1189] = ~(layer3_outputs[2093]);
    assign layer4_outputs[1190] = 1'b0;
    assign layer4_outputs[1191] = (layer3_outputs[3468]) & ~(layer3_outputs[4335]);
    assign layer4_outputs[1192] = ~(layer3_outputs[2336]);
    assign layer4_outputs[1193] = layer3_outputs[1564];
    assign layer4_outputs[1194] = ~(layer3_outputs[4855]);
    assign layer4_outputs[1195] = (layer3_outputs[4255]) & ~(layer3_outputs[4386]);
    assign layer4_outputs[1196] = ~(layer3_outputs[2582]);
    assign layer4_outputs[1197] = ~(layer3_outputs[4224]);
    assign layer4_outputs[1198] = ~((layer3_outputs[1348]) | (layer3_outputs[3278]));
    assign layer4_outputs[1199] = ~((layer3_outputs[908]) & (layer3_outputs[4240]));
    assign layer4_outputs[1200] = ~(layer3_outputs[678]) | (layer3_outputs[988]);
    assign layer4_outputs[1201] = layer3_outputs[504];
    assign layer4_outputs[1202] = (layer3_outputs[2395]) ^ (layer3_outputs[3772]);
    assign layer4_outputs[1203] = ~((layer3_outputs[4074]) | (layer3_outputs[3536]));
    assign layer4_outputs[1204] = (layer3_outputs[184]) | (layer3_outputs[3972]);
    assign layer4_outputs[1205] = layer3_outputs[1366];
    assign layer4_outputs[1206] = (layer3_outputs[3779]) & ~(layer3_outputs[4991]);
    assign layer4_outputs[1207] = layer3_outputs[2108];
    assign layer4_outputs[1208] = layer3_outputs[1396];
    assign layer4_outputs[1209] = layer3_outputs[4037];
    assign layer4_outputs[1210] = 1'b0;
    assign layer4_outputs[1211] = layer3_outputs[1615];
    assign layer4_outputs[1212] = layer3_outputs[1612];
    assign layer4_outputs[1213] = ~(layer3_outputs[3037]) | (layer3_outputs[4841]);
    assign layer4_outputs[1214] = 1'b1;
    assign layer4_outputs[1215] = ~(layer3_outputs[3544]);
    assign layer4_outputs[1216] = layer3_outputs[937];
    assign layer4_outputs[1217] = ~((layer3_outputs[3658]) | (layer3_outputs[2467]));
    assign layer4_outputs[1218] = (layer3_outputs[584]) & ~(layer3_outputs[1158]);
    assign layer4_outputs[1219] = (layer3_outputs[2999]) & ~(layer3_outputs[3454]);
    assign layer4_outputs[1220] = ~(layer3_outputs[25]);
    assign layer4_outputs[1221] = ~(layer3_outputs[3291]);
    assign layer4_outputs[1222] = ~((layer3_outputs[1128]) | (layer3_outputs[2689]));
    assign layer4_outputs[1223] = layer3_outputs[1094];
    assign layer4_outputs[1224] = ~(layer3_outputs[1988]);
    assign layer4_outputs[1225] = ~(layer3_outputs[1796]);
    assign layer4_outputs[1226] = layer3_outputs[3498];
    assign layer4_outputs[1227] = 1'b1;
    assign layer4_outputs[1228] = layer3_outputs[4530];
    assign layer4_outputs[1229] = (layer3_outputs[4713]) & ~(layer3_outputs[337]);
    assign layer4_outputs[1230] = ~(layer3_outputs[13]);
    assign layer4_outputs[1231] = layer3_outputs[4477];
    assign layer4_outputs[1232] = (layer3_outputs[3343]) & (layer3_outputs[4423]);
    assign layer4_outputs[1233] = ~(layer3_outputs[739]);
    assign layer4_outputs[1234] = layer3_outputs[2970];
    assign layer4_outputs[1235] = (layer3_outputs[2428]) & ~(layer3_outputs[4039]);
    assign layer4_outputs[1236] = ~(layer3_outputs[594]);
    assign layer4_outputs[1237] = ~((layer3_outputs[4961]) & (layer3_outputs[2804]));
    assign layer4_outputs[1238] = (layer3_outputs[4908]) & ~(layer3_outputs[4957]);
    assign layer4_outputs[1239] = layer3_outputs[4525];
    assign layer4_outputs[1240] = ~((layer3_outputs[977]) & (layer3_outputs[4729]));
    assign layer4_outputs[1241] = ~(layer3_outputs[2001]);
    assign layer4_outputs[1242] = layer3_outputs[4129];
    assign layer4_outputs[1243] = ~(layer3_outputs[346]);
    assign layer4_outputs[1244] = ~((layer3_outputs[1381]) & (layer3_outputs[2647]));
    assign layer4_outputs[1245] = (layer3_outputs[453]) ^ (layer3_outputs[812]);
    assign layer4_outputs[1246] = ~(layer3_outputs[4030]);
    assign layer4_outputs[1247] = ~(layer3_outputs[1100]);
    assign layer4_outputs[1248] = ~((layer3_outputs[2836]) | (layer3_outputs[3576]));
    assign layer4_outputs[1249] = ~((layer3_outputs[3650]) | (layer3_outputs[2937]));
    assign layer4_outputs[1250] = layer3_outputs[1451];
    assign layer4_outputs[1251] = (layer3_outputs[2103]) & ~(layer3_outputs[2192]);
    assign layer4_outputs[1252] = 1'b0;
    assign layer4_outputs[1253] = (layer3_outputs[1274]) & (layer3_outputs[850]);
    assign layer4_outputs[1254] = ~((layer3_outputs[3561]) & (layer3_outputs[3152]));
    assign layer4_outputs[1255] = 1'b0;
    assign layer4_outputs[1256] = ~(layer3_outputs[4220]);
    assign layer4_outputs[1257] = layer3_outputs[932];
    assign layer4_outputs[1258] = ~(layer3_outputs[2406]);
    assign layer4_outputs[1259] = ~(layer3_outputs[150]) | (layer3_outputs[4588]);
    assign layer4_outputs[1260] = (layer3_outputs[1646]) & (layer3_outputs[2708]);
    assign layer4_outputs[1261] = ~(layer3_outputs[266]);
    assign layer4_outputs[1262] = ~((layer3_outputs[1294]) | (layer3_outputs[3113]));
    assign layer4_outputs[1263] = ~(layer3_outputs[2694]);
    assign layer4_outputs[1264] = ~((layer3_outputs[2684]) | (layer3_outputs[1713]));
    assign layer4_outputs[1265] = ~(layer3_outputs[996]);
    assign layer4_outputs[1266] = ~((layer3_outputs[280]) ^ (layer3_outputs[2986]));
    assign layer4_outputs[1267] = 1'b0;
    assign layer4_outputs[1268] = 1'b0;
    assign layer4_outputs[1269] = ~(layer3_outputs[677]);
    assign layer4_outputs[1270] = ~(layer3_outputs[4779]);
    assign layer4_outputs[1271] = 1'b0;
    assign layer4_outputs[1272] = ~(layer3_outputs[1764]) | (layer3_outputs[2854]);
    assign layer4_outputs[1273] = layer3_outputs[1053];
    assign layer4_outputs[1274] = (layer3_outputs[4442]) & (layer3_outputs[3548]);
    assign layer4_outputs[1275] = 1'b0;
    assign layer4_outputs[1276] = (layer3_outputs[3052]) & ~(layer3_outputs[4340]);
    assign layer4_outputs[1277] = ~(layer3_outputs[729]) | (layer3_outputs[1136]);
    assign layer4_outputs[1278] = (layer3_outputs[4344]) | (layer3_outputs[1345]);
    assign layer4_outputs[1279] = layer3_outputs[1387];
    assign layer4_outputs[1280] = layer3_outputs[4104];
    assign layer4_outputs[1281] = (layer3_outputs[3617]) | (layer3_outputs[1527]);
    assign layer4_outputs[1282] = 1'b1;
    assign layer4_outputs[1283] = ~(layer3_outputs[4352]);
    assign layer4_outputs[1284] = (layer3_outputs[2055]) & ~(layer3_outputs[5059]);
    assign layer4_outputs[1285] = (layer3_outputs[2565]) & ~(layer3_outputs[4286]);
    assign layer4_outputs[1286] = ~(layer3_outputs[388]);
    assign layer4_outputs[1287] = (layer3_outputs[4825]) & ~(layer3_outputs[975]);
    assign layer4_outputs[1288] = ~((layer3_outputs[4699]) & (layer3_outputs[4391]));
    assign layer4_outputs[1289] = 1'b1;
    assign layer4_outputs[1290] = ~((layer3_outputs[1474]) | (layer3_outputs[1924]));
    assign layer4_outputs[1291] = ~(layer3_outputs[4803]) | (layer3_outputs[262]);
    assign layer4_outputs[1292] = (layer3_outputs[3216]) & ~(layer3_outputs[3515]);
    assign layer4_outputs[1293] = (layer3_outputs[331]) & ~(layer3_outputs[4333]);
    assign layer4_outputs[1294] = layer3_outputs[2482];
    assign layer4_outputs[1295] = ~(layer3_outputs[878]);
    assign layer4_outputs[1296] = ~(layer3_outputs[830]);
    assign layer4_outputs[1297] = ~((layer3_outputs[1077]) ^ (layer3_outputs[424]));
    assign layer4_outputs[1298] = ~(layer3_outputs[3223]);
    assign layer4_outputs[1299] = ~(layer3_outputs[3525]);
    assign layer4_outputs[1300] = (layer3_outputs[104]) | (layer3_outputs[2065]);
    assign layer4_outputs[1301] = 1'b1;
    assign layer4_outputs[1302] = layer3_outputs[580];
    assign layer4_outputs[1303] = (layer3_outputs[2746]) & ~(layer3_outputs[2818]);
    assign layer4_outputs[1304] = ~(layer3_outputs[2691]);
    assign layer4_outputs[1305] = ~((layer3_outputs[1903]) & (layer3_outputs[3103]));
    assign layer4_outputs[1306] = layer3_outputs[4174];
    assign layer4_outputs[1307] = (layer3_outputs[641]) | (layer3_outputs[2323]);
    assign layer4_outputs[1308] = (layer3_outputs[1292]) & (layer3_outputs[3066]);
    assign layer4_outputs[1309] = layer3_outputs[2926];
    assign layer4_outputs[1310] = layer3_outputs[4529];
    assign layer4_outputs[1311] = (layer3_outputs[3887]) & ~(layer3_outputs[382]);
    assign layer4_outputs[1312] = ~(layer3_outputs[132]);
    assign layer4_outputs[1313] = layer3_outputs[4334];
    assign layer4_outputs[1314] = ~((layer3_outputs[3512]) | (layer3_outputs[3993]));
    assign layer4_outputs[1315] = 1'b1;
    assign layer4_outputs[1316] = layer3_outputs[2473];
    assign layer4_outputs[1317] = ~((layer3_outputs[3232]) ^ (layer3_outputs[2426]));
    assign layer4_outputs[1318] = (layer3_outputs[3723]) & (layer3_outputs[2009]);
    assign layer4_outputs[1319] = layer3_outputs[1604];
    assign layer4_outputs[1320] = layer3_outputs[2969];
    assign layer4_outputs[1321] = layer3_outputs[4263];
    assign layer4_outputs[1322] = 1'b0;
    assign layer4_outputs[1323] = ~(layer3_outputs[383]);
    assign layer4_outputs[1324] = (layer3_outputs[5079]) & (layer3_outputs[3705]);
    assign layer4_outputs[1325] = 1'b1;
    assign layer4_outputs[1326] = (layer3_outputs[2111]) & (layer3_outputs[2966]);
    assign layer4_outputs[1327] = 1'b0;
    assign layer4_outputs[1328] = 1'b1;
    assign layer4_outputs[1329] = ~(layer3_outputs[32]) | (layer3_outputs[998]);
    assign layer4_outputs[1330] = ~(layer3_outputs[2922]);
    assign layer4_outputs[1331] = ~((layer3_outputs[1039]) ^ (layer3_outputs[4329]));
    assign layer4_outputs[1332] = ~(layer3_outputs[1688]) | (layer3_outputs[3709]);
    assign layer4_outputs[1333] = 1'b0;
    assign layer4_outputs[1334] = ~(layer3_outputs[1880]) | (layer3_outputs[3994]);
    assign layer4_outputs[1335] = ~(layer3_outputs[2715]);
    assign layer4_outputs[1336] = 1'b0;
    assign layer4_outputs[1337] = ~((layer3_outputs[597]) | (layer3_outputs[3438]));
    assign layer4_outputs[1338] = ~((layer3_outputs[2343]) | (layer3_outputs[1931]));
    assign layer4_outputs[1339] = ~(layer3_outputs[2608]) | (layer3_outputs[3316]);
    assign layer4_outputs[1340] = (layer3_outputs[786]) & (layer3_outputs[3860]);
    assign layer4_outputs[1341] = layer3_outputs[2763];
    assign layer4_outputs[1342] = (layer3_outputs[2706]) & ~(layer3_outputs[4569]);
    assign layer4_outputs[1343] = 1'b0;
    assign layer4_outputs[1344] = ~(layer3_outputs[4266]);
    assign layer4_outputs[1345] = ~(layer3_outputs[1784]);
    assign layer4_outputs[1346] = layer3_outputs[3732];
    assign layer4_outputs[1347] = layer3_outputs[2425];
    assign layer4_outputs[1348] = layer3_outputs[3469];
    assign layer4_outputs[1349] = ~((layer3_outputs[4226]) ^ (layer3_outputs[113]));
    assign layer4_outputs[1350] = (layer3_outputs[247]) | (layer3_outputs[2450]);
    assign layer4_outputs[1351] = (layer3_outputs[4509]) | (layer3_outputs[213]);
    assign layer4_outputs[1352] = (layer3_outputs[3575]) & ~(layer3_outputs[4868]);
    assign layer4_outputs[1353] = ~((layer3_outputs[618]) & (layer3_outputs[2676]));
    assign layer4_outputs[1354] = (layer3_outputs[903]) | (layer3_outputs[3905]);
    assign layer4_outputs[1355] = (layer3_outputs[1373]) ^ (layer3_outputs[2283]);
    assign layer4_outputs[1356] = layer3_outputs[2258];
    assign layer4_outputs[1357] = layer3_outputs[910];
    assign layer4_outputs[1358] = ~(layer3_outputs[771]);
    assign layer4_outputs[1359] = ~(layer3_outputs[1218]) | (layer3_outputs[3944]);
    assign layer4_outputs[1360] = ~(layer3_outputs[3706]) | (layer3_outputs[2549]);
    assign layer4_outputs[1361] = layer3_outputs[2110];
    assign layer4_outputs[1362] = ~((layer3_outputs[4032]) ^ (layer3_outputs[750]));
    assign layer4_outputs[1363] = ~(layer3_outputs[2235]);
    assign layer4_outputs[1364] = ~(layer3_outputs[3836]);
    assign layer4_outputs[1365] = ~(layer3_outputs[4492]);
    assign layer4_outputs[1366] = ~(layer3_outputs[3392]);
    assign layer4_outputs[1367] = ~(layer3_outputs[1275]) | (layer3_outputs[2433]);
    assign layer4_outputs[1368] = ~(layer3_outputs[2630]) | (layer3_outputs[1120]);
    assign layer4_outputs[1369] = layer3_outputs[4349];
    assign layer4_outputs[1370] = 1'b0;
    assign layer4_outputs[1371] = (layer3_outputs[1150]) & (layer3_outputs[4168]);
    assign layer4_outputs[1372] = ~(layer3_outputs[233]);
    assign layer4_outputs[1373] = layer3_outputs[4610];
    assign layer4_outputs[1374] = ~(layer3_outputs[3932]) | (layer3_outputs[1125]);
    assign layer4_outputs[1375] = ~(layer3_outputs[159]) | (layer3_outputs[1169]);
    assign layer4_outputs[1376] = layer3_outputs[4710];
    assign layer4_outputs[1377] = ~((layer3_outputs[843]) & (layer3_outputs[2800]));
    assign layer4_outputs[1378] = 1'b1;
    assign layer4_outputs[1379] = ~(layer3_outputs[177]) | (layer3_outputs[1402]);
    assign layer4_outputs[1380] = 1'b1;
    assign layer4_outputs[1381] = ~((layer3_outputs[366]) ^ (layer3_outputs[1427]));
    assign layer4_outputs[1382] = (layer3_outputs[4436]) | (layer3_outputs[2351]);
    assign layer4_outputs[1383] = layer3_outputs[3619];
    assign layer4_outputs[1384] = ~(layer3_outputs[1608]);
    assign layer4_outputs[1385] = (layer3_outputs[3125]) & ~(layer3_outputs[2973]);
    assign layer4_outputs[1386] = (layer3_outputs[4204]) ^ (layer3_outputs[3180]);
    assign layer4_outputs[1387] = layer3_outputs[1209];
    assign layer4_outputs[1388] = layer3_outputs[403];
    assign layer4_outputs[1389] = ~(layer3_outputs[4149]);
    assign layer4_outputs[1390] = 1'b0;
    assign layer4_outputs[1391] = layer3_outputs[2089];
    assign layer4_outputs[1392] = ~((layer3_outputs[1299]) | (layer3_outputs[3758]));
    assign layer4_outputs[1393] = ~(layer3_outputs[1620]);
    assign layer4_outputs[1394] = (layer3_outputs[3225]) & ~(layer3_outputs[2670]);
    assign layer4_outputs[1395] = ~(layer3_outputs[3026]);
    assign layer4_outputs[1396] = ~(layer3_outputs[416]);
    assign layer4_outputs[1397] = ~((layer3_outputs[1184]) & (layer3_outputs[4654]));
    assign layer4_outputs[1398] = 1'b1;
    assign layer4_outputs[1399] = layer3_outputs[4076];
    assign layer4_outputs[1400] = layer3_outputs[4695];
    assign layer4_outputs[1401] = ~(layer3_outputs[1271]);
    assign layer4_outputs[1402] = 1'b1;
    assign layer4_outputs[1403] = ~((layer3_outputs[3358]) & (layer3_outputs[3450]));
    assign layer4_outputs[1404] = 1'b0;
    assign layer4_outputs[1405] = ~(layer3_outputs[3835]);
    assign layer4_outputs[1406] = ~(layer3_outputs[4400]) | (layer3_outputs[1757]);
    assign layer4_outputs[1407] = (layer3_outputs[3461]) & (layer3_outputs[3678]);
    assign layer4_outputs[1408] = layer3_outputs[1777];
    assign layer4_outputs[1409] = ~(layer3_outputs[4748]);
    assign layer4_outputs[1410] = ~(layer3_outputs[3597]);
    assign layer4_outputs[1411] = ~((layer3_outputs[4143]) | (layer3_outputs[434]));
    assign layer4_outputs[1412] = (layer3_outputs[4091]) & ~(layer3_outputs[4478]);
    assign layer4_outputs[1413] = ~(layer3_outputs[4845]) | (layer3_outputs[3762]);
    assign layer4_outputs[1414] = layer3_outputs[2753];
    assign layer4_outputs[1415] = ~(layer3_outputs[502]);
    assign layer4_outputs[1416] = layer3_outputs[1758];
    assign layer4_outputs[1417] = ~(layer3_outputs[509]);
    assign layer4_outputs[1418] = (layer3_outputs[1538]) & ~(layer3_outputs[462]);
    assign layer4_outputs[1419] = (layer3_outputs[1040]) & (layer3_outputs[1891]);
    assign layer4_outputs[1420] = ~((layer3_outputs[3364]) & (layer3_outputs[2175]));
    assign layer4_outputs[1421] = ~((layer3_outputs[456]) & (layer3_outputs[284]));
    assign layer4_outputs[1422] = 1'b1;
    assign layer4_outputs[1423] = ~((layer3_outputs[1859]) & (layer3_outputs[1521]));
    assign layer4_outputs[1424] = ~((layer3_outputs[251]) | (layer3_outputs[806]));
    assign layer4_outputs[1425] = ~(layer3_outputs[2236]) | (layer3_outputs[4284]);
    assign layer4_outputs[1426] = ~((layer3_outputs[3266]) | (layer3_outputs[2226]));
    assign layer4_outputs[1427] = 1'b0;
    assign layer4_outputs[1428] = ~((layer3_outputs[4894]) & (layer3_outputs[4317]));
    assign layer4_outputs[1429] = 1'b0;
    assign layer4_outputs[1430] = (layer3_outputs[753]) & ~(layer3_outputs[3483]);
    assign layer4_outputs[1431] = (layer3_outputs[2047]) & ~(layer3_outputs[2052]);
    assign layer4_outputs[1432] = ~(layer3_outputs[3159]);
    assign layer4_outputs[1433] = layer3_outputs[2830];
    assign layer4_outputs[1434] = layer3_outputs[1044];
    assign layer4_outputs[1435] = ~(layer3_outputs[1241]) | (layer3_outputs[3029]);
    assign layer4_outputs[1436] = layer3_outputs[3767];
    assign layer4_outputs[1437] = (layer3_outputs[887]) & (layer3_outputs[2987]);
    assign layer4_outputs[1438] = (layer3_outputs[3497]) & ~(layer3_outputs[3240]);
    assign layer4_outputs[1439] = ~(layer3_outputs[3821]);
    assign layer4_outputs[1440] = ~((layer3_outputs[336]) | (layer3_outputs[1661]));
    assign layer4_outputs[1441] = ~((layer3_outputs[2326]) ^ (layer3_outputs[541]));
    assign layer4_outputs[1442] = layer3_outputs[319];
    assign layer4_outputs[1443] = (layer3_outputs[625]) ^ (layer3_outputs[2115]);
    assign layer4_outputs[1444] = ~(layer3_outputs[594]);
    assign layer4_outputs[1445] = (layer3_outputs[4460]) & (layer3_outputs[3570]);
    assign layer4_outputs[1446] = ~(layer3_outputs[2126]) | (layer3_outputs[4862]);
    assign layer4_outputs[1447] = ~(layer3_outputs[3011]) | (layer3_outputs[2051]);
    assign layer4_outputs[1448] = layer3_outputs[1409];
    assign layer4_outputs[1449] = ~(layer3_outputs[3126]);
    assign layer4_outputs[1450] = ~(layer3_outputs[3121]);
    assign layer4_outputs[1451] = layer3_outputs[1805];
    assign layer4_outputs[1452] = layer3_outputs[264];
    assign layer4_outputs[1453] = layer3_outputs[4153];
    assign layer4_outputs[1454] = ~(layer3_outputs[2186]);
    assign layer4_outputs[1455] = (layer3_outputs[2292]) & ~(layer3_outputs[3296]);
    assign layer4_outputs[1456] = ~(layer3_outputs[4309]);
    assign layer4_outputs[1457] = ~(layer3_outputs[943]);
    assign layer4_outputs[1458] = (layer3_outputs[3393]) & (layer3_outputs[4777]);
    assign layer4_outputs[1459] = layer3_outputs[476];
    assign layer4_outputs[1460] = ~(layer3_outputs[3254]) | (layer3_outputs[902]);
    assign layer4_outputs[1461] = (layer3_outputs[2895]) & ~(layer3_outputs[2664]);
    assign layer4_outputs[1462] = (layer3_outputs[2330]) & ~(layer3_outputs[389]);
    assign layer4_outputs[1463] = 1'b0;
    assign layer4_outputs[1464] = ~(layer3_outputs[2444]);
    assign layer4_outputs[1465] = ~(layer3_outputs[2173]);
    assign layer4_outputs[1466] = ~(layer3_outputs[774]);
    assign layer4_outputs[1467] = (layer3_outputs[4784]) & (layer3_outputs[4267]);
    assign layer4_outputs[1468] = 1'b0;
    assign layer4_outputs[1469] = ~((layer3_outputs[609]) ^ (layer3_outputs[245]));
    assign layer4_outputs[1470] = layer3_outputs[1705];
    assign layer4_outputs[1471] = (layer3_outputs[3060]) & ~(layer3_outputs[3103]);
    assign layer4_outputs[1472] = ~((layer3_outputs[1560]) | (layer3_outputs[737]));
    assign layer4_outputs[1473] = ~(layer3_outputs[4006]);
    assign layer4_outputs[1474] = ~(layer3_outputs[522]);
    assign layer4_outputs[1475] = ~((layer3_outputs[3416]) | (layer3_outputs[524]));
    assign layer4_outputs[1476] = (layer3_outputs[4604]) & ~(layer3_outputs[1839]);
    assign layer4_outputs[1477] = (layer3_outputs[91]) & ~(layer3_outputs[3422]);
    assign layer4_outputs[1478] = (layer3_outputs[1914]) & (layer3_outputs[3459]);
    assign layer4_outputs[1479] = (layer3_outputs[3061]) & (layer3_outputs[2724]);
    assign layer4_outputs[1480] = ~((layer3_outputs[4285]) & (layer3_outputs[3194]));
    assign layer4_outputs[1481] = ~(layer3_outputs[1207]) | (layer3_outputs[3029]);
    assign layer4_outputs[1482] = (layer3_outputs[2527]) & (layer3_outputs[3361]);
    assign layer4_outputs[1483] = ~((layer3_outputs[1522]) ^ (layer3_outputs[4066]));
    assign layer4_outputs[1484] = (layer3_outputs[2840]) & ~(layer3_outputs[1265]);
    assign layer4_outputs[1485] = layer3_outputs[1671];
    assign layer4_outputs[1486] = layer3_outputs[344];
    assign layer4_outputs[1487] = ~(layer3_outputs[5015]);
    assign layer4_outputs[1488] = ~((layer3_outputs[918]) | (layer3_outputs[4242]));
    assign layer4_outputs[1489] = ~(layer3_outputs[956]);
    assign layer4_outputs[1490] = layer3_outputs[2299];
    assign layer4_outputs[1491] = 1'b1;
    assign layer4_outputs[1492] = ~(layer3_outputs[726]);
    assign layer4_outputs[1493] = ~(layer3_outputs[4054]);
    assign layer4_outputs[1494] = (layer3_outputs[1273]) & (layer3_outputs[4691]);
    assign layer4_outputs[1495] = 1'b1;
    assign layer4_outputs[1496] = ~(layer3_outputs[4768]) | (layer3_outputs[3410]);
    assign layer4_outputs[1497] = ~(layer3_outputs[1659]) | (layer3_outputs[2922]);
    assign layer4_outputs[1498] = ~((layer3_outputs[1295]) ^ (layer3_outputs[3867]));
    assign layer4_outputs[1499] = (layer3_outputs[1527]) & ~(layer3_outputs[4487]);
    assign layer4_outputs[1500] = (layer3_outputs[4101]) | (layer3_outputs[4950]);
    assign layer4_outputs[1501] = ~(layer3_outputs[4361]) | (layer3_outputs[3334]);
    assign layer4_outputs[1502] = (layer3_outputs[4499]) | (layer3_outputs[631]);
    assign layer4_outputs[1503] = ~(layer3_outputs[1551]) | (layer3_outputs[2937]);
    assign layer4_outputs[1504] = layer3_outputs[3464];
    assign layer4_outputs[1505] = (layer3_outputs[825]) | (layer3_outputs[770]);
    assign layer4_outputs[1506] = ~((layer3_outputs[2669]) & (layer3_outputs[921]));
    assign layer4_outputs[1507] = ~((layer3_outputs[2532]) & (layer3_outputs[866]));
    assign layer4_outputs[1508] = 1'b0;
    assign layer4_outputs[1509] = ~(layer3_outputs[4458]) | (layer3_outputs[555]);
    assign layer4_outputs[1510] = layer3_outputs[4170];
    assign layer4_outputs[1511] = ~(layer3_outputs[3104]);
    assign layer4_outputs[1512] = (layer3_outputs[187]) ^ (layer3_outputs[2005]);
    assign layer4_outputs[1513] = ~(layer3_outputs[4686]);
    assign layer4_outputs[1514] = layer3_outputs[4079];
    assign layer4_outputs[1515] = (layer3_outputs[411]) & ~(layer3_outputs[2412]);
    assign layer4_outputs[1516] = layer3_outputs[3606];
    assign layer4_outputs[1517] = 1'b1;
    assign layer4_outputs[1518] = layer3_outputs[3460];
    assign layer4_outputs[1519] = layer3_outputs[4295];
    assign layer4_outputs[1520] = 1'b0;
    assign layer4_outputs[1521] = ~(layer3_outputs[4532]) | (layer3_outputs[1408]);
    assign layer4_outputs[1522] = ~(layer3_outputs[328]);
    assign layer4_outputs[1523] = (layer3_outputs[1120]) & ~(layer3_outputs[2961]);
    assign layer4_outputs[1524] = ~((layer3_outputs[543]) & (layer3_outputs[325]));
    assign layer4_outputs[1525] = layer3_outputs[4082];
    assign layer4_outputs[1526] = ~(layer3_outputs[4169]);
    assign layer4_outputs[1527] = ~(layer3_outputs[3538]) | (layer3_outputs[2929]);
    assign layer4_outputs[1528] = 1'b0;
    assign layer4_outputs[1529] = ~(layer3_outputs[1140]);
    assign layer4_outputs[1530] = ~((layer3_outputs[2644]) ^ (layer3_outputs[2626]));
    assign layer4_outputs[1531] = ~(layer3_outputs[3380]);
    assign layer4_outputs[1532] = (layer3_outputs[1312]) & ~(layer3_outputs[1706]);
    assign layer4_outputs[1533] = (layer3_outputs[1271]) & ~(layer3_outputs[1469]);
    assign layer4_outputs[1534] = layer3_outputs[3891];
    assign layer4_outputs[1535] = ~(layer3_outputs[3344]);
    assign layer4_outputs[1536] = ~(layer3_outputs[4536]);
    assign layer4_outputs[1537] = ~(layer3_outputs[1887]);
    assign layer4_outputs[1538] = layer3_outputs[3825];
    assign layer4_outputs[1539] = ~(layer3_outputs[1802]);
    assign layer4_outputs[1540] = (layer3_outputs[1897]) & ~(layer3_outputs[4477]);
    assign layer4_outputs[1541] = 1'b0;
    assign layer4_outputs[1542] = (layer3_outputs[3596]) & (layer3_outputs[2377]);
    assign layer4_outputs[1543] = layer3_outputs[689];
    assign layer4_outputs[1544] = 1'b1;
    assign layer4_outputs[1545] = ~(layer3_outputs[969]);
    assign layer4_outputs[1546] = (layer3_outputs[527]) ^ (layer3_outputs[97]);
    assign layer4_outputs[1547] = ~(layer3_outputs[1980]);
    assign layer4_outputs[1548] = ~(layer3_outputs[157]) | (layer3_outputs[2368]);
    assign layer4_outputs[1549] = ~(layer3_outputs[3146]);
    assign layer4_outputs[1550] = layer3_outputs[841];
    assign layer4_outputs[1551] = layer3_outputs[343];
    assign layer4_outputs[1552] = ~(layer3_outputs[2375]) | (layer3_outputs[2095]);
    assign layer4_outputs[1553] = layer3_outputs[2701];
    assign layer4_outputs[1554] = ~(layer3_outputs[3249]);
    assign layer4_outputs[1555] = (layer3_outputs[4879]) | (layer3_outputs[1543]);
    assign layer4_outputs[1556] = (layer3_outputs[2749]) & (layer3_outputs[292]);
    assign layer4_outputs[1557] = 1'b1;
    assign layer4_outputs[1558] = ~(layer3_outputs[2667]);
    assign layer4_outputs[1559] = ~(layer3_outputs[1892]);
    assign layer4_outputs[1560] = ~(layer3_outputs[1969]);
    assign layer4_outputs[1561] = 1'b0;
    assign layer4_outputs[1562] = (layer3_outputs[740]) ^ (layer3_outputs[2674]);
    assign layer4_outputs[1563] = (layer3_outputs[3098]) & ~(layer3_outputs[1516]);
    assign layer4_outputs[1564] = layer3_outputs[811];
    assign layer4_outputs[1565] = ~((layer3_outputs[849]) | (layer3_outputs[4224]));
    assign layer4_outputs[1566] = (layer3_outputs[3601]) & ~(layer3_outputs[744]);
    assign layer4_outputs[1567] = ~((layer3_outputs[4619]) | (layer3_outputs[2744]));
    assign layer4_outputs[1568] = (layer3_outputs[2768]) & (layer3_outputs[4474]);
    assign layer4_outputs[1569] = (layer3_outputs[2141]) & ~(layer3_outputs[3065]);
    assign layer4_outputs[1570] = ~((layer3_outputs[1245]) & (layer3_outputs[3425]));
    assign layer4_outputs[1571] = layer3_outputs[2984];
    assign layer4_outputs[1572] = ~((layer3_outputs[3174]) ^ (layer3_outputs[3581]));
    assign layer4_outputs[1573] = ~(layer3_outputs[1761]);
    assign layer4_outputs[1574] = 1'b0;
    assign layer4_outputs[1575] = ~(layer3_outputs[2732]);
    assign layer4_outputs[1576] = layer3_outputs[3159];
    assign layer4_outputs[1577] = ~((layer3_outputs[4322]) | (layer3_outputs[4489]));
    assign layer4_outputs[1578] = layer3_outputs[573];
    assign layer4_outputs[1579] = layer3_outputs[3373];
    assign layer4_outputs[1580] = ~((layer3_outputs[4397]) ^ (layer3_outputs[2583]));
    assign layer4_outputs[1581] = 1'b1;
    assign layer4_outputs[1582] = (layer3_outputs[1355]) & ~(layer3_outputs[1140]);
    assign layer4_outputs[1583] = ~((layer3_outputs[1457]) | (layer3_outputs[3454]));
    assign layer4_outputs[1584] = ~(layer3_outputs[2206]);
    assign layer4_outputs[1585] = ~(layer3_outputs[4399]) | (layer3_outputs[1974]);
    assign layer4_outputs[1586] = (layer3_outputs[43]) & ~(layer3_outputs[179]);
    assign layer4_outputs[1587] = (layer3_outputs[2471]) ^ (layer3_outputs[5042]);
    assign layer4_outputs[1588] = (layer3_outputs[2209]) & ~(layer3_outputs[2743]);
    assign layer4_outputs[1589] = (layer3_outputs[3696]) & (layer3_outputs[3863]);
    assign layer4_outputs[1590] = (layer3_outputs[337]) & ~(layer3_outputs[841]);
    assign layer4_outputs[1591] = layer3_outputs[3059];
    assign layer4_outputs[1592] = ~(layer3_outputs[2404]);
    assign layer4_outputs[1593] = layer3_outputs[766];
    assign layer4_outputs[1594] = ~(layer3_outputs[1694]) | (layer3_outputs[4931]);
    assign layer4_outputs[1595] = (layer3_outputs[2586]) & ~(layer3_outputs[1370]);
    assign layer4_outputs[1596] = layer3_outputs[1156];
    assign layer4_outputs[1597] = 1'b0;
    assign layer4_outputs[1598] = ~(layer3_outputs[4893]);
    assign layer4_outputs[1599] = layer3_outputs[4451];
    assign layer4_outputs[1600] = layer3_outputs[1829];
    assign layer4_outputs[1601] = ~(layer3_outputs[3066]);
    assign layer4_outputs[1602] = (layer3_outputs[669]) & ~(layer3_outputs[802]);
    assign layer4_outputs[1603] = ~(layer3_outputs[2349]) | (layer3_outputs[955]);
    assign layer4_outputs[1604] = layer3_outputs[3637];
    assign layer4_outputs[1605] = ~(layer3_outputs[4938]);
    assign layer4_outputs[1606] = 1'b1;
    assign layer4_outputs[1607] = (layer3_outputs[5035]) & ~(layer3_outputs[489]);
    assign layer4_outputs[1608] = ~((layer3_outputs[351]) & (layer3_outputs[2222]));
    assign layer4_outputs[1609] = ~(layer3_outputs[2454]);
    assign layer4_outputs[1610] = layer3_outputs[3781];
    assign layer4_outputs[1611] = ~((layer3_outputs[1607]) & (layer3_outputs[1342]));
    assign layer4_outputs[1612] = ~(layer3_outputs[653]);
    assign layer4_outputs[1613] = (layer3_outputs[3409]) | (layer3_outputs[3120]);
    assign layer4_outputs[1614] = (layer3_outputs[3440]) & (layer3_outputs[4473]);
    assign layer4_outputs[1615] = layer3_outputs[4296];
    assign layer4_outputs[1616] = ~(layer3_outputs[4636]);
    assign layer4_outputs[1617] = ~(layer3_outputs[2116]);
    assign layer4_outputs[1618] = ~((layer3_outputs[3950]) | (layer3_outputs[4453]));
    assign layer4_outputs[1619] = ~(layer3_outputs[1297]);
    assign layer4_outputs[1620] = 1'b0;
    assign layer4_outputs[1621] = ~(layer3_outputs[426]);
    assign layer4_outputs[1622] = (layer3_outputs[2712]) & ~(layer3_outputs[10]);
    assign layer4_outputs[1623] = 1'b1;
    assign layer4_outputs[1624] = ~(layer3_outputs[318]) | (layer3_outputs[689]);
    assign layer4_outputs[1625] = layer3_outputs[4885];
    assign layer4_outputs[1626] = (layer3_outputs[1701]) & ~(layer3_outputs[1874]);
    assign layer4_outputs[1627] = ~(layer3_outputs[40]);
    assign layer4_outputs[1628] = ~(layer3_outputs[1462]);
    assign layer4_outputs[1629] = (layer3_outputs[1841]) & (layer3_outputs[1807]);
    assign layer4_outputs[1630] = layer3_outputs[4793];
    assign layer4_outputs[1631] = ~(layer3_outputs[713]) | (layer3_outputs[3765]);
    assign layer4_outputs[1632] = layer3_outputs[1284];
    assign layer4_outputs[1633] = ~((layer3_outputs[3499]) ^ (layer3_outputs[4027]));
    assign layer4_outputs[1634] = ~(layer3_outputs[33]) | (layer3_outputs[1203]);
    assign layer4_outputs[1635] = (layer3_outputs[1252]) & (layer3_outputs[259]);
    assign layer4_outputs[1636] = (layer3_outputs[1714]) & (layer3_outputs[5049]);
    assign layer4_outputs[1637] = (layer3_outputs[2920]) & ~(layer3_outputs[1298]);
    assign layer4_outputs[1638] = layer3_outputs[4593];
    assign layer4_outputs[1639] = layer3_outputs[4536];
    assign layer4_outputs[1640] = ~(layer3_outputs[2240]);
    assign layer4_outputs[1641] = layer3_outputs[739];
    assign layer4_outputs[1642] = ~(layer3_outputs[410]);
    assign layer4_outputs[1643] = layer3_outputs[1611];
    assign layer4_outputs[1644] = ~(layer3_outputs[655]) | (layer3_outputs[798]);
    assign layer4_outputs[1645] = layer3_outputs[1393];
    assign layer4_outputs[1646] = ~((layer3_outputs[5078]) | (layer3_outputs[3996]));
    assign layer4_outputs[1647] = layer3_outputs[2496];
    assign layer4_outputs[1648] = 1'b0;
    assign layer4_outputs[1649] = layer3_outputs[3799];
    assign layer4_outputs[1650] = layer3_outputs[408];
    assign layer4_outputs[1651] = 1'b1;
    assign layer4_outputs[1652] = (layer3_outputs[2967]) & ~(layer3_outputs[2651]);
    assign layer4_outputs[1653] = ~((layer3_outputs[1637]) | (layer3_outputs[3383]));
    assign layer4_outputs[1654] = ~((layer3_outputs[688]) | (layer3_outputs[3195]));
    assign layer4_outputs[1655] = ~(layer3_outputs[679]) | (layer3_outputs[1545]);
    assign layer4_outputs[1656] = ~((layer3_outputs[296]) ^ (layer3_outputs[35]));
    assign layer4_outputs[1657] = layer3_outputs[1832];
    assign layer4_outputs[1658] = layer3_outputs[23];
    assign layer4_outputs[1659] = 1'b1;
    assign layer4_outputs[1660] = ~(layer3_outputs[1552]);
    assign layer4_outputs[1661] = (layer3_outputs[212]) ^ (layer3_outputs[2968]);
    assign layer4_outputs[1662] = ~(layer3_outputs[2924]) | (layer3_outputs[3998]);
    assign layer4_outputs[1663] = ~((layer3_outputs[3603]) ^ (layer3_outputs[1693]));
    assign layer4_outputs[1664] = ~((layer3_outputs[5044]) | (layer3_outputs[4757]));
    assign layer4_outputs[1665] = ~((layer3_outputs[1574]) & (layer3_outputs[4853]));
    assign layer4_outputs[1666] = layer3_outputs[2662];
    assign layer4_outputs[1667] = (layer3_outputs[1494]) & ~(layer3_outputs[4697]);
    assign layer4_outputs[1668] = (layer3_outputs[2430]) & ~(layer3_outputs[2635]);
    assign layer4_outputs[1669] = layer3_outputs[728];
    assign layer4_outputs[1670] = (layer3_outputs[3247]) ^ (layer3_outputs[3866]);
    assign layer4_outputs[1671] = ~(layer3_outputs[1683]);
    assign layer4_outputs[1672] = layer3_outputs[2653];
    assign layer4_outputs[1673] = 1'b0;
    assign layer4_outputs[1674] = ~(layer3_outputs[3182]) | (layer3_outputs[4812]);
    assign layer4_outputs[1675] = ~((layer3_outputs[2513]) ^ (layer3_outputs[3871]));
    assign layer4_outputs[1676] = ~(layer3_outputs[1342]);
    assign layer4_outputs[1677] = layer3_outputs[1221];
    assign layer4_outputs[1678] = layer3_outputs[2698];
    assign layer4_outputs[1679] = (layer3_outputs[1703]) & ~(layer3_outputs[4012]);
    assign layer4_outputs[1680] = ~((layer3_outputs[1834]) | (layer3_outputs[2799]));
    assign layer4_outputs[1681] = layer3_outputs[2268];
    assign layer4_outputs[1682] = ~(layer3_outputs[1267]);
    assign layer4_outputs[1683] = (layer3_outputs[2381]) & ~(layer3_outputs[4304]);
    assign layer4_outputs[1684] = (layer3_outputs[2275]) & ~(layer3_outputs[1153]);
    assign layer4_outputs[1685] = layer3_outputs[2864];
    assign layer4_outputs[1686] = ~(layer3_outputs[3604]) | (layer3_outputs[4999]);
    assign layer4_outputs[1687] = ~(layer3_outputs[2231]);
    assign layer4_outputs[1688] = ~(layer3_outputs[2615]);
    assign layer4_outputs[1689] = ~((layer3_outputs[1809]) & (layer3_outputs[430]));
    assign layer4_outputs[1690] = layer3_outputs[4437];
    assign layer4_outputs[1691] = (layer3_outputs[2392]) & (layer3_outputs[649]);
    assign layer4_outputs[1692] = ~(layer3_outputs[4352]);
    assign layer4_outputs[1693] = (layer3_outputs[216]) | (layer3_outputs[1723]);
    assign layer4_outputs[1694] = (layer3_outputs[2358]) | (layer3_outputs[2403]);
    assign layer4_outputs[1695] = layer3_outputs[2366];
    assign layer4_outputs[1696] = (layer3_outputs[3804]) & ~(layer3_outputs[2094]);
    assign layer4_outputs[1697] = (layer3_outputs[2950]) & ~(layer3_outputs[970]);
    assign layer4_outputs[1698] = (layer3_outputs[2935]) & (layer3_outputs[2018]);
    assign layer4_outputs[1699] = ~(layer3_outputs[1594]);
    assign layer4_outputs[1700] = (layer3_outputs[2618]) ^ (layer3_outputs[2910]);
    assign layer4_outputs[1701] = (layer3_outputs[4667]) & ~(layer3_outputs[2996]);
    assign layer4_outputs[1702] = (layer3_outputs[2902]) ^ (layer3_outputs[3601]);
    assign layer4_outputs[1703] = ~(layer3_outputs[3241]);
    assign layer4_outputs[1704] = layer3_outputs[2481];
    assign layer4_outputs[1705] = 1'b0;
    assign layer4_outputs[1706] = ~(layer3_outputs[4144]);
    assign layer4_outputs[1707] = ~(layer3_outputs[50]);
    assign layer4_outputs[1708] = ~(layer3_outputs[2140]);
    assign layer4_outputs[1709] = ~(layer3_outputs[293]) | (layer3_outputs[2494]);
    assign layer4_outputs[1710] = ~(layer3_outputs[370]);
    assign layer4_outputs[1711] = ~(layer3_outputs[1886]);
    assign layer4_outputs[1712] = ~(layer3_outputs[4075]);
    assign layer4_outputs[1713] = (layer3_outputs[3531]) & (layer3_outputs[4664]);
    assign layer4_outputs[1714] = layer3_outputs[2032];
    assign layer4_outputs[1715] = (layer3_outputs[3887]) | (layer3_outputs[577]);
    assign layer4_outputs[1716] = ~((layer3_outputs[2594]) ^ (layer3_outputs[2051]));
    assign layer4_outputs[1717] = ~(layer3_outputs[1838]);
    assign layer4_outputs[1718] = layer3_outputs[57];
    assign layer4_outputs[1719] = ~(layer3_outputs[926]);
    assign layer4_outputs[1720] = layer3_outputs[1396];
    assign layer4_outputs[1721] = ~(layer3_outputs[3424]) | (layer3_outputs[360]);
    assign layer4_outputs[1722] = ~((layer3_outputs[4146]) & (layer3_outputs[3387]));
    assign layer4_outputs[1723] = layer3_outputs[1723];
    assign layer4_outputs[1724] = (layer3_outputs[3978]) & (layer3_outputs[4614]);
    assign layer4_outputs[1725] = (layer3_outputs[212]) ^ (layer3_outputs[2878]);
    assign layer4_outputs[1726] = ~(layer3_outputs[3145]);
    assign layer4_outputs[1727] = ~(layer3_outputs[3162]) | (layer3_outputs[513]);
    assign layer4_outputs[1728] = (layer3_outputs[1779]) & (layer3_outputs[2563]);
    assign layer4_outputs[1729] = (layer3_outputs[512]) & (layer3_outputs[2423]);
    assign layer4_outputs[1730] = ~(layer3_outputs[859]);
    assign layer4_outputs[1731] = (layer3_outputs[4717]) & ~(layer3_outputs[3328]);
    assign layer4_outputs[1732] = layer3_outputs[3461];
    assign layer4_outputs[1733] = ~(layer3_outputs[566]) | (layer3_outputs[3415]);
    assign layer4_outputs[1734] = layer3_outputs[1163];
    assign layer4_outputs[1735] = ~(layer3_outputs[5083]);
    assign layer4_outputs[1736] = ~(layer3_outputs[1076]);
    assign layer4_outputs[1737] = ~((layer3_outputs[3341]) | (layer3_outputs[4362]));
    assign layer4_outputs[1738] = layer3_outputs[4826];
    assign layer4_outputs[1739] = ~((layer3_outputs[4082]) ^ (layer3_outputs[376]));
    assign layer4_outputs[1740] = ~((layer3_outputs[1756]) | (layer3_outputs[3288]));
    assign layer4_outputs[1741] = ~(layer3_outputs[2236]);
    assign layer4_outputs[1742] = ~((layer3_outputs[1460]) & (layer3_outputs[3238]));
    assign layer4_outputs[1743] = (layer3_outputs[1948]) & ~(layer3_outputs[4438]);
    assign layer4_outputs[1744] = 1'b1;
    assign layer4_outputs[1745] = 1'b0;
    assign layer4_outputs[1746] = ~(layer3_outputs[4926]);
    assign layer4_outputs[1747] = ~((layer3_outputs[2851]) & (layer3_outputs[5005]));
    assign layer4_outputs[1748] = layer3_outputs[1501];
    assign layer4_outputs[1749] = ~(layer3_outputs[3761]);
    assign layer4_outputs[1750] = ~((layer3_outputs[4809]) | (layer3_outputs[2428]));
    assign layer4_outputs[1751] = 1'b1;
    assign layer4_outputs[1752] = ~(layer3_outputs[1340]);
    assign layer4_outputs[1753] = (layer3_outputs[3292]) | (layer3_outputs[772]);
    assign layer4_outputs[1754] = 1'b0;
    assign layer4_outputs[1755] = ~(layer3_outputs[3912]);
    assign layer4_outputs[1756] = ~(layer3_outputs[4167]);
    assign layer4_outputs[1757] = layer3_outputs[2478];
    assign layer4_outputs[1758] = (layer3_outputs[3654]) ^ (layer3_outputs[2365]);
    assign layer4_outputs[1759] = layer3_outputs[3418];
    assign layer4_outputs[1760] = ~(layer3_outputs[1247]);
    assign layer4_outputs[1761] = layer3_outputs[4159];
    assign layer4_outputs[1762] = (layer3_outputs[163]) & (layer3_outputs[4631]);
    assign layer4_outputs[1763] = layer3_outputs[4618];
    assign layer4_outputs[1764] = ~(layer3_outputs[1537]);
    assign layer4_outputs[1765] = layer3_outputs[2273];
    assign layer4_outputs[1766] = (layer3_outputs[1616]) & (layer3_outputs[3437]);
    assign layer4_outputs[1767] = (layer3_outputs[2668]) & ~(layer3_outputs[4843]);
    assign layer4_outputs[1768] = ~(layer3_outputs[764]) | (layer3_outputs[254]);
    assign layer4_outputs[1769] = layer3_outputs[748];
    assign layer4_outputs[1770] = ~((layer3_outputs[4572]) ^ (layer3_outputs[524]));
    assign layer4_outputs[1771] = (layer3_outputs[1912]) & ~(layer3_outputs[1063]);
    assign layer4_outputs[1772] = ~(layer3_outputs[4835]);
    assign layer4_outputs[1773] = layer3_outputs[2259];
    assign layer4_outputs[1774] = ~(layer3_outputs[3566]) | (layer3_outputs[4535]);
    assign layer4_outputs[1775] = (layer3_outputs[3692]) ^ (layer3_outputs[1068]);
    assign layer4_outputs[1776] = ~((layer3_outputs[4396]) | (layer3_outputs[2785]));
    assign layer4_outputs[1777] = ~(layer3_outputs[2588]);
    assign layer4_outputs[1778] = 1'b0;
    assign layer4_outputs[1779] = layer3_outputs[2969];
    assign layer4_outputs[1780] = ~((layer3_outputs[1205]) ^ (layer3_outputs[5006]));
    assign layer4_outputs[1781] = 1'b0;
    assign layer4_outputs[1782] = (layer3_outputs[135]) & ~(layer3_outputs[1464]);
    assign layer4_outputs[1783] = layer3_outputs[3770];
    assign layer4_outputs[1784] = 1'b1;
    assign layer4_outputs[1785] = 1'b1;
    assign layer4_outputs[1786] = ~(layer3_outputs[1103]) | (layer3_outputs[2874]);
    assign layer4_outputs[1787] = ~(layer3_outputs[4479]);
    assign layer4_outputs[1788] = (layer3_outputs[1204]) ^ (layer3_outputs[217]);
    assign layer4_outputs[1789] = ~(layer3_outputs[620]);
    assign layer4_outputs[1790] = layer3_outputs[2999];
    assign layer4_outputs[1791] = layer3_outputs[700];
    assign layer4_outputs[1792] = (layer3_outputs[636]) & ~(layer3_outputs[4376]);
    assign layer4_outputs[1793] = (layer3_outputs[4213]) & (layer3_outputs[3407]);
    assign layer4_outputs[1794] = ~(layer3_outputs[2187]) | (layer3_outputs[185]);
    assign layer4_outputs[1795] = ~((layer3_outputs[66]) | (layer3_outputs[4605]));
    assign layer4_outputs[1796] = layer3_outputs[4018];
    assign layer4_outputs[1797] = ~(layer3_outputs[2456]);
    assign layer4_outputs[1798] = ~((layer3_outputs[136]) & (layer3_outputs[1947]));
    assign layer4_outputs[1799] = 1'b1;
    assign layer4_outputs[1800] = 1'b0;
    assign layer4_outputs[1801] = (layer3_outputs[4621]) & (layer3_outputs[4549]);
    assign layer4_outputs[1802] = ~((layer3_outputs[3848]) | (layer3_outputs[4972]));
    assign layer4_outputs[1803] = (layer3_outputs[3000]) & (layer3_outputs[4670]);
    assign layer4_outputs[1804] = layer3_outputs[93];
    assign layer4_outputs[1805] = (layer3_outputs[4113]) & ~(layer3_outputs[1335]);
    assign layer4_outputs[1806] = layer3_outputs[4192];
    assign layer4_outputs[1807] = ~(layer3_outputs[2127]);
    assign layer4_outputs[1808] = ~(layer3_outputs[328]) | (layer3_outputs[1229]);
    assign layer4_outputs[1809] = (layer3_outputs[4466]) & ~(layer3_outputs[2316]);
    assign layer4_outputs[1810] = 1'b1;
    assign layer4_outputs[1811] = ~(layer3_outputs[1655]) | (layer3_outputs[2522]);
    assign layer4_outputs[1812] = ~(layer3_outputs[720]);
    assign layer4_outputs[1813] = 1'b0;
    assign layer4_outputs[1814] = ~(layer3_outputs[2219]);
    assign layer4_outputs[1815] = ~(layer3_outputs[4707]) | (layer3_outputs[4377]);
    assign layer4_outputs[1816] = (layer3_outputs[293]) & ~(layer3_outputs[860]);
    assign layer4_outputs[1817] = ~((layer3_outputs[736]) | (layer3_outputs[4832]));
    assign layer4_outputs[1818] = (layer3_outputs[4377]) | (layer3_outputs[5051]);
    assign layer4_outputs[1819] = ~((layer3_outputs[2358]) | (layer3_outputs[1860]));
    assign layer4_outputs[1820] = (layer3_outputs[4959]) ^ (layer3_outputs[1371]);
    assign layer4_outputs[1821] = (layer3_outputs[894]) & (layer3_outputs[454]);
    assign layer4_outputs[1822] = layer3_outputs[2985];
    assign layer4_outputs[1823] = ~(layer3_outputs[4112]);
    assign layer4_outputs[1824] = ~(layer3_outputs[3864]) | (layer3_outputs[402]);
    assign layer4_outputs[1825] = ~((layer3_outputs[4267]) & (layer3_outputs[4411]));
    assign layer4_outputs[1826] = (layer3_outputs[1432]) & ~(layer3_outputs[3134]);
    assign layer4_outputs[1827] = (layer3_outputs[1123]) & (layer3_outputs[1266]);
    assign layer4_outputs[1828] = ~((layer3_outputs[137]) & (layer3_outputs[2714]));
    assign layer4_outputs[1829] = layer3_outputs[5036];
    assign layer4_outputs[1830] = (layer3_outputs[640]) & ~(layer3_outputs[411]);
    assign layer4_outputs[1831] = (layer3_outputs[5010]) & (layer3_outputs[4254]);
    assign layer4_outputs[1832] = 1'b0;
    assign layer4_outputs[1833] = (layer3_outputs[378]) & ~(layer3_outputs[2526]);
    assign layer4_outputs[1834] = layer3_outputs[987];
    assign layer4_outputs[1835] = 1'b1;
    assign layer4_outputs[1836] = 1'b1;
    assign layer4_outputs[1837] = (layer3_outputs[488]) | (layer3_outputs[279]);
    assign layer4_outputs[1838] = (layer3_outputs[5012]) & (layer3_outputs[2144]);
    assign layer4_outputs[1839] = ~((layer3_outputs[2726]) | (layer3_outputs[2997]));
    assign layer4_outputs[1840] = ~(layer3_outputs[1490]) | (layer3_outputs[4828]);
    assign layer4_outputs[1841] = 1'b1;
    assign layer4_outputs[1842] = ~(layer3_outputs[18]);
    assign layer4_outputs[1843] = ~((layer3_outputs[2638]) & (layer3_outputs[1332]));
    assign layer4_outputs[1844] = ~(layer3_outputs[1950]) | (layer3_outputs[648]);
    assign layer4_outputs[1845] = (layer3_outputs[974]) | (layer3_outputs[2633]);
    assign layer4_outputs[1846] = (layer3_outputs[288]) & ~(layer3_outputs[2136]);
    assign layer4_outputs[1847] = ~((layer3_outputs[712]) & (layer3_outputs[3488]));
    assign layer4_outputs[1848] = 1'b1;
    assign layer4_outputs[1849] = ~(layer3_outputs[2580]);
    assign layer4_outputs[1850] = ~(layer3_outputs[2348]);
    assign layer4_outputs[1851] = layer3_outputs[710];
    assign layer4_outputs[1852] = ~(layer3_outputs[4167]);
    assign layer4_outputs[1853] = ~(layer3_outputs[4913]) | (layer3_outputs[3884]);
    assign layer4_outputs[1854] = 1'b0;
    assign layer4_outputs[1855] = ~((layer3_outputs[4974]) & (layer3_outputs[784]));
    assign layer4_outputs[1856] = ~((layer3_outputs[2086]) | (layer3_outputs[2322]));
    assign layer4_outputs[1857] = ~(layer3_outputs[4814]);
    assign layer4_outputs[1858] = 1'b0;
    assign layer4_outputs[1859] = layer3_outputs[5105];
    assign layer4_outputs[1860] = (layer3_outputs[3670]) & ~(layer3_outputs[3046]);
    assign layer4_outputs[1861] = (layer3_outputs[3569]) & ~(layer3_outputs[3990]);
    assign layer4_outputs[1862] = (layer3_outputs[2434]) ^ (layer3_outputs[616]);
    assign layer4_outputs[1863] = ~(layer3_outputs[1136]);
    assign layer4_outputs[1864] = (layer3_outputs[1857]) & ~(layer3_outputs[3054]);
    assign layer4_outputs[1865] = (layer3_outputs[4878]) | (layer3_outputs[2890]);
    assign layer4_outputs[1866] = layer3_outputs[899];
    assign layer4_outputs[1867] = layer3_outputs[2978];
    assign layer4_outputs[1868] = ~(layer3_outputs[1446]);
    assign layer4_outputs[1869] = ~(layer3_outputs[1792]);
    assign layer4_outputs[1870] = (layer3_outputs[1724]) & (layer3_outputs[1070]);
    assign layer4_outputs[1871] = (layer3_outputs[3338]) & (layer3_outputs[1075]);
    assign layer4_outputs[1872] = layer3_outputs[4880];
    assign layer4_outputs[1873] = layer3_outputs[2961];
    assign layer4_outputs[1874] = (layer3_outputs[3005]) & ~(layer3_outputs[461]);
    assign layer4_outputs[1875] = (layer3_outputs[2390]) & ~(layer3_outputs[3181]);
    assign layer4_outputs[1876] = layer3_outputs[868];
    assign layer4_outputs[1877] = layer3_outputs[1039];
    assign layer4_outputs[1878] = ~(layer3_outputs[511]);
    assign layer4_outputs[1879] = (layer3_outputs[1566]) & ~(layer3_outputs[1134]);
    assign layer4_outputs[1880] = ~((layer3_outputs[897]) | (layer3_outputs[1184]));
    assign layer4_outputs[1881] = ~((layer3_outputs[1126]) & (layer3_outputs[4499]));
    assign layer4_outputs[1882] = ~((layer3_outputs[4602]) & (layer3_outputs[897]));
    assign layer4_outputs[1883] = ~(layer3_outputs[1154]) | (layer3_outputs[317]);
    assign layer4_outputs[1884] = 1'b0;
    assign layer4_outputs[1885] = (layer3_outputs[3649]) & ~(layer3_outputs[891]);
    assign layer4_outputs[1886] = layer3_outputs[4454];
    assign layer4_outputs[1887] = ~(layer3_outputs[59]);
    assign layer4_outputs[1888] = ~(layer3_outputs[4869]);
    assign layer4_outputs[1889] = layer3_outputs[1306];
    assign layer4_outputs[1890] = ~((layer3_outputs[895]) | (layer3_outputs[1514]));
    assign layer4_outputs[1891] = ~(layer3_outputs[3649]);
    assign layer4_outputs[1892] = 1'b0;
    assign layer4_outputs[1893] = (layer3_outputs[3016]) ^ (layer3_outputs[1677]);
    assign layer4_outputs[1894] = (layer3_outputs[4440]) | (layer3_outputs[932]);
    assign layer4_outputs[1895] = (layer3_outputs[5070]) | (layer3_outputs[985]);
    assign layer4_outputs[1896] = ~((layer3_outputs[3641]) | (layer3_outputs[4671]));
    assign layer4_outputs[1897] = layer3_outputs[637];
    assign layer4_outputs[1898] = ~(layer3_outputs[4115]);
    assign layer4_outputs[1899] = layer3_outputs[3625];
    assign layer4_outputs[1900] = layer3_outputs[621];
    assign layer4_outputs[1901] = ~(layer3_outputs[4127]);
    assign layer4_outputs[1902] = ~(layer3_outputs[3780]);
    assign layer4_outputs[1903] = 1'b1;
    assign layer4_outputs[1904] = ~(layer3_outputs[1024]);
    assign layer4_outputs[1905] = layer3_outputs[1466];
    assign layer4_outputs[1906] = layer3_outputs[4858];
    assign layer4_outputs[1907] = ~((layer3_outputs[196]) | (layer3_outputs[5116]));
    assign layer4_outputs[1908] = ~(layer3_outputs[3992]);
    assign layer4_outputs[1909] = layer3_outputs[3443];
    assign layer4_outputs[1910] = 1'b1;
    assign layer4_outputs[1911] = ~((layer3_outputs[3547]) ^ (layer3_outputs[4930]));
    assign layer4_outputs[1912] = (layer3_outputs[4334]) & ~(layer3_outputs[98]);
    assign layer4_outputs[1913] = (layer3_outputs[2521]) & ~(layer3_outputs[4776]);
    assign layer4_outputs[1914] = layer3_outputs[63];
    assign layer4_outputs[1915] = ~(layer3_outputs[2121]) | (layer3_outputs[3745]);
    assign layer4_outputs[1916] = ~((layer3_outputs[1697]) ^ (layer3_outputs[2812]));
    assign layer4_outputs[1917] = 1'b1;
    assign layer4_outputs[1918] = 1'b0;
    assign layer4_outputs[1919] = ~(layer3_outputs[2679]);
    assign layer4_outputs[1920] = ~((layer3_outputs[1293]) & (layer3_outputs[4529]));
    assign layer4_outputs[1921] = ~((layer3_outputs[2034]) ^ (layer3_outputs[4674]));
    assign layer4_outputs[1922] = ~((layer3_outputs[1793]) | (layer3_outputs[37]));
    assign layer4_outputs[1923] = (layer3_outputs[1777]) & (layer3_outputs[3296]);
    assign layer4_outputs[1924] = ~(layer3_outputs[2931]) | (layer3_outputs[1802]);
    assign layer4_outputs[1925] = ~(layer3_outputs[4216]);
    assign layer4_outputs[1926] = ~(layer3_outputs[3100]) | (layer3_outputs[4009]);
    assign layer4_outputs[1927] = ~(layer3_outputs[4293]) | (layer3_outputs[2307]);
    assign layer4_outputs[1928] = ~(layer3_outputs[3275]) | (layer3_outputs[3357]);
    assign layer4_outputs[1929] = layer3_outputs[4280];
    assign layer4_outputs[1930] = ~(layer3_outputs[511]);
    assign layer4_outputs[1931] = (layer3_outputs[3467]) & ~(layer3_outputs[2938]);
    assign layer4_outputs[1932] = (layer3_outputs[4392]) & ~(layer3_outputs[1569]);
    assign layer4_outputs[1933] = ~(layer3_outputs[4181]) | (layer3_outputs[3614]);
    assign layer4_outputs[1934] = 1'b1;
    assign layer4_outputs[1935] = (layer3_outputs[3770]) & ~(layer3_outputs[1579]);
    assign layer4_outputs[1936] = layer3_outputs[2422];
    assign layer4_outputs[1937] = ~((layer3_outputs[2553]) & (layer3_outputs[582]));
    assign layer4_outputs[1938] = (layer3_outputs[2584]) & ~(layer3_outputs[1851]);
    assign layer4_outputs[1939] = ~((layer3_outputs[1124]) | (layer3_outputs[4939]));
    assign layer4_outputs[1940] = ~(layer3_outputs[3582]) | (layer3_outputs[2013]);
    assign layer4_outputs[1941] = ~(layer3_outputs[4055]);
    assign layer4_outputs[1942] = 1'b1;
    assign layer4_outputs[1943] = layer3_outputs[3384];
    assign layer4_outputs[1944] = (layer3_outputs[3302]) & ~(layer3_outputs[5093]);
    assign layer4_outputs[1945] = (layer3_outputs[1925]) & ~(layer3_outputs[4427]);
    assign layer4_outputs[1946] = layer3_outputs[4014];
    assign layer4_outputs[1947] = ~(layer3_outputs[3915]);
    assign layer4_outputs[1948] = ~((layer3_outputs[1391]) ^ (layer3_outputs[4389]));
    assign layer4_outputs[1949] = layer3_outputs[1233];
    assign layer4_outputs[1950] = ~(layer3_outputs[3339]);
    assign layer4_outputs[1951] = 1'b0;
    assign layer4_outputs[1952] = (layer3_outputs[4775]) ^ (layer3_outputs[4520]);
    assign layer4_outputs[1953] = ~((layer3_outputs[696]) ^ (layer3_outputs[1309]));
    assign layer4_outputs[1954] = ~((layer3_outputs[24]) ^ (layer3_outputs[6]));
    assign layer4_outputs[1955] = (layer3_outputs[2776]) | (layer3_outputs[3214]);
    assign layer4_outputs[1956] = ~(layer3_outputs[3431]);
    assign layer4_outputs[1957] = layer3_outputs[3514];
    assign layer4_outputs[1958] = layer3_outputs[1244];
    assign layer4_outputs[1959] = (layer3_outputs[3990]) & ~(layer3_outputs[4537]);
    assign layer4_outputs[1960] = 1'b1;
    assign layer4_outputs[1961] = (layer3_outputs[4409]) & ~(layer3_outputs[271]);
    assign layer4_outputs[1962] = ~(layer3_outputs[1849]) | (layer3_outputs[3859]);
    assign layer4_outputs[1963] = ~(layer3_outputs[3533]) | (layer3_outputs[151]);
    assign layer4_outputs[1964] = ~(layer3_outputs[2313]) | (layer3_outputs[3096]);
    assign layer4_outputs[1965] = ~(layer3_outputs[4904]) | (layer3_outputs[4283]);
    assign layer4_outputs[1966] = layer3_outputs[1122];
    assign layer4_outputs[1967] = 1'b0;
    assign layer4_outputs[1968] = ~((layer3_outputs[565]) ^ (layer3_outputs[2460]));
    assign layer4_outputs[1969] = (layer3_outputs[3253]) & ~(layer3_outputs[4033]);
    assign layer4_outputs[1970] = (layer3_outputs[4665]) & ~(layer3_outputs[1828]);
    assign layer4_outputs[1971] = ~((layer3_outputs[2327]) | (layer3_outputs[5092]));
    assign layer4_outputs[1972] = (layer3_outputs[1146]) & ~(layer3_outputs[4985]);
    assign layer4_outputs[1973] = (layer3_outputs[2123]) & ~(layer3_outputs[5061]);
    assign layer4_outputs[1974] = layer3_outputs[3634];
    assign layer4_outputs[1975] = 1'b0;
    assign layer4_outputs[1976] = layer3_outputs[844];
    assign layer4_outputs[1977] = (layer3_outputs[2698]) ^ (layer3_outputs[361]);
    assign layer4_outputs[1978] = ~((layer3_outputs[2599]) & (layer3_outputs[3527]));
    assign layer4_outputs[1979] = ~((layer3_outputs[3327]) & (layer3_outputs[3511]));
    assign layer4_outputs[1980] = (layer3_outputs[1734]) & (layer3_outputs[4319]);
    assign layer4_outputs[1981] = layer3_outputs[4609];
    assign layer4_outputs[1982] = ~(layer3_outputs[3370]) | (layer3_outputs[1917]);
    assign layer4_outputs[1983] = ~((layer3_outputs[2479]) | (layer3_outputs[5039]));
    assign layer4_outputs[1984] = (layer3_outputs[3375]) & ~(layer3_outputs[1459]);
    assign layer4_outputs[1985] = ~(layer3_outputs[3801]);
    assign layer4_outputs[1986] = 1'b0;
    assign layer4_outputs[1987] = ~(layer3_outputs[1093]) | (layer3_outputs[4122]);
    assign layer4_outputs[1988] = layer3_outputs[3222];
    assign layer4_outputs[1989] = layer3_outputs[4538];
    assign layer4_outputs[1990] = ~(layer3_outputs[4866]);
    assign layer4_outputs[1991] = layer3_outputs[1248];
    assign layer4_outputs[1992] = ~(layer3_outputs[5115]);
    assign layer4_outputs[1993] = ~(layer3_outputs[4399]);
    assign layer4_outputs[1994] = layer3_outputs[4681];
    assign layer4_outputs[1995] = ~((layer3_outputs[2149]) & (layer3_outputs[1834]));
    assign layer4_outputs[1996] = ~((layer3_outputs[14]) | (layer3_outputs[1543]));
    assign layer4_outputs[1997] = layer3_outputs[1647];
    assign layer4_outputs[1998] = layer3_outputs[2747];
    assign layer4_outputs[1999] = (layer3_outputs[3617]) & ~(layer3_outputs[4951]);
    assign layer4_outputs[2000] = layer3_outputs[4762];
    assign layer4_outputs[2001] = ~(layer3_outputs[2367]);
    assign layer4_outputs[2002] = 1'b0;
    assign layer4_outputs[2003] = (layer3_outputs[1437]) & (layer3_outputs[4327]);
    assign layer4_outputs[2004] = layer3_outputs[2286];
    assign layer4_outputs[2005] = ~(layer3_outputs[701]);
    assign layer4_outputs[2006] = layer3_outputs[2078];
    assign layer4_outputs[2007] = (layer3_outputs[1453]) | (layer3_outputs[3435]);
    assign layer4_outputs[2008] = (layer3_outputs[3897]) & ~(layer3_outputs[4645]);
    assign layer4_outputs[2009] = layer3_outputs[2680];
    assign layer4_outputs[2010] = (layer3_outputs[4575]) & ~(layer3_outputs[2359]);
    assign layer4_outputs[2011] = ~(layer3_outputs[608]);
    assign layer4_outputs[2012] = (layer3_outputs[1005]) ^ (layer3_outputs[313]);
    assign layer4_outputs[2013] = ~((layer3_outputs[1840]) & (layer3_outputs[1425]));
    assign layer4_outputs[2014] = ~((layer3_outputs[619]) & (layer3_outputs[115]));
    assign layer4_outputs[2015] = ~(layer3_outputs[4893]);
    assign layer4_outputs[2016] = ~(layer3_outputs[4533]) | (layer3_outputs[4243]);
    assign layer4_outputs[2017] = ~(layer3_outputs[1159]) | (layer3_outputs[3943]);
    assign layer4_outputs[2018] = ~(layer3_outputs[3578]);
    assign layer4_outputs[2019] = ~(layer3_outputs[476]) | (layer3_outputs[1400]);
    assign layer4_outputs[2020] = (layer3_outputs[1656]) & ~(layer3_outputs[4916]);
    assign layer4_outputs[2021] = (layer3_outputs[4679]) | (layer3_outputs[5005]);
    assign layer4_outputs[2022] = ~(layer3_outputs[3292]) | (layer3_outputs[2844]);
    assign layer4_outputs[2023] = ~(layer3_outputs[4998]);
    assign layer4_outputs[2024] = (layer3_outputs[1284]) & ~(layer3_outputs[3982]);
    assign layer4_outputs[2025] = 1'b0;
    assign layer4_outputs[2026] = layer3_outputs[582];
    assign layer4_outputs[2027] = (layer3_outputs[4287]) & ~(layer3_outputs[3330]);
    assign layer4_outputs[2028] = ~((layer3_outputs[2153]) & (layer3_outputs[1940]));
    assign layer4_outputs[2029] = layer3_outputs[42];
    assign layer4_outputs[2030] = ~(layer3_outputs[1486]);
    assign layer4_outputs[2031] = (layer3_outputs[2903]) & ~(layer3_outputs[380]);
    assign layer4_outputs[2032] = ~((layer3_outputs[4989]) | (layer3_outputs[4384]));
    assign layer4_outputs[2033] = (layer3_outputs[3829]) | (layer3_outputs[2861]);
    assign layer4_outputs[2034] = ~(layer3_outputs[2307]);
    assign layer4_outputs[2035] = layer3_outputs[4191];
    assign layer4_outputs[2036] = ~((layer3_outputs[165]) & (layer3_outputs[1422]));
    assign layer4_outputs[2037] = ~(layer3_outputs[875]);
    assign layer4_outputs[2038] = ~(layer3_outputs[2587]);
    assign layer4_outputs[2039] = ~((layer3_outputs[987]) ^ (layer3_outputs[362]));
    assign layer4_outputs[2040] = ~((layer3_outputs[2843]) | (layer3_outputs[5019]));
    assign layer4_outputs[2041] = ~((layer3_outputs[475]) | (layer3_outputs[1138]));
    assign layer4_outputs[2042] = layer3_outputs[4778];
    assign layer4_outputs[2043] = ~(layer3_outputs[1395]) | (layer3_outputs[1971]);
    assign layer4_outputs[2044] = ~(layer3_outputs[4997]);
    assign layer4_outputs[2045] = ~((layer3_outputs[2754]) & (layer3_outputs[1637]));
    assign layer4_outputs[2046] = (layer3_outputs[3209]) | (layer3_outputs[4072]);
    assign layer4_outputs[2047] = ~(layer3_outputs[3496]) | (layer3_outputs[1649]);
    assign layer4_outputs[2048] = ~(layer3_outputs[1769]) | (layer3_outputs[4861]);
    assign layer4_outputs[2049] = layer3_outputs[4819];
    assign layer4_outputs[2050] = layer3_outputs[3982];
    assign layer4_outputs[2051] = ~(layer3_outputs[3002]) | (layer3_outputs[1878]);
    assign layer4_outputs[2052] = ~((layer3_outputs[2779]) & (layer3_outputs[4]));
    assign layer4_outputs[2053] = 1'b1;
    assign layer4_outputs[2054] = layer3_outputs[1959];
    assign layer4_outputs[2055] = ~(layer3_outputs[3018]);
    assign layer4_outputs[2056] = layer3_outputs[251];
    assign layer4_outputs[2057] = 1'b1;
    assign layer4_outputs[2058] = layer3_outputs[4094];
    assign layer4_outputs[2059] = ~(layer3_outputs[4941]) | (layer3_outputs[452]);
    assign layer4_outputs[2060] = ~((layer3_outputs[859]) | (layer3_outputs[2145]));
    assign layer4_outputs[2061] = ~(layer3_outputs[295]);
    assign layer4_outputs[2062] = ~(layer3_outputs[2445]);
    assign layer4_outputs[2063] = ~((layer3_outputs[4640]) ^ (layer3_outputs[4870]));
    assign layer4_outputs[2064] = ~(layer3_outputs[1670]) | (layer3_outputs[1455]);
    assign layer4_outputs[2065] = ~(layer3_outputs[2511]) | (layer3_outputs[5020]);
    assign layer4_outputs[2066] = (layer3_outputs[4052]) & ~(layer3_outputs[1101]);
    assign layer4_outputs[2067] = ~(layer3_outputs[2866]);
    assign layer4_outputs[2068] = layer3_outputs[3467];
    assign layer4_outputs[2069] = ~((layer3_outputs[3812]) & (layer3_outputs[3236]));
    assign layer4_outputs[2070] = layer3_outputs[255];
    assign layer4_outputs[2071] = layer3_outputs[1290];
    assign layer4_outputs[2072] = (layer3_outputs[3724]) & ~(layer3_outputs[1855]);
    assign layer4_outputs[2073] = 1'b0;
    assign layer4_outputs[2074] = layer3_outputs[3445];
    assign layer4_outputs[2075] = layer3_outputs[2694];
    assign layer4_outputs[2076] = ~(layer3_outputs[4028]) | (layer3_outputs[2146]);
    assign layer4_outputs[2077] = ~(layer3_outputs[1051]);
    assign layer4_outputs[2078] = (layer3_outputs[3254]) ^ (layer3_outputs[4140]);
    assign layer4_outputs[2079] = ~(layer3_outputs[3524]);
    assign layer4_outputs[2080] = (layer3_outputs[2578]) | (layer3_outputs[3285]);
    assign layer4_outputs[2081] = ~((layer3_outputs[2349]) ^ (layer3_outputs[584]));
    assign layer4_outputs[2082] = (layer3_outputs[1360]) & ~(layer3_outputs[3593]);
    assign layer4_outputs[2083] = ~((layer3_outputs[3375]) ^ (layer3_outputs[4088]));
    assign layer4_outputs[2084] = (layer3_outputs[2695]) | (layer3_outputs[4990]);
    assign layer4_outputs[2085] = layer3_outputs[1711];
    assign layer4_outputs[2086] = layer3_outputs[4425];
    assign layer4_outputs[2087] = ~(layer3_outputs[2666]);
    assign layer4_outputs[2088] = 1'b1;
    assign layer4_outputs[2089] = 1'b0;
    assign layer4_outputs[2090] = layer3_outputs[5054];
    assign layer4_outputs[2091] = layer3_outputs[2364];
    assign layer4_outputs[2092] = (layer3_outputs[2875]) & (layer3_outputs[4916]);
    assign layer4_outputs[2093] = layer3_outputs[1029];
    assign layer4_outputs[2094] = layer3_outputs[189];
    assign layer4_outputs[2095] = 1'b0;
    assign layer4_outputs[2096] = ~(layer3_outputs[653]);
    assign layer4_outputs[2097] = layer3_outputs[4632];
    assign layer4_outputs[2098] = (layer3_outputs[4821]) & ~(layer3_outputs[316]);
    assign layer4_outputs[2099] = (layer3_outputs[1607]) ^ (layer3_outputs[2853]);
    assign layer4_outputs[2100] = (layer3_outputs[1060]) & ~(layer3_outputs[2939]);
    assign layer4_outputs[2101] = ~(layer3_outputs[231]);
    assign layer4_outputs[2102] = (layer3_outputs[1803]) & ~(layer3_outputs[2978]);
    assign layer4_outputs[2103] = ~((layer3_outputs[2930]) & (layer3_outputs[3816]));
    assign layer4_outputs[2104] = ~(layer3_outputs[2576]) | (layer3_outputs[2063]);
    assign layer4_outputs[2105] = (layer3_outputs[1739]) ^ (layer3_outputs[2244]);
    assign layer4_outputs[2106] = ~(layer3_outputs[1775]);
    assign layer4_outputs[2107] = (layer3_outputs[1480]) & ~(layer3_outputs[11]);
    assign layer4_outputs[2108] = ~(layer3_outputs[3941]) | (layer3_outputs[1450]);
    assign layer4_outputs[2109] = ~(layer3_outputs[1547]);
    assign layer4_outputs[2110] = ~(layer3_outputs[354]);
    assign layer4_outputs[2111] = (layer3_outputs[1632]) ^ (layer3_outputs[447]);
    assign layer4_outputs[2112] = ~((layer3_outputs[591]) | (layer3_outputs[1506]));
    assign layer4_outputs[2113] = ~(layer3_outputs[4111]);
    assign layer4_outputs[2114] = ~((layer3_outputs[2155]) & (layer3_outputs[738]));
    assign layer4_outputs[2115] = (layer3_outputs[2080]) & (layer3_outputs[2013]);
    assign layer4_outputs[2116] = 1'b0;
    assign layer4_outputs[2117] = ~(layer3_outputs[2703]);
    assign layer4_outputs[2118] = ~(layer3_outputs[3938]) | (layer3_outputs[985]);
    assign layer4_outputs[2119] = (layer3_outputs[386]) & (layer3_outputs[4553]);
    assign layer4_outputs[2120] = layer3_outputs[3260];
    assign layer4_outputs[2121] = ~(layer3_outputs[3555]) | (layer3_outputs[2865]);
    assign layer4_outputs[2122] = (layer3_outputs[1108]) | (layer3_outputs[4157]);
    assign layer4_outputs[2123] = (layer3_outputs[4095]) & ~(layer3_outputs[3920]);
    assign layer4_outputs[2124] = layer3_outputs[2468];
    assign layer4_outputs[2125] = ~(layer3_outputs[2490]) | (layer3_outputs[1439]);
    assign layer4_outputs[2126] = layer3_outputs[2180];
    assign layer4_outputs[2127] = ~((layer3_outputs[1965]) ^ (layer3_outputs[1499]));
    assign layer4_outputs[2128] = (layer3_outputs[3861]) & (layer3_outputs[604]);
    assign layer4_outputs[2129] = ~(layer3_outputs[580]);
    assign layer4_outputs[2130] = 1'b0;
    assign layer4_outputs[2131] = ~(layer3_outputs[1980]);
    assign layer4_outputs[2132] = ~((layer3_outputs[296]) & (layer3_outputs[2475]));
    assign layer4_outputs[2133] = ~((layer3_outputs[1439]) | (layer3_outputs[2956]));
    assign layer4_outputs[2134] = layer3_outputs[2192];
    assign layer4_outputs[2135] = ~(layer3_outputs[138]);
    assign layer4_outputs[2136] = ~(layer3_outputs[1324]);
    assign layer4_outputs[2137] = ~((layer3_outputs[2591]) ^ (layer3_outputs[769]));
    assign layer4_outputs[2138] = layer3_outputs[1984];
    assign layer4_outputs[2139] = ~(layer3_outputs[2916]);
    assign layer4_outputs[2140] = ~(layer3_outputs[5046]) | (layer3_outputs[531]);
    assign layer4_outputs[2141] = layer3_outputs[1051];
    assign layer4_outputs[2142] = ~((layer3_outputs[2792]) & (layer3_outputs[435]));
    assign layer4_outputs[2143] = ~(layer3_outputs[3509]) | (layer3_outputs[38]);
    assign layer4_outputs[2144] = (layer3_outputs[4625]) & ~(layer3_outputs[4446]);
    assign layer4_outputs[2145] = (layer3_outputs[2565]) & (layer3_outputs[1954]);
    assign layer4_outputs[2146] = ~((layer3_outputs[554]) & (layer3_outputs[1521]));
    assign layer4_outputs[2147] = ~((layer3_outputs[4510]) | (layer3_outputs[1361]));
    assign layer4_outputs[2148] = (layer3_outputs[2455]) | (layer3_outputs[238]);
    assign layer4_outputs[2149] = layer3_outputs[1580];
    assign layer4_outputs[2150] = layer3_outputs[2797];
    assign layer4_outputs[2151] = ~((layer3_outputs[4161]) ^ (layer3_outputs[1623]));
    assign layer4_outputs[2152] = 1'b0;
    assign layer4_outputs[2153] = (layer3_outputs[2933]) & ~(layer3_outputs[1194]);
    assign layer4_outputs[2154] = 1'b1;
    assign layer4_outputs[2155] = layer3_outputs[1471];
    assign layer4_outputs[2156] = layer3_outputs[3970];
    assign layer4_outputs[2157] = ~((layer3_outputs[2634]) & (layer3_outputs[3803]));
    assign layer4_outputs[2158] = ~(layer3_outputs[2738]) | (layer3_outputs[3937]);
    assign layer4_outputs[2159] = layer3_outputs[2796];
    assign layer4_outputs[2160] = layer3_outputs[2076];
    assign layer4_outputs[2161] = layer3_outputs[895];
    assign layer4_outputs[2162] = (layer3_outputs[4804]) ^ (layer3_outputs[3568]);
    assign layer4_outputs[2163] = layer3_outputs[3272];
    assign layer4_outputs[2164] = (layer3_outputs[4119]) ^ (layer3_outputs[2891]);
    assign layer4_outputs[2165] = (layer3_outputs[2137]) & (layer3_outputs[2177]);
    assign layer4_outputs[2166] = ~(layer3_outputs[3881]) | (layer3_outputs[3329]);
    assign layer4_outputs[2167] = ~((layer3_outputs[3116]) & (layer3_outputs[494]));
    assign layer4_outputs[2168] = ~((layer3_outputs[1513]) & (layer3_outputs[3810]));
    assign layer4_outputs[2169] = (layer3_outputs[1708]) & (layer3_outputs[2197]);
    assign layer4_outputs[2170] = (layer3_outputs[1351]) & ~(layer3_outputs[3248]);
    assign layer4_outputs[2171] = ~(layer3_outputs[1821]);
    assign layer4_outputs[2172] = ~(layer3_outputs[4002]);
    assign layer4_outputs[2173] = layer3_outputs[1159];
    assign layer4_outputs[2174] = ~(layer3_outputs[480]);
    assign layer4_outputs[2175] = (layer3_outputs[55]) & ~(layer3_outputs[3047]);
    assign layer4_outputs[2176] = ~((layer3_outputs[557]) | (layer3_outputs[720]));
    assign layer4_outputs[2177] = layer3_outputs[4718];
    assign layer4_outputs[2178] = ~((layer3_outputs[1781]) | (layer3_outputs[3017]));
    assign layer4_outputs[2179] = layer3_outputs[4230];
    assign layer4_outputs[2180] = layer3_outputs[5023];
    assign layer4_outputs[2181] = ~(layer3_outputs[1349]);
    assign layer4_outputs[2182] = (layer3_outputs[2596]) & ~(layer3_outputs[2752]);
    assign layer4_outputs[2183] = 1'b0;
    assign layer4_outputs[2184] = (layer3_outputs[285]) & ~(layer3_outputs[4712]);
    assign layer4_outputs[2185] = (layer3_outputs[2681]) & ~(layer3_outputs[5026]);
    assign layer4_outputs[2186] = ~(layer3_outputs[1089]);
    assign layer4_outputs[2187] = ~((layer3_outputs[2444]) & (layer3_outputs[3778]));
    assign layer4_outputs[2188] = (layer3_outputs[805]) ^ (layer3_outputs[1212]);
    assign layer4_outputs[2189] = layer3_outputs[2790];
    assign layer4_outputs[2190] = ~((layer3_outputs[2570]) & (layer3_outputs[1498]));
    assign layer4_outputs[2191] = (layer3_outputs[3654]) & ~(layer3_outputs[2857]);
    assign layer4_outputs[2192] = layer3_outputs[610];
    assign layer4_outputs[2193] = ~(layer3_outputs[2468]) | (layer3_outputs[4701]);
    assign layer4_outputs[2194] = ~(layer3_outputs[3451]);
    assign layer4_outputs[2195] = ~(layer3_outputs[634]);
    assign layer4_outputs[2196] = ~(layer3_outputs[796]);
    assign layer4_outputs[2197] = (layer3_outputs[4330]) | (layer3_outputs[4329]);
    assign layer4_outputs[2198] = layer3_outputs[601];
    assign layer4_outputs[2199] = (layer3_outputs[2419]) & ~(layer3_outputs[4915]);
    assign layer4_outputs[2200] = ~(layer3_outputs[3877]);
    assign layer4_outputs[2201] = layer3_outputs[4247];
    assign layer4_outputs[2202] = ~(layer3_outputs[3631]) | (layer3_outputs[3402]);
    assign layer4_outputs[2203] = layer3_outputs[3698];
    assign layer4_outputs[2204] = ~(layer3_outputs[4876]) | (layer3_outputs[463]);
    assign layer4_outputs[2205] = ~(layer3_outputs[3611]) | (layer3_outputs[3]);
    assign layer4_outputs[2206] = layer3_outputs[1279];
    assign layer4_outputs[2207] = ~(layer3_outputs[3473]);
    assign layer4_outputs[2208] = (layer3_outputs[2442]) & (layer3_outputs[2422]);
    assign layer4_outputs[2209] = ~(layer3_outputs[4761]);
    assign layer4_outputs[2210] = ~((layer3_outputs[4586]) ^ (layer3_outputs[106]));
    assign layer4_outputs[2211] = layer3_outputs[5037];
    assign layer4_outputs[2212] = (layer3_outputs[70]) & (layer3_outputs[4093]);
    assign layer4_outputs[2213] = (layer3_outputs[4545]) & ~(layer3_outputs[2541]);
    assign layer4_outputs[2214] = (layer3_outputs[2510]) & ~(layer3_outputs[4806]);
    assign layer4_outputs[2215] = (layer3_outputs[4679]) | (layer3_outputs[1519]);
    assign layer4_outputs[2216] = ~(layer3_outputs[4336]) | (layer3_outputs[1591]);
    assign layer4_outputs[2217] = layer3_outputs[1553];
    assign layer4_outputs[2218] = ~((layer3_outputs[4053]) | (layer3_outputs[363]));
    assign layer4_outputs[2219] = ~((layer3_outputs[2361]) | (layer3_outputs[733]));
    assign layer4_outputs[2220] = layer3_outputs[1228];
    assign layer4_outputs[2221] = ~(layer3_outputs[4952]);
    assign layer4_outputs[2222] = ~(layer3_outputs[1048]);
    assign layer4_outputs[2223] = (layer3_outputs[4623]) & ~(layer3_outputs[2822]);
    assign layer4_outputs[2224] = 1'b1;
    assign layer4_outputs[2225] = ~((layer3_outputs[3762]) | (layer3_outputs[196]));
    assign layer4_outputs[2226] = ~((layer3_outputs[2300]) & (layer3_outputs[2962]));
    assign layer4_outputs[2227] = (layer3_outputs[1072]) & (layer3_outputs[3519]);
    assign layer4_outputs[2228] = (layer3_outputs[4801]) & ~(layer3_outputs[4628]);
    assign layer4_outputs[2229] = ~(layer3_outputs[821]);
    assign layer4_outputs[2230] = ~(layer3_outputs[4045]) | (layer3_outputs[2590]);
    assign layer4_outputs[2231] = layer3_outputs[1658];
    assign layer4_outputs[2232] = ~((layer3_outputs[173]) & (layer3_outputs[3947]));
    assign layer4_outputs[2233] = ~(layer3_outputs[220]);
    assign layer4_outputs[2234] = layer3_outputs[1203];
    assign layer4_outputs[2235] = 1'b0;
    assign layer4_outputs[2236] = 1'b1;
    assign layer4_outputs[2237] = (layer3_outputs[1239]) & (layer3_outputs[1520]);
    assign layer4_outputs[2238] = layer3_outputs[3138];
    assign layer4_outputs[2239] = layer3_outputs[801];
    assign layer4_outputs[2240] = ~(layer3_outputs[3085]) | (layer3_outputs[2537]);
    assign layer4_outputs[2241] = (layer3_outputs[1141]) & ~(layer3_outputs[4969]);
    assign layer4_outputs[2242] = (layer3_outputs[3101]) & ~(layer3_outputs[1440]);
    assign layer4_outputs[2243] = layer3_outputs[574];
    assign layer4_outputs[2244] = layer3_outputs[530];
    assign layer4_outputs[2245] = layer3_outputs[4726];
    assign layer4_outputs[2246] = (layer3_outputs[534]) ^ (layer3_outputs[1535]);
    assign layer4_outputs[2247] = ~((layer3_outputs[2727]) | (layer3_outputs[2882]));
    assign layer4_outputs[2248] = ~(layer3_outputs[2654]) | (layer3_outputs[3458]);
    assign layer4_outputs[2249] = (layer3_outputs[4774]) ^ (layer3_outputs[314]);
    assign layer4_outputs[2250] = layer3_outputs[188];
    assign layer4_outputs[2251] = (layer3_outputs[1059]) & (layer3_outputs[1710]);
    assign layer4_outputs[2252] = ~(layer3_outputs[4557]);
    assign layer4_outputs[2253] = layer3_outputs[915];
    assign layer4_outputs[2254] = layer3_outputs[1014];
    assign layer4_outputs[2255] = (layer3_outputs[4745]) ^ (layer3_outputs[1800]);
    assign layer4_outputs[2256] = ~((layer3_outputs[728]) & (layer3_outputs[1706]));
    assign layer4_outputs[2257] = 1'b0;
    assign layer4_outputs[2258] = ~((layer3_outputs[216]) | (layer3_outputs[113]));
    assign layer4_outputs[2259] = (layer3_outputs[3624]) & ~(layer3_outputs[5102]);
    assign layer4_outputs[2260] = layer3_outputs[4808];
    assign layer4_outputs[2261] = (layer3_outputs[3322]) & ~(layer3_outputs[3808]);
    assign layer4_outputs[2262] = layer3_outputs[3100];
    assign layer4_outputs[2263] = layer3_outputs[3599];
    assign layer4_outputs[2264] = ~(layer3_outputs[5107]) | (layer3_outputs[3480]);
    assign layer4_outputs[2265] = ~((layer3_outputs[824]) & (layer3_outputs[4570]));
    assign layer4_outputs[2266] = (layer3_outputs[3376]) & ~(layer3_outputs[2112]);
    assign layer4_outputs[2267] = layer3_outputs[2097];
    assign layer4_outputs[2268] = layer3_outputs[3268];
    assign layer4_outputs[2269] = layer3_outputs[3310];
    assign layer4_outputs[2270] = ~(layer3_outputs[2003]);
    assign layer4_outputs[2271] = 1'b1;
    assign layer4_outputs[2272] = layer3_outputs[957];
    assign layer4_outputs[2273] = ~(layer3_outputs[3900]);
    assign layer4_outputs[2274] = ~(layer3_outputs[4101]) | (layer3_outputs[2411]);
    assign layer4_outputs[2275] = 1'b1;
    assign layer4_outputs[2276] = (layer3_outputs[3715]) & (layer3_outputs[3664]);
    assign layer4_outputs[2277] = 1'b1;
    assign layer4_outputs[2278] = (layer3_outputs[2996]) & (layer3_outputs[3847]);
    assign layer4_outputs[2279] = 1'b1;
    assign layer4_outputs[2280] = ~(layer3_outputs[1407]);
    assign layer4_outputs[2281] = (layer3_outputs[137]) & ~(layer3_outputs[1759]);
    assign layer4_outputs[2282] = layer3_outputs[1463];
    assign layer4_outputs[2283] = ~(layer3_outputs[3287]);
    assign layer4_outputs[2284] = ~((layer3_outputs[2214]) & (layer3_outputs[2982]));
    assign layer4_outputs[2285] = (layer3_outputs[630]) & ~(layer3_outputs[838]);
    assign layer4_outputs[2286] = (layer3_outputs[2974]) & ~(layer3_outputs[208]);
    assign layer4_outputs[2287] = (layer3_outputs[3130]) & ~(layer3_outputs[1105]);
    assign layer4_outputs[2288] = 1'b1;
    assign layer4_outputs[2289] = ~(layer3_outputs[685]);
    assign layer4_outputs[2290] = 1'b1;
    assign layer4_outputs[2291] = ~((layer3_outputs[3268]) & (layer3_outputs[680]));
    assign layer4_outputs[2292] = ~((layer3_outputs[2030]) & (layer3_outputs[3367]));
    assign layer4_outputs[2293] = (layer3_outputs[3748]) & ~(layer3_outputs[1435]);
    assign layer4_outputs[2294] = ~(layer3_outputs[535]);
    assign layer4_outputs[2295] = ~(layer3_outputs[4095]);
    assign layer4_outputs[2296] = layer3_outputs[4541];
    assign layer4_outputs[2297] = (layer3_outputs[2545]) ^ (layer3_outputs[3807]);
    assign layer4_outputs[2298] = ~((layer3_outputs[2072]) | (layer3_outputs[1722]));
    assign layer4_outputs[2299] = 1'b1;
    assign layer4_outputs[2300] = 1'b1;
    assign layer4_outputs[2301] = layer3_outputs[1852];
    assign layer4_outputs[2302] = layer3_outputs[2018];
    assign layer4_outputs[2303] = (layer3_outputs[330]) & (layer3_outputs[775]);
    assign layer4_outputs[2304] = ~(layer3_outputs[3342]);
    assign layer4_outputs[2305] = 1'b0;
    assign layer4_outputs[2306] = ~(layer3_outputs[2540]);
    assign layer4_outputs[2307] = (layer3_outputs[541]) & (layer3_outputs[256]);
    assign layer4_outputs[2308] = (layer3_outputs[3732]) | (layer3_outputs[3067]);
    assign layer4_outputs[2309] = ~(layer3_outputs[1928]);
    assign layer4_outputs[2310] = 1'b1;
    assign layer4_outputs[2311] = ~(layer3_outputs[3806]) | (layer3_outputs[5073]);
    assign layer4_outputs[2312] = layer3_outputs[3904];
    assign layer4_outputs[2313] = layer3_outputs[581];
    assign layer4_outputs[2314] = ~((layer3_outputs[3169]) ^ (layer3_outputs[1889]));
    assign layer4_outputs[2315] = layer3_outputs[1091];
    assign layer4_outputs[2316] = layer3_outputs[3728];
    assign layer4_outputs[2317] = ~(layer3_outputs[3427]);
    assign layer4_outputs[2318] = layer3_outputs[4753];
    assign layer4_outputs[2319] = ~(layer3_outputs[4097]);
    assign layer4_outputs[2320] = layer3_outputs[486];
    assign layer4_outputs[2321] = ~(layer3_outputs[4785]);
    assign layer4_outputs[2322] = ~(layer3_outputs[999]);
    assign layer4_outputs[2323] = ~(layer3_outputs[4782]) | (layer3_outputs[3151]);
    assign layer4_outputs[2324] = ~(layer3_outputs[2102]) | (layer3_outputs[2862]);
    assign layer4_outputs[2325] = layer3_outputs[4430];
    assign layer4_outputs[2326] = 1'b0;
    assign layer4_outputs[2327] = (layer3_outputs[1326]) & ~(layer3_outputs[4425]);
    assign layer4_outputs[2328] = layer3_outputs[2793];
    assign layer4_outputs[2329] = ~(layer3_outputs[2113]);
    assign layer4_outputs[2330] = (layer3_outputs[4147]) & (layer3_outputs[1047]);
    assign layer4_outputs[2331] = ~(layer3_outputs[4148]);
    assign layer4_outputs[2332] = ~(layer3_outputs[2389]) | (layer3_outputs[3513]);
    assign layer4_outputs[2333] = ~((layer3_outputs[1514]) ^ (layer3_outputs[1742]));
    assign layer4_outputs[2334] = ~((layer3_outputs[5118]) & (layer3_outputs[1127]));
    assign layer4_outputs[2335] = layer3_outputs[4059];
    assign layer4_outputs[2336] = layer3_outputs[1664];
    assign layer4_outputs[2337] = (layer3_outputs[4476]) ^ (layer3_outputs[4892]);
    assign layer4_outputs[2338] = ~(layer3_outputs[4254]);
    assign layer4_outputs[2339] = layer3_outputs[2734];
    assign layer4_outputs[2340] = (layer3_outputs[4735]) & ~(layer3_outputs[1102]);
    assign layer4_outputs[2341] = ~((layer3_outputs[4937]) ^ (layer3_outputs[4766]));
    assign layer4_outputs[2342] = layer3_outputs[2533];
    assign layer4_outputs[2343] = (layer3_outputs[2781]) & (layer3_outputs[4706]);
    assign layer4_outputs[2344] = ~(layer3_outputs[4467]);
    assign layer4_outputs[2345] = ~(layer3_outputs[1098]);
    assign layer4_outputs[2346] = layer3_outputs[1736];
    assign layer4_outputs[2347] = ~((layer3_outputs[3384]) & (layer3_outputs[2067]));
    assign layer4_outputs[2348] = (layer3_outputs[3005]) ^ (layer3_outputs[705]);
    assign layer4_outputs[2349] = (layer3_outputs[4852]) & (layer3_outputs[41]);
    assign layer4_outputs[2350] = layer3_outputs[482];
    assign layer4_outputs[2351] = layer3_outputs[549];
    assign layer4_outputs[2352] = (layer3_outputs[2851]) & ~(layer3_outputs[3647]);
    assign layer4_outputs[2353] = (layer3_outputs[4784]) | (layer3_outputs[2225]);
    assign layer4_outputs[2354] = (layer3_outputs[3209]) & ~(layer3_outputs[4321]);
    assign layer4_outputs[2355] = ~(layer3_outputs[310]);
    assign layer4_outputs[2356] = layer3_outputs[5065];
    assign layer4_outputs[2357] = ~(layer3_outputs[1227]) | (layer3_outputs[2098]);
    assign layer4_outputs[2358] = ~(layer3_outputs[1758]);
    assign layer4_outputs[2359] = ~(layer3_outputs[842]);
    assign layer4_outputs[2360] = layer3_outputs[3616];
    assign layer4_outputs[2361] = 1'b1;
    assign layer4_outputs[2362] = ~(layer3_outputs[1004]) | (layer3_outputs[2646]);
    assign layer4_outputs[2363] = ~(layer3_outputs[4452]);
    assign layer4_outputs[2364] = ~(layer3_outputs[3509]);
    assign layer4_outputs[2365] = ~(layer3_outputs[3748]) | (layer3_outputs[210]);
    assign layer4_outputs[2366] = ~(layer3_outputs[2503]) | (layer3_outputs[2528]);
    assign layer4_outputs[2367] = (layer3_outputs[90]) | (layer3_outputs[930]);
    assign layer4_outputs[2368] = ~((layer3_outputs[2670]) | (layer3_outputs[981]));
    assign layer4_outputs[2369] = ~(layer3_outputs[3567]) | (layer3_outputs[4656]);
    assign layer4_outputs[2370] = ~((layer3_outputs[2944]) ^ (layer3_outputs[1885]));
    assign layer4_outputs[2371] = (layer3_outputs[1152]) & (layer3_outputs[886]);
    assign layer4_outputs[2372] = (layer3_outputs[2041]) & (layer3_outputs[4324]);
    assign layer4_outputs[2373] = ~((layer3_outputs[1931]) ^ (layer3_outputs[3323]));
    assign layer4_outputs[2374] = layer3_outputs[3628];
    assign layer4_outputs[2375] = ~(layer3_outputs[4239]) | (layer3_outputs[4831]);
    assign layer4_outputs[2376] = layer3_outputs[866];
    assign layer4_outputs[2377] = ~((layer3_outputs[3124]) & (layer3_outputs[1459]));
    assign layer4_outputs[2378] = 1'b0;
    assign layer4_outputs[2379] = layer3_outputs[2374];
    assign layer4_outputs[2380] = ~(layer3_outputs[3766]) | (layer3_outputs[1845]);
    assign layer4_outputs[2381] = layer3_outputs[1017];
    assign layer4_outputs[2382] = ~(layer3_outputs[107]);
    assign layer4_outputs[2383] = ~(layer3_outputs[356]);
    assign layer4_outputs[2384] = ~(layer3_outputs[207]);
    assign layer4_outputs[2385] = (layer3_outputs[4994]) & (layer3_outputs[958]);
    assign layer4_outputs[2386] = ~(layer3_outputs[2707]) | (layer3_outputs[3776]);
    assign layer4_outputs[2387] = ~(layer3_outputs[1171]);
    assign layer4_outputs[2388] = 1'b1;
    assign layer4_outputs[2389] = ~((layer3_outputs[1902]) ^ (layer3_outputs[1838]));
    assign layer4_outputs[2390] = (layer3_outputs[4125]) & ~(layer3_outputs[189]);
    assign layer4_outputs[2391] = ~(layer3_outputs[4767]);
    assign layer4_outputs[2392] = (layer3_outputs[833]) ^ (layer3_outputs[2717]);
    assign layer4_outputs[2393] = (layer3_outputs[303]) & ~(layer3_outputs[1288]);
    assign layer4_outputs[2394] = ~(layer3_outputs[506]) | (layer3_outputs[894]);
    assign layer4_outputs[2395] = ~((layer3_outputs[1965]) | (layer3_outputs[4356]));
    assign layer4_outputs[2396] = (layer3_outputs[3465]) & (layer3_outputs[83]);
    assign layer4_outputs[2397] = (layer3_outputs[3144]) | (layer3_outputs[335]);
    assign layer4_outputs[2398] = (layer3_outputs[529]) ^ (layer3_outputs[4628]);
    assign layer4_outputs[2399] = (layer3_outputs[1092]) & ~(layer3_outputs[4230]);
    assign layer4_outputs[2400] = layer3_outputs[458];
    assign layer4_outputs[2401] = 1'b1;
    assign layer4_outputs[2402] = (layer3_outputs[2006]) | (layer3_outputs[4600]);
    assign layer4_outputs[2403] = (layer3_outputs[4024]) ^ (layer3_outputs[3410]);
    assign layer4_outputs[2404] = ~((layer3_outputs[5082]) | (layer3_outputs[3820]));
    assign layer4_outputs[2405] = (layer3_outputs[4818]) & ~(layer3_outputs[352]);
    assign layer4_outputs[2406] = (layer3_outputs[1026]) & ~(layer3_outputs[4898]);
    assign layer4_outputs[2407] = ~((layer3_outputs[3401]) | (layer3_outputs[3810]));
    assign layer4_outputs[2408] = layer3_outputs[254];
    assign layer4_outputs[2409] = (layer3_outputs[1409]) ^ (layer3_outputs[3433]);
    assign layer4_outputs[2410] = ~(layer3_outputs[3257]);
    assign layer4_outputs[2411] = ~((layer3_outputs[1234]) | (layer3_outputs[4318]));
    assign layer4_outputs[2412] = ~(layer3_outputs[2558]) | (layer3_outputs[96]);
    assign layer4_outputs[2413] = ~(layer3_outputs[19]) | (layer3_outputs[843]);
    assign layer4_outputs[2414] = ~((layer3_outputs[5114]) & (layer3_outputs[2129]));
    assign layer4_outputs[2415] = 1'b0;
    assign layer4_outputs[2416] = (layer3_outputs[374]) | (layer3_outputs[3472]);
    assign layer4_outputs[2417] = layer3_outputs[1496];
    assign layer4_outputs[2418] = layer3_outputs[1700];
    assign layer4_outputs[2419] = ~(layer3_outputs[1766]) | (layer3_outputs[3685]);
    assign layer4_outputs[2420] = (layer3_outputs[30]) & (layer3_outputs[2965]);
    assign layer4_outputs[2421] = 1'b1;
    assign layer4_outputs[2422] = (layer3_outputs[698]) & (layer3_outputs[3991]);
    assign layer4_outputs[2423] = ~(layer3_outputs[1605]) | (layer3_outputs[876]);
    assign layer4_outputs[2424] = layer3_outputs[4657];
    assign layer4_outputs[2425] = (layer3_outputs[3724]) & (layer3_outputs[5006]);
    assign layer4_outputs[2426] = ~(layer3_outputs[3518]);
    assign layer4_outputs[2427] = (layer3_outputs[3906]) ^ (layer3_outputs[646]);
    assign layer4_outputs[2428] = (layer3_outputs[3185]) | (layer3_outputs[1323]);
    assign layer4_outputs[2429] = ~(layer3_outputs[2621]);
    assign layer4_outputs[2430] = ~(layer3_outputs[2556]);
    assign layer4_outputs[2431] = layer3_outputs[3712];
    assign layer4_outputs[2432] = layer3_outputs[4839];
    assign layer4_outputs[2433] = 1'b0;
    assign layer4_outputs[2434] = ~(layer3_outputs[4290]);
    assign layer4_outputs[2435] = layer3_outputs[2484];
    assign layer4_outputs[2436] = layer3_outputs[116];
    assign layer4_outputs[2437] = ~(layer3_outputs[4398]);
    assign layer4_outputs[2438] = 1'b0;
    assign layer4_outputs[2439] = ~(layer3_outputs[4683]);
    assign layer4_outputs[2440] = 1'b0;
    assign layer4_outputs[2441] = (layer3_outputs[4544]) | (layer3_outputs[4542]);
    assign layer4_outputs[2442] = (layer3_outputs[2143]) | (layer3_outputs[4370]);
    assign layer4_outputs[2443] = ~(layer3_outputs[4732]) | (layer3_outputs[975]);
    assign layer4_outputs[2444] = ~((layer3_outputs[478]) & (layer3_outputs[3633]));
    assign layer4_outputs[2445] = ~((layer3_outputs[3550]) | (layer3_outputs[4945]));
    assign layer4_outputs[2446] = 1'b0;
    assign layer4_outputs[2447] = ~(layer3_outputs[2520]);
    assign layer4_outputs[2448] = ~(layer3_outputs[3621]);
    assign layer4_outputs[2449] = (layer3_outputs[4383]) ^ (layer3_outputs[780]);
    assign layer4_outputs[2450] = ~(layer3_outputs[1325]);
    assign layer4_outputs[2451] = ~(layer3_outputs[3845]);
    assign layer4_outputs[2452] = ~(layer3_outputs[5040]);
    assign layer4_outputs[2453] = (layer3_outputs[4347]) & (layer3_outputs[1752]);
    assign layer4_outputs[2454] = layer3_outputs[4933];
    assign layer4_outputs[2455] = layer3_outputs[2250];
    assign layer4_outputs[2456] = layer3_outputs[1453];
    assign layer4_outputs[2457] = layer3_outputs[1486];
    assign layer4_outputs[2458] = ~(layer3_outputs[2467]);
    assign layer4_outputs[2459] = ~(layer3_outputs[3759]);
    assign layer4_outputs[2460] = ~((layer3_outputs[3439]) & (layer3_outputs[2421]));
    assign layer4_outputs[2461] = (layer3_outputs[344]) & ~(layer3_outputs[1789]);
    assign layer4_outputs[2462] = ~(layer3_outputs[174]) | (layer3_outputs[129]);
    assign layer4_outputs[2463] = layer3_outputs[446];
    assign layer4_outputs[2464] = (layer3_outputs[3563]) & (layer3_outputs[629]);
    assign layer4_outputs[2465] = ~((layer3_outputs[3862]) & (layer3_outputs[5104]));
    assign layer4_outputs[2466] = layer3_outputs[4076];
    assign layer4_outputs[2467] = ~(layer3_outputs[814]);
    assign layer4_outputs[2468] = layer3_outputs[2205];
    assign layer4_outputs[2469] = ~((layer3_outputs[1259]) | (layer3_outputs[1321]));
    assign layer4_outputs[2470] = (layer3_outputs[4013]) & ~(layer3_outputs[3184]);
    assign layer4_outputs[2471] = ~(layer3_outputs[100]) | (layer3_outputs[1781]);
    assign layer4_outputs[2472] = layer3_outputs[1183];
    assign layer4_outputs[2473] = (layer3_outputs[1054]) & (layer3_outputs[2132]);
    assign layer4_outputs[2474] = ~(layer3_outputs[77]) | (layer3_outputs[795]);
    assign layer4_outputs[2475] = (layer3_outputs[1863]) | (layer3_outputs[3131]);
    assign layer4_outputs[2476] = layer3_outputs[4172];
    assign layer4_outputs[2477] = ~(layer3_outputs[1227]) | (layer3_outputs[1223]);
    assign layer4_outputs[2478] = (layer3_outputs[3237]) & ~(layer3_outputs[2214]);
    assign layer4_outputs[2479] = ~(layer3_outputs[2240]);
    assign layer4_outputs[2480] = (layer3_outputs[4539]) & ~(layer3_outputs[1574]);
    assign layer4_outputs[2481] = ~(layer3_outputs[4724]);
    assign layer4_outputs[2482] = layer3_outputs[92];
    assign layer4_outputs[2483] = ~(layer3_outputs[1369]);
    assign layer4_outputs[2484] = ~(layer3_outputs[2062]);
    assign layer4_outputs[2485] = ~((layer3_outputs[2796]) | (layer3_outputs[3076]));
    assign layer4_outputs[2486] = (layer3_outputs[1470]) & ~(layer3_outputs[4640]);
    assign layer4_outputs[2487] = (layer3_outputs[3093]) ^ (layer3_outputs[2338]);
    assign layer4_outputs[2488] = ~((layer3_outputs[2879]) ^ (layer3_outputs[1095]));
    assign layer4_outputs[2489] = 1'b0;
    assign layer4_outputs[2490] = ~((layer3_outputs[1483]) ^ (layer3_outputs[1008]));
    assign layer4_outputs[2491] = ~(layer3_outputs[499]);
    assign layer4_outputs[2492] = ~(layer3_outputs[1890]);
    assign layer4_outputs[2493] = ~(layer3_outputs[4677]);
    assign layer4_outputs[2494] = ~(layer3_outputs[3710]);
    assign layer4_outputs[2495] = ~((layer3_outputs[3577]) & (layer3_outputs[533]));
    assign layer4_outputs[2496] = layer3_outputs[2105];
    assign layer4_outputs[2497] = (layer3_outputs[2631]) ^ (layer3_outputs[4211]);
    assign layer4_outputs[2498] = ~(layer3_outputs[4428]);
    assign layer4_outputs[2499] = (layer3_outputs[3983]) & ~(layer3_outputs[4460]);
    assign layer4_outputs[2500] = ~((layer3_outputs[3289]) & (layer3_outputs[282]));
    assign layer4_outputs[2501] = layer3_outputs[4970];
    assign layer4_outputs[2502] = layer3_outputs[2418];
    assign layer4_outputs[2503] = ~(layer3_outputs[3775]);
    assign layer4_outputs[2504] = 1'b1;
    assign layer4_outputs[2505] = ~((layer3_outputs[3935]) & (layer3_outputs[497]));
    assign layer4_outputs[2506] = (layer3_outputs[4071]) & (layer3_outputs[3795]);
    assign layer4_outputs[2507] = layer3_outputs[2470];
    assign layer4_outputs[2508] = ~((layer3_outputs[4692]) ^ (layer3_outputs[168]));
    assign layer4_outputs[2509] = layer3_outputs[1660];
    assign layer4_outputs[2510] = ~(layer3_outputs[2393]) | (layer3_outputs[3274]);
    assign layer4_outputs[2511] = ~(layer3_outputs[4211]);
    assign layer4_outputs[2512] = (layer3_outputs[4468]) ^ (layer3_outputs[4759]);
    assign layer4_outputs[2513] = ~(layer3_outputs[2919]);
    assign layer4_outputs[2514] = ~(layer3_outputs[2560]);
    assign layer4_outputs[2515] = (layer3_outputs[675]) & ~(layer3_outputs[2498]);
    assign layer4_outputs[2516] = ~(layer3_outputs[723]) | (layer3_outputs[887]);
    assign layer4_outputs[2517] = (layer3_outputs[306]) | (layer3_outputs[4917]);
    assign layer4_outputs[2518] = ~(layer3_outputs[3933]) | (layer3_outputs[606]);
    assign layer4_outputs[2519] = 1'b0;
    assign layer4_outputs[2520] = 1'b1;
    assign layer4_outputs[2521] = layer3_outputs[3068];
    assign layer4_outputs[2522] = 1'b1;
    assign layer4_outputs[2523] = ~(layer3_outputs[3366]);
    assign layer4_outputs[2524] = layer3_outputs[27];
    assign layer4_outputs[2525] = ~(layer3_outputs[2773]) | (layer3_outputs[2472]);
    assign layer4_outputs[2526] = 1'b1;
    assign layer4_outputs[2527] = (layer3_outputs[3545]) ^ (layer3_outputs[350]);
    assign layer4_outputs[2528] = layer3_outputs[1053];
    assign layer4_outputs[2529] = layer3_outputs[978];
    assign layer4_outputs[2530] = (layer3_outputs[3108]) ^ (layer3_outputs[1402]);
    assign layer4_outputs[2531] = ~((layer3_outputs[3677]) ^ (layer3_outputs[3738]));
    assign layer4_outputs[2532] = ~(layer3_outputs[4851]) | (layer3_outputs[4402]);
    assign layer4_outputs[2533] = ~((layer3_outputs[2924]) & (layer3_outputs[4877]));
    assign layer4_outputs[2534] = layer3_outputs[3072];
    assign layer4_outputs[2535] = ~(layer3_outputs[1610]);
    assign layer4_outputs[2536] = ~(layer3_outputs[1475]) | (layer3_outputs[4570]);
    assign layer4_outputs[2537] = ~(layer3_outputs[4368]);
    assign layer4_outputs[2538] = layer3_outputs[3270];
    assign layer4_outputs[2539] = ~((layer3_outputs[2053]) & (layer3_outputs[1382]));
    assign layer4_outputs[2540] = ~(layer3_outputs[1283]);
    assign layer4_outputs[2541] = layer3_outputs[956];
    assign layer4_outputs[2542] = 1'b1;
    assign layer4_outputs[2543] = ~(layer3_outputs[3600]);
    assign layer4_outputs[2544] = ~(layer3_outputs[2682]);
    assign layer4_outputs[2545] = ~((layer3_outputs[2632]) | (layer3_outputs[3446]));
    assign layer4_outputs[2546] = ~(layer3_outputs[2559]) | (layer3_outputs[1532]);
    assign layer4_outputs[2547] = layer3_outputs[721];
    assign layer4_outputs[2548] = layer3_outputs[1009];
    assign layer4_outputs[2549] = layer3_outputs[4576];
    assign layer4_outputs[2550] = (layer3_outputs[4795]) & ~(layer3_outputs[5072]);
    assign layer4_outputs[2551] = (layer3_outputs[3329]) & ~(layer3_outputs[2633]);
    assign layer4_outputs[2552] = ~((layer3_outputs[4531]) | (layer3_outputs[4978]));
    assign layer4_outputs[2553] = layer3_outputs[1910];
    assign layer4_outputs[2554] = ~(layer3_outputs[3556]);
    assign layer4_outputs[2555] = (layer3_outputs[4550]) & ~(layer3_outputs[2828]);
    assign layer4_outputs[2556] = layer3_outputs[1847];
    assign layer4_outputs[2557] = layer3_outputs[3869];
    assign layer4_outputs[2558] = 1'b0;
    assign layer4_outputs[2559] = ~(layer3_outputs[3846]) | (layer3_outputs[4944]);
    assign layer4_outputs[2560] = 1'b1;
    assign layer4_outputs[2561] = (layer3_outputs[1457]) & ~(layer3_outputs[2020]);
    assign layer4_outputs[2562] = (layer3_outputs[624]) & ~(layer3_outputs[2776]);
    assign layer4_outputs[2563] = layer3_outputs[3473];
    assign layer4_outputs[2564] = layer3_outputs[816];
    assign layer4_outputs[2565] = (layer3_outputs[590]) & ~(layer3_outputs[1357]);
    assign layer4_outputs[2566] = ~(layer3_outputs[2341]) | (layer3_outputs[576]);
    assign layer4_outputs[2567] = (layer3_outputs[2850]) & ~(layer3_outputs[1433]);
    assign layer4_outputs[2568] = layer3_outputs[2012];
    assign layer4_outputs[2569] = ~((layer3_outputs[3795]) ^ (layer3_outputs[940]));
    assign layer4_outputs[2570] = ~(layer3_outputs[1611]);
    assign layer4_outputs[2571] = layer3_outputs[5030];
    assign layer4_outputs[2572] = ~(layer3_outputs[3012]) | (layer3_outputs[3957]);
    assign layer4_outputs[2573] = ~(layer3_outputs[2894]);
    assign layer4_outputs[2574] = ~(layer3_outputs[4121]);
    assign layer4_outputs[2575] = (layer3_outputs[2364]) & ~(layer3_outputs[2230]);
    assign layer4_outputs[2576] = layer3_outputs[2239];
    assign layer4_outputs[2577] = ~(layer3_outputs[141]);
    assign layer4_outputs[2578] = layer3_outputs[983];
    assign layer4_outputs[2579] = ~(layer3_outputs[1581]);
    assign layer4_outputs[2580] = (layer3_outputs[743]) & ~(layer3_outputs[4643]);
    assign layer4_outputs[2581] = ~((layer3_outputs[2751]) ^ (layer3_outputs[1696]));
    assign layer4_outputs[2582] = (layer3_outputs[1890]) | (layer3_outputs[2769]);
    assign layer4_outputs[2583] = (layer3_outputs[510]) & (layer3_outputs[4007]);
    assign layer4_outputs[2584] = (layer3_outputs[1976]) ^ (layer3_outputs[989]);
    assign layer4_outputs[2585] = ~(layer3_outputs[3975]) | (layer3_outputs[1119]);
    assign layer4_outputs[2586] = ~(layer3_outputs[2028]);
    assign layer4_outputs[2587] = ~(layer3_outputs[1743]) | (layer3_outputs[2660]);
    assign layer4_outputs[2588] = layer3_outputs[2193];
    assign layer4_outputs[2589] = 1'b1;
    assign layer4_outputs[2590] = ~(layer3_outputs[2331]);
    assign layer4_outputs[2591] = ~((layer3_outputs[24]) ^ (layer3_outputs[4176]));
    assign layer4_outputs[2592] = (layer3_outputs[4526]) ^ (layer3_outputs[4824]);
    assign layer4_outputs[2593] = ~((layer3_outputs[107]) ^ (layer3_outputs[2437]));
    assign layer4_outputs[2594] = (layer3_outputs[2267]) | (layer3_outputs[2178]);
    assign layer4_outputs[2595] = ~((layer3_outputs[831]) | (layer3_outputs[1213]));
    assign layer4_outputs[2596] = layer3_outputs[313];
    assign layer4_outputs[2597] = layer3_outputs[4748];
    assign layer4_outputs[2598] = layer3_outputs[2341];
    assign layer4_outputs[2599] = (layer3_outputs[545]) | (layer3_outputs[2339]);
    assign layer4_outputs[2600] = ~(layer3_outputs[3220]);
    assign layer4_outputs[2601] = ~(layer3_outputs[464]) | (layer3_outputs[3421]);
    assign layer4_outputs[2602] = ~(layer3_outputs[1148]);
    assign layer4_outputs[2603] = (layer3_outputs[2593]) | (layer3_outputs[4059]);
    assign layer4_outputs[2604] = 1'b1;
    assign layer4_outputs[2605] = ~(layer3_outputs[456]);
    assign layer4_outputs[2606] = ~(layer3_outputs[1103]);
    assign layer4_outputs[2607] = layer3_outputs[230];
    assign layer4_outputs[2608] = (layer3_outputs[4219]) & ~(layer3_outputs[3796]);
    assign layer4_outputs[2609] = (layer3_outputs[438]) & (layer3_outputs[3142]);
    assign layer4_outputs[2610] = layer3_outputs[1465];
    assign layer4_outputs[2611] = ~((layer3_outputs[1872]) | (layer3_outputs[3031]));
    assign layer4_outputs[2612] = ~(layer3_outputs[2926]);
    assign layer4_outputs[2613] = (layer3_outputs[4948]) & (layer3_outputs[3925]);
    assign layer4_outputs[2614] = ~(layer3_outputs[882]);
    assign layer4_outputs[2615] = (layer3_outputs[890]) & ~(layer3_outputs[3635]);
    assign layer4_outputs[2616] = ~(layer3_outputs[84]);
    assign layer4_outputs[2617] = ~(layer3_outputs[1794]);
    assign layer4_outputs[2618] = ~(layer3_outputs[3482]);
    assign layer4_outputs[2619] = (layer3_outputs[152]) & ~(layer3_outputs[4023]);
    assign layer4_outputs[2620] = ~((layer3_outputs[905]) & (layer3_outputs[1954]));
    assign layer4_outputs[2621] = (layer3_outputs[221]) | (layer3_outputs[3734]);
    assign layer4_outputs[2622] = ~(layer3_outputs[2134]) | (layer3_outputs[1142]);
    assign layer4_outputs[2623] = (layer3_outputs[4138]) | (layer3_outputs[1445]);
    assign layer4_outputs[2624] = ~((layer3_outputs[350]) & (layer3_outputs[4073]));
    assign layer4_outputs[2625] = (layer3_outputs[5081]) & ~(layer3_outputs[1124]);
    assign layer4_outputs[2626] = ~((layer3_outputs[1944]) | (layer3_outputs[1165]));
    assign layer4_outputs[2627] = 1'b0;
    assign layer4_outputs[2628] = layer3_outputs[1951];
    assign layer4_outputs[2629] = ~(layer3_outputs[3429]) | (layer3_outputs[4171]);
    assign layer4_outputs[2630] = ~(layer3_outputs[1970]);
    assign layer4_outputs[2631] = layer3_outputs[4698];
    assign layer4_outputs[2632] = 1'b0;
    assign layer4_outputs[2633] = (layer3_outputs[3360]) ^ (layer3_outputs[4719]);
    assign layer4_outputs[2634] = ~(layer3_outputs[3466]);
    assign layer4_outputs[2635] = layer3_outputs[553];
    assign layer4_outputs[2636] = ~((layer3_outputs[1181]) & (layer3_outputs[3864]));
    assign layer4_outputs[2637] = layer3_outputs[4522];
    assign layer4_outputs[2638] = 1'b1;
    assign layer4_outputs[2639] = layer3_outputs[1546];
    assign layer4_outputs[2640] = layer3_outputs[635];
    assign layer4_outputs[2641] = ~(layer3_outputs[3053]);
    assign layer4_outputs[2642] = (layer3_outputs[1046]) & ~(layer3_outputs[4195]);
    assign layer4_outputs[2643] = layer3_outputs[2291];
    assign layer4_outputs[2644] = ~(layer3_outputs[4993]);
    assign layer4_outputs[2645] = ~(layer3_outputs[3311]) | (layer3_outputs[75]);
    assign layer4_outputs[2646] = (layer3_outputs[3099]) & ~(layer3_outputs[480]);
    assign layer4_outputs[2647] = (layer3_outputs[2973]) & ~(layer3_outputs[3875]);
    assign layer4_outputs[2648] = 1'b0;
    assign layer4_outputs[2649] = ~(layer3_outputs[422]);
    assign layer4_outputs[2650] = ~((layer3_outputs[991]) | (layer3_outputs[272]));
    assign layer4_outputs[2651] = (layer3_outputs[2805]) | (layer3_outputs[236]);
    assign layer4_outputs[2652] = (layer3_outputs[1429]) & ~(layer3_outputs[4623]);
    assign layer4_outputs[2653] = layer3_outputs[3946];
    assign layer4_outputs[2654] = ~(layer3_outputs[3475]);
    assign layer4_outputs[2655] = (layer3_outputs[1938]) & ~(layer3_outputs[2761]);
    assign layer4_outputs[2656] = layer3_outputs[1094];
    assign layer4_outputs[2657] = (layer3_outputs[5091]) | (layer3_outputs[2709]);
    assign layer4_outputs[2658] = (layer3_outputs[1114]) & (layer3_outputs[4308]);
    assign layer4_outputs[2659] = ~((layer3_outputs[3377]) & (layer3_outputs[1174]));
    assign layer4_outputs[2660] = ~(layer3_outputs[3305]) | (layer3_outputs[692]);
    assign layer4_outputs[2661] = ~((layer3_outputs[3669]) & (layer3_outputs[3926]));
    assign layer4_outputs[2662] = ~(layer3_outputs[2564]) | (layer3_outputs[2846]);
    assign layer4_outputs[2663] = (layer3_outputs[2524]) | (layer3_outputs[1955]);
    assign layer4_outputs[2664] = (layer3_outputs[4660]) | (layer3_outputs[3199]);
    assign layer4_outputs[2665] = layer3_outputs[1176];
    assign layer4_outputs[2666] = (layer3_outputs[539]) | (layer3_outputs[441]);
    assign layer4_outputs[2667] = layer3_outputs[2918];
    assign layer4_outputs[2668] = 1'b1;
    assign layer4_outputs[2669] = ~(layer3_outputs[3957]);
    assign layer4_outputs[2670] = layer3_outputs[1960];
    assign layer4_outputs[2671] = ~((layer3_outputs[4704]) | (layer3_outputs[242]));
    assign layer4_outputs[2672] = ~(layer3_outputs[2282]) | (layer3_outputs[4965]);
    assign layer4_outputs[2673] = layer3_outputs[5029];
    assign layer4_outputs[2674] = (layer3_outputs[2068]) | (layer3_outputs[1559]);
    assign layer4_outputs[2675] = ~(layer3_outputs[1683]);
    assign layer4_outputs[2676] = ~((layer3_outputs[3283]) ^ (layer3_outputs[3623]));
    assign layer4_outputs[2677] = layer3_outputs[1962];
    assign layer4_outputs[2678] = layer3_outputs[974];
    assign layer4_outputs[2679] = layer3_outputs[2379];
    assign layer4_outputs[2680] = layer3_outputs[2338];
    assign layer4_outputs[2681] = ~(layer3_outputs[3119]) | (layer3_outputs[788]);
    assign layer4_outputs[2682] = ~(layer3_outputs[3863]);
    assign layer4_outputs[2683] = ~((layer3_outputs[2709]) & (layer3_outputs[3667]));
    assign layer4_outputs[2684] = ~(layer3_outputs[468]) | (layer3_outputs[3693]);
    assign layer4_outputs[2685] = ~(layer3_outputs[2409]);
    assign layer4_outputs[2686] = ~(layer3_outputs[2652]);
    assign layer4_outputs[2687] = (layer3_outputs[703]) ^ (layer3_outputs[1258]);
    assign layer4_outputs[2688] = layer3_outputs[1322];
    assign layer4_outputs[2689] = ~((layer3_outputs[3278]) ^ (layer3_outputs[1649]));
    assign layer4_outputs[2690] = ~(layer3_outputs[3925]);
    assign layer4_outputs[2691] = (layer3_outputs[1680]) | (layer3_outputs[2556]);
    assign layer4_outputs[2692] = ~(layer3_outputs[2544]);
    assign layer4_outputs[2693] = ~(layer3_outputs[3643]) | (layer3_outputs[2837]);
    assign layer4_outputs[2694] = (layer3_outputs[3453]) & (layer3_outputs[1810]);
    assign layer4_outputs[2695] = layer3_outputs[3224];
    assign layer4_outputs[2696] = ~(layer3_outputs[4963]);
    assign layer4_outputs[2697] = ~(layer3_outputs[4156]) | (layer3_outputs[3630]);
    assign layer4_outputs[2698] = (layer3_outputs[62]) | (layer3_outputs[4728]);
    assign layer4_outputs[2699] = ~(layer3_outputs[2477]);
    assign layer4_outputs[2700] = ~((layer3_outputs[4598]) ^ (layer3_outputs[1481]));
    assign layer4_outputs[2701] = ~(layer3_outputs[225]);
    assign layer4_outputs[2702] = (layer3_outputs[3405]) & ~(layer3_outputs[2554]);
    assign layer4_outputs[2703] = ~((layer3_outputs[436]) | (layer3_outputs[2906]));
    assign layer4_outputs[2704] = ~(layer3_outputs[3080]) | (layer3_outputs[2737]);
    assign layer4_outputs[2705] = (layer3_outputs[2005]) & ~(layer3_outputs[1000]);
    assign layer4_outputs[2706] = ~(layer3_outputs[238]);
    assign layer4_outputs[2707] = ~((layer3_outputs[2147]) & (layer3_outputs[359]));
    assign layer4_outputs[2708] = layer3_outputs[1908];
    assign layer4_outputs[2709] = layer3_outputs[816];
    assign layer4_outputs[2710] = (layer3_outputs[202]) & ~(layer3_outputs[3003]);
    assign layer4_outputs[2711] = ~((layer3_outputs[183]) | (layer3_outputs[5038]));
    assign layer4_outputs[2712] = ~((layer3_outputs[2221]) | (layer3_outputs[4479]));
    assign layer4_outputs[2713] = ~((layer3_outputs[3746]) | (layer3_outputs[1248]));
    assign layer4_outputs[2714] = ~((layer3_outputs[3234]) | (layer3_outputs[3385]));
    assign layer4_outputs[2715] = ~(layer3_outputs[2994]) | (layer3_outputs[3377]);
    assign layer4_outputs[2716] = layer3_outputs[3769];
    assign layer4_outputs[2717] = (layer3_outputs[926]) ^ (layer3_outputs[3256]);
    assign layer4_outputs[2718] = (layer3_outputs[3962]) & ~(layer3_outputs[4364]);
    assign layer4_outputs[2719] = ~(layer3_outputs[244]) | (layer3_outputs[5022]);
    assign layer4_outputs[2720] = ~(layer3_outputs[4534]);
    assign layer4_outputs[2721] = (layer3_outputs[4895]) & (layer3_outputs[3495]);
    assign layer4_outputs[2722] = ~(layer3_outputs[202]);
    assign layer4_outputs[2723] = 1'b1;
    assign layer4_outputs[2724] = ~(layer3_outputs[2028]);
    assign layer4_outputs[2725] = (layer3_outputs[3514]) ^ (layer3_outputs[1638]);
    assign layer4_outputs[2726] = ~(layer3_outputs[466]);
    assign layer4_outputs[2727] = 1'b1;
    assign layer4_outputs[2728] = (layer3_outputs[3988]) ^ (layer3_outputs[2669]);
    assign layer4_outputs[2729] = layer3_outputs[1823];
    assign layer4_outputs[2730] = 1'b1;
    assign layer4_outputs[2731] = ~(layer3_outputs[718]);
    assign layer4_outputs[2732] = ~(layer3_outputs[1388]);
    assign layer4_outputs[2733] = (layer3_outputs[71]) & ~(layer3_outputs[4541]);
    assign layer4_outputs[2734] = ~(layer3_outputs[5090]) | (layer3_outputs[664]);
    assign layer4_outputs[2735] = layer3_outputs[1046];
    assign layer4_outputs[2736] = (layer3_outputs[1989]) & (layer3_outputs[4264]);
    assign layer4_outputs[2737] = layer3_outputs[3105];
    assign layer4_outputs[2738] = ~((layer3_outputs[2055]) & (layer3_outputs[1603]));
    assign layer4_outputs[2739] = ~(layer3_outputs[2995]);
    assign layer4_outputs[2740] = layer3_outputs[2561];
    assign layer4_outputs[2741] = ~((layer3_outputs[2147]) | (layer3_outputs[4843]));
    assign layer4_outputs[2742] = ~((layer3_outputs[2515]) & (layer3_outputs[3399]));
    assign layer4_outputs[2743] = layer3_outputs[4912];
    assign layer4_outputs[2744] = ~(layer3_outputs[2310]);
    assign layer4_outputs[2745] = ~(layer3_outputs[795]);
    assign layer4_outputs[2746] = layer3_outputs[4292];
    assign layer4_outputs[2747] = layer3_outputs[3211];
    assign layer4_outputs[2748] = (layer3_outputs[3777]) | (layer3_outputs[4178]);
    assign layer4_outputs[2749] = layer3_outputs[2017];
    assign layer4_outputs[2750] = layer3_outputs[3851];
    assign layer4_outputs[2751] = ~(layer3_outputs[2612]) | (layer3_outputs[3610]);
    assign layer4_outputs[2752] = (layer3_outputs[1796]) & (layer3_outputs[3874]);
    assign layer4_outputs[2753] = ~(layer3_outputs[397]) | (layer3_outputs[2542]);
    assign layer4_outputs[2754] = layer3_outputs[1700];
    assign layer4_outputs[2755] = 1'b0;
    assign layer4_outputs[2756] = 1'b0;
    assign layer4_outputs[2757] = layer3_outputs[1705];
    assign layer4_outputs[2758] = 1'b0;
    assign layer4_outputs[2759] = (layer3_outputs[3965]) | (layer3_outputs[1079]);
    assign layer4_outputs[2760] = ~(layer3_outputs[3841]);
    assign layer4_outputs[2761] = ~(layer3_outputs[2856]);
    assign layer4_outputs[2762] = (layer3_outputs[1741]) & (layer3_outputs[4789]);
    assign layer4_outputs[2763] = layer3_outputs[5027];
    assign layer4_outputs[2764] = (layer3_outputs[4622]) & (layer3_outputs[3825]);
    assign layer4_outputs[2765] = (layer3_outputs[3557]) | (layer3_outputs[3015]);
    assign layer4_outputs[2766] = ~(layer3_outputs[3635]);
    assign layer4_outputs[2767] = (layer3_outputs[708]) ^ (layer3_outputs[250]);
    assign layer4_outputs[2768] = (layer3_outputs[4741]) | (layer3_outputs[777]);
    assign layer4_outputs[2769] = (layer3_outputs[4244]) & ~(layer3_outputs[2928]);
    assign layer4_outputs[2770] = ~(layer3_outputs[4199]);
    assign layer4_outputs[2771] = layer3_outputs[205];
    assign layer4_outputs[2772] = (layer3_outputs[4958]) | (layer3_outputs[481]);
    assign layer4_outputs[2773] = ~(layer3_outputs[4771]) | (layer3_outputs[4881]);
    assign layer4_outputs[2774] = 1'b0;
    assign layer4_outputs[2775] = ~(layer3_outputs[3043]);
    assign layer4_outputs[2776] = (layer3_outputs[401]) & ~(layer3_outputs[1941]);
    assign layer4_outputs[2777] = ~(layer3_outputs[2653]);
    assign layer4_outputs[2778] = ~((layer3_outputs[4751]) & (layer3_outputs[2061]));
    assign layer4_outputs[2779] = (layer3_outputs[2917]) & ~(layer3_outputs[2288]);
    assign layer4_outputs[2780] = ~(layer3_outputs[597]);
    assign layer4_outputs[2781] = layer3_outputs[2168];
    assign layer4_outputs[2782] = ~(layer3_outputs[3954]);
    assign layer4_outputs[2783] = 1'b0;
    assign layer4_outputs[2784] = 1'b1;
    assign layer4_outputs[2785] = layer3_outputs[4774];
    assign layer4_outputs[2786] = 1'b1;
    assign layer4_outputs[2787] = ~(layer3_outputs[4867]);
    assign layer4_outputs[2788] = (layer3_outputs[2083]) & (layer3_outputs[3000]);
    assign layer4_outputs[2789] = ~(layer3_outputs[834]) | (layer3_outputs[155]);
    assign layer4_outputs[2790] = 1'b1;
    assign layer4_outputs[2791] = (layer3_outputs[560]) ^ (layer3_outputs[2775]);
    assign layer4_outputs[2792] = (layer3_outputs[417]) | (layer3_outputs[2980]);
    assign layer4_outputs[2793] = ~(layer3_outputs[1344]);
    assign layer4_outputs[2794] = layer3_outputs[5003];
    assign layer4_outputs[2795] = (layer3_outputs[2646]) & ~(layer3_outputs[3059]);
    assign layer4_outputs[2796] = layer3_outputs[4647];
    assign layer4_outputs[2797] = layer3_outputs[4353];
    assign layer4_outputs[2798] = layer3_outputs[3028];
    assign layer4_outputs[2799] = layer3_outputs[4759];
    assign layer4_outputs[2800] = ~(layer3_outputs[3726]);
    assign layer4_outputs[2801] = (layer3_outputs[4404]) | (layer3_outputs[3133]);
    assign layer4_outputs[2802] = 1'b1;
    assign layer4_outputs[2803] = ~(layer3_outputs[909]);
    assign layer4_outputs[2804] = (layer3_outputs[4452]) | (layer3_outputs[2400]);
    assign layer4_outputs[2805] = ~(layer3_outputs[1555]);
    assign layer4_outputs[2806] = layer3_outputs[213];
    assign layer4_outputs[2807] = layer3_outputs[5080];
    assign layer4_outputs[2808] = (layer3_outputs[2525]) & (layer3_outputs[4763]);
    assign layer4_outputs[2809] = (layer3_outputs[1335]) & ~(layer3_outputs[4739]);
    assign layer4_outputs[2810] = layer3_outputs[4180];
    assign layer4_outputs[2811] = ~((layer3_outputs[2579]) ^ (layer3_outputs[1472]));
    assign layer4_outputs[2812] = ~(layer3_outputs[76]);
    assign layer4_outputs[2813] = ~((layer3_outputs[4168]) | (layer3_outputs[1725]));
    assign layer4_outputs[2814] = ~(layer3_outputs[2687]) | (layer3_outputs[466]);
    assign layer4_outputs[2815] = (layer3_outputs[3126]) & ~(layer3_outputs[205]);
    assign layer4_outputs[2816] = ~(layer3_outputs[4859]) | (layer3_outputs[244]);
    assign layer4_outputs[2817] = ~(layer3_outputs[551]) | (layer3_outputs[1305]);
    assign layer4_outputs[2818] = (layer3_outputs[654]) | (layer3_outputs[3048]);
    assign layer4_outputs[2819] = layer3_outputs[2004];
    assign layer4_outputs[2820] = layer3_outputs[3701];
    assign layer4_outputs[2821] = layer3_outputs[3667];
    assign layer4_outputs[2822] = 1'b0;
    assign layer4_outputs[2823] = ~((layer3_outputs[2888]) | (layer3_outputs[1586]));
    assign layer4_outputs[2824] = layer3_outputs[4441];
    assign layer4_outputs[2825] = layer3_outputs[914];
    assign layer4_outputs[2826] = layer3_outputs[2906];
    assign layer4_outputs[2827] = ~((layer3_outputs[2456]) ^ (layer3_outputs[2067]));
    assign layer4_outputs[2828] = 1'b0;
    assign layer4_outputs[2829] = layer3_outputs[2898];
    assign layer4_outputs[2830] = ~((layer3_outputs[1372]) | (layer3_outputs[246]));
    assign layer4_outputs[2831] = 1'b0;
    assign layer4_outputs[2832] = (layer3_outputs[692]) ^ (layer3_outputs[4210]);
    assign layer4_outputs[2833] = (layer3_outputs[3245]) & ~(layer3_outputs[2716]);
    assign layer4_outputs[2834] = ~((layer3_outputs[2402]) & (layer3_outputs[2257]));
    assign layer4_outputs[2835] = layer3_outputs[2174];
    assign layer4_outputs[2836] = layer3_outputs[607];
    assign layer4_outputs[2837] = (layer3_outputs[1755]) | (layer3_outputs[3756]);
    assign layer4_outputs[2838] = ~(layer3_outputs[2815]);
    assign layer4_outputs[2839] = (layer3_outputs[1737]) & (layer3_outputs[1982]);
    assign layer4_outputs[2840] = (layer3_outputs[74]) & (layer3_outputs[388]);
    assign layer4_outputs[2841] = ~((layer3_outputs[4270]) & (layer3_outputs[136]));
    assign layer4_outputs[2842] = ~((layer3_outputs[2500]) & (layer3_outputs[2509]));
    assign layer4_outputs[2843] = layer3_outputs[4792];
    assign layer4_outputs[2844] = (layer3_outputs[3323]) & ~(layer3_outputs[1007]);
    assign layer4_outputs[2845] = 1'b0;
    assign layer4_outputs[2846] = (layer3_outputs[156]) & (layer3_outputs[1131]);
    assign layer4_outputs[2847] = ~(layer3_outputs[1319]) | (layer3_outputs[835]);
    assign layer4_outputs[2848] = ~(layer3_outputs[1730]) | (layer3_outputs[1064]);
    assign layer4_outputs[2849] = ~(layer3_outputs[4330]);
    assign layer4_outputs[2850] = (layer3_outputs[608]) & ~(layer3_outputs[1588]);
    assign layer4_outputs[2851] = (layer3_outputs[2492]) | (layer3_outputs[622]);
    assign layer4_outputs[2852] = 1'b1;
    assign layer4_outputs[2853] = ~((layer3_outputs[2393]) | (layer3_outputs[2954]));
    assign layer4_outputs[2854] = (layer3_outputs[1468]) & (layer3_outputs[4743]);
    assign layer4_outputs[2855] = layer3_outputs[5058];
    assign layer4_outputs[2856] = (layer3_outputs[3149]) | (layer3_outputs[3153]);
    assign layer4_outputs[2857] = layer3_outputs[4592];
    assign layer4_outputs[2858] = (layer3_outputs[2941]) & ~(layer3_outputs[120]);
    assign layer4_outputs[2859] = layer3_outputs[3611];
    assign layer4_outputs[2860] = 1'b0;
    assign layer4_outputs[2861] = (layer3_outputs[4482]) & (layer3_outputs[3101]);
    assign layer4_outputs[2862] = 1'b1;
    assign layer4_outputs[2863] = ~(layer3_outputs[4001]);
    assign layer4_outputs[2864] = layer3_outputs[3055];
    assign layer4_outputs[2865] = ~((layer3_outputs[2203]) & (layer3_outputs[4424]));
    assign layer4_outputs[2866] = ~(layer3_outputs[2228]) | (layer3_outputs[3782]);
    assign layer4_outputs[2867] = ~((layer3_outputs[474]) & (layer3_outputs[945]));
    assign layer4_outputs[2868] = ~(layer3_outputs[2432]);
    assign layer4_outputs[2869] = ~((layer3_outputs[4300]) | (layer3_outputs[2968]));
    assign layer4_outputs[2870] = ~(layer3_outputs[3075]);
    assign layer4_outputs[2871] = ~(layer3_outputs[4544]);
    assign layer4_outputs[2872] = ~(layer3_outputs[2841]) | (layer3_outputs[2672]);
    assign layer4_outputs[2873] = (layer3_outputs[3333]) ^ (layer3_outputs[951]);
    assign layer4_outputs[2874] = 1'b1;
    assign layer4_outputs[2875] = layer3_outputs[1687];
    assign layer4_outputs[2876] = layer3_outputs[2639];
    assign layer4_outputs[2877] = (layer3_outputs[1799]) & ~(layer3_outputs[3013]);
    assign layer4_outputs[2878] = (layer3_outputs[1292]) & ~(layer3_outputs[1192]);
    assign layer4_outputs[2879] = (layer3_outputs[4608]) ^ (layer3_outputs[1707]);
    assign layer4_outputs[2880] = ~(layer3_outputs[2798]);
    assign layer4_outputs[2881] = 1'b1;
    assign layer4_outputs[2882] = ~(layer3_outputs[587]);
    assign layer4_outputs[2883] = ~(layer3_outputs[557]) | (layer3_outputs[3219]);
    assign layer4_outputs[2884] = (layer3_outputs[2770]) & ~(layer3_outputs[1197]);
    assign layer4_outputs[2885] = (layer3_outputs[1287]) & ~(layer3_outputs[4508]);
    assign layer4_outputs[2886] = layer3_outputs[3475];
    assign layer4_outputs[2887] = (layer3_outputs[1109]) & (layer3_outputs[2688]);
    assign layer4_outputs[2888] = (layer3_outputs[4328]) | (layer3_outputs[1392]);
    assign layer4_outputs[2889] = ~(layer3_outputs[1445]);
    assign layer4_outputs[2890] = ~((layer3_outputs[4688]) | (layer3_outputs[1293]));
    assign layer4_outputs[2891] = (layer3_outputs[671]) & ~(layer3_outputs[297]);
    assign layer4_outputs[2892] = layer3_outputs[1199];
    assign layer4_outputs[2893] = ~(layer3_outputs[4661]) | (layer3_outputs[3452]);
    assign layer4_outputs[2894] = (layer3_outputs[2146]) & ~(layer3_outputs[1412]);
    assign layer4_outputs[2895] = (layer3_outputs[488]) & (layer3_outputs[4611]);
    assign layer4_outputs[2896] = (layer3_outputs[1688]) & ~(layer3_outputs[5013]);
    assign layer4_outputs[2897] = ~(layer3_outputs[963]);
    assign layer4_outputs[2898] = layer3_outputs[3686];
    assign layer4_outputs[2899] = layer3_outputs[4023];
    assign layer4_outputs[2900] = ~(layer3_outputs[680]) | (layer3_outputs[2813]);
    assign layer4_outputs[2901] = ~(layer3_outputs[4323]);
    assign layer4_outputs[2902] = ~((layer3_outputs[4324]) | (layer3_outputs[268]));
    assign layer4_outputs[2903] = (layer3_outputs[3378]) ^ (layer3_outputs[170]);
    assign layer4_outputs[2904] = layer3_outputs[426];
    assign layer4_outputs[2905] = layer3_outputs[3511];
    assign layer4_outputs[2906] = ~(layer3_outputs[5046]) | (layer3_outputs[5064]);
    assign layer4_outputs[2907] = layer3_outputs[4625];
    assign layer4_outputs[2908] = (layer3_outputs[2853]) | (layer3_outputs[5108]);
    assign layer4_outputs[2909] = layer3_outputs[307];
    assign layer4_outputs[2910] = ~(layer3_outputs[429]) | (layer3_outputs[5036]);
    assign layer4_outputs[2911] = ~(layer3_outputs[4651]) | (layer3_outputs[2485]);
    assign layer4_outputs[2912] = ~((layer3_outputs[3186]) | (layer3_outputs[4312]));
    assign layer4_outputs[2913] = ~((layer3_outputs[3584]) & (layer3_outputs[3014]));
    assign layer4_outputs[2914] = (layer3_outputs[3836]) & ~(layer3_outputs[3840]);
    assign layer4_outputs[2915] = (layer3_outputs[2949]) & ~(layer3_outputs[1251]);
    assign layer4_outputs[2916] = (layer3_outputs[517]) | (layer3_outputs[2914]);
    assign layer4_outputs[2917] = (layer3_outputs[1097]) & (layer3_outputs[1460]);
    assign layer4_outputs[2918] = 1'b0;
    assign layer4_outputs[2919] = (layer3_outputs[2384]) ^ (layer3_outputs[586]);
    assign layer4_outputs[2920] = layer3_outputs[1520];
    assign layer4_outputs[2921] = 1'b1;
    assign layer4_outputs[2922] = (layer3_outputs[4333]) & ~(layer3_outputs[664]);
    assign layer4_outputs[2923] = ~((layer3_outputs[3682]) & (layer3_outputs[2530]));
    assign layer4_outputs[2924] = layer3_outputs[4038];
    assign layer4_outputs[2925] = ~(layer3_outputs[2224]);
    assign layer4_outputs[2926] = ~(layer3_outputs[857]) | (layer3_outputs[4215]);
    assign layer4_outputs[2927] = ~(layer3_outputs[2863]) | (layer3_outputs[5018]);
    assign layer4_outputs[2928] = ~(layer3_outputs[1596]) | (layer3_outputs[2601]);
    assign layer4_outputs[2929] = ~(layer3_outputs[2859]);
    assign layer4_outputs[2930] = (layer3_outputs[858]) | (layer3_outputs[3746]);
    assign layer4_outputs[2931] = (layer3_outputs[361]) | (layer3_outputs[747]);
    assign layer4_outputs[2932] = layer3_outputs[3792];
    assign layer4_outputs[2933] = layer3_outputs[4554];
    assign layer4_outputs[2934] = layer3_outputs[1012];
    assign layer4_outputs[2935] = layer3_outputs[4068];
    assign layer4_outputs[2936] = 1'b0;
    assign layer4_outputs[2937] = ~(layer3_outputs[3200]) | (layer3_outputs[2413]);
    assign layer4_outputs[2938] = 1'b0;
    assign layer4_outputs[2939] = ~(layer3_outputs[1005]);
    assign layer4_outputs[2940] = (layer3_outputs[4491]) & ~(layer3_outputs[2946]);
    assign layer4_outputs[2941] = (layer3_outputs[2317]) & ~(layer3_outputs[4214]);
    assign layer4_outputs[2942] = (layer3_outputs[1613]) ^ (layer3_outputs[2380]);
    assign layer4_outputs[2943] = ~(layer3_outputs[2499]);
    assign layer4_outputs[2944] = layer3_outputs[5002];
    assign layer4_outputs[2945] = ~(layer3_outputs[3855]) | (layer3_outputs[3269]);
    assign layer4_outputs[2946] = (layer3_outputs[1185]) | (layer3_outputs[4733]);
    assign layer4_outputs[2947] = ~((layer3_outputs[4869]) | (layer3_outputs[1454]));
    assign layer4_outputs[2948] = (layer3_outputs[2663]) & ~(layer3_outputs[1630]);
    assign layer4_outputs[2949] = ~(layer3_outputs[5025]);
    assign layer4_outputs[2950] = layer3_outputs[4697];
    assign layer4_outputs[2951] = ~((layer3_outputs[2639]) | (layer3_outputs[3349]));
    assign layer4_outputs[2952] = layer3_outputs[3110];
    assign layer4_outputs[2953] = (layer3_outputs[781]) & ~(layer3_outputs[877]);
    assign layer4_outputs[2954] = ~(layer3_outputs[4546]);
    assign layer4_outputs[2955] = 1'b1;
    assign layer4_outputs[2956] = ~(layer3_outputs[2243]);
    assign layer4_outputs[2957] = layer3_outputs[1820];
    assign layer4_outputs[2958] = ~(layer3_outputs[222]);
    assign layer4_outputs[2959] = layer3_outputs[3730];
    assign layer4_outputs[2960] = layer3_outputs[4208];
    assign layer4_outputs[2961] = (layer3_outputs[146]) ^ (layer3_outputs[3165]);
    assign layer4_outputs[2962] = (layer3_outputs[2491]) & ~(layer3_outputs[3264]);
    assign layer4_outputs[2963] = ~(layer3_outputs[2825]);
    assign layer4_outputs[2964] = 1'b1;
    assign layer4_outputs[2965] = ~((layer3_outputs[5054]) | (layer3_outputs[2290]));
    assign layer4_outputs[2966] = ~(layer3_outputs[659]);
    assign layer4_outputs[2967] = layer3_outputs[1467];
    assign layer4_outputs[2968] = ~(layer3_outputs[1813]) | (layer3_outputs[1853]);
    assign layer4_outputs[2969] = ~(layer3_outputs[516]);
    assign layer4_outputs[2970] = ~(layer3_outputs[292]);
    assign layer4_outputs[2971] = layer3_outputs[708];
    assign layer4_outputs[2972] = layer3_outputs[852];
    assign layer4_outputs[2973] = ~(layer3_outputs[3550]);
    assign layer4_outputs[2974] = (layer3_outputs[1999]) | (layer3_outputs[5038]);
    assign layer4_outputs[2975] = ~(layer3_outputs[1525]) | (layer3_outputs[3281]);
    assign layer4_outputs[2976] = ~(layer3_outputs[1240]);
    assign layer4_outputs[2977] = ~((layer3_outputs[1145]) & (layer3_outputs[2873]));
    assign layer4_outputs[2978] = (layer3_outputs[265]) ^ (layer3_outputs[326]);
    assign layer4_outputs[2979] = ~(layer3_outputs[67]);
    assign layer4_outputs[2980] = ~(layer3_outputs[1461]);
    assign layer4_outputs[2981] = ~(layer3_outputs[2910]);
    assign layer4_outputs[2982] = ~(layer3_outputs[1604]);
    assign layer4_outputs[2983] = ~((layer3_outputs[2812]) ^ (layer3_outputs[1202]));
    assign layer4_outputs[2984] = ~(layer3_outputs[3150]) | (layer3_outputs[510]);
    assign layer4_outputs[2985] = layer3_outputs[2921];
    assign layer4_outputs[2986] = ~(layer3_outputs[1188]);
    assign layer4_outputs[2987] = (layer3_outputs[4577]) & ~(layer3_outputs[4606]);
    assign layer4_outputs[2988] = (layer3_outputs[1636]) ^ (layer3_outputs[4126]);
    assign layer4_outputs[2989] = ~(layer3_outputs[1987]) | (layer3_outputs[4564]);
    assign layer4_outputs[2990] = ~(layer3_outputs[1173]);
    assign layer4_outputs[2991] = ~(layer3_outputs[4833]) | (layer3_outputs[870]);
    assign layer4_outputs[2992] = layer3_outputs[2683];
    assign layer4_outputs[2993] = ~(layer3_outputs[4811]) | (layer3_outputs[4359]);
    assign layer4_outputs[2994] = (layer3_outputs[1313]) & ~(layer3_outputs[3397]);
    assign layer4_outputs[2995] = layer3_outputs[3913];
    assign layer4_outputs[2996] = layer3_outputs[2563];
    assign layer4_outputs[2997] = ~(layer3_outputs[4245]);
    assign layer4_outputs[2998] = layer3_outputs[1230];
    assign layer4_outputs[2999] = ~(layer3_outputs[3017]);
    assign layer4_outputs[3000] = ~((layer3_outputs[3783]) | (layer3_outputs[599]));
    assign layer4_outputs[3001] = ~((layer3_outputs[186]) & (layer3_outputs[4057]));
    assign layer4_outputs[3002] = layer3_outputs[4585];
    assign layer4_outputs[3003] = ~((layer3_outputs[4553]) | (layer3_outputs[5114]));
    assign layer4_outputs[3004] = layer3_outputs[1044];
    assign layer4_outputs[3005] = (layer3_outputs[3996]) & (layer3_outputs[5101]);
    assign layer4_outputs[3006] = layer3_outputs[1082];
    assign layer4_outputs[3007] = ~((layer3_outputs[4155]) ^ (layer3_outputs[1372]));
    assign layer4_outputs[3008] = layer3_outputs[517];
    assign layer4_outputs[3009] = layer3_outputs[1691];
    assign layer4_outputs[3010] = 1'b0;
    assign layer4_outputs[3011] = ~(layer3_outputs[3510]);
    assign layer4_outputs[3012] = ~((layer3_outputs[4547]) & (layer3_outputs[3583]));
    assign layer4_outputs[3013] = (layer3_outputs[1338]) | (layer3_outputs[2617]);
    assign layer4_outputs[3014] = ~((layer3_outputs[941]) ^ (layer3_outputs[2665]));
    assign layer4_outputs[3015] = layer3_outputs[2465];
    assign layer4_outputs[3016] = (layer3_outputs[2241]) ^ (layer3_outputs[445]);
    assign layer4_outputs[3017] = (layer3_outputs[1570]) & ~(layer3_outputs[1883]);
    assign layer4_outputs[3018] = ~(layer3_outputs[3639]);
    assign layer4_outputs[3019] = layer3_outputs[3147];
    assign layer4_outputs[3020] = ~((layer3_outputs[3681]) & (layer3_outputs[2509]));
    assign layer4_outputs[3021] = ~(layer3_outputs[2588]);
    assign layer4_outputs[3022] = ~(layer3_outputs[1308]);
    assign layer4_outputs[3023] = ~((layer3_outputs[515]) & (layer3_outputs[2964]));
    assign layer4_outputs[3024] = layer3_outputs[2607];
    assign layer4_outputs[3025] = ~(layer3_outputs[4812]);
    assign layer4_outputs[3026] = layer3_outputs[4778];
    assign layer4_outputs[3027] = (layer3_outputs[3006]) ^ (layer3_outputs[125]);
    assign layer4_outputs[3028] = 1'b0;
    assign layer4_outputs[3029] = ~(layer3_outputs[2432]);
    assign layer4_outputs[3030] = layer3_outputs[1717];
    assign layer4_outputs[3031] = (layer3_outputs[1645]) ^ (layer3_outputs[1141]);
    assign layer4_outputs[3032] = ~(layer3_outputs[3326]);
    assign layer4_outputs[3033] = layer3_outputs[1509];
    assign layer4_outputs[3034] = layer3_outputs[2483];
    assign layer4_outputs[3035] = layer3_outputs[1408];
    assign layer4_outputs[3036] = ~(layer3_outputs[3305]);
    assign layer4_outputs[3037] = (layer3_outputs[2628]) | (layer3_outputs[4094]);
    assign layer4_outputs[3038] = layer3_outputs[4674];
    assign layer4_outputs[3039] = ~(layer3_outputs[298]) | (layer3_outputs[789]);
    assign layer4_outputs[3040] = layer3_outputs[3432];
    assign layer4_outputs[3041] = (layer3_outputs[2439]) & ~(layer3_outputs[4852]);
    assign layer4_outputs[3042] = (layer3_outputs[1589]) | (layer3_outputs[1010]);
    assign layer4_outputs[3043] = ~(layer3_outputs[4419]);
    assign layer4_outputs[3044] = ~(layer3_outputs[2725]);
    assign layer4_outputs[3045] = ~(layer3_outputs[4085]) | (layer3_outputs[2121]);
    assign layer4_outputs[3046] = ~((layer3_outputs[4314]) & (layer3_outputs[1272]));
    assign layer4_outputs[3047] = (layer3_outputs[669]) & (layer3_outputs[3478]);
    assign layer4_outputs[3048] = layer3_outputs[4303];
    assign layer4_outputs[3049] = (layer3_outputs[1077]) ^ (layer3_outputs[223]);
    assign layer4_outputs[3050] = ~((layer3_outputs[1661]) | (layer3_outputs[4822]));
    assign layer4_outputs[3051] = (layer3_outputs[1078]) & (layer3_outputs[2097]);
    assign layer4_outputs[3052] = ~(layer3_outputs[3446]);
    assign layer4_outputs[3053] = ~(layer3_outputs[3917]);
    assign layer4_outputs[3054] = ~(layer3_outputs[4594]);
    assign layer4_outputs[3055] = ~(layer3_outputs[443]) | (layer3_outputs[949]);
    assign layer4_outputs[3056] = 1'b1;
    assign layer4_outputs[3057] = layer3_outputs[528];
    assign layer4_outputs[3058] = ~(layer3_outputs[699]) | (layer3_outputs[804]);
    assign layer4_outputs[3059] = layer3_outputs[536];
    assign layer4_outputs[3060] = (layer3_outputs[369]) & (layer3_outputs[3051]);
    assign layer4_outputs[3061] = layer3_outputs[4714];
    assign layer4_outputs[3062] = layer3_outputs[1033];
    assign layer4_outputs[3063] = ~(layer3_outputs[4928]);
    assign layer4_outputs[3064] = ~(layer3_outputs[2987]);
    assign layer4_outputs[3065] = (layer3_outputs[405]) | (layer3_outputs[384]);
    assign layer4_outputs[3066] = (layer3_outputs[4661]) & ~(layer3_outputs[3379]);
    assign layer4_outputs[3067] = ~((layer3_outputs[4022]) | (layer3_outputs[4666]));
    assign layer4_outputs[3068] = ~(layer3_outputs[310]);
    assign layer4_outputs[3069] = (layer3_outputs[3394]) & (layer3_outputs[4143]);
    assign layer4_outputs[3070] = ~((layer3_outputs[394]) & (layer3_outputs[4089]));
    assign layer4_outputs[3071] = 1'b0;
    assign layer4_outputs[3072] = ~(layer3_outputs[1403]) | (layer3_outputs[3793]);
    assign layer4_outputs[3073] = layer3_outputs[2212];
    assign layer4_outputs[3074] = layer3_outputs[4055];
    assign layer4_outputs[3075] = (layer3_outputs[1742]) & ~(layer3_outputs[867]);
    assign layer4_outputs[3076] = ~(layer3_outputs[4574]);
    assign layer4_outputs[3077] = ~((layer3_outputs[1577]) | (layer3_outputs[3170]));
    assign layer4_outputs[3078] = ~(layer3_outputs[243]) | (layer3_outputs[751]);
    assign layer4_outputs[3079] = layer3_outputs[2905];
    assign layer4_outputs[3080] = (layer3_outputs[4882]) & ~(layer3_outputs[142]);
    assign layer4_outputs[3081] = ~((layer3_outputs[162]) & (layer3_outputs[2932]));
    assign layer4_outputs[3082] = 1'b1;
    assign layer4_outputs[3083] = ~((layer3_outputs[2399]) | (layer3_outputs[3898]));
    assign layer4_outputs[3084] = ~((layer3_outputs[721]) | (layer3_outputs[2841]));
    assign layer4_outputs[3085] = (layer3_outputs[3636]) & (layer3_outputs[2582]);
    assign layer4_outputs[3086] = ~((layer3_outputs[3333]) & (layer3_outputs[1577]));
    assign layer4_outputs[3087] = ~((layer3_outputs[3886]) | (layer3_outputs[28]));
    assign layer4_outputs[3088] = (layer3_outputs[2845]) ^ (layer3_outputs[3935]);
    assign layer4_outputs[3089] = ~(layer3_outputs[3597]) | (layer3_outputs[2252]);
    assign layer4_outputs[3090] = layer3_outputs[1426];
    assign layer4_outputs[3091] = ~(layer3_outputs[2178]);
    assign layer4_outputs[3092] = ~(layer3_outputs[1201]) | (layer3_outputs[2736]);
    assign layer4_outputs[3093] = ~(layer3_outputs[3729]) | (layer3_outputs[442]);
    assign layer4_outputs[3094] = 1'b0;
    assign layer4_outputs[3095] = ~((layer3_outputs[2947]) | (layer3_outputs[4675]));
    assign layer4_outputs[3096] = layer3_outputs[2457];
    assign layer4_outputs[3097] = layer3_outputs[2203];
    assign layer4_outputs[3098] = layer3_outputs[4441];
    assign layer4_outputs[3099] = ~(layer3_outputs[825]);
    assign layer4_outputs[3100] = layer3_outputs[4934];
    assign layer4_outputs[3101] = (layer3_outputs[4074]) | (layer3_outputs[3409]);
    assign layer4_outputs[3102] = (layer3_outputs[3694]) & ~(layer3_outputs[2152]);
    assign layer4_outputs[3103] = ~((layer3_outputs[4468]) | (layer3_outputs[4403]));
    assign layer4_outputs[3104] = (layer3_outputs[2309]) ^ (layer3_outputs[2089]);
    assign layer4_outputs[3105] = ~(layer3_outputs[2154]) | (layer3_outputs[2675]);
    assign layer4_outputs[3106] = (layer3_outputs[176]) & ~(layer3_outputs[3408]);
    assign layer4_outputs[3107] = layer3_outputs[340];
    assign layer4_outputs[3108] = ~(layer3_outputs[2058]);
    assign layer4_outputs[3109] = layer3_outputs[1922];
    assign layer4_outputs[3110] = layer3_outputs[2700];
    assign layer4_outputs[3111] = (layer3_outputs[250]) & ~(layer3_outputs[3092]);
    assign layer4_outputs[3112] = ~(layer3_outputs[2723]);
    assign layer4_outputs[3113] = ~((layer3_outputs[2440]) & (layer3_outputs[620]));
    assign layer4_outputs[3114] = layer3_outputs[1072];
    assign layer4_outputs[3115] = ~(layer3_outputs[2466]) | (layer3_outputs[622]);
    assign layer4_outputs[3116] = layer3_outputs[3726];
    assign layer4_outputs[3117] = (layer3_outputs[2945]) & (layer3_outputs[1484]);
    assign layer4_outputs[3118] = (layer3_outputs[3494]) & ~(layer3_outputs[4201]);
    assign layer4_outputs[3119] = ~((layer3_outputs[2135]) | (layer3_outputs[4339]));
    assign layer4_outputs[3120] = ~(layer3_outputs[4431]);
    assign layer4_outputs[3121] = 1'b0;
    assign layer4_outputs[3122] = ~((layer3_outputs[1983]) & (layer3_outputs[2729]));
    assign layer4_outputs[3123] = ~(layer3_outputs[3541]) | (layer3_outputs[2069]);
    assign layer4_outputs[3124] = ~((layer3_outputs[1942]) & (layer3_outputs[5055]));
    assign layer4_outputs[3125] = (layer3_outputs[3609]) | (layer3_outputs[4964]);
    assign layer4_outputs[3126] = ~(layer3_outputs[3819]);
    assign layer4_outputs[3127] = (layer3_outputs[4827]) & ~(layer3_outputs[943]);
    assign layer4_outputs[3128] = layer3_outputs[421];
    assign layer4_outputs[3129] = layer3_outputs[3847];
    assign layer4_outputs[3130] = (layer3_outputs[674]) & ~(layer3_outputs[1331]);
    assign layer4_outputs[3131] = ~(layer3_outputs[4835]);
    assign layer4_outputs[3132] = layer3_outputs[2557];
    assign layer4_outputs[3133] = (layer3_outputs[715]) & (layer3_outputs[1247]);
    assign layer4_outputs[3134] = layer3_outputs[4811];
    assign layer4_outputs[3135] = ~(layer3_outputs[3885]);
    assign layer4_outputs[3136] = ~((layer3_outputs[3718]) & (layer3_outputs[3899]));
    assign layer4_outputs[3137] = ~((layer3_outputs[1181]) ^ (layer3_outputs[291]));
    assign layer4_outputs[3138] = (layer3_outputs[758]) & ~(layer3_outputs[4051]);
    assign layer4_outputs[3139] = (layer3_outputs[2819]) & (layer3_outputs[294]);
    assign layer4_outputs[3140] = layer3_outputs[2929];
    assign layer4_outputs[3141] = ~(layer3_outputs[4581]);
    assign layer4_outputs[3142] = ~((layer3_outputs[4900]) & (layer3_outputs[4532]));
    assign layer4_outputs[3143] = (layer3_outputs[1343]) | (layer3_outputs[4725]);
    assign layer4_outputs[3144] = layer3_outputs[3901];
    assign layer4_outputs[3145] = layer3_outputs[1791];
    assign layer4_outputs[3146] = ~(layer3_outputs[4834]) | (layer3_outputs[2232]);
    assign layer4_outputs[3147] = ~(layer3_outputs[2046]);
    assign layer4_outputs[3148] = ~(layer3_outputs[1395]);
    assign layer4_outputs[3149] = (layer3_outputs[5026]) & ~(layer3_outputs[3894]);
    assign layer4_outputs[3150] = (layer3_outputs[4560]) ^ (layer3_outputs[2971]);
    assign layer4_outputs[3151] = ~(layer3_outputs[1272]) | (layer3_outputs[3507]);
    assign layer4_outputs[3152] = (layer3_outputs[3934]) | (layer3_outputs[4815]);
    assign layer4_outputs[3153] = layer3_outputs[1354];
    assign layer4_outputs[3154] = ~((layer3_outputs[2751]) & (layer3_outputs[3248]));
    assign layer4_outputs[3155] = ~(layer3_outputs[2747]) | (layer3_outputs[4891]);
    assign layer4_outputs[3156] = ~((layer3_outputs[3411]) | (layer3_outputs[3350]));
    assign layer4_outputs[3157] = layer3_outputs[3730];
    assign layer4_outputs[3158] = ~(layer3_outputs[4369]);
    assign layer4_outputs[3159] = (layer3_outputs[4265]) ^ (layer3_outputs[783]);
    assign layer4_outputs[3160] = 1'b0;
    assign layer4_outputs[3161] = layer3_outputs[1083];
    assign layer4_outputs[3162] = layer3_outputs[4727];
    assign layer4_outputs[3163] = (layer3_outputs[1170]) & (layer3_outputs[1387]);
    assign layer4_outputs[3164] = ~(layer3_outputs[4469]) | (layer3_outputs[4217]);
    assign layer4_outputs[3165] = ~((layer3_outputs[4534]) | (layer3_outputs[2638]));
    assign layer4_outputs[3166] = layer3_outputs[4886];
    assign layer4_outputs[3167] = layer3_outputs[3951];
    assign layer4_outputs[3168] = (layer3_outputs[4485]) ^ (layer3_outputs[544]);
    assign layer4_outputs[3169] = ~(layer3_outputs[3039]) | (layer3_outputs[3788]);
    assign layer4_outputs[3170] = 1'b1;
    assign layer4_outputs[3171] = ~((layer3_outputs[4302]) | (layer3_outputs[1343]));
    assign layer4_outputs[3172] = (layer3_outputs[826]) ^ (layer3_outputs[1444]);
    assign layer4_outputs[3173] = ~((layer3_outputs[4291]) & (layer3_outputs[5010]));
    assign layer4_outputs[3174] = (layer3_outputs[3970]) ^ (layer3_outputs[547]);
    assign layer4_outputs[3175] = ~(layer3_outputs[2786]) | (layer3_outputs[595]);
    assign layer4_outputs[3176] = 1'b1;
    assign layer4_outputs[3177] = layer3_outputs[3731];
    assign layer4_outputs[3178] = ~((layer3_outputs[3620]) | (layer3_outputs[82]));
    assign layer4_outputs[3179] = (layer3_outputs[4238]) | (layer3_outputs[911]);
    assign layer4_outputs[3180] = layer3_outputs[4657];
    assign layer4_outputs[3181] = layer3_outputs[2015];
    assign layer4_outputs[3182] = layer3_outputs[2825];
    assign layer4_outputs[3183] = 1'b1;
    assign layer4_outputs[3184] = ~((layer3_outputs[5073]) | (layer3_outputs[4445]));
    assign layer4_outputs[3185] = (layer3_outputs[3907]) & ~(layer3_outputs[2788]);
    assign layer4_outputs[3186] = ~((layer3_outputs[3335]) ^ (layer3_outputs[4683]));
    assign layer4_outputs[3187] = layer3_outputs[3137];
    assign layer4_outputs[3188] = 1'b1;
    assign layer4_outputs[3189] = ~((layer3_outputs[204]) | (layer3_outputs[315]));
    assign layer4_outputs[3190] = layer3_outputs[1912];
    assign layer4_outputs[3191] = ~(layer3_outputs[3985]) | (layer3_outputs[4014]);
    assign layer4_outputs[3192] = ~(layer3_outputs[3888]);
    assign layer4_outputs[3193] = ~(layer3_outputs[1430]) | (layer3_outputs[3671]);
    assign layer4_outputs[3194] = ~((layer3_outputs[4102]) & (layer3_outputs[3826]));
    assign layer4_outputs[3195] = layer3_outputs[3289];
    assign layer4_outputs[3196] = 1'b0;
    assign layer4_outputs[3197] = ~(layer3_outputs[3259]);
    assign layer4_outputs[3198] = 1'b1;
    assign layer4_outputs[3199] = ~(layer3_outputs[5029]);
    assign layer4_outputs[3200] = (layer3_outputs[84]) & ~(layer3_outputs[4568]);
    assign layer4_outputs[3201] = 1'b0;
    assign layer4_outputs[3202] = ~(layer3_outputs[936]);
    assign layer4_outputs[3203] = ~((layer3_outputs[395]) ^ (layer3_outputs[3660]));
    assign layer4_outputs[3204] = ~(layer3_outputs[155]) | (layer3_outputs[2990]);
    assign layer4_outputs[3205] = ~(layer3_outputs[907]) | (layer3_outputs[984]);
    assign layer4_outputs[3206] = ~(layer3_outputs[2256]) | (layer3_outputs[1193]);
    assign layer4_outputs[3207] = ~(layer3_outputs[5103]);
    assign layer4_outputs[3208] = (layer3_outputs[4526]) & ~(layer3_outputs[641]);
    assign layer4_outputs[3209] = ~(layer3_outputs[307]);
    assign layer4_outputs[3210] = ~(layer3_outputs[2060]);
    assign layer4_outputs[3211] = ~(layer3_outputs[2441]) | (layer3_outputs[1968]);
    assign layer4_outputs[3212] = ~(layer3_outputs[4798]);
    assign layer4_outputs[3213] = ~(layer3_outputs[725]) | (layer3_outputs[3057]);
    assign layer4_outputs[3214] = (layer3_outputs[2957]) | (layer3_outputs[2037]);
    assign layer4_outputs[3215] = (layer3_outputs[1873]) | (layer3_outputs[5074]);
    assign layer4_outputs[3216] = ~((layer3_outputs[3021]) ^ (layer3_outputs[2860]));
    assign layer4_outputs[3217] = ~(layer3_outputs[3817]);
    assign layer4_outputs[3218] = (layer3_outputs[339]) | (layer3_outputs[2433]);
    assign layer4_outputs[3219] = ~(layer3_outputs[1932]) | (layer3_outputs[3656]);
    assign layer4_outputs[3220] = ~(layer3_outputs[4663]);
    assign layer4_outputs[3221] = (layer3_outputs[1052]) & ~(layer3_outputs[3750]);
    assign layer4_outputs[3222] = ~(layer3_outputs[2244]) | (layer3_outputs[915]);
    assign layer4_outputs[3223] = (layer3_outputs[3879]) & (layer3_outputs[503]);
    assign layer4_outputs[3224] = 1'b0;
    assign layer4_outputs[3225] = ~(layer3_outputs[1920]);
    assign layer4_outputs[3226] = ~(layer3_outputs[359]);
    assign layer4_outputs[3227] = (layer3_outputs[1298]) & (layer3_outputs[3376]);
    assign layer4_outputs[3228] = ~(layer3_outputs[4769]) | (layer3_outputs[4182]);
    assign layer4_outputs[3229] = layer3_outputs[1310];
    assign layer4_outputs[3230] = 1'b0;
    assign layer4_outputs[3231] = layer3_outputs[277];
    assign layer4_outputs[3232] = (layer3_outputs[1083]) & (layer3_outputs[1087]);
    assign layer4_outputs[3233] = layer3_outputs[449];
    assign layer4_outputs[3234] = (layer3_outputs[7]) & ~(layer3_outputs[1326]);
    assign layer4_outputs[3235] = ~(layer3_outputs[2892]);
    assign layer4_outputs[3236] = (layer3_outputs[2153]) ^ (layer3_outputs[2857]);
    assign layer4_outputs[3237] = 1'b1;
    assign layer4_outputs[3238] = ~(layer3_outputs[3240]);
    assign layer4_outputs[3239] = ~(layer3_outputs[3040]) | (layer3_outputs[3923]);
    assign layer4_outputs[3240] = layer3_outputs[2142];
    assign layer4_outputs[3241] = (layer3_outputs[440]) ^ (layer3_outputs[1026]);
    assign layer4_outputs[3242] = layer3_outputs[3354];
    assign layer4_outputs[3243] = (layer3_outputs[1253]) ^ (layer3_outputs[3715]);
    assign layer4_outputs[3244] = (layer3_outputs[1302]) & (layer3_outputs[2671]);
    assign layer4_outputs[3245] = layer3_outputs[1736];
    assign layer4_outputs[3246] = ~(layer3_outputs[1673]);
    assign layer4_outputs[3247] = layer3_outputs[2581];
    assign layer4_outputs[3248] = (layer3_outputs[2469]) & (layer3_outputs[181]);
    assign layer4_outputs[3249] = layer3_outputs[4462];
    assign layer4_outputs[3250] = ~(layer3_outputs[3555]) | (layer3_outputs[2032]);
    assign layer4_outputs[3251] = layer3_outputs[2863];
    assign layer4_outputs[3252] = ~(layer3_outputs[2123]);
    assign layer4_outputs[3253] = ~(layer3_outputs[2748]);
    assign layer4_outputs[3254] = (layer3_outputs[4817]) & ~(layer3_outputs[4509]);
    assign layer4_outputs[3255] = (layer3_outputs[5068]) | (layer3_outputs[3372]);
    assign layer4_outputs[3256] = layer3_outputs[3365];
    assign layer4_outputs[3257] = layer3_outputs[2185];
    assign layer4_outputs[3258] = (layer3_outputs[2503]) | (layer3_outputs[1196]);
    assign layer4_outputs[3259] = ~((layer3_outputs[283]) & (layer3_outputs[3679]));
    assign layer4_outputs[3260] = layer3_outputs[1032];
    assign layer4_outputs[3261] = layer3_outputs[2193];
    assign layer4_outputs[3262] = layer3_outputs[3079];
    assign layer4_outputs[3263] = layer3_outputs[671];
    assign layer4_outputs[3264] = layer3_outputs[4947];
    assign layer4_outputs[3265] = (layer3_outputs[2699]) ^ (layer3_outputs[2010]);
    assign layer4_outputs[3266] = ~(layer3_outputs[4037]) | (layer3_outputs[799]);
    assign layer4_outputs[3267] = 1'b1;
    assign layer4_outputs[3268] = layer3_outputs[2122];
    assign layer4_outputs[3269] = layer3_outputs[4638];
    assign layer4_outputs[3270] = layer3_outputs[5106];
    assign layer4_outputs[3271] = ~(layer3_outputs[2452]) | (layer3_outputs[35]);
    assign layer4_outputs[3272] = ~((layer3_outputs[4413]) ^ (layer3_outputs[2485]));
    assign layer4_outputs[3273] = ~(layer3_outputs[1513]);
    assign layer4_outputs[3274] = (layer3_outputs[639]) | (layer3_outputs[1622]);
    assign layer4_outputs[3275] = ~(layer3_outputs[1806]);
    assign layer4_outputs[3276] = ~((layer3_outputs[363]) | (layer3_outputs[3821]));
    assign layer4_outputs[3277] = ~(layer3_outputs[2166]);
    assign layer4_outputs[3278] = layer3_outputs[2347];
    assign layer4_outputs[3279] = layer3_outputs[749];
    assign layer4_outputs[3280] = layer3_outputs[1568];
    assign layer4_outputs[3281] = ~(layer3_outputs[3012]);
    assign layer4_outputs[3282] = layer3_outputs[4608];
    assign layer4_outputs[3283] = ~(layer3_outputs[267]);
    assign layer4_outputs[3284] = ~(layer3_outputs[2021]) | (layer3_outputs[1881]);
    assign layer4_outputs[3285] = ~(layer3_outputs[3319]);
    assign layer4_outputs[3286] = 1'b1;
    assign layer4_outputs[3287] = ~(layer3_outputs[2769]);
    assign layer4_outputs[3288] = ~(layer3_outputs[2370]);
    assign layer4_outputs[3289] = ~(layer3_outputs[2103]);
    assign layer4_outputs[3290] = ~(layer3_outputs[1364]);
    assign layer4_outputs[3291] = ~(layer3_outputs[1334]) | (layer3_outputs[1842]);
    assign layer4_outputs[3292] = (layer3_outputs[1189]) & (layer3_outputs[390]);
    assign layer4_outputs[3293] = layer3_outputs[4982];
    assign layer4_outputs[3294] = ~(layer3_outputs[4580]);
    assign layer4_outputs[3295] = ~(layer3_outputs[5088]);
    assign layer4_outputs[3296] = ~(layer3_outputs[1773]);
    assign layer4_outputs[3297] = ~(layer3_outputs[4232]);
    assign layer4_outputs[3298] = ~((layer3_outputs[3608]) | (layer3_outputs[686]));
    assign layer4_outputs[3299] = layer3_outputs[1263];
    assign layer4_outputs[3300] = ~((layer3_outputs[960]) & (layer3_outputs[2955]));
    assign layer4_outputs[3301] = ~(layer3_outputs[377]) | (layer3_outputs[1390]);
    assign layer4_outputs[3302] = (layer3_outputs[496]) & (layer3_outputs[1602]);
    assign layer4_outputs[3303] = layer3_outputs[55];
    assign layer4_outputs[3304] = (layer3_outputs[682]) & ~(layer3_outputs[612]);
    assign layer4_outputs[3305] = ~(layer3_outputs[3669]);
    assign layer4_outputs[3306] = layer3_outputs[2838];
    assign layer4_outputs[3307] = ~((layer3_outputs[2604]) | (layer3_outputs[302]));
    assign layer4_outputs[3308] = layer3_outputs[3711];
    assign layer4_outputs[3309] = ~(layer3_outputs[3690]);
    assign layer4_outputs[3310] = ~(layer3_outputs[2944]);
    assign layer4_outputs[3311] = (layer3_outputs[2253]) & (layer3_outputs[1436]);
    assign layer4_outputs[3312] = ~(layer3_outputs[4194]) | (layer3_outputs[36]);
    assign layer4_outputs[3313] = ~((layer3_outputs[2729]) ^ (layer3_outputs[2174]));
    assign layer4_outputs[3314] = layer3_outputs[3946];
    assign layer4_outputs[3315] = layer3_outputs[1766];
    assign layer4_outputs[3316] = layer3_outputs[4735];
    assign layer4_outputs[3317] = layer3_outputs[4417];
    assign layer4_outputs[3318] = (layer3_outputs[651]) ^ (layer3_outputs[2862]);
    assign layer4_outputs[3319] = ~(layer3_outputs[3744]);
    assign layer4_outputs[3320] = ~(layer3_outputs[4235]) | (layer3_outputs[3160]);
    assign layer4_outputs[3321] = ~(layer3_outputs[1769]) | (layer3_outputs[880]);
    assign layer4_outputs[3322] = 1'b1;
    assign layer4_outputs[3323] = layer3_outputs[1466];
    assign layer4_outputs[3324] = ~((layer3_outputs[3573]) ^ (layer3_outputs[367]));
    assign layer4_outputs[3325] = 1'b1;
    assign layer4_outputs[3326] = (layer3_outputs[3524]) & ~(layer3_outputs[4666]);
    assign layer4_outputs[3327] = (layer3_outputs[815]) & ~(layer3_outputs[1594]);
    assign layer4_outputs[3328] = layer3_outputs[1360];
    assign layer4_outputs[3329] = (layer3_outputs[4315]) & ~(layer3_outputs[1665]);
    assign layer4_outputs[3330] = (layer3_outputs[4647]) & (layer3_outputs[3022]);
    assign layer4_outputs[3331] = layer3_outputs[2953];
    assign layer4_outputs[3332] = ~(layer3_outputs[3038]);
    assign layer4_outputs[3333] = layer3_outputs[4351];
    assign layer4_outputs[3334] = (layer3_outputs[979]) & (layer3_outputs[3695]);
    assign layer4_outputs[3335] = ~(layer3_outputs[4317]);
    assign layer4_outputs[3336] = ~(layer3_outputs[4865]);
    assign layer4_outputs[3337] = layer3_outputs[3883];
    assign layer4_outputs[3338] = (layer3_outputs[3457]) & (layer3_outputs[4199]);
    assign layer4_outputs[3339] = ~(layer3_outputs[1500]) | (layer3_outputs[519]);
    assign layer4_outputs[3340] = ~(layer3_outputs[3138]);
    assign layer4_outputs[3341] = ~(layer3_outputs[1379]) | (layer3_outputs[4307]);
    assign layer4_outputs[3342] = ~(layer3_outputs[3156]);
    assign layer4_outputs[3343] = ~(layer3_outputs[3275]) | (layer3_outputs[492]);
    assign layer4_outputs[3344] = ~(layer3_outputs[228]) | (layer3_outputs[2852]);
    assign layer4_outputs[3345] = ~((layer3_outputs[3256]) ^ (layer3_outputs[1771]));
    assign layer4_outputs[3346] = layer3_outputs[1542];
    assign layer4_outputs[3347] = ~(layer3_outputs[5041]) | (layer3_outputs[504]);
    assign layer4_outputs[3348] = layer3_outputs[4150];
    assign layer4_outputs[3349] = ~((layer3_outputs[2226]) & (layer3_outputs[2204]));
    assign layer4_outputs[3350] = ~((layer3_outputs[299]) | (layer3_outputs[2900]));
    assign layer4_outputs[3351] = ~(layer3_outputs[1505]);
    assign layer4_outputs[3352] = (layer3_outputs[3637]) & ~(layer3_outputs[2489]);
    assign layer4_outputs[3353] = (layer3_outputs[1585]) & ~(layer3_outputs[316]);
    assign layer4_outputs[3354] = layer3_outputs[4220];
    assign layer4_outputs[3355] = (layer3_outputs[6]) & (layer3_outputs[3468]);
    assign layer4_outputs[3356] = layer3_outputs[3386];
    assign layer4_outputs[3357] = (layer3_outputs[4856]) | (layer3_outputs[2524]);
    assign layer4_outputs[3358] = layer3_outputs[5113];
    assign layer4_outputs[3359] = (layer3_outputs[2045]) & ~(layer3_outputs[1225]);
    assign layer4_outputs[3360] = ~(layer3_outputs[5119]) | (layer3_outputs[1926]);
    assign layer4_outputs[3361] = layer3_outputs[4043];
    assign layer4_outputs[3362] = ~(layer3_outputs[4819]);
    assign layer4_outputs[3363] = ~(layer3_outputs[324]);
    assign layer4_outputs[3364] = ~(layer3_outputs[2280]);
    assign layer4_outputs[3365] = 1'b1;
    assign layer4_outputs[3366] = ~(layer3_outputs[1857]) | (layer3_outputs[3675]);
    assign layer4_outputs[3367] = ~(layer3_outputs[917]);
    assign layer4_outputs[3368] = ~(layer3_outputs[3132]);
    assign layer4_outputs[3369] = ~(layer3_outputs[408]);
    assign layer4_outputs[3370] = layer3_outputs[4009];
    assign layer4_outputs[3371] = layer3_outputs[2463];
    assign layer4_outputs[3372] = ~(layer3_outputs[2480]);
    assign layer4_outputs[3373] = ~(layer3_outputs[5043]);
    assign layer4_outputs[3374] = (layer3_outputs[4004]) & ~(layer3_outputs[2320]);
    assign layer4_outputs[3375] = ~(layer3_outputs[2654]);
    assign layer4_outputs[3376] = ~((layer3_outputs[2090]) ^ (layer3_outputs[3064]));
    assign layer4_outputs[3377] = 1'b0;
    assign layer4_outputs[3378] = 1'b1;
    assign layer4_outputs[3379] = ~(layer3_outputs[2847]);
    assign layer4_outputs[3380] = ~(layer3_outputs[1090]) | (layer3_outputs[4113]);
    assign layer4_outputs[3381] = layer3_outputs[1812];
    assign layer4_outputs[3382] = layer3_outputs[4779];
    assign layer4_outputs[3383] = (layer3_outputs[1240]) & ~(layer3_outputs[3090]);
    assign layer4_outputs[3384] = ~(layer3_outputs[2399]) | (layer3_outputs[1625]);
    assign layer4_outputs[3385] = ~(layer3_outputs[2384]);
    assign layer4_outputs[3386] = ~(layer3_outputs[3036]) | (layer3_outputs[1666]);
    assign layer4_outputs[3387] = (layer3_outputs[194]) & ~(layer3_outputs[3709]);
    assign layer4_outputs[3388] = 1'b0;
    assign layer4_outputs[3389] = layer3_outputs[2842];
    assign layer4_outputs[3390] = ~(layer3_outputs[4783]) | (layer3_outputs[1175]);
    assign layer4_outputs[3391] = (layer3_outputs[2066]) & ~(layer3_outputs[1067]);
    assign layer4_outputs[3392] = ~(layer3_outputs[4740]);
    assign layer4_outputs[3393] = layer3_outputs[3131];
    assign layer4_outputs[3394] = ~(layer3_outputs[1082]);
    assign layer4_outputs[3395] = 1'b1;
    assign layer4_outputs[3396] = ~(layer3_outputs[4669]) | (layer3_outputs[788]);
    assign layer4_outputs[3397] = ~(layer3_outputs[886]) | (layer3_outputs[4932]);
    assign layer4_outputs[3398] = layer3_outputs[4450];
    assign layer4_outputs[3399] = (layer3_outputs[2353]) ^ (layer3_outputs[278]);
    assign layer4_outputs[3400] = (layer3_outputs[1255]) | (layer3_outputs[1624]);
    assign layer4_outputs[3401] = layer3_outputs[4691];
    assign layer4_outputs[3402] = ~((layer3_outputs[146]) & (layer3_outputs[0]));
    assign layer4_outputs[3403] = layer3_outputs[1990];
    assign layer4_outputs[3404] = ~(layer3_outputs[1668]) | (layer3_outputs[1405]);
    assign layer4_outputs[3405] = layer3_outputs[704];
    assign layer4_outputs[3406] = layer3_outputs[1180];
    assign layer4_outputs[3407] = ~((layer3_outputs[4906]) & (layer3_outputs[4139]));
    assign layer4_outputs[3408] = ~(layer3_outputs[1655]);
    assign layer4_outputs[3409] = ~(layer3_outputs[1991]) | (layer3_outputs[2720]);
    assign layer4_outputs[3410] = (layer3_outputs[3259]) & ~(layer3_outputs[759]);
    assign layer4_outputs[3411] = ~(layer3_outputs[3862]) | (layer3_outputs[39]);
    assign layer4_outputs[3412] = ~((layer3_outputs[509]) | (layer3_outputs[390]));
    assign layer4_outputs[3413] = (layer3_outputs[4241]) ^ (layer3_outputs[4035]);
    assign layer4_outputs[3414] = ~((layer3_outputs[2933]) & (layer3_outputs[4036]));
    assign layer4_outputs[3415] = layer3_outputs[3370];
    assign layer4_outputs[3416] = (layer3_outputs[2154]) & ~(layer3_outputs[3518]);
    assign layer4_outputs[3417] = ~(layer3_outputs[2573]);
    assign layer4_outputs[3418] = ~(layer3_outputs[195]);
    assign layer4_outputs[3419] = (layer3_outputs[1375]) & (layer3_outputs[4726]);
    assign layer4_outputs[3420] = ~(layer3_outputs[294]) | (layer3_outputs[2622]);
    assign layer4_outputs[3421] = ~(layer3_outputs[1138]);
    assign layer4_outputs[3422] = (layer3_outputs[4836]) & ~(layer3_outputs[51]);
    assign layer4_outputs[3423] = ~(layer3_outputs[3237]) | (layer3_outputs[3253]);
    assign layer4_outputs[3424] = ~(layer3_outputs[1629]) | (layer3_outputs[172]);
    assign layer4_outputs[3425] = 1'b0;
    assign layer4_outputs[3426] = layer3_outputs[4252];
    assign layer4_outputs[3427] = (layer3_outputs[4086]) | (layer3_outputs[2611]);
    assign layer4_outputs[3428] = layer3_outputs[4467];
    assign layer4_outputs[3429] = layer3_outputs[2942];
    assign layer4_outputs[3430] = layer3_outputs[270];
    assign layer4_outputs[3431] = layer3_outputs[3425];
    assign layer4_outputs[3432] = ~(layer3_outputs[2504]);
    assign layer4_outputs[3433] = 1'b0;
    assign layer4_outputs[3434] = ~((layer3_outputs[1542]) ^ (layer3_outputs[1808]));
    assign layer4_outputs[3435] = layer3_outputs[3713];
    assign layer4_outputs[3436] = ~(layer3_outputs[3958]);
    assign layer4_outputs[3437] = ~((layer3_outputs[3914]) & (layer3_outputs[4849]));
    assign layer4_outputs[3438] = (layer3_outputs[4744]) & (layer3_outputs[1892]);
    assign layer4_outputs[3439] = ~((layer3_outputs[291]) ^ (layer3_outputs[2718]));
    assign layer4_outputs[3440] = ~(layer3_outputs[904]);
    assign layer4_outputs[3441] = ~(layer3_outputs[4987]);
    assign layer4_outputs[3442] = (layer3_outputs[3868]) & ~(layer3_outputs[2424]);
    assign layer4_outputs[3443] = ~(layer3_outputs[3966]);
    assign layer4_outputs[3444] = ~(layer3_outputs[4695]) | (layer3_outputs[3680]);
    assign layer4_outputs[3445] = ~(layer3_outputs[1458]) | (layer3_outputs[3828]);
    assign layer4_outputs[3446] = layer3_outputs[958];
    assign layer4_outputs[3447] = ~(layer3_outputs[2837]);
    assign layer4_outputs[3448] = ~((layer3_outputs[3346]) ^ (layer3_outputs[3564]));
    assign layer4_outputs[3449] = layer3_outputs[3699];
    assign layer4_outputs[3450] = ~((layer3_outputs[2979]) ^ (layer3_outputs[3326]));
    assign layer4_outputs[3451] = layer3_outputs[948];
    assign layer4_outputs[3452] = ~(layer3_outputs[3830]) | (layer3_outputs[526]);
    assign layer4_outputs[3453] = (layer3_outputs[3927]) & ~(layer3_outputs[2883]);
    assign layer4_outputs[3454] = (layer3_outputs[2574]) & (layer3_outputs[4680]);
    assign layer4_outputs[3455] = ~((layer3_outputs[2372]) | (layer3_outputs[3421]));
    assign layer4_outputs[3456] = (layer3_outputs[1551]) & ~(layer3_outputs[4234]);
    assign layer4_outputs[3457] = ~((layer3_outputs[4219]) & (layer3_outputs[2]));
    assign layer4_outputs[3458] = layer3_outputs[4587];
    assign layer4_outputs[3459] = 1'b1;
    assign layer4_outputs[3460] = (layer3_outputs[3951]) | (layer3_outputs[1951]);
    assign layer4_outputs[3461] = ~(layer3_outputs[2469]) | (layer3_outputs[1668]);
    assign layer4_outputs[3462] = ~(layer3_outputs[2054]) | (layer3_outputs[2135]);
    assign layer4_outputs[3463] = (layer3_outputs[2651]) & ~(layer3_outputs[2414]);
    assign layer4_outputs[3464] = ~((layer3_outputs[971]) | (layer3_outputs[3215]));
    assign layer4_outputs[3465] = layer3_outputs[3035];
    assign layer4_outputs[3466] = ~((layer3_outputs[3163]) | (layer3_outputs[4395]));
    assign layer4_outputs[3467] = 1'b0;
    assign layer4_outputs[3468] = layer3_outputs[3105];
    assign layer4_outputs[3469] = ~((layer3_outputs[4867]) | (layer3_outputs[1773]));
    assign layer4_outputs[3470] = 1'b1;
    assign layer4_outputs[3471] = (layer3_outputs[97]) ^ (layer3_outputs[3419]);
    assign layer4_outputs[3472] = ~(layer3_outputs[2636]) | (layer3_outputs[1318]);
    assign layer4_outputs[3473] = ~((layer3_outputs[4639]) | (layer3_outputs[2279]));
    assign layer4_outputs[3474] = ~(layer3_outputs[104]);
    assign layer4_outputs[3475] = ~((layer3_outputs[1887]) ^ (layer3_outputs[4261]));
    assign layer4_outputs[3476] = ~((layer3_outputs[206]) & (layer3_outputs[3800]));
    assign layer4_outputs[3477] = ~(layer3_outputs[2408]);
    assign layer4_outputs[3478] = layer3_outputs[3528];
    assign layer4_outputs[3479] = ~(layer3_outputs[3930]);
    assign layer4_outputs[3480] = ~(layer3_outputs[1287]);
    assign layer4_outputs[3481] = (layer3_outputs[4418]) & ~(layer3_outputs[114]);
    assign layer4_outputs[3482] = layer3_outputs[3883];
    assign layer4_outputs[3483] = ~((layer3_outputs[1966]) ^ (layer3_outputs[2357]));
    assign layer4_outputs[3484] = ~(layer3_outputs[4204]) | (layer3_outputs[551]);
    assign layer4_outputs[3485] = ~((layer3_outputs[2533]) | (layer3_outputs[735]));
    assign layer4_outputs[3486] = (layer3_outputs[2023]) & (layer3_outputs[3992]);
    assign layer4_outputs[3487] = ~((layer3_outputs[4339]) | (layer3_outputs[3094]));
    assign layer4_outputs[3488] = ~(layer3_outputs[2466]) | (layer3_outputs[3484]);
    assign layer4_outputs[3489] = layer3_outputs[2081];
    assign layer4_outputs[3490] = ~(layer3_outputs[2975]);
    assign layer4_outputs[3491] = (layer3_outputs[1033]) & (layer3_outputs[1969]);
    assign layer4_outputs[3492] = 1'b0;
    assign layer4_outputs[3493] = (layer3_outputs[4264]) & ~(layer3_outputs[4231]);
    assign layer4_outputs[3494] = ~(layer3_outputs[2807]);
    assign layer4_outputs[3495] = (layer3_outputs[626]) & (layer3_outputs[1407]);
    assign layer4_outputs[3496] = (layer3_outputs[3097]) & (layer3_outputs[2256]);
    assign layer4_outputs[3497] = ~(layer3_outputs[1986]);
    assign layer4_outputs[3498] = layer3_outputs[1032];
    assign layer4_outputs[3499] = ~((layer3_outputs[2834]) | (layer3_outputs[1632]));
    assign layer4_outputs[3500] = ~((layer3_outputs[4]) | (layer3_outputs[2027]));
    assign layer4_outputs[3501] = layer3_outputs[4422];
    assign layer4_outputs[3502] = layer3_outputs[3714];
    assign layer4_outputs[3503] = ~((layer3_outputs[3707]) ^ (layer3_outputs[2427]));
    assign layer4_outputs[3504] = ~(layer3_outputs[4103]) | (layer3_outputs[1862]);
    assign layer4_outputs[3505] = layer3_outputs[2645];
    assign layer4_outputs[3506] = ~(layer3_outputs[143]);
    assign layer4_outputs[3507] = (layer3_outputs[776]) | (layer3_outputs[3622]);
    assign layer4_outputs[3508] = layer3_outputs[3504];
    assign layer4_outputs[3509] = ~((layer3_outputs[142]) ^ (layer3_outputs[4119]));
    assign layer4_outputs[3510] = layer3_outputs[121];
    assign layer4_outputs[3511] = layer3_outputs[4607];
    assign layer4_outputs[3512] = (layer3_outputs[3503]) | (layer3_outputs[3203]);
    assign layer4_outputs[3513] = ~(layer3_outputs[658]);
    assign layer4_outputs[3514] = (layer3_outputs[3842]) & ~(layer3_outputs[820]);
    assign layer4_outputs[3515] = ~(layer3_outputs[4688]);
    assign layer4_outputs[3516] = ~(layer3_outputs[2526]);
    assign layer4_outputs[3517] = layer3_outputs[1739];
    assign layer4_outputs[3518] = (layer3_outputs[1237]) ^ (layer3_outputs[1805]);
    assign layer4_outputs[3519] = ~((layer3_outputs[2637]) | (layer3_outputs[3700]));
    assign layer4_outputs[3520] = ~((layer3_outputs[2833]) | (layer3_outputs[3659]));
    assign layer4_outputs[3521] = layer3_outputs[1047];
    assign layer4_outputs[3522] = (layer3_outputs[1695]) & ~(layer3_outputs[2846]);
    assign layer4_outputs[3523] = ~(layer3_outputs[827]) | (layer3_outputs[1049]);
    assign layer4_outputs[3524] = ~(layer3_outputs[3245]) | (layer3_outputs[3655]);
    assign layer4_outputs[3525] = (layer3_outputs[3666]) & (layer3_outputs[2886]);
    assign layer4_outputs[3526] = layer3_outputs[2684];
    assign layer4_outputs[3527] = (layer3_outputs[2220]) & (layer3_outputs[3758]);
    assign layer4_outputs[3528] = 1'b0;
    assign layer4_outputs[3529] = ~(layer3_outputs[1899]);
    assign layer4_outputs[3530] = layer3_outputs[4096];
    assign layer4_outputs[3531] = layer3_outputs[42];
    assign layer4_outputs[3532] = layer3_outputs[1856];
    assign layer4_outputs[3533] = layer3_outputs[2439];
    assign layer4_outputs[3534] = 1'b0;
    assign layer4_outputs[3535] = (layer3_outputs[1036]) ^ (layer3_outputs[1775]);
    assign layer4_outputs[3536] = ~((layer3_outputs[4029]) & (layer3_outputs[1985]));
    assign layer4_outputs[3537] = ~(layer3_outputs[2960]);
    assign layer4_outputs[3538] = ~(layer3_outputs[4552]);
    assign layer4_outputs[3539] = ~(layer3_outputs[4874]);
    assign layer4_outputs[3540] = (layer3_outputs[1276]) & (layer3_outputs[1567]);
    assign layer4_outputs[3541] = (layer3_outputs[1351]) | (layer3_outputs[5117]);
    assign layer4_outputs[3542] = layer3_outputs[3106];
    assign layer4_outputs[3543] = ~(layer3_outputs[4725]);
    assign layer4_outputs[3544] = ~((layer3_outputs[3221]) | (layer3_outputs[2132]));
    assign layer4_outputs[3545] = 1'b0;
    assign layer4_outputs[3546] = ~(layer3_outputs[438]);
    assign layer4_outputs[3547] = ~(layer3_outputs[3503]);
    assign layer4_outputs[3548] = layer3_outputs[4402];
    assign layer4_outputs[3549] = layer3_outputs[3876];
    assign layer4_outputs[3550] = ~(layer3_outputs[2266]);
    assign layer4_outputs[3551] = ~(layer3_outputs[4004]);
    assign layer4_outputs[3552] = (layer3_outputs[4235]) & (layer3_outputs[1029]);
    assign layer4_outputs[3553] = (layer3_outputs[2162]) & (layer3_outputs[138]);
    assign layer4_outputs[3554] = ~(layer3_outputs[4270]);
    assign layer4_outputs[3555] = ~(layer3_outputs[2443]);
    assign layer4_outputs[3556] = ~(layer3_outputs[1934]);
    assign layer4_outputs[3557] = ~((layer3_outputs[2376]) | (layer3_outputs[367]));
    assign layer4_outputs[3558] = ~(layer3_outputs[21]);
    assign layer4_outputs[3559] = layer3_outputs[2395];
    assign layer4_outputs[3560] = ~(layer3_outputs[4114]);
    assign layer4_outputs[3561] = layer3_outputs[1555];
    assign layer4_outputs[3562] = ~(layer3_outputs[5067]);
    assign layer4_outputs[3563] = ~(layer3_outputs[851]);
    assign layer4_outputs[3564] = ~(layer3_outputs[1827]) | (layer3_outputs[4562]);
    assign layer4_outputs[3565] = ~(layer3_outputs[379]);
    assign layer4_outputs[3566] = ~((layer3_outputs[3052]) | (layer3_outputs[2854]));
    assign layer4_outputs[3567] = (layer3_outputs[2394]) ^ (layer3_outputs[345]);
    assign layer4_outputs[3568] = (layer3_outputs[118]) & (layer3_outputs[3349]);
    assign layer4_outputs[3569] = ~(layer3_outputs[4825]) | (layer3_outputs[1863]);
    assign layer4_outputs[3570] = ~(layer3_outputs[2314]);
    assign layer4_outputs[3571] = ~(layer3_outputs[281]);
    assign layer4_outputs[3572] = ~(layer3_outputs[604]) | (layer3_outputs[87]);
    assign layer4_outputs[3573] = ~(layer3_outputs[939]) | (layer3_outputs[3271]);
    assign layer4_outputs[3574] = (layer3_outputs[777]) ^ (layer3_outputs[3119]);
    assign layer4_outputs[3575] = ~(layer3_outputs[5027]);
    assign layer4_outputs[3576] = layer3_outputs[2791];
    assign layer4_outputs[3577] = ~(layer3_outputs[2173]) | (layer3_outputs[4015]);
    assign layer4_outputs[3578] = (layer3_outputs[3781]) & (layer3_outputs[3226]);
    assign layer4_outputs[3579] = layer3_outputs[4791];
    assign layer4_outputs[3580] = ~((layer3_outputs[3144]) & (layer3_outputs[3155]));
    assign layer4_outputs[3581] = layer3_outputs[1349];
    assign layer4_outputs[3582] = layer3_outputs[1307];
    assign layer4_outputs[3583] = (layer3_outputs[501]) & (layer3_outputs[3487]);
    assign layer4_outputs[3584] = ~(layer3_outputs[4491]);
    assign layer4_outputs[3585] = ~((layer3_outputs[2707]) ^ (layer3_outputs[227]));
    assign layer4_outputs[3586] = ~((layer3_outputs[327]) & (layer3_outputs[4063]));
    assign layer4_outputs[3587] = (layer3_outputs[2605]) & ~(layer3_outputs[1030]);
    assign layer4_outputs[3588] = ~(layer3_outputs[4942]);
    assign layer4_outputs[3589] = (layer3_outputs[3583]) & ~(layer3_outputs[806]);
    assign layer4_outputs[3590] = (layer3_outputs[4724]) & ~(layer3_outputs[1566]);
    assign layer4_outputs[3591] = layer3_outputs[1786];
    assign layer4_outputs[3592] = layer3_outputs[4127];
    assign layer4_outputs[3593] = ~((layer3_outputs[3219]) & (layer3_outputs[2905]));
    assign layer4_outputs[3594] = ~((layer3_outputs[1043]) & (layer3_outputs[2040]));
    assign layer4_outputs[3595] = 1'b1;
    assign layer4_outputs[3596] = (layer3_outputs[5032]) & (layer3_outputs[4162]);
    assign layer4_outputs[3597] = layer3_outputs[4178];
    assign layer4_outputs[3598] = layer3_outputs[1767];
    assign layer4_outputs[3599] = layer3_outputs[4543];
    assign layer4_outputs[3600] = ~((layer3_outputs[2622]) & (layer3_outputs[1081]));
    assign layer4_outputs[3601] = layer3_outputs[891];
    assign layer4_outputs[3602] = 1'b1;
    assign layer4_outputs[3603] = ~(layer3_outputs[4153]);
    assign layer4_outputs[3604] = (layer3_outputs[4313]) & ~(layer3_outputs[3859]);
    assign layer4_outputs[3605] = layer3_outputs[494];
    assign layer4_outputs[3606] = layer3_outputs[1057];
    assign layer4_outputs[3607] = ~(layer3_outputs[3577]);
    assign layer4_outputs[3608] = ~((layer3_outputs[2595]) | (layer3_outputs[767]));
    assign layer4_outputs[3609] = ~((layer3_outputs[3494]) ^ (layer3_outputs[22]));
    assign layer4_outputs[3610] = ~(layer3_outputs[4305]);
    assign layer4_outputs[3611] = ~(layer3_outputs[1710]);
    assign layer4_outputs[3612] = (layer3_outputs[1018]) & ~(layer3_outputs[3940]);
    assign layer4_outputs[3613] = ~(layer3_outputs[1150]) | (layer3_outputs[3045]);
    assign layer4_outputs[3614] = ~(layer3_outputs[2407]);
    assign layer4_outputs[3615] = layer3_outputs[884];
    assign layer4_outputs[3616] = ~(layer3_outputs[4277]);
    assign layer4_outputs[3617] = ~(layer3_outputs[665]) | (layer3_outputs[885]);
    assign layer4_outputs[3618] = (layer3_outputs[4445]) & ~(layer3_outputs[4337]);
    assign layer4_outputs[3619] = ~(layer3_outputs[3845]);
    assign layer4_outputs[3620] = 1'b1;
    assign layer4_outputs[3621] = ~(layer3_outputs[2703]);
    assign layer4_outputs[3622] = 1'b0;
    assign layer4_outputs[3623] = (layer3_outputs[1780]) & ~(layer3_outputs[3340]);
    assign layer4_outputs[3624] = (layer3_outputs[4391]) & ~(layer3_outputs[4016]);
    assign layer4_outputs[3625] = ~(layer3_outputs[3517]) | (layer3_outputs[3800]);
    assign layer4_outputs[3626] = ~((layer3_outputs[3083]) & (layer3_outputs[1943]));
    assign layer4_outputs[3627] = layer3_outputs[2258];
    assign layer4_outputs[3628] = layer3_outputs[3312];
    assign layer4_outputs[3629] = (layer3_outputs[2429]) & ~(layer3_outputs[1675]);
    assign layer4_outputs[3630] = ~((layer3_outputs[4591]) | (layer3_outputs[725]));
    assign layer4_outputs[3631] = (layer3_outputs[2673]) & ~(layer3_outputs[797]);
    assign layer4_outputs[3632] = (layer3_outputs[4760]) ^ (layer3_outputs[487]);
    assign layer4_outputs[3633] = ~(layer3_outputs[981]) | (layer3_outputs[2139]);
    assign layer4_outputs[3634] = layer3_outputs[2303];
    assign layer4_outputs[3635] = ~(layer3_outputs[2289]) | (layer3_outputs[650]);
    assign layer4_outputs[3636] = layer3_outputs[598];
    assign layer4_outputs[3637] = layer3_outputs[4939];
    assign layer4_outputs[3638] = ~(layer3_outputs[3418]);
    assign layer4_outputs[3639] = ~(layer3_outputs[3455]);
    assign layer4_outputs[3640] = ~(layer3_outputs[957]) | (layer3_outputs[1681]);
    assign layer4_outputs[3641] = ~((layer3_outputs[4830]) & (layer3_outputs[4593]));
    assign layer4_outputs[3642] = ~(layer3_outputs[3173]);
    assign layer4_outputs[3643] = 1'b1;
    assign layer4_outputs[3644] = 1'b0;
    assign layer4_outputs[3645] = (layer3_outputs[2882]) | (layer3_outputs[3488]);
    assign layer4_outputs[3646] = layer3_outputs[1058];
    assign layer4_outputs[3647] = layer3_outputs[3252];
    assign layer4_outputs[3648] = ~(layer3_outputs[3167]);
    assign layer4_outputs[3649] = layer3_outputs[2918];
    assign layer4_outputs[3650] = ~(layer3_outputs[357]);
    assign layer4_outputs[3651] = (layer3_outputs[4420]) & ~(layer3_outputs[4776]);
    assign layer4_outputs[3652] = (layer3_outputs[2318]) & (layer3_outputs[1541]);
    assign layer4_outputs[3653] = (layer3_outputs[2329]) & ~(layer3_outputs[1810]);
    assign layer4_outputs[3654] = ~(layer3_outputs[224]);
    assign layer4_outputs[3655] = ~((layer3_outputs[51]) & (layer3_outputs[4746]));
    assign layer4_outputs[3656] = (layer3_outputs[1957]) | (layer3_outputs[2295]);
    assign layer4_outputs[3657] = (layer3_outputs[1236]) & ~(layer3_outputs[3943]);
    assign layer4_outputs[3658] = layer3_outputs[1774];
    assign layer4_outputs[3659] = (layer3_outputs[539]) | (layer3_outputs[2387]);
    assign layer4_outputs[3660] = 1'b0;
    assign layer4_outputs[3661] = ~(layer3_outputs[1282]) | (layer3_outputs[237]);
    assign layer4_outputs[3662] = ~(layer3_outputs[4979]);
    assign layer4_outputs[3663] = ~(layer3_outputs[13]);
    assign layer4_outputs[3664] = ~(layer3_outputs[174]);
    assign layer4_outputs[3665] = ~(layer3_outputs[3767]);
    assign layer4_outputs[3666] = layer3_outputs[3716];
    assign layer4_outputs[3667] = ~(layer3_outputs[832]);
    assign layer4_outputs[3668] = ~((layer3_outputs[4067]) & (layer3_outputs[166]));
    assign layer4_outputs[3669] = 1'b1;
    assign layer4_outputs[3670] = 1'b1;
    assign layer4_outputs[3671] = ~(layer3_outputs[2992]);
    assign layer4_outputs[3672] = ~(layer3_outputs[3262]);
    assign layer4_outputs[3673] = 1'b1;
    assign layer4_outputs[3674] = layer3_outputs[1913];
    assign layer4_outputs[3675] = (layer3_outputs[2900]) & ~(layer3_outputs[719]);
    assign layer4_outputs[3676] = ~((layer3_outputs[4555]) | (layer3_outputs[1879]));
    assign layer4_outputs[3677] = (layer3_outputs[235]) & (layer3_outputs[4021]);
    assign layer4_outputs[3678] = ~(layer3_outputs[4704]) | (layer3_outputs[2150]);
    assign layer4_outputs[3679] = layer3_outputs[3048];
    assign layer4_outputs[3680] = ~(layer3_outputs[861]);
    assign layer4_outputs[3681] = ~(layer3_outputs[1449]) | (layer3_outputs[2665]);
    assign layer4_outputs[3682] = layer3_outputs[4546];
    assign layer4_outputs[3683] = layer3_outputs[1726];
    assign layer4_outputs[3684] = 1'b1;
    assign layer4_outputs[3685] = 1'b1;
    assign layer4_outputs[3686] = ~(layer3_outputs[1066]);
    assign layer4_outputs[3687] = ~((layer3_outputs[2038]) & (layer3_outputs[1062]));
    assign layer4_outputs[3688] = (layer3_outputs[1860]) | (layer3_outputs[500]);
    assign layer4_outputs[3689] = 1'b1;
    assign layer4_outputs[3690] = ~(layer3_outputs[3986]);
    assign layer4_outputs[3691] = ~(layer3_outputs[4618]) | (layer3_outputs[170]);
    assign layer4_outputs[3692] = (layer3_outputs[2238]) & ~(layer3_outputs[2238]);
    assign layer4_outputs[3693] = 1'b0;
    assign layer4_outputs[3694] = layer3_outputs[1703];
    assign layer4_outputs[3695] = layer3_outputs[1202];
    assign layer4_outputs[3696] = ~(layer3_outputs[4180]);
    assign layer4_outputs[3697] = ~(layer3_outputs[1399]);
    assign layer4_outputs[3698] = layer3_outputs[1025];
    assign layer4_outputs[3699] = (layer3_outputs[1034]) | (layer3_outputs[3163]);
    assign layer4_outputs[3700] = ~((layer3_outputs[1174]) & (layer3_outputs[4803]));
    assign layer4_outputs[3701] = ~((layer3_outputs[2794]) | (layer3_outputs[1533]));
    assign layer4_outputs[3702] = ~(layer3_outputs[4728]);
    assign layer4_outputs[3703] = layer3_outputs[1899];
    assign layer4_outputs[3704] = ~(layer3_outputs[2447]);
    assign layer4_outputs[3705] = ~(layer3_outputs[4793]);
    assign layer4_outputs[3706] = 1'b0;
    assign layer4_outputs[3707] = layer3_outputs[2577];
    assign layer4_outputs[3708] = ~(layer3_outputs[2323]) | (layer3_outputs[4699]);
    assign layer4_outputs[3709] = 1'b0;
    assign layer4_outputs[3710] = ~(layer3_outputs[74]);
    assign layer4_outputs[3711] = layer3_outputs[3050];
    assign layer4_outputs[3712] = ~(layer3_outputs[1648]) | (layer3_outputs[150]);
    assign layer4_outputs[3713] = layer3_outputs[2867];
    assign layer4_outputs[3714] = ~(layer3_outputs[1786]);
    assign layer4_outputs[3715] = ~(layer3_outputs[636]);
    assign layer4_outputs[3716] = layer3_outputs[2571];
    assign layer4_outputs[3717] = ~(layer3_outputs[1276]);
    assign layer4_outputs[3718] = (layer3_outputs[3872]) & (layer3_outputs[994]);
    assign layer4_outputs[3719] = ~((layer3_outputs[2680]) & (layer3_outputs[3498]));
    assign layer4_outputs[3720] = ~(layer3_outputs[2755]) | (layer3_outputs[4482]);
    assign layer4_outputs[3721] = (layer3_outputs[3201]) ^ (layer3_outputs[5047]);
    assign layer4_outputs[3722] = layer3_outputs[1187];
    assign layer4_outputs[3723] = layer3_outputs[912];
    assign layer4_outputs[3724] = ~(layer3_outputs[2177]);
    assign layer4_outputs[3725] = (layer3_outputs[941]) & ~(layer3_outputs[85]);
    assign layer4_outputs[3726] = ~(layer3_outputs[2405]);
    assign layer4_outputs[3727] = ~(layer3_outputs[3342]);
    assign layer4_outputs[3728] = ~((layer3_outputs[4685]) & (layer3_outputs[2211]));
    assign layer4_outputs[3729] = ~(layer3_outputs[2521]);
    assign layer4_outputs[3730] = layer3_outputs[907];
    assign layer4_outputs[3731] = 1'b1;
    assign layer4_outputs[3732] = ~((layer3_outputs[2281]) ^ (layer3_outputs[3442]));
    assign layer4_outputs[3733] = (layer3_outputs[1464]) & ~(layer3_outputs[4972]);
    assign layer4_outputs[3734] = (layer3_outputs[381]) & (layer3_outputs[1631]);
    assign layer4_outputs[3735] = ~((layer3_outputs[3930]) ^ (layer3_outputs[3392]));
    assign layer4_outputs[3736] = ~((layer3_outputs[2505]) ^ (layer3_outputs[3803]));
    assign layer4_outputs[3737] = ~(layer3_outputs[1650]);
    assign layer4_outputs[3738] = (layer3_outputs[4503]) ^ (layer3_outputs[2723]);
    assign layer4_outputs[3739] = ~(layer3_outputs[2325]);
    assign layer4_outputs[3740] = ~(layer3_outputs[585]);
    assign layer4_outputs[3741] = ~((layer3_outputs[2401]) & (layer3_outputs[3865]));
    assign layer4_outputs[3742] = layer3_outputs[602];
    assign layer4_outputs[3743] = ~((layer3_outputs[1432]) & (layer3_outputs[674]));
    assign layer4_outputs[3744] = ~((layer3_outputs[1908]) & (layer3_outputs[3735]));
    assign layer4_outputs[3745] = ~(layer3_outputs[3544]);
    assign layer4_outputs[3746] = ~(layer3_outputs[4538]);
    assign layer4_outputs[3747] = (layer3_outputs[4145]) & ~(layer3_outputs[2277]);
    assign layer4_outputs[3748] = layer3_outputs[4633];
    assign layer4_outputs[3749] = ~(layer3_outputs[4016]) | (layer3_outputs[5094]);
    assign layer4_outputs[3750] = ~(layer3_outputs[2297]);
    assign layer4_outputs[3751] = ~(layer3_outputs[4286]);
    assign layer4_outputs[3752] = (layer3_outputs[4948]) & ~(layer3_outputs[1811]);
    assign layer4_outputs[3753] = ~(layer3_outputs[2381]) | (layer3_outputs[483]);
    assign layer4_outputs[3754] = ~(layer3_outputs[4299]);
    assign layer4_outputs[3755] = (layer3_outputs[2022]) & (layer3_outputs[3704]);
    assign layer4_outputs[3756] = (layer3_outputs[2927]) & ~(layer3_outputs[3814]);
    assign layer4_outputs[3757] = (layer3_outputs[1780]) & ~(layer3_outputs[3335]);
    assign layer4_outputs[3758] = ~((layer3_outputs[1304]) ^ (layer3_outputs[1143]));
    assign layer4_outputs[3759] = ~(layer3_outputs[3479]);
    assign layer4_outputs[3760] = ~(layer3_outputs[925]);
    assign layer4_outputs[3761] = layer3_outputs[2695];
    assign layer4_outputs[3762] = ~(layer3_outputs[4858]) | (layer3_outputs[1347]);
    assign layer4_outputs[3763] = layer3_outputs[3391];
    assign layer4_outputs[3764] = (layer3_outputs[1973]) & ~(layer3_outputs[5084]);
    assign layer4_outputs[3765] = ~(layer3_outputs[5062]) | (layer3_outputs[4371]);
    assign layer4_outputs[3766] = ~(layer3_outputs[4412]);
    assign layer4_outputs[3767] = ~(layer3_outputs[3909]) | (layer3_outputs[4954]);
    assign layer4_outputs[3768] = ~(layer3_outputs[1411]) | (layer3_outputs[2229]);
    assign layer4_outputs[3769] = (layer3_outputs[4419]) | (layer3_outputs[640]);
    assign layer4_outputs[3770] = (layer3_outputs[5034]) & ~(layer3_outputs[457]);
    assign layer4_outputs[3771] = ~(layer3_outputs[2859]);
    assign layer4_outputs[3772] = ~(layer3_outputs[4417]);
    assign layer4_outputs[3773] = ~(layer3_outputs[4738]);
    assign layer4_outputs[3774] = layer3_outputs[2142];
    assign layer4_outputs[3775] = ~((layer3_outputs[3974]) | (layer3_outputs[2091]));
    assign layer4_outputs[3776] = layer3_outputs[4447];
    assign layer4_outputs[3777] = (layer3_outputs[3440]) & ~(layer3_outputs[209]);
    assign layer4_outputs[3778] = ~(layer3_outputs[1826]);
    assign layer4_outputs[3779] = ~(layer3_outputs[1680]) | (layer3_outputs[1177]);
    assign layer4_outputs[3780] = ~((layer3_outputs[615]) | (layer3_outputs[2273]));
    assign layer4_outputs[3781] = (layer3_outputs[1231]) & (layer3_outputs[1547]);
    assign layer4_outputs[3782] = ~(layer3_outputs[5064]);
    assign layer4_outputs[3783] = 1'b1;
    assign layer4_outputs[3784] = ~(layer3_outputs[4470]) | (layer3_outputs[1774]);
    assign layer4_outputs[3785] = layer3_outputs[2659];
    assign layer4_outputs[3786] = layer3_outputs[1261];
    assign layer4_outputs[3787] = ~(layer3_outputs[3227]) | (layer3_outputs[397]);
    assign layer4_outputs[3788] = ~((layer3_outputs[4276]) & (layer3_outputs[3395]));
    assign layer4_outputs[3789] = 1'b1;
    assign layer4_outputs[3790] = (layer3_outputs[3317]) & ~(layer3_outputs[2170]);
    assign layer4_outputs[3791] = ~((layer3_outputs[2578]) & (layer3_outputs[944]));
    assign layer4_outputs[3792] = ~(layer3_outputs[1832]);
    assign layer4_outputs[3793] = 1'b0;
    assign layer4_outputs[3794] = ~(layer3_outputs[5025]) | (layer3_outputs[4681]);
    assign layer4_outputs[3795] = (layer3_outputs[5081]) & ~(layer3_outputs[1848]);
    assign layer4_outputs[3796] = layer3_outputs[2734];
    assign layer4_outputs[3797] = (layer3_outputs[1799]) & ~(layer3_outputs[3973]);
    assign layer4_outputs[3798] = ~((layer3_outputs[619]) & (layer3_outputs[4092]));
    assign layer4_outputs[3799] = (layer3_outputs[2077]) | (layer3_outputs[2696]);
    assign layer4_outputs[3800] = (layer3_outputs[2403]) & ~(layer3_outputs[4945]);
    assign layer4_outputs[3801] = ~((layer3_outputs[4213]) & (layer3_outputs[1183]));
    assign layer4_outputs[3802] = (layer3_outputs[3258]) & ~(layer3_outputs[3884]);
    assign layer4_outputs[3803] = (layer3_outputs[3741]) & ~(layer3_outputs[2881]);
    assign layer4_outputs[3804] = (layer3_outputs[497]) ^ (layer3_outputs[542]);
    assign layer4_outputs[3805] = (layer3_outputs[4147]) & ~(layer3_outputs[896]);
    assign layer4_outputs[3806] = ~(layer3_outputs[258]) | (layer3_outputs[870]);
    assign layer4_outputs[3807] = ~((layer3_outputs[2431]) & (layer3_outputs[1367]));
    assign layer4_outputs[3808] = (layer3_outputs[1924]) & (layer3_outputs[2495]);
    assign layer4_outputs[3809] = ~(layer3_outputs[352]) | (layer3_outputs[78]);
    assign layer4_outputs[3810] = 1'b1;
    assign layer4_outputs[3811] = layer3_outputs[1383];
    assign layer4_outputs[3812] = ~(layer3_outputs[3491]);
    assign layer4_outputs[3813] = 1'b1;
    assign layer4_outputs[3814] = ~(layer3_outputs[4806]);
    assign layer4_outputs[3815] = ~((layer3_outputs[1421]) & (layer3_outputs[2415]));
    assign layer4_outputs[3816] = ~((layer3_outputs[1588]) | (layer3_outputs[4375]));
    assign layer4_outputs[3817] = layer3_outputs[2597];
    assign layer4_outputs[3818] = ~(layer3_outputs[3590]) | (layer3_outputs[3702]);
    assign layer4_outputs[3819] = ~((layer3_outputs[4839]) | (layer3_outputs[3589]));
    assign layer4_outputs[3820] = 1'b0;
    assign layer4_outputs[3821] = ~((layer3_outputs[896]) | (layer3_outputs[2346]));
    assign layer4_outputs[3822] = ~(layer3_outputs[1977]) | (layer3_outputs[4379]);
    assign layer4_outputs[3823] = ~((layer3_outputs[4411]) & (layer3_outputs[1517]));
    assign layer4_outputs[3824] = layer3_outputs[5053];
    assign layer4_outputs[3825] = (layer3_outputs[5066]) & ~(layer3_outputs[4190]);
    assign layer4_outputs[3826] = 1'b0;
    assign layer4_outputs[3827] = ~(layer3_outputs[1782]);
    assign layer4_outputs[3828] = ~((layer3_outputs[3365]) ^ (layer3_outputs[3090]));
    assign layer4_outputs[3829] = ~((layer3_outputs[3330]) & (layer3_outputs[45]));
    assign layer4_outputs[3830] = layer3_outputs[1728];
    assign layer4_outputs[3831] = ~(layer3_outputs[269]);
    assign layer4_outputs[3832] = 1'b0;
    assign layer4_outputs[3833] = ~(layer3_outputs[431]);
    assign layer4_outputs[3834] = 1'b0;
    assign layer4_outputs[3835] = layer3_outputs[2278];
    assign layer4_outputs[3836] = 1'b1;
    assign layer4_outputs[3837] = ~((layer3_outputs[4736]) | (layer3_outputs[1695]));
    assign layer4_outputs[3838] = ~(layer3_outputs[1903]);
    assign layer4_outputs[3839] = (layer3_outputs[3791]) | (layer3_outputs[547]);
    assign layer4_outputs[3840] = 1'b1;
    assign layer4_outputs[3841] = ~(layer3_outputs[2782]);
    assign layer4_outputs[3842] = (layer3_outputs[2860]) ^ (layer3_outputs[774]);
    assign layer4_outputs[3843] = ~(layer3_outputs[1040]) | (layer3_outputs[2604]);
    assign layer4_outputs[3844] = (layer3_outputs[5033]) & ~(layer3_outputs[1242]);
    assign layer4_outputs[3845] = ~((layer3_outputs[3885]) | (layer3_outputs[4663]));
    assign layer4_outputs[3846] = layer3_outputs[3932];
    assign layer4_outputs[3847] = ~((layer3_outputs[1881]) & (layer3_outputs[1790]));
    assign layer4_outputs[3848] = ~(layer3_outputs[381]);
    assign layer4_outputs[3849] = ~(layer3_outputs[2023]);
    assign layer4_outputs[3850] = layer3_outputs[3490];
    assign layer4_outputs[3851] = ~((layer3_outputs[2006]) | (layer3_outputs[5053]));
    assign layer4_outputs[3852] = ~((layer3_outputs[472]) ^ (layer3_outputs[3865]));
    assign layer4_outputs[3853] = layer3_outputs[760];
    assign layer4_outputs[3854] = (layer3_outputs[1505]) & ~(layer3_outputs[2515]);
    assign layer4_outputs[3855] = (layer3_outputs[2976]) | (layer3_outputs[3563]);
    assign layer4_outputs[3856] = ~(layer3_outputs[479]) | (layer3_outputs[1546]);
    assign layer4_outputs[3857] = ~(layer3_outputs[4611]);
    assign layer4_outputs[3858] = layer3_outputs[1257];
    assign layer4_outputs[3859] = ~(layer3_outputs[153]);
    assign layer4_outputs[3860] = ~(layer3_outputs[3324]) | (layer3_outputs[4600]);
    assign layer4_outputs[3861] = layer3_outputs[924];
    assign layer4_outputs[3862] = ~(layer3_outputs[4763]);
    assign layer4_outputs[3863] = ~(layer3_outputs[422]);
    assign layer4_outputs[3864] = ~(layer3_outputs[3797]);
    assign layer4_outputs[3865] = ~(layer3_outputs[3035]) | (layer3_outputs[1508]);
    assign layer4_outputs[3866] = (layer3_outputs[3060]) & (layer3_outputs[3175]);
    assign layer4_outputs[3867] = ~(layer3_outputs[3890]);
    assign layer4_outputs[3868] = ~(layer3_outputs[440]) | (layer3_outputs[867]);
    assign layer4_outputs[3869] = layer3_outputs[1712];
    assign layer4_outputs[3870] = ~((layer3_outputs[3991]) ^ (layer3_outputs[4463]));
    assign layer4_outputs[3871] = 1'b0;
    assign layer4_outputs[3872] = ~((layer3_outputs[3784]) & (layer3_outputs[4904]));
    assign layer4_outputs[3873] = (layer3_outputs[1263]) & (layer3_outputs[1743]);
    assign layer4_outputs[3874] = ~(layer3_outputs[1697]) | (layer3_outputs[931]);
    assign layer4_outputs[3875] = (layer3_outputs[3684]) ^ (layer3_outputs[1482]);
    assign layer4_outputs[3876] = ~(layer3_outputs[4344]);
    assign layer4_outputs[3877] = ~((layer3_outputs[161]) | (layer3_outputs[1895]));
    assign layer4_outputs[3878] = (layer3_outputs[537]) | (layer3_outputs[4680]);
    assign layer4_outputs[3879] = 1'b0;
    assign layer4_outputs[3880] = ~(layer3_outputs[3725]);
    assign layer4_outputs[3881] = ~(layer3_outputs[3042]) | (layer3_outputs[4874]);
    assign layer4_outputs[3882] = ~(layer3_outputs[991]);
    assign layer4_outputs[3883] = (layer3_outputs[857]) & ~(layer3_outputs[4988]);
    assign layer4_outputs[3884] = (layer3_outputs[4136]) & ~(layer3_outputs[3389]);
    assign layer4_outputs[3885] = ~(layer3_outputs[4993]);
    assign layer4_outputs[3886] = (layer3_outputs[1502]) ^ (layer3_outputs[415]);
    assign layer4_outputs[3887] = layer3_outputs[4222];
    assign layer4_outputs[3888] = ~(layer3_outputs[824]);
    assign layer4_outputs[3889] = ~(layer3_outputs[4420]);
    assign layer4_outputs[3890] = layer3_outputs[218];
    assign layer4_outputs[3891] = ~(layer3_outputs[762]) | (layer3_outputs[3554]);
    assign layer4_outputs[3892] = (layer3_outputs[4957]) & ~(layer3_outputs[592]);
    assign layer4_outputs[3893] = layer3_outputs[1707];
    assign layer4_outputs[3894] = ~((layer3_outputs[4906]) & (layer3_outputs[3796]));
    assign layer4_outputs[3895] = (layer3_outputs[1759]) & ~(layer3_outputs[829]);
    assign layer4_outputs[3896] = ~((layer3_outputs[1037]) & (layer3_outputs[1689]));
    assign layer4_outputs[3897] = ~(layer3_outputs[2615]);
    assign layer4_outputs[3898] = (layer3_outputs[4985]) & (layer3_outputs[3882]);
    assign layer4_outputs[3899] = ~(layer3_outputs[3692]);
    assign layer4_outputs[3900] = ~(layer3_outputs[4393]);
    assign layer4_outputs[3901] = ~((layer3_outputs[4021]) | (layer3_outputs[4745]));
    assign layer4_outputs[3902] = layer3_outputs[1829];
    assign layer4_outputs[3903] = 1'b1;
    assign layer4_outputs[3904] = ~(layer3_outputs[1045]) | (layer3_outputs[3071]);
    assign layer4_outputs[3905] = ~(layer3_outputs[1994]);
    assign layer4_outputs[3906] = layer3_outputs[2762];
    assign layer4_outputs[3907] = ~((layer3_outputs[2274]) | (layer3_outputs[3588]));
    assign layer4_outputs[3908] = layer3_outputs[837];
    assign layer4_outputs[3909] = 1'b1;
    assign layer4_outputs[3910] = layer3_outputs[2408];
    assign layer4_outputs[3911] = (layer3_outputs[423]) & ~(layer3_outputs[405]);
    assign layer4_outputs[3912] = (layer3_outputs[1972]) | (layer3_outputs[3513]);
    assign layer4_outputs[3913] = ~(layer3_outputs[3814]);
    assign layer4_outputs[3914] = layer3_outputs[935];
    assign layer4_outputs[3915] = (layer3_outputs[3243]) & ~(layer3_outputs[2088]);
    assign layer4_outputs[3916] = ~(layer3_outputs[3711]);
    assign layer4_outputs[3917] = (layer3_outputs[4307]) & ~(layer3_outputs[2868]);
    assign layer4_outputs[3918] = (layer3_outputs[3369]) & ~(layer3_outputs[4817]);
    assign layer4_outputs[3919] = (layer3_outputs[1156]) & ~(layer3_outputs[3001]);
    assign layer4_outputs[3920] = (layer3_outputs[2350]) & ~(layer3_outputs[758]);
    assign layer4_outputs[3921] = (layer3_outputs[707]) | (layer3_outputs[2301]);
    assign layer4_outputs[3922] = ~((layer3_outputs[4967]) & (layer3_outputs[3282]));
    assign layer4_outputs[3923] = layer3_outputs[3356];
    assign layer4_outputs[3924] = layer3_outputs[1392];
    assign layer4_outputs[3925] = ~((layer3_outputs[4786]) | (layer3_outputs[2925]));
    assign layer4_outputs[3926] = 1'b1;
    assign layer4_outputs[3927] = ~(layer3_outputs[3340]);
    assign layer4_outputs[3928] = ~(layer3_outputs[607]) | (layer3_outputs[167]);
    assign layer4_outputs[3929] = ~((layer3_outputs[105]) | (layer3_outputs[2056]));
    assign layer4_outputs[3930] = 1'b1;
    assign layer4_outputs[3931] = ~(layer3_outputs[3728]) | (layer3_outputs[685]);
    assign layer4_outputs[3932] = (layer3_outputs[4653]) & ~(layer3_outputs[2216]);
    assign layer4_outputs[3933] = ~(layer3_outputs[1213]);
    assign layer4_outputs[3934] = (layer3_outputs[4775]) & ~(layer3_outputs[1557]);
    assign layer4_outputs[3935] = ~(layer3_outputs[1831]);
    assign layer4_outputs[3936] = layer3_outputs[682];
    assign layer4_outputs[3937] = (layer3_outputs[3282]) | (layer3_outputs[4301]);
    assign layer4_outputs[3938] = layer3_outputs[263];
    assign layer4_outputs[3939] = ~(layer3_outputs[980]);
    assign layer4_outputs[3940] = ~(layer3_outputs[5050]);
    assign layer4_outputs[3941] = layer3_outputs[901];
    assign layer4_outputs[3942] = ~(layer3_outputs[811]);
    assign layer4_outputs[3943] = layer3_outputs[803];
    assign layer4_outputs[3944] = ~((layer3_outputs[1641]) & (layer3_outputs[2267]));
    assign layer4_outputs[3945] = ~(layer3_outputs[717]) | (layer3_outputs[1585]);
    assign layer4_outputs[3946] = ~((layer3_outputs[845]) & (layer3_outputs[4208]));
    assign layer4_outputs[3947] = ~((layer3_outputs[1215]) & (layer3_outputs[4188]));
    assign layer4_outputs[3948] = ~((layer3_outputs[4573]) | (layer3_outputs[2625]));
    assign layer4_outputs[3949] = layer3_outputs[2185];
    assign layer4_outputs[3950] = (layer3_outputs[2095]) | (layer3_outputs[4511]);
    assign layer4_outputs[3951] = layer3_outputs[2988];
    assign layer4_outputs[3952] = ~(layer3_outputs[823]);
    assign layer4_outputs[3953] = 1'b0;
    assign layer4_outputs[3954] = ~(layer3_outputs[2271]);
    assign layer4_outputs[3955] = ~(layer3_outputs[3179]);
    assign layer4_outputs[3956] = ~(layer3_outputs[3046]);
    assign layer4_outputs[3957] = ~(layer3_outputs[3024]);
    assign layer4_outputs[3958] = layer3_outputs[2131];
    assign layer4_outputs[3959] = ~((layer3_outputs[4137]) & (layer3_outputs[846]));
    assign layer4_outputs[3960] = ~(layer3_outputs[2148]);
    assign layer4_outputs[3961] = ~(layer3_outputs[1558]);
    assign layer4_outputs[3962] = (layer3_outputs[127]) | (layer3_outputs[4627]);
    assign layer4_outputs[3963] = (layer3_outputs[2379]) ^ (layer3_outputs[2901]);
    assign layer4_outputs[3964] = layer3_outputs[1831];
    assign layer4_outputs[3965] = (layer3_outputs[2187]) & ~(layer3_outputs[2916]);
    assign layer4_outputs[3966] = ~(layer3_outputs[2199]) | (layer3_outputs[960]);
    assign layer4_outputs[3967] = ~((layer3_outputs[3203]) & (layer3_outputs[3618]));
    assign layer4_outputs[3968] = (layer3_outputs[314]) ^ (layer3_outputs[3362]);
    assign layer4_outputs[3969] = ~(layer3_outputs[3463]);
    assign layer4_outputs[3970] = ~(layer3_outputs[1201]) | (layer3_outputs[4713]);
    assign layer4_outputs[3971] = (layer3_outputs[2068]) ^ (layer3_outputs[5018]);
    assign layer4_outputs[3972] = ~(layer3_outputs[2655]);
    assign layer4_outputs[3973] = ~(layer3_outputs[1672]);
    assign layer4_outputs[3974] = (layer3_outputs[403]) & ~(layer3_outputs[2285]);
    assign layer4_outputs[3975] = 1'b0;
    assign layer4_outputs[3976] = ~((layer3_outputs[1337]) ^ (layer3_outputs[3789]));
    assign layer4_outputs[3977] = (layer3_outputs[1749]) & (layer3_outputs[3955]);
    assign layer4_outputs[3978] = layer3_outputs[2685];
    assign layer4_outputs[3979] = ~(layer3_outputs[2402]);
    assign layer4_outputs[3980] = ~(layer3_outputs[1041]);
    assign layer4_outputs[3981] = (layer3_outputs[4535]) | (layer3_outputs[4331]);
    assign layer4_outputs[3982] = ~(layer3_outputs[4163]) | (layer3_outputs[4944]);
    assign layer4_outputs[3983] = layer3_outputs[545];
    assign layer4_outputs[3984] = layer3_outputs[4217];
    assign layer4_outputs[3985] = ~((layer3_outputs[4599]) ^ (layer3_outputs[3490]));
    assign layer4_outputs[3986] = layer3_outputs[1826];
    assign layer4_outputs[3987] = layer3_outputs[3794];
    assign layer4_outputs[3988] = layer3_outputs[3661];
    assign layer4_outputs[3989] = ~((layer3_outputs[1463]) | (layer3_outputs[4071]));
    assign layer4_outputs[3990] = layer3_outputs[5016];
    assign layer4_outputs[3991] = (layer3_outputs[1473]) & ~(layer3_outputs[4008]);
    assign layer4_outputs[3992] = ~(layer3_outputs[4814]);
    assign layer4_outputs[3993] = ~((layer3_outputs[1111]) & (layer3_outputs[2602]));
    assign layer4_outputs[3994] = ~((layer3_outputs[2019]) | (layer3_outputs[498]));
    assign layer4_outputs[3995] = ~(layer3_outputs[52]);
    assign layer4_outputs[3996] = ~((layer3_outputs[2993]) & (layer3_outputs[2330]));
    assign layer4_outputs[3997] = ~(layer3_outputs[5009]);
    assign layer4_outputs[3998] = (layer3_outputs[1143]) & ~(layer3_outputs[190]);
    assign layer4_outputs[3999] = layer3_outputs[1516];
    assign layer4_outputs[4000] = 1'b0;
    assign layer4_outputs[4001] = ~(layer3_outputs[2165]);
    assign layer4_outputs[4002] = (layer3_outputs[82]) ^ (layer3_outputs[4251]);
    assign layer4_outputs[4003] = 1'b0;
    assign layer4_outputs[4004] = (layer3_outputs[210]) | (layer3_outputs[498]);
    assign layer4_outputs[4005] = (layer3_outputs[5023]) & ~(layer3_outputs[614]);
    assign layer4_outputs[4006] = ~(layer3_outputs[5069]) | (layer3_outputs[4878]);
    assign layer4_outputs[4007] = (layer3_outputs[1469]) ^ (layer3_outputs[3164]);
    assign layer4_outputs[4008] = layer3_outputs[3019];
    assign layer4_outputs[4009] = ~(layer3_outputs[2442]);
    assign layer4_outputs[4010] = (layer3_outputs[4437]) ^ (layer3_outputs[737]);
    assign layer4_outputs[4011] = layer3_outputs[1894];
    assign layer4_outputs[4012] = (layer3_outputs[3522]) & (layer3_outputs[3612]);
    assign layer4_outputs[4013] = ~(layer3_outputs[3246]) | (layer3_outputs[404]);
    assign layer4_outputs[4014] = 1'b1;
    assign layer4_outputs[4015] = ~(layer3_outputs[2269]) | (layer3_outputs[3999]);
    assign layer4_outputs[4016] = (layer3_outputs[753]) & ~(layer3_outputs[3157]);
    assign layer4_outputs[4017] = layer3_outputs[2719];
    assign layer4_outputs[4018] = ~(layer3_outputs[1412]) | (layer3_outputs[1677]);
    assign layer4_outputs[4019] = (layer3_outputs[2356]) & ~(layer3_outputs[507]);
    assign layer4_outputs[4020] = layer3_outputs[4698];
    assign layer4_outputs[4021] = ~(layer3_outputs[1999]);
    assign layer4_outputs[4022] = 1'b1;
    assign layer4_outputs[4023] = ~((layer3_outputs[3214]) & (layer3_outputs[856]));
    assign layer4_outputs[4024] = ~(layer3_outputs[9]);
    assign layer4_outputs[4025] = (layer3_outputs[4409]) | (layer3_outputs[4822]);
    assign layer4_outputs[4026] = ~((layer3_outputs[4141]) & (layer3_outputs[2396]));
    assign layer4_outputs[4027] = ~(layer3_outputs[4889]) | (layer3_outputs[578]);
    assign layer4_outputs[4028] = (layer3_outputs[1564]) | (layer3_outputs[1512]);
    assign layer4_outputs[4029] = (layer3_outputs[661]) & ~(layer3_outputs[2414]);
    assign layer4_outputs[4030] = ~((layer3_outputs[505]) & (layer3_outputs[88]));
    assign layer4_outputs[4031] = ~(layer3_outputs[4520]);
    assign layer4_outputs[4032] = layer3_outputs[4262];
    assign layer4_outputs[4033] = ~(layer3_outputs[3620]);
    assign layer4_outputs[4034] = layer3_outputs[1948];
    assign layer4_outputs[4035] = ~((layer3_outputs[971]) | (layer3_outputs[1153]));
    assign layer4_outputs[4036] = ~(layer3_outputs[4489]) | (layer3_outputs[1975]);
    assign layer4_outputs[4037] = ~(layer3_outputs[450]) | (layer3_outputs[1277]);
    assign layer4_outputs[4038] = 1'b1;
    assign layer4_outputs[4039] = (layer3_outputs[2744]) & (layer3_outputs[4312]);
    assign layer4_outputs[4040] = ~((layer3_outputs[1417]) & (layer3_outputs[4316]));
    assign layer4_outputs[4041] = layer3_outputs[3374];
    assign layer4_outputs[4042] = (layer3_outputs[2107]) ^ (layer3_outputs[1038]);
    assign layer4_outputs[4043] = ~(layer3_outputs[342]) | (layer3_outputs[670]);
    assign layer4_outputs[4044] = ~(layer3_outputs[5001]);
    assign layer4_outputs[4045] = layer3_outputs[4871];
    assign layer4_outputs[4046] = layer3_outputs[1642];
    assign layer4_outputs[4047] = ~(layer3_outputs[1506]);
    assign layer4_outputs[4048] = ~((layer3_outputs[585]) | (layer3_outputs[2446]));
    assign layer4_outputs[4049] = layer3_outputs[3229];
    assign layer4_outputs[4050] = ~((layer3_outputs[349]) | (layer3_outputs[925]));
    assign layer4_outputs[4051] = layer3_outputs[4246];
    assign layer4_outputs[4052] = layer3_outputs[4848];
    assign layer4_outputs[4053] = (layer3_outputs[1544]) ^ (layer3_outputs[4562]);
    assign layer4_outputs[4054] = layer3_outputs[4253];
    assign layer4_outputs[4055] = ~(layer3_outputs[1624]);
    assign layer4_outputs[4056] = layer3_outputs[888];
    assign layer4_outputs[4057] = ~(layer3_outputs[637]);
    assign layer4_outputs[4058] = layer3_outputs[1216];
    assign layer4_outputs[4059] = (layer3_outputs[4070]) & ~(layer3_outputs[3619]);
    assign layer4_outputs[4060] = 1'b0;
    assign layer4_outputs[4061] = layer3_outputs[1717];
    assign layer4_outputs[4062] = (layer3_outputs[2096]) & ~(layer3_outputs[3206]);
    assign layer4_outputs[4063] = layer3_outputs[2278];
    assign layer4_outputs[4064] = ~(layer3_outputs[3557]);
    assign layer4_outputs[4065] = ~((layer3_outputs[2038]) | (layer3_outputs[3261]));
    assign layer4_outputs[4066] = ~(layer3_outputs[1865]);
    assign layer4_outputs[4067] = (layer3_outputs[3727]) & ~(layer3_outputs[4629]);
    assign layer4_outputs[4068] = ~((layer3_outputs[1610]) | (layer3_outputs[1801]));
    assign layer4_outputs[4069] = ~((layer3_outputs[2397]) ^ (layer3_outputs[1378]));
    assign layer4_outputs[4070] = ~(layer3_outputs[4028]);
    assign layer4_outputs[4071] = ~(layer3_outputs[1905]);
    assign layer4_outputs[4072] = (layer3_outputs[2801]) & ~(layer3_outputs[852]);
    assign layer4_outputs[4073] = ~(layer3_outputs[235]);
    assign layer4_outputs[4074] = (layer3_outputs[305]) & ~(layer3_outputs[2824]);
    assign layer4_outputs[4075] = (layer3_outputs[11]) & (layer3_outputs[4652]);
    assign layer4_outputs[4076] = (layer3_outputs[345]) & ~(layer3_outputs[4130]);
    assign layer4_outputs[4077] = (layer3_outputs[2843]) | (layer3_outputs[1332]);
    assign layer4_outputs[4078] = (layer3_outputs[1768]) & ~(layer3_outputs[996]);
    assign layer4_outputs[4079] = ~(layer3_outputs[790]) | (layer3_outputs[1871]);
    assign layer4_outputs[4080] = ~((layer3_outputs[3027]) | (layer3_outputs[3896]));
    assign layer4_outputs[4081] = (layer3_outputs[309]) | (layer3_outputs[2155]);
    assign layer4_outputs[4082] = layer3_outputs[3332];
    assign layer4_outputs[4083] = ~(layer3_outputs[1495]);
    assign layer4_outputs[4084] = (layer3_outputs[4703]) | (layer3_outputs[1936]);
    assign layer4_outputs[4085] = ~(layer3_outputs[4110]) | (layer3_outputs[1728]);
    assign layer4_outputs[4086] = ~(layer3_outputs[1019]) | (layer3_outputs[627]);
    assign layer4_outputs[4087] = (layer3_outputs[613]) | (layer3_outputs[3013]);
    assign layer4_outputs[4088] = ~((layer3_outputs[3345]) | (layer3_outputs[4393]));
    assign layer4_outputs[4089] = (layer3_outputs[1224]) | (layer3_outputs[3102]);
    assign layer4_outputs[4090] = ~(layer3_outputs[4375]);
    assign layer4_outputs[4091] = layer3_outputs[1116];
    assign layer4_outputs[4092] = ~((layer3_outputs[2234]) | (layer3_outputs[848]));
    assign layer4_outputs[4093] = (layer3_outputs[4291]) ^ (layer3_outputs[3381]);
    assign layer4_outputs[4094] = ~(layer3_outputs[1994]) | (layer3_outputs[209]);
    assign layer4_outputs[4095] = ~(layer3_outputs[2772]);
    assign layer4_outputs[4096] = layer3_outputs[4360];
    assign layer4_outputs[4097] = layer3_outputs[2711];
    assign layer4_outputs[4098] = 1'b0;
    assign layer4_outputs[4099] = layer3_outputs[507];
    assign layer4_outputs[4100] = layer3_outputs[1318];
    assign layer4_outputs[4101] = (layer3_outputs[810]) & (layer3_outputs[1652]);
    assign layer4_outputs[4102] = (layer3_outputs[676]) | (layer3_outputs[518]);
    assign layer4_outputs[4103] = layer3_outputs[1971];
    assign layer4_outputs[4104] = (layer3_outputs[260]) & ~(layer3_outputs[4578]);
    assign layer4_outputs[4105] = layer3_outputs[3610];
    assign layer4_outputs[4106] = ~(layer3_outputs[3752]) | (layer3_outputs[2355]);
    assign layer4_outputs[4107] = (layer3_outputs[1102]) ^ (layer3_outputs[652]);
    assign layer4_outputs[4108] = ~(layer3_outputs[3486]);
    assign layer4_outputs[4109] = (layer3_outputs[2025]) & ~(layer3_outputs[1434]);
    assign layer4_outputs[4110] = (layer3_outputs[5072]) ^ (layer3_outputs[970]);
    assign layer4_outputs[4111] = (layer3_outputs[4607]) & ~(layer3_outputs[3107]);
    assign layer4_outputs[4112] = layer3_outputs[4591];
    assign layer4_outputs[4113] = ~(layer3_outputs[4935]) | (layer3_outputs[2876]);
    assign layer4_outputs[4114] = (layer3_outputs[2832]) | (layer3_outputs[3807]);
    assign layer4_outputs[4115] = 1'b1;
    assign layer4_outputs[4116] = (layer3_outputs[3733]) | (layer3_outputs[5051]);
    assign layer4_outputs[4117] = layer3_outputs[249];
    assign layer4_outputs[4118] = (layer3_outputs[4320]) & ~(layer3_outputs[1927]);
    assign layer4_outputs[4119] = (layer3_outputs[1477]) & (layer3_outputs[2567]);
    assign layer4_outputs[4120] = ~(layer3_outputs[2352]) | (layer3_outputs[3722]);
    assign layer4_outputs[4121] = ~((layer3_outputs[276]) | (layer3_outputs[91]));
    assign layer4_outputs[4122] = ~(layer3_outputs[2721]);
    assign layer4_outputs[4123] = (layer3_outputs[3078]) | (layer3_outputs[973]);
    assign layer4_outputs[4124] = (layer3_outputs[4694]) & (layer3_outputs[2315]);
    assign layer4_outputs[4125] = ~(layer3_outputs[2216]) | (layer3_outputs[2191]);
    assign layer4_outputs[4126] = ~(layer3_outputs[2907]);
    assign layer4_outputs[4127] = ~(layer3_outputs[4598]);
    assign layer4_outputs[4128] = ~(layer3_outputs[1749]);
    assign layer4_outputs[4129] = (layer3_outputs[4921]) | (layer3_outputs[1397]);
    assign layer4_outputs[4130] = ~((layer3_outputs[4621]) ^ (layer3_outputs[2138]));
    assign layer4_outputs[4131] = layer3_outputs[3678];
    assign layer4_outputs[4132] = (layer3_outputs[1901]) & (layer3_outputs[126]);
    assign layer4_outputs[4133] = layer3_outputs[4975];
    assign layer4_outputs[4134] = ~((layer3_outputs[3665]) & (layer3_outputs[3572]));
    assign layer4_outputs[4135] = ~(layer3_outputs[2034]);
    assign layer4_outputs[4136] = ~(layer3_outputs[1421]);
    assign layer4_outputs[4137] = layer3_outputs[2809];
    assign layer4_outputs[4138] = layer3_outputs[2953];
    assign layer4_outputs[4139] = ~((layer3_outputs[2148]) | (layer3_outputs[3691]));
    assign layer4_outputs[4140] = (layer3_outputs[2642]) & ~(layer3_outputs[3804]);
    assign layer4_outputs[4141] = ~(layer3_outputs[265]);
    assign layer4_outputs[4142] = ~(layer3_outputs[4935]);
    assign layer4_outputs[4143] = (layer3_outputs[3750]) & (layer3_outputs[3135]);
    assign layer4_outputs[4144] = ~(layer3_outputs[4069]) | (layer3_outputs[219]);
    assign layer4_outputs[4145] = layer3_outputs[668];
    assign layer4_outputs[4146] = layer3_outputs[691];
    assign layer4_outputs[4147] = 1'b0;
    assign layer4_outputs[4148] = (layer3_outputs[206]) & (layer3_outputs[298]);
    assign layer4_outputs[4149] = ~(layer3_outputs[2464]);
    assign layer4_outputs[4150] = ~(layer3_outputs[4777]);
    assign layer4_outputs[4151] = ~(layer3_outputs[550]) | (layer3_outputs[3984]);
    assign layer4_outputs[4152] = (layer3_outputs[4236]) & ~(layer3_outputs[2061]);
    assign layer4_outputs[4153] = (layer3_outputs[1709]) & ~(layer3_outputs[2728]);
    assign layer4_outputs[4154] = ~(layer3_outputs[2879]);
    assign layer4_outputs[4155] = ~(layer3_outputs[449]);
    assign layer4_outputs[4156] = 1'b1;
    assign layer4_outputs[4157] = ~(layer3_outputs[1021]) | (layer3_outputs[1757]);
    assign layer4_outputs[4158] = (layer3_outputs[188]) ^ (layer3_outputs[3811]);
    assign layer4_outputs[4159] = ~((layer3_outputs[2376]) ^ (layer3_outputs[2348]));
    assign layer4_outputs[4160] = 1'b0;
    assign layer4_outputs[4161] = (layer3_outputs[2548]) ^ (layer3_outputs[4200]);
    assign layer4_outputs[4162] = layer3_outputs[4669];
    assign layer4_outputs[4163] = ~(layer3_outputs[3453]);
    assign layer4_outputs[4164] = ~(layer3_outputs[769]);
    assign layer4_outputs[4165] = ~((layer3_outputs[3280]) | (layer3_outputs[4764]));
    assign layer4_outputs[4166] = (layer3_outputs[1347]) | (layer3_outputs[1596]);
    assign layer4_outputs[4167] = (layer3_outputs[4079]) & ~(layer3_outputs[3585]);
    assign layer4_outputs[4168] = ~(layer3_outputs[5077]) | (layer3_outputs[2625]);
    assign layer4_outputs[4169] = ~(layer3_outputs[1187]);
    assign layer4_outputs[4170] = ~(layer3_outputs[2180]) | (layer3_outputs[23]);
    assign layer4_outputs[4171] = 1'b0;
    assign layer4_outputs[4172] = ~(layer3_outputs[1377]);
    assign layer4_outputs[4173] = (layer3_outputs[3227]) & ~(layer3_outputs[2811]);
    assign layer4_outputs[4174] = ~((layer3_outputs[2489]) | (layer3_outputs[936]));
    assign layer4_outputs[4175] = (layer3_outputs[658]) & (layer3_outputs[2912]);
    assign layer4_outputs[4176] = ~(layer3_outputs[2915]) | (layer3_outputs[1643]);
    assign layer4_outputs[4177] = ~(layer3_outputs[3381]);
    assign layer4_outputs[4178] = (layer3_outputs[2304]) | (layer3_outputs[779]);
    assign layer4_outputs[4179] = ~(layer3_outputs[1101]) | (layer3_outputs[4986]);
    assign layer4_outputs[4180] = ~(layer3_outputs[3325]);
    assign layer4_outputs[4181] = ~((layer3_outputs[18]) & (layer3_outputs[819]));
    assign layer4_outputs[4182] = layer3_outputs[2536];
    assign layer4_outputs[4183] = (layer3_outputs[2696]) & ~(layer3_outputs[4145]);
    assign layer4_outputs[4184] = ~((layer3_outputs[2607]) & (layer3_outputs[4453]));
    assign layer4_outputs[4185] = (layer3_outputs[1341]) & ~(layer3_outputs[885]);
    assign layer4_outputs[4186] = ~(layer3_outputs[1913]);
    assign layer4_outputs[4187] = ~(layer3_outputs[2436]) | (layer3_outputs[357]);
    assign layer4_outputs[4188] = layer3_outputs[4258];
    assign layer4_outputs[4189] = ~(layer3_outputs[3955]);
    assign layer4_outputs[4190] = ~(layer3_outputs[2480]) | (layer3_outputs[998]);
    assign layer4_outputs[4191] = (layer3_outputs[3561]) ^ (layer3_outputs[747]);
    assign layer4_outputs[4192] = ~(layer3_outputs[4381]);
    assign layer4_outputs[4193] = ~((layer3_outputs[2870]) ^ (layer3_outputs[3449]));
    assign layer4_outputs[4194] = layer3_outputs[1696];
    assign layer4_outputs[4195] = ~(layer3_outputs[561]);
    assign layer4_outputs[4196] = ~(layer3_outputs[2946]);
    assign layer4_outputs[4197] = ~((layer3_outputs[2378]) | (layer3_outputs[2025]));
    assign layer4_outputs[4198] = layer3_outputs[2959];
    assign layer4_outputs[4199] = (layer3_outputs[3222]) ^ (layer3_outputs[3967]);
    assign layer4_outputs[4200] = ~(layer3_outputs[3537]) | (layer3_outputs[320]);
    assign layer4_outputs[4201] = ~(layer3_outputs[3831]) | (layer3_outputs[3179]);
    assign layer4_outputs[4202] = (layer3_outputs[4846]) | (layer3_outputs[239]);
    assign layer4_outputs[4203] = ~(layer3_outputs[3058]);
    assign layer4_outputs[4204] = ~(layer3_outputs[528]);
    assign layer4_outputs[4205] = layer3_outputs[4296];
    assign layer4_outputs[4206] = layer3_outputs[2758];
    assign layer4_outputs[4207] = ~((layer3_outputs[1186]) & (layer3_outputs[2592]));
    assign layer4_outputs[4208] = layer3_outputs[2877];
    assign layer4_outputs[4209] = (layer3_outputs[4901]) | (layer3_outputs[2623]);
    assign layer4_outputs[4210] = ~(layer3_outputs[2283]) | (layer3_outputs[1004]);
    assign layer4_outputs[4211] = ~(layer3_outputs[1716]);
    assign layer4_outputs[4212] = ~(layer3_outputs[1686]) | (layer3_outputs[1754]);
    assign layer4_outputs[4213] = ~(layer3_outputs[2159]);
    assign layer4_outputs[4214] = ~((layer3_outputs[2650]) | (layer3_outputs[4651]));
    assign layer4_outputs[4215] = layer3_outputs[3521];
    assign layer4_outputs[4216] = ~(layer3_outputs[4374]);
    assign layer4_outputs[4217] = ~(layer3_outputs[1162]);
    assign layer4_outputs[4218] = ~(layer3_outputs[3607]);
    assign layer4_outputs[4219] = 1'b1;
    assign layer4_outputs[4220] = (layer3_outputs[815]) & ~(layer3_outputs[2806]);
    assign layer4_outputs[4221] = ~((layer3_outputs[1623]) & (layer3_outputs[3136]));
    assign layer4_outputs[4222] = ~(layer3_outputs[4592]) | (layer3_outputs[3202]);
    assign layer4_outputs[4223] = (layer3_outputs[4186]) & ~(layer3_outputs[4758]);
    assign layer4_outputs[4224] = (layer3_outputs[465]) & (layer3_outputs[2247]);
    assign layer4_outputs[4225] = ~(layer3_outputs[2075]) | (layer3_outputs[336]);
    assign layer4_outputs[4226] = (layer3_outputs[4771]) | (layer3_outputs[1237]);
    assign layer4_outputs[4227] = ~(layer3_outputs[1065]);
    assign layer4_outputs[4228] = 1'b0;
    assign layer4_outputs[4229] = ~((layer3_outputs[3571]) | (layer3_outputs[1450]));
    assign layer4_outputs[4230] = ~((layer3_outputs[4073]) & (layer3_outputs[1949]));
    assign layer4_outputs[4231] = ~(layer3_outputs[4923]) | (layer3_outputs[882]);
    assign layer4_outputs[4232] = ~((layer3_outputs[2458]) ^ (layer3_outputs[413]));
    assign layer4_outputs[4233] = (layer3_outputs[4925]) | (layer3_outputs[1751]);
    assign layer4_outputs[4234] = ~((layer3_outputs[1576]) & (layer3_outputs[1301]));
    assign layer4_outputs[4235] = (layer3_outputs[455]) & ~(layer3_outputs[1944]);
    assign layer4_outputs[4236] = layer3_outputs[2603];
    assign layer4_outputs[4237] = ~(layer3_outputs[1836]) | (layer3_outputs[259]);
    assign layer4_outputs[4238] = (layer3_outputs[1363]) | (layer3_outputs[830]);
    assign layer4_outputs[4239] = ~((layer3_outputs[4646]) | (layer3_outputs[3351]));
    assign layer4_outputs[4240] = ~(layer3_outputs[3893]);
    assign layer4_outputs[4241] = (layer3_outputs[2760]) & ~(layer3_outputs[3424]);
    assign layer4_outputs[4242] = ~((layer3_outputs[2855]) ^ (layer3_outputs[2181]));
    assign layer4_outputs[4243] = ~(layer3_outputs[2767]);
    assign layer4_outputs[4244] = (layer3_outputs[1985]) & (layer3_outputs[1578]);
    assign layer4_outputs[4245] = ~(layer3_outputs[4595]);
    assign layer4_outputs[4246] = ~(layer3_outputs[4297]);
    assign layer4_outputs[4247] = ~(layer3_outputs[2803]);
    assign layer4_outputs[4248] = layer3_outputs[4172];
    assign layer4_outputs[4249] = (layer3_outputs[2892]) & (layer3_outputs[3197]);
    assign layer4_outputs[4250] = ~(layer3_outputs[321]);
    assign layer4_outputs[4251] = (layer3_outputs[110]) | (layer3_outputs[1406]);
    assign layer4_outputs[4252] = layer3_outputs[691];
    assign layer4_outputs[4253] = layer3_outputs[3912];
    assign layer4_outputs[4254] = layer3_outputs[3435];
    assign layer4_outputs[4255] = (layer3_outputs[69]) | (layer3_outputs[3304]);
    assign layer4_outputs[4256] = (layer3_outputs[4962]) & ~(layer3_outputs[2997]);
    assign layer4_outputs[4257] = ~((layer3_outputs[1481]) & (layer3_outputs[2975]));
    assign layer4_outputs[4258] = ~((layer3_outputs[2789]) | (layer3_outputs[2508]));
    assign layer4_outputs[4259] = (layer3_outputs[1896]) | (layer3_outputs[3395]);
    assign layer4_outputs[4260] = (layer3_outputs[2058]) ^ (layer3_outputs[4085]);
    assign layer4_outputs[4261] = 1'b0;
    assign layer4_outputs[4262] = layer3_outputs[3924];
    assign layer4_outputs[4263] = ~(layer3_outputs[364]) | (layer3_outputs[3010]);
    assign layer4_outputs[4264] = layer3_outputs[4462];
    assign layer4_outputs[4265] = (layer3_outputs[3042]) & (layer3_outputs[50]);
    assign layer4_outputs[4266] = layer3_outputs[2538];
    assign layer4_outputs[4267] = layer3_outputs[182];
    assign layer4_outputs[4268] = ~(layer3_outputs[4755]) | (layer3_outputs[3747]);
    assign layer4_outputs[4269] = layer3_outputs[1264];
    assign layer4_outputs[4270] = layer3_outputs[4134];
    assign layer4_outputs[4271] = (layer3_outputs[4483]) & ~(layer3_outputs[2963]);
    assign layer4_outputs[4272] = layer3_outputs[2217];
    assign layer4_outputs[4273] = ~(layer3_outputs[4407]);
    assign layer4_outputs[4274] = (layer3_outputs[3535]) & (layer3_outputs[2624]);
    assign layer4_outputs[4275] = layer3_outputs[4956];
    assign layer4_outputs[4276] = ~(layer3_outputs[2532]) | (layer3_outputs[713]);
    assign layer4_outputs[4277] = layer3_outputs[4289];
    assign layer4_outputs[4278] = layer3_outputs[134];
    assign layer4_outputs[4279] = ~(layer3_outputs[2496]) | (layer3_outputs[105]);
    assign layer4_outputs[4280] = (layer3_outputs[4278]) & (layer3_outputs[3876]);
    assign layer4_outputs[4281] = 1'b1;
    assign layer4_outputs[4282] = ~(layer3_outputs[3255]) | (layer3_outputs[4316]);
    assign layer4_outputs[4283] = (layer3_outputs[3916]) | (layer3_outputs[853]);
    assign layer4_outputs[4284] = (layer3_outputs[950]) | (layer3_outputs[156]);
    assign layer4_outputs[4285] = ~(layer3_outputs[110]) | (layer3_outputs[3529]);
    assign layer4_outputs[4286] = ~(layer3_outputs[39]) | (layer3_outputs[4685]);
    assign layer4_outputs[4287] = layer3_outputs[1220];
    assign layer4_outputs[4288] = layer3_outputs[1333];
    assign layer4_outputs[4289] = layer3_outputs[5012];
    assign layer4_outputs[4290] = ~(layer3_outputs[3193]) | (layer3_outputs[2775]);
    assign layer4_outputs[4291] = (layer3_outputs[4347]) | (layer3_outputs[4102]);
    assign layer4_outputs[4292] = (layer3_outputs[2691]) & ~(layer3_outputs[3641]);
    assign layer4_outputs[4293] = ~(layer3_outputs[3166]);
    assign layer4_outputs[4294] = (layer3_outputs[1386]) & ~(layer3_outputs[2893]);
    assign layer4_outputs[4295] = ~(layer3_outputs[4358]) | (layer3_outputs[4466]);
    assign layer4_outputs[4296] = (layer3_outputs[228]) ^ (layer3_outputs[644]);
    assign layer4_outputs[4297] = (layer3_outputs[2535]) & (layer3_outputs[952]);
    assign layer4_outputs[4298] = ~((layer3_outputs[1565]) & (layer3_outputs[4709]));
    assign layer4_outputs[4299] = ~((layer3_outputs[1662]) ^ (layer3_outputs[3717]));
    assign layer4_outputs[4300] = ~(layer3_outputs[2991]);
    assign layer4_outputs[4301] = ~((layer3_outputs[323]) | (layer3_outputs[2543]));
    assign layer4_outputs[4302] = ~((layer3_outputs[1084]) & (layer3_outputs[3729]));
    assign layer4_outputs[4303] = layer3_outputs[1833];
    assign layer4_outputs[4304] = 1'b1;
    assign layer4_outputs[4305] = layer3_outputs[757];
    assign layer4_outputs[4306] = 1'b0;
    assign layer4_outputs[4307] = ~(layer3_outputs[280]) | (layer3_outputs[4414]);
    assign layer4_outputs[4308] = 1'b0;
    assign layer4_outputs[4309] = ~(layer3_outputs[638]) | (layer3_outputs[2255]);
    assign layer4_outputs[4310] = ~(layer3_outputs[4684]);
    assign layer4_outputs[4311] = ~(layer3_outputs[4225]);
    assign layer4_outputs[4312] = layer3_outputs[4589];
    assign layer4_outputs[4313] = ~((layer3_outputs[3290]) | (layer3_outputs[2971]));
    assign layer4_outputs[4314] = (layer3_outputs[3128]) & ~(layer3_outputs[448]);
    assign layer4_outputs[4315] = layer3_outputs[4866];
    assign layer4_outputs[4316] = ~(layer3_outputs[4298]);
    assign layer4_outputs[4317] = (layer3_outputs[4476]) & ~(layer3_outputs[2836]);
    assign layer4_outputs[4318] = (layer3_outputs[4459]) & ~(layer3_outputs[2073]);
    assign layer4_outputs[4319] = layer3_outputs[2874];
    assign layer4_outputs[4320] = layer3_outputs[145];
    assign layer4_outputs[4321] = layer3_outputs[5077];
    assign layer4_outputs[4322] = 1'b0;
    assign layer4_outputs[4323] = (layer3_outputs[1419]) & ~(layer3_outputs[2271]);
    assign layer4_outputs[4324] = (layer3_outputs[881]) & (layer3_outputs[4115]);
    assign layer4_outputs[4325] = (layer3_outputs[3786]) & (layer3_outputs[2705]);
    assign layer4_outputs[4326] = ~(layer3_outputs[3979]) | (layer3_outputs[4596]);
    assign layer4_outputs[4327] = (layer3_outputs[4733]) & ~(layer3_outputs[1411]);
    assign layer4_outputs[4328] = layer3_outputs[2325];
    assign layer4_outputs[4329] = layer3_outputs[776];
    assign layer4_outputs[4330] = ~((layer3_outputs[4363]) | (layer3_outputs[4354]));
    assign layer4_outputs[4331] = 1'b0;
    assign layer4_outputs[4332] = layer3_outputs[3102];
    assign layer4_outputs[4333] = (layer3_outputs[995]) & ~(layer3_outputs[2923]);
    assign layer4_outputs[4334] = layer3_outputs[5];
    assign layer4_outputs[4335] = ~((layer3_outputs[5088]) & (layer3_outputs[4118]));
    assign layer4_outputs[4336] = ~(layer3_outputs[2743]);
    assign layer4_outputs[4337] = layer3_outputs[5090];
    assign layer4_outputs[4338] = 1'b1;
    assign layer4_outputs[4339] = ~(layer3_outputs[1503]);
    assign layer4_outputs[4340] = ~(layer3_outputs[4921]);
    assign layer4_outputs[4341] = (layer3_outputs[626]) & ~(layer3_outputs[1587]);
    assign layer4_outputs[4342] = ~(layer3_outputs[1085]) | (layer3_outputs[2114]);
    assign layer4_outputs[4343] = layer3_outputs[660];
    assign layer4_outputs[4344] = ~((layer3_outputs[4610]) | (layer3_outputs[4432]));
    assign layer4_outputs[4345] = (layer3_outputs[3306]) & ~(layer3_outputs[1819]);
    assign layer4_outputs[4346] = ~(layer3_outputs[3693]);
    assign layer4_outputs[4347] = ~(layer3_outputs[3680]);
    assign layer4_outputs[4348] = ~(layer3_outputs[3239]);
    assign layer4_outputs[4349] = (layer3_outputs[3873]) ^ (layer3_outputs[4350]);
    assign layer4_outputs[4350] = 1'b0;
    assign layer4_outputs[4351] = layer3_outputs[1310];
    assign layer4_outputs[4352] = layer3_outputs[2561];
    assign layer4_outputs[4353] = (layer3_outputs[53]) & (layer3_outputs[4946]);
    assign layer4_outputs[4354] = (layer3_outputs[3515]) ^ (layer3_outputs[1235]);
    assign layer4_outputs[4355] = ~(layer3_outputs[746]) | (layer3_outputs[1601]);
    assign layer4_outputs[4356] = (layer3_outputs[4198]) & ~(layer3_outputs[2739]);
    assign layer4_outputs[4357] = 1'b1;
    assign layer4_outputs[4358] = layer3_outputs[1635];
    assign layer4_outputs[4359] = (layer3_outputs[4044]) & (layer3_outputs[1535]);
    assign layer4_outputs[4360] = ~((layer3_outputs[103]) & (layer3_outputs[2808]));
    assign layer4_outputs[4361] = layer3_outputs[4566];
    assign layer4_outputs[4362] = layer3_outputs[1984];
    assign layer4_outputs[4363] = (layer3_outputs[1157]) & ~(layer3_outputs[5096]);
    assign layer4_outputs[4364] = ~(layer3_outputs[3813]);
    assign layer4_outputs[4365] = ~(layer3_outputs[4613]) | (layer3_outputs[4523]);
    assign layer4_outputs[4366] = ~((layer3_outputs[5067]) & (layer3_outputs[554]));
    assign layer4_outputs[4367] = 1'b0;
    assign layer4_outputs[4368] = (layer3_outputs[4956]) | (layer3_outputs[4933]);
    assign layer4_outputs[4369] = layer3_outputs[124];
    assign layer4_outputs[4370] = ~(layer3_outputs[1117]);
    assign layer4_outputs[4371] = ~(layer3_outputs[4851]);
    assign layer4_outputs[4372] = 1'b1;
    assign layer4_outputs[4373] = ~(layer3_outputs[3643]);
    assign layer4_outputs[4374] = ~(layer3_outputs[3156]);
    assign layer4_outputs[4375] = (layer3_outputs[1239]) ^ (layer3_outputs[2977]);
    assign layer4_outputs[4376] = layer3_outputs[968];
    assign layer4_outputs[4377] = ~(layer3_outputs[599]);
    assign layer4_outputs[4378] = ~((layer3_outputs[2400]) & (layer3_outputs[2225]));
    assign layer4_outputs[4379] = layer3_outputs[215];
    assign layer4_outputs[4380] = ~(layer3_outputs[1329]) | (layer3_outputs[398]);
    assign layer4_outputs[4381] = layer3_outputs[2183];
    assign layer4_outputs[4382] = ~(layer3_outputs[2529]);
    assign layer4_outputs[4383] = ~(layer3_outputs[391]) | (layer3_outputs[2677]);
    assign layer4_outputs[4384] = (layer3_outputs[540]) ^ (layer3_outputs[4934]);
    assign layer4_outputs[4385] = (layer3_outputs[4282]) & ~(layer3_outputs[382]);
    assign layer4_outputs[4386] = ~(layer3_outputs[1488]);
    assign layer4_outputs[4387] = ~((layer3_outputs[5059]) | (layer3_outputs[4770]));
    assign layer4_outputs[4388] = 1'b0;
    assign layer4_outputs[4389] = ~((layer3_outputs[4910]) & (layer3_outputs[634]));
    assign layer4_outputs[4390] = ~(layer3_outputs[4873]);
    assign layer4_outputs[4391] = ~(layer3_outputs[3230]) | (layer3_outputs[755]);
    assign layer4_outputs[4392] = ~(layer3_outputs[4849]) | (layer3_outputs[3079]);
    assign layer4_outputs[4393] = ~(layer3_outputs[1265]);
    assign layer4_outputs[4394] = ~(layer3_outputs[4673]);
    assign layer4_outputs[4395] = layer3_outputs[2031];
    assign layer4_outputs[4396] = ~(layer3_outputs[2573]);
    assign layer4_outputs[4397] = layer3_outputs[1945];
    assign layer4_outputs[4398] = ~((layer3_outputs[3592]) ^ (layer3_outputs[976]));
    assign layer4_outputs[4399] = ~(layer3_outputs[4644]);
    assign layer4_outputs[4400] = layer3_outputs[1702];
    assign layer4_outputs[4401] = ~(layer3_outputs[642]) | (layer3_outputs[3063]);
    assign layer4_outputs[4402] = ~(layer3_outputs[3543]);
    assign layer4_outputs[4403] = ~(layer3_outputs[2175]) | (layer3_outputs[1848]);
    assign layer4_outputs[4404] = ~((layer3_outputs[4552]) ^ (layer3_outputs[1532]));
    assign layer4_outputs[4405] = ~(layer3_outputs[1813]);
    assign layer4_outputs[4406] = ~(layer3_outputs[2179]);
    assign layer4_outputs[4407] = ~(layer3_outputs[4478]) | (layer3_outputs[3714]);
    assign layer4_outputs[4408] = ~(layer3_outputs[4711]);
    assign layer4_outputs[4409] = 1'b1;
    assign layer4_outputs[4410] = layer3_outputs[3872];
    assign layer4_outputs[4411] = layer3_outputs[131];
    assign layer4_outputs[4412] = layer3_outputs[192];
    assign layer4_outputs[4413] = layer3_outputs[4831];
    assign layer4_outputs[4414] = (layer3_outputs[4872]) | (layer3_outputs[3073]);
    assign layer4_outputs[4415] = (layer3_outputs[4586]) & ~(layer3_outputs[72]);
    assign layer4_outputs[4416] = layer3_outputs[1907];
    assign layer4_outputs[4417] = (layer3_outputs[3444]) & ~(layer3_outputs[2043]);
    assign layer4_outputs[4418] = ~(layer3_outputs[139]) | (layer3_outputs[2755]);
    assign layer4_outputs[4419] = ~((layer3_outputs[4277]) & (layer3_outputs[1015]));
    assign layer4_outputs[4420] = (layer3_outputs[3787]) & (layer3_outputs[2692]);
    assign layer4_outputs[4421] = 1'b1;
    assign layer4_outputs[4422] = (layer3_outputs[2079]) & ~(layer3_outputs[214]);
    assign layer4_outputs[4423] = layer3_outputs[1730];
    assign layer4_outputs[4424] = (layer3_outputs[4064]) & ~(layer3_outputs[3651]);
    assign layer4_outputs[4425] = layer3_outputs[3145];
    assign layer4_outputs[4426] = (layer3_outputs[2022]) & (layer3_outputs[948]);
    assign layer4_outputs[4427] = (layer3_outputs[4216]) & ~(layer3_outputs[3107]);
    assign layer4_outputs[4428] = layer3_outputs[112];
    assign layer4_outputs[4429] = layer3_outputs[160];
    assign layer4_outputs[4430] = layer3_outputs[535];
    assign layer4_outputs[4431] = ~(layer3_outputs[4561]);
    assign layer4_outputs[4432] = ~((layer3_outputs[627]) & (layer3_outputs[3353]));
    assign layer4_outputs[4433] = 1'b0;
    assign layer4_outputs[4434] = (layer3_outputs[460]) & ~(layer3_outputs[2951]);
    assign layer4_outputs[4435] = (layer3_outputs[2538]) ^ (layer3_outputs[1748]);
    assign layer4_outputs[4436] = (layer3_outputs[695]) & ~(layer3_outputs[693]);
    assign layer4_outputs[4437] = (layer3_outputs[2907]) | (layer3_outputs[1550]);
    assign layer4_outputs[4438] = 1'b0;
    assign layer4_outputs[4439] = (layer3_outputs[2460]) | (layer3_outputs[755]);
    assign layer4_outputs[4440] = (layer3_outputs[4548]) ^ (layer3_outputs[874]);
    assign layer4_outputs[4441] = layer3_outputs[3280];
    assign layer4_outputs[4442] = ~((layer3_outputs[733]) & (layer3_outputs[129]));
    assign layer4_outputs[4443] = ~(layer3_outputs[1698]);
    assign layer4_outputs[4444] = ~(layer3_outputs[837]);
    assign layer4_outputs[4445] = (layer3_outputs[1629]) & ~(layer3_outputs[4281]);
    assign layer4_outputs[4446] = 1'b0;
    assign layer4_outputs[4447] = (layer3_outputs[2014]) | (layer3_outputs[893]);
    assign layer4_outputs[4448] = ~(layer3_outputs[3058]);
    assign layer4_outputs[4449] = layer3_outputs[888];
    assign layer4_outputs[4450] = ~(layer3_outputs[2771]);
    assign layer4_outputs[4451] = ~(layer3_outputs[3185]);
    assign layer4_outputs[4452] = ~(layer3_outputs[874]) | (layer3_outputs[632]);
    assign layer4_outputs[4453] = ~(layer3_outputs[1782]);
    assign layer4_outputs[4454] = (layer3_outputs[3997]) & ~(layer3_outputs[2864]);
    assign layer4_outputs[4455] = (layer3_outputs[4631]) & (layer3_outputs[3749]);
    assign layer4_outputs[4456] = (layer3_outputs[2246]) | (layer3_outputs[17]);
    assign layer4_outputs[4457] = ~(layer3_outputs[1149]);
    assign layer4_outputs[4458] = ~(layer3_outputs[3858]);
    assign layer4_outputs[4459] = layer3_outputs[3223];
    assign layer4_outputs[4460] = ~(layer3_outputs[414]);
    assign layer4_outputs[4461] = (layer3_outputs[973]) & ~(layer3_outputs[2327]);
    assign layer4_outputs[4462] = (layer3_outputs[347]) & (layer3_outputs[4187]);
    assign layer4_outputs[4463] = ~(layer3_outputs[4961]);
    assign layer4_outputs[4464] = ~(layer3_outputs[302]);
    assign layer4_outputs[4465] = (layer3_outputs[384]) & ~(layer3_outputs[2725]);
    assign layer4_outputs[4466] = ~(layer3_outputs[5089]);
    assign layer4_outputs[4467] = 1'b1;
    assign layer4_outputs[4468] = ~(layer3_outputs[1583]);
    assign layer4_outputs[4469] = ~(layer3_outputs[1904]) | (layer3_outputs[2475]);
    assign layer4_outputs[4470] = ~(layer3_outputs[3217]);
    assign layer4_outputs[4471] = (layer3_outputs[2015]) & ~(layer3_outputs[4872]);
    assign layer4_outputs[4472] = ~((layer3_outputs[8]) | (layer3_outputs[4207]));
    assign layer4_outputs[4473] = layer3_outputs[2585];
    assign layer4_outputs[4474] = ~((layer3_outputs[4092]) | (layer3_outputs[3177]));
    assign layer4_outputs[4475] = layer3_outputs[687];
    assign layer4_outputs[4476] = (layer3_outputs[1850]) & (layer3_outputs[1447]);
    assign layer4_outputs[4477] = 1'b0;
    assign layer4_outputs[4478] = layer3_outputs[3290];
    assign layer4_outputs[4479] = ~(layer3_outputs[1401]);
    assign layer4_outputs[4480] = ~((layer3_outputs[527]) & (layer3_outputs[835]));
    assign layer4_outputs[4481] = ~(layer3_outputs[5119]);
    assign layer4_outputs[4482] = layer3_outputs[693];
    assign layer4_outputs[4483] = layer3_outputs[628];
    assign layer4_outputs[4484] = 1'b0;
    assign layer4_outputs[4485] = ~(layer3_outputs[1019]);
    assign layer4_outputs[4486] = 1'b0;
    assign layer4_outputs[4487] = ~(layer3_outputs[3712]);
    assign layer4_outputs[4488] = (layer3_outputs[3023]) & (layer3_outputs[3050]);
    assign layer4_outputs[4489] = (layer3_outputs[2777]) & ~(layer3_outputs[2629]);
    assign layer4_outputs[4490] = layer3_outputs[2749];
    assign layer4_outputs[4491] = ~(layer3_outputs[1657]);
    assign layer4_outputs[4492] = (layer3_outputs[3529]) ^ (layer3_outputs[48]);
    assign layer4_outputs[4493] = (layer3_outputs[2113]) | (layer3_outputs[3303]);
    assign layer4_outputs[4494] = (layer3_outputs[3535]) | (layer3_outputs[1050]);
    assign layer4_outputs[4495] = ~(layer3_outputs[4838]) | (layer3_outputs[1978]);
    assign layer4_outputs[4496] = layer3_outputs[4268];
    assign layer4_outputs[4497] = ~(layer3_outputs[2790]);
    assign layer4_outputs[4498] = layer3_outputs[2413];
    assign layer4_outputs[4499] = ~(layer3_outputs[2943]) | (layer3_outputs[2035]);
    assign layer4_outputs[4500] = layer3_outputs[4027];
    assign layer4_outputs[4501] = ~((layer3_outputs[2010]) | (layer3_outputs[2506]));
    assign layer4_outputs[4502] = (layer3_outputs[2791]) & ~(layer3_outputs[4619]);
    assign layer4_outputs[4503] = layer3_outputs[2370];
    assign layer4_outputs[4504] = layer3_outputs[4288];
    assign layer4_outputs[4505] = 1'b0;
    assign layer4_outputs[4506] = (layer3_outputs[3291]) | (layer3_outputs[1603]);
    assign layer4_outputs[4507] = (layer3_outputs[3404]) ^ (layer3_outputs[1926]);
    assign layer4_outputs[4508] = ~((layer3_outputs[4865]) | (layer3_outputs[3075]));
    assign layer4_outputs[4509] = 1'b0;
    assign layer4_outputs[4510] = 1'b0;
    assign layer4_outputs[4511] = ~(layer3_outputs[871]);
    assign layer4_outputs[4512] = layer3_outputs[1509];
    assign layer4_outputs[4513] = ~(layer3_outputs[684]);
    assign layer4_outputs[4514] = ~(layer3_outputs[3673]);
    assign layer4_outputs[4515] = layer3_outputs[3150];
    assign layer4_outputs[4516] = (layer3_outputs[1561]) ^ (layer3_outputs[1296]);
    assign layer4_outputs[4517] = ~(layer3_outputs[1950]);
    assign layer4_outputs[4518] = (layer3_outputs[3604]) & ~(layer3_outputs[4241]);
    assign layer4_outputs[4519] = ~(layer3_outputs[4430]);
    assign layer4_outputs[4520] = ~(layer3_outputs[2501]);
    assign layer4_outputs[4521] = (layer3_outputs[4047]) & (layer3_outputs[869]);
    assign layer4_outputs[4522] = (layer3_outputs[4471]) ^ (layer3_outputs[1590]);
    assign layer4_outputs[4523] = ~(layer3_outputs[2539]);
    assign layer4_outputs[4524] = ~((layer3_outputs[4080]) & (layer3_outputs[2599]));
    assign layer4_outputs[4525] = ~(layer3_outputs[3833]);
    assign layer4_outputs[4526] = ~((layer3_outputs[2626]) | (layer3_outputs[1346]));
    assign layer4_outputs[4527] = ~(layer3_outputs[3530]);
    assign layer4_outputs[4528] = layer3_outputs[1056];
    assign layer4_outputs[4529] = ~(layer3_outputs[3157]) | (layer3_outputs[4456]);
    assign layer4_outputs[4530] = (layer3_outputs[3575]) & ~(layer3_outputs[1977]);
    assign layer4_outputs[4531] = 1'b0;
    assign layer4_outputs[4532] = (layer3_outputs[1268]) & (layer3_outputs[2233]);
    assign layer4_outputs[4533] = ~((layer3_outputs[1282]) | (layer3_outputs[1224]));
    assign layer4_outputs[4534] = (layer3_outputs[1711]) & ~(layer3_outputs[2869]);
    assign layer4_outputs[4535] = ~(layer3_outputs[124]);
    assign layer4_outputs[4536] = (layer3_outputs[3401]) & ~(layer3_outputs[4805]);
    assign layer4_outputs[4537] = ~(layer3_outputs[4166]);
    assign layer4_outputs[4538] = (layer3_outputs[1399]) & ~(layer3_outputs[3599]);
    assign layer4_outputs[4539] = layer3_outputs[1957];
    assign layer4_outputs[4540] = 1'b1;
    assign layer4_outputs[4541] = layer3_outputs[4279];
    assign layer4_outputs[4542] = ~((layer3_outputs[4648]) | (layer3_outputs[3215]));
    assign layer4_outputs[4543] = ~(layer3_outputs[4756]);
    assign layer4_outputs[4544] = layer3_outputs[2923];
    assign layer4_outputs[4545] = ~(layer3_outputs[1719]);
    assign layer4_outputs[4546] = ~(layer3_outputs[2434]);
    assign layer4_outputs[4547] = ~(layer3_outputs[3448]) | (layer3_outputs[1217]);
    assign layer4_outputs[4548] = ~((layer3_outputs[940]) | (layer3_outputs[4433]));
    assign layer4_outputs[4549] = ~(layer3_outputs[3033]);
    assign layer4_outputs[4550] = ~((layer3_outputs[3644]) & (layer3_outputs[4397]));
    assign layer4_outputs[4551] = (layer3_outputs[2041]) & ~(layer3_outputs[122]);
    assign layer4_outputs[4552] = ~(layer3_outputs[5096]) | (layer3_outputs[851]);
    assign layer4_outputs[4553] = ~((layer3_outputs[3902]) & (layer3_outputs[2852]));
    assign layer4_outputs[4554] = 1'b0;
    assign layer4_outputs[4555] = (layer3_outputs[4138]) ^ (layer3_outputs[1978]);
    assign layer4_outputs[4556] = ~(layer3_outputs[4617]);
    assign layer4_outputs[4557] = ~(layer3_outputs[1443]) | (layer3_outputs[2682]);
    assign layer4_outputs[4558] = ~(layer3_outputs[4981]);
    assign layer4_outputs[4559] = (layer3_outputs[1021]) | (layer3_outputs[1267]);
    assign layer4_outputs[4560] = ~(layer3_outputs[4644]);
    assign layer4_outputs[4561] = (layer3_outputs[3388]) ^ (layer3_outputs[5084]);
    assign layer4_outputs[4562] = (layer3_outputs[659]) & ~(layer3_outputs[4772]);
    assign layer4_outputs[4563] = (layer3_outputs[1879]) | (layer3_outputs[2835]);
    assign layer4_outputs[4564] = (layer3_outputs[2091]) & ~(layer3_outputs[2766]);
    assign layer4_outputs[4565] = ~(layer3_outputs[3321]);
    assign layer4_outputs[4566] = 1'b0;
    assign layer4_outputs[4567] = (layer3_outputs[2815]) & ~(layer3_outputs[3744]);
    assign layer4_outputs[4568] = layer3_outputs[1388];
    assign layer4_outputs[4569] = layer3_outputs[3534];
    assign layer4_outputs[4570] = layer3_outputs[2249];
    assign layer4_outputs[4571] = ~(layer3_outputs[207]) | (layer3_outputs[2398]);
    assign layer4_outputs[4572] = ~((layer3_outputs[3420]) | (layer3_outputs[4373]));
    assign layer4_outputs[4573] = (layer3_outputs[4897]) & (layer3_outputs[4561]);
    assign layer4_outputs[4574] = ~(layer3_outputs[119]);
    assign layer4_outputs[4575] = 1'b1;
    assign layer4_outputs[4576] = (layer3_outputs[3838]) ^ (layer3_outputs[4550]);
    assign layer4_outputs[4577] = 1'b0;
    assign layer4_outputs[4578] = ~(layer3_outputs[530]);
    assign layer4_outputs[4579] = ~((layer3_outputs[4665]) ^ (layer3_outputs[2501]));
    assign layer4_outputs[4580] = (layer3_outputs[7]) | (layer3_outputs[2360]);
    assign layer4_outputs[4581] = layer3_outputs[4029];
    assign layer4_outputs[4582] = (layer3_outputs[3505]) & ~(layer3_outputs[371]);
    assign layer4_outputs[4583] = layer3_outputs[4248];
    assign layer4_outputs[4584] = ~(layer3_outputs[2292]) | (layer3_outputs[1137]);
    assign layer4_outputs[4585] = layer3_outputs[1650];
    assign layer4_outputs[4586] = (layer3_outputs[1576]) & (layer3_outputs[3317]);
    assign layer4_outputs[4587] = ~(layer3_outputs[3672]) | (layer3_outputs[4331]);
    assign layer4_outputs[4588] = ~(layer3_outputs[1718]) | (layer3_outputs[2373]);
    assign layer4_outputs[4589] = ~(layer3_outputs[605]);
    assign layer4_outputs[4590] = ~(layer3_outputs[450]);
    assign layer4_outputs[4591] = layer3_outputs[1112];
    assign layer4_outputs[4592] = (layer3_outputs[4185]) & ~(layer3_outputs[1288]);
    assign layer4_outputs[4593] = layer3_outputs[2934];
    assign layer4_outputs[4594] = layer3_outputs[2473];
    assign layer4_outputs[4595] = (layer3_outputs[3579]) | (layer3_outputs[1761]);
    assign layer4_outputs[4596] = 1'b0;
    assign layer4_outputs[4597] = layer3_outputs[3530];
    assign layer4_outputs[4598] = ~(layer3_outputs[3106]);
    assign layer4_outputs[4599] = ~(layer3_outputs[792]);
    assign layer4_outputs[4600] = ~(layer3_outputs[1571]);
    assign layer4_outputs[4601] = layer3_outputs[3995];
    assign layer4_outputs[4602] = ~(layer3_outputs[635]) | (layer3_outputs[1640]);
    assign layer4_outputs[4603] = 1'b1;
    assign layer4_outputs[4604] = layer3_outputs[2700];
    assign layer4_outputs[4605] = ~(layer3_outputs[3974]) | (layer3_outputs[3589]);
    assign layer4_outputs[4606] = (layer3_outputs[3648]) & ~(layer3_outputs[2201]);
    assign layer4_outputs[4607] = ~((layer3_outputs[3336]) & (layer3_outputs[2080]));
    assign layer4_outputs[4608] = ~(layer3_outputs[3673]) | (layer3_outputs[4108]);
    assign layer4_outputs[4609] = (layer3_outputs[2591]) & ~(layer3_outputs[4976]);
    assign layer4_outputs[4610] = ~(layer3_outputs[1938]);
    assign layer4_outputs[4611] = ~(layer3_outputs[239]) | (layer3_outputs[1363]);
    assign layer4_outputs[4612] = ~(layer3_outputs[3104]) | (layer3_outputs[570]);
    assign layer4_outputs[4613] = layer3_outputs[2585];
    assign layer4_outputs[4614] = ~(layer3_outputs[166]);
    assign layer4_outputs[4615] = (layer3_outputs[3123]) & (layer3_outputs[4820]);
    assign layer4_outputs[4616] = (layer3_outputs[2248]) & (layer3_outputs[2581]);
    assign layer4_outputs[4617] = layer3_outputs[3592];
    assign layer4_outputs[4618] = ~((layer3_outputs[889]) & (layer3_outputs[3926]));
    assign layer4_outputs[4619] = (layer3_outputs[4708]) & ~(layer3_outputs[4932]);
    assign layer4_outputs[4620] = 1'b1;
    assign layer4_outputs[4621] = ~(layer3_outputs[2528]) | (layer3_outputs[2306]);
    assign layer4_outputs[4622] = (layer3_outputs[5080]) & ~(layer3_outputs[1715]);
    assign layer4_outputs[4623] = layer3_outputs[791];
    assign layer4_outputs[4624] = (layer3_outputs[2003]) & ~(layer3_outputs[1800]);
    assign layer4_outputs[4625] = (layer3_outputs[1628]) | (layer3_outputs[1130]);
    assign layer4_outputs[4626] = layer3_outputs[3001];
    assign layer4_outputs[4627] = layer3_outputs[1941];
    assign layer4_outputs[4628] = ~(layer3_outputs[3360]);
    assign layer4_outputs[4629] = ~((layer3_outputs[4590]) | (layer3_outputs[4864]));
    assign layer4_outputs[4630] = layer3_outputs[4510];
    assign layer4_outputs[4631] = ~((layer3_outputs[1471]) | (layer3_outputs[1311]));
    assign layer4_outputs[4632] = ~((layer3_outputs[4929]) & (layer3_outputs[1037]));
    assign layer4_outputs[4633] = (layer3_outputs[2982]) & ~(layer3_outputs[756]);
    assign layer4_outputs[4634] = layer3_outputs[4991];
    assign layer4_outputs[4635] = 1'b0;
    assign layer4_outputs[4636] = (layer3_outputs[4348]) & (layer3_outputs[2976]);
    assign layer4_outputs[4637] = 1'b0;
    assign layer4_outputs[4638] = ~((layer3_outputs[3284]) ^ (layer3_outputs[169]));
    assign layer4_outputs[4639] = ~(layer3_outputs[409]) | (layer3_outputs[2992]);
    assign layer4_outputs[4640] = layer3_outputs[4617];
    assign layer4_outputs[4641] = (layer3_outputs[1844]) | (layer3_outputs[4407]);
    assign layer4_outputs[4642] = ~(layer3_outputs[3257]);
    assign layer4_outputs[4643] = 1'b1;
    assign layer4_outputs[4644] = ~(layer3_outputs[4207]) | (layer3_outputs[2122]);
    assign layer4_outputs[4645] = (layer3_outputs[1034]) | (layer3_outputs[3371]);
    assign layer4_outputs[4646] = ~(layer3_outputs[4632]) | (layer3_outputs[4385]);
    assign layer4_outputs[4647] = ~(layer3_outputs[376]) | (layer3_outputs[3703]);
    assign layer4_outputs[4648] = layer3_outputs[3629];
    assign layer4_outputs[4649] = ~((layer3_outputs[3298]) & (layer3_outputs[4638]));
    assign layer4_outputs[4650] = ~(layer3_outputs[621]);
    assign layer4_outputs[4651] = (layer3_outputs[3902]) | (layer3_outputs[2221]);
    assign layer4_outputs[4652] = 1'b1;
    assign layer4_outputs[4653] = ~(layer3_outputs[1497]) | (layer3_outputs[903]);
    assign layer4_outputs[4654] = (layer3_outputs[241]) & ~(layer3_outputs[575]);
    assign layer4_outputs[4655] = ~(layer3_outputs[2985]) | (layer3_outputs[1313]);
    assign layer4_outputs[4656] = layer3_outputs[4501];
    assign layer4_outputs[4657] = ~(layer3_outputs[942]);
    assign layer4_outputs[4658] = ~((layer3_outputs[1028]) | (layer3_outputs[845]));
    assign layer4_outputs[4659] = 1'b0;
    assign layer4_outputs[4660] = ~(layer3_outputs[2569]);
    assign layer4_outputs[4661] = ~(layer3_outputs[1245]) | (layer3_outputs[1791]);
    assign layer4_outputs[4662] = ~(layer3_outputs[3947]);
    assign layer4_outputs[4663] = layer3_outputs[1208];
    assign layer4_outputs[4664] = ~(layer3_outputs[2936]) | (layer3_outputs[1249]);
    assign layer4_outputs[4665] = layer3_outputs[3854];
    assign layer4_outputs[4666] = layer3_outputs[672];
    assign layer4_outputs[4667] = ~((layer3_outputs[1109]) & (layer3_outputs[484]));
    assign layer4_outputs[4668] = ~(layer3_outputs[132]) | (layer3_outputs[2092]);
    assign layer4_outputs[4669] = (layer3_outputs[1088]) ^ (layer3_outputs[3697]);
    assign layer4_outputs[4670] = layer3_outputs[2959];
    assign layer4_outputs[4671] = (layer3_outputs[1952]) & ~(layer3_outputs[3794]);
    assign layer4_outputs[4672] = (layer3_outputs[2765]) & ~(layer3_outputs[1945]);
    assign layer4_outputs[4673] = ~(layer3_outputs[1654]);
    assign layer4_outputs[4674] = layer3_outputs[2374];
    assign layer4_outputs[4675] = (layer3_outputs[1979]) | (layer3_outputs[2305]);
    assign layer4_outputs[4676] = ~(layer3_outputs[2254]) | (layer3_outputs[3901]);
    assign layer4_outputs[4677] = ~(layer3_outputs[3133]);
    assign layer4_outputs[4678] = (layer3_outputs[3526]) & ~(layer3_outputs[27]);
    assign layer4_outputs[4679] = (layer3_outputs[475]) ^ (layer3_outputs[1727]);
    assign layer4_outputs[4680] = layer3_outputs[4780];
    assign layer4_outputs[4681] = ~((layer3_outputs[955]) ^ (layer3_outputs[3785]));
    assign layer4_outputs[4682] = 1'b1;
    assign layer4_outputs[4683] = (layer3_outputs[3452]) & ~(layer3_outputs[3069]);
    assign layer4_outputs[4684] = ~(layer3_outputs[1536]) | (layer3_outputs[2314]);
    assign layer4_outputs[4685] = ~(layer3_outputs[3591]);
    assign layer4_outputs[4686] = ~(layer3_outputs[1917]);
    assign layer4_outputs[4687] = layer3_outputs[1485];
    assign layer4_outputs[4688] = layer3_outputs[3238];
    assign layer4_outputs[4689] = ~(layer3_outputs[2354]);
    assign layer4_outputs[4690] = (layer3_outputs[4615]) & ~(layer3_outputs[2109]);
    assign layer4_outputs[4691] = ~(layer3_outputs[1397]);
    assign layer4_outputs[4692] = layer3_outputs[1858];
    assign layer4_outputs[4693] = ~((layer3_outputs[3772]) & (layer3_outputs[3696]));
    assign layer4_outputs[4694] = (layer3_outputs[1302]) | (layer3_outputs[1640]);
    assign layer4_outputs[4695] = (layer3_outputs[3398]) ^ (layer3_outputs[2044]);
    assign layer4_outputs[4696] = ~((layer3_outputs[3208]) | (layer3_outputs[419]));
    assign layer4_outputs[4697] = layer3_outputs[4976];
    assign layer4_outputs[4698] = (layer3_outputs[3924]) & (layer3_outputs[1195]);
    assign layer4_outputs[4699] = layer3_outputs[3414];
    assign layer4_outputs[4700] = (layer3_outputs[2254]) & ~(layer3_outputs[1232]);
    assign layer4_outputs[4701] = ~(layer3_outputs[253]);
    assign layer4_outputs[4702] = (layer3_outputs[3602]) & (layer3_outputs[2461]);
    assign layer4_outputs[4703] = ~(layer3_outputs[1441]);
    assign layer4_outputs[4704] = ~(layer3_outputs[4051]);
    assign layer4_outputs[4705] = ~(layer3_outputs[3908]) | (layer3_outputs[1222]);
    assign layer4_outputs[4706] = (layer3_outputs[4398]) & ~(layer3_outputs[1324]);
    assign layer4_outputs[4707] = layer3_outputs[5112];
    assign layer4_outputs[4708] = ~(layer3_outputs[2219]);
    assign layer4_outputs[4709] = (layer3_outputs[2296]) & ~(layer3_outputs[2207]);
    assign layer4_outputs[4710] = ~((layer3_outputs[4888]) | (layer3_outputs[2243]));
    assign layer4_outputs[4711] = ~(layer3_outputs[183]);
    assign layer4_outputs[4712] = (layer3_outputs[1366]) | (layer3_outputs[3588]);
    assign layer4_outputs[4713] = ~((layer3_outputs[5022]) & (layer3_outputs[4788]));
    assign layer4_outputs[4714] = 1'b1;
    assign layer4_outputs[4715] = ~(layer3_outputs[1315]);
    assign layer4_outputs[4716] = ~((layer3_outputs[4142]) & (layer3_outputs[4682]));
    assign layer4_outputs[4717] = (layer3_outputs[1595]) & (layer3_outputs[4088]);
    assign layer4_outputs[4718] = (layer3_outputs[1179]) & ~(layer3_outputs[2764]);
    assign layer4_outputs[4719] = ~((layer3_outputs[2406]) | (layer3_outputs[2614]));
    assign layer4_outputs[4720] = ~((layer3_outputs[3294]) | (layer3_outputs[2483]));
    assign layer4_outputs[4721] = ~(layer3_outputs[3171]) | (layer3_outputs[93]);
    assign layer4_outputs[4722] = ~((layer3_outputs[5000]) & (layer3_outputs[2036]));
    assign layer4_outputs[4723] = layer3_outputs[4183];
    assign layer4_outputs[4724] = ~((layer3_outputs[3603]) ^ (layer3_outputs[855]));
    assign layer4_outputs[4725] = ~(layer3_outputs[2247]);
    assign layer4_outputs[4726] = ~(layer3_outputs[1572]);
    assign layer4_outputs[4727] = (layer3_outputs[485]) & ~(layer3_outputs[3184]);
    assign layer4_outputs[4728] = (layer3_outputs[2689]) ^ (layer3_outputs[2935]);
    assign layer4_outputs[4729] = ~(layer3_outputs[4571]);
    assign layer4_outputs[4730] = layer3_outputs[3510];
    assign layer4_outputs[4731] = (layer3_outputs[20]) | (layer3_outputs[1634]);
    assign layer4_outputs[4732] = (layer3_outputs[4498]) & (layer3_outputs[2362]);
    assign layer4_outputs[4733] = ~(layer3_outputs[4457]);
    assign layer4_outputs[4734] = ~(layer3_outputs[4928]);
    assign layer4_outputs[4735] = (layer3_outputs[2880]) & (layer3_outputs[2981]);
    assign layer4_outputs[4736] = layer3_outputs[1368];
    assign layer4_outputs[4737] = layer3_outputs[717];
    assign layer4_outputs[4738] = 1'b0;
    assign layer4_outputs[4739] = layer3_outputs[4807];
    assign layer4_outputs[4740] = layer3_outputs[4973];
    assign layer4_outputs[4741] = ~(layer3_outputs[4011]);
    assign layer4_outputs[4742] = ~((layer3_outputs[603]) & (layer3_outputs[2227]));
    assign layer4_outputs[4743] = (layer3_outputs[4563]) & ~(layer3_outputs[1018]);
    assign layer4_outputs[4744] = 1'b1;
    assign layer4_outputs[4745] = layer3_outputs[4303];
    assign layer4_outputs[4746] = ~((layer3_outputs[1871]) | (layer3_outputs[1087]));
    assign layer4_outputs[4747] = (layer3_outputs[2641]) | (layer3_outputs[1621]);
    assign layer4_outputs[4748] = ~(layer3_outputs[1104]);
    assign layer4_outputs[4749] = ~(layer3_outputs[4031]);
    assign layer4_outputs[4750] = (layer3_outputs[219]) ^ (layer3_outputs[3596]);
    assign layer4_outputs[4751] = ~((layer3_outputs[3155]) ^ (layer3_outputs[87]));
    assign layer4_outputs[4752] = (layer3_outputs[1548]) | (layer3_outputs[4907]);
    assign layer4_outputs[4753] = ~(layer3_outputs[765]);
    assign layer4_outputs[4754] = ~(layer3_outputs[290]);
    assign layer4_outputs[4755] = (layer3_outputs[3520]) & ~(layer3_outputs[1178]);
    assign layer4_outputs[4756] = ~(layer3_outputs[2850]);
    assign layer4_outputs[4757] = layer3_outputs[3470];
    assign layer4_outputs[4758] = ~((layer3_outputs[1221]) ^ (layer3_outputs[3299]));
    assign layer4_outputs[4759] = layer3_outputs[2810];
    assign layer4_outputs[4760] = ~((layer3_outputs[1166]) | (layer3_outputs[197]));
    assign layer4_outputs[4761] = (layer3_outputs[4155]) & (layer3_outputs[986]);
    assign layer4_outputs[4762] = ~(layer3_outputs[3301]);
    assign layer4_outputs[4763] = ~((layer3_outputs[3496]) & (layer3_outputs[3677]));
    assign layer4_outputs[4764] = ~(layer3_outputs[3411]);
    assign layer4_outputs[4765] = ~(layer3_outputs[1815]);
    assign layer4_outputs[4766] = (layer3_outputs[135]) | (layer3_outputs[2182]);
    assign layer4_outputs[4767] = ~(layer3_outputs[2730]);
    assign layer4_outputs[4768] = ~(layer3_outputs[1251]) | (layer3_outputs[1855]);
    assign layer4_outputs[4769] = layer3_outputs[4310];
    assign layer4_outputs[4770] = (layer3_outputs[1982]) & ~(layer3_outputs[731]);
    assign layer4_outputs[4771] = ~(layer3_outputs[1667]);
    assign layer4_outputs[4772] = (layer3_outputs[4276]) ^ (layer3_outputs[4915]);
    assign layer4_outputs[4773] = layer3_outputs[770];
    assign layer4_outputs[4774] = layer3_outputs[402];
    assign layer4_outputs[4775] = ~(layer3_outputs[4185]);
    assign layer4_outputs[4776] = layer3_outputs[2397];
    assign layer4_outputs[4777] = ~((layer3_outputs[1511]) & (layer3_outputs[2502]));
    assign layer4_outputs[4778] = ~((layer3_outputs[930]) ^ (layer3_outputs[4885]));
    assign layer4_outputs[4779] = layer3_outputs[1824];
    assign layer4_outputs[4780] = layer3_outputs[3390];
    assign layer4_outputs[4781] = layer3_outputs[4084];
    assign layer4_outputs[4782] = ~(layer3_outputs[203]);
    assign layer4_outputs[4783] = ~(layer3_outputs[5015]) | (layer3_outputs[4559]);
    assign layer4_outputs[4784] = ~((layer3_outputs[3041]) ^ (layer3_outputs[521]));
    assign layer4_outputs[4785] = layer3_outputs[2890];
    assign layer4_outputs[4786] = layer3_outputs[2134];
    assign layer4_outputs[4787] = ~(layer3_outputs[4829]) | (layer3_outputs[2066]);
    assign layer4_outputs[4788] = ~(layer3_outputs[1167]);
    assign layer4_outputs[4789] = (layer3_outputs[2021]) ^ (layer3_outputs[2876]);
    assign layer4_outputs[4790] = (layer3_outputs[2145]) & ~(layer3_outputs[4338]);
    assign layer4_outputs[4791] = ~((layer3_outputs[1648]) & (layer3_outputs[4864]));
    assign layer4_outputs[4792] = (layer3_outputs[4162]) & ~(layer3_outputs[3193]);
    assign layer4_outputs[4793] = (layer3_outputs[1013]) & ~(layer3_outputs[875]);
    assign layer4_outputs[4794] = (layer3_outputs[3878]) & (layer3_outputs[232]);
    assign layer4_outputs[4795] = ~(layer3_outputs[3485]);
    assign layer4_outputs[4796] = ~((layer3_outputs[3232]) | (layer3_outputs[3965]));
    assign layer4_outputs[4797] = layer3_outputs[334];
    assign layer4_outputs[4798] = (layer3_outputs[4612]) ^ (layer3_outputs[1843]);
    assign layer4_outputs[4799] = ~(layer3_outputs[1299]);
    assign layer4_outputs[4800] = ~(layer3_outputs[2294]);
    assign layer4_outputs[4801] = ~(layer3_outputs[1017]);
    assign layer4_outputs[4802] = layer3_outputs[4714];
    assign layer4_outputs[4803] = (layer3_outputs[790]) ^ (layer3_outputs[4637]);
    assign layer4_outputs[4804] = (layer3_outputs[2335]) & (layer3_outputs[261]);
    assign layer4_outputs[4805] = layer3_outputs[1375];
    assign layer4_outputs[4806] = (layer3_outputs[3216]) & ~(layer3_outputs[616]);
    assign layer4_outputs[4807] = layer3_outputs[436];
    assign layer4_outputs[4808] = layer3_outputs[3161];
    assign layer4_outputs[4809] = ~((layer3_outputs[1964]) ^ (layer3_outputs[112]));
    assign layer4_outputs[4810] = ~(layer3_outputs[1339]);
    assign layer4_outputs[4811] = ~((layer3_outputs[1465]) | (layer3_outputs[990]));
    assign layer4_outputs[4812] = (layer3_outputs[3606]) & ~(layer3_outputs[3345]);
    assign layer4_outputs[4813] = layer3_outputs[439];
    assign layer4_outputs[4814] = ~(layer3_outputs[1429]);
    assign layer4_outputs[4815] = layer3_outputs[1553];
    assign layer4_outputs[4816] = ~((layer3_outputs[2277]) | (layer3_outputs[3328]));
    assign layer4_outputs[4817] = layer3_outputs[4884];
    assign layer4_outputs[4818] = ~(layer3_outputs[4521]);
    assign layer4_outputs[4819] = (layer3_outputs[4117]) & ~(layer3_outputs[2059]);
    assign layer4_outputs[4820] = ~(layer3_outputs[1118]);
    assign layer4_outputs[4821] = layer3_outputs[4151];
    assign layer4_outputs[4822] = ~(layer3_outputs[4112]);
    assign layer4_outputs[4823] = (layer3_outputs[2390]) ^ (layer3_outputs[703]);
    assign layer4_outputs[4824] = (layer3_outputs[4335]) ^ (layer3_outputs[3790]);
    assign layer4_outputs[4825] = ~(layer3_outputs[1618]);
    assign layer4_outputs[4826] = ~(layer3_outputs[1768]);
    assign layer4_outputs[4827] = (layer3_outputs[1165]) ^ (layer3_outputs[1285]);
    assign layer4_outputs[4828] = (layer3_outputs[1825]) | (layer3_outputs[1741]);
    assign layer4_outputs[4829] = ~((layer3_outputs[2774]) | (layer3_outputs[4637]));
    assign layer4_outputs[4830] = (layer3_outputs[1211]) & ~(layer3_outputs[1003]);
    assign layer4_outputs[4831] = ~((layer3_outputs[738]) ^ (layer3_outputs[1572]));
    assign layer4_outputs[4832] = (layer3_outputs[329]) | (layer3_outputs[386]);
    assign layer4_outputs[4833] = layer3_outputs[2802];
    assign layer4_outputs[4834] = layer3_outputs[5079];
    assign layer4_outputs[4835] = ~(layer3_outputs[3056]) | (layer3_outputs[4256]);
    assign layer4_outputs[4836] = ~(layer3_outputs[4720]);
    assign layer4_outputs[4837] = layer3_outputs[3146];
    assign layer4_outputs[4838] = ~(layer3_outputs[5011]) | (layer3_outputs[4752]);
    assign layer4_outputs[4839] = ~(layer3_outputs[3018]) | (layer3_outputs[3258]);
    assign layer4_outputs[4840] = (layer3_outputs[2293]) & ~(layer3_outputs[2652]);
    assign layer4_outputs[4841] = ~(layer3_outputs[2569]);
    assign layer4_outputs[4842] = ~((layer3_outputs[3049]) & (layer3_outputs[2911]));
    assign layer4_outputs[4843] = layer3_outputs[3713];
    assign layer4_outputs[4844] = ~(layer3_outputs[4272]);
    assign layer4_outputs[4845] = layer3_outputs[2780];
    assign layer4_outputs[4846] = (layer3_outputs[533]) | (layer3_outputs[1548]);
    assign layer4_outputs[4847] = (layer3_outputs[1772]) & (layer3_outputs[1583]);
    assign layer4_outputs[4848] = layer3_outputs[791];
    assign layer4_outputs[4849] = 1'b1;
    assign layer4_outputs[4850] = layer3_outputs[873];
    assign layer4_outputs[4851] = ~(layer3_outputs[3595]) | (layer3_outputs[1179]);
    assign layer4_outputs[4852] = (layer3_outputs[4860]) | (layer3_outputs[2001]);
    assign layer4_outputs[4853] = ~(layer3_outputs[46]);
    assign layer4_outputs[4854] = ~(layer3_outputs[3959]) | (layer3_outputs[3565]);
    assign layer4_outputs[4855] = layer3_outputs[1233];
    assign layer4_outputs[4856] = ~(layer3_outputs[439]) | (layer3_outputs[4260]);
    assign layer4_outputs[4857] = (layer3_outputs[982]) & ~(layer3_outputs[3071]);
    assign layer4_outputs[4858] = (layer3_outputs[3162]) & ~(layer3_outputs[1030]);
    assign layer4_outputs[4859] = ~(layer3_outputs[3431]);
    assign layer4_outputs[4860] = layer3_outputs[2008];
    assign layer4_outputs[4861] = (layer3_outputs[4149]) & ~(layer3_outputs[1549]);
    assign layer4_outputs[4862] = (layer3_outputs[4415]) | (layer3_outputs[2312]);
    assign layer4_outputs[4863] = ~(layer3_outputs[3911]);
    assign layer4_outputs[4864] = layer3_outputs[4346];
    assign layer4_outputs[4865] = layer3_outputs[1352];
    assign layer4_outputs[4866] = layer3_outputs[3502];
    assign layer4_outputs[4867] = ~(layer3_outputs[1633]);
    assign layer4_outputs[4868] = ~(layer3_outputs[3607]);
    assign layer4_outputs[4869] = layer3_outputs[4244];
    assign layer4_outputs[4870] = (layer3_outputs[4895]) & ~(layer3_outputs[3683]);
    assign layer4_outputs[4871] = layer3_outputs[2909];
    assign layer4_outputs[4872] = 1'b1;
    assign layer4_outputs[4873] = ~((layer3_outputs[3413]) | (layer3_outputs[2881]));
    assign layer4_outputs[4874] = layer3_outputs[2685];
    assign layer4_outputs[4875] = ~(layer3_outputs[1634]);
    assign layer4_outputs[4876] = (layer3_outputs[4001]) | (layer3_outputs[1277]);
    assign layer4_outputs[4877] = ~(layer3_outputs[876]);
    assign layer4_outputs[4878] = ~(layer3_outputs[483]) | (layer3_outputs[372]);
    assign layer4_outputs[4879] = ~(layer3_outputs[667]);
    assign layer4_outputs[4880] = (layer3_outputs[1296]) & ~(layer3_outputs[4760]);
    assign layer4_outputs[4881] = layer3_outputs[4257];
    assign layer4_outputs[4882] = ~((layer3_outputs[4833]) | (layer3_outputs[617]));
    assign layer4_outputs[4883] = (layer3_outputs[3231]) & (layer3_outputs[2462]);
    assign layer4_outputs[4884] = ~(layer3_outputs[562]);
    assign layer4_outputs[4885] = ~(layer3_outputs[1286]);
    assign layer4_outputs[4886] = ~(layer3_outputs[2188]) | (layer3_outputs[2378]);
    assign layer4_outputs[4887] = ~(layer3_outputs[1261]);
    assign layer4_outputs[4888] = (layer3_outputs[3880]) | (layer3_outputs[4925]);
    assign layer4_outputs[4889] = ~((layer3_outputs[1413]) | (layer3_outputs[3615]));
    assign layer4_outputs[4890] = ~(layer3_outputs[2131]);
    assign layer4_outputs[4891] = layer3_outputs[3559];
    assign layer4_outputs[4892] = (layer3_outputs[192]) & (layer3_outputs[379]);
    assign layer4_outputs[4893] = ~(layer3_outputs[3833]) | (layer3_outputs[657]);
    assign layer4_outputs[4894] = ~((layer3_outputs[3605]) & (layer3_outputs[586]));
    assign layer4_outputs[4895] = layer3_outputs[4557];
    assign layer4_outputs[4896] = ~(layer3_outputs[1818]);
    assign layer4_outputs[4897] = layer3_outputs[2079];
    assign layer4_outputs[4898] = layer3_outputs[3578];
    assign layer4_outputs[4899] = (layer3_outputs[715]) ^ (layer3_outputs[1732]);
    assign layer4_outputs[4900] = ~(layer3_outputs[3979]) | (layer3_outputs[3880]);
    assign layer4_outputs[4901] = (layer3_outputs[3500]) & ~(layer3_outputs[2598]);
    assign layer4_outputs[4902] = (layer3_outputs[589]) & ~(layer3_outputs[3956]);
    assign layer4_outputs[4903] = layer3_outputs[3747];
    assign layer4_outputs[4904] = (layer3_outputs[3441]) & ~(layer3_outputs[1923]);
    assign layer4_outputs[4905] = layer3_outputs[768];
    assign layer4_outputs[4906] = ~(layer3_outputs[1418]);
    assign layer4_outputs[4907] = ~(layer3_outputs[2630]) | (layer3_outputs[2057]);
    assign layer4_outputs[4908] = (layer3_outputs[1394]) & ~(layer3_outputs[3211]);
    assign layer4_outputs[4909] = (layer3_outputs[743]) & ~(layer3_outputs[4690]);
    assign layer4_outputs[4910] = 1'b0;
    assign layer4_outputs[4911] = ~(layer3_outputs[5113]) | (layer3_outputs[3067]);
    assign layer4_outputs[4912] = ~((layer3_outputs[831]) & (layer3_outputs[3141]));
    assign layer4_outputs[4913] = (layer3_outputs[756]) & (layer3_outputs[670]);
    assign layer4_outputs[4914] = layer3_outputs[83];
    assign layer4_outputs[4915] = ~(layer3_outputs[3826]);
    assign layer4_outputs[4916] = ~((layer3_outputs[995]) & (layer3_outputs[3823]));
    assign layer4_outputs[4917] = ~(layer3_outputs[2037]) | (layer3_outputs[211]);
    assign layer4_outputs[4918] = (layer3_outputs[1013]) & ~(layer3_outputs[3743]);
    assign layer4_outputs[4919] = layer3_outputs[1997];
    assign layer4_outputs[4920] = (layer3_outputs[3764]) & ~(layer3_outputs[3895]);
    assign layer4_outputs[4921] = ~(layer3_outputs[1257]);
    assign layer4_outputs[4922] = (layer3_outputs[2024]) & ~(layer3_outputs[2380]);
    assign layer4_outputs[4923] = ~((layer3_outputs[4190]) | (layer3_outputs[4978]));
    assign layer4_outputs[4924] = ~(layer3_outputs[690]);
    assign layer4_outputs[4925] = layer3_outputs[2272];
    assign layer4_outputs[4926] = ~(layer3_outputs[1320]) | (layer3_outputs[3481]);
    assign layer4_outputs[4927] = ~(layer3_outputs[3931]);
    assign layer4_outputs[4928] = ~(layer3_outputs[3134]);
    assign layer4_outputs[4929] = (layer3_outputs[2832]) | (layer3_outputs[4090]);
    assign layer4_outputs[4930] = layer3_outputs[778];
    assign layer4_outputs[4931] = ~(layer3_outputs[4642]);
    assign layer4_outputs[4932] = layer3_outputs[647];
    assign layer4_outputs[4933] = ~((layer3_outputs[4249]) & (layer3_outputs[1185]));
    assign layer4_outputs[4934] = ~(layer3_outputs[5076]) | (layer3_outputs[3789]);
    assign layer4_outputs[4935] = ~(layer3_outputs[3548]);
    assign layer4_outputs[4936] = (layer3_outputs[4747]) | (layer3_outputs[12]);
    assign layer4_outputs[4937] = layer3_outputs[3739];
    assign layer4_outputs[4938] = layer3_outputs[2921];
    assign layer4_outputs[4939] = layer3_outputs[3187];
    assign layer4_outputs[4940] = (layer3_outputs[4981]) & ~(layer3_outputs[605]);
    assign layer4_outputs[4941] = (layer3_outputs[2294]) ^ (layer3_outputs[3225]);
    assign layer4_outputs[4942] = 1'b1;
    assign layer4_outputs[4943] = layer3_outputs[3367];
    assign layer4_outputs[4944] = 1'b1;
    assign layer4_outputs[4945] = 1'b0;
    assign layer4_outputs[4946] = ~(layer3_outputs[2877]);
    assign layer4_outputs[4947] = ~((layer3_outputs[2649]) & (layer3_outputs[2885]));
    assign layer4_outputs[4948] = ~(layer3_outputs[4871]);
    assign layer4_outputs[4949] = ~((layer3_outputs[1142]) ^ (layer3_outputs[461]));
    assign layer4_outputs[4950] = (layer3_outputs[4480]) & (layer3_outputs[3065]);
    assign layer4_outputs[4951] = ~(layer3_outputs[1764]);
    assign layer4_outputs[4952] = (layer3_outputs[4318]) & ~(layer3_outputs[1552]);
    assign layer4_outputs[4953] = 1'b1;
    assign layer4_outputs[4954] = layer3_outputs[4924];
    assign layer4_outputs[4955] = (layer3_outputs[4583]) & ~(layer3_outputs[1898]);
    assign layer4_outputs[4956] = layer3_outputs[808];
    assign layer4_outputs[4957] = ~((layer3_outputs[562]) ^ (layer3_outputs[2733]));
    assign layer4_outputs[4958] = layer3_outputs[4313];
    assign layer4_outputs[4959] = layer3_outputs[2613];
    assign layer4_outputs[4960] = layer3_outputs[1253];
    assign layer4_outputs[4961] = ~(layer3_outputs[4767]) | (layer3_outputs[2382]);
    assign layer4_outputs[4962] = layer3_outputs[1674];
    assign layer4_outputs[4963] = (layer3_outputs[1828]) & (layer3_outputs[111]);
    assign layer4_outputs[4964] = 1'b1;
    assign layer4_outputs[4965] = ~(layer3_outputs[544]);
    assign layer4_outputs[4966] = layer3_outputs[953];
    assign layer4_outputs[4967] = layer3_outputs[4025];
    assign layer4_outputs[4968] = 1'b0;
    assign layer4_outputs[4969] = ~((layer3_outputs[2453]) | (layer3_outputs[3520]));
    assign layer4_outputs[4970] = layer3_outputs[131];
    assign layer4_outputs[4971] = 1'b1;
    assign layer4_outputs[4972] = (layer3_outputs[4179]) & (layer3_outputs[559]);
    assign layer4_outputs[4973] = (layer3_outputs[165]) ^ (layer3_outputs[4306]);
    assign layer4_outputs[4974] = layer3_outputs[3311];
    assign layer4_outputs[4975] = layer3_outputs[3694];
    assign layer4_outputs[4976] = layer3_outputs[1825];
    assign layer4_outputs[4977] = 1'b1;
    assign layer4_outputs[4978] = 1'b1;
    assign layer4_outputs[4979] = (layer3_outputs[1357]) & ~(layer3_outputs[3458]);
    assign layer4_outputs[4980] = ~(layer3_outputs[1676]);
    assign layer4_outputs[4981] = 1'b0;
    assign layer4_outputs[4982] = layer3_outputs[64];
    assign layer4_outputs[4983] = ~(layer3_outputs[4218]) | (layer3_outputs[4210]);
    assign layer4_outputs[4984] = (layer3_outputs[4903]) | (layer3_outputs[3271]);
    assign layer4_outputs[4985] = 1'b1;
    assign layer4_outputs[4986] = ~((layer3_outputs[248]) & (layer3_outputs[2144]));
    assign layer4_outputs[4987] = ~(layer3_outputs[2789]) | (layer3_outputs[4287]);
    assign layer4_outputs[4988] = layer3_outputs[4636];
    assign layer4_outputs[4989] = 1'b1;
    assign layer4_outputs[4990] = ~(layer3_outputs[1609]);
    assign layer4_outputs[4991] = ~((layer3_outputs[1853]) | (layer3_outputs[243]));
    assign layer4_outputs[4992] = ~((layer3_outputs[1933]) & (layer3_outputs[29]));
    assign layer4_outputs[4993] = ~(layer3_outputs[57]);
    assign layer4_outputs[4994] = 1'b0;
    assign layer4_outputs[4995] = 1'b0;
    assign layer4_outputs[4996] = ~(layer3_outputs[2782]);
    assign layer4_outputs[4997] = (layer3_outputs[3857]) | (layer3_outputs[2644]);
    assign layer4_outputs[4998] = ~(layer3_outputs[2643]);
    assign layer4_outputs[4999] = (layer3_outputs[4157]) ^ (layer3_outputs[4749]);
    assign layer4_outputs[5000] = ~(layer3_outputs[1868]) | (layer3_outputs[4967]);
    assign layer4_outputs[5001] = (layer3_outputs[1510]) & (layer3_outputs[2245]);
    assign layer4_outputs[5002] = (layer3_outputs[499]) | (layer3_outputs[2568]);
    assign layer4_outputs[5003] = layer3_outputs[2313];
    assign layer4_outputs[5004] = ~(layer3_outputs[4710]);
    assign layer4_outputs[5005] = (layer3_outputs[3552]) & ~(layer3_outputs[4379]);
    assign layer4_outputs[5006] = ~(layer3_outputs[312]);
    assign layer4_outputs[5007] = ~(layer3_outputs[4209]);
    assign layer4_outputs[5008] = 1'b0;
    assign layer4_outputs[5009] = ~(layer3_outputs[375]);
    assign layer4_outputs[5010] = layer3_outputs[2161];
    assign layer4_outputs[5011] = layer3_outputs[3949];
    assign layer4_outputs[5012] = ~(layer3_outputs[3983]);
    assign layer4_outputs[5013] = ~(layer3_outputs[4214]);
    assign layer4_outputs[5014] = (layer3_outputs[4227]) & (layer3_outputs[3347]);
    assign layer4_outputs[5015] = ~(layer3_outputs[4563]) | (layer3_outputs[4106]);
    assign layer4_outputs[5016] = ~(layer3_outputs[1206]);
    assign layer4_outputs[5017] = ~(layer3_outputs[2543]);
    assign layer4_outputs[5018] = ~((layer3_outputs[125]) | (layer3_outputs[1438]));
    assign layer4_outputs[5019] = (layer3_outputs[949]) & (layer3_outputs[4588]);
    assign layer4_outputs[5020] = ~(layer3_outputs[892]);
    assign layer4_outputs[5021] = (layer3_outputs[0]) & (layer3_outputs[2450]);
    assign layer4_outputs[5022] = ~(layer3_outputs[1842]);
    assign layer4_outputs[5023] = ~(layer3_outputs[1423]);
    assign layer4_outputs[5024] = layer3_outputs[4894];
    assign layer4_outputs[5025] = (layer3_outputs[2141]) & ~(layer3_outputs[15]);
    assign layer4_outputs[5026] = ~(layer3_outputs[99]) | (layer3_outputs[4821]);
    assign layer4_outputs[5027] = ~(layer3_outputs[901]);
    assign layer4_outputs[5028] = ~((layer3_outputs[1016]) ^ (layer3_outputs[1107]));
    assign layer4_outputs[5029] = (layer3_outputs[3363]) ^ (layer3_outputs[1216]);
    assign layer4_outputs[5030] = (layer3_outputs[718]) & ~(layer3_outputs[3700]);
    assign layer4_outputs[5031] = ~(layer3_outputs[963]);
    assign layer4_outputs[5032] = layer3_outputs[148];
    assign layer4_outputs[5033] = (layer3_outputs[49]) ^ (layer3_outputs[2738]);
    assign layer4_outputs[5034] = ~(layer3_outputs[2941]);
    assign layer4_outputs[5035] = ~(layer3_outputs[3743]);
    assign layer4_outputs[5036] = ~(layer3_outputs[3839]);
    assign layer4_outputs[5037] = ~(layer3_outputs[2459]);
    assign layer4_outputs[5038] = ~(layer3_outputs[3176]);
    assign layer4_outputs[5039] = ~(layer3_outputs[1533]) | (layer3_outputs[4754]);
    assign layer4_outputs[5040] = (layer3_outputs[273]) & ~(layer3_outputs[4188]);
    assign layer4_outputs[5041] = layer3_outputs[3350];
    assign layer4_outputs[5042] = 1'b0;
    assign layer4_outputs[5043] = (layer3_outputs[1404]) & ~(layer3_outputs[1933]);
    assign layer4_outputs[5044] = layer3_outputs[2409];
    assign layer4_outputs[5045] = ~(layer3_outputs[4261]) | (layer3_outputs[3314]);
    assign layer4_outputs[5046] = ~(layer3_outputs[3194]) | (layer3_outputs[1241]);
    assign layer4_outputs[5047] = ~(layer3_outputs[1210]) | (layer3_outputs[4376]);
    assign layer4_outputs[5048] = ~(layer3_outputs[4712]) | (layer3_outputs[2405]);
    assign layer4_outputs[5049] = (layer3_outputs[3095]) & (layer3_outputs[4451]);
    assign layer4_outputs[5050] = 1'b1;
    assign layer4_outputs[5051] = layer3_outputs[1041];
    assign layer4_outputs[5052] = layer3_outputs[1379];
    assign layer4_outputs[5053] = layer3_outputs[2824];
    assign layer4_outputs[5054] = ~(layer3_outputs[374]);
    assign layer4_outputs[5055] = (layer3_outputs[3129]) & ~(layer3_outputs[301]);
    assign layer4_outputs[5056] = ~(layer3_outputs[3674]) | (layer3_outputs[4443]);
    assign layer4_outputs[5057] = ~(layer3_outputs[4650]);
    assign layer4_outputs[5058] = (layer3_outputs[3903]) & (layer3_outputs[4794]);
    assign layer4_outputs[5059] = ~((layer3_outputs[175]) ^ (layer3_outputs[3626]));
    assign layer4_outputs[5060] = (layer3_outputs[4165]) | (layer3_outputs[3949]);
    assign layer4_outputs[5061] = ~((layer3_outputs[4652]) & (layer3_outputs[3922]));
    assign layer4_outputs[5062] = ~(layer3_outputs[1031]);
    assign layer4_outputs[5063] = (layer3_outputs[4448]) ^ (layer3_outputs[3759]);
    assign layer4_outputs[5064] = layer3_outputs[906];
    assign layer4_outputs[5065] = ~((layer3_outputs[2359]) & (layer3_outputs[4659]));
    assign layer4_outputs[5066] = ~(layer3_outputs[3704]);
    assign layer4_outputs[5067] = (layer3_outputs[4483]) ^ (layer3_outputs[2576]);
    assign layer4_outputs[5068] = (layer3_outputs[2514]) & ~(layer3_outputs[2575]);
    assign layer4_outputs[5069] = 1'b0;
    assign layer4_outputs[5070] = (layer3_outputs[2828]) ^ (layer3_outputs[2321]);
    assign layer4_outputs[5071] = ~(layer3_outputs[871]);
    assign layer4_outputs[5072] = ~((layer3_outputs[4979]) ^ (layer3_outputs[645]));
    assign layer4_outputs[5073] = ~(layer3_outputs[3426]);
    assign layer4_outputs[5074] = layer3_outputs[4555];
    assign layer4_outputs[5075] = layer3_outputs[2064];
    assign layer4_outputs[5076] = (layer3_outputs[3668]) ^ (layer3_outputs[3993]);
    assign layer4_outputs[5077] = ~((layer3_outputs[2092]) & (layer3_outputs[4832]));
    assign layer4_outputs[5078] = layer3_outputs[4826];
    assign layer4_outputs[5079] = layer3_outputs[3043];
    assign layer4_outputs[5080] = (layer3_outputs[4422]) | (layer3_outputs[2741]);
    assign layer4_outputs[5081] = (layer3_outputs[3099]) | (layer3_outputs[923]);
    assign layer4_outputs[5082] = 1'b0;
    assign layer4_outputs[5083] = ~(layer3_outputs[1738]);
    assign layer4_outputs[5084] = layer3_outputs[3310];
    assign layer4_outputs[5085] = ~(layer3_outputs[4868]) | (layer3_outputs[3936]);
    assign layer4_outputs[5086] = layer3_outputs[4884];
    assign layer4_outputs[5087] = 1'b1;
    assign layer4_outputs[5088] = ~(layer3_outputs[4061]) | (layer3_outputs[1882]);
    assign layer4_outputs[5089] = layer3_outputs[4500];
    assign layer4_outputs[5090] = layer3_outputs[4292];
    assign layer4_outputs[5091] = ~(layer3_outputs[3756]);
    assign layer4_outputs[5092] = layer3_outputs[1058];
    assign layer4_outputs[5093] = ~(layer3_outputs[46]);
    assign layer4_outputs[5094] = layer3_outputs[5089];
    assign layer4_outputs[5095] = ~(layer3_outputs[4053]);
    assign layer4_outputs[5096] = ~(layer3_outputs[130]) | (layer3_outputs[2491]);
    assign layer4_outputs[5097] = 1'b0;
    assign layer4_outputs[5098] = ~(layer3_outputs[2800]) | (layer3_outputs[3952]);
    assign layer4_outputs[5099] = 1'b1;
    assign layer4_outputs[5100] = (layer3_outputs[723]) & (layer3_outputs[1562]);
    assign layer4_outputs[5101] = ~(layer3_outputs[2610]);
    assign layer4_outputs[5102] = ~(layer3_outputs[1928]) | (layer3_outputs[4846]);
    assign layer4_outputs[5103] = ~(layer3_outputs[3436]);
    assign layer4_outputs[5104] = (layer3_outputs[565]) & ~(layer3_outputs[4903]);
    assign layer4_outputs[5105] = ~(layer3_outputs[3569]) | (layer3_outputs[1584]);
    assign layer4_outputs[5106] = layer3_outputs[1384];
    assign layer4_outputs[5107] = (layer3_outputs[4613]) & ~(layer3_outputs[30]);
    assign layer4_outputs[5108] = (layer3_outputs[846]) | (layer3_outputs[362]);
    assign layer4_outputs[5109] = layer3_outputs[2156];
    assign layer4_outputs[5110] = (layer3_outputs[3348]) ^ (layer3_outputs[927]);
    assign layer4_outputs[5111] = (layer3_outputs[442]) ^ (layer3_outputs[180]);
    assign layer4_outputs[5112] = ~(layer3_outputs[3387]);
    assign layer4_outputs[5113] = ~((layer3_outputs[3852]) ^ (layer3_outputs[4121]));
    assign layer4_outputs[5114] = (layer3_outputs[702]) | (layer3_outputs[3844]);
    assign layer4_outputs[5115] = ~(layer3_outputs[2220]) | (layer3_outputs[804]);
    assign layer4_outputs[5116] = layer3_outputs[4863];
    assign layer4_outputs[5117] = ~(layer3_outputs[2350]);
    assign layer4_outputs[5118] = (layer3_outputs[5102]) ^ (layer3_outputs[1476]);
    assign layer4_outputs[5119] = ~(layer3_outputs[3956]);
    assign layer5_outputs[0] = layer4_outputs[497];
    assign layer5_outputs[1] = layer4_outputs[3317];
    assign layer5_outputs[2] = layer4_outputs[4878];
    assign layer5_outputs[3] = ~((layer4_outputs[121]) & (layer4_outputs[1952]));
    assign layer5_outputs[4] = ~(layer4_outputs[2389]) | (layer4_outputs[3084]);
    assign layer5_outputs[5] = ~((layer4_outputs[1789]) ^ (layer4_outputs[1722]));
    assign layer5_outputs[6] = ~(layer4_outputs[4063]);
    assign layer5_outputs[7] = (layer4_outputs[5062]) | (layer4_outputs[2115]);
    assign layer5_outputs[8] = ~(layer4_outputs[476]);
    assign layer5_outputs[9] = layer4_outputs[1607];
    assign layer5_outputs[10] = layer4_outputs[2173];
    assign layer5_outputs[11] = ~(layer4_outputs[2419]) | (layer4_outputs[2667]);
    assign layer5_outputs[12] = ~((layer4_outputs[4141]) ^ (layer4_outputs[3310]));
    assign layer5_outputs[13] = (layer4_outputs[4906]) & ~(layer4_outputs[327]);
    assign layer5_outputs[14] = ~(layer4_outputs[3718]) | (layer4_outputs[2526]);
    assign layer5_outputs[15] = layer4_outputs[2690];
    assign layer5_outputs[16] = ~((layer4_outputs[3160]) ^ (layer4_outputs[3902]));
    assign layer5_outputs[17] = layer4_outputs[4411];
    assign layer5_outputs[18] = ~(layer4_outputs[1894]);
    assign layer5_outputs[19] = (layer4_outputs[4960]) | (layer4_outputs[2427]);
    assign layer5_outputs[20] = ~(layer4_outputs[127]);
    assign layer5_outputs[21] = (layer4_outputs[4263]) & ~(layer4_outputs[2391]);
    assign layer5_outputs[22] = ~(layer4_outputs[2835]);
    assign layer5_outputs[23] = layer4_outputs[3721];
    assign layer5_outputs[24] = (layer4_outputs[5068]) ^ (layer4_outputs[4058]);
    assign layer5_outputs[25] = layer4_outputs[3355];
    assign layer5_outputs[26] = 1'b1;
    assign layer5_outputs[27] = (layer4_outputs[4075]) | (layer4_outputs[3766]);
    assign layer5_outputs[28] = layer4_outputs[224];
    assign layer5_outputs[29] = layer4_outputs[3274];
    assign layer5_outputs[30] = ~(layer4_outputs[4925]) | (layer4_outputs[3375]);
    assign layer5_outputs[31] = layer4_outputs[1661];
    assign layer5_outputs[32] = ~(layer4_outputs[4736]) | (layer4_outputs[2988]);
    assign layer5_outputs[33] = ~((layer4_outputs[3518]) | (layer4_outputs[3181]));
    assign layer5_outputs[34] = ~(layer4_outputs[691]);
    assign layer5_outputs[35] = ~(layer4_outputs[1816]) | (layer4_outputs[1209]);
    assign layer5_outputs[36] = layer4_outputs[761];
    assign layer5_outputs[37] = ~(layer4_outputs[476]);
    assign layer5_outputs[38] = ~((layer4_outputs[3292]) | (layer4_outputs[3000]));
    assign layer5_outputs[39] = ~((layer4_outputs[3139]) ^ (layer4_outputs[2263]));
    assign layer5_outputs[40] = (layer4_outputs[2308]) & ~(layer4_outputs[4182]);
    assign layer5_outputs[41] = ~(layer4_outputs[4984]);
    assign layer5_outputs[42] = layer4_outputs[1436];
    assign layer5_outputs[43] = layer4_outputs[795];
    assign layer5_outputs[44] = ~(layer4_outputs[56]);
    assign layer5_outputs[45] = (layer4_outputs[1174]) & ~(layer4_outputs[169]);
    assign layer5_outputs[46] = ~(layer4_outputs[673]);
    assign layer5_outputs[47] = layer4_outputs[2096];
    assign layer5_outputs[48] = layer4_outputs[5047];
    assign layer5_outputs[49] = ~(layer4_outputs[1645]);
    assign layer5_outputs[50] = (layer4_outputs[4880]) & ~(layer4_outputs[2072]);
    assign layer5_outputs[51] = 1'b0;
    assign layer5_outputs[52] = (layer4_outputs[2637]) & ~(layer4_outputs[1011]);
    assign layer5_outputs[53] = ~((layer4_outputs[841]) & (layer4_outputs[4580]));
    assign layer5_outputs[54] = ~((layer4_outputs[4751]) & (layer4_outputs[1410]));
    assign layer5_outputs[55] = (layer4_outputs[1395]) | (layer4_outputs[422]);
    assign layer5_outputs[56] = ~(layer4_outputs[272]) | (layer4_outputs[1535]);
    assign layer5_outputs[57] = (layer4_outputs[5107]) ^ (layer4_outputs[4514]);
    assign layer5_outputs[58] = (layer4_outputs[4783]) & ~(layer4_outputs[648]);
    assign layer5_outputs[59] = 1'b0;
    assign layer5_outputs[60] = (layer4_outputs[4524]) & ~(layer4_outputs[2695]);
    assign layer5_outputs[61] = 1'b0;
    assign layer5_outputs[62] = ~(layer4_outputs[2844]);
    assign layer5_outputs[63] = ~(layer4_outputs[229]);
    assign layer5_outputs[64] = layer4_outputs[3766];
    assign layer5_outputs[65] = (layer4_outputs[1289]) & ~(layer4_outputs[374]);
    assign layer5_outputs[66] = (layer4_outputs[3667]) & ~(layer4_outputs[4447]);
    assign layer5_outputs[67] = (layer4_outputs[4351]) & ~(layer4_outputs[1698]);
    assign layer5_outputs[68] = (layer4_outputs[1180]) | (layer4_outputs[3477]);
    assign layer5_outputs[69] = ~(layer4_outputs[347]);
    assign layer5_outputs[70] = ~((layer4_outputs[2693]) ^ (layer4_outputs[4545]));
    assign layer5_outputs[71] = ~(layer4_outputs[1746]);
    assign layer5_outputs[72] = (layer4_outputs[523]) ^ (layer4_outputs[3319]);
    assign layer5_outputs[73] = ~((layer4_outputs[2735]) & (layer4_outputs[3999]));
    assign layer5_outputs[74] = (layer4_outputs[2743]) & ~(layer4_outputs[645]);
    assign layer5_outputs[75] = ~(layer4_outputs[2012]);
    assign layer5_outputs[76] = ~(layer4_outputs[1357]) | (layer4_outputs[4855]);
    assign layer5_outputs[77] = layer4_outputs[4307];
    assign layer5_outputs[78] = layer4_outputs[3513];
    assign layer5_outputs[79] = (layer4_outputs[4203]) & (layer4_outputs[2212]);
    assign layer5_outputs[80] = ~(layer4_outputs[2173]);
    assign layer5_outputs[81] = (layer4_outputs[2932]) & ~(layer4_outputs[1342]);
    assign layer5_outputs[82] = layer4_outputs[3210];
    assign layer5_outputs[83] = ~(layer4_outputs[4448]) | (layer4_outputs[1424]);
    assign layer5_outputs[84] = layer4_outputs[2048];
    assign layer5_outputs[85] = layer4_outputs[1876];
    assign layer5_outputs[86] = 1'b0;
    assign layer5_outputs[87] = ~(layer4_outputs[4059]);
    assign layer5_outputs[88] = (layer4_outputs[4446]) & ~(layer4_outputs[2034]);
    assign layer5_outputs[89] = 1'b0;
    assign layer5_outputs[90] = ~((layer4_outputs[4857]) & (layer4_outputs[2722]));
    assign layer5_outputs[91] = (layer4_outputs[4065]) & ~(layer4_outputs[842]);
    assign layer5_outputs[92] = 1'b0;
    assign layer5_outputs[93] = 1'b0;
    assign layer5_outputs[94] = ~((layer4_outputs[3735]) & (layer4_outputs[2971]));
    assign layer5_outputs[95] = 1'b1;
    assign layer5_outputs[96] = ~(layer4_outputs[4900]);
    assign layer5_outputs[97] = ~(layer4_outputs[2688]);
    assign layer5_outputs[98] = ~(layer4_outputs[3804]);
    assign layer5_outputs[99] = ~(layer4_outputs[110]) | (layer4_outputs[3503]);
    assign layer5_outputs[100] = ~(layer4_outputs[2029]);
    assign layer5_outputs[101] = ~(layer4_outputs[709]) | (layer4_outputs[828]);
    assign layer5_outputs[102] = layer4_outputs[913];
    assign layer5_outputs[103] = (layer4_outputs[2091]) | (layer4_outputs[883]);
    assign layer5_outputs[104] = ~(layer4_outputs[21]);
    assign layer5_outputs[105] = (layer4_outputs[2035]) & ~(layer4_outputs[4174]);
    assign layer5_outputs[106] = (layer4_outputs[2228]) ^ (layer4_outputs[1854]);
    assign layer5_outputs[107] = ~(layer4_outputs[4382]);
    assign layer5_outputs[108] = (layer4_outputs[818]) & (layer4_outputs[2407]);
    assign layer5_outputs[109] = ~((layer4_outputs[2515]) | (layer4_outputs[4693]));
    assign layer5_outputs[110] = ~(layer4_outputs[1813]);
    assign layer5_outputs[111] = layer4_outputs[3061];
    assign layer5_outputs[112] = layer4_outputs[942];
    assign layer5_outputs[113] = ~(layer4_outputs[750]) | (layer4_outputs[1787]);
    assign layer5_outputs[114] = layer4_outputs[4020];
    assign layer5_outputs[115] = ~(layer4_outputs[4537]);
    assign layer5_outputs[116] = layer4_outputs[2893];
    assign layer5_outputs[117] = ~((layer4_outputs[2919]) ^ (layer4_outputs[2255]));
    assign layer5_outputs[118] = layer4_outputs[1389];
    assign layer5_outputs[119] = ~((layer4_outputs[1430]) & (layer4_outputs[983]));
    assign layer5_outputs[120] = (layer4_outputs[3406]) & ~(layer4_outputs[4430]);
    assign layer5_outputs[121] = ~(layer4_outputs[54]);
    assign layer5_outputs[122] = layer4_outputs[4311];
    assign layer5_outputs[123] = (layer4_outputs[3178]) | (layer4_outputs[271]);
    assign layer5_outputs[124] = (layer4_outputs[4756]) | (layer4_outputs[4731]);
    assign layer5_outputs[125] = 1'b0;
    assign layer5_outputs[126] = ~(layer4_outputs[15]);
    assign layer5_outputs[127] = 1'b1;
    assign layer5_outputs[128] = ~(layer4_outputs[2828]);
    assign layer5_outputs[129] = ~(layer4_outputs[2643]);
    assign layer5_outputs[130] = ~(layer4_outputs[1408]);
    assign layer5_outputs[131] = layer4_outputs[2671];
    assign layer5_outputs[132] = (layer4_outputs[4370]) ^ (layer4_outputs[4500]);
    assign layer5_outputs[133] = layer4_outputs[4164];
    assign layer5_outputs[134] = ~(layer4_outputs[3837]);
    assign layer5_outputs[135] = layer4_outputs[484];
    assign layer5_outputs[136] = 1'b1;
    assign layer5_outputs[137] = layer4_outputs[1619];
    assign layer5_outputs[138] = ~(layer4_outputs[3972]);
    assign layer5_outputs[139] = (layer4_outputs[31]) ^ (layer4_outputs[1515]);
    assign layer5_outputs[140] = ~((layer4_outputs[2457]) ^ (layer4_outputs[4467]));
    assign layer5_outputs[141] = 1'b0;
    assign layer5_outputs[142] = (layer4_outputs[4025]) & ~(layer4_outputs[173]);
    assign layer5_outputs[143] = (layer4_outputs[75]) ^ (layer4_outputs[1919]);
    assign layer5_outputs[144] = ~(layer4_outputs[3845]);
    assign layer5_outputs[145] = layer4_outputs[3120];
    assign layer5_outputs[146] = layer4_outputs[4797];
    assign layer5_outputs[147] = ~(layer4_outputs[4891]);
    assign layer5_outputs[148] = (layer4_outputs[3520]) ^ (layer4_outputs[2808]);
    assign layer5_outputs[149] = 1'b1;
    assign layer5_outputs[150] = ~(layer4_outputs[1844]);
    assign layer5_outputs[151] = ~(layer4_outputs[833]);
    assign layer5_outputs[152] = ~((layer4_outputs[4]) & (layer4_outputs[2335]));
    assign layer5_outputs[153] = ~(layer4_outputs[4512]) | (layer4_outputs[2861]);
    assign layer5_outputs[154] = layer4_outputs[1793];
    assign layer5_outputs[155] = 1'b0;
    assign layer5_outputs[156] = ~(layer4_outputs[3219]);
    assign layer5_outputs[157] = layer4_outputs[3007];
    assign layer5_outputs[158] = ~(layer4_outputs[447]);
    assign layer5_outputs[159] = ~((layer4_outputs[3005]) & (layer4_outputs[483]));
    assign layer5_outputs[160] = ~(layer4_outputs[1182]);
    assign layer5_outputs[161] = (layer4_outputs[1898]) & (layer4_outputs[1363]);
    assign layer5_outputs[162] = ~(layer4_outputs[3787]);
    assign layer5_outputs[163] = (layer4_outputs[1568]) ^ (layer4_outputs[2007]);
    assign layer5_outputs[164] = ~(layer4_outputs[1198]);
    assign layer5_outputs[165] = (layer4_outputs[3001]) & ~(layer4_outputs[81]);
    assign layer5_outputs[166] = layer4_outputs[3376];
    assign layer5_outputs[167] = ~((layer4_outputs[2570]) ^ (layer4_outputs[1519]));
    assign layer5_outputs[168] = ~((layer4_outputs[2927]) | (layer4_outputs[4730]));
    assign layer5_outputs[169] = ~((layer4_outputs[3551]) ^ (layer4_outputs[3642]));
    assign layer5_outputs[170] = (layer4_outputs[3294]) | (layer4_outputs[4560]);
    assign layer5_outputs[171] = ~((layer4_outputs[4829]) & (layer4_outputs[2609]));
    assign layer5_outputs[172] = ~(layer4_outputs[2351]) | (layer4_outputs[4633]);
    assign layer5_outputs[173] = layer4_outputs[3773];
    assign layer5_outputs[174] = layer4_outputs[5050];
    assign layer5_outputs[175] = 1'b1;
    assign layer5_outputs[176] = ~(layer4_outputs[187]);
    assign layer5_outputs[177] = ~(layer4_outputs[4526]);
    assign layer5_outputs[178] = ~(layer4_outputs[3323]);
    assign layer5_outputs[179] = ~(layer4_outputs[4323]);
    assign layer5_outputs[180] = ~(layer4_outputs[1622]);
    assign layer5_outputs[181] = ~((layer4_outputs[4586]) & (layer4_outputs[2032]));
    assign layer5_outputs[182] = ~(layer4_outputs[265]);
    assign layer5_outputs[183] = (layer4_outputs[111]) & ~(layer4_outputs[3943]);
    assign layer5_outputs[184] = ~(layer4_outputs[4774]);
    assign layer5_outputs[185] = (layer4_outputs[5067]) & ~(layer4_outputs[3647]);
    assign layer5_outputs[186] = ~((layer4_outputs[3539]) | (layer4_outputs[1750]));
    assign layer5_outputs[187] = layer4_outputs[1621];
    assign layer5_outputs[188] = (layer4_outputs[4709]) & ~(layer4_outputs[4377]);
    assign layer5_outputs[189] = layer4_outputs[2215];
    assign layer5_outputs[190] = layer4_outputs[1150];
    assign layer5_outputs[191] = layer4_outputs[3763];
    assign layer5_outputs[192] = ~((layer4_outputs[2595]) & (layer4_outputs[4707]));
    assign layer5_outputs[193] = (layer4_outputs[3243]) & ~(layer4_outputs[3068]);
    assign layer5_outputs[194] = ~(layer4_outputs[4527]);
    assign layer5_outputs[195] = ~(layer4_outputs[3790]);
    assign layer5_outputs[196] = layer4_outputs[223];
    assign layer5_outputs[197] = (layer4_outputs[1875]) & ~(layer4_outputs[478]);
    assign layer5_outputs[198] = ~(layer4_outputs[2510]);
    assign layer5_outputs[199] = ~(layer4_outputs[1800]);
    assign layer5_outputs[200] = 1'b0;
    assign layer5_outputs[201] = ~(layer4_outputs[3578]) | (layer4_outputs[1320]);
    assign layer5_outputs[202] = ~(layer4_outputs[5030]);
    assign layer5_outputs[203] = layer4_outputs[3331];
    assign layer5_outputs[204] = (layer4_outputs[1889]) & ~(layer4_outputs[3059]);
    assign layer5_outputs[205] = layer4_outputs[2664];
    assign layer5_outputs[206] = ~((layer4_outputs[570]) ^ (layer4_outputs[2304]));
    assign layer5_outputs[207] = (layer4_outputs[4163]) | (layer4_outputs[2375]);
    assign layer5_outputs[208] = layer4_outputs[1981];
    assign layer5_outputs[209] = ~(layer4_outputs[1471]);
    assign layer5_outputs[210] = (layer4_outputs[3184]) & ~(layer4_outputs[3973]);
    assign layer5_outputs[211] = ~(layer4_outputs[2726]);
    assign layer5_outputs[212] = (layer4_outputs[2896]) & ~(layer4_outputs[1778]);
    assign layer5_outputs[213] = ~(layer4_outputs[4514]);
    assign layer5_outputs[214] = (layer4_outputs[2294]) & (layer4_outputs[4027]);
    assign layer5_outputs[215] = ~((layer4_outputs[1191]) & (layer4_outputs[2049]));
    assign layer5_outputs[216] = 1'b1;
    assign layer5_outputs[217] = ~((layer4_outputs[4378]) | (layer4_outputs[4242]));
    assign layer5_outputs[218] = ~(layer4_outputs[1869]);
    assign layer5_outputs[219] = layer4_outputs[2419];
    assign layer5_outputs[220] = (layer4_outputs[2302]) & ~(layer4_outputs[3011]);
    assign layer5_outputs[221] = (layer4_outputs[3018]) & (layer4_outputs[1583]);
    assign layer5_outputs[222] = layer4_outputs[1230];
    assign layer5_outputs[223] = ~(layer4_outputs[391]);
    assign layer5_outputs[224] = layer4_outputs[557];
    assign layer5_outputs[225] = layer4_outputs[1186];
    assign layer5_outputs[226] = ~(layer4_outputs[2115]) | (layer4_outputs[1050]);
    assign layer5_outputs[227] = (layer4_outputs[3468]) & ~(layer4_outputs[3662]);
    assign layer5_outputs[228] = layer4_outputs[1474];
    assign layer5_outputs[229] = ~(layer4_outputs[4680]);
    assign layer5_outputs[230] = 1'b1;
    assign layer5_outputs[231] = ~(layer4_outputs[460]);
    assign layer5_outputs[232] = ~(layer4_outputs[1742]);
    assign layer5_outputs[233] = layer4_outputs[4215];
    assign layer5_outputs[234] = layer4_outputs[1199];
    assign layer5_outputs[235] = (layer4_outputs[4729]) & (layer4_outputs[3595]);
    assign layer5_outputs[236] = ~(layer4_outputs[1511]);
    assign layer5_outputs[237] = layer4_outputs[3131];
    assign layer5_outputs[238] = layer4_outputs[3391];
    assign layer5_outputs[239] = ~(layer4_outputs[3658]);
    assign layer5_outputs[240] = ~(layer4_outputs[2544]) | (layer4_outputs[1943]);
    assign layer5_outputs[241] = layer4_outputs[53];
    assign layer5_outputs[242] = 1'b0;
    assign layer5_outputs[243] = ~((layer4_outputs[3613]) & (layer4_outputs[2529]));
    assign layer5_outputs[244] = layer4_outputs[2574];
    assign layer5_outputs[245] = ~((layer4_outputs[2403]) ^ (layer4_outputs[855]));
    assign layer5_outputs[246] = ~(layer4_outputs[2019]);
    assign layer5_outputs[247] = layer4_outputs[339];
    assign layer5_outputs[248] = layer4_outputs[2650];
    assign layer5_outputs[249] = layer4_outputs[1175];
    assign layer5_outputs[250] = layer4_outputs[4336];
    assign layer5_outputs[251] = ~(layer4_outputs[662]);
    assign layer5_outputs[252] = ~(layer4_outputs[5119]) | (layer4_outputs[4804]);
    assign layer5_outputs[253] = ~(layer4_outputs[2439]);
    assign layer5_outputs[254] = ~(layer4_outputs[4718]) | (layer4_outputs[1076]);
    assign layer5_outputs[255] = ~((layer4_outputs[783]) | (layer4_outputs[678]));
    assign layer5_outputs[256] = (layer4_outputs[5041]) ^ (layer4_outputs[3314]);
    assign layer5_outputs[257] = (layer4_outputs[2060]) & ~(layer4_outputs[1693]);
    assign layer5_outputs[258] = layer4_outputs[508];
    assign layer5_outputs[259] = ~((layer4_outputs[3908]) ^ (layer4_outputs[1890]));
    assign layer5_outputs[260] = (layer4_outputs[2106]) & (layer4_outputs[1190]);
    assign layer5_outputs[261] = ~(layer4_outputs[3734]);
    assign layer5_outputs[262] = ~(layer4_outputs[3374]);
    assign layer5_outputs[263] = (layer4_outputs[470]) & (layer4_outputs[3048]);
    assign layer5_outputs[264] = ~(layer4_outputs[571]);
    assign layer5_outputs[265] = 1'b0;
    assign layer5_outputs[266] = ~(layer4_outputs[2954]);
    assign layer5_outputs[267] = ~(layer4_outputs[4003]);
    assign layer5_outputs[268] = layer4_outputs[3287];
    assign layer5_outputs[269] = ~(layer4_outputs[1779]);
    assign layer5_outputs[270] = (layer4_outputs[2857]) & ~(layer4_outputs[4521]);
    assign layer5_outputs[271] = (layer4_outputs[2992]) & (layer4_outputs[207]);
    assign layer5_outputs[272] = 1'b0;
    assign layer5_outputs[273] = ~(layer4_outputs[1571]);
    assign layer5_outputs[274] = layer4_outputs[2203];
    assign layer5_outputs[275] = (layer4_outputs[3123]) & ~(layer4_outputs[3899]);
    assign layer5_outputs[276] = layer4_outputs[724];
    assign layer5_outputs[277] = ~(layer4_outputs[2849]);
    assign layer5_outputs[278] = (layer4_outputs[3294]) | (layer4_outputs[3405]);
    assign layer5_outputs[279] = ~(layer4_outputs[4362]) | (layer4_outputs[2438]);
    assign layer5_outputs[280] = ~(layer4_outputs[764]) | (layer4_outputs[4507]);
    assign layer5_outputs[281] = layer4_outputs[4045];
    assign layer5_outputs[282] = (layer4_outputs[3394]) & ~(layer4_outputs[71]);
    assign layer5_outputs[283] = ~(layer4_outputs[3937]);
    assign layer5_outputs[284] = ~(layer4_outputs[1731]);
    assign layer5_outputs[285] = layer4_outputs[2820];
    assign layer5_outputs[286] = (layer4_outputs[665]) ^ (layer4_outputs[1468]);
    assign layer5_outputs[287] = layer4_outputs[1505];
    assign layer5_outputs[288] = (layer4_outputs[4738]) & ~(layer4_outputs[1288]);
    assign layer5_outputs[289] = (layer4_outputs[4668]) | (layer4_outputs[4768]);
    assign layer5_outputs[290] = ~(layer4_outputs[2693]) | (layer4_outputs[2282]);
    assign layer5_outputs[291] = (layer4_outputs[704]) ^ (layer4_outputs[2044]);
    assign layer5_outputs[292] = layer4_outputs[3614];
    assign layer5_outputs[293] = ~(layer4_outputs[4812]) | (layer4_outputs[837]);
    assign layer5_outputs[294] = ~(layer4_outputs[1407]);
    assign layer5_outputs[295] = layer4_outputs[434];
    assign layer5_outputs[296] = layer4_outputs[2605];
    assign layer5_outputs[297] = layer4_outputs[905];
    assign layer5_outputs[298] = ~((layer4_outputs[393]) ^ (layer4_outputs[3452]));
    assign layer5_outputs[299] = ~(layer4_outputs[2922]) | (layer4_outputs[1273]);
    assign layer5_outputs[300] = ~((layer4_outputs[2543]) | (layer4_outputs[3805]));
    assign layer5_outputs[301] = ~(layer4_outputs[1449]);
    assign layer5_outputs[302] = layer4_outputs[4998];
    assign layer5_outputs[303] = layer4_outputs[551];
    assign layer5_outputs[304] = ~(layer4_outputs[3632]);
    assign layer5_outputs[305] = 1'b0;
    assign layer5_outputs[306] = (layer4_outputs[595]) & ~(layer4_outputs[2999]);
    assign layer5_outputs[307] = layer4_outputs[2338];
    assign layer5_outputs[308] = 1'b1;
    assign layer5_outputs[309] = ~(layer4_outputs[3152]);
    assign layer5_outputs[310] = (layer4_outputs[1083]) & (layer4_outputs[1832]);
    assign layer5_outputs[311] = ~(layer4_outputs[2352]);
    assign layer5_outputs[312] = (layer4_outputs[2867]) & ~(layer4_outputs[2013]);
    assign layer5_outputs[313] = ~(layer4_outputs[2721]) | (layer4_outputs[5106]);
    assign layer5_outputs[314] = ~((layer4_outputs[4138]) ^ (layer4_outputs[4281]));
    assign layer5_outputs[315] = ~(layer4_outputs[2026]);
    assign layer5_outputs[316] = (layer4_outputs[1804]) & ~(layer4_outputs[1904]);
    assign layer5_outputs[317] = (layer4_outputs[2863]) & (layer4_outputs[4089]);
    assign layer5_outputs[318] = (layer4_outputs[473]) & ~(layer4_outputs[5000]);
    assign layer5_outputs[319] = layer4_outputs[528];
    assign layer5_outputs[320] = (layer4_outputs[1552]) & (layer4_outputs[2729]);
    assign layer5_outputs[321] = layer4_outputs[1302];
    assign layer5_outputs[322] = layer4_outputs[92];
    assign layer5_outputs[323] = ~((layer4_outputs[3622]) ^ (layer4_outputs[823]));
    assign layer5_outputs[324] = (layer4_outputs[5119]) | (layer4_outputs[2182]);
    assign layer5_outputs[325] = (layer4_outputs[3215]) & ~(layer4_outputs[4755]);
    assign layer5_outputs[326] = layer4_outputs[2493];
    assign layer5_outputs[327] = ~(layer4_outputs[2662]);
    assign layer5_outputs[328] = ~(layer4_outputs[658]) | (layer4_outputs[3775]);
    assign layer5_outputs[329] = ~((layer4_outputs[216]) | (layer4_outputs[1394]));
    assign layer5_outputs[330] = ~(layer4_outputs[3229]);
    assign layer5_outputs[331] = ~(layer4_outputs[4235]) | (layer4_outputs[3523]);
    assign layer5_outputs[332] = ~((layer4_outputs[3206]) & (layer4_outputs[1760]));
    assign layer5_outputs[333] = layer4_outputs[1241];
    assign layer5_outputs[334] = (layer4_outputs[1802]) & ~(layer4_outputs[2585]);
    assign layer5_outputs[335] = layer4_outputs[3729];
    assign layer5_outputs[336] = ~(layer4_outputs[3826]) | (layer4_outputs[1766]);
    assign layer5_outputs[337] = ~(layer4_outputs[2608]);
    assign layer5_outputs[338] = ~((layer4_outputs[4049]) ^ (layer4_outputs[4500]));
    assign layer5_outputs[339] = ~(layer4_outputs[568]);
    assign layer5_outputs[340] = layer4_outputs[9];
    assign layer5_outputs[341] = layer4_outputs[4868];
    assign layer5_outputs[342] = (layer4_outputs[2225]) & ~(layer4_outputs[2911]);
    assign layer5_outputs[343] = ~((layer4_outputs[2730]) | (layer4_outputs[4021]));
    assign layer5_outputs[344] = ~(layer4_outputs[1928]);
    assign layer5_outputs[345] = layer4_outputs[433];
    assign layer5_outputs[346] = (layer4_outputs[4497]) & ~(layer4_outputs[59]);
    assign layer5_outputs[347] = (layer4_outputs[3569]) ^ (layer4_outputs[2675]);
    assign layer5_outputs[348] = (layer4_outputs[4519]) & ~(layer4_outputs[3698]);
    assign layer5_outputs[349] = layer4_outputs[3988];
    assign layer5_outputs[350] = (layer4_outputs[1141]) | (layer4_outputs[992]);
    assign layer5_outputs[351] = ~(layer4_outputs[543]);
    assign layer5_outputs[352] = ~(layer4_outputs[1357]);
    assign layer5_outputs[353] = ~(layer4_outputs[1444]) | (layer4_outputs[3630]);
    assign layer5_outputs[354] = ~((layer4_outputs[4110]) & (layer4_outputs[2599]));
    assign layer5_outputs[355] = layer4_outputs[3583];
    assign layer5_outputs[356] = (layer4_outputs[177]) ^ (layer4_outputs[369]);
    assign layer5_outputs[357] = ~((layer4_outputs[1829]) & (layer4_outputs[3101]));
    assign layer5_outputs[358] = ~(layer4_outputs[160]);
    assign layer5_outputs[359] = ~((layer4_outputs[3314]) ^ (layer4_outputs[4384]));
    assign layer5_outputs[360] = 1'b0;
    assign layer5_outputs[361] = layer4_outputs[1396];
    assign layer5_outputs[362] = ~(layer4_outputs[417]) | (layer4_outputs[731]);
    assign layer5_outputs[363] = (layer4_outputs[4821]) | (layer4_outputs[398]);
    assign layer5_outputs[364] = ~(layer4_outputs[1576]) | (layer4_outputs[3480]);
    assign layer5_outputs[365] = ~(layer4_outputs[1245]);
    assign layer5_outputs[366] = layer4_outputs[453];
    assign layer5_outputs[367] = ~(layer4_outputs[4922]);
    assign layer5_outputs[368] = layer4_outputs[1885];
    assign layer5_outputs[369] = (layer4_outputs[4713]) ^ (layer4_outputs[302]);
    assign layer5_outputs[370] = ~((layer4_outputs[593]) | (layer4_outputs[1280]));
    assign layer5_outputs[371] = (layer4_outputs[211]) ^ (layer4_outputs[185]);
    assign layer5_outputs[372] = ~(layer4_outputs[2872]);
    assign layer5_outputs[373] = ~(layer4_outputs[3701]);
    assign layer5_outputs[374] = ~(layer4_outputs[4884]) | (layer4_outputs[3782]);
    assign layer5_outputs[375] = ~((layer4_outputs[543]) | (layer4_outputs[4976]));
    assign layer5_outputs[376] = ~((layer4_outputs[2489]) ^ (layer4_outputs[901]));
    assign layer5_outputs[377] = ~(layer4_outputs[4743]) | (layer4_outputs[3801]);
    assign layer5_outputs[378] = (layer4_outputs[2357]) & ~(layer4_outputs[1919]);
    assign layer5_outputs[379] = layer4_outputs[2639];
    assign layer5_outputs[380] = ~(layer4_outputs[1511]);
    assign layer5_outputs[381] = ~(layer4_outputs[3731]) | (layer4_outputs[2481]);
    assign layer5_outputs[382] = layer4_outputs[3798];
    assign layer5_outputs[383] = ~(layer4_outputs[699]);
    assign layer5_outputs[384] = (layer4_outputs[4197]) & ~(layer4_outputs[2237]);
    assign layer5_outputs[385] = layer4_outputs[3052];
    assign layer5_outputs[386] = layer4_outputs[4561];
    assign layer5_outputs[387] = ~(layer4_outputs[165]) | (layer4_outputs[1653]);
    assign layer5_outputs[388] = (layer4_outputs[355]) & (layer4_outputs[2025]);
    assign layer5_outputs[389] = ~(layer4_outputs[2319]);
    assign layer5_outputs[390] = layer4_outputs[1755];
    assign layer5_outputs[391] = ~(layer4_outputs[18]) | (layer4_outputs[1963]);
    assign layer5_outputs[392] = ~(layer4_outputs[2748]);
    assign layer5_outputs[393] = layer4_outputs[2750];
    assign layer5_outputs[394] = ~((layer4_outputs[4978]) ^ (layer4_outputs[4706]));
    assign layer5_outputs[395] = ~(layer4_outputs[1276]) | (layer4_outputs[1882]);
    assign layer5_outputs[396] = layer4_outputs[2980];
    assign layer5_outputs[397] = (layer4_outputs[3697]) & (layer4_outputs[1703]);
    assign layer5_outputs[398] = ~(layer4_outputs[3744]);
    assign layer5_outputs[399] = layer4_outputs[717];
    assign layer5_outputs[400] = ~(layer4_outputs[4305]);
    assign layer5_outputs[401] = (layer4_outputs[2826]) & (layer4_outputs[4817]);
    assign layer5_outputs[402] = ~(layer4_outputs[4504]);
    assign layer5_outputs[403] = ~(layer4_outputs[2029]);
    assign layer5_outputs[404] = layer4_outputs[2050];
    assign layer5_outputs[405] = ~(layer4_outputs[533]);
    assign layer5_outputs[406] = (layer4_outputs[3826]) & ~(layer4_outputs[296]);
    assign layer5_outputs[407] = ~(layer4_outputs[259]);
    assign layer5_outputs[408] = layer4_outputs[1116];
    assign layer5_outputs[409] = ~((layer4_outputs[2752]) & (layer4_outputs[2523]));
    assign layer5_outputs[410] = layer4_outputs[3045];
    assign layer5_outputs[411] = ~(layer4_outputs[2554]);
    assign layer5_outputs[412] = layer4_outputs[317];
    assign layer5_outputs[413] = ~(layer4_outputs[2916]);
    assign layer5_outputs[414] = ~(layer4_outputs[3329]);
    assign layer5_outputs[415] = ~(layer4_outputs[4752]) | (layer4_outputs[3677]);
    assign layer5_outputs[416] = ~(layer4_outputs[1771]) | (layer4_outputs[960]);
    assign layer5_outputs[417] = layer4_outputs[2492];
    assign layer5_outputs[418] = (layer4_outputs[3364]) & (layer4_outputs[3506]);
    assign layer5_outputs[419] = (layer4_outputs[2339]) & ~(layer4_outputs[3677]);
    assign layer5_outputs[420] = (layer4_outputs[897]) ^ (layer4_outputs[1117]);
    assign layer5_outputs[421] = ~(layer4_outputs[837]);
    assign layer5_outputs[422] = ~((layer4_outputs[4764]) & (layer4_outputs[1500]));
    assign layer5_outputs[423] = ~(layer4_outputs[3389]);
    assign layer5_outputs[424] = ~(layer4_outputs[3037]) | (layer4_outputs[1371]);
    assign layer5_outputs[425] = ~((layer4_outputs[5100]) | (layer4_outputs[3869]));
    assign layer5_outputs[426] = ~(layer4_outputs[1601]);
    assign layer5_outputs[427] = ~(layer4_outputs[1655]);
    assign layer5_outputs[428] = layer4_outputs[3947];
    assign layer5_outputs[429] = ~((layer4_outputs[1643]) & (layer4_outputs[4724]));
    assign layer5_outputs[430] = ~((layer4_outputs[4237]) ^ (layer4_outputs[3785]));
    assign layer5_outputs[431] = layer4_outputs[121];
    assign layer5_outputs[432] = ~(layer4_outputs[466]);
    assign layer5_outputs[433] = layer4_outputs[4467];
    assign layer5_outputs[434] = ~(layer4_outputs[2997]);
    assign layer5_outputs[435] = ~(layer4_outputs[1417]);
    assign layer5_outputs[436] = layer4_outputs[2859];
    assign layer5_outputs[437] = layer4_outputs[2863];
    assign layer5_outputs[438] = (layer4_outputs[2030]) | (layer4_outputs[1102]);
    assign layer5_outputs[439] = (layer4_outputs[2213]) ^ (layer4_outputs[1166]);
    assign layer5_outputs[440] = 1'b1;
    assign layer5_outputs[441] = ~(layer4_outputs[566]);
    assign layer5_outputs[442] = (layer4_outputs[5056]) ^ (layer4_outputs[2544]);
    assign layer5_outputs[443] = (layer4_outputs[767]) & ~(layer4_outputs[4587]);
    assign layer5_outputs[444] = 1'b1;
    assign layer5_outputs[445] = layer4_outputs[568];
    assign layer5_outputs[446] = layer4_outputs[479];
    assign layer5_outputs[447] = (layer4_outputs[4377]) & (layer4_outputs[4417]);
    assign layer5_outputs[448] = (layer4_outputs[1715]) | (layer4_outputs[3612]);
    assign layer5_outputs[449] = 1'b1;
    assign layer5_outputs[450] = layer4_outputs[222];
    assign layer5_outputs[451] = (layer4_outputs[675]) & (layer4_outputs[392]);
    assign layer5_outputs[452] = ~(layer4_outputs[654]);
    assign layer5_outputs[453] = (layer4_outputs[1069]) ^ (layer4_outputs[1490]);
    assign layer5_outputs[454] = layer4_outputs[4198];
    assign layer5_outputs[455] = ~((layer4_outputs[4625]) ^ (layer4_outputs[3499]));
    assign layer5_outputs[456] = layer4_outputs[3087];
    assign layer5_outputs[457] = ~(layer4_outputs[4597]);
    assign layer5_outputs[458] = layer4_outputs[3973];
    assign layer5_outputs[459] = layer4_outputs[4720];
    assign layer5_outputs[460] = layer4_outputs[699];
    assign layer5_outputs[461] = layer4_outputs[341];
    assign layer5_outputs[462] = layer4_outputs[4453];
    assign layer5_outputs[463] = ~(layer4_outputs[625]);
    assign layer5_outputs[464] = layer4_outputs[3249];
    assign layer5_outputs[465] = layer4_outputs[3107];
    assign layer5_outputs[466] = ~(layer4_outputs[627]);
    assign layer5_outputs[467] = layer4_outputs[1656];
    assign layer5_outputs[468] = 1'b1;
    assign layer5_outputs[469] = (layer4_outputs[4850]) ^ (layer4_outputs[3072]);
    assign layer5_outputs[470] = 1'b1;
    assign layer5_outputs[471] = layer4_outputs[3498];
    assign layer5_outputs[472] = ~(layer4_outputs[378]);
    assign layer5_outputs[473] = ~(layer4_outputs[3626]);
    assign layer5_outputs[474] = ~((layer4_outputs[49]) | (layer4_outputs[4040]));
    assign layer5_outputs[475] = ~(layer4_outputs[2591]);
    assign layer5_outputs[476] = ~((layer4_outputs[14]) & (layer4_outputs[3399]));
    assign layer5_outputs[477] = (layer4_outputs[2648]) & ~(layer4_outputs[4986]);
    assign layer5_outputs[478] = layer4_outputs[2897];
    assign layer5_outputs[479] = layer4_outputs[4828];
    assign layer5_outputs[480] = (layer4_outputs[2624]) & (layer4_outputs[1238]);
    assign layer5_outputs[481] = layer4_outputs[409];
    assign layer5_outputs[482] = ~(layer4_outputs[484]) | (layer4_outputs[726]);
    assign layer5_outputs[483] = 1'b0;
    assign layer5_outputs[484] = (layer4_outputs[4390]) & ~(layer4_outputs[3508]);
    assign layer5_outputs[485] = ~(layer4_outputs[2587]);
    assign layer5_outputs[486] = ~(layer4_outputs[1539]);
    assign layer5_outputs[487] = ~((layer4_outputs[2159]) | (layer4_outputs[963]));
    assign layer5_outputs[488] = (layer4_outputs[440]) & ~(layer4_outputs[3058]);
    assign layer5_outputs[489] = layer4_outputs[2396];
    assign layer5_outputs[490] = (layer4_outputs[2625]) & (layer4_outputs[4741]);
    assign layer5_outputs[491] = ~((layer4_outputs[2581]) ^ (layer4_outputs[3456]));
    assign layer5_outputs[492] = (layer4_outputs[1274]) & (layer4_outputs[3060]);
    assign layer5_outputs[493] = ~((layer4_outputs[1383]) | (layer4_outputs[356]));
    assign layer5_outputs[494] = layer4_outputs[3658];
    assign layer5_outputs[495] = ~(layer4_outputs[3270]) | (layer4_outputs[1946]);
    assign layer5_outputs[496] = ~(layer4_outputs[1294]);
    assign layer5_outputs[497] = ~(layer4_outputs[1564]) | (layer4_outputs[4888]);
    assign layer5_outputs[498] = 1'b1;
    assign layer5_outputs[499] = layer4_outputs[4765];
    assign layer5_outputs[500] = ~((layer4_outputs[3254]) & (layer4_outputs[4239]));
    assign layer5_outputs[501] = ~((layer4_outputs[2959]) & (layer4_outputs[113]));
    assign layer5_outputs[502] = ~(layer4_outputs[2009]);
    assign layer5_outputs[503] = (layer4_outputs[2450]) & (layer4_outputs[4428]);
    assign layer5_outputs[504] = ~(layer4_outputs[1005]);
    assign layer5_outputs[505] = ~(layer4_outputs[3117]);
    assign layer5_outputs[506] = ~(layer4_outputs[3262]);
    assign layer5_outputs[507] = (layer4_outputs[1723]) ^ (layer4_outputs[4327]);
    assign layer5_outputs[508] = ~(layer4_outputs[4866]);
    assign layer5_outputs[509] = ~(layer4_outputs[2628]);
    assign layer5_outputs[510] = ~(layer4_outputs[4578]);
    assign layer5_outputs[511] = layer4_outputs[2534];
    assign layer5_outputs[512] = (layer4_outputs[4661]) ^ (layer4_outputs[3221]);
    assign layer5_outputs[513] = layer4_outputs[854];
    assign layer5_outputs[514] = ~(layer4_outputs[890]);
    assign layer5_outputs[515] = layer4_outputs[3533];
    assign layer5_outputs[516] = (layer4_outputs[3625]) ^ (layer4_outputs[76]);
    assign layer5_outputs[517] = (layer4_outputs[4543]) & ~(layer4_outputs[4619]);
    assign layer5_outputs[518] = ~(layer4_outputs[2518]);
    assign layer5_outputs[519] = (layer4_outputs[751]) | (layer4_outputs[3088]);
    assign layer5_outputs[520] = ~(layer4_outputs[5037]) | (layer4_outputs[208]);
    assign layer5_outputs[521] = (layer4_outputs[2986]) ^ (layer4_outputs[4234]);
    assign layer5_outputs[522] = ~(layer4_outputs[1905]) | (layer4_outputs[3717]);
    assign layer5_outputs[523] = layer4_outputs[862];
    assign layer5_outputs[524] = ~((layer4_outputs[3092]) ^ (layer4_outputs[1172]));
    assign layer5_outputs[525] = (layer4_outputs[906]) & (layer4_outputs[1227]);
    assign layer5_outputs[526] = ~((layer4_outputs[1666]) ^ (layer4_outputs[4010]));
    assign layer5_outputs[527] = (layer4_outputs[925]) | (layer4_outputs[1915]);
    assign layer5_outputs[528] = layer4_outputs[1470];
    assign layer5_outputs[529] = ~(layer4_outputs[3489]);
    assign layer5_outputs[530] = layer4_outputs[1464];
    assign layer5_outputs[531] = (layer4_outputs[968]) & (layer4_outputs[173]);
    assign layer5_outputs[532] = layer4_outputs[3944];
    assign layer5_outputs[533] = layer4_outputs[2482];
    assign layer5_outputs[534] = layer4_outputs[4398];
    assign layer5_outputs[535] = (layer4_outputs[5067]) & ~(layer4_outputs[4472]);
    assign layer5_outputs[536] = ~(layer4_outputs[5090]);
    assign layer5_outputs[537] = ~(layer4_outputs[3910]);
    assign layer5_outputs[538] = (layer4_outputs[2879]) ^ (layer4_outputs[1384]);
    assign layer5_outputs[539] = (layer4_outputs[3224]) & (layer4_outputs[3033]);
    assign layer5_outputs[540] = ~(layer4_outputs[1064]) | (layer4_outputs[1155]);
    assign layer5_outputs[541] = layer4_outputs[2595];
    assign layer5_outputs[542] = ~((layer4_outputs[3899]) ^ (layer4_outputs[3999]));
    assign layer5_outputs[543] = layer4_outputs[3990];
    assign layer5_outputs[544] = ~(layer4_outputs[1521]);
    assign layer5_outputs[545] = (layer4_outputs[4715]) ^ (layer4_outputs[727]);
    assign layer5_outputs[546] = ~(layer4_outputs[2191]);
    assign layer5_outputs[547] = ~(layer4_outputs[2661]) | (layer4_outputs[710]);
    assign layer5_outputs[548] = layer4_outputs[4452];
    assign layer5_outputs[549] = layer4_outputs[3290];
    assign layer5_outputs[550] = 1'b0;
    assign layer5_outputs[551] = ~(layer4_outputs[3681]);
    assign layer5_outputs[552] = layer4_outputs[4047];
    assign layer5_outputs[553] = ~(layer4_outputs[720]) | (layer4_outputs[3968]);
    assign layer5_outputs[554] = ~(layer4_outputs[4245]);
    assign layer5_outputs[555] = (layer4_outputs[4364]) & ~(layer4_outputs[2004]);
    assign layer5_outputs[556] = (layer4_outputs[3661]) & ~(layer4_outputs[132]);
    assign layer5_outputs[557] = (layer4_outputs[1691]) & ~(layer4_outputs[2157]);
    assign layer5_outputs[558] = 1'b1;
    assign layer5_outputs[559] = (layer4_outputs[547]) | (layer4_outputs[3958]);
    assign layer5_outputs[560] = ~((layer4_outputs[3255]) ^ (layer4_outputs[2982]));
    assign layer5_outputs[561] = ~((layer4_outputs[2707]) & (layer4_outputs[2925]));
    assign layer5_outputs[562] = ~(layer4_outputs[3269]);
    assign layer5_outputs[563] = ~((layer4_outputs[412]) ^ (layer4_outputs[515]));
    assign layer5_outputs[564] = ~(layer4_outputs[4159]);
    assign layer5_outputs[565] = layer4_outputs[3063];
    assign layer5_outputs[566] = ~(layer4_outputs[1534]);
    assign layer5_outputs[567] = ~(layer4_outputs[2399]);
    assign layer5_outputs[568] = (layer4_outputs[3921]) & ~(layer4_outputs[3006]);
    assign layer5_outputs[569] = (layer4_outputs[1096]) & (layer4_outputs[2468]);
    assign layer5_outputs[570] = ~(layer4_outputs[989]);
    assign layer5_outputs[571] = layer4_outputs[95];
    assign layer5_outputs[572] = 1'b1;
    assign layer5_outputs[573] = (layer4_outputs[4436]) & ~(layer4_outputs[1587]);
    assign layer5_outputs[574] = ~(layer4_outputs[1037]) | (layer4_outputs[3648]);
    assign layer5_outputs[575] = (layer4_outputs[2044]) & ~(layer4_outputs[4663]);
    assign layer5_outputs[576] = ~((layer4_outputs[2006]) ^ (layer4_outputs[2674]));
    assign layer5_outputs[577] = (layer4_outputs[158]) & (layer4_outputs[1129]);
    assign layer5_outputs[578] = layer4_outputs[4749];
    assign layer5_outputs[579] = ~(layer4_outputs[3208]);
    assign layer5_outputs[580] = layer4_outputs[927];
    assign layer5_outputs[581] = ~(layer4_outputs[942]);
    assign layer5_outputs[582] = (layer4_outputs[4819]) ^ (layer4_outputs[905]);
    assign layer5_outputs[583] = ~((layer4_outputs[2466]) | (layer4_outputs[3277]));
    assign layer5_outputs[584] = ~(layer4_outputs[853]);
    assign layer5_outputs[585] = ~(layer4_outputs[4900]);
    assign layer5_outputs[586] = ~(layer4_outputs[1935]);
    assign layer5_outputs[587] = (layer4_outputs[2517]) & ~(layer4_outputs[5098]);
    assign layer5_outputs[588] = layer4_outputs[152];
    assign layer5_outputs[589] = (layer4_outputs[4299]) ^ (layer4_outputs[4795]);
    assign layer5_outputs[590] = ~(layer4_outputs[2796]);
    assign layer5_outputs[591] = (layer4_outputs[3049]) & ~(layer4_outputs[310]);
    assign layer5_outputs[592] = ~(layer4_outputs[4833]);
    assign layer5_outputs[593] = (layer4_outputs[4604]) & (layer4_outputs[461]);
    assign layer5_outputs[594] = (layer4_outputs[3772]) & (layer4_outputs[799]);
    assign layer5_outputs[595] = ~((layer4_outputs[169]) | (layer4_outputs[3669]));
    assign layer5_outputs[596] = 1'b0;
    assign layer5_outputs[597] = ~(layer4_outputs[502]);
    assign layer5_outputs[598] = (layer4_outputs[86]) & ~(layer4_outputs[2715]);
    assign layer5_outputs[599] = (layer4_outputs[4659]) & ~(layer4_outputs[923]);
    assign layer5_outputs[600] = 1'b1;
    assign layer5_outputs[601] = layer4_outputs[3662];
    assign layer5_outputs[602] = ~(layer4_outputs[4258]);
    assign layer5_outputs[603] = (layer4_outputs[1275]) & ~(layer4_outputs[4432]);
    assign layer5_outputs[604] = ~(layer4_outputs[2207]);
    assign layer5_outputs[605] = ~(layer4_outputs[335]) | (layer4_outputs[4764]);
    assign layer5_outputs[606] = ~(layer4_outputs[1535]);
    assign layer5_outputs[607] = (layer4_outputs[3309]) & (layer4_outputs[1633]);
    assign layer5_outputs[608] = (layer4_outputs[4702]) & ~(layer4_outputs[4983]);
    assign layer5_outputs[609] = ~((layer4_outputs[1196]) & (layer4_outputs[2320]));
    assign layer5_outputs[610] = ~((layer4_outputs[4800]) & (layer4_outputs[2326]));
    assign layer5_outputs[611] = ~((layer4_outputs[4577]) ^ (layer4_outputs[1337]));
    assign layer5_outputs[612] = ~(layer4_outputs[4670]);
    assign layer5_outputs[613] = layer4_outputs[3216];
    assign layer5_outputs[614] = layer4_outputs[4496];
    assign layer5_outputs[615] = ~(layer4_outputs[3742]);
    assign layer5_outputs[616] = (layer4_outputs[4315]) | (layer4_outputs[1086]);
    assign layer5_outputs[617] = ~(layer4_outputs[1364]) | (layer4_outputs[2498]);
    assign layer5_outputs[618] = (layer4_outputs[3142]) ^ (layer4_outputs[3043]);
    assign layer5_outputs[619] = (layer4_outputs[3179]) ^ (layer4_outputs[2248]);
    assign layer5_outputs[620] = ~(layer4_outputs[4636]) | (layer4_outputs[572]);
    assign layer5_outputs[621] = (layer4_outputs[4294]) & (layer4_outputs[3866]);
    assign layer5_outputs[622] = ~(layer4_outputs[3409]);
    assign layer5_outputs[623] = ~(layer4_outputs[4847]) | (layer4_outputs[444]);
    assign layer5_outputs[624] = layer4_outputs[808];
    assign layer5_outputs[625] = ~((layer4_outputs[640]) & (layer4_outputs[2583]));
    assign layer5_outputs[626] = (layer4_outputs[2768]) & ~(layer4_outputs[1979]);
    assign layer5_outputs[627] = ~(layer4_outputs[4867]);
    assign layer5_outputs[628] = ~(layer4_outputs[3379]);
    assign layer5_outputs[629] = (layer4_outputs[2100]) & ~(layer4_outputs[2799]);
    assign layer5_outputs[630] = 1'b1;
    assign layer5_outputs[631] = (layer4_outputs[3616]) | (layer4_outputs[3749]);
    assign layer5_outputs[632] = layer4_outputs[3026];
    assign layer5_outputs[633] = ~(layer4_outputs[4664]);
    assign layer5_outputs[634] = (layer4_outputs[4266]) & ~(layer4_outputs[4296]);
    assign layer5_outputs[635] = (layer4_outputs[3377]) & ~(layer4_outputs[3629]);
    assign layer5_outputs[636] = ~((layer4_outputs[1672]) & (layer4_outputs[3830]));
    assign layer5_outputs[637] = ~((layer4_outputs[2781]) & (layer4_outputs[157]));
    assign layer5_outputs[638] = (layer4_outputs[4944]) & ~(layer4_outputs[3302]);
    assign layer5_outputs[639] = layer4_outputs[869];
    assign layer5_outputs[640] = layer4_outputs[1305];
    assign layer5_outputs[641] = (layer4_outputs[2418]) & ~(layer4_outputs[3864]);
    assign layer5_outputs[642] = (layer4_outputs[1454]) | (layer4_outputs[3574]);
    assign layer5_outputs[643] = (layer4_outputs[186]) & ~(layer4_outputs[1176]);
    assign layer5_outputs[644] = (layer4_outputs[2566]) & (layer4_outputs[2895]);
    assign layer5_outputs[645] = layer4_outputs[2269];
    assign layer5_outputs[646] = ~((layer4_outputs[2989]) & (layer4_outputs[89]));
    assign layer5_outputs[647] = ~((layer4_outputs[2920]) & (layer4_outputs[1]));
    assign layer5_outputs[648] = layer4_outputs[2149];
    assign layer5_outputs[649] = ~(layer4_outputs[1839]);
    assign layer5_outputs[650] = ~((layer4_outputs[365]) | (layer4_outputs[4691]));
    assign layer5_outputs[651] = ~((layer4_outputs[1047]) & (layer4_outputs[633]));
    assign layer5_outputs[652] = layer4_outputs[4425];
    assign layer5_outputs[653] = layer4_outputs[3907];
    assign layer5_outputs[654] = ~(layer4_outputs[4591]) | (layer4_outputs[3494]);
    assign layer5_outputs[655] = ~(layer4_outputs[3256]);
    assign layer5_outputs[656] = ~(layer4_outputs[45]);
    assign layer5_outputs[657] = 1'b0;
    assign layer5_outputs[658] = ~((layer4_outputs[4968]) & (layer4_outputs[4897]));
    assign layer5_outputs[659] = ~(layer4_outputs[437]) | (layer4_outputs[282]);
    assign layer5_outputs[660] = (layer4_outputs[3820]) ^ (layer4_outputs[396]);
    assign layer5_outputs[661] = (layer4_outputs[1173]) & (layer4_outputs[3370]);
    assign layer5_outputs[662] = (layer4_outputs[4107]) & (layer4_outputs[3993]);
    assign layer5_outputs[663] = layer4_outputs[4225];
    assign layer5_outputs[664] = ~(layer4_outputs[1586]);
    assign layer5_outputs[665] = layer4_outputs[1161];
    assign layer5_outputs[666] = 1'b1;
    assign layer5_outputs[667] = ~(layer4_outputs[1510]);
    assign layer5_outputs[668] = (layer4_outputs[2016]) & ~(layer4_outputs[759]);
    assign layer5_outputs[669] = 1'b1;
    assign layer5_outputs[670] = (layer4_outputs[2589]) & ~(layer4_outputs[2887]);
    assign layer5_outputs[671] = layer4_outputs[3310];
    assign layer5_outputs[672] = layer4_outputs[2129];
    assign layer5_outputs[673] = layer4_outputs[5064];
    assign layer5_outputs[674] = layer4_outputs[5111];
    assign layer5_outputs[675] = layer4_outputs[4415];
    assign layer5_outputs[676] = ~(layer4_outputs[2963]) | (layer4_outputs[909]);
    assign layer5_outputs[677] = (layer4_outputs[10]) & ~(layer4_outputs[562]);
    assign layer5_outputs[678] = ~(layer4_outputs[134]);
    assign layer5_outputs[679] = layer4_outputs[61];
    assign layer5_outputs[680] = ~(layer4_outputs[303]) | (layer4_outputs[4068]);
    assign layer5_outputs[681] = ~(layer4_outputs[3598]) | (layer4_outputs[1299]);
    assign layer5_outputs[682] = ~(layer4_outputs[2166]);
    assign layer5_outputs[683] = ~(layer4_outputs[535]);
    assign layer5_outputs[684] = ~((layer4_outputs[596]) & (layer4_outputs[1595]));
    assign layer5_outputs[685] = ~((layer4_outputs[3831]) | (layer4_outputs[763]));
    assign layer5_outputs[686] = ~(layer4_outputs[585]) | (layer4_outputs[1605]);
    assign layer5_outputs[687] = ~(layer4_outputs[830]);
    assign layer5_outputs[688] = (layer4_outputs[4987]) & (layer4_outputs[1995]);
    assign layer5_outputs[689] = (layer4_outputs[3717]) & ~(layer4_outputs[2847]);
    assign layer5_outputs[690] = ~((layer4_outputs[872]) | (layer4_outputs[3600]));
    assign layer5_outputs[691] = ~(layer4_outputs[2135]);
    assign layer5_outputs[692] = layer4_outputs[4922];
    assign layer5_outputs[693] = ~((layer4_outputs[4044]) & (layer4_outputs[3363]));
    assign layer5_outputs[694] = 1'b1;
    assign layer5_outputs[695] = layer4_outputs[3647];
    assign layer5_outputs[696] = ~(layer4_outputs[1762]);
    assign layer5_outputs[697] = layer4_outputs[1066];
    assign layer5_outputs[698] = layer4_outputs[4831];
    assign layer5_outputs[699] = layer4_outputs[2238];
    assign layer5_outputs[700] = (layer4_outputs[2106]) | (layer4_outputs[3034]);
    assign layer5_outputs[701] = ~((layer4_outputs[2983]) & (layer4_outputs[84]));
    assign layer5_outputs[702] = ~(layer4_outputs[2441]);
    assign layer5_outputs[703] = ~((layer4_outputs[4016]) | (layer4_outputs[1591]));
    assign layer5_outputs[704] = 1'b0;
    assign layer5_outputs[705] = ~(layer4_outputs[3656]) | (layer4_outputs[3102]);
    assign layer5_outputs[706] = ~((layer4_outputs[4566]) | (layer4_outputs[1401]));
    assign layer5_outputs[707] = layer4_outputs[916];
    assign layer5_outputs[708] = ~(layer4_outputs[4042]);
    assign layer5_outputs[709] = (layer4_outputs[2674]) & ~(layer4_outputs[4447]);
    assign layer5_outputs[710] = (layer4_outputs[4712]) & (layer4_outputs[4209]);
    assign layer5_outputs[711] = layer4_outputs[3958];
    assign layer5_outputs[712] = ~(layer4_outputs[312]);
    assign layer5_outputs[713] = ~(layer4_outputs[3741]);
    assign layer5_outputs[714] = layer4_outputs[3582];
    assign layer5_outputs[715] = ~((layer4_outputs[1038]) ^ (layer4_outputs[1866]));
    assign layer5_outputs[716] = (layer4_outputs[3659]) ^ (layer4_outputs[1868]);
    assign layer5_outputs[717] = (layer4_outputs[651]) ^ (layer4_outputs[1340]);
    assign layer5_outputs[718] = (layer4_outputs[1781]) ^ (layer4_outputs[4145]);
    assign layer5_outputs[719] = ~(layer4_outputs[2571]) | (layer4_outputs[1622]);
    assign layer5_outputs[720] = 1'b0;
    assign layer5_outputs[721] = (layer4_outputs[1988]) ^ (layer4_outputs[2378]);
    assign layer5_outputs[722] = ~(layer4_outputs[4081]) | (layer4_outputs[1421]);
    assign layer5_outputs[723] = 1'b0;
    assign layer5_outputs[724] = ~(layer4_outputs[1264]);
    assign layer5_outputs[725] = ~(layer4_outputs[217]);
    assign layer5_outputs[726] = ~(layer4_outputs[636]);
    assign layer5_outputs[727] = layer4_outputs[758];
    assign layer5_outputs[728] = (layer4_outputs[2803]) & ~(layer4_outputs[4600]);
    assign layer5_outputs[729] = (layer4_outputs[4820]) & ~(layer4_outputs[4754]);
    assign layer5_outputs[730] = ~(layer4_outputs[3259]);
    assign layer5_outputs[731] = (layer4_outputs[591]) & ~(layer4_outputs[490]);
    assign layer5_outputs[732] = ~(layer4_outputs[3303]);
    assign layer5_outputs[733] = ~(layer4_outputs[649]) | (layer4_outputs[4013]);
    assign layer5_outputs[734] = layer4_outputs[1104];
    assign layer5_outputs[735] = ~(layer4_outputs[1679]);
    assign layer5_outputs[736] = layer4_outputs[3131];
    assign layer5_outputs[737] = (layer4_outputs[2714]) & ~(layer4_outputs[1697]);
    assign layer5_outputs[738] = ~(layer4_outputs[3141]);
    assign layer5_outputs[739] = ~((layer4_outputs[1055]) | (layer4_outputs[3977]));
    assign layer5_outputs[740] = ~(layer4_outputs[1495]);
    assign layer5_outputs[741] = ~(layer4_outputs[3458]);
    assign layer5_outputs[742] = ~(layer4_outputs[1639]);
    assign layer5_outputs[743] = (layer4_outputs[1724]) ^ (layer4_outputs[412]);
    assign layer5_outputs[744] = (layer4_outputs[3540]) & ~(layer4_outputs[2355]);
    assign layer5_outputs[745] = 1'b0;
    assign layer5_outputs[746] = (layer4_outputs[3492]) & (layer4_outputs[3443]);
    assign layer5_outputs[747] = ~((layer4_outputs[4927]) ^ (layer4_outputs[3770]));
    assign layer5_outputs[748] = ~(layer4_outputs[2772]);
    assign layer5_outputs[749] = ~((layer4_outputs[3098]) ^ (layer4_outputs[3566]));
    assign layer5_outputs[750] = ~(layer4_outputs[4055]);
    assign layer5_outputs[751] = ~((layer4_outputs[3245]) & (layer4_outputs[4582]));
    assign layer5_outputs[752] = 1'b0;
    assign layer5_outputs[753] = layer4_outputs[5029];
    assign layer5_outputs[754] = layer4_outputs[1257];
    assign layer5_outputs[755] = layer4_outputs[3814];
    assign layer5_outputs[756] = ~(layer4_outputs[253]);
    assign layer5_outputs[757] = layer4_outputs[2331];
    assign layer5_outputs[758] = layer4_outputs[257];
    assign layer5_outputs[759] = layer4_outputs[185];
    assign layer5_outputs[760] = layer4_outputs[3758];
    assign layer5_outputs[761] = layer4_outputs[4611];
    assign layer5_outputs[762] = (layer4_outputs[3687]) & ~(layer4_outputs[3747]);
    assign layer5_outputs[763] = ~((layer4_outputs[3486]) & (layer4_outputs[3035]));
    assign layer5_outputs[764] = (layer4_outputs[149]) | (layer4_outputs[332]);
    assign layer5_outputs[765] = ~((layer4_outputs[4856]) | (layer4_outputs[4486]));
    assign layer5_outputs[766] = ~(layer4_outputs[1234]);
    assign layer5_outputs[767] = (layer4_outputs[813]) & (layer4_outputs[3132]);
    assign layer5_outputs[768] = (layer4_outputs[4745]) ^ (layer4_outputs[1267]);
    assign layer5_outputs[769] = (layer4_outputs[4317]) ^ (layer4_outputs[2645]);
    assign layer5_outputs[770] = (layer4_outputs[3040]) & ~(layer4_outputs[2503]);
    assign layer5_outputs[771] = ~(layer4_outputs[700]);
    assign layer5_outputs[772] = layer4_outputs[2363];
    assign layer5_outputs[773] = ~(layer4_outputs[3438]);
    assign layer5_outputs[774] = ~(layer4_outputs[1122]);
    assign layer5_outputs[775] = layer4_outputs[2788];
    assign layer5_outputs[776] = ~(layer4_outputs[3989]);
    assign layer5_outputs[777] = ~((layer4_outputs[2198]) & (layer4_outputs[3122]));
    assign layer5_outputs[778] = (layer4_outputs[737]) & ~(layer4_outputs[2382]);
    assign layer5_outputs[779] = (layer4_outputs[4098]) | (layer4_outputs[4644]);
    assign layer5_outputs[780] = (layer4_outputs[5048]) | (layer4_outputs[3759]);
    assign layer5_outputs[781] = layer4_outputs[2363];
    assign layer5_outputs[782] = 1'b0;
    assign layer5_outputs[783] = 1'b1;
    assign layer5_outputs[784] = 1'b1;
    assign layer5_outputs[785] = ~(layer4_outputs[3267]);
    assign layer5_outputs[786] = 1'b1;
    assign layer5_outputs[787] = layer4_outputs[1638];
    assign layer5_outputs[788] = layer4_outputs[2043];
    assign layer5_outputs[789] = layer4_outputs[3135];
    assign layer5_outputs[790] = ~((layer4_outputs[2758]) & (layer4_outputs[3243]));
    assign layer5_outputs[791] = ~(layer4_outputs[4759]);
    assign layer5_outputs[792] = ~(layer4_outputs[5035]);
    assign layer5_outputs[793] = 1'b1;
    assign layer5_outputs[794] = layer4_outputs[4613];
    assign layer5_outputs[795] = layer4_outputs[4332];
    assign layer5_outputs[796] = layer4_outputs[3825];
    assign layer5_outputs[797] = ~(layer4_outputs[2107]);
    assign layer5_outputs[798] = ~(layer4_outputs[424]) | (layer4_outputs[4056]);
    assign layer5_outputs[799] = ~((layer4_outputs[2353]) & (layer4_outputs[4015]));
    assign layer5_outputs[800] = layer4_outputs[871];
    assign layer5_outputs[801] = layer4_outputs[2347];
    assign layer5_outputs[802] = (layer4_outputs[5021]) ^ (layer4_outputs[2223]);
    assign layer5_outputs[803] = ~(layer4_outputs[5061]);
    assign layer5_outputs[804] = ~(layer4_outputs[4874]);
    assign layer5_outputs[805] = (layer4_outputs[4575]) ^ (layer4_outputs[3241]);
    assign layer5_outputs[806] = ~((layer4_outputs[689]) | (layer4_outputs[1473]));
    assign layer5_outputs[807] = (layer4_outputs[2041]) & ~(layer4_outputs[3204]);
    assign layer5_outputs[808] = ~(layer4_outputs[3768]);
    assign layer5_outputs[809] = ~(layer4_outputs[4959]) | (layer4_outputs[2770]);
    assign layer5_outputs[810] = layer4_outputs[631];
    assign layer5_outputs[811] = layer4_outputs[1931];
    assign layer5_outputs[812] = 1'b0;
    assign layer5_outputs[813] = layer4_outputs[437];
    assign layer5_outputs[814] = layer4_outputs[1541];
    assign layer5_outputs[815] = ~((layer4_outputs[474]) | (layer4_outputs[1402]));
    assign layer5_outputs[816] = ~(layer4_outputs[248]);
    assign layer5_outputs[817] = layer4_outputs[2481];
    assign layer5_outputs[818] = layer4_outputs[4557];
    assign layer5_outputs[819] = 1'b0;
    assign layer5_outputs[820] = (layer4_outputs[337]) | (layer4_outputs[3190]);
    assign layer5_outputs[821] = ~((layer4_outputs[5082]) | (layer4_outputs[461]));
    assign layer5_outputs[822] = ~(layer4_outputs[2435]);
    assign layer5_outputs[823] = ~((layer4_outputs[4757]) | (layer4_outputs[2855]));
    assign layer5_outputs[824] = ~(layer4_outputs[932]) | (layer4_outputs[658]);
    assign layer5_outputs[825] = ~((layer4_outputs[2434]) & (layer4_outputs[3250]));
    assign layer5_outputs[826] = layer4_outputs[4636];
    assign layer5_outputs[827] = ~((layer4_outputs[2949]) | (layer4_outputs[855]));
    assign layer5_outputs[828] = ~(layer4_outputs[3342]);
    assign layer5_outputs[829] = ~(layer4_outputs[480]);
    assign layer5_outputs[830] = layer4_outputs[4666];
    assign layer5_outputs[831] = (layer4_outputs[3247]) & ~(layer4_outputs[1008]);
    assign layer5_outputs[832] = (layer4_outputs[2107]) & (layer4_outputs[872]);
    assign layer5_outputs[833] = ~(layer4_outputs[352]) | (layer4_outputs[2065]);
    assign layer5_outputs[834] = ~(layer4_outputs[4343]);
    assign layer5_outputs[835] = ~(layer4_outputs[5103]);
    assign layer5_outputs[836] = (layer4_outputs[1648]) ^ (layer4_outputs[1881]);
    assign layer5_outputs[837] = ~(layer4_outputs[4726]);
    assign layer5_outputs[838] = layer4_outputs[4881];
    assign layer5_outputs[839] = ~(layer4_outputs[3555]);
    assign layer5_outputs[840] = layer4_outputs[183];
    assign layer5_outputs[841] = ~((layer4_outputs[2420]) & (layer4_outputs[743]));
    assign layer5_outputs[842] = ~(layer4_outputs[4729]);
    assign layer5_outputs[843] = ~(layer4_outputs[4730]) | (layer4_outputs[4116]);
    assign layer5_outputs[844] = ~(layer4_outputs[1306]);
    assign layer5_outputs[845] = 1'b0;
    assign layer5_outputs[846] = ~(layer4_outputs[4921]);
    assign layer5_outputs[847] = ~(layer4_outputs[5031]);
    assign layer5_outputs[848] = (layer4_outputs[4681]) & ~(layer4_outputs[911]);
    assign layer5_outputs[849] = 1'b1;
    assign layer5_outputs[850] = ~(layer4_outputs[3105]) | (layer4_outputs[4603]);
    assign layer5_outputs[851] = (layer4_outputs[2836]) & ~(layer4_outputs[3281]);
    assign layer5_outputs[852] = ~((layer4_outputs[2423]) ^ (layer4_outputs[2325]));
    assign layer5_outputs[853] = (layer4_outputs[2424]) & ~(layer4_outputs[3923]);
    assign layer5_outputs[854] = ~(layer4_outputs[4107]);
    assign layer5_outputs[855] = layer4_outputs[1022];
    assign layer5_outputs[856] = (layer4_outputs[2564]) & ~(layer4_outputs[252]);
    assign layer5_outputs[857] = 1'b0;
    assign layer5_outputs[858] = ~(layer4_outputs[2556]);
    assign layer5_outputs[859] = ~((layer4_outputs[39]) & (layer4_outputs[1898]));
    assign layer5_outputs[860] = (layer4_outputs[76]) | (layer4_outputs[4947]);
    assign layer5_outputs[861] = ~((layer4_outputs[4104]) ^ (layer4_outputs[1562]));
    assign layer5_outputs[862] = (layer4_outputs[2536]) | (layer4_outputs[3976]);
    assign layer5_outputs[863] = (layer4_outputs[3352]) & (layer4_outputs[806]);
    assign layer5_outputs[864] = ~(layer4_outputs[5082]);
    assign layer5_outputs[865] = ~((layer4_outputs[1540]) | (layer4_outputs[3797]));
    assign layer5_outputs[866] = ~(layer4_outputs[1081]);
    assign layer5_outputs[867] = 1'b1;
    assign layer5_outputs[868] = (layer4_outputs[524]) & ~(layer4_outputs[4697]);
    assign layer5_outputs[869] = ~(layer4_outputs[3421]);
    assign layer5_outputs[870] = ~(layer4_outputs[2045]);
    assign layer5_outputs[871] = layer4_outputs[99];
    assign layer5_outputs[872] = ~((layer4_outputs[324]) | (layer4_outputs[4033]));
    assign layer5_outputs[873] = ~(layer4_outputs[2104]);
    assign layer5_outputs[874] = layer4_outputs[2771];
    assign layer5_outputs[875] = ~((layer4_outputs[3004]) & (layer4_outputs[1379]));
    assign layer5_outputs[876] = layer4_outputs[1765];
    assign layer5_outputs[877] = ~(layer4_outputs[141]);
    assign layer5_outputs[878] = layer4_outputs[3187];
    assign layer5_outputs[879] = layer4_outputs[540];
    assign layer5_outputs[880] = ~((layer4_outputs[3714]) ^ (layer4_outputs[3832]));
    assign layer5_outputs[881] = ~(layer4_outputs[2377]);
    assign layer5_outputs[882] = 1'b0;
    assign layer5_outputs[883] = ~(layer4_outputs[442]);
    assign layer5_outputs[884] = (layer4_outputs[847]) & (layer4_outputs[2553]);
    assign layer5_outputs[885] = ~(layer4_outputs[4907]);
    assign layer5_outputs[886] = 1'b0;
    assign layer5_outputs[887] = ~(layer4_outputs[4252]);
    assign layer5_outputs[888] = ~(layer4_outputs[3610]);
    assign layer5_outputs[889] = ~(layer4_outputs[4338]);
    assign layer5_outputs[890] = (layer4_outputs[349]) ^ (layer4_outputs[3515]);
    assign layer5_outputs[891] = (layer4_outputs[2834]) | (layer4_outputs[3963]);
    assign layer5_outputs[892] = (layer4_outputs[3286]) & ~(layer4_outputs[770]);
    assign layer5_outputs[893] = (layer4_outputs[200]) & ~(layer4_outputs[4240]);
    assign layer5_outputs[894] = ~((layer4_outputs[4206]) | (layer4_outputs[1496]));
    assign layer5_outputs[895] = (layer4_outputs[4460]) & ~(layer4_outputs[1177]);
    assign layer5_outputs[896] = ~((layer4_outputs[4761]) | (layer4_outputs[4792]));
    assign layer5_outputs[897] = (layer4_outputs[3634]) ^ (layer4_outputs[676]);
    assign layer5_outputs[898] = (layer4_outputs[604]) | (layer4_outputs[363]);
    assign layer5_outputs[899] = layer4_outputs[1543];
    assign layer5_outputs[900] = ~((layer4_outputs[3589]) | (layer4_outputs[1917]));
    assign layer5_outputs[901] = ~(layer4_outputs[1292]);
    assign layer5_outputs[902] = ~((layer4_outputs[4980]) & (layer4_outputs[2475]));
    assign layer5_outputs[903] = layer4_outputs[222];
    assign layer5_outputs[904] = layer4_outputs[4642];
    assign layer5_outputs[905] = layer4_outputs[723];
    assign layer5_outputs[906] = layer4_outputs[951];
    assign layer5_outputs[907] = (layer4_outputs[4038]) | (layer4_outputs[4940]);
    assign layer5_outputs[908] = layer4_outputs[2965];
    assign layer5_outputs[909] = layer4_outputs[2379];
    assign layer5_outputs[910] = layer4_outputs[488];
    assign layer5_outputs[911] = layer4_outputs[4703];
    assign layer5_outputs[912] = layer4_outputs[1154];
    assign layer5_outputs[913] = (layer4_outputs[921]) & ~(layer4_outputs[3347]);
    assign layer5_outputs[914] = (layer4_outputs[2386]) & ~(layer4_outputs[2511]);
    assign layer5_outputs[915] = ~(layer4_outputs[64]);
    assign layer5_outputs[916] = (layer4_outputs[4385]) & (layer4_outputs[2831]);
    assign layer5_outputs[917] = (layer4_outputs[3487]) & ~(layer4_outputs[3056]);
    assign layer5_outputs[918] = layer4_outputs[4399];
    assign layer5_outputs[919] = (layer4_outputs[3019]) & (layer4_outputs[3191]);
    assign layer5_outputs[920] = layer4_outputs[4996];
    assign layer5_outputs[921] = (layer4_outputs[1534]) & (layer4_outputs[3186]);
    assign layer5_outputs[922] = ~(layer4_outputs[477]);
    assign layer5_outputs[923] = (layer4_outputs[774]) | (layer4_outputs[3499]);
    assign layer5_outputs[924] = ~((layer4_outputs[3983]) & (layer4_outputs[4508]));
    assign layer5_outputs[925] = ~(layer4_outputs[1187]);
    assign layer5_outputs[926] = ~((layer4_outputs[3395]) ^ (layer4_outputs[2620]));
    assign layer5_outputs[927] = (layer4_outputs[2656]) & (layer4_outputs[1518]);
    assign layer5_outputs[928] = layer4_outputs[248];
    assign layer5_outputs[929] = (layer4_outputs[5061]) ^ (layer4_outputs[3016]);
    assign layer5_outputs[930] = ~(layer4_outputs[786]);
    assign layer5_outputs[931] = ~(layer4_outputs[1019]);
    assign layer5_outputs[932] = layer4_outputs[586];
    assign layer5_outputs[933] = layer4_outputs[2990];
    assign layer5_outputs[934] = layer4_outputs[4562];
    assign layer5_outputs[935] = layer4_outputs[1350];
    assign layer5_outputs[936] = (layer4_outputs[203]) & ~(layer4_outputs[2699]);
    assign layer5_outputs[937] = layer4_outputs[3019];
    assign layer5_outputs[938] = ~(layer4_outputs[4482]);
    assign layer5_outputs[939] = ~(layer4_outputs[4521]);
    assign layer5_outputs[940] = 1'b1;
    assign layer5_outputs[941] = layer4_outputs[1223];
    assign layer5_outputs[942] = layer4_outputs[5019];
    assign layer5_outputs[943] = ~((layer4_outputs[903]) | (layer4_outputs[2908]));
    assign layer5_outputs[944] = layer4_outputs[607];
    assign layer5_outputs[945] = ~((layer4_outputs[1469]) | (layer4_outputs[5024]));
    assign layer5_outputs[946] = ~(layer4_outputs[1717]);
    assign layer5_outputs[947] = layer4_outputs[4223];
    assign layer5_outputs[948] = ~(layer4_outputs[3772]);
    assign layer5_outputs[949] = ~(layer4_outputs[2458]) | (layer4_outputs[386]);
    assign layer5_outputs[950] = ~(layer4_outputs[849]) | (layer4_outputs[1113]);
    assign layer5_outputs[951] = layer4_outputs[1623];
    assign layer5_outputs[952] = 1'b1;
    assign layer5_outputs[953] = 1'b1;
    assign layer5_outputs[954] = (layer4_outputs[1447]) ^ (layer4_outputs[2895]);
    assign layer5_outputs[955] = layer4_outputs[1700];
    assign layer5_outputs[956] = ~(layer4_outputs[1450]);
    assign layer5_outputs[957] = layer4_outputs[2313];
    assign layer5_outputs[958] = ~(layer4_outputs[2503]);
    assign layer5_outputs[959] = layer4_outputs[730];
    assign layer5_outputs[960] = (layer4_outputs[4280]) & ~(layer4_outputs[2727]);
    assign layer5_outputs[961] = ~((layer4_outputs[4756]) & (layer4_outputs[3852]));
    assign layer5_outputs[962] = layer4_outputs[2832];
    assign layer5_outputs[963] = ~(layer4_outputs[1409]);
    assign layer5_outputs[964] = ~(layer4_outputs[4797]);
    assign layer5_outputs[965] = (layer4_outputs[802]) & ~(layer4_outputs[4761]);
    assign layer5_outputs[966] = ~((layer4_outputs[4202]) ^ (layer4_outputs[3232]));
    assign layer5_outputs[967] = ~(layer4_outputs[1958]) | (layer4_outputs[1747]);
    assign layer5_outputs[968] = layer4_outputs[533];
    assign layer5_outputs[969] = (layer4_outputs[1444]) ^ (layer4_outputs[4558]);
    assign layer5_outputs[970] = layer4_outputs[2188];
    assign layer5_outputs[971] = ~(layer4_outputs[3333]);
    assign layer5_outputs[972] = ~((layer4_outputs[2577]) & (layer4_outputs[1145]));
    assign layer5_outputs[973] = 1'b0;
    assign layer5_outputs[974] = 1'b1;
    assign layer5_outputs[975] = (layer4_outputs[3275]) & ~(layer4_outputs[1226]);
    assign layer5_outputs[976] = ~(layer4_outputs[4974]);
    assign layer5_outputs[977] = ~(layer4_outputs[4395]);
    assign layer5_outputs[978] = ~((layer4_outputs[2466]) | (layer4_outputs[4270]));
    assign layer5_outputs[979] = layer4_outputs[1289];
    assign layer5_outputs[980] = (layer4_outputs[605]) ^ (layer4_outputs[3465]);
    assign layer5_outputs[981] = ~(layer4_outputs[1162]) | (layer4_outputs[1448]);
    assign layer5_outputs[982] = 1'b1;
    assign layer5_outputs[983] = (layer4_outputs[3379]) ^ (layer4_outputs[1389]);
    assign layer5_outputs[984] = (layer4_outputs[2380]) | (layer4_outputs[1705]);
    assign layer5_outputs[985] = layer4_outputs[1452];
    assign layer5_outputs[986] = layer4_outputs[927];
    assign layer5_outputs[987] = (layer4_outputs[3361]) | (layer4_outputs[1767]);
    assign layer5_outputs[988] = layer4_outputs[4162];
    assign layer5_outputs[989] = ~(layer4_outputs[4917]);
    assign layer5_outputs[990] = (layer4_outputs[4457]) | (layer4_outputs[3301]);
    assign layer5_outputs[991] = layer4_outputs[1987];
    assign layer5_outputs[992] = ~(layer4_outputs[1416]);
    assign layer5_outputs[993] = ~(layer4_outputs[1714]);
    assign layer5_outputs[994] = ~(layer4_outputs[4245]);
    assign layer5_outputs[995] = layer4_outputs[1956];
    assign layer5_outputs[996] = ~(layer4_outputs[485]);
    assign layer5_outputs[997] = layer4_outputs[659];
    assign layer5_outputs[998] = ~(layer4_outputs[1106]);
    assign layer5_outputs[999] = ~(layer4_outputs[4931]);
    assign layer5_outputs[1000] = (layer4_outputs[4277]) | (layer4_outputs[1066]);
    assign layer5_outputs[1001] = ~(layer4_outputs[1592]) | (layer4_outputs[3152]);
    assign layer5_outputs[1002] = layer4_outputs[2328];
    assign layer5_outputs[1003] = (layer4_outputs[3231]) | (layer4_outputs[2925]);
    assign layer5_outputs[1004] = ~((layer4_outputs[1397]) & (layer4_outputs[5020]));
    assign layer5_outputs[1005] = layer4_outputs[641];
    assign layer5_outputs[1006] = ~(layer4_outputs[1465]);
    assign layer5_outputs[1007] = ~(layer4_outputs[465]);
    assign layer5_outputs[1008] = layer4_outputs[929];
    assign layer5_outputs[1009] = layer4_outputs[739];
    assign layer5_outputs[1010] = ~(layer4_outputs[1222]) | (layer4_outputs[3580]);
    assign layer5_outputs[1011] = (layer4_outputs[2086]) & (layer4_outputs[5074]);
    assign layer5_outputs[1012] = ~((layer4_outputs[1099]) | (layer4_outputs[1799]));
    assign layer5_outputs[1013] = ~(layer4_outputs[1213]);
    assign layer5_outputs[1014] = 1'b0;
    assign layer5_outputs[1015] = ~((layer4_outputs[931]) ^ (layer4_outputs[4176]));
    assign layer5_outputs[1016] = layer4_outputs[680];
    assign layer5_outputs[1017] = 1'b0;
    assign layer5_outputs[1018] = layer4_outputs[3657];
    assign layer5_outputs[1019] = (layer4_outputs[3097]) & ~(layer4_outputs[1270]);
    assign layer5_outputs[1020] = (layer4_outputs[1325]) | (layer4_outputs[277]);
    assign layer5_outputs[1021] = ~(layer4_outputs[3284]);
    assign layer5_outputs[1022] = layer4_outputs[3786];
    assign layer5_outputs[1023] = layer4_outputs[1713];
    assign layer5_outputs[1024] = layer4_outputs[2537];
    assign layer5_outputs[1025] = ~(layer4_outputs[2459]) | (layer4_outputs[2824]);
    assign layer5_outputs[1026] = ~(layer4_outputs[1233]);
    assign layer5_outputs[1027] = ~((layer4_outputs[3289]) ^ (layer4_outputs[1328]));
    assign layer5_outputs[1028] = layer4_outputs[3824];
    assign layer5_outputs[1029] = ~((layer4_outputs[3156]) & (layer4_outputs[2698]));
    assign layer5_outputs[1030] = ~(layer4_outputs[749]);
    assign layer5_outputs[1031] = ~(layer4_outputs[4309]) | (layer4_outputs[303]);
    assign layer5_outputs[1032] = layer4_outputs[3902];
    assign layer5_outputs[1033] = ~(layer4_outputs[518]);
    assign layer5_outputs[1034] = layer4_outputs[705];
    assign layer5_outputs[1035] = (layer4_outputs[3963]) & ~(layer4_outputs[1968]);
    assign layer5_outputs[1036] = ~(layer4_outputs[1584]);
    assign layer5_outputs[1037] = ~(layer4_outputs[4609]) | (layer4_outputs[4810]);
    assign layer5_outputs[1038] = ~(layer4_outputs[2637]);
    assign layer5_outputs[1039] = (layer4_outputs[3775]) | (layer4_outputs[2726]);
    assign layer5_outputs[1040] = layer4_outputs[2773];
    assign layer5_outputs[1041] = (layer4_outputs[366]) & (layer4_outputs[2566]);
    assign layer5_outputs[1042] = 1'b1;
    assign layer5_outputs[1043] = ~(layer4_outputs[1489]);
    assign layer5_outputs[1044] = layer4_outputs[717];
    assign layer5_outputs[1045] = layer4_outputs[4482];
    assign layer5_outputs[1046] = layer4_outputs[2046];
    assign layer5_outputs[1047] = layer4_outputs[1405];
    assign layer5_outputs[1048] = ~(layer4_outputs[788]) | (layer4_outputs[1664]);
    assign layer5_outputs[1049] = layer4_outputs[2785];
    assign layer5_outputs[1050] = (layer4_outputs[838]) & (layer4_outputs[1812]);
    assign layer5_outputs[1051] = layer4_outputs[1662];
    assign layer5_outputs[1052] = ~(layer4_outputs[2661]);
    assign layer5_outputs[1053] = ~(layer4_outputs[733]);
    assign layer5_outputs[1054] = layer4_outputs[3479];
    assign layer5_outputs[1055] = layer4_outputs[684];
    assign layer5_outputs[1056] = (layer4_outputs[1329]) & ~(layer4_outputs[2237]);
    assign layer5_outputs[1057] = (layer4_outputs[3610]) ^ (layer4_outputs[4644]);
    assign layer5_outputs[1058] = (layer4_outputs[3195]) & ~(layer4_outputs[4256]);
    assign layer5_outputs[1059] = layer4_outputs[3469];
    assign layer5_outputs[1060] = (layer4_outputs[1254]) ^ (layer4_outputs[452]);
    assign layer5_outputs[1061] = ~((layer4_outputs[4034]) | (layer4_outputs[1803]));
    assign layer5_outputs[1062] = ~(layer4_outputs[1876]);
    assign layer5_outputs[1063] = ~(layer4_outputs[1269]);
    assign layer5_outputs[1064] = ~(layer4_outputs[2839]);
    assign layer5_outputs[1065] = ~((layer4_outputs[2502]) ^ (layer4_outputs[686]));
    assign layer5_outputs[1066] = ~(layer4_outputs[97]) | (layer4_outputs[4187]);
    assign layer5_outputs[1067] = (layer4_outputs[1523]) | (layer4_outputs[1652]);
    assign layer5_outputs[1068] = ~((layer4_outputs[3910]) ^ (layer4_outputs[2415]));
    assign layer5_outputs[1069] = ~(layer4_outputs[1415]);
    assign layer5_outputs[1070] = (layer4_outputs[4393]) & ~(layer4_outputs[3653]);
    assign layer5_outputs[1071] = 1'b1;
    assign layer5_outputs[1072] = (layer4_outputs[1872]) ^ (layer4_outputs[2672]);
    assign layer5_outputs[1073] = layer4_outputs[1888];
    assign layer5_outputs[1074] = ~(layer4_outputs[3289]);
    assign layer5_outputs[1075] = (layer4_outputs[4166]) & (layer4_outputs[4139]);
    assign layer5_outputs[1076] = ~(layer4_outputs[3290]);
    assign layer5_outputs[1077] = ~(layer4_outputs[1730]);
    assign layer5_outputs[1078] = layer4_outputs[1017];
    assign layer5_outputs[1079] = layer4_outputs[4459];
    assign layer5_outputs[1080] = layer4_outputs[3346];
    assign layer5_outputs[1081] = layer4_outputs[372];
    assign layer5_outputs[1082] = (layer4_outputs[2815]) & ~(layer4_outputs[3230]);
    assign layer5_outputs[1083] = (layer4_outputs[2922]) & (layer4_outputs[2998]);
    assign layer5_outputs[1084] = (layer4_outputs[1480]) ^ (layer4_outputs[2904]);
    assign layer5_outputs[1085] = ~(layer4_outputs[1917]);
    assign layer5_outputs[1086] = layer4_outputs[1069];
    assign layer5_outputs[1087] = ~(layer4_outputs[3351]);
    assign layer5_outputs[1088] = layer4_outputs[421];
    assign layer5_outputs[1089] = (layer4_outputs[1548]) & ~(layer4_outputs[2528]);
    assign layer5_outputs[1090] = ~((layer4_outputs[4861]) | (layer4_outputs[2162]));
    assign layer5_outputs[1091] = layer4_outputs[3729];
    assign layer5_outputs[1092] = layer4_outputs[1804];
    assign layer5_outputs[1093] = ~(layer4_outputs[4136]) | (layer4_outputs[491]);
    assign layer5_outputs[1094] = ~(layer4_outputs[159]) | (layer4_outputs[4190]);
    assign layer5_outputs[1095] = ~(layer4_outputs[1686]);
    assign layer5_outputs[1096] = layer4_outputs[3484];
    assign layer5_outputs[1097] = ~(layer4_outputs[1973]);
    assign layer5_outputs[1098] = layer4_outputs[4939];
    assign layer5_outputs[1099] = ~((layer4_outputs[3195]) ^ (layer4_outputs[1891]));
    assign layer5_outputs[1100] = ~(layer4_outputs[851]) | (layer4_outputs[4559]);
    assign layer5_outputs[1101] = ~(layer4_outputs[4119]);
    assign layer5_outputs[1102] = ~((layer4_outputs[2508]) | (layer4_outputs[3192]));
    assign layer5_outputs[1103] = (layer4_outputs[3818]) & ~(layer4_outputs[4704]);
    assign layer5_outputs[1104] = ~((layer4_outputs[4771]) ^ (layer4_outputs[2557]));
    assign layer5_outputs[1105] = (layer4_outputs[4412]) & ~(layer4_outputs[447]);
    assign layer5_outputs[1106] = (layer4_outputs[5007]) & ~(layer4_outputs[2974]);
    assign layer5_outputs[1107] = ~((layer4_outputs[4493]) | (layer4_outputs[991]));
    assign layer5_outputs[1108] = (layer4_outputs[4298]) ^ (layer4_outputs[1195]);
    assign layer5_outputs[1109] = (layer4_outputs[3184]) | (layer4_outputs[3961]);
    assign layer5_outputs[1110] = (layer4_outputs[2227]) ^ (layer4_outputs[1481]);
    assign layer5_outputs[1111] = 1'b0;
    assign layer5_outputs[1112] = (layer4_outputs[2170]) & ~(layer4_outputs[3082]);
    assign layer5_outputs[1113] = 1'b1;
    assign layer5_outputs[1114] = layer4_outputs[81];
    assign layer5_outputs[1115] = ~((layer4_outputs[675]) | (layer4_outputs[316]));
    assign layer5_outputs[1116] = ~((layer4_outputs[5108]) & (layer4_outputs[3298]));
    assign layer5_outputs[1117] = 1'b1;
    assign layer5_outputs[1118] = ~((layer4_outputs[982]) & (layer4_outputs[4945]));
    assign layer5_outputs[1119] = ~(layer4_outputs[4321]);
    assign layer5_outputs[1120] = 1'b1;
    assign layer5_outputs[1121] = (layer4_outputs[980]) ^ (layer4_outputs[3060]);
    assign layer5_outputs[1122] = ~(layer4_outputs[1944]);
    assign layer5_outputs[1123] = layer4_outputs[416];
    assign layer5_outputs[1124] = layer4_outputs[4918];
    assign layer5_outputs[1125] = ~(layer4_outputs[2633]);
    assign layer5_outputs[1126] = (layer4_outputs[2606]) ^ (layer4_outputs[4635]);
    assign layer5_outputs[1127] = ~((layer4_outputs[3997]) | (layer4_outputs[3812]));
    assign layer5_outputs[1128] = ~(layer4_outputs[4260]) | (layer4_outputs[4564]);
    assign layer5_outputs[1129] = 1'b0;
    assign layer5_outputs[1130] = ~(layer4_outputs[1462]) | (layer4_outputs[4742]);
    assign layer5_outputs[1131] = ~(layer4_outputs[4033]) | (layer4_outputs[4640]);
    assign layer5_outputs[1132] = ~(layer4_outputs[233]) | (layer4_outputs[757]);
    assign layer5_outputs[1133] = layer4_outputs[1199];
    assign layer5_outputs[1134] = layer4_outputs[536];
    assign layer5_outputs[1135] = ~(layer4_outputs[4806]) | (layer4_outputs[4545]);
    assign layer5_outputs[1136] = layer4_outputs[394];
    assign layer5_outputs[1137] = ~(layer4_outputs[2435]);
    assign layer5_outputs[1138] = (layer4_outputs[3205]) ^ (layer4_outputs[3030]);
    assign layer5_outputs[1139] = ~((layer4_outputs[1482]) & (layer4_outputs[164]));
    assign layer5_outputs[1140] = ~(layer4_outputs[1003]) | (layer4_outputs[577]);
    assign layer5_outputs[1141] = (layer4_outputs[3309]) | (layer4_outputs[1036]);
    assign layer5_outputs[1142] = (layer4_outputs[3957]) & (layer4_outputs[300]);
    assign layer5_outputs[1143] = 1'b1;
    assign layer5_outputs[1144] = ~(layer4_outputs[4083]) | (layer4_outputs[4145]);
    assign layer5_outputs[1145] = (layer4_outputs[3489]) | (layer4_outputs[362]);
    assign layer5_outputs[1146] = (layer4_outputs[3860]) & ~(layer4_outputs[3086]);
    assign layer5_outputs[1147] = layer4_outputs[1640];
    assign layer5_outputs[1148] = layer4_outputs[4391];
    assign layer5_outputs[1149] = layer4_outputs[1434];
    assign layer5_outputs[1150] = layer4_outputs[3582];
    assign layer5_outputs[1151] = (layer4_outputs[3313]) | (layer4_outputs[2425]);
    assign layer5_outputs[1152] = ~(layer4_outputs[4360]);
    assign layer5_outputs[1153] = (layer4_outputs[3497]) & ~(layer4_outputs[4499]);
    assign layer5_outputs[1154] = ~(layer4_outputs[44]);
    assign layer5_outputs[1155] = ~(layer4_outputs[2965]);
    assign layer5_outputs[1156] = ~(layer4_outputs[4902]) | (layer4_outputs[1126]);
    assign layer5_outputs[1157] = ~(layer4_outputs[590]);
    assign layer5_outputs[1158] = ~(layer4_outputs[858]) | (layer4_outputs[970]);
    assign layer5_outputs[1159] = layer4_outputs[4352];
    assign layer5_outputs[1160] = layer4_outputs[756];
    assign layer5_outputs[1161] = (layer4_outputs[5007]) & (layer4_outputs[3163]);
    assign layer5_outputs[1162] = layer4_outputs[2263];
    assign layer5_outputs[1163] = layer4_outputs[2287];
    assign layer5_outputs[1164] = ~(layer4_outputs[297]);
    assign layer5_outputs[1165] = ~(layer4_outputs[2473]);
    assign layer5_outputs[1166] = (layer4_outputs[2278]) & ~(layer4_outputs[2548]);
    assign layer5_outputs[1167] = ~(layer4_outputs[3802]);
    assign layer5_outputs[1168] = ~(layer4_outputs[4091]);
    assign layer5_outputs[1169] = (layer4_outputs[1227]) & (layer4_outputs[4865]);
    assign layer5_outputs[1170] = ~(layer4_outputs[1945]);
    assign layer5_outputs[1171] = ~((layer4_outputs[3321]) & (layer4_outputs[1862]));
    assign layer5_outputs[1172] = 1'b1;
    assign layer5_outputs[1173] = ~(layer4_outputs[3801]);
    assign layer5_outputs[1174] = layer4_outputs[2384];
    assign layer5_outputs[1175] = ~((layer4_outputs[2039]) | (layer4_outputs[3091]));
    assign layer5_outputs[1176] = ~(layer4_outputs[4796]) | (layer4_outputs[4852]);
    assign layer5_outputs[1177] = layer4_outputs[1103];
    assign layer5_outputs[1178] = layer4_outputs[3110];
    assign layer5_outputs[1179] = (layer4_outputs[2745]) & ~(layer4_outputs[3214]);
    assign layer5_outputs[1180] = (layer4_outputs[2843]) & ~(layer4_outputs[3324]);
    assign layer5_outputs[1181] = ~((layer4_outputs[2127]) ^ (layer4_outputs[2846]));
    assign layer5_outputs[1182] = ~(layer4_outputs[4593]) | (layer4_outputs[4154]);
    assign layer5_outputs[1183] = layer4_outputs[3781];
    assign layer5_outputs[1184] = layer4_outputs[2252];
    assign layer5_outputs[1185] = layer4_outputs[3757];
    assign layer5_outputs[1186] = (layer4_outputs[2117]) ^ (layer4_outputs[46]);
    assign layer5_outputs[1187] = layer4_outputs[4666];
    assign layer5_outputs[1188] = ~(layer4_outputs[301]);
    assign layer5_outputs[1189] = layer4_outputs[2977];
    assign layer5_outputs[1190] = 1'b1;
    assign layer5_outputs[1191] = ~((layer4_outputs[2516]) | (layer4_outputs[632]));
    assign layer5_outputs[1192] = layer4_outputs[3062];
    assign layer5_outputs[1193] = (layer4_outputs[606]) & ~(layer4_outputs[3700]);
    assign layer5_outputs[1194] = 1'b0;
    assign layer5_outputs[1195] = (layer4_outputs[4439]) & (layer4_outputs[956]);
    assign layer5_outputs[1196] = (layer4_outputs[1284]) ^ (layer4_outputs[2734]);
    assign layer5_outputs[1197] = (layer4_outputs[146]) & ~(layer4_outputs[38]);
    assign layer5_outputs[1198] = ~((layer4_outputs[2978]) ^ (layer4_outputs[2127]));
    assign layer5_outputs[1199] = ~((layer4_outputs[4559]) ^ (layer4_outputs[2690]));
    assign layer5_outputs[1200] = (layer4_outputs[545]) & ~(layer4_outputs[2444]);
    assign layer5_outputs[1201] = ~((layer4_outputs[2404]) ^ (layer4_outputs[5009]));
    assign layer5_outputs[1202] = ~(layer4_outputs[3081]);
    assign layer5_outputs[1203] = (layer4_outputs[5101]) & ~(layer4_outputs[304]);
    assign layer5_outputs[1204] = (layer4_outputs[4579]) & ~(layer4_outputs[4071]);
    assign layer5_outputs[1205] = layer4_outputs[3473];
    assign layer5_outputs[1206] = ~((layer4_outputs[1115]) & (layer4_outputs[4890]));
    assign layer5_outputs[1207] = ~((layer4_outputs[1114]) | (layer4_outputs[353]));
    assign layer5_outputs[1208] = (layer4_outputs[2002]) & ~(layer4_outputs[3279]);
    assign layer5_outputs[1209] = (layer4_outputs[2508]) ^ (layer4_outputs[22]);
    assign layer5_outputs[1210] = ~(layer4_outputs[1372]);
    assign layer5_outputs[1211] = layer4_outputs[1304];
    assign layer5_outputs[1212] = ~((layer4_outputs[420]) & (layer4_outputs[3159]));
    assign layer5_outputs[1213] = ~(layer4_outputs[3173]);
    assign layer5_outputs[1214] = layer4_outputs[867];
    assign layer5_outputs[1215] = ~(layer4_outputs[3199]) | (layer4_outputs[1767]);
    assign layer5_outputs[1216] = ~((layer4_outputs[1248]) ^ (layer4_outputs[1100]));
    assign layer5_outputs[1217] = ~(layer4_outputs[4527]) | (layer4_outputs[4608]);
    assign layer5_outputs[1218] = (layer4_outputs[641]) & (layer4_outputs[721]);
    assign layer5_outputs[1219] = layer4_outputs[864];
    assign layer5_outputs[1220] = ~(layer4_outputs[219]);
    assign layer5_outputs[1221] = ~(layer4_outputs[393]);
    assign layer5_outputs[1222] = (layer4_outputs[1058]) & (layer4_outputs[228]);
    assign layer5_outputs[1223] = layer4_outputs[5112];
    assign layer5_outputs[1224] = (layer4_outputs[2083]) & ~(layer4_outputs[2298]);
    assign layer5_outputs[1225] = layer4_outputs[4005];
    assign layer5_outputs[1226] = 1'b0;
    assign layer5_outputs[1227] = ~(layer4_outputs[2488]) | (layer4_outputs[4938]);
    assign layer5_outputs[1228] = (layer4_outputs[4301]) ^ (layer4_outputs[417]);
    assign layer5_outputs[1229] = ~(layer4_outputs[3441]) | (layer4_outputs[1518]);
    assign layer5_outputs[1230] = (layer4_outputs[3884]) & ~(layer4_outputs[3950]);
    assign layer5_outputs[1231] = (layer4_outputs[3115]) & (layer4_outputs[4537]);
    assign layer5_outputs[1232] = ~((layer4_outputs[1319]) & (layer4_outputs[74]));
    assign layer5_outputs[1233] = (layer4_outputs[3769]) & (layer4_outputs[4574]);
    assign layer5_outputs[1234] = ~((layer4_outputs[1822]) & (layer4_outputs[1892]));
    assign layer5_outputs[1235] = (layer4_outputs[1753]) & ~(layer4_outputs[2094]);
    assign layer5_outputs[1236] = ~((layer4_outputs[1913]) | (layer4_outputs[1253]));
    assign layer5_outputs[1237] = ~((layer4_outputs[2930]) & (layer4_outputs[3755]));
    assign layer5_outputs[1238] = ~((layer4_outputs[1427]) | (layer4_outputs[5079]));
    assign layer5_outputs[1239] = ~(layer4_outputs[1437]) | (layer4_outputs[4981]);
    assign layer5_outputs[1240] = layer4_outputs[3428];
    assign layer5_outputs[1241] = (layer4_outputs[1758]) & ~(layer4_outputs[4163]);
    assign layer5_outputs[1242] = (layer4_outputs[294]) & ~(layer4_outputs[1383]);
    assign layer5_outputs[1243] = (layer4_outputs[3634]) & ~(layer4_outputs[2666]);
    assign layer5_outputs[1244] = layer4_outputs[2141];
    assign layer5_outputs[1245] = ~((layer4_outputs[1546]) | (layer4_outputs[822]));
    assign layer5_outputs[1246] = ~(layer4_outputs[3097]);
    assign layer5_outputs[1247] = ~(layer4_outputs[2920]);
    assign layer5_outputs[1248] = layer4_outputs[3304];
    assign layer5_outputs[1249] = ~(layer4_outputs[2626]);
    assign layer5_outputs[1250] = ~(layer4_outputs[2634]);
    assign layer5_outputs[1251] = layer4_outputs[2742];
    assign layer5_outputs[1252] = 1'b0;
    assign layer5_outputs[1253] = layer4_outputs[2070];
    assign layer5_outputs[1254] = 1'b1;
    assign layer5_outputs[1255] = (layer4_outputs[1647]) & ~(layer4_outputs[2593]);
    assign layer5_outputs[1256] = (layer4_outputs[4680]) ^ (layer4_outputs[4721]);
    assign layer5_outputs[1257] = ~((layer4_outputs[1615]) ^ (layer4_outputs[3282]));
    assign layer5_outputs[1258] = ~((layer4_outputs[3931]) | (layer4_outputs[2759]));
    assign layer5_outputs[1259] = (layer4_outputs[779]) & ~(layer4_outputs[4552]);
    assign layer5_outputs[1260] = layer4_outputs[1719];
    assign layer5_outputs[1261] = ~(layer4_outputs[2345]);
    assign layer5_outputs[1262] = layer4_outputs[789];
    assign layer5_outputs[1263] = layer4_outputs[722];
    assign layer5_outputs[1264] = (layer4_outputs[3507]) & ~(layer4_outputs[3252]);
    assign layer5_outputs[1265] = layer4_outputs[3436];
    assign layer5_outputs[1266] = layer4_outputs[907];
    assign layer5_outputs[1267] = 1'b0;
    assign layer5_outputs[1268] = (layer4_outputs[2118]) & ~(layer4_outputs[908]);
    assign layer5_outputs[1269] = ~((layer4_outputs[2111]) | (layer4_outputs[2881]));
    assign layer5_outputs[1270] = (layer4_outputs[1378]) & (layer4_outputs[3387]);
    assign layer5_outputs[1271] = layer4_outputs[1001];
    assign layer5_outputs[1272] = ~(layer4_outputs[2323]);
    assign layer5_outputs[1273] = ~(layer4_outputs[3038]);
    assign layer5_outputs[1274] = ~(layer4_outputs[2673]);
    assign layer5_outputs[1275] = ~(layer4_outputs[3796]);
    assign layer5_outputs[1276] = 1'b1;
    assign layer5_outputs[1277] = ~(layer4_outputs[4946]);
    assign layer5_outputs[1278] = layer4_outputs[1812];
    assign layer5_outputs[1279] = ~(layer4_outputs[3423]) | (layer4_outputs[2871]);
    assign layer5_outputs[1280] = ~(layer4_outputs[783]);
    assign layer5_outputs[1281] = ~(layer4_outputs[3008]);
    assign layer5_outputs[1282] = (layer4_outputs[4816]) | (layer4_outputs[2491]);
    assign layer5_outputs[1283] = ~((layer4_outputs[4113]) & (layer4_outputs[702]));
    assign layer5_outputs[1284] = (layer4_outputs[3085]) & ~(layer4_outputs[4593]);
    assign layer5_outputs[1285] = ~(layer4_outputs[997]) | (layer4_outputs[4576]);
    assign layer5_outputs[1286] = ~(layer4_outputs[989]) | (layer4_outputs[1493]);
    assign layer5_outputs[1287] = (layer4_outputs[2111]) & ~(layer4_outputs[3562]);
    assign layer5_outputs[1288] = (layer4_outputs[1055]) & (layer4_outputs[2841]);
    assign layer5_outputs[1289] = ~(layer4_outputs[68]);
    assign layer5_outputs[1290] = (layer4_outputs[4039]) ^ (layer4_outputs[2533]);
    assign layer5_outputs[1291] = (layer4_outputs[390]) & (layer4_outputs[1485]);
    assign layer5_outputs[1292] = ~(layer4_outputs[1582]);
    assign layer5_outputs[1293] = layer4_outputs[5025];
    assign layer5_outputs[1294] = ~(layer4_outputs[3972]);
    assign layer5_outputs[1295] = ~((layer4_outputs[1330]) | (layer4_outputs[4173]));
    assign layer5_outputs[1296] = layer4_outputs[132];
    assign layer5_outputs[1297] = layer4_outputs[3765];
    assign layer5_outputs[1298] = layer4_outputs[382];
    assign layer5_outputs[1299] = ~(layer4_outputs[4375]);
    assign layer5_outputs[1300] = layer4_outputs[3556];
    assign layer5_outputs[1301] = ~(layer4_outputs[193]);
    assign layer5_outputs[1302] = layer4_outputs[4525];
    assign layer5_outputs[1303] = 1'b0;
    assign layer5_outputs[1304] = ~((layer4_outputs[602]) & (layer4_outputs[2599]));
    assign layer5_outputs[1305] = ~(layer4_outputs[278]);
    assign layer5_outputs[1306] = ~(layer4_outputs[2994]) | (layer4_outputs[513]);
    assign layer5_outputs[1307] = layer4_outputs[4142];
    assign layer5_outputs[1308] = ~(layer4_outputs[3849]);
    assign layer5_outputs[1309] = layer4_outputs[2557];
    assign layer5_outputs[1310] = (layer4_outputs[1814]) & ~(layer4_outputs[2876]);
    assign layer5_outputs[1311] = layer4_outputs[2780];
    assign layer5_outputs[1312] = ~(layer4_outputs[1909]) | (layer4_outputs[4170]);
    assign layer5_outputs[1313] = ~(layer4_outputs[2933]) | (layer4_outputs[3894]);
    assign layer5_outputs[1314] = (layer4_outputs[4118]) & (layer4_outputs[3227]);
    assign layer5_outputs[1315] = ~((layer4_outputs[1417]) | (layer4_outputs[79]));
    assign layer5_outputs[1316] = ~((layer4_outputs[815]) | (layer4_outputs[3218]));
    assign layer5_outputs[1317] = ~((layer4_outputs[3522]) ^ (layer4_outputs[3285]));
    assign layer5_outputs[1318] = 1'b1;
    assign layer5_outputs[1319] = (layer4_outputs[3827]) | (layer4_outputs[4903]);
    assign layer5_outputs[1320] = ~((layer4_outputs[1004]) & (layer4_outputs[2945]));
    assign layer5_outputs[1321] = layer4_outputs[4734];
    assign layer5_outputs[1322] = layer4_outputs[4443];
    assign layer5_outputs[1323] = ~(layer4_outputs[4969]) | (layer4_outputs[55]);
    assign layer5_outputs[1324] = 1'b1;
    assign layer5_outputs[1325] = (layer4_outputs[4097]) & (layer4_outputs[3202]);
    assign layer5_outputs[1326] = layer4_outputs[1009];
    assign layer5_outputs[1327] = (layer4_outputs[2485]) | (layer4_outputs[402]);
    assign layer5_outputs[1328] = ~(layer4_outputs[3251]);
    assign layer5_outputs[1329] = layer4_outputs[375];
    assign layer5_outputs[1330] = ~(layer4_outputs[0]);
    assign layer5_outputs[1331] = layer4_outputs[1605];
    assign layer5_outputs[1332] = ~((layer4_outputs[3009]) & (layer4_outputs[3397]));
    assign layer5_outputs[1333] = ~(layer4_outputs[745]) | (layer4_outputs[3196]);
    assign layer5_outputs[1334] = layer4_outputs[2121];
    assign layer5_outputs[1335] = ~(layer4_outputs[3093]);
    assign layer5_outputs[1336] = (layer4_outputs[2061]) | (layer4_outputs[206]);
    assign layer5_outputs[1337] = layer4_outputs[3079];
    assign layer5_outputs[1338] = ~(layer4_outputs[1539]);
    assign layer5_outputs[1339] = (layer4_outputs[4443]) & ~(layer4_outputs[4278]);
    assign layer5_outputs[1340] = layer4_outputs[1977];
    assign layer5_outputs[1341] = ~(layer4_outputs[4737]);
    assign layer5_outputs[1342] = ~(layer4_outputs[3696]);
    assign layer5_outputs[1343] = (layer4_outputs[279]) | (layer4_outputs[1983]);
    assign layer5_outputs[1344] = layer4_outputs[4491];
    assign layer5_outputs[1345] = ~((layer4_outputs[3711]) & (layer4_outputs[3427]));
    assign layer5_outputs[1346] = (layer4_outputs[507]) & (layer4_outputs[467]);
    assign layer5_outputs[1347] = ~(layer4_outputs[902]);
    assign layer5_outputs[1348] = (layer4_outputs[2131]) ^ (layer4_outputs[601]);
    assign layer5_outputs[1349] = layer4_outputs[4841];
    assign layer5_outputs[1350] = (layer4_outputs[2525]) ^ (layer4_outputs[4746]);
    assign layer5_outputs[1351] = layer4_outputs[63];
    assign layer5_outputs[1352] = (layer4_outputs[2273]) & ~(layer4_outputs[797]);
    assign layer5_outputs[1353] = layer4_outputs[3807];
    assign layer5_outputs[1354] = (layer4_outputs[2369]) & (layer4_outputs[4807]);
    assign layer5_outputs[1355] = (layer4_outputs[3422]) & ~(layer4_outputs[1951]);
    assign layer5_outputs[1356] = ~(layer4_outputs[2699]);
    assign layer5_outputs[1357] = ~((layer4_outputs[4212]) & (layer4_outputs[1140]));
    assign layer5_outputs[1358] = layer4_outputs[237];
    assign layer5_outputs[1359] = (layer4_outputs[1221]) ^ (layer4_outputs[1904]);
    assign layer5_outputs[1360] = ~((layer4_outputs[4007]) | (layer4_outputs[3896]));
    assign layer5_outputs[1361] = ~(layer4_outputs[2531]);
    assign layer5_outputs[1362] = ~(layer4_outputs[416]);
    assign layer5_outputs[1363] = ~(layer4_outputs[2385]);
    assign layer5_outputs[1364] = (layer4_outputs[4541]) | (layer4_outputs[4130]);
    assign layer5_outputs[1365] = layer4_outputs[3361];
    assign layer5_outputs[1366] = layer4_outputs[3892];
    assign layer5_outputs[1367] = ~(layer4_outputs[3284]);
    assign layer5_outputs[1368] = 1'b1;
    assign layer5_outputs[1369] = ~(layer4_outputs[1683]);
    assign layer5_outputs[1370] = (layer4_outputs[5038]) & ~(layer4_outputs[2358]);
    assign layer5_outputs[1371] = layer4_outputs[3750];
    assign layer5_outputs[1372] = ~(layer4_outputs[4789]) | (layer4_outputs[2655]);
    assign layer5_outputs[1373] = ~(layer4_outputs[1916]) | (layer4_outputs[1504]);
    assign layer5_outputs[1374] = ~(layer4_outputs[2074]) | (layer4_outputs[1557]);
    assign layer5_outputs[1375] = (layer4_outputs[4929]) | (layer4_outputs[2288]);
    assign layer5_outputs[1376] = layer4_outputs[1077];
    assign layer5_outputs[1377] = ~(layer4_outputs[4247]);
    assign layer5_outputs[1378] = (layer4_outputs[4319]) | (layer4_outputs[3584]);
    assign layer5_outputs[1379] = layer4_outputs[4123];
    assign layer5_outputs[1380] = layer4_outputs[2513];
    assign layer5_outputs[1381] = ~((layer4_outputs[2761]) & (layer4_outputs[172]));
    assign layer5_outputs[1382] = (layer4_outputs[634]) & ~(layer4_outputs[2]);
    assign layer5_outputs[1383] = ~((layer4_outputs[2538]) & (layer4_outputs[796]));
    assign layer5_outputs[1384] = ~((layer4_outputs[4454]) & (layer4_outputs[4573]));
    assign layer5_outputs[1385] = layer4_outputs[4086];
    assign layer5_outputs[1386] = layer4_outputs[2694];
    assign layer5_outputs[1387] = ~(layer4_outputs[360]);
    assign layer5_outputs[1388] = 1'b1;
    assign layer5_outputs[1389] = ~(layer4_outputs[455]);
    assign layer5_outputs[1390] = (layer4_outputs[742]) & ~(layer4_outputs[4010]);
    assign layer5_outputs[1391] = ~((layer4_outputs[4743]) ^ (layer4_outputs[728]));
    assign layer5_outputs[1392] = (layer4_outputs[2073]) ^ (layer4_outputs[4125]);
    assign layer5_outputs[1393] = ~(layer4_outputs[2089]) | (layer4_outputs[2076]);
    assign layer5_outputs[1394] = layer4_outputs[2422];
    assign layer5_outputs[1395] = ~(layer4_outputs[1861]) | (layer4_outputs[14]);
    assign layer5_outputs[1396] = 1'b1;
    assign layer5_outputs[1397] = ~(layer4_outputs[1326]);
    assign layer5_outputs[1398] = ~((layer4_outputs[4440]) ^ (layer4_outputs[2254]));
    assign layer5_outputs[1399] = ~(layer4_outputs[3462]);
    assign layer5_outputs[1400] = layer4_outputs[4444];
    assign layer5_outputs[1401] = 1'b1;
    assign layer5_outputs[1402] = ~(layer4_outputs[298]);
    assign layer5_outputs[1403] = ~(layer4_outputs[1991]) | (layer4_outputs[4073]);
    assign layer5_outputs[1404] = layer4_outputs[4529];
    assign layer5_outputs[1405] = layer4_outputs[1409];
    assign layer5_outputs[1406] = ~((layer4_outputs[1843]) | (layer4_outputs[1630]));
    assign layer5_outputs[1407] = ~(layer4_outputs[3964]);
    assign layer5_outputs[1408] = (layer4_outputs[2377]) & (layer4_outputs[1811]);
    assign layer5_outputs[1409] = (layer4_outputs[1171]) & ~(layer4_outputs[428]);
    assign layer5_outputs[1410] = 1'b1;
    assign layer5_outputs[1411] = ~(layer4_outputs[3415]) | (layer4_outputs[3491]);
    assign layer5_outputs[1412] = (layer4_outputs[3584]) ^ (layer4_outputs[1242]);
    assign layer5_outputs[1413] = ~((layer4_outputs[3890]) & (layer4_outputs[4140]));
    assign layer5_outputs[1414] = (layer4_outputs[2069]) | (layer4_outputs[1777]);
    assign layer5_outputs[1415] = ~((layer4_outputs[4838]) & (layer4_outputs[3569]));
    assign layer5_outputs[1416] = ~(layer4_outputs[431]);
    assign layer5_outputs[1417] = layer4_outputs[3];
    assign layer5_outputs[1418] = ~(layer4_outputs[3811]);
    assign layer5_outputs[1419] = ~((layer4_outputs[2976]) | (layer4_outputs[3956]));
    assign layer5_outputs[1420] = ~(layer4_outputs[2696]);
    assign layer5_outputs[1421] = layer4_outputs[3616];
    assign layer5_outputs[1422] = ~(layer4_outputs[1525]);
    assign layer5_outputs[1423] = ~(layer4_outputs[1457]) | (layer4_outputs[49]);
    assign layer5_outputs[1424] = layer4_outputs[3240];
    assign layer5_outputs[1425] = layer4_outputs[246];
    assign layer5_outputs[1426] = layer4_outputs[439];
    assign layer5_outputs[1427] = ~(layer4_outputs[2658]);
    assign layer5_outputs[1428] = ~(layer4_outputs[494]);
    assign layer5_outputs[1429] = ~(layer4_outputs[58]) | (layer4_outputs[1390]);
    assign layer5_outputs[1430] = 1'b1;
    assign layer5_outputs[1431] = layer4_outputs[329];
    assign layer5_outputs[1432] = layer4_outputs[2886];
    assign layer5_outputs[1433] = (layer4_outputs[77]) & ~(layer4_outputs[4264]);
    assign layer5_outputs[1434] = layer4_outputs[2168];
    assign layer5_outputs[1435] = (layer4_outputs[4435]) | (layer4_outputs[805]);
    assign layer5_outputs[1436] = (layer4_outputs[2455]) & ~(layer4_outputs[2223]);
    assign layer5_outputs[1437] = layer4_outputs[112];
    assign layer5_outputs[1438] = ~(layer4_outputs[2809]) | (layer4_outputs[2715]);
    assign layer5_outputs[1439] = (layer4_outputs[1352]) ^ (layer4_outputs[1828]);
    assign layer5_outputs[1440] = ~((layer4_outputs[4267]) ^ (layer4_outputs[1078]));
    assign layer5_outputs[1441] = ~(layer4_outputs[5010]);
    assign layer5_outputs[1442] = layer4_outputs[414];
    assign layer5_outputs[1443] = layer4_outputs[1374];
    assign layer5_outputs[1444] = ~(layer4_outputs[788]);
    assign layer5_outputs[1445] = layer4_outputs[999];
    assign layer5_outputs[1446] = layer4_outputs[3510];
    assign layer5_outputs[1447] = (layer4_outputs[2749]) & (layer4_outputs[1670]);
    assign layer5_outputs[1448] = layer4_outputs[4723];
    assign layer5_outputs[1449] = ~((layer4_outputs[2494]) & (layer4_outputs[3679]));
    assign layer5_outputs[1450] = layer4_outputs[4374];
    assign layer5_outputs[1451] = layer4_outputs[3200];
    assign layer5_outputs[1452] = (layer4_outputs[2266]) ^ (layer4_outputs[427]);
    assign layer5_outputs[1453] = ~((layer4_outputs[3613]) & (layer4_outputs[358]));
    assign layer5_outputs[1454] = (layer4_outputs[3378]) ^ (layer4_outputs[1042]);
    assign layer5_outputs[1455] = (layer4_outputs[2600]) & ~(layer4_outputs[1744]);
    assign layer5_outputs[1456] = ~(layer4_outputs[2815]);
    assign layer5_outputs[1457] = ~(layer4_outputs[2030]) | (layer4_outputs[3407]);
    assign layer5_outputs[1458] = ~((layer4_outputs[1092]) ^ (layer4_outputs[4157]));
    assign layer5_outputs[1459] = layer4_outputs[3981];
    assign layer5_outputs[1460] = layer4_outputs[1997];
    assign layer5_outputs[1461] = layer4_outputs[3877];
    assign layer5_outputs[1462] = (layer4_outputs[496]) & ~(layer4_outputs[186]);
    assign layer5_outputs[1463] = layer4_outputs[2181];
    assign layer5_outputs[1464] = ~(layer4_outputs[2866]);
    assign layer5_outputs[1465] = ~(layer4_outputs[4066]);
    assign layer5_outputs[1466] = ~(layer4_outputs[3261]);
    assign layer5_outputs[1467] = ~(layer4_outputs[3398]);
    assign layer5_outputs[1468] = ~((layer4_outputs[4346]) | (layer4_outputs[3611]));
    assign layer5_outputs[1469] = 1'b0;
    assign layer5_outputs[1470] = (layer4_outputs[3448]) & (layer4_outputs[3707]);
    assign layer5_outputs[1471] = ~(layer4_outputs[4766]) | (layer4_outputs[2217]);
    assign layer5_outputs[1472] = layer4_outputs[5109];
    assign layer5_outputs[1473] = (layer4_outputs[4997]) ^ (layer4_outputs[1252]);
    assign layer5_outputs[1474] = layer4_outputs[1017];
    assign layer5_outputs[1475] = ~(layer4_outputs[1266]);
    assign layer5_outputs[1476] = ~(layer4_outputs[4200]);
    assign layer5_outputs[1477] = ~(layer4_outputs[1589]);
    assign layer5_outputs[1478] = ~(layer4_outputs[1312]);
    assign layer5_outputs[1479] = (layer4_outputs[1005]) & ~(layer4_outputs[179]);
    assign layer5_outputs[1480] = 1'b0;
    assign layer5_outputs[1481] = ~(layer4_outputs[2380]) | (layer4_outputs[112]);
    assign layer5_outputs[1482] = layer4_outputs[400];
    assign layer5_outputs[1483] = (layer4_outputs[3912]) & (layer4_outputs[2057]);
    assign layer5_outputs[1484] = layer4_outputs[5005];
    assign layer5_outputs[1485] = ~(layer4_outputs[4564]);
    assign layer5_outputs[1486] = layer4_outputs[1618];
    assign layer5_outputs[1487] = (layer4_outputs[600]) & ~(layer4_outputs[1651]);
    assign layer5_outputs[1488] = ~(layer4_outputs[1259]) | (layer4_outputs[4860]);
    assign layer5_outputs[1489] = (layer4_outputs[4551]) & ~(layer4_outputs[4662]);
    assign layer5_outputs[1490] = layer4_outputs[4459];
    assign layer5_outputs[1491] = ~(layer4_outputs[4955]);
    assign layer5_outputs[1492] = layer4_outputs[256];
    assign layer5_outputs[1493] = (layer4_outputs[3316]) & ~(layer4_outputs[5071]);
    assign layer5_outputs[1494] = ~(layer4_outputs[1262]) | (layer4_outputs[2322]);
    assign layer5_outputs[1495] = layer4_outputs[2827];
    assign layer5_outputs[1496] = layer4_outputs[3693];
    assign layer5_outputs[1497] = ~((layer4_outputs[2592]) ^ (layer4_outputs[3891]));
    assign layer5_outputs[1498] = (layer4_outputs[4074]) & ~(layer4_outputs[1846]);
    assign layer5_outputs[1499] = ~(layer4_outputs[171]);
    assign layer5_outputs[1500] = (layer4_outputs[4572]) & ~(layer4_outputs[284]);
    assign layer5_outputs[1501] = ~((layer4_outputs[4747]) & (layer4_outputs[1437]));
    assign layer5_outputs[1502] = layer4_outputs[327];
    assign layer5_outputs[1503] = (layer4_outputs[3182]) & ~(layer4_outputs[1179]);
    assign layer5_outputs[1504] = ~((layer4_outputs[1033]) & (layer4_outputs[3908]));
    assign layer5_outputs[1505] = (layer4_outputs[1484]) & ~(layer4_outputs[4382]);
    assign layer5_outputs[1506] = (layer4_outputs[2060]) & (layer4_outputs[3194]);
    assign layer5_outputs[1507] = (layer4_outputs[2311]) | (layer4_outputs[3157]);
    assign layer5_outputs[1508] = 1'b0;
    assign layer5_outputs[1509] = (layer4_outputs[4986]) ^ (layer4_outputs[3467]);
    assign layer5_outputs[1510] = layer4_outputs[189];
    assign layer5_outputs[1511] = ~(layer4_outputs[1188]);
    assign layer5_outputs[1512] = ~((layer4_outputs[2823]) ^ (layer4_outputs[3618]));
    assign layer5_outputs[1513] = ~(layer4_outputs[3526]);
    assign layer5_outputs[1514] = layer4_outputs[897];
    assign layer5_outputs[1515] = ~((layer4_outputs[1065]) | (layer4_outputs[139]));
    assign layer5_outputs[1516] = (layer4_outputs[1701]) & ~(layer4_outputs[4249]);
    assign layer5_outputs[1517] = ~(layer4_outputs[1456]);
    assign layer5_outputs[1518] = (layer4_outputs[661]) | (layer4_outputs[2085]);
    assign layer5_outputs[1519] = ~((layer4_outputs[1428]) ^ (layer4_outputs[2446]));
    assign layer5_outputs[1520] = ~(layer4_outputs[3590]);
    assign layer5_outputs[1521] = ~((layer4_outputs[3716]) & (layer4_outputs[4926]));
    assign layer5_outputs[1522] = (layer4_outputs[3955]) & (layer4_outputs[1309]);
    assign layer5_outputs[1523] = layer4_outputs[1023];
    assign layer5_outputs[1524] = (layer4_outputs[1737]) & ~(layer4_outputs[4213]);
    assign layer5_outputs[1525] = ~((layer4_outputs[3674]) | (layer4_outputs[4544]));
    assign layer5_outputs[1526] = ~(layer4_outputs[42]) | (layer4_outputs[4006]);
    assign layer5_outputs[1527] = ~(layer4_outputs[433]);
    assign layer5_outputs[1528] = 1'b1;
    assign layer5_outputs[1529] = ~((layer4_outputs[3347]) | (layer4_outputs[2638]));
    assign layer5_outputs[1530] = layer4_outputs[2196];
    assign layer5_outputs[1531] = (layer4_outputs[2610]) & ~(layer4_outputs[549]);
    assign layer5_outputs[1532] = layer4_outputs[249];
    assign layer5_outputs[1533] = 1'b1;
    assign layer5_outputs[1534] = ~(layer4_outputs[2954]);
    assign layer5_outputs[1535] = layer4_outputs[150];
    assign layer5_outputs[1536] = (layer4_outputs[1700]) | (layer4_outputs[2610]);
    assign layer5_outputs[1537] = layer4_outputs[2186];
    assign layer5_outputs[1538] = 1'b0;
    assign layer5_outputs[1539] = ~((layer4_outputs[4000]) ^ (layer4_outputs[4613]));
    assign layer5_outputs[1540] = 1'b0;
    assign layer5_outputs[1541] = ~(layer4_outputs[2379]);
    assign layer5_outputs[1542] = (layer4_outputs[4004]) ^ (layer4_outputs[506]);
    assign layer5_outputs[1543] = ~((layer4_outputs[2204]) ^ (layer4_outputs[397]));
    assign layer5_outputs[1544] = ~(layer4_outputs[3542]);
    assign layer5_outputs[1545] = ~(layer4_outputs[3830]);
    assign layer5_outputs[1546] = (layer4_outputs[2612]) | (layer4_outputs[2710]);
    assign layer5_outputs[1547] = ~(layer4_outputs[3099]);
    assign layer5_outputs[1548] = ~(layer4_outputs[4851]) | (layer4_outputs[987]);
    assign layer5_outputs[1549] = (layer4_outputs[3127]) & (layer4_outputs[523]);
    assign layer5_outputs[1550] = layer4_outputs[1234];
    assign layer5_outputs[1551] = (layer4_outputs[2428]) & ~(layer4_outputs[617]);
    assign layer5_outputs[1552] = layer4_outputs[4892];
    assign layer5_outputs[1553] = ~((layer4_outputs[3920]) ^ (layer4_outputs[3885]));
    assign layer5_outputs[1554] = ~(layer4_outputs[1889]);
    assign layer5_outputs[1555] = ~(layer4_outputs[1617]);
    assign layer5_outputs[1556] = (layer4_outputs[3833]) ^ (layer4_outputs[4618]);
    assign layer5_outputs[1557] = ~(layer4_outputs[3200]) | (layer4_outputs[2880]);
    assign layer5_outputs[1558] = ~(layer4_outputs[103]);
    assign layer5_outputs[1559] = (layer4_outputs[432]) | (layer4_outputs[3133]);
    assign layer5_outputs[1560] = (layer4_outputs[2075]) & (layer4_outputs[1847]);
    assign layer5_outputs[1561] = layer4_outputs[2969];
    assign layer5_outputs[1562] = ~(layer4_outputs[3225]);
    assign layer5_outputs[1563] = ~(layer4_outputs[59]);
    assign layer5_outputs[1564] = (layer4_outputs[2777]) | (layer4_outputs[617]);
    assign layer5_outputs[1565] = 1'b0;
    assign layer5_outputs[1566] = ~((layer4_outputs[1122]) | (layer4_outputs[1315]));
    assign layer5_outputs[1567] = ~(layer4_outputs[1543]) | (layer4_outputs[911]);
    assign layer5_outputs[1568] = layer4_outputs[4307];
    assign layer5_outputs[1569] = layer4_outputs[2096];
    assign layer5_outputs[1570] = layer4_outputs[1958];
    assign layer5_outputs[1571] = ~(layer4_outputs[4064]) | (layer4_outputs[2066]);
    assign layer5_outputs[1572] = ~(layer4_outputs[2805]);
    assign layer5_outputs[1573] = ~(layer4_outputs[4099]);
    assign layer5_outputs[1574] = layer4_outputs[3517];
    assign layer5_outputs[1575] = (layer4_outputs[3002]) | (layer4_outputs[560]);
    assign layer5_outputs[1576] = layer4_outputs[850];
    assign layer5_outputs[1577] = layer4_outputs[922];
    assign layer5_outputs[1578] = ~(layer4_outputs[4311]);
    assign layer5_outputs[1579] = ~(layer4_outputs[3969]);
    assign layer5_outputs[1580] = ~((layer4_outputs[4211]) ^ (layer4_outputs[3663]));
    assign layer5_outputs[1581] = 1'b1;
    assign layer5_outputs[1582] = ~(layer4_outputs[939]) | (layer4_outputs[3039]);
    assign layer5_outputs[1583] = ~(layer4_outputs[2013]);
    assign layer5_outputs[1584] = (layer4_outputs[1882]) & ~(layer4_outputs[2850]);
    assign layer5_outputs[1585] = layer4_outputs[4071];
    assign layer5_outputs[1586] = ~((layer4_outputs[3161]) & (layer4_outputs[3765]));
    assign layer5_outputs[1587] = (layer4_outputs[4329]) & ~(layer4_outputs[3018]);
    assign layer5_outputs[1588] = ~(layer4_outputs[1549]);
    assign layer5_outputs[1589] = ~(layer4_outputs[2397]);
    assign layer5_outputs[1590] = ~(layer4_outputs[3966]);
    assign layer5_outputs[1591] = (layer4_outputs[1716]) ^ (layer4_outputs[376]);
    assign layer5_outputs[1592] = ~(layer4_outputs[2890]) | (layer4_outputs[2559]);
    assign layer5_outputs[1593] = layer4_outputs[1991];
    assign layer5_outputs[1594] = ~(layer4_outputs[1204]);
    assign layer5_outputs[1595] = ~((layer4_outputs[2669]) & (layer4_outputs[2430]));
    assign layer5_outputs[1596] = (layer4_outputs[263]) | (layer4_outputs[2267]);
    assign layer5_outputs[1597] = layer4_outputs[2132];
    assign layer5_outputs[1598] = ~(layer4_outputs[2411]) | (layer4_outputs[4827]);
    assign layer5_outputs[1599] = 1'b1;
    assign layer5_outputs[1600] = layer4_outputs[3101];
    assign layer5_outputs[1601] = layer4_outputs[3277];
    assign layer5_outputs[1602] = ~((layer4_outputs[798]) ^ (layer4_outputs[2159]));
    assign layer5_outputs[1603] = ~((layer4_outputs[478]) & (layer4_outputs[3978]));
    assign layer5_outputs[1604] = ~(layer4_outputs[3813]);
    assign layer5_outputs[1605] = ~(layer4_outputs[2031]);
    assign layer5_outputs[1606] = ~(layer4_outputs[2407]);
    assign layer5_outputs[1607] = (layer4_outputs[1482]) & ~(layer4_outputs[4976]);
    assign layer5_outputs[1608] = layer4_outputs[736];
    assign layer5_outputs[1609] = (layer4_outputs[757]) ^ (layer4_outputs[1277]);
    assign layer5_outputs[1610] = ~(layer4_outputs[3177]);
    assign layer5_outputs[1611] = (layer4_outputs[1106]) & ~(layer4_outputs[3480]);
    assign layer5_outputs[1612] = ~(layer4_outputs[4842]);
    assign layer5_outputs[1613] = ~(layer4_outputs[3881]);
    assign layer5_outputs[1614] = layer4_outputs[3945];
    assign layer5_outputs[1615] = (layer4_outputs[898]) | (layer4_outputs[3011]);
    assign layer5_outputs[1616] = ~((layer4_outputs[4389]) & (layer4_outputs[379]));
    assign layer5_outputs[1617] = ~((layer4_outputs[4174]) | (layer4_outputs[584]));
    assign layer5_outputs[1618] = (layer4_outputs[1366]) ^ (layer4_outputs[3145]);
    assign layer5_outputs[1619] = ~(layer4_outputs[105]);
    assign layer5_outputs[1620] = ~(layer4_outputs[2565]) | (layer4_outputs[1218]);
    assign layer5_outputs[1621] = ~(layer4_outputs[3901]);
    assign layer5_outputs[1622] = (layer4_outputs[3773]) & ~(layer4_outputs[1996]);
    assign layer5_outputs[1623] = (layer4_outputs[4947]) & (layer4_outputs[2652]);
    assign layer5_outputs[1624] = layer4_outputs[1139];
    assign layer5_outputs[1625] = (layer4_outputs[2680]) & ~(layer4_outputs[323]);
    assign layer5_outputs[1626] = layer4_outputs[4275];
    assign layer5_outputs[1627] = ~((layer4_outputs[3158]) | (layer4_outputs[375]));
    assign layer5_outputs[1628] = ~(layer4_outputs[1850]);
    assign layer5_outputs[1629] = ~(layer4_outputs[2579]);
    assign layer5_outputs[1630] = (layer4_outputs[408]) & ~(layer4_outputs[448]);
    assign layer5_outputs[1631] = layer4_outputs[4468];
    assign layer5_outputs[1632] = layer4_outputs[1503];
    assign layer5_outputs[1633] = (layer4_outputs[1984]) & (layer4_outputs[513]);
    assign layer5_outputs[1634] = ~(layer4_outputs[3106]) | (layer4_outputs[1940]);
    assign layer5_outputs[1635] = 1'b1;
    assign layer5_outputs[1636] = ~(layer4_outputs[4283]);
    assign layer5_outputs[1637] = (layer4_outputs[156]) | (layer4_outputs[2408]);
    assign layer5_outputs[1638] = ~(layer4_outputs[2623]);
    assign layer5_outputs[1639] = ~(layer4_outputs[612]);
    assign layer5_outputs[1640] = ~(layer4_outputs[4611]);
    assign layer5_outputs[1641] = (layer4_outputs[3726]) & ~(layer4_outputs[1689]);
    assign layer5_outputs[1642] = ~(layer4_outputs[2780]);
    assign layer5_outputs[1643] = ~((layer4_outputs[1634]) | (layer4_outputs[1589]));
    assign layer5_outputs[1644] = (layer4_outputs[2158]) & ~(layer4_outputs[1873]);
    assign layer5_outputs[1645] = (layer4_outputs[4094]) ^ (layer4_outputs[4399]);
    assign layer5_outputs[1646] = 1'b0;
    assign layer5_outputs[1647] = (layer4_outputs[2782]) | (layer4_outputs[4228]);
    assign layer5_outputs[1648] = ~(layer4_outputs[61]);
    assign layer5_outputs[1649] = layer4_outputs[4078];
    assign layer5_outputs[1650] = ~(layer4_outputs[2511]);
    assign layer5_outputs[1651] = (layer4_outputs[4945]) & ~(layer4_outputs[3305]);
    assign layer5_outputs[1652] = 1'b1;
    assign layer5_outputs[1653] = ~((layer4_outputs[1835]) | (layer4_outputs[4049]));
    assign layer5_outputs[1654] = layer4_outputs[3880];
    assign layer5_outputs[1655] = (layer4_outputs[2353]) & ~(layer4_outputs[1432]);
    assign layer5_outputs[1656] = ~(layer4_outputs[4919]);
    assign layer5_outputs[1657] = layer4_outputs[962];
    assign layer5_outputs[1658] = ~(layer4_outputs[2553]) | (layer4_outputs[1885]);
    assign layer5_outputs[1659] = 1'b1;
    assign layer5_outputs[1660] = (layer4_outputs[3650]) | (layer4_outputs[165]);
    assign layer5_outputs[1661] = ~(layer4_outputs[1952]);
    assign layer5_outputs[1662] = (layer4_outputs[1501]) & (layer4_outputs[4849]);
    assign layer5_outputs[1663] = (layer4_outputs[3037]) & (layer4_outputs[2810]);
    assign layer5_outputs[1664] = (layer4_outputs[3149]) & ~(layer4_outputs[1692]);
    assign layer5_outputs[1665] = (layer4_outputs[2593]) & ~(layer4_outputs[1285]);
    assign layer5_outputs[1666] = layer4_outputs[4687];
    assign layer5_outputs[1667] = 1'b1;
    assign layer5_outputs[1668] = ~((layer4_outputs[2763]) | (layer4_outputs[3750]));
    assign layer5_outputs[1669] = (layer4_outputs[3788]) & (layer4_outputs[3903]);
    assign layer5_outputs[1670] = ~(layer4_outputs[4711]) | (layer4_outputs[2884]);
    assign layer5_outputs[1671] = (layer4_outputs[3260]) & (layer4_outputs[2486]);
    assign layer5_outputs[1672] = (layer4_outputs[2806]) | (layer4_outputs[2114]);
    assign layer5_outputs[1673] = (layer4_outputs[2874]) & (layer4_outputs[4889]);
    assign layer5_outputs[1674] = (layer4_outputs[737]) & ~(layer4_outputs[3133]);
    assign layer5_outputs[1675] = 1'b1;
    assign layer5_outputs[1676] = layer4_outputs[3589];
    assign layer5_outputs[1677] = layer4_outputs[4031];
    assign layer5_outputs[1678] = (layer4_outputs[618]) | (layer4_outputs[3991]);
    assign layer5_outputs[1679] = ~(layer4_outputs[2333]) | (layer4_outputs[4971]);
    assign layer5_outputs[1680] = ~((layer4_outputs[3148]) ^ (layer4_outputs[1201]));
    assign layer5_outputs[1681] = (layer4_outputs[2571]) ^ (layer4_outputs[601]);
    assign layer5_outputs[1682] = ~(layer4_outputs[2700]);
    assign layer5_outputs[1683] = (layer4_outputs[2856]) & ~(layer4_outputs[1916]);
    assign layer5_outputs[1684] = ~(layer4_outputs[3539]);
    assign layer5_outputs[1685] = layer4_outputs[2026];
    assign layer5_outputs[1686] = ~(layer4_outputs[2921]);
    assign layer5_outputs[1687] = ~((layer4_outputs[3979]) & (layer4_outputs[2837]));
    assign layer5_outputs[1688] = (layer4_outputs[313]) & ~(layer4_outputs[4532]);
    assign layer5_outputs[1689] = ~((layer4_outputs[1057]) ^ (layer4_outputs[4719]));
    assign layer5_outputs[1690] = (layer4_outputs[2383]) & (layer4_outputs[145]);
    assign layer5_outputs[1691] = ~(layer4_outputs[766]);
    assign layer5_outputs[1692] = ~((layer4_outputs[1580]) ^ (layer4_outputs[2838]));
    assign layer5_outputs[1693] = (layer4_outputs[754]) ^ (layer4_outputs[1798]);
    assign layer5_outputs[1694] = (layer4_outputs[776]) | (layer4_outputs[526]);
    assign layer5_outputs[1695] = (layer4_outputs[1273]) ^ (layer4_outputs[4477]);
    assign layer5_outputs[1696] = ~((layer4_outputs[3568]) ^ (layer4_outputs[1101]));
    assign layer5_outputs[1697] = (layer4_outputs[3064]) & ~(layer4_outputs[1388]);
    assign layer5_outputs[1698] = ~(layer4_outputs[4655]);
    assign layer5_outputs[1699] = ~(layer4_outputs[3615]);
    assign layer5_outputs[1700] = ~(layer4_outputs[868]);
    assign layer5_outputs[1701] = (layer4_outputs[2456]) ^ (layer4_outputs[954]);
    assign layer5_outputs[1702] = ~(layer4_outputs[984]);
    assign layer5_outputs[1703] = (layer4_outputs[4518]) & (layer4_outputs[2887]);
    assign layer5_outputs[1704] = (layer4_outputs[3280]) | (layer4_outputs[4998]);
    assign layer5_outputs[1705] = ~(layer4_outputs[4092]) | (layer4_outputs[3954]);
    assign layer5_outputs[1706] = ~((layer4_outputs[3100]) ^ (layer4_outputs[3079]));
    assign layer5_outputs[1707] = (layer4_outputs[1251]) & ~(layer4_outputs[1034]);
    assign layer5_outputs[1708] = layer4_outputs[4323];
    assign layer5_outputs[1709] = ~((layer4_outputs[4925]) ^ (layer4_outputs[760]));
    assign layer5_outputs[1710] = (layer4_outputs[2413]) ^ (layer4_outputs[541]);
    assign layer5_outputs[1711] = layer4_outputs[391];
    assign layer5_outputs[1712] = (layer4_outputs[130]) & (layer4_outputs[909]);
    assign layer5_outputs[1713] = ~(layer4_outputs[2130]);
    assign layer5_outputs[1714] = ~((layer4_outputs[1987]) & (layer4_outputs[4017]));
    assign layer5_outputs[1715] = layer4_outputs[2775];
    assign layer5_outputs[1716] = ~((layer4_outputs[4417]) & (layer4_outputs[767]));
    assign layer5_outputs[1717] = (layer4_outputs[4517]) & ~(layer4_outputs[4982]);
    assign layer5_outputs[1718] = ~(layer4_outputs[1901]);
    assign layer5_outputs[1719] = ~((layer4_outputs[2119]) ^ (layer4_outputs[2614]));
    assign layer5_outputs[1720] = ~((layer4_outputs[2308]) | (layer4_outputs[308]));
    assign layer5_outputs[1721] = ~(layer4_outputs[333]) | (layer4_outputs[1365]);
    assign layer5_outputs[1722] = layer4_outputs[75];
    assign layer5_outputs[1723] = ~((layer4_outputs[2109]) & (layer4_outputs[4303]));
    assign layer5_outputs[1724] = (layer4_outputs[4117]) & ~(layer4_outputs[2612]);
    assign layer5_outputs[1725] = ~(layer4_outputs[3272]);
    assign layer5_outputs[1726] = ~((layer4_outputs[554]) | (layer4_outputs[2542]));
    assign layer5_outputs[1727] = layer4_outputs[3593];
    assign layer5_outputs[1728] = ~(layer4_outputs[182]) | (layer4_outputs[1425]);
    assign layer5_outputs[1729] = ~((layer4_outputs[4531]) ^ (layer4_outputs[2909]));
    assign layer5_outputs[1730] = layer4_outputs[3604];
    assign layer5_outputs[1731] = ~(layer4_outputs[4939]);
    assign layer5_outputs[1732] = layer4_outputs[3278];
    assign layer5_outputs[1733] = ~(layer4_outputs[4930]);
    assign layer5_outputs[1734] = ~(layer4_outputs[1918]) | (layer4_outputs[3478]);
    assign layer5_outputs[1735] = (layer4_outputs[4617]) & ~(layer4_outputs[2611]);
    assign layer5_outputs[1736] = ~(layer4_outputs[4019]) | (layer4_outputs[3508]);
    assign layer5_outputs[1737] = ~(layer4_outputs[3029]);
    assign layer5_outputs[1738] = ~((layer4_outputs[4909]) ^ (layer4_outputs[3135]));
    assign layer5_outputs[1739] = ~(layer4_outputs[775]);
    assign layer5_outputs[1740] = (layer4_outputs[5086]) & ~(layer4_outputs[2283]);
    assign layer5_outputs[1741] = (layer4_outputs[3940]) & ~(layer4_outputs[4260]);
    assign layer5_outputs[1742] = 1'b0;
    assign layer5_outputs[1743] = ~(layer4_outputs[3741]) | (layer4_outputs[4112]);
    assign layer5_outputs[1744] = layer4_outputs[528];
    assign layer5_outputs[1745] = layer4_outputs[1696];
    assign layer5_outputs[1746] = ~(layer4_outputs[4082]);
    assign layer5_outputs[1747] = ~(layer4_outputs[2201]);
    assign layer5_outputs[1748] = 1'b1;
    assign layer5_outputs[1749] = ~(layer4_outputs[1852]);
    assign layer5_outputs[1750] = ~(layer4_outputs[2070]);
    assign layer5_outputs[1751] = (layer4_outputs[4964]) ^ (layer4_outputs[3714]);
    assign layer5_outputs[1752] = ~(layer4_outputs[1953]) | (layer4_outputs[247]);
    assign layer5_outputs[1753] = ~(layer4_outputs[4638]);
    assign layer5_outputs[1754] = ~((layer4_outputs[756]) ^ (layer4_outputs[3783]));
    assign layer5_outputs[1755] = ~(layer4_outputs[1655]);
    assign layer5_outputs[1756] = (layer4_outputs[4773]) & ~(layer4_outputs[287]);
    assign layer5_outputs[1757] = (layer4_outputs[4865]) & ~(layer4_outputs[1324]);
    assign layer5_outputs[1758] = layer4_outputs[4648];
    assign layer5_outputs[1759] = ~((layer4_outputs[3795]) & (layer4_outputs[826]));
    assign layer5_outputs[1760] = ~(layer4_outputs[3829]);
    assign layer5_outputs[1761] = layer4_outputs[4152];
    assign layer5_outputs[1762] = layer4_outputs[1178];
    assign layer5_outputs[1763] = layer4_outputs[2137];
    assign layer5_outputs[1764] = 1'b0;
    assign layer5_outputs[1765] = (layer4_outputs[288]) | (layer4_outputs[1128]);
    assign layer5_outputs[1766] = ~(layer4_outputs[3385]);
    assign layer5_outputs[1767] = ~(layer4_outputs[2020]) | (layer4_outputs[1974]);
    assign layer5_outputs[1768] = 1'b0;
    assign layer5_outputs[1769] = layer4_outputs[4131];
    assign layer5_outputs[1770] = (layer4_outputs[3266]) & ~(layer4_outputs[1439]);
    assign layer5_outputs[1771] = ~((layer4_outputs[124]) ^ (layer4_outputs[3220]));
    assign layer5_outputs[1772] = (layer4_outputs[4744]) & ~(layer4_outputs[1322]);
    assign layer5_outputs[1773] = ~(layer4_outputs[3362]);
    assign layer5_outputs[1774] = ~((layer4_outputs[1146]) | (layer4_outputs[4530]));
    assign layer5_outputs[1775] = ~(layer4_outputs[3763]) | (layer4_outputs[1036]);
    assign layer5_outputs[1776] = (layer4_outputs[1854]) | (layer4_outputs[2003]);
    assign layer5_outputs[1777] = (layer4_outputs[1421]) & (layer4_outputs[1632]);
    assign layer5_outputs[1778] = layer4_outputs[2984];
    assign layer5_outputs[1779] = (layer4_outputs[3417]) & (layer4_outputs[34]);
    assign layer5_outputs[1780] = layer4_outputs[4054];
    assign layer5_outputs[1781] = (layer4_outputs[3269]) & ~(layer4_outputs[811]);
    assign layer5_outputs[1782] = layer4_outputs[3405];
    assign layer5_outputs[1783] = ~(layer4_outputs[1256]);
    assign layer5_outputs[1784] = ~(layer4_outputs[2779]) | (layer4_outputs[3521]);
    assign layer5_outputs[1785] = ~(layer4_outputs[4641]);
    assign layer5_outputs[1786] = ~(layer4_outputs[2061]) | (layer4_outputs[2591]);
    assign layer5_outputs[1787] = layer4_outputs[2596];
    assign layer5_outputs[1788] = ~((layer4_outputs[407]) | (layer4_outputs[4269]));
    assign layer5_outputs[1789] = ~((layer4_outputs[3388]) ^ (layer4_outputs[3044]));
    assign layer5_outputs[1790] = layer4_outputs[10];
    assign layer5_outputs[1791] = ~(layer4_outputs[2889]);
    assign layer5_outputs[1792] = ~(layer4_outputs[4008]);
    assign layer5_outputs[1793] = ~((layer4_outputs[2827]) | (layer4_outputs[2944]));
    assign layer5_outputs[1794] = layer4_outputs[3993];
    assign layer5_outputs[1795] = ~((layer4_outputs[1640]) & (layer4_outputs[2268]));
    assign layer5_outputs[1796] = ~(layer4_outputs[4405]);
    assign layer5_outputs[1797] = layer4_outputs[2929];
    assign layer5_outputs[1798] = ~(layer4_outputs[4966]);
    assign layer5_outputs[1799] = layer4_outputs[3904];
    assign layer5_outputs[1800] = (layer4_outputs[2499]) | (layer4_outputs[2432]);
    assign layer5_outputs[1801] = ~(layer4_outputs[4190]);
    assign layer5_outputs[1802] = ~((layer4_outputs[37]) | (layer4_outputs[2412]));
    assign layer5_outputs[1803] = ~((layer4_outputs[4740]) & (layer4_outputs[196]));
    assign layer5_outputs[1804] = ~(layer4_outputs[2243]);
    assign layer5_outputs[1805] = ~(layer4_outputs[1658]) | (layer4_outputs[2865]);
    assign layer5_outputs[1806] = layer4_outputs[3679];
    assign layer5_outputs[1807] = layer4_outputs[692];
    assign layer5_outputs[1808] = (layer4_outputs[4995]) & ~(layer4_outputs[3045]);
    assign layer5_outputs[1809] = ~(layer4_outputs[1772]);
    assign layer5_outputs[1810] = ~((layer4_outputs[1613]) & (layer4_outputs[1114]));
    assign layer5_outputs[1811] = (layer4_outputs[3925]) & ~(layer4_outputs[685]);
    assign layer5_outputs[1812] = 1'b0;
    assign layer5_outputs[1813] = layer4_outputs[2638];
    assign layer5_outputs[1814] = (layer4_outputs[1022]) & ~(layer4_outputs[1837]);
    assign layer5_outputs[1815] = layer4_outputs[4585];
    assign layer5_outputs[1816] = layer4_outputs[4519];
    assign layer5_outputs[1817] = ~(layer4_outputs[3708]);
    assign layer5_outputs[1818] = layer4_outputs[3252];
    assign layer5_outputs[1819] = ~(layer4_outputs[4184]);
    assign layer5_outputs[1820] = (layer4_outputs[3697]) ^ (layer4_outputs[1296]);
    assign layer5_outputs[1821] = layer4_outputs[3916];
    assign layer5_outputs[1822] = layer4_outputs[1193];
    assign layer5_outputs[1823] = ~((layer4_outputs[2296]) ^ (layer4_outputs[4194]));
    assign layer5_outputs[1824] = layer4_outputs[2793];
    assign layer5_outputs[1825] = layer4_outputs[3512];
    assign layer5_outputs[1826] = ~(layer4_outputs[432]);
    assign layer5_outputs[1827] = ~((layer4_outputs[2778]) ^ (layer4_outputs[1908]));
    assign layer5_outputs[1828] = layer4_outputs[1246];
    assign layer5_outputs[1829] = ~(layer4_outputs[281]);
    assign layer5_outputs[1830] = layer4_outputs[1806];
    assign layer5_outputs[1831] = layer4_outputs[1350];
    assign layer5_outputs[1832] = (layer4_outputs[633]) & ~(layer4_outputs[664]);
    assign layer5_outputs[1833] = ~(layer4_outputs[1206]);
    assign layer5_outputs[1834] = ~((layer4_outputs[3438]) & (layer4_outputs[3588]));
    assign layer5_outputs[1835] = (layer4_outputs[187]) & ~(layer4_outputs[1492]);
    assign layer5_outputs[1836] = ~(layer4_outputs[4536]);
    assign layer5_outputs[1837] = ~(layer4_outputs[4748]);
    assign layer5_outputs[1838] = ~(layer4_outputs[340]) | (layer4_outputs[2213]);
    assign layer5_outputs[1839] = ~(layer4_outputs[4576]) | (layer4_outputs[939]);
    assign layer5_outputs[1840] = ~(layer4_outputs[1626]);
    assign layer5_outputs[1841] = (layer4_outputs[1327]) & ~(layer4_outputs[325]);
    assign layer5_outputs[1842] = ~((layer4_outputs[2275]) | (layer4_outputs[1578]));
    assign layer5_outputs[1843] = (layer4_outputs[3334]) & ~(layer4_outputs[125]);
    assign layer5_outputs[1844] = layer4_outputs[4341];
    assign layer5_outputs[1845] = ~(layer4_outputs[3676]);
    assign layer5_outputs[1846] = (layer4_outputs[8]) & ~(layer4_outputs[4257]);
    assign layer5_outputs[1847] = ~(layer4_outputs[1138]) | (layer4_outputs[1051]);
    assign layer5_outputs[1848] = ~(layer4_outputs[3435]);
    assign layer5_outputs[1849] = (layer4_outputs[4649]) & (layer4_outputs[4152]);
    assign layer5_outputs[1850] = layer4_outputs[3073];
    assign layer5_outputs[1851] = ~(layer4_outputs[1025]);
    assign layer5_outputs[1852] = layer4_outputs[2396];
    assign layer5_outputs[1853] = layer4_outputs[4859];
    assign layer5_outputs[1854] = layer4_outputs[5059];
    assign layer5_outputs[1855] = (layer4_outputs[4229]) & ~(layer4_outputs[435]);
    assign layer5_outputs[1856] = ~(layer4_outputs[3186]) | (layer4_outputs[3288]);
    assign layer5_outputs[1857] = ~(layer4_outputs[90]) | (layer4_outputs[4961]);
    assign layer5_outputs[1858] = (layer4_outputs[1156]) & ~(layer4_outputs[2417]);
    assign layer5_outputs[1859] = (layer4_outputs[1654]) ^ (layer4_outputs[1922]);
    assign layer5_outputs[1860] = layer4_outputs[4742];
    assign layer5_outputs[1861] = 1'b1;
    assign layer5_outputs[1862] = (layer4_outputs[1390]) & ~(layer4_outputs[3457]);
    assign layer5_outputs[1863] = ~((layer4_outputs[2513]) | (layer4_outputs[29]));
    assign layer5_outputs[1864] = layer4_outputs[3144];
    assign layer5_outputs[1865] = (layer4_outputs[4388]) | (layer4_outputs[1472]);
    assign layer5_outputs[1866] = layer4_outputs[492];
    assign layer5_outputs[1867] = ~(layer4_outputs[1970]);
    assign layer5_outputs[1868] = (layer4_outputs[3349]) & (layer4_outputs[4779]);
    assign layer5_outputs[1869] = 1'b1;
    assign layer5_outputs[1870] = ~(layer4_outputs[582]) | (layer4_outputs[1769]);
    assign layer5_outputs[1871] = (layer4_outputs[1687]) & ~(layer4_outputs[4546]);
    assign layer5_outputs[1872] = (layer4_outputs[1512]) ^ (layer4_outputs[4217]);
    assign layer5_outputs[1873] = (layer4_outputs[384]) ^ (layer4_outputs[4124]);
    assign layer5_outputs[1874] = (layer4_outputs[3459]) & ~(layer4_outputs[2972]);
    assign layer5_outputs[1875] = ~(layer4_outputs[2091]);
    assign layer5_outputs[1876] = layer4_outputs[5051];
    assign layer5_outputs[1877] = layer4_outputs[2889];
    assign layer5_outputs[1878] = ~(layer4_outputs[1968]);
    assign layer5_outputs[1879] = ~(layer4_outputs[3882]) | (layer4_outputs[4077]);
    assign layer5_outputs[1880] = (layer4_outputs[4061]) & ~(layer4_outputs[1851]);
    assign layer5_outputs[1881] = ~(layer4_outputs[236]);
    assign layer5_outputs[1882] = ~(layer4_outputs[4604]);
    assign layer5_outputs[1883] = ~((layer4_outputs[2023]) & (layer4_outputs[965]));
    assign layer5_outputs[1884] = ~(layer4_outputs[1475]);
    assign layer5_outputs[1885] = ~((layer4_outputs[3940]) ^ (layer4_outputs[1261]));
    assign layer5_outputs[1886] = (layer4_outputs[940]) & ~(layer4_outputs[2078]);
    assign layer5_outputs[1887] = ~(layer4_outputs[3016]);
    assign layer5_outputs[1888] = ~(layer4_outputs[266]) | (layer4_outputs[4013]);
    assign layer5_outputs[1889] = 1'b0;
    assign layer5_outputs[1890] = layer4_outputs[628];
    assign layer5_outputs[1891] = layer4_outputs[2445];
    assign layer5_outputs[1892] = layer4_outputs[1867];
    assign layer5_outputs[1893] = layer4_outputs[3883];
    assign layer5_outputs[1894] = ~(layer4_outputs[4106]);
    assign layer5_outputs[1895] = layer4_outputs[2080];
    assign layer5_outputs[1896] = ~((layer4_outputs[283]) ^ (layer4_outputs[4873]));
    assign layer5_outputs[1897] = ~(layer4_outputs[5063]);
    assign layer5_outputs[1898] = ~(layer4_outputs[3581]);
    assign layer5_outputs[1899] = layer4_outputs[4870];
    assign layer5_outputs[1900] = ~(layer4_outputs[4815]) | (layer4_outputs[3572]);
    assign layer5_outputs[1901] = layer4_outputs[891];
    assign layer5_outputs[1902] = layer4_outputs[302];
    assign layer5_outputs[1903] = layer4_outputs[3645];
    assign layer5_outputs[1904] = ~(layer4_outputs[5095]);
    assign layer5_outputs[1905] = 1'b0;
    assign layer5_outputs[1906] = ~(layer4_outputs[1466]);
    assign layer5_outputs[1907] = ~((layer4_outputs[469]) ^ (layer4_outputs[72]));
    assign layer5_outputs[1908] = 1'b1;
    assign layer5_outputs[1909] = layer4_outputs[1161];
    assign layer5_outputs[1910] = ~((layer4_outputs[4188]) & (layer4_outputs[834]));
    assign layer5_outputs[1911] = ~(layer4_outputs[4392]);
    assign layer5_outputs[1912] = ~(layer4_outputs[1900]);
    assign layer5_outputs[1913] = ~(layer4_outputs[846]);
    assign layer5_outputs[1914] = (layer4_outputs[340]) & ~(layer4_outputs[2390]);
    assign layer5_outputs[1915] = (layer4_outputs[3922]) & ~(layer4_outputs[614]);
    assign layer5_outputs[1916] = (layer4_outputs[1834]) & (layer4_outputs[4754]);
    assign layer5_outputs[1917] = ~(layer4_outputs[4887]) | (layer4_outputs[378]);
    assign layer5_outputs[1918] = (layer4_outputs[1314]) & (layer4_outputs[992]);
    assign layer5_outputs[1919] = ~((layer4_outputs[762]) & (layer4_outputs[4850]));
    assign layer5_outputs[1920] = ~(layer4_outputs[4927]);
    assign layer5_outputs[1921] = (layer4_outputs[3872]) | (layer4_outputs[1270]);
    assign layer5_outputs[1922] = ~(layer4_outputs[2385]) | (layer4_outputs[2113]);
    assign layer5_outputs[1923] = ~(layer4_outputs[2062]) | (layer4_outputs[2259]);
    assign layer5_outputs[1924] = ~(layer4_outputs[3415]);
    assign layer5_outputs[1925] = layer4_outputs[2740];
    assign layer5_outputs[1926] = (layer4_outputs[3223]) & ~(layer4_outputs[1557]);
    assign layer5_outputs[1927] = ~(layer4_outputs[3760]);
    assign layer5_outputs[1928] = ~(layer4_outputs[3493]);
    assign layer5_outputs[1929] = ~((layer4_outputs[1038]) & (layer4_outputs[2349]));
    assign layer5_outputs[1930] = ~(layer4_outputs[4696]);
    assign layer5_outputs[1931] = layer4_outputs[3559];
    assign layer5_outputs[1932] = layer4_outputs[3412];
    assign layer5_outputs[1933] = ~(layer4_outputs[5]);
    assign layer5_outputs[1934] = (layer4_outputs[2844]) & (layer4_outputs[937]);
    assign layer5_outputs[1935] = layer4_outputs[3036];
    assign layer5_outputs[1936] = ~((layer4_outputs[4836]) ^ (layer4_outputs[2156]));
    assign layer5_outputs[1937] = 1'b0;
    assign layer5_outputs[1938] = (layer4_outputs[966]) & ~(layer4_outputs[1823]);
    assign layer5_outputs[1939] = layer4_outputs[2720];
    assign layer5_outputs[1940] = (layer4_outputs[4844]) & ~(layer4_outputs[4250]);
    assign layer5_outputs[1941] = ~(layer4_outputs[2112]);
    assign layer5_outputs[1942] = ~(layer4_outputs[672]);
    assign layer5_outputs[1943] = layer4_outputs[5003];
    assign layer5_outputs[1944] = ~((layer4_outputs[1523]) | (layer4_outputs[1674]));
    assign layer5_outputs[1945] = ~(layer4_outputs[2391]) | (layer4_outputs[3687]);
    assign layer5_outputs[1946] = ~(layer4_outputs[4869]);
    assign layer5_outputs[1947] = (layer4_outputs[1291]) | (layer4_outputs[3668]);
    assign layer5_outputs[1948] = ~(layer4_outputs[803]);
    assign layer5_outputs[1949] = ~((layer4_outputs[846]) | (layer4_outputs[3402]));
    assign layer5_outputs[1950] = (layer4_outputs[175]) ^ (layer4_outputs[4533]);
    assign layer5_outputs[1951] = layer4_outputs[3623];
    assign layer5_outputs[1952] = ~(layer4_outputs[4168]) | (layer4_outputs[1733]);
    assign layer5_outputs[1953] = ~(layer4_outputs[3942]);
    assign layer5_outputs[1954] = (layer4_outputs[1245]) | (layer4_outputs[3876]);
    assign layer5_outputs[1955] = ~(layer4_outputs[943]) | (layer4_outputs[2036]);
    assign layer5_outputs[1956] = (layer4_outputs[3878]) & ~(layer4_outputs[3870]);
    assign layer5_outputs[1957] = ~((layer4_outputs[2198]) ^ (layer4_outputs[1880]));
    assign layer5_outputs[1958] = ~((layer4_outputs[4758]) ^ (layer4_outputs[4717]));
    assign layer5_outputs[1959] = (layer4_outputs[923]) ^ (layer4_outputs[4209]);
    assign layer5_outputs[1960] = ~((layer4_outputs[2792]) & (layer4_outputs[1770]));
    assign layer5_outputs[1961] = (layer4_outputs[4627]) & (layer4_outputs[1132]);
    assign layer5_outputs[1962] = ~(layer4_outputs[4956]) | (layer4_outputs[644]);
    assign layer5_outputs[1963] = layer4_outputs[2344];
    assign layer5_outputs[1964] = layer4_outputs[1392];
    assign layer5_outputs[1965] = ~(layer4_outputs[379]);
    assign layer5_outputs[1966] = ~(layer4_outputs[3271]);
    assign layer5_outputs[1967] = ~((layer4_outputs[668]) | (layer4_outputs[4176]));
    assign layer5_outputs[1968] = layer4_outputs[1551];
    assign layer5_outputs[1969] = ~(layer4_outputs[4657]);
    assign layer5_outputs[1970] = ~((layer4_outputs[4731]) ^ (layer4_outputs[4828]));
    assign layer5_outputs[1971] = ~((layer4_outputs[1158]) ^ (layer4_outputs[3621]));
    assign layer5_outputs[1972] = ~(layer4_outputs[4808]);
    assign layer5_outputs[1973] = ~(layer4_outputs[4623]);
    assign layer5_outputs[1974] = ~(layer4_outputs[232]);
    assign layer5_outputs[1975] = layer4_outputs[1684];
    assign layer5_outputs[1976] = (layer4_outputs[1278]) & (layer4_outputs[995]);
    assign layer5_outputs[1977] = ~((layer4_outputs[280]) & (layer4_outputs[3829]));
    assign layer5_outputs[1978] = 1'b1;
    assign layer5_outputs[1979] = (layer4_outputs[1746]) ^ (layer4_outputs[886]);
    assign layer5_outputs[1980] = ~(layer4_outputs[3319]);
    assign layer5_outputs[1981] = ~(layer4_outputs[1504]) | (layer4_outputs[2679]);
    assign layer5_outputs[1982] = ~((layer4_outputs[162]) & (layer4_outputs[944]));
    assign layer5_outputs[1983] = layer4_outputs[998];
    assign layer5_outputs[1984] = ~(layer4_outputs[1341]);
    assign layer5_outputs[1985] = ~((layer4_outputs[3636]) & (layer4_outputs[1441]));
    assign layer5_outputs[1986] = ~((layer4_outputs[1649]) | (layer4_outputs[550]));
    assign layer5_outputs[1987] = ~(layer4_outputs[626]);
    assign layer5_outputs[1988] = ~((layer4_outputs[2387]) & (layer4_outputs[4606]));
    assign layer5_outputs[1989] = 1'b0;
    assign layer5_outputs[1990] = ~((layer4_outputs[2801]) | (layer4_outputs[4476]));
    assign layer5_outputs[1991] = 1'b0;
    assign layer5_outputs[1992] = ~(layer4_outputs[4431]) | (layer4_outputs[1688]);
    assign layer5_outputs[1993] = ~(layer4_outputs[3874]) | (layer4_outputs[3855]);
    assign layer5_outputs[1994] = layer4_outputs[1732];
    assign layer5_outputs[1995] = ~((layer4_outputs[445]) | (layer4_outputs[4567]));
    assign layer5_outputs[1996] = layer4_outputs[3142];
    assign layer5_outputs[1997] = (layer4_outputs[3341]) & ~(layer4_outputs[1851]);
    assign layer5_outputs[1998] = ~((layer4_outputs[1792]) & (layer4_outputs[1345]));
    assign layer5_outputs[1999] = layer4_outputs[299];
    assign layer5_outputs[2000] = ~(layer4_outputs[1630]);
    assign layer5_outputs[2001] = layer4_outputs[3761];
    assign layer5_outputs[2002] = (layer4_outputs[2195]) ^ (layer4_outputs[1033]);
    assign layer5_outputs[2003] = (layer4_outputs[4199]) ^ (layer4_outputs[888]);
    assign layer5_outputs[2004] = ~(layer4_outputs[3433]) | (layer4_outputs[4584]);
    assign layer5_outputs[2005] = 1'b0;
    assign layer5_outputs[2006] = (layer4_outputs[5076]) | (layer4_outputs[4393]);
    assign layer5_outputs[2007] = layer4_outputs[951];
    assign layer5_outputs[2008] = ~((layer4_outputs[5077]) | (layer4_outputs[2974]));
    assign layer5_outputs[2009] = 1'b1;
    assign layer5_outputs[2010] = ~((layer4_outputs[57]) & (layer4_outputs[4698]));
    assign layer5_outputs[2011] = layer4_outputs[4883];
    assign layer5_outputs[2012] = (layer4_outputs[3914]) & (layer4_outputs[2575]);
    assign layer5_outputs[2013] = 1'b0;
    assign layer5_outputs[2014] = ~(layer4_outputs[3698]);
    assign layer5_outputs[2015] = layer4_outputs[2547];
    assign layer5_outputs[2016] = ~((layer4_outputs[4298]) | (layer4_outputs[1686]));
    assign layer5_outputs[2017] = ~((layer4_outputs[3561]) & (layer4_outputs[4215]));
    assign layer5_outputs[2018] = ~(layer4_outputs[807]);
    assign layer5_outputs[2019] = (layer4_outputs[4320]) & (layer4_outputs[1763]);
    assign layer5_outputs[2020] = ~((layer4_outputs[3551]) | (layer4_outputs[3941]));
    assign layer5_outputs[2021] = layer4_outputs[2293];
    assign layer5_outputs[2022] = layer4_outputs[1149];
    assign layer5_outputs[2023] = (layer4_outputs[1654]) & ~(layer4_outputs[3490]);
    assign layer5_outputs[2024] = ~((layer4_outputs[4242]) | (layer4_outputs[613]));
    assign layer5_outputs[2025] = ~((layer4_outputs[3831]) | (layer4_outputs[2221]));
    assign layer5_outputs[2026] = ~(layer4_outputs[1197]);
    assign layer5_outputs[2027] = 1'b1;
    assign layer5_outputs[2028] = ~(layer4_outputs[2573]);
    assign layer5_outputs[2029] = layer4_outputs[882];
    assign layer5_outputs[2030] = ~(layer4_outputs[1503]);
    assign layer5_outputs[2031] = ~(layer4_outputs[4776]);
    assign layer5_outputs[2032] = ~(layer4_outputs[2806]);
    assign layer5_outputs[2033] = (layer4_outputs[591]) & ~(layer4_outputs[3437]);
    assign layer5_outputs[2034] = (layer4_outputs[444]) ^ (layer4_outputs[3534]);
    assign layer5_outputs[2035] = ~((layer4_outputs[4306]) & (layer4_outputs[4696]));
    assign layer5_outputs[2036] = ~(layer4_outputs[2731]);
    assign layer5_outputs[2037] = ~(layer4_outputs[2410]);
    assign layer5_outputs[2038] = ~(layer4_outputs[1551]);
    assign layer5_outputs[2039] = (layer4_outputs[1167]) & (layer4_outputs[2463]);
    assign layer5_outputs[2040] = (layer4_outputs[3203]) | (layer4_outputs[294]);
    assign layer5_outputs[2041] = 1'b0;
    assign layer5_outputs[2042] = ~(layer4_outputs[4032]) | (layer4_outputs[866]);
    assign layer5_outputs[2043] = layer4_outputs[1501];
    assign layer5_outputs[2044] = layer4_outputs[3661];
    assign layer5_outputs[2045] = (layer4_outputs[2189]) ^ (layer4_outputs[1476]);
    assign layer5_outputs[2046] = ~(layer4_outputs[3575]) | (layer4_outputs[4161]);
    assign layer5_outputs[2047] = layer4_outputs[335];
    assign layer5_outputs[2048] = 1'b1;
    assign layer5_outputs[2049] = ~(layer4_outputs[5101]);
    assign layer5_outputs[2050] = layer4_outputs[2946];
    assign layer5_outputs[2051] = ~(layer4_outputs[2272]);
    assign layer5_outputs[2052] = ~(layer4_outputs[4712]) | (layer4_outputs[3376]);
    assign layer5_outputs[2053] = ~((layer4_outputs[1608]) ^ (layer4_outputs[3014]));
    assign layer5_outputs[2054] = layer4_outputs[4772];
    assign layer5_outputs[2055] = (layer4_outputs[2255]) ^ (layer4_outputs[849]);
    assign layer5_outputs[2056] = (layer4_outputs[4169]) & (layer4_outputs[276]);
    assign layer5_outputs[2057] = (layer4_outputs[1317]) ^ (layer4_outputs[2703]);
    assign layer5_outputs[2058] = ~(layer4_outputs[3920]);
    assign layer5_outputs[2059] = ~(layer4_outputs[1661]) | (layer4_outputs[1298]);
    assign layer5_outputs[2060] = ~((layer4_outputs[2136]) ^ (layer4_outputs[4144]));
    assign layer5_outputs[2061] = ~(layer4_outputs[3719]);
    assign layer5_outputs[2062] = layer4_outputs[2789];
    assign layer5_outputs[2063] = layer4_outputs[1193];
    assign layer5_outputs[2064] = ~(layer4_outputs[4915]);
    assign layer5_outputs[2065] = layer4_outputs[2003];
    assign layer5_outputs[2066] = (layer4_outputs[2231]) & (layer4_outputs[985]);
    assign layer5_outputs[2067] = ~(layer4_outputs[3631]);
    assign layer5_outputs[2068] = ~(layer4_outputs[1018]);
    assign layer5_outputs[2069] = ~((layer4_outputs[3134]) | (layer4_outputs[2497]));
    assign layer5_outputs[2070] = ~((layer4_outputs[2239]) | (layer4_outputs[1299]));
    assign layer5_outputs[2071] = layer4_outputs[3245];
    assign layer5_outputs[2072] = ~(layer4_outputs[4358]) | (layer4_outputs[1950]);
    assign layer5_outputs[2073] = layer4_outputs[2635];
    assign layer5_outputs[2074] = (layer4_outputs[1872]) ^ (layer4_outputs[674]);
    assign layer5_outputs[2075] = (layer4_outputs[3585]) & (layer4_outputs[3863]);
    assign layer5_outputs[2076] = (layer4_outputs[3192]) & ~(layer4_outputs[2010]);
    assign layer5_outputs[2077] = (layer4_outputs[3456]) & ~(layer4_outputs[2168]);
    assign layer5_outputs[2078] = ~(layer4_outputs[188]);
    assign layer5_outputs[2079] = ~(layer4_outputs[4052]);
    assign layer5_outputs[2080] = layer4_outputs[1624];
    assign layer5_outputs[2081] = layer4_outputs[5040];
    assign layer5_outputs[2082] = 1'b1;
    assign layer5_outputs[2083] = layer4_outputs[1158];
    assign layer5_outputs[2084] = (layer4_outputs[4353]) ^ (layer4_outputs[4621]);
    assign layer5_outputs[2085] = (layer4_outputs[784]) & (layer4_outputs[881]);
    assign layer5_outputs[2086] = ~((layer4_outputs[3787]) & (layer4_outputs[3924]));
    assign layer5_outputs[2087] = ~(layer4_outputs[1293]) | (layer4_outputs[4588]);
    assign layer5_outputs[2088] = layer4_outputs[4638];
    assign layer5_outputs[2089] = ~(layer4_outputs[1095]);
    assign layer5_outputs[2090] = layer4_outputs[2051];
    assign layer5_outputs[2091] = layer4_outputs[1407];
    assign layer5_outputs[2092] = ~(layer4_outputs[4280]);
    assign layer5_outputs[2093] = ~(layer4_outputs[2331]);
    assign layer5_outputs[2094] = layer4_outputs[3597];
    assign layer5_outputs[2095] = ~((layer4_outputs[1000]) | (layer4_outputs[1842]));
    assign layer5_outputs[2096] = ~(layer4_outputs[3169]);
    assign layer5_outputs[2097] = (layer4_outputs[2831]) ^ (layer4_outputs[700]);
    assign layer5_outputs[2098] = ~((layer4_outputs[2165]) ^ (layer4_outputs[4703]));
    assign layer5_outputs[2099] = (layer4_outputs[3987]) & (layer4_outputs[1061]);
    assign layer5_outputs[2100] = ~(layer4_outputs[4346]);
    assign layer5_outputs[2101] = layer4_outputs[2984];
    assign layer5_outputs[2102] = ~(layer4_outputs[4120]) | (layer4_outputs[564]);
    assign layer5_outputs[2103] = ~(layer4_outputs[1418]) | (layer4_outputs[1942]);
    assign layer5_outputs[2104] = ~((layer4_outputs[1202]) & (layer4_outputs[3078]));
    assign layer5_outputs[2105] = layer4_outputs[3998];
    assign layer5_outputs[2106] = ~(layer4_outputs[4232]) | (layer4_outputs[1626]);
    assign layer5_outputs[2107] = (layer4_outputs[2539]) & ~(layer4_outputs[4263]);
    assign layer5_outputs[2108] = layer4_outputs[1499];
    assign layer5_outputs[2109] = ~(layer4_outputs[5116]);
    assign layer5_outputs[2110] = ~(layer4_outputs[1295]);
    assign layer5_outputs[2111] = 1'b0;
    assign layer5_outputs[2112] = ~(layer4_outputs[2389]);
    assign layer5_outputs[2113] = (layer4_outputs[1560]) & ~(layer4_outputs[3082]);
    assign layer5_outputs[2114] = (layer4_outputs[2245]) ^ (layer4_outputs[3358]);
    assign layer5_outputs[2115] = ~(layer4_outputs[5016]);
    assign layer5_outputs[2116] = (layer4_outputs[1920]) & ~(layer4_outputs[3651]);
    assign layer5_outputs[2117] = ~((layer4_outputs[4621]) & (layer4_outputs[2356]));
    assign layer5_outputs[2118] = ~(layer4_outputs[465]);
    assign layer5_outputs[2119] = ~(layer4_outputs[2429]);
    assign layer5_outputs[2120] = ~((layer4_outputs[1302]) | (layer4_outputs[1232]));
    assign layer5_outputs[2121] = (layer4_outputs[4938]) ^ (layer4_outputs[4457]);
    assign layer5_outputs[2122] = layer4_outputs[1853];
    assign layer5_outputs[2123] = layer4_outputs[1165];
    assign layer5_outputs[2124] = layer4_outputs[4760];
    assign layer5_outputs[2125] = (layer4_outputs[1628]) & ~(layer4_outputs[2347]);
    assign layer5_outputs[2126] = layer4_outputs[3193];
    assign layer5_outputs[2127] = layer4_outputs[588];
    assign layer5_outputs[2128] = ~((layer4_outputs[671]) | (layer4_outputs[3663]));
    assign layer5_outputs[2129] = layer4_outputs[4664];
    assign layer5_outputs[2130] = ~((layer4_outputs[1387]) ^ (layer4_outputs[2936]));
    assign layer5_outputs[2131] = ~((layer4_outputs[2001]) & (layer4_outputs[990]));
    assign layer5_outputs[2132] = (layer4_outputs[578]) | (layer4_outputs[2720]);
    assign layer5_outputs[2133] = ~(layer4_outputs[4074]);
    assign layer5_outputs[2134] = (layer4_outputs[505]) & ~(layer4_outputs[1974]);
    assign layer5_outputs[2135] = ~((layer4_outputs[4662]) | (layer4_outputs[3690]));
    assign layer5_outputs[2136] = ~(layer4_outputs[3728]) | (layer4_outputs[2680]);
    assign layer5_outputs[2137] = ~(layer4_outputs[2484]) | (layer4_outputs[2716]);
    assign layer5_outputs[2138] = layer4_outputs[4567];
    assign layer5_outputs[2139] = ~((layer4_outputs[2600]) & (layer4_outputs[239]));
    assign layer5_outputs[2140] = (layer4_outputs[4762]) & ~(layer4_outputs[3693]);
    assign layer5_outputs[2141] = layer4_outputs[2194];
    assign layer5_outputs[2142] = ~((layer4_outputs[687]) ^ (layer4_outputs[1070]));
    assign layer5_outputs[2143] = 1'b1;
    assign layer5_outputs[2144] = ~((layer4_outputs[4186]) & (layer4_outputs[3012]));
    assign layer5_outputs[2145] = layer4_outputs[1996];
    assign layer5_outputs[2146] = ~(layer4_outputs[4890]);
    assign layer5_outputs[2147] = ~(layer4_outputs[4336]) | (layer4_outputs[646]);
    assign layer5_outputs[2148] = layer4_outputs[2736];
    assign layer5_outputs[2149] = (layer4_outputs[2387]) | (layer4_outputs[977]);
    assign layer5_outputs[2150] = ~(layer4_outputs[3733]);
    assign layer5_outputs[2151] = ~(layer4_outputs[3280]);
    assign layer5_outputs[2152] = ~(layer4_outputs[2669]);
    assign layer5_outputs[2153] = layer4_outputs[4070];
    assign layer5_outputs[2154] = layer4_outputs[4175];
    assign layer5_outputs[2155] = (layer4_outputs[1627]) | (layer4_outputs[3291]);
    assign layer5_outputs[2156] = layer4_outputs[3531];
    assign layer5_outputs[2157] = (layer4_outputs[4825]) ^ (layer4_outputs[2315]);
    assign layer5_outputs[2158] = layer4_outputs[1188];
    assign layer5_outputs[2159] = (layer4_outputs[2636]) | (layer4_outputs[4175]);
    assign layer5_outputs[2160] = layer4_outputs[3129];
    assign layer5_outputs[2161] = ~(layer4_outputs[4226]);
    assign layer5_outputs[2162] = ~(layer4_outputs[3126]);
    assign layer5_outputs[2163] = layer4_outputs[414];
    assign layer5_outputs[2164] = 1'b1;
    assign layer5_outputs[2165] = 1'b0;
    assign layer5_outputs[2166] = layer4_outputs[4676];
    assign layer5_outputs[2167] = (layer4_outputs[3167]) | (layer4_outputs[492]);
    assign layer5_outputs[2168] = (layer4_outputs[835]) | (layer4_outputs[5114]);
    assign layer5_outputs[2169] = layer4_outputs[1146];
    assign layer5_outputs[2170] = layer4_outputs[3675];
    assign layer5_outputs[2171] = ~(layer4_outputs[1899]) | (layer4_outputs[1782]);
    assign layer5_outputs[2172] = ~(layer4_outputs[1900]);
    assign layer5_outputs[2173] = ~(layer4_outputs[740]);
    assign layer5_outputs[2174] = ~((layer4_outputs[1698]) ^ (layer4_outputs[996]));
    assign layer5_outputs[2175] = ~((layer4_outputs[697]) | (layer4_outputs[4780]));
    assign layer5_outputs[2176] = ~(layer4_outputs[1781]);
    assign layer5_outputs[2177] = ~(layer4_outputs[2975]) | (layer4_outputs[4774]);
    assign layer5_outputs[2178] = (layer4_outputs[1256]) | (layer4_outputs[269]);
    assign layer5_outputs[2179] = (layer4_outputs[4661]) & (layer4_outputs[2146]);
    assign layer5_outputs[2180] = ~(layer4_outputs[4216]);
    assign layer5_outputs[2181] = layer4_outputs[4631];
    assign layer5_outputs[2182] = (layer4_outputs[1455]) & ~(layer4_outputs[4284]);
    assign layer5_outputs[2183] = ~(layer4_outputs[4329]);
    assign layer5_outputs[2184] = (layer4_outputs[4750]) & (layer4_outputs[4693]);
    assign layer5_outputs[2185] = ~(layer4_outputs[2619]);
    assign layer5_outputs[2186] = ~((layer4_outputs[1030]) & (layer4_outputs[3371]));
    assign layer5_outputs[2187] = layer4_outputs[587];
    assign layer5_outputs[2188] = ~(layer4_outputs[3389]);
    assign layer5_outputs[2189] = ~(layer4_outputs[2836]);
    assign layer5_outputs[2190] = layer4_outputs[1111];
    assign layer5_outputs[2191] = layer4_outputs[1718];
    assign layer5_outputs[2192] = (layer4_outputs[2592]) & ~(layer4_outputs[1355]);
    assign layer5_outputs[2193] = ~(layer4_outputs[4406]) | (layer4_outputs[5099]);
    assign layer5_outputs[2194] = ~(layer4_outputs[33]);
    assign layer5_outputs[2195] = (layer4_outputs[1662]) & (layer4_outputs[4429]);
    assign layer5_outputs[2196] = ~(layer4_outputs[2660]);
    assign layer5_outputs[2197] = (layer4_outputs[1834]) ^ (layer4_outputs[2101]);
    assign layer5_outputs[2198] = ~(layer4_outputs[2177]);
    assign layer5_outputs[2199] = layer4_outputs[2501];
    assign layer5_outputs[2200] = layer4_outputs[4317];
    assign layer5_outputs[2201] = ~(layer4_outputs[2244]);
    assign layer5_outputs[2202] = 1'b1;
    assign layer5_outputs[2203] = layer4_outputs[1347];
    assign layer5_outputs[2204] = ~(layer4_outputs[4802]);
    assign layer5_outputs[2205] = ~(layer4_outputs[117]);
    assign layer5_outputs[2206] = 1'b1;
    assign layer5_outputs[2207] = layer4_outputs[2443];
    assign layer5_outputs[2208] = ~((layer4_outputs[126]) ^ (layer4_outputs[2133]));
    assign layer5_outputs[2209] = ~((layer4_outputs[2303]) & (layer4_outputs[3161]));
    assign layer5_outputs[2210] = ~(layer4_outputs[3565]) | (layer4_outputs[3120]);
    assign layer5_outputs[2211] = (layer4_outputs[281]) ^ (layer4_outputs[2209]);
    assign layer5_outputs[2212] = ~(layer4_outputs[312]);
    assign layer5_outputs[2213] = layer4_outputs[4266];
    assign layer5_outputs[2214] = layer4_outputs[4121];
    assign layer5_outputs[2215] = layer4_outputs[1224];
    assign layer5_outputs[2216] = (layer4_outputs[1043]) & ~(layer4_outputs[3946]);
    assign layer5_outputs[2217] = ~(layer4_outputs[4622]);
    assign layer5_outputs[2218] = ~((layer4_outputs[4381]) | (layer4_outputs[5083]));
    assign layer5_outputs[2219] = (layer4_outputs[147]) | (layer4_outputs[1840]);
    assign layer5_outputs[2220] = ~(layer4_outputs[3875]) | (layer4_outputs[794]);
    assign layer5_outputs[2221] = ~(layer4_outputs[3615]) | (layer4_outputs[2400]);
    assign layer5_outputs[2222] = ~(layer4_outputs[2649]);
    assign layer5_outputs[2223] = ~(layer4_outputs[4547]) | (layer4_outputs[1810]);
    assign layer5_outputs[2224] = layer4_outputs[4874];
    assign layer5_outputs[2225] = (layer4_outputs[4111]) ^ (layer4_outputs[3809]);
    assign layer5_outputs[2226] = ~(layer4_outputs[1224]);
    assign layer5_outputs[2227] = layer4_outputs[2412];
    assign layer5_outputs[2228] = layer4_outputs[899];
    assign layer5_outputs[2229] = (layer4_outputs[4543]) ^ (layer4_outputs[3682]);
    assign layer5_outputs[2230] = ~((layer4_outputs[4005]) ^ (layer4_outputs[4577]));
    assign layer5_outputs[2231] = layer4_outputs[3118];
    assign layer5_outputs[2232] = (layer4_outputs[2659]) ^ (layer4_outputs[3835]);
    assign layer5_outputs[2233] = (layer4_outputs[2576]) ^ (layer4_outputs[2064]);
    assign layer5_outputs[2234] = ~(layer4_outputs[1317]);
    assign layer5_outputs[2235] = layer4_outputs[5081];
    assign layer5_outputs[2236] = ~(layer4_outputs[4476]) | (layer4_outputs[1821]);
    assign layer5_outputs[2237] = layer4_outputs[3881];
    assign layer5_outputs[2238] = ~(layer4_outputs[3848]);
    assign layer5_outputs[2239] = layer4_outputs[3159];
    assign layer5_outputs[2240] = 1'b0;
    assign layer5_outputs[2241] = (layer4_outputs[4834]) & (layer4_outputs[3735]);
    assign layer5_outputs[2242] = ~((layer4_outputs[4038]) | (layer4_outputs[2000]));
    assign layer5_outputs[2243] = (layer4_outputs[4148]) & ~(layer4_outputs[3464]);
    assign layer5_outputs[2244] = (layer4_outputs[1046]) | (layer4_outputs[1808]);
    assign layer5_outputs[2245] = (layer4_outputs[4984]) ^ (layer4_outputs[4624]);
    assign layer5_outputs[2246] = 1'b0;
    assign layer5_outputs[2247] = layer4_outputs[4451];
    assign layer5_outputs[2248] = ~(layer4_outputs[374]);
    assign layer5_outputs[2249] = ~(layer4_outputs[3147]);
    assign layer5_outputs[2250] = (layer4_outputs[322]) & ~(layer4_outputs[2813]);
    assign layer5_outputs[2251] = ~(layer4_outputs[2644]) | (layer4_outputs[2059]);
    assign layer5_outputs[2252] = layer4_outputs[4964];
    assign layer5_outputs[2253] = layer4_outputs[4974];
    assign layer5_outputs[2254] = (layer4_outputs[2160]) & ~(layer4_outputs[317]);
    assign layer5_outputs[2255] = 1'b1;
    assign layer5_outputs[2256] = ~((layer4_outputs[4445]) & (layer4_outputs[2509]));
    assign layer5_outputs[2257] = ~(layer4_outputs[1519]) | (layer4_outputs[4531]);
    assign layer5_outputs[2258] = ~((layer4_outputs[1745]) | (layer4_outputs[4588]));
    assign layer5_outputs[2259] = ~(layer4_outputs[4843]);
    assign layer5_outputs[2260] = (layer4_outputs[4687]) & ~(layer4_outputs[1147]);
    assign layer5_outputs[2261] = layer4_outputs[4539];
    assign layer5_outputs[2262] = layer4_outputs[3962];
    assign layer5_outputs[2263] = ~(layer4_outputs[5064]);
    assign layer5_outputs[2264] = ~((layer4_outputs[5056]) ^ (layer4_outputs[424]));
    assign layer5_outputs[2265] = ~(layer4_outputs[1311]);
    assign layer5_outputs[2266] = (layer4_outputs[1253]) & ~(layer4_outputs[3181]);
    assign layer5_outputs[2267] = (layer4_outputs[2479]) & (layer4_outputs[481]);
    assign layer5_outputs[2268] = (layer4_outputs[2093]) ^ (layer4_outputs[1326]);
    assign layer5_outputs[2269] = 1'b1;
    assign layer5_outputs[2270] = (layer4_outputs[5009]) | (layer4_outputs[1838]);
    assign layer5_outputs[2271] = ~((layer4_outputs[2752]) | (layer4_outputs[986]));
    assign layer5_outputs[2272] = ~(layer4_outputs[1144]);
    assign layer5_outputs[2273] = ~(layer4_outputs[3234]) | (layer4_outputs[534]);
    assign layer5_outputs[2274] = ~(layer4_outputs[4818]) | (layer4_outputs[2787]);
    assign layer5_outputs[2275] = ~((layer4_outputs[5104]) | (layer4_outputs[1935]));
    assign layer5_outputs[2276] = (layer4_outputs[4753]) | (layer4_outputs[959]);
    assign layer5_outputs[2277] = ~(layer4_outputs[2882]);
    assign layer5_outputs[2278] = ~((layer4_outputs[2858]) & (layer4_outputs[1128]));
    assign layer5_outputs[2279] = layer4_outputs[4498];
    assign layer5_outputs[2280] = layer4_outputs[4634];
    assign layer5_outputs[2281] = ~((layer4_outputs[2232]) ^ (layer4_outputs[326]));
    assign layer5_outputs[2282] = ~(layer4_outputs[2260]);
    assign layer5_outputs[2283] = layer4_outputs[4775];
    assign layer5_outputs[2284] = (layer4_outputs[3212]) ^ (layer4_outputs[2289]);
    assign layer5_outputs[2285] = (layer4_outputs[118]) & ~(layer4_outputs[2793]);
    assign layer5_outputs[2286] = ~((layer4_outputs[3917]) & (layer4_outputs[760]));
    assign layer5_outputs[2287] = ~((layer4_outputs[4583]) ^ (layer4_outputs[1115]));
    assign layer5_outputs[2288] = (layer4_outputs[2073]) ^ (layer4_outputs[1318]);
    assign layer5_outputs[2289] = layer4_outputs[443];
    assign layer5_outputs[2290] = ~((layer4_outputs[3137]) | (layer4_outputs[4650]));
    assign layer5_outputs[2291] = ~((layer4_outputs[1776]) | (layer4_outputs[1868]));
    assign layer5_outputs[2292] = ~((layer4_outputs[3755]) & (layer4_outputs[3460]));
    assign layer5_outputs[2293] = (layer4_outputs[300]) ^ (layer4_outputs[4233]);
    assign layer5_outputs[2294] = layer4_outputs[4515];
    assign layer5_outputs[2295] = ~((layer4_outputs[2944]) ^ (layer4_outputs[1978]));
    assign layer5_outputs[2296] = layer4_outputs[2151];
    assign layer5_outputs[2297] = ~(layer4_outputs[3880]);
    assign layer5_outputs[2298] = layer4_outputs[4208];
    assign layer5_outputs[2299] = layer4_outputs[4727];
    assign layer5_outputs[2300] = layer4_outputs[3168];
    assign layer5_outputs[2301] = ~(layer4_outputs[2468]);
    assign layer5_outputs[2302] = ~(layer4_outputs[4975]);
    assign layer5_outputs[2303] = ~((layer4_outputs[3596]) & (layer4_outputs[2757]));
    assign layer5_outputs[2304] = layer4_outputs[4897];
    assign layer5_outputs[2305] = ~(layer4_outputs[471]);
    assign layer5_outputs[2306] = (layer4_outputs[4541]) ^ (layer4_outputs[4413]);
    assign layer5_outputs[2307] = ~(layer4_outputs[3715]);
    assign layer5_outputs[2308] = ~((layer4_outputs[4505]) ^ (layer4_outputs[3096]));
    assign layer5_outputs[2309] = (layer4_outputs[567]) | (layer4_outputs[715]);
    assign layer5_outputs[2310] = ~(layer4_outputs[177]);
    assign layer5_outputs[2311] = ~(layer4_outputs[3068]);
    assign layer5_outputs[2312] = (layer4_outputs[2409]) | (layer4_outputs[4030]);
    assign layer5_outputs[2313] = layer4_outputs[4348];
    assign layer5_outputs[2314] = layer4_outputs[1712];
    assign layer5_outputs[2315] = (layer4_outputs[3346]) & ~(layer4_outputs[3511]);
    assign layer5_outputs[2316] = layer4_outputs[611];
    assign layer5_outputs[2317] = ~(layer4_outputs[4858]);
    assign layer5_outputs[2318] = layer4_outputs[315];
    assign layer5_outputs[2319] = layer4_outputs[4358];
    assign layer5_outputs[2320] = layer4_outputs[5006];
    assign layer5_outputs[2321] = layer4_outputs[4127];
    assign layer5_outputs[2322] = layer4_outputs[3446];
    assign layer5_outputs[2323] = (layer4_outputs[5020]) & (layer4_outputs[3730]);
    assign layer5_outputs[2324] = (layer4_outputs[3225]) | (layer4_outputs[1477]);
    assign layer5_outputs[2325] = (layer4_outputs[195]) & ~(layer4_outputs[237]);
    assign layer5_outputs[2326] = layer4_outputs[3873];
    assign layer5_outputs[2327] = layer4_outputs[1594];
    assign layer5_outputs[2328] = ~(layer4_outputs[1711]);
    assign layer5_outputs[2329] = ~(layer4_outputs[935]);
    assign layer5_outputs[2330] = ~(layer4_outputs[4836]);
    assign layer5_outputs[2331] = (layer4_outputs[3420]) | (layer4_outputs[157]);
    assign layer5_outputs[2332] = 1'b1;
    assign layer5_outputs[2333] = ~(layer4_outputs[5044]);
    assign layer5_outputs[2334] = ~((layer4_outputs[1648]) & (layer4_outputs[2195]));
    assign layer5_outputs[2335] = ~((layer4_outputs[3013]) | (layer4_outputs[1864]));
    assign layer5_outputs[2336] = ~(layer4_outputs[987]);
    assign layer5_outputs[2337] = (layer4_outputs[1362]) ^ (layer4_outputs[4122]);
    assign layer5_outputs[2338] = (layer4_outputs[5063]) & ~(layer4_outputs[1041]);
    assign layer5_outputs[2339] = ~(layer4_outputs[500]);
    assign layer5_outputs[2340] = (layer4_outputs[4122]) ^ (layer4_outputs[4568]);
    assign layer5_outputs[2341] = layer4_outputs[2777];
    assign layer5_outputs[2342] = layer4_outputs[766];
    assign layer5_outputs[2343] = ~(layer4_outputs[538]) | (layer4_outputs[1936]);
    assign layer5_outputs[2344] = ~(layer4_outputs[1967]);
    assign layer5_outputs[2345] = ~((layer4_outputs[4675]) | (layer4_outputs[3865]));
    assign layer5_outputs[2346] = layer4_outputs[3512];
    assign layer5_outputs[2347] = ~(layer4_outputs[1922]);
    assign layer5_outputs[2348] = ~((layer4_outputs[3343]) & (layer4_outputs[1721]));
    assign layer5_outputs[2349] = 1'b1;
    assign layer5_outputs[2350] = ~((layer4_outputs[2037]) | (layer4_outputs[2339]));
    assign layer5_outputs[2351] = ~(layer4_outputs[3632]) | (layer4_outputs[4806]);
    assign layer5_outputs[2352] = ~(layer4_outputs[1007]) | (layer4_outputs[1112]);
    assign layer5_outputs[2353] = ~(layer4_outputs[4172]);
    assign layer5_outputs[2354] = ~((layer4_outputs[4766]) & (layer4_outputs[2359]));
    assign layer5_outputs[2355] = ~(layer4_outputs[1964]);
    assign layer5_outputs[2356] = (layer4_outputs[1006]) & ~(layer4_outputs[820]);
    assign layer5_outputs[2357] = 1'b0;
    assign layer5_outputs[2358] = layer4_outputs[1925];
    assign layer5_outputs[2359] = ~(layer4_outputs[3798]);
    assign layer5_outputs[2360] = layer4_outputs[4273];
    assign layer5_outputs[2361] = layer4_outputs[1565];
    assign layer5_outputs[2362] = layer4_outputs[2338];
    assign layer5_outputs[2363] = layer4_outputs[425];
    assign layer5_outputs[2364] = layer4_outputs[5078];
    assign layer5_outputs[2365] = ~(layer4_outputs[2207]);
    assign layer5_outputs[2366] = ~((layer4_outputs[3561]) ^ (layer4_outputs[2668]));
    assign layer5_outputs[2367] = ~(layer4_outputs[2306]);
    assign layer5_outputs[2368] = ~((layer4_outputs[4852]) ^ (layer4_outputs[4410]));
    assign layer5_outputs[2369] = layer4_outputs[3799];
    assign layer5_outputs[2370] = ~(layer4_outputs[2687]);
    assign layer5_outputs[2371] = (layer4_outputs[4091]) ^ (layer4_outputs[1673]);
    assign layer5_outputs[2372] = ~(layer4_outputs[3078]);
    assign layer5_outputs[2373] = (layer4_outputs[310]) & ~(layer4_outputs[308]);
    assign layer5_outputs[2374] = (layer4_outputs[2787]) & ~(layer4_outputs[1011]);
    assign layer5_outputs[2375] = (layer4_outputs[4688]) & ~(layer4_outputs[3785]);
    assign layer5_outputs[2376] = ~(layer4_outputs[3927]);
    assign layer5_outputs[2377] = layer4_outputs[4859];
    assign layer5_outputs[2378] = ~(layer4_outputs[3982]);
    assign layer5_outputs[2379] = (layer4_outputs[1690]) & ~(layer4_outputs[2421]);
    assign layer5_outputs[2380] = layer4_outputs[1796];
    assign layer5_outputs[2381] = ~(layer4_outputs[3542]);
    assign layer5_outputs[2382] = layer4_outputs[5010];
    assign layer5_outputs[2383] = ~(layer4_outputs[2952]);
    assign layer5_outputs[2384] = (layer4_outputs[745]) ^ (layer4_outputs[4787]);
    assign layer5_outputs[2385] = layer4_outputs[1075];
    assign layer5_outputs[2386] = layer4_outputs[4397];
    assign layer5_outputs[2387] = ~((layer4_outputs[1447]) & (layer4_outputs[2916]));
    assign layer5_outputs[2388] = layer4_outputs[565];
    assign layer5_outputs[2389] = ~(layer4_outputs[3933]) | (layer4_outputs[4302]);
    assign layer5_outputs[2390] = ~(layer4_outputs[1298]);
    assign layer5_outputs[2391] = ~(layer4_outputs[3838]);
    assign layer5_outputs[2392] = (layer4_outputs[3003]) ^ (layer4_outputs[2256]);
    assign layer5_outputs[2393] = layer4_outputs[1572];
    assign layer5_outputs[2394] = layer4_outputs[3567];
    assign layer5_outputs[2395] = (layer4_outputs[1753]) & (layer4_outputs[4678]);
    assign layer5_outputs[2396] = (layer4_outputs[144]) | (layer4_outputs[3553]);
    assign layer5_outputs[2397] = ~(layer4_outputs[3263]);
    assign layer5_outputs[2398] = (layer4_outputs[4087]) | (layer4_outputs[367]);
    assign layer5_outputs[2399] = ~(layer4_outputs[5116]);
    assign layer5_outputs[2400] = ~(layer4_outputs[1130]);
    assign layer5_outputs[2401] = ~((layer4_outputs[968]) & (layer4_outputs[2692]));
    assign layer5_outputs[2402] = ~(layer4_outputs[3239]) | (layer4_outputs[1653]);
    assign layer5_outputs[2403] = layer4_outputs[2058];
    assign layer5_outputs[2404] = layer4_outputs[4973];
    assign layer5_outputs[2405] = layer4_outputs[3752];
    assign layer5_outputs[2406] = (layer4_outputs[545]) ^ (layer4_outputs[3559]);
    assign layer5_outputs[2407] = ~(layer4_outputs[1827]);
    assign layer5_outputs[2408] = layer4_outputs[524];
    assign layer5_outputs[2409] = ~(layer4_outputs[3791]);
    assign layer5_outputs[2410] = (layer4_outputs[3844]) & ~(layer4_outputs[3176]);
    assign layer5_outputs[2411] = ~(layer4_outputs[1927]) | (layer4_outputs[1803]);
    assign layer5_outputs[2412] = (layer4_outputs[4854]) | (layer4_outputs[116]);
    assign layer5_outputs[2413] = 1'b1;
    assign layer5_outputs[2414] = ~((layer4_outputs[66]) ^ (layer4_outputs[82]));
    assign layer5_outputs[2415] = ~((layer4_outputs[4373]) & (layer4_outputs[3945]));
    assign layer5_outputs[2416] = ~(layer4_outputs[2082]);
    assign layer5_outputs[2417] = ~(layer4_outputs[4435]) | (layer4_outputs[3154]);
    assign layer5_outputs[2418] = (layer4_outputs[1191]) & (layer4_outputs[5072]);
    assign layer5_outputs[2419] = ~(layer4_outputs[48]);
    assign layer5_outputs[2420] = ~((layer4_outputs[3308]) | (layer4_outputs[4506]));
    assign layer5_outputs[2421] = (layer4_outputs[4405]) | (layer4_outputs[5080]);
    assign layer5_outputs[2422] = 1'b0;
    assign layer5_outputs[2423] = 1'b0;
    assign layer5_outputs[2424] = layer4_outputs[4124];
    assign layer5_outputs[2425] = layer4_outputs[3671];
    assign layer5_outputs[2426] = ~(layer4_outputs[3737]);
    assign layer5_outputs[2427] = layer4_outputs[3064];
    assign layer5_outputs[2428] = 1'b1;
    assign layer5_outputs[2429] = ~(layer4_outputs[4285]) | (layer4_outputs[3059]);
    assign layer5_outputs[2430] = layer4_outputs[287];
    assign layer5_outputs[2431] = layer4_outputs[1239];
    assign layer5_outputs[2432] = ~(layer4_outputs[1208]);
    assign layer5_outputs[2433] = layer4_outputs[4581];
    assign layer5_outputs[2434] = layer4_outputs[1119];
    assign layer5_outputs[2435] = layer4_outputs[4179];
    assign layer5_outputs[2436] = layer4_outputs[1403];
    assign layer5_outputs[2437] = ~((layer4_outputs[1028]) ^ (layer4_outputs[1088]));
    assign layer5_outputs[2438] = (layer4_outputs[1214]) ^ (layer4_outputs[3995]);
    assign layer5_outputs[2439] = layer4_outputs[2400];
    assign layer5_outputs[2440] = ~(layer4_outputs[1513]);
    assign layer5_outputs[2441] = ~(layer4_outputs[4826]);
    assign layer5_outputs[2442] = (layer4_outputs[1506]) & ~(layer4_outputs[78]);
    assign layer5_outputs[2443] = layer4_outputs[2917];
    assign layer5_outputs[2444] = (layer4_outputs[2814]) | (layer4_outputs[3806]);
    assign layer5_outputs[2445] = (layer4_outputs[2076]) ^ (layer4_outputs[2751]);
    assign layer5_outputs[2446] = (layer4_outputs[4674]) & ~(layer4_outputs[4247]);
    assign layer5_outputs[2447] = ~((layer4_outputs[283]) & (layer4_outputs[491]));
    assign layer5_outputs[2448] = (layer4_outputs[1060]) & ~(layer4_outputs[1494]);
    assign layer5_outputs[2449] = 1'b0;
    assign layer5_outputs[2450] = layer4_outputs[3929];
    assign layer5_outputs[2451] = layer4_outputs[870];
    assign layer5_outputs[2452] = layer4_outputs[2249];
    assign layer5_outputs[2453] = layer4_outputs[2683];
    assign layer5_outputs[2454] = ~(layer4_outputs[4004]);
    assign layer5_outputs[2455] = ~((layer4_outputs[4297]) | (layer4_outputs[2222]));
    assign layer5_outputs[2456] = ~(layer4_outputs[1470]);
    assign layer5_outputs[2457] = layer4_outputs[3230];
    assign layer5_outputs[2458] = ~(layer4_outputs[4396]);
    assign layer5_outputs[2459] = (layer4_outputs[3795]) ^ (layer4_outputs[1718]);
    assign layer5_outputs[2460] = (layer4_outputs[453]) & (layer4_outputs[974]);
    assign layer5_outputs[2461] = (layer4_outputs[4426]) | (layer4_outputs[714]);
    assign layer5_outputs[2462] = ~(layer4_outputs[2923]) | (layer4_outputs[320]);
    assign layer5_outputs[2463] = ~((layer4_outputs[54]) | (layer4_outputs[1031]));
    assign layer5_outputs[2464] = 1'b0;
    assign layer5_outputs[2465] = layer4_outputs[3022];
    assign layer5_outputs[2466] = ~(layer4_outputs[2028]) | (layer4_outputs[4885]);
    assign layer5_outputs[2467] = ~(layer4_outputs[1497]);
    assign layer5_outputs[2468] = ~(layer4_outputs[2691]);
    assign layer5_outputs[2469] = ~(layer4_outputs[2312]);
    assign layer5_outputs[2470] = ~((layer4_outputs[1915]) ^ (layer4_outputs[3626]));
    assign layer5_outputs[2471] = (layer4_outputs[4632]) & (layer4_outputs[2430]);
    assign layer5_outputs[2472] = ~(layer4_outputs[2926]);
    assign layer5_outputs[2473] = ~(layer4_outputs[67]) | (layer4_outputs[2968]);
    assign layer5_outputs[2474] = layer4_outputs[2616];
    assign layer5_outputs[2475] = ~(layer4_outputs[2708]);
    assign layer5_outputs[2476] = (layer4_outputs[326]) & (layer4_outputs[4423]);
    assign layer5_outputs[2477] = (layer4_outputs[4276]) & (layer4_outputs[1726]);
    assign layer5_outputs[2478] = ~(layer4_outputs[3345]);
    assign layer5_outputs[2479] = layer4_outputs[5015];
    assign layer5_outputs[2480] = layer4_outputs[3948];
    assign layer5_outputs[2481] = ~((layer4_outputs[3067]) & (layer4_outputs[2490]));
    assign layer5_outputs[2482] = layer4_outputs[360];
    assign layer5_outputs[2483] = ~((layer4_outputs[3937]) & (layer4_outputs[2205]));
    assign layer5_outputs[2484] = ~((layer4_outputs[4658]) & (layer4_outputs[124]));
    assign layer5_outputs[2485] = ~(layer4_outputs[1914]);
    assign layer5_outputs[2486] = layer4_outputs[397];
    assign layer5_outputs[2487] = ~(layer4_outputs[5110]);
    assign layer5_outputs[2488] = (layer4_outputs[4344]) & ~(layer4_outputs[787]);
    assign layer5_outputs[2489] = ~(layer4_outputs[2457]);
    assign layer5_outputs[2490] = ~((layer4_outputs[1633]) ^ (layer4_outputs[4863]));
    assign layer5_outputs[2491] = 1'b1;
    assign layer5_outputs[2492] = ~(layer4_outputs[3335]);
    assign layer5_outputs[2493] = ~(layer4_outputs[2797]);
    assign layer5_outputs[2494] = (layer4_outputs[1045]) & (layer4_outputs[260]);
    assign layer5_outputs[2495] = ~((layer4_outputs[16]) & (layer4_outputs[3215]));
    assign layer5_outputs[2496] = (layer4_outputs[366]) & ~(layer4_outputs[895]);
    assign layer5_outputs[2497] = ~((layer4_outputs[900]) | (layer4_outputs[2811]));
    assign layer5_outputs[2498] = ~(layer4_outputs[2340]);
    assign layer5_outputs[2499] = (layer4_outputs[3466]) & ~(layer4_outputs[4522]);
    assign layer5_outputs[2500] = layer4_outputs[1497];
    assign layer5_outputs[2501] = (layer4_outputs[3419]) ^ (layer4_outputs[4055]);
    assign layer5_outputs[2502] = ~(layer4_outputs[4759]);
    assign layer5_outputs[2503] = (layer4_outputs[4952]) & ~(layer4_outputs[1807]);
    assign layer5_outputs[2504] = ~(layer4_outputs[4173]);
    assign layer5_outputs[2505] = ~(layer4_outputs[3024]) | (layer4_outputs[3080]);
    assign layer5_outputs[2506] = layer4_outputs[3827];
    assign layer5_outputs[2507] = ~(layer4_outputs[1725]);
    assign layer5_outputs[2508] = (layer4_outputs[4445]) & (layer4_outputs[1399]);
    assign layer5_outputs[2509] = ~(layer4_outputs[2657]);
    assign layer5_outputs[2510] = ~(layer4_outputs[3936]);
    assign layer5_outputs[2511] = ~((layer4_outputs[1349]) | (layer4_outputs[4025]));
    assign layer5_outputs[2512] = (layer4_outputs[2654]) & ~(layer4_outputs[3293]);
    assign layer5_outputs[2513] = layer4_outputs[1165];
    assign layer5_outputs[2514] = (layer4_outputs[192]) | (layer4_outputs[4295]);
    assign layer5_outputs[2515] = ~(layer4_outputs[4227]);
    assign layer5_outputs[2516] = (layer4_outputs[551]) & (layer4_outputs[4609]);
    assign layer5_outputs[2517] = (layer4_outputs[2522]) & (layer4_outputs[2853]);
    assign layer5_outputs[2518] = layer4_outputs[936];
    assign layer5_outputs[2519] = layer4_outputs[2211];
    assign layer5_outputs[2520] = (layer4_outputs[2937]) & ~(layer4_outputs[3248]);
    assign layer5_outputs[2521] = layer4_outputs[1550];
    assign layer5_outputs[2522] = (layer4_outputs[3835]) & ~(layer4_outputs[3364]);
    assign layer5_outputs[2523] = (layer4_outputs[1658]) & ~(layer4_outputs[4700]);
    assign layer5_outputs[2524] = layer4_outputs[32];
    assign layer5_outputs[2525] = (layer4_outputs[1924]) ^ (layer4_outputs[17]);
    assign layer5_outputs[2526] = (layer4_outputs[172]) ^ (layer4_outputs[685]);
    assign layer5_outputs[2527] = ~((layer4_outputs[3620]) ^ (layer4_outputs[1027]));
    assign layer5_outputs[2528] = ~(layer4_outputs[718]);
    assign layer5_outputs[2529] = ~(layer4_outputs[3951]);
    assign layer5_outputs[2530] = (layer4_outputs[4924]) & ~(layer4_outputs[3654]);
    assign layer5_outputs[2531] = 1'b0;
    assign layer5_outputs[2532] = (layer4_outputs[79]) & (layer4_outputs[4689]);
    assign layer5_outputs[2533] = ~(layer4_outputs[1891]);
    assign layer5_outputs[2534] = ~(layer4_outputs[1282]) | (layer4_outputs[2541]);
    assign layer5_outputs[2535] = layer4_outputs[2771];
    assign layer5_outputs[2536] = ~(layer4_outputs[1067]);
    assign layer5_outputs[2537] = ~(layer4_outputs[3088]);
    assign layer5_outputs[2538] = ~(layer4_outputs[2090]);
    assign layer5_outputs[2539] = (layer4_outputs[3366]) & (layer4_outputs[4189]);
    assign layer5_outputs[2540] = (layer4_outputs[1720]) & ~(layer4_outputs[4936]);
    assign layer5_outputs[2541] = (layer4_outputs[85]) & ~(layer4_outputs[4155]);
    assign layer5_outputs[2542] = layer4_outputs[3643];
    assign layer5_outputs[2543] = ~(layer4_outputs[3695]) | (layer4_outputs[2480]);
    assign layer5_outputs[2544] = ~(layer4_outputs[28]) | (layer4_outputs[922]);
    assign layer5_outputs[2545] = layer4_outputs[1682];
    assign layer5_outputs[2546] = 1'b1;
    assign layer5_outputs[2547] = layer4_outputs[2547];
    assign layer5_outputs[2548] = layer4_outputs[582];
    assign layer5_outputs[2549] = ~((layer4_outputs[2180]) & (layer4_outputs[957]));
    assign layer5_outputs[2550] = layer4_outputs[456];
    assign layer5_outputs[2551] = ~((layer4_outputs[4934]) | (layer4_outputs[106]));
    assign layer5_outputs[2552] = ~(layer4_outputs[3234]) | (layer4_outputs[695]);
    assign layer5_outputs[2553] = layer4_outputs[2318];
    assign layer5_outputs[2554] = ~(layer4_outputs[4686]);
    assign layer5_outputs[2555] = (layer4_outputs[2129]) & ~(layer4_outputs[1411]);
    assign layer5_outputs[2556] = layer4_outputs[902];
    assign layer5_outputs[2557] = (layer4_outputs[4222]) | (layer4_outputs[2205]);
    assign layer5_outputs[2558] = ~(layer4_outputs[4530]);
    assign layer5_outputs[2559] = layer4_outputs[1221];
    assign layer5_outputs[2560] = (layer4_outputs[1597]) & ~(layer4_outputs[4244]);
    assign layer5_outputs[2561] = layer4_outputs[866];
    assign layer5_outputs[2562] = ~(layer4_outputs[3601]) | (layer4_outputs[2945]);
    assign layer5_outputs[2563] = (layer4_outputs[3718]) ^ (layer4_outputs[1824]);
    assign layer5_outputs[2564] = (layer4_outputs[4779]) & ~(layer4_outputs[4040]);
    assign layer5_outputs[2565] = ~(layer4_outputs[174]);
    assign layer5_outputs[2566] = ~((layer4_outputs[160]) | (layer4_outputs[3030]));
    assign layer5_outputs[2567] = ~((layer4_outputs[1818]) ^ (layer4_outputs[306]));
    assign layer5_outputs[2568] = (layer4_outputs[410]) | (layer4_outputs[5118]);
    assign layer5_outputs[2569] = ~(layer4_outputs[259]);
    assign layer5_outputs[2570] = layer4_outputs[2337];
    assign layer5_outputs[2571] = ~(layer4_outputs[2306]);
    assign layer5_outputs[2572] = layer4_outputs[1331];
    assign layer5_outputs[2573] = ~(layer4_outputs[3948]);
    assign layer5_outputs[2574] = layer4_outputs[3983];
    assign layer5_outputs[2575] = ~(layer4_outputs[2071]);
    assign layer5_outputs[2576] = layer4_outputs[1874];
    assign layer5_outputs[2577] = ~((layer4_outputs[4908]) | (layer4_outputs[3373]));
    assign layer5_outputs[2578] = 1'b1;
    assign layer5_outputs[2579] = layer4_outputs[4052];
    assign layer5_outputs[2580] = ~(layer4_outputs[2996]) | (layer4_outputs[2234]);
    assign layer5_outputs[2581] = ~((layer4_outputs[982]) ^ (layer4_outputs[493]));
    assign layer5_outputs[2582] = ~((layer4_outputs[2829]) & (layer4_outputs[1701]));
    assign layer5_outputs[2583] = (layer4_outputs[1031]) & (layer4_outputs[4465]);
    assign layer5_outputs[2584] = (layer4_outputs[3686]) & ~(layer4_outputs[824]);
    assign layer5_outputs[2585] = ~((layer4_outputs[1835]) | (layer4_outputs[3375]));
    assign layer5_outputs[2586] = (layer4_outputs[2616]) ^ (layer4_outputs[1284]);
    assign layer5_outputs[2587] = ~(layer4_outputs[143]);
    assign layer5_outputs[2588] = layer4_outputs[3502];
    assign layer5_outputs[2589] = (layer4_outputs[3355]) & ~(layer4_outputs[1864]);
    assign layer5_outputs[2590] = layer4_outputs[2360];
    assign layer5_outputs[2591] = (layer4_outputs[558]) & ~(layer4_outputs[2733]);
    assign layer5_outputs[2592] = layer4_outputs[2728];
    assign layer5_outputs[2593] = layer4_outputs[975];
    assign layer5_outputs[2594] = layer4_outputs[3335];
    assign layer5_outputs[2595] = ~((layer4_outputs[2894]) | (layer4_outputs[4506]));
    assign layer5_outputs[2596] = layer4_outputs[2681];
    assign layer5_outputs[2597] = layer4_outputs[4528];
    assign layer5_outputs[2598] = ~((layer4_outputs[3399]) | (layer4_outputs[262]));
    assign layer5_outputs[2599] = ~(layer4_outputs[2742]) | (layer4_outputs[2246]);
    assign layer5_outputs[2600] = (layer4_outputs[4286]) & ~(layer4_outputs[2436]);
    assign layer5_outputs[2601] = ~(layer4_outputs[3760]);
    assign layer5_outputs[2602] = ~(layer4_outputs[3095]);
    assign layer5_outputs[2603] = ~((layer4_outputs[665]) ^ (layer4_outputs[1528]));
    assign layer5_outputs[2604] = ~(layer4_outputs[2769]);
    assign layer5_outputs[2605] = layer4_outputs[3529];
    assign layer5_outputs[2606] = layer4_outputs[3316];
    assign layer5_outputs[2607] = layer4_outputs[663];
    assign layer5_outputs[2608] = (layer4_outputs[2365]) ^ (layer4_outputs[1488]);
    assign layer5_outputs[2609] = ~((layer4_outputs[2131]) | (layer4_outputs[1905]));
    assign layer5_outputs[2610] = layer4_outputs[3986];
    assign layer5_outputs[2611] = (layer4_outputs[3263]) & ~(layer4_outputs[4276]);
    assign layer5_outputs[2612] = layer4_outputs[3865];
    assign layer5_outputs[2613] = ~(layer4_outputs[2402]);
    assign layer5_outputs[2614] = (layer4_outputs[4057]) & ~(layer4_outputs[5057]);
    assign layer5_outputs[2615] = (layer4_outputs[4924]) & (layer4_outputs[2008]);
    assign layer5_outputs[2616] = ~(layer4_outputs[3371]);
    assign layer5_outputs[2617] = layer4_outputs[2767];
    assign layer5_outputs[2618] = ~(layer4_outputs[1883]) | (layer4_outputs[2975]);
    assign layer5_outputs[2619] = (layer4_outputs[3922]) ^ (layer4_outputs[1858]);
    assign layer5_outputs[2620] = layer4_outputs[4248];
    assign layer5_outputs[2621] = (layer4_outputs[3797]) & ~(layer4_outputs[801]);
    assign layer5_outputs[2622] = ~((layer4_outputs[4448]) | (layer4_outputs[38]));
    assign layer5_outputs[2623] = layer4_outputs[4906];
    assign layer5_outputs[2624] = (layer4_outputs[647]) ^ (layer4_outputs[3478]);
    assign layer5_outputs[2625] = ~((layer4_outputs[1545]) & (layer4_outputs[1378]));
    assign layer5_outputs[2626] = layer4_outputs[851];
    assign layer5_outputs[2627] = layer4_outputs[907];
    assign layer5_outputs[2628] = (layer4_outputs[4603]) ^ (layer4_outputs[1596]);
    assign layer5_outputs[2629] = ~(layer4_outputs[2348]) | (layer4_outputs[517]);
    assign layer5_outputs[2630] = ~(layer4_outputs[2187]);
    assign layer5_outputs[2631] = ~(layer4_outputs[4092]);
    assign layer5_outputs[2632] = (layer4_outputs[26]) & ~(layer4_outputs[1754]);
    assign layer5_outputs[2633] = layer4_outputs[674];
    assign layer5_outputs[2634] = ~(layer4_outputs[4929]);
    assign layer5_outputs[2635] = ~(layer4_outputs[1849]);
    assign layer5_outputs[2636] = layer4_outputs[3296];
    assign layer5_outputs[2637] = ~((layer4_outputs[1385]) | (layer4_outputs[1024]));
    assign layer5_outputs[2638] = layer4_outputs[3362];
    assign layer5_outputs[2639] = ~(layer4_outputs[4340]);
    assign layer5_outputs[2640] = layer4_outputs[2392];
    assign layer5_outputs[2641] = (layer4_outputs[4156]) & (layer4_outputs[2454]);
    assign layer5_outputs[2642] = ~((layer4_outputs[4487]) ^ (layer4_outputs[3368]));
    assign layer5_outputs[2643] = (layer4_outputs[2979]) | (layer4_outputs[4571]);
    assign layer5_outputs[2644] = ~(layer4_outputs[5003]);
    assign layer5_outputs[2645] = ~((layer4_outputs[765]) | (layer4_outputs[687]));
    assign layer5_outputs[2646] = 1'b0;
    assign layer5_outputs[2647] = (layer4_outputs[4550]) ^ (layer4_outputs[1452]);
    assign layer5_outputs[2648] = ~(layer4_outputs[4402]);
    assign layer5_outputs[2649] = ~(layer4_outputs[4146]);
    assign layer5_outputs[2650] = (layer4_outputs[5]) ^ (layer4_outputs[3913]);
    assign layer5_outputs[2651] = layer4_outputs[1393];
    assign layer5_outputs[2652] = 1'b1;
    assign layer5_outputs[2653] = layer4_outputs[2655];
    assign layer5_outputs[2654] = layer4_outputs[5090];
    assign layer5_outputs[2655] = (layer4_outputs[206]) & ~(layer4_outputs[1877]);
    assign layer5_outputs[2656] = layer4_outputs[4578];
    assign layer5_outputs[2657] = layer4_outputs[2628];
    assign layer5_outputs[2658] = (layer4_outputs[2778]) & ~(layer4_outputs[1453]);
    assign layer5_outputs[2659] = layer4_outputs[3428];
    assign layer5_outputs[2660] = (layer4_outputs[2658]) & (layer4_outputs[2580]);
    assign layer5_outputs[2661] = ~((layer4_outputs[2652]) | (layer4_outputs[3111]));
    assign layer5_outputs[2662] = ~((layer4_outputs[1592]) & (layer4_outputs[1241]));
    assign layer5_outputs[2663] = ~(layer4_outputs[1442]);
    assign layer5_outputs[2664] = ~(layer4_outputs[1538]);
    assign layer5_outputs[2665] = ~(layer4_outputs[595]);
    assign layer5_outputs[2666] = (layer4_outputs[1694]) | (layer4_outputs[4862]);
    assign layer5_outputs[2667] = 1'b1;
    assign layer5_outputs[2668] = ~((layer4_outputs[2450]) & (layer4_outputs[3065]));
    assign layer5_outputs[2669] = (layer4_outputs[3353]) & (layer4_outputs[3649]);
    assign layer5_outputs[2670] = 1'b1;
    assign layer5_outputs[2671] = ~(layer4_outputs[4103]);
    assign layer5_outputs[2672] = ~(layer4_outputs[510]);
    assign layer5_outputs[2673] = ~(layer4_outputs[1773]);
    assign layer5_outputs[2674] = ~(layer4_outputs[119]);
    assign layer5_outputs[2675] = ~((layer4_outputs[1649]) | (layer4_outputs[4627]));
    assign layer5_outputs[2676] = ~(layer4_outputs[5015]) | (layer4_outputs[4371]);
    assign layer5_outputs[2677] = (layer4_outputs[2325]) & ~(layer4_outputs[1035]);
    assign layer5_outputs[2678] = ~(layer4_outputs[1903]) | (layer4_outputs[3624]);
    assign layer5_outputs[2679] = ~(layer4_outputs[2416]);
    assign layer5_outputs[2680] = layer4_outputs[4361];
    assign layer5_outputs[2681] = layer4_outputs[4704];
    assign layer5_outputs[2682] = ~((layer4_outputs[1422]) & (layer4_outputs[755]));
    assign layer5_outputs[2683] = ~(layer4_outputs[119]);
    assign layer5_outputs[2684] = ~(layer4_outputs[1969]);
    assign layer5_outputs[2685] = (layer4_outputs[1075]) ^ (layer4_outputs[4099]);
    assign layer5_outputs[2686] = layer4_outputs[4826];
    assign layer5_outputs[2687] = layer4_outputs[311];
    assign layer5_outputs[2688] = ~(layer4_outputs[207]);
    assign layer5_outputs[2689] = (layer4_outputs[3146]) & (layer4_outputs[637]);
    assign layer5_outputs[2690] = (layer4_outputs[1166]) & ~(layer4_outputs[831]);
    assign layer5_outputs[2691] = (layer4_outputs[2124]) & ~(layer4_outputs[3279]);
    assign layer5_outputs[2692] = ~(layer4_outputs[542]);
    assign layer5_outputs[2693] = ~(layer4_outputs[3138]);
    assign layer5_outputs[2694] = ~((layer4_outputs[263]) & (layer4_outputs[3791]));
    assign layer5_outputs[2695] = (layer4_outputs[2221]) & ~(layer4_outputs[180]);
    assign layer5_outputs[2696] = layer4_outputs[1430];
    assign layer5_outputs[2697] = ~((layer4_outputs[1738]) ^ (layer4_outputs[2297]));
    assign layer5_outputs[2698] = 1'b0;
    assign layer5_outputs[2699] = ~((layer4_outputs[516]) | (layer4_outputs[4520]));
    assign layer5_outputs[2700] = (layer4_outputs[80]) & (layer4_outputs[589]);
    assign layer5_outputs[2701] = ~((layer4_outputs[2340]) ^ (layer4_outputs[4021]));
    assign layer5_outputs[2702] = (layer4_outputs[3453]) ^ (layer4_outputs[2145]);
    assign layer5_outputs[2703] = layer4_outputs[3430];
    assign layer5_outputs[2704] = ~((layer4_outputs[1837]) ^ (layer4_outputs[419]));
    assign layer5_outputs[2705] = ~(layer4_outputs[648]);
    assign layer5_outputs[2706] = layer4_outputs[3404];
    assign layer5_outputs[2707] = ~((layer4_outputs[3752]) ^ (layer4_outputs[1989]));
    assign layer5_outputs[2708] = ~(layer4_outputs[4228]);
    assign layer5_outputs[2709] = ~(layer4_outputs[2740]);
    assign layer5_outputs[2710] = ~(layer4_outputs[825]);
    assign layer5_outputs[2711] = layer4_outputs[4418];
    assign layer5_outputs[2712] = ~(layer4_outputs[2665]) | (layer4_outputs[1848]);
    assign layer5_outputs[2713] = ~(layer4_outputs[5023]);
    assign layer5_outputs[2714] = layer4_outputs[5042];
    assign layer5_outputs[2715] = ~(layer4_outputs[4279]);
    assign layer5_outputs[2716] = ~(layer4_outputs[4064]);
    assign layer5_outputs[2717] = (layer4_outputs[4509]) & ~(layer4_outputs[1134]);
    assign layer5_outputs[2718] = (layer4_outputs[56]) & ~(layer4_outputs[4485]);
    assign layer5_outputs[2719] = ~(layer4_outputs[650]);
    assign layer5_outputs[2720] = ~(layer4_outputs[2621]) | (layer4_outputs[2449]);
    assign layer5_outputs[2721] = ~(layer4_outputs[2795]);
    assign layer5_outputs[2722] = ~(layer4_outputs[958]);
    assign layer5_outputs[2723] = ~(layer4_outputs[3744]);
    assign layer5_outputs[2724] = layer4_outputs[857];
    assign layer5_outputs[2725] = ~(layer4_outputs[3402]);
    assign layer5_outputs[2726] = layer4_outputs[894];
    assign layer5_outputs[2727] = ~(layer4_outputs[903]) | (layer4_outputs[2613]);
    assign layer5_outputs[2728] = ~(layer4_outputs[2909]);
    assign layer5_outputs[2729] = layer4_outputs[732];
    assign layer5_outputs[2730] = (layer4_outputs[2270]) | (layer4_outputs[3545]);
    assign layer5_outputs[2731] = layer4_outputs[3318];
    assign layer5_outputs[2732] = layer4_outputs[473];
    assign layer5_outputs[2733] = ~(layer4_outputs[170]);
    assign layer5_outputs[2734] = (layer4_outputs[3010]) ^ (layer4_outputs[670]);
    assign layer5_outputs[2735] = ~(layer4_outputs[2153]) | (layer4_outputs[3124]);
    assign layer5_outputs[2736] = ~(layer4_outputs[4183]) | (layer4_outputs[2330]);
    assign layer5_outputs[2737] = ~((layer4_outputs[4327]) & (layer4_outputs[1124]));
    assign layer5_outputs[2738] = ~(layer4_outputs[3425]) | (layer4_outputs[2444]);
    assign layer5_outputs[2739] = ~(layer4_outputs[5004]);
    assign layer5_outputs[2740] = ~(layer4_outputs[2420]);
    assign layer5_outputs[2741] = ~(layer4_outputs[3893]);
    assign layer5_outputs[2742] = ~(layer4_outputs[2082]);
    assign layer5_outputs[2743] = ~(layer4_outputs[735]);
    assign layer5_outputs[2744] = 1'b1;
    assign layer5_outputs[2745] = ~(layer4_outputs[446]) | (layer4_outputs[4975]);
    assign layer5_outputs[2746] = (layer4_outputs[840]) ^ (layer4_outputs[3975]);
    assign layer5_outputs[2747] = ~(layer4_outputs[1499]);
    assign layer5_outputs[2748] = ~(layer4_outputs[3636]) | (layer4_outputs[740]);
    assign layer5_outputs[2749] = (layer4_outputs[2977]) ^ (layer4_outputs[2562]);
    assign layer5_outputs[2750] = layer4_outputs[3025];
    assign layer5_outputs[2751] = (layer4_outputs[3995]) & (layer4_outputs[747]);
    assign layer5_outputs[2752] = (layer4_outputs[2147]) | (layer4_outputs[3756]);
    assign layer5_outputs[2753] = (layer4_outputs[1926]) & (layer4_outputs[2428]);
    assign layer5_outputs[2754] = layer4_outputs[4463];
    assign layer5_outputs[2755] = layer4_outputs[662];
    assign layer5_outputs[2756] = (layer4_outputs[4056]) & (layer4_outputs[2285]);
    assign layer5_outputs[2757] = layer4_outputs[2549];
    assign layer5_outputs[2758] = layer4_outputs[4646];
    assign layer5_outputs[2759] = ~(layer4_outputs[522]) | (layer4_outputs[2382]);
    assign layer5_outputs[2760] = layer4_outputs[1784];
    assign layer5_outputs[2761] = ~(layer4_outputs[3283]);
    assign layer5_outputs[2762] = ~((layer4_outputs[2297]) | (layer4_outputs[4552]));
    assign layer5_outputs[2763] = ~((layer4_outputs[1143]) ^ (layer4_outputs[4138]));
    assign layer5_outputs[2764] = ~(layer4_outputs[320]);
    assign layer5_outputs[2765] = ~(layer4_outputs[2684]) | (layer4_outputs[616]);
    assign layer5_outputs[2766] = ~(layer4_outputs[1129]);
    assign layer5_outputs[2767] = ~(layer4_outputs[893]);
    assign layer5_outputs[2768] = ~((layer4_outputs[4794]) | (layer4_outputs[4823]));
    assign layer5_outputs[2769] = (layer4_outputs[3177]) & ~(layer4_outputs[1336]);
    assign layer5_outputs[2770] = ~(layer4_outputs[607]) | (layer4_outputs[1442]);
    assign layer5_outputs[2771] = ~(layer4_outputs[3628]);
    assign layer5_outputs[2772] = ~(layer4_outputs[2120]);
    assign layer5_outputs[2773] = (layer4_outputs[4486]) & ~(layer4_outputs[1226]);
    assign layer5_outputs[2774] = layer4_outputs[1567];
    assign layer5_outputs[2775] = (layer4_outputs[3356]) | (layer4_outputs[789]);
    assign layer5_outputs[2776] = (layer4_outputs[3273]) & ~(layer4_outputs[4734]);
    assign layer5_outputs[2777] = ~((layer4_outputs[1956]) ^ (layer4_outputs[1583]));
    assign layer5_outputs[2778] = (layer4_outputs[2896]) & ~(layer4_outputs[4131]);
    assign layer5_outputs[2779] = ~((layer4_outputs[3822]) | (layer4_outputs[1244]));
    assign layer5_outputs[2780] = layer4_outputs[451];
    assign layer5_outputs[2781] = ~((layer4_outputs[225]) | (layer4_outputs[1761]));
    assign layer5_outputs[2782] = ~(layer4_outputs[3883]);
    assign layer5_outputs[2783] = ~(layer4_outputs[5039]);
    assign layer5_outputs[2784] = (layer4_outputs[3562]) & ~(layer4_outputs[4705]);
    assign layer5_outputs[2785] = ~(layer4_outputs[1086]) | (layer4_outputs[226]);
    assign layer5_outputs[2786] = ~(layer4_outputs[1240]);
    assign layer5_outputs[2787] = (layer4_outputs[3918]) & ~(layer4_outputs[2155]);
    assign layer5_outputs[2788] = layer4_outputs[1206];
    assign layer5_outputs[2789] = ~((layer4_outputs[4635]) ^ (layer4_outputs[1536]));
    assign layer5_outputs[2790] = (layer4_outputs[3171]) | (layer4_outputs[1481]);
    assign layer5_outputs[2791] = ~((layer4_outputs[382]) & (layer4_outputs[1190]));
    assign layer5_outputs[2792] = (layer4_outputs[3792]) & ~(layer4_outputs[1340]);
    assign layer5_outputs[2793] = layer4_outputs[3608];
    assign layer5_outputs[2794] = ~(layer4_outputs[2507]);
    assign layer5_outputs[2795] = ~(layer4_outputs[4594]);
    assign layer5_outputs[2796] = 1'b1;
    assign layer5_outputs[2797] = ~(layer4_outputs[1795]) | (layer4_outputs[4376]);
    assign layer5_outputs[2798] = layer4_outputs[230];
    assign layer5_outputs[2799] = ~((layer4_outputs[4408]) & (layer4_outputs[4812]));
    assign layer5_outputs[2800] = ~(layer4_outputs[961]);
    assign layer5_outputs[2801] = ~(layer4_outputs[1982]);
    assign layer5_outputs[2802] = ~(layer4_outputs[630]);
    assign layer5_outputs[2803] = (layer4_outputs[4141]) & ~(layer4_outputs[4401]);
    assign layer5_outputs[2804] = 1'b1;
    assign layer5_outputs[2805] = 1'b1;
    assign layer5_outputs[2806] = (layer4_outputs[1927]) & (layer4_outputs[3089]);
    assign layer5_outputs[2807] = (layer4_outputs[407]) ^ (layer4_outputs[3633]);
    assign layer5_outputs[2808] = ~(layer4_outputs[1370]);
    assign layer5_outputs[2809] = (layer4_outputs[4996]) & (layer4_outputs[2951]);
    assign layer5_outputs[2810] = ~((layer4_outputs[3904]) | (layer4_outputs[4557]));
    assign layer5_outputs[2811] = layer4_outputs[290];
    assign layer5_outputs[2812] = layer4_outputs[3400];
    assign layer5_outputs[2813] = layer4_outputs[380];
    assign layer5_outputs[2814] = (layer4_outputs[3071]) & ~(layer4_outputs[4076]);
    assign layer5_outputs[2815] = ~(layer4_outputs[1345]);
    assign layer5_outputs[2816] = ~((layer4_outputs[4830]) ^ (layer4_outputs[4394]));
    assign layer5_outputs[2817] = (layer4_outputs[3808]) & ~(layer4_outputs[4236]);
    assign layer5_outputs[2818] = layer4_outputs[1930];
    assign layer5_outputs[2819] = ~(layer4_outputs[1163]);
    assign layer5_outputs[2820] = 1'b1;
    assign layer5_outputs[2821] = ~(layer4_outputs[4085]);
    assign layer5_outputs[2822] = ~(layer4_outputs[2570]) | (layer4_outputs[4007]);
    assign layer5_outputs[2823] = ~((layer4_outputs[2296]) ^ (layer4_outputs[1558]));
    assign layer5_outputs[2824] = ~(layer4_outputs[1775]);
    assign layer5_outputs[2825] = ~(layer4_outputs[1794]) | (layer4_outputs[4534]);
    assign layer5_outputs[2826] = ~(layer4_outputs[2808]);
    assign layer5_outputs[2827] = ~((layer4_outputs[3305]) ^ (layer4_outputs[4191]));
    assign layer5_outputs[2828] = ~(layer4_outputs[3702]);
    assign layer5_outputs[2829] = (layer4_outputs[2383]) & ~(layer4_outputs[9]);
    assign layer5_outputs[2830] = (layer4_outputs[4909]) & ~(layer4_outputs[2875]);
    assign layer5_outputs[2831] = layer4_outputs[514];
    assign layer5_outputs[2832] = layer4_outputs[197];
    assign layer5_outputs[2833] = ~(layer4_outputs[4686]);
    assign layer5_outputs[2834] = ~((layer4_outputs[1406]) & (layer4_outputs[1998]));
    assign layer5_outputs[2835] = ~((layer4_outputs[2816]) ^ (layer4_outputs[3541]));
    assign layer5_outputs[2836] = (layer4_outputs[2322]) & ~(layer4_outputs[776]);
    assign layer5_outputs[2837] = layer4_outputs[3832];
    assign layer5_outputs[2838] = ~(layer4_outputs[1983]) | (layer4_outputs[1082]);
    assign layer5_outputs[2839] = layer4_outputs[4066];
    assign layer5_outputs[2840] = (layer4_outputs[3789]) & (layer4_outputs[1858]);
    assign layer5_outputs[2841] = ~((layer4_outputs[5114]) | (layer4_outputs[247]));
    assign layer5_outputs[2842] = layer4_outputs[3354];
    assign layer5_outputs[2843] = 1'b0;
    assign layer5_outputs[2844] = ~((layer4_outputs[4213]) | (layer4_outputs[4825]));
    assign layer5_outputs[2845] = (layer4_outputs[171]) & (layer4_outputs[1912]);
    assign layer5_outputs[2846] = (layer4_outputs[748]) & ~(layer4_outputs[3872]);
    assign layer5_outputs[2847] = 1'b1;
    assign layer5_outputs[2848] = 1'b1;
    assign layer5_outputs[2849] = layer4_outputs[4291];
    assign layer5_outputs[2850] = ~(layer4_outputs[4210]);
    assign layer5_outputs[2851] = (layer4_outputs[2621]) ^ (layer4_outputs[475]);
    assign layer5_outputs[2852] = (layer4_outputs[413]) & (layer4_outputs[3100]);
    assign layer5_outputs[2853] = ~(layer4_outputs[3889]);
    assign layer5_outputs[2854] = 1'b1;
    assign layer5_outputs[2855] = layer4_outputs[3627];
    assign layer5_outputs[2856] = layer4_outputs[1339];
    assign layer5_outputs[2857] = (layer4_outputs[2762]) & ~(layer4_outputs[1435]);
    assign layer5_outputs[2858] = ~((layer4_outputs[2963]) | (layer4_outputs[1024]));
    assign layer5_outputs[2859] = (layer4_outputs[3951]) | (layer4_outputs[2454]);
    assign layer5_outputs[2860] = ~(layer4_outputs[1121]) | (layer4_outputs[115]);
    assign layer5_outputs[2861] = ~(layer4_outputs[180]);
    assign layer5_outputs[2862] = ~(layer4_outputs[1533]);
    assign layer5_outputs[2863] = ~(layer4_outputs[2092]);
    assign layer5_outputs[2864] = ~(layer4_outputs[4315]);
    assign layer5_outputs[2865] = layer4_outputs[406];
    assign layer5_outputs[2866] = ~(layer4_outputs[86]);
    assign layer5_outputs[2867] = layer4_outputs[5075];
    assign layer5_outputs[2868] = ~((layer4_outputs[4877]) & (layer4_outputs[4011]));
    assign layer5_outputs[2869] = (layer4_outputs[4285]) & ~(layer4_outputs[1810]);
    assign layer5_outputs[2870] = ~(layer4_outputs[669]);
    assign layer5_outputs[2871] = layer4_outputs[2822];
    assign layer5_outputs[2872] = (layer4_outputs[781]) & ~(layer4_outputs[976]);
    assign layer5_outputs[2873] = ~(layer4_outputs[4017]) | (layer4_outputs[4289]);
    assign layer5_outputs[2874] = ~((layer4_outputs[4722]) | (layer4_outputs[2079]));
    assign layer5_outputs[2875] = (layer4_outputs[3262]) ^ (layer4_outputs[4255]);
    assign layer5_outputs[2876] = ~((layer4_outputs[4316]) & (layer4_outputs[852]));
    assign layer5_outputs[2877] = ~((layer4_outputs[4566]) | (layer4_outputs[3168]));
    assign layer5_outputs[2878] = ~(layer4_outputs[1579]);
    assign layer5_outputs[2879] = ~(layer4_outputs[4708]);
    assign layer5_outputs[2880] = layer4_outputs[4466];
    assign layer5_outputs[2881] = (layer4_outputs[3264]) ^ (layer4_outputs[3839]);
    assign layer5_outputs[2882] = ~((layer4_outputs[4350]) & (layer4_outputs[869]));
    assign layer5_outputs[2883] = ~(layer4_outputs[2848]) | (layer4_outputs[3110]);
    assign layer5_outputs[2884] = layer4_outputs[2883];
    assign layer5_outputs[2885] = layer4_outputs[1433];
    assign layer5_outputs[2886] = ~(layer4_outputs[2372]);
    assign layer5_outputs[2887] = ~(layer4_outputs[2848]);
    assign layer5_outputs[2888] = (layer4_outputs[3568]) & (layer4_outputs[1715]);
    assign layer5_outputs[2889] = ~((layer4_outputs[953]) ^ (layer4_outputs[1568]));
    assign layer5_outputs[2890] = layer4_outputs[4413];
    assign layer5_outputs[2891] = layer4_outputs[3235];
    assign layer5_outputs[2892] = (layer4_outputs[1213]) | (layer4_outputs[1211]);
    assign layer5_outputs[2893] = (layer4_outputs[3303]) ^ (layer4_outputs[2763]);
    assign layer5_outputs[2894] = (layer4_outputs[2892]) & (layer4_outputs[3783]);
    assign layer5_outputs[2895] = ~(layer4_outputs[5022]);
    assign layer5_outputs[2896] = 1'b1;
    assign layer5_outputs[2897] = ~(layer4_outputs[4972]);
    assign layer5_outputs[2898] = layer4_outputs[1026];
    assign layer5_outputs[2899] = layer4_outputs[108];
    assign layer5_outputs[2900] = layer4_outputs[3004];
    assign layer5_outputs[2901] = layer4_outputs[3209];
    assign layer5_outputs[2902] = (layer4_outputs[5062]) & ~(layer4_outputs[2706]);
    assign layer5_outputs[2903] = ~((layer4_outputs[1598]) & (layer4_outputs[383]));
    assign layer5_outputs[2904] = ~(layer4_outputs[1401]);
    assign layer5_outputs[2905] = (layer4_outputs[2326]) ^ (layer4_outputs[4880]);
    assign layer5_outputs[2906] = 1'b0;
    assign layer5_outputs[2907] = ~(layer4_outputs[231]);
    assign layer5_outputs[2908] = layer4_outputs[4012];
    assign layer5_outputs[2909] = (layer4_outputs[3180]) | (layer4_outputs[985]);
    assign layer5_outputs[2910] = layer4_outputs[4149];
    assign layer5_outputs[2911] = ~(layer4_outputs[109]);
    assign layer5_outputs[2912] = ~((layer4_outputs[4271]) ^ (layer4_outputs[4303]));
    assign layer5_outputs[2913] = ~(layer4_outputs[5073]);
    assign layer5_outputs[2914] = ~(layer4_outputs[4999]);
    assign layer5_outputs[2915] = (layer4_outputs[796]) & ~(layer4_outputs[4940]);
    assign layer5_outputs[2916] = ~(layer4_outputs[3180]);
    assign layer5_outputs[2917] = ~((layer4_outputs[5089]) ^ (layer4_outputs[865]));
    assign layer5_outputs[2918] = ~(layer4_outputs[894]);
    assign layer5_outputs[2919] = (layer4_outputs[2957]) & (layer4_outputs[2733]);
    assign layer5_outputs[2920] = ~(layer4_outputs[2294]);
    assign layer5_outputs[2921] = 1'b1;
    assign layer5_outputs[2922] = layer4_outputs[1021];
    assign layer5_outputs[2923] = layer4_outputs[3506];
    assign layer5_outputs[2924] = ~(layer4_outputs[2681]) | (layer4_outputs[4786]);
    assign layer5_outputs[2925] = ~(layer4_outputs[4781]);
    assign layer5_outputs[2926] = ~((layer4_outputs[1283]) | (layer4_outputs[4035]));
    assign layer5_outputs[2927] = (layer4_outputs[4170]) | (layer4_outputs[2500]);
    assign layer5_outputs[2928] = layer4_outputs[3451];
    assign layer5_outputs[2929] = ~(layer4_outputs[2888]);
    assign layer5_outputs[2930] = layer4_outputs[1554];
    assign layer5_outputs[2931] = layer4_outputs[1722];
    assign layer5_outputs[2932] = layer4_outputs[2704];
    assign layer5_outputs[2933] = ~(layer4_outputs[2581]) | (layer4_outputs[153]);
    assign layer5_outputs[2934] = ~(layer4_outputs[164]);
    assign layer5_outputs[2935] = layer4_outputs[4705];
    assign layer5_outputs[2936] = (layer4_outputs[2215]) & ~(layer4_outputs[4932]);
    assign layer5_outputs[2937] = layer4_outputs[1764];
    assign layer5_outputs[2938] = layer4_outputs[1763];
    assign layer5_outputs[2939] = layer4_outputs[323];
    assign layer5_outputs[2940] = layer4_outputs[1014];
    assign layer5_outputs[2941] = (layer4_outputs[2476]) & (layer4_outputs[1281]);
    assign layer5_outputs[2942] = layer4_outputs[4485];
    assign layer5_outputs[2943] = ~((layer4_outputs[2047]) ^ (layer4_outputs[2141]));
    assign layer5_outputs[2944] = (layer4_outputs[3401]) & (layer4_outputs[245]);
    assign layer5_outputs[2945] = ~(layer4_outputs[1181]);
    assign layer5_outputs[2946] = ~(layer4_outputs[2770]);
    assign layer5_outputs[2947] = layer4_outputs[4397];
    assign layer5_outputs[2948] = (layer4_outputs[398]) & (layer4_outputs[7]);
    assign layer5_outputs[2949] = layer4_outputs[2265];
    assign layer5_outputs[2950] = layer4_outputs[1673];
    assign layer5_outputs[2951] = ~(layer4_outputs[2104]);
    assign layer5_outputs[2952] = layer4_outputs[3297];
    assign layer5_outputs[2953] = ~(layer4_outputs[2110]);
    assign layer5_outputs[2954] = ~((layer4_outputs[1271]) | (layer4_outputs[350]));
    assign layer5_outputs[2955] = ~(layer4_outputs[722]);
    assign layer5_outputs[2956] = ~(layer4_outputs[784]) | (layer4_outputs[3716]);
    assign layer5_outputs[2957] = ~((layer4_outputs[2760]) ^ (layer4_outputs[3838]));
    assign layer5_outputs[2958] = ~(layer4_outputs[1207]);
    assign layer5_outputs[2959] = ~(layer4_outputs[4269]);
    assign layer5_outputs[2960] = (layer4_outputs[2324]) & ~(layer4_outputs[759]);
    assign layer5_outputs[2961] = ~(layer4_outputs[1105]);
    assign layer5_outputs[2962] = ~(layer4_outputs[2422]);
    assign layer5_outputs[2963] = ~((layer4_outputs[2487]) | (layer4_outputs[5096]));
    assign layer5_outputs[2964] = (layer4_outputs[3023]) & ~(layer4_outputs[4264]);
    assign layer5_outputs[2965] = layer4_outputs[4823];
    assign layer5_outputs[2966] = (layer4_outputs[2031]) & (layer4_outputs[2890]);
    assign layer5_outputs[2967] = layer4_outputs[899];
    assign layer5_outputs[2968] = (layer4_outputs[1237]) & (layer4_outputs[2137]);
    assign layer5_outputs[2969] = (layer4_outputs[4000]) & (layer4_outputs[516]);
    assign layer5_outputs[2970] = ~(layer4_outputs[3162]);
    assign layer5_outputs[2971] = ~((layer4_outputs[1170]) & (layer4_outputs[3055]));
    assign layer5_outputs[2972] = (layer4_outputs[181]) & (layer4_outputs[1168]);
    assign layer5_outputs[2973] = layer4_outputs[4105];
    assign layer5_outputs[2974] = layer4_outputs[1729];
    assign layer5_outputs[2975] = (layer4_outputs[3119]) & ~(layer4_outputs[1615]);
    assign layer5_outputs[2976] = ~(layer4_outputs[4673]);
    assign layer5_outputs[2977] = ~(layer4_outputs[1893]) | (layer4_outputs[3654]);
    assign layer5_outputs[2978] = 1'b1;
    assign layer5_outputs[2979] = layer4_outputs[1913];
    assign layer5_outputs[2980] = ~(layer4_outputs[2134]);
    assign layer5_outputs[2981] = ~(layer4_outputs[5113]);
    assign layer5_outputs[2982] = (layer4_outputs[1728]) & ~(layer4_outputs[2364]);
    assign layer5_outputs[2983] = (layer4_outputs[1745]) & ~(layer4_outputs[4372]);
    assign layer5_outputs[2984] = (layer4_outputs[2561]) | (layer4_outputs[1367]);
    assign layer5_outputs[2985] = (layer4_outputs[3038]) & (layer4_outputs[1928]);
    assign layer5_outputs[2986] = layer4_outputs[1756];
    assign layer5_outputs[2987] = ~((layer4_outputs[2381]) & (layer4_outputs[1067]));
    assign layer5_outputs[2988] = ~(layer4_outputs[1950]);
    assign layer5_outputs[2989] = (layer4_outputs[1569]) | (layer4_outputs[2578]);
    assign layer5_outputs[2990] = (layer4_outputs[3471]) | (layer4_outputs[2572]);
    assign layer5_outputs[2991] = ~(layer4_outputs[4287]);
    assign layer5_outputs[2992] = 1'b1;
    assign layer5_outputs[2993] = (layer4_outputs[3211]) & ~(layer4_outputs[2196]);
    assign layer5_outputs[2994] = ~((layer4_outputs[3445]) | (layer4_outputs[4889]));
    assign layer5_outputs[2995] = (layer4_outputs[2546]) & (layer4_outputs[3492]);
    assign layer5_outputs[2996] = ~(layer4_outputs[2873]) | (layer4_outputs[4651]);
    assign layer5_outputs[2997] = 1'b1;
    assign layer5_outputs[2998] = ~(layer4_outputs[852]);
    assign layer5_outputs[2999] = (layer4_outputs[3892]) ^ (layer4_outputs[2177]);
    assign layer5_outputs[3000] = (layer4_outputs[3777]) & ~(layer4_outputs[771]);
    assign layer5_outputs[3001] = (layer4_outputs[969]) | (layer4_outputs[1591]);
    assign layer5_outputs[3002] = ~((layer4_outputs[3001]) | (layer4_outputs[318]));
    assign layer5_outputs[3003] = layer4_outputs[355];
    assign layer5_outputs[3004] = ~(layer4_outputs[2549]);
    assign layer5_outputs[3005] = ~(layer4_outputs[4822]);
    assign layer5_outputs[3006] = layer4_outputs[1994];
    assign layer5_outputs[3007] = 1'b0;
    assign layer5_outputs[3008] = ~(layer4_outputs[2587]);
    assign layer5_outputs[3009] = (layer4_outputs[3665]) | (layer4_outputs[1469]);
    assign layer5_outputs[3010] = layer4_outputs[4782];
    assign layer5_outputs[3011] = (layer4_outputs[4334]) & ~(layer4_outputs[1637]);
    assign layer5_outputs[3012] = layer4_outputs[113];
    assign layer5_outputs[3013] = ~(layer4_outputs[1348]);
    assign layer5_outputs[3014] = ~(layer4_outputs[4908]);
    assign layer5_outputs[3015] = layer4_outputs[597];
    assign layer5_outputs[3016] = ~(layer4_outputs[1547]);
    assign layer5_outputs[3017] = ~((layer4_outputs[4497]) & (layer4_outputs[4356]));
    assign layer5_outputs[3018] = 1'b0;
    assign layer5_outputs[3019] = (layer4_outputs[2862]) | (layer4_outputs[515]);
    assign layer5_outputs[3020] = layer4_outputs[73];
    assign layer5_outputs[3021] = layer4_outputs[750];
    assign layer5_outputs[3022] = ~(layer4_outputs[4129]);
    assign layer5_outputs[3023] = (layer4_outputs[539]) ^ (layer4_outputs[4286]);
    assign layer5_outputs[3024] = ~(layer4_outputs[4047]);
    assign layer5_outputs[3025] = ~(layer4_outputs[2995]);
    assign layer5_outputs[3026] = ~(layer4_outputs[1400]);
    assign layer5_outputs[3027] = 1'b1;
    assign layer5_outputs[3028] = (layer4_outputs[1878]) & ~(layer4_outputs[4600]);
    assign layer5_outputs[3029] = ~(layer4_outputs[3043]);
    assign layer5_outputs[3030] = layer4_outputs[336];
    assign layer5_outputs[3031] = ~((layer4_outputs[2943]) | (layer4_outputs[3339]));
    assign layer5_outputs[3032] = layer4_outputs[3921];
    assign layer5_outputs[3033] = (layer4_outputs[459]) ^ (layer4_outputs[5084]);
    assign layer5_outputs[3034] = (layer4_outputs[1225]) & ~(layer4_outputs[969]);
    assign layer5_outputs[3035] = 1'b1;
    assign layer5_outputs[3036] = layer4_outputs[1152];
    assign layer5_outputs[3037] = layer4_outputs[2314];
    assign layer5_outputs[3038] = 1'b0;
    assign layer5_outputs[3039] = (layer4_outputs[917]) & (layer4_outputs[2607]);
    assign layer5_outputs[3040] = layer4_outputs[4189];
    assign layer5_outputs[3041] = layer4_outputs[480];
    assign layer5_outputs[3042] = ~(layer4_outputs[3502]);
    assign layer5_outputs[3043] = layer4_outputs[2507];
    assign layer5_outputs[3044] = ~(layer4_outputs[4679]) | (layer4_outputs[210]);
    assign layer5_outputs[3045] = layer4_outputs[1765];
    assign layer5_outputs[3046] = ~(layer4_outputs[2142]) | (layer4_outputs[4219]);
    assign layer5_outputs[3047] = 1'b0;
    assign layer5_outputs[3048] = (layer4_outputs[4725]) & (layer4_outputs[3650]);
    assign layer5_outputs[3049] = (layer4_outputs[1556]) & (layer4_outputs[941]);
    assign layer5_outputs[3050] = ~((layer4_outputs[935]) & (layer4_outputs[4011]));
    assign layer5_outputs[3051] = layer4_outputs[4972];
    assign layer5_outputs[3052] = (layer4_outputs[3605]) & (layer4_outputs[228]);
    assign layer5_outputs[3053] = ~(layer4_outputs[1374]) | (layer4_outputs[2697]);
    assign layer5_outputs[3054] = ~(layer4_outputs[2835]);
    assign layer5_outputs[3055] = (layer4_outputs[422]) & ~(layer4_outputs[741]);
    assign layer5_outputs[3056] = ~(layer4_outputs[1660]) | (layer4_outputs[3573]);
    assign layer5_outputs[3057] = ~(layer4_outputs[4683]);
    assign layer5_outputs[3058] = ~(layer4_outputs[3013]) | (layer4_outputs[2200]);
    assign layer5_outputs[3059] = layer4_outputs[1748];
    assign layer5_outputs[3060] = layer4_outputs[2212];
    assign layer5_outputs[3061] = layer4_outputs[322];
    assign layer5_outputs[3062] = layer4_outputs[4114];
    assign layer5_outputs[3063] = ~(layer4_outputs[3743]);
    assign layer5_outputs[3064] = 1'b1;
    assign layer5_outputs[3065] = 1'b1;
    assign layer5_outputs[3066] = (layer4_outputs[1616]) ^ (layer4_outputs[387]);
    assign layer5_outputs[3067] = ~(layer4_outputs[938]);
    assign layer5_outputs[3068] = ~(layer4_outputs[1059]);
    assign layer5_outputs[3069] = 1'b1;
    assign layer5_outputs[3070] = ~((layer4_outputs[2761]) ^ (layer4_outputs[4008]));
    assign layer5_outputs[3071] = layer4_outputs[3986];
    assign layer5_outputs[3072] = ~(layer4_outputs[4595]);
    assign layer5_outputs[3073] = (layer4_outputs[4277]) | (layer4_outputs[4672]);
    assign layer5_outputs[3074] = ~((layer4_outputs[4471]) | (layer4_outputs[2234]));
    assign layer5_outputs[3075] = ~(layer4_outputs[2194]);
    assign layer5_outputs[3076] = ~((layer4_outputs[3862]) ^ (layer4_outputs[4195]));
    assign layer5_outputs[3077] = layer4_outputs[4184];
    assign layer5_outputs[3078] = ~(layer4_outputs[41]);
    assign layer5_outputs[3079] = ~(layer4_outputs[971]) | (layer4_outputs[2718]);
    assign layer5_outputs[3080] = ~(layer4_outputs[791]) | (layer4_outputs[3917]);
    assign layer5_outputs[3081] = ~((layer4_outputs[4267]) | (layer4_outputs[3450]));
    assign layer5_outputs[3082] = (layer4_outputs[1555]) & (layer4_outputs[3570]);
    assign layer5_outputs[3083] = 1'b0;
    assign layer5_outputs[3084] = layer4_outputs[4400];
    assign layer5_outputs[3085] = ~(layer4_outputs[635]) | (layer4_outputs[4069]);
    assign layer5_outputs[3086] = (layer4_outputs[4135]) ^ (layer4_outputs[3709]);
    assign layer5_outputs[3087] = layer4_outputs[880];
    assign layer5_outputs[3088] = layer4_outputs[3122];
    assign layer5_outputs[3089] = ~((layer4_outputs[279]) ^ (layer4_outputs[203]));
    assign layer5_outputs[3090] = ~(layer4_outputs[3891]);
    assign layer5_outputs[3091] = (layer4_outputs[4408]) | (layer4_outputs[1312]);
    assign layer5_outputs[3092] = (layer4_outputs[3604]) & ~(layer4_outputs[2373]);
    assign layer5_outputs[3093] = (layer4_outputs[2636]) & ~(layer4_outputs[243]);
    assign layer5_outputs[3094] = 1'b1;
    assign layer5_outputs[3095] = layer4_outputs[3106];
    assign layer5_outputs[3096] = ~(layer4_outputs[1098]);
    assign layer5_outputs[3097] = layer4_outputs[4660];
    assign layer5_outputs[3098] = (layer4_outputs[2856]) | (layer4_outputs[2240]);
    assign layer5_outputs[3099] = (layer4_outputs[496]) & ~(layer4_outputs[4123]);
    assign layer5_outputs[3100] = ~((layer4_outputs[4278]) ^ (layer4_outputs[4364]));
    assign layer5_outputs[3101] = ~(layer4_outputs[2994]);
    assign layer5_outputs[3102] = ~(layer4_outputs[3488]);
    assign layer5_outputs[3103] = ~(layer4_outputs[2113]);
    assign layer5_outputs[3104] = layer4_outputs[430];
    assign layer5_outputs[3105] = (layer4_outputs[2949]) & ~(layer4_outputs[1372]);
    assign layer5_outputs[3106] = ~((layer4_outputs[538]) | (layer4_outputs[368]));
    assign layer5_outputs[3107] = (layer4_outputs[4624]) & (layer4_outputs[1431]);
    assign layer5_outputs[3108] = ~(layer4_outputs[1657]);
    assign layer5_outputs[3109] = layer4_outputs[3069];
    assign layer5_outputs[3110] = ~(layer4_outputs[4934]);
    assign layer5_outputs[3111] = layer4_outputs[3703];
    assign layer5_outputs[3112] = ~((layer4_outputs[282]) ^ (layer4_outputs[1028]));
    assign layer5_outputs[3113] = 1'b1;
    assign layer5_outputs[3114] = layer4_outputs[2369];
    assign layer5_outputs[3115] = layer4_outputs[660];
    assign layer5_outputs[3116] = ~(layer4_outputs[4851]) | (layer4_outputs[2818]);
    assign layer5_outputs[3117] = ~(layer4_outputs[1385]);
    assign layer5_outputs[3118] = ~((layer4_outputs[3116]) ^ (layer4_outputs[4688]));
    assign layer5_outputs[3119] = layer4_outputs[1720];
    assign layer5_outputs[3120] = ~(layer4_outputs[2433]) | (layer4_outputs[39]);
    assign layer5_outputs[3121] = ~(layer4_outputs[1369]) | (layer4_outputs[3537]);
    assign layer5_outputs[3122] = layer4_outputs[2253];
    assign layer5_outputs[3123] = (layer4_outputs[3926]) & ~(layer4_outputs[2046]);
    assign layer5_outputs[3124] = (layer4_outputs[2923]) & ~(layer4_outputs[3984]);
    assign layer5_outputs[3125] = ~((layer4_outputs[3725]) ^ (layer4_outputs[3982]));
    assign layer5_outputs[3126] = layer4_outputs[592];
    assign layer5_outputs[3127] = 1'b1;
    assign layer5_outputs[3128] = (layer4_outputs[5065]) & ~(layer4_outputs[1290]);
    assign layer5_outputs[3129] = ~(layer4_outputs[4710]) | (layer4_outputs[4236]);
    assign layer5_outputs[3130] = ~(layer4_outputs[752]);
    assign layer5_outputs[3131] = (layer4_outputs[4239]) & ~(layer4_outputs[4483]);
    assign layer5_outputs[3132] = (layer4_outputs[1584]) & (layer4_outputs[2365]);
    assign layer5_outputs[3133] = ~(layer4_outputs[2574]);
    assign layer5_outputs[3134] = layer4_outputs[4885];
    assign layer5_outputs[3135] = 1'b0;
    assign layer5_outputs[3136] = ~(layer4_outputs[1684]) | (layer4_outputs[3684]);
    assign layer5_outputs[3137] = ~(layer4_outputs[53]);
    assign layer5_outputs[3138] = ~((layer4_outputs[1113]) ^ (layer4_outputs[3381]));
    assign layer5_outputs[3139] = ~(layer4_outputs[158]) | (layer4_outputs[719]);
    assign layer5_outputs[3140] = ~(layer4_outputs[1436]);
    assign layer5_outputs[3141] = ~(layer4_outputs[2802]);
    assign layer5_outputs[3142] = ~(layer4_outputs[701]);
    assign layer5_outputs[3143] = ~((layer4_outputs[4018]) & (layer4_outputs[254]));
    assign layer5_outputs[3144] = layer4_outputs[1250];
    assign layer5_outputs[3145] = (layer4_outputs[4042]) & ~(layer4_outputs[834]);
    assign layer5_outputs[3146] = (layer4_outputs[2884]) ^ (layer4_outputs[3804]);
    assign layer5_outputs[3147] = layer4_outputs[4326];
    assign layer5_outputs[3148] = ~(layer4_outputs[4273]) | (layer4_outputs[3936]);
    assign layer5_outputs[3149] = ~(layer4_outputs[2704]) | (layer4_outputs[2754]);
    assign layer5_outputs[3150] = ~((layer4_outputs[1297]) ^ (layer4_outputs[4268]));
    assign layer5_outputs[3151] = ~((layer4_outputs[2900]) & (layer4_outputs[3715]));
    assign layer5_outputs[3152] = (layer4_outputs[3550]) ^ (layer4_outputs[4811]);
    assign layer5_outputs[3153] = (layer4_outputs[4341]) ^ (layer4_outputs[1073]);
    assign layer5_outputs[3154] = layer4_outputs[1524];
    assign layer5_outputs[3155] = layer4_outputs[5001];
    assign layer5_outputs[3156] = 1'b0;
    assign layer5_outputs[3157] = ~(layer4_outputs[3619]);
    assign layer5_outputs[3158] = layer4_outputs[3274];
    assign layer5_outputs[3159] = layer4_outputs[3333];
    assign layer5_outputs[3160] = ~(layer4_outputs[3205]) | (layer4_outputs[285]);
    assign layer5_outputs[3161] = layer4_outputs[70];
    assign layer5_outputs[3162] = (layer4_outputs[2929]) & (layer4_outputs[1096]);
    assign layer5_outputs[3163] = ~((layer4_outputs[1724]) & (layer4_outputs[4994]));
    assign layer5_outputs[3164] = ~((layer4_outputs[1600]) ^ (layer4_outputs[3509]));
    assign layer5_outputs[3165] = layer4_outputs[4914];
    assign layer5_outputs[3166] = layer4_outputs[1356];
    assign layer5_outputs[3167] = ~((layer4_outputs[4522]) & (layer4_outputs[4423]));
    assign layer5_outputs[3168] = (layer4_outputs[1580]) & (layer4_outputs[3894]);
    assign layer5_outputs[3169] = ~((layer4_outputs[2823]) & (layer4_outputs[4400]));
    assign layer5_outputs[3170] = ~((layer4_outputs[1907]) & (layer4_outputs[2542]));
    assign layer5_outputs[3171] = ~((layer4_outputs[4499]) & (layer4_outputs[806]));
    assign layer5_outputs[3172] = layer4_outputs[3590];
    assign layer5_outputs[3173] = ~(layer4_outputs[1797]) | (layer4_outputs[2114]);
    assign layer5_outputs[3174] = layer4_outputs[569];
    assign layer5_outputs[3175] = ~(layer4_outputs[782]);
    assign layer5_outputs[3176] = 1'b0;
    assign layer5_outputs[3177] = layer4_outputs[1118];
    assign layer5_outputs[3178] = ~(layer4_outputs[1475]);
    assign layer5_outputs[3179] = layer4_outputs[710];
    assign layer5_outputs[3180] = ~((layer4_outputs[3648]) | (layer4_outputs[4450]));
    assign layer5_outputs[3181] = layer4_outputs[3552];
    assign layer5_outputs[3182] = ~((layer4_outputs[4893]) ^ (layer4_outputs[552]));
    assign layer5_outputs[3183] = layer4_outputs[563];
    assign layer5_outputs[3184] = ~(layer4_outputs[594]);
    assign layer5_outputs[3185] = layer4_outputs[2077];
    assign layer5_outputs[3186] = ~(layer4_outputs[2225]);
    assign layer5_outputs[3187] = (layer4_outputs[937]) ^ (layer4_outputs[5029]);
    assign layer5_outputs[3188] = layer4_outputs[307];
    assign layer5_outputs[3189] = (layer4_outputs[5052]) ^ (layer4_outputs[2689]);
    assign layer5_outputs[3190] = ~(layer4_outputs[3491]) | (layer4_outputs[3723]);
    assign layer5_outputs[3191] = (layer4_outputs[3857]) & ~(layer4_outputs[126]);
    assign layer5_outputs[3192] = ~((layer4_outputs[4748]) | (layer4_outputs[234]));
    assign layer5_outputs[3193] = layer4_outputs[1652];
    assign layer5_outputs[3194] = (layer4_outputs[2746]) ^ (layer4_outputs[635]);
    assign layer5_outputs[3195] = (layer4_outputs[532]) ^ (layer4_outputs[1282]);
    assign layer5_outputs[3196] = layer4_outputs[1200];
    assign layer5_outputs[3197] = ~(layer4_outputs[4078]);
    assign layer5_outputs[3198] = ~(layer4_outputs[3155]);
    assign layer5_outputs[3199] = ~((layer4_outputs[5087]) ^ (layer4_outputs[3579]));
    assign layer5_outputs[3200] = ~(layer4_outputs[993]);
    assign layer5_outputs[3201] = (layer4_outputs[4369]) | (layer4_outputs[1163]);
    assign layer5_outputs[3202] = ~((layer4_outputs[832]) & (layer4_outputs[1532]));
    assign layer5_outputs[3203] = (layer4_outputs[2348]) & ~(layer4_outputs[2366]);
    assign layer5_outputs[3204] = (layer4_outputs[3989]) & (layer4_outputs[3359]);
    assign layer5_outputs[3205] = ~(layer4_outputs[743]) | (layer4_outputs[5075]);
    assign layer5_outputs[3206] = ~(layer4_outputs[3048]) | (layer4_outputs[3888]);
    assign layer5_outputs[3207] = (layer4_outputs[4740]) & ~(layer4_outputs[6]);
    assign layer5_outputs[3208] = ~(layer4_outputs[4679]) | (layer4_outputs[3057]);
    assign layer5_outputs[3209] = (layer4_outputs[128]) ^ (layer4_outputs[3745]);
    assign layer5_outputs[3210] = ~((layer4_outputs[955]) ^ (layer4_outputs[351]));
    assign layer5_outputs[3211] = (layer4_outputs[2931]) ^ (layer4_outputs[2386]);
    assign layer5_outputs[3212] = ~((layer4_outputs[1932]) ^ (layer4_outputs[2812]));
    assign layer5_outputs[3213] = (layer4_outputs[2410]) & (layer4_outputs[1228]);
    assign layer5_outputs[3214] = (layer4_outputs[4410]) & (layer4_outputs[2885]);
    assign layer5_outputs[3215] = ~(layer4_outputs[1914]);
    assign layer5_outputs[3216] = ~((layer4_outputs[2328]) & (layer4_outputs[1703]));
    assign layer5_outputs[3217] = (layer4_outputs[4488]) | (layer4_outputs[2817]);
    assign layer5_outputs[3218] = layer4_outputs[1478];
    assign layer5_outputs[3219] = ~(layer4_outputs[3598]);
    assign layer5_outputs[3220] = ~(layer4_outputs[138]);
    assign layer5_outputs[3221] = (layer4_outputs[2406]) | (layer4_outputs[2665]);
    assign layer5_outputs[3222] = layer4_outputs[870];
    assign layer5_outputs[3223] = ~(layer4_outputs[3635]) | (layer4_outputs[2857]);
    assign layer5_outputs[3224] = ~(layer4_outputs[3591]);
    assign layer5_outputs[3225] = layer4_outputs[1613];
    assign layer5_outputs[3226] = (layer4_outputs[3112]) & ~(layer4_outputs[1367]);
    assign layer5_outputs[3227] = layer4_outputs[307];
    assign layer5_outputs[3228] = ~((layer4_outputs[4794]) ^ (layer4_outputs[2270]));
    assign layer5_outputs[3229] = layer4_outputs[981];
    assign layer5_outputs[3230] = layer4_outputs[2321];
    assign layer5_outputs[3231] = layer4_outputs[692];
    assign layer5_outputs[3232] = layer4_outputs[4419];
    assign layer5_outputs[3233] = layer4_outputs[1865];
    assign layer5_outputs[3234] = (layer4_outputs[4919]) & ~(layer4_outputs[2071]);
    assign layer5_outputs[3235] = (layer4_outputs[1627]) | (layer4_outputs[4395]);
    assign layer5_outputs[3236] = layer4_outputs[5086];
    assign layer5_outputs[3237] = ~(layer4_outputs[486]);
    assign layer5_outputs[3238] = 1'b0;
    assign layer5_outputs[3239] = layer4_outputs[3984];
    assign layer5_outputs[3240] = ~(layer4_outputs[3585]);
    assign layer5_outputs[3241] = ~(layer4_outputs[3046]) | (layer4_outputs[329]);
    assign layer5_outputs[3242] = ~((layer4_outputs[3579]) ^ (layer4_outputs[2626]));
    assign layer5_outputs[3243] = ~(layer4_outputs[1059]);
    assign layer5_outputs[3244] = layer4_outputs[3295];
    assign layer5_outputs[3245] = layer4_outputs[2448];
    assign layer5_outputs[3246] = ~(layer4_outputs[3646]);
    assign layer5_outputs[3247] = ~(layer4_outputs[245]);
    assign layer5_outputs[3248] = ~((layer4_outputs[98]) & (layer4_outputs[2957]));
    assign layer5_outputs[3249] = ~(layer4_outputs[1721]) | (layer4_outputs[3644]);
    assign layer5_outputs[3250] = ~(layer4_outputs[3071]);
    assign layer5_outputs[3251] = ~(layer4_outputs[1628]);
    assign layer5_outputs[3252] = (layer4_outputs[4689]) & ~(layer4_outputs[2224]);
    assign layer5_outputs[3253] = ~(layer4_outputs[2042]);
    assign layer5_outputs[3254] = layer4_outputs[4719];
    assign layer5_outputs[3255] = (layer4_outputs[3895]) & ~(layer4_outputs[878]);
    assign layer5_outputs[3256] = (layer4_outputs[2103]) ^ (layer4_outputs[421]);
    assign layer5_outputs[3257] = (layer4_outputs[99]) & ~(layer4_outputs[3074]);
    assign layer5_outputs[3258] = layer4_outputs[1487];
    assign layer5_outputs[3259] = ~(layer4_outputs[5000]);
    assign layer5_outputs[3260] = ~(layer4_outputs[4365]);
    assign layer5_outputs[3261] = ~(layer4_outputs[4379]);
    assign layer5_outputs[3262] = ~((layer4_outputs[2892]) & (layer4_outputs[1010]));
    assign layer5_outputs[3263] = layer4_outputs[1820];
    assign layer5_outputs[3264] = (layer4_outputs[3348]) & (layer4_outputs[4433]);
    assign layer5_outputs[3265] = ~(layer4_outputs[1965]);
    assign layer5_outputs[3266] = ~((layer4_outputs[4169]) | (layer4_outputs[4886]));
    assign layer5_outputs[3267] = ~(layer4_outputs[2644]);
    assign layer5_outputs[3268] = layer4_outputs[2472];
    assign layer5_outputs[3269] = ~(layer4_outputs[3853]);
    assign layer5_outputs[3270] = 1'b0;
    assign layer5_outputs[3271] = ~(layer4_outputs[5012]);
    assign layer5_outputs[3272] = (layer4_outputs[3817]) | (layer4_outputs[2230]);
    assign layer5_outputs[3273] = (layer4_outputs[4598]) & ~(layer4_outputs[876]);
    assign layer5_outputs[3274] = layer4_outputs[2799];
    assign layer5_outputs[3275] = layer4_outputs[895];
    assign layer5_outputs[3276] = (layer4_outputs[3089]) & ~(layer4_outputs[4827]);
    assign layer5_outputs[3277] = (layer4_outputs[3736]) & ~(layer4_outputs[4750]);
    assign layer5_outputs[3278] = 1'b0;
    assign layer5_outputs[3279] = layer4_outputs[4154];
    assign layer5_outputs[3280] = ~((layer4_outputs[4837]) & (layer4_outputs[1110]));
    assign layer5_outputs[3281] = layer4_outputs[2243];
    assign layer5_outputs[3282] = ~(layer4_outputs[4556]) | (layer4_outputs[2729]);
    assign layer5_outputs[3283] = (layer4_outputs[2602]) & ~(layer4_outputs[4259]);
    assign layer5_outputs[3284] = ~(layer4_outputs[4328]);
    assign layer5_outputs[3285] = ~((layer4_outputs[3118]) | (layer4_outputs[4149]));
    assign layer5_outputs[3286] = layer4_outputs[4660];
    assign layer5_outputs[3287] = (layer4_outputs[4095]) & ~(layer4_outputs[2899]);
    assign layer5_outputs[3288] = layer4_outputs[4820];
    assign layer5_outputs[3289] = ~(layer4_outputs[1249]);
    assign layer5_outputs[3290] = (layer4_outputs[2940]) ^ (layer4_outputs[4407]);
    assign layer5_outputs[3291] = (layer4_outputs[62]) & (layer4_outputs[947]);
    assign layer5_outputs[3292] = layer4_outputs[2846];
    assign layer5_outputs[3293] = (layer4_outputs[4322]) & (layer4_outputs[5073]);
    assign layer5_outputs[3294] = layer4_outputs[2011];
    assign layer5_outputs[3295] = ~(layer4_outputs[3337]);
    assign layer5_outputs[3296] = (layer4_outputs[4297]) ^ (layer4_outputs[4044]);
    assign layer5_outputs[3297] = ~(layer4_outputs[4991]) | (layer4_outputs[4027]);
    assign layer5_outputs[3298] = (layer4_outputs[2700]) | (layer4_outputs[3049]);
    assign layer5_outputs[3299] = (layer4_outputs[4773]) & ~(layer4_outputs[4862]);
    assign layer5_outputs[3300] = ~(layer4_outputs[2051]);
    assign layer5_outputs[3301] = ~(layer4_outputs[2719]);
    assign layer5_outputs[3302] = layer4_outputs[2573];
    assign layer5_outputs[3303] = 1'b0;
    assign layer5_outputs[3304] = ~(layer4_outputs[2022]);
    assign layer5_outputs[3305] = (layer4_outputs[3391]) & (layer4_outputs[489]);
    assign layer5_outputs[3306] = layer4_outputs[1461];
    assign layer5_outputs[3307] = ~((layer4_outputs[1774]) ^ (layer4_outputs[2191]));
    assign layer5_outputs[3308] = (layer4_outputs[4321]) & ~(layer4_outputs[2864]);
    assign layer5_outputs[3309] = ~(layer4_outputs[1599]);
    assign layer5_outputs[3310] = ~(layer4_outputs[1822]) | (layer4_outputs[2486]);
    assign layer5_outputs[3311] = (layer4_outputs[4839]) & (layer4_outputs[1042]);
    assign layer5_outputs[3312] = ~(layer4_outputs[4147]) | (layer4_outputs[3817]);
    assign layer5_outputs[3313] = ~(layer4_outputs[2333]);
    assign layer5_outputs[3314] = layer4_outputs[2985];
    assign layer5_outputs[3315] = ~((layer4_outputs[149]) & (layer4_outputs[4045]));
    assign layer5_outputs[3316] = layer4_outputs[3694];
    assign layer5_outputs[3317] = ~(layer4_outputs[2336]);
    assign layer5_outputs[3318] = layer4_outputs[2766];
    assign layer5_outputs[3319] = layer4_outputs[4657];
    assign layer5_outputs[3320] = ~(layer4_outputs[3708]) | (layer4_outputs[1454]);
    assign layer5_outputs[3321] = (layer4_outputs[1052]) & ~(layer4_outputs[2952]);
    assign layer5_outputs[3322] = layer4_outputs[3301];
    assign layer5_outputs[3323] = layer4_outputs[2452];
    assign layer5_outputs[3324] = layer4_outputs[1897];
    assign layer5_outputs[3325] = layer4_outputs[5001];
    assign layer5_outputs[3326] = 1'b0;
    assign layer5_outputs[3327] = ~(layer4_outputs[972]);
    assign layer5_outputs[3328] = ~(layer4_outputs[4428]);
    assign layer5_outputs[3329] = layer4_outputs[2056];
    assign layer5_outputs[3330] = layer4_outputs[1806];
    assign layer5_outputs[3331] = (layer4_outputs[1388]) ^ (layer4_outputs[385]);
    assign layer5_outputs[3332] = ~((layer4_outputs[4218]) & (layer4_outputs[3828]));
    assign layer5_outputs[3333] = layer4_outputs[2192];
    assign layer5_outputs[3334] = ~(layer4_outputs[2533]) | (layer4_outputs[1533]);
    assign layer5_outputs[3335] = ~((layer4_outputs[4810]) | (layer4_outputs[3171]));
    assign layer5_outputs[3336] = ~(layer4_outputs[4882]);
    assign layer5_outputs[3337] = layer4_outputs[4815];
    assign layer5_outputs[3338] = ~(layer4_outputs[1330]);
    assign layer5_outputs[3339] = (layer4_outputs[1237]) ^ (layer4_outputs[2469]);
    assign layer5_outputs[3340] = ~((layer4_outputs[4294]) ^ (layer4_outputs[2]));
    assign layer5_outputs[3341] = (layer4_outputs[226]) ^ (layer4_outputs[3834]);
    assign layer5_outputs[3342] = (layer4_outputs[1961]) & ~(layer4_outputs[696]);
    assign layer5_outputs[3343] = layer4_outputs[3446];
    assign layer5_outputs[3344] = (layer4_outputs[2686]) ^ (layer4_outputs[3472]);
    assign layer5_outputs[3345] = 1'b1;
    assign layer5_outputs[3346] = (layer4_outputs[4330]) & (layer4_outputs[4901]);
    assign layer5_outputs[3347] = ~(layer4_outputs[4048]);
    assign layer5_outputs[3348] = (layer4_outputs[2143]) & ~(layer4_outputs[4656]);
    assign layer5_outputs[3349] = ~(layer4_outputs[1263]);
    assign layer5_outputs[3350] = ~((layer4_outputs[1338]) | (layer4_outputs[4954]));
    assign layer5_outputs[3351] = ~(layer4_outputs[1164]);
    assign layer5_outputs[3352] = layer4_outputs[4814];
    assign layer5_outputs[3353] = (layer4_outputs[3538]) & ~(layer4_outputs[4758]);
    assign layer5_outputs[3354] = ~(layer4_outputs[940]) | (layer4_outputs[1645]);
    assign layer5_outputs[3355] = ~(layer4_outputs[3764]);
    assign layer5_outputs[3356] = ~(layer4_outputs[751]) | (layer4_outputs[268]);
    assign layer5_outputs[3357] = (layer4_outputs[3394]) | (layer4_outputs[2915]);
    assign layer5_outputs[3358] = ~(layer4_outputs[3164]);
    assign layer5_outputs[3359] = ~((layer4_outputs[2282]) | (layer4_outputs[2186]));
    assign layer5_outputs[3360] = ~(layer4_outputs[2406]);
    assign layer5_outputs[3361] = (layer4_outputs[919]) & ~(layer4_outputs[2564]);
    assign layer5_outputs[3362] = ~(layer4_outputs[4692]) | (layer4_outputs[713]);
    assign layer5_outputs[3363] = layer4_outputs[1878];
    assign layer5_outputs[3364] = ~(layer4_outputs[1416]) | (layer4_outputs[4941]);
    assign layer5_outputs[3365] = ~((layer4_outputs[1356]) & (layer4_outputs[1279]));
    assign layer5_outputs[3366] = layer4_outputs[3320];
    assign layer5_outputs[3367] = (layer4_outputs[511]) & (layer4_outputs[1175]);
    assign layer5_outputs[3368] = layer4_outputs[3847];
    assign layer5_outputs[3369] = ~(layer4_outputs[91]) | (layer4_outputs[1427]);
    assign layer5_outputs[3370] = (layer4_outputs[334]) ^ (layer4_outputs[643]);
    assign layer5_outputs[3371] = ~((layer4_outputs[2238]) | (layer4_outputs[3962]));
    assign layer5_outputs[3372] = (layer4_outputs[4414]) | (layer4_outputs[4380]);
    assign layer5_outputs[3373] = 1'b1;
    assign layer5_outputs[3374] = 1'b0;
    assign layer5_outputs[3375] = ~(layer4_outputs[1564]);
    assign layer5_outputs[3376] = ~(layer4_outputs[3426]);
    assign layer5_outputs[3377] = ~(layer4_outputs[5032]) | (layer4_outputs[403]);
    assign layer5_outputs[3378] = ~(layer4_outputs[4840]);
    assign layer5_outputs[3379] = ~((layer4_outputs[2143]) & (layer4_outputs[413]));
    assign layer5_outputs[3380] = (layer4_outputs[238]) & (layer4_outputs[555]);
    assign layer5_outputs[3381] = (layer4_outputs[223]) ^ (layer4_outputs[3054]);
    assign layer5_outputs[3382] = layer4_outputs[2316];
    assign layer5_outputs[3383] = (layer4_outputs[3350]) & (layer4_outputs[3871]);
    assign layer5_outputs[3384] = ~(layer4_outputs[4132]) | (layer4_outputs[1676]);
    assign layer5_outputs[3385] = layer4_outputs[1817];
    assign layer5_outputs[3386] = layer4_outputs[3083];
    assign layer5_outputs[3387] = layer4_outputs[1026];
    assign layer5_outputs[3388] = (layer4_outputs[3764]) | (layer4_outputs[1573]);
    assign layer5_outputs[3389] = ~(layer4_outputs[3678]);
    assign layer5_outputs[3390] = layer4_outputs[1418];
    assign layer5_outputs[3391] = ~((layer4_outputs[4334]) | (layer4_outputs[2005]));
    assign layer5_outputs[3392] = ~(layer4_outputs[3994]);
    assign layer5_outputs[3393] = ~((layer4_outputs[1954]) ^ (layer4_outputs[3027]));
    assign layer5_outputs[3394] = ~((layer4_outputs[4478]) | (layer4_outputs[3985]));
    assign layer5_outputs[3395] = ~(layer4_outputs[3592]) | (layer4_outputs[2272]);
    assign layer5_outputs[3396] = ~(layer4_outputs[1949]);
    assign layer5_outputs[3397] = (layer4_outputs[1242]) | (layer4_outputs[1109]);
    assign layer5_outputs[3398] = ~(layer4_outputs[691]);
    assign layer5_outputs[3399] = layer4_outputs[682];
    assign layer5_outputs[3400] = 1'b0;
    assign layer5_outputs[3401] = layer4_outputs[2560];
    assign layer5_outputs[3402] = ~((layer4_outputs[5014]) ^ (layer4_outputs[1310]));
    assign layer5_outputs[3403] = ~((layer4_outputs[4864]) & (layer4_outputs[3689]));
    assign layer5_outputs[3404] = ~(layer4_outputs[1064]);
    assign layer5_outputs[3405] = (layer4_outputs[4449]) & ~(layer4_outputs[1371]);
    assign layer5_outputs[3406] = ~(layer4_outputs[4523]);
    assign layer5_outputs[3407] = ~(layer4_outputs[3220]);
    assign layer5_outputs[3408] = (layer4_outputs[1020]) & ~(layer4_outputs[4676]);
    assign layer5_outputs[3409] = ~(layer4_outputs[4767]);
    assign layer5_outputs[3410] = (layer4_outputs[3762]) & ~(layer4_outputs[1484]);
    assign layer5_outputs[3411] = (layer4_outputs[2722]) & ~(layer4_outputs[69]);
    assign layer5_outputs[3412] = layer4_outputs[4845];
    assign layer5_outputs[3413] = (layer4_outputs[3108]) & ~(layer4_outputs[2935]);
    assign layer5_outputs[3414] = layer4_outputs[151];
    assign layer5_outputs[3415] = ~(layer4_outputs[4997]);
    assign layer5_outputs[3416] = (layer4_outputs[816]) ^ (layer4_outputs[3977]);
    assign layer5_outputs[3417] = ~(layer4_outputs[1483]) | (layer4_outputs[2847]);
    assign layer5_outputs[3418] = ~((layer4_outputs[4834]) ^ (layer4_outputs[3738]));
    assign layer5_outputs[3419] = layer4_outputs[1152];
    assign layer5_outputs[3420] = layer4_outputs[5070];
    assign layer5_outputs[3421] = (layer4_outputs[2239]) & (layer4_outputs[613]);
    assign layer5_outputs[3422] = ~(layer4_outputs[138]) | (layer4_outputs[949]);
    assign layer5_outputs[3423] = ~((layer4_outputs[4]) | (layer4_outputs[19]));
    assign layer5_outputs[3424] = (layer4_outputs[2496]) & ~(layer4_outputs[3782]);
    assign layer5_outputs[3425] = (layer4_outputs[471]) & (layer4_outputs[3338]);
    assign layer5_outputs[3426] = layer4_outputs[291];
    assign layer5_outputs[3427] = ~(layer4_outputs[3386]) | (layer4_outputs[3020]);
    assign layer5_outputs[3428] = ~(layer4_outputs[2292]);
    assign layer5_outputs[3429] = (layer4_outputs[4035]) ^ (layer4_outputs[377]);
    assign layer5_outputs[3430] = (layer4_outputs[1756]) & (layer4_outputs[790]);
    assign layer5_outputs[3431] = layer4_outputs[202];
    assign layer5_outputs[3432] = ~(layer4_outputs[4904]);
    assign layer5_outputs[3433] = layer4_outputs[2941];
    assign layer5_outputs[3434] = ~(layer4_outputs[1716]) | (layer4_outputs[4193]);
    assign layer5_outputs[3435] = (layer4_outputs[1062]) ^ (layer4_outputs[3246]);
    assign layer5_outputs[3436] = ~(layer4_outputs[1216]);
    assign layer5_outputs[3437] = 1'b0;
    assign layer5_outputs[3438] = ~((layer4_outputs[871]) & (layer4_outputs[4829]));
    assign layer5_outputs[3439] = layer4_outputs[3510];
    assign layer5_outputs[3440] = layer4_outputs[2488];
    assign layer5_outputs[3441] = (layer4_outputs[4304]) & (layer4_outputs[2523]);
    assign layer5_outputs[3442] = ~(layer4_outputs[4305]);
    assign layer5_outputs[3443] = layer4_outputs[2081];
    assign layer5_outputs[3444] = ~(layer4_outputs[2120]);
    assign layer5_outputs[3445] = layer4_outputs[125];
    assign layer5_outputs[3446] = layer4_outputs[449];
    assign layer5_outputs[3447] = ~(layer4_outputs[4090]);
    assign layer5_outputs[3448] = ~(layer4_outputs[4374]);
    assign layer5_outputs[3449] = ~(layer4_outputs[3461]);
    assign layer5_outputs[3450] = ~(layer4_outputs[3805]);
    assign layer5_outputs[3451] = ~(layer4_outputs[3605]);
    assign layer5_outputs[3452] = (layer4_outputs[2249]) & (layer4_outputs[4628]);
    assign layer5_outputs[3453] = layer4_outputs[3621];
    assign layer5_outputs[3454] = layer4_outputs[3695];
    assign layer5_outputs[3455] = (layer4_outputs[3083]) & (layer4_outputs[2332]);
    assign layer5_outputs[3456] = layer4_outputs[583];
    assign layer5_outputs[3457] = ~(layer4_outputs[5008]);
    assign layer5_outputs[3458] = ~((layer4_outputs[273]) & (layer4_outputs[3069]));
    assign layer5_outputs[3459] = 1'b0;
    assign layer5_outputs[3460] = layer4_outputs[550];
    assign layer5_outputs[3461] = layer4_outputs[4958];
    assign layer5_outputs[3462] = ~(layer4_outputs[3167]);
    assign layer5_outputs[3463] = layer4_outputs[2873];
    assign layer5_outputs[3464] = ~(layer4_outputs[848]) | (layer4_outputs[4846]);
    assign layer5_outputs[3465] = layer4_outputs[884];
    assign layer5_outputs[3466] = ~((layer4_outputs[4969]) | (layer4_outputs[4196]));
    assign layer5_outputs[3467] = (layer4_outputs[4288]) | (layer4_outputs[2981]);
    assign layer5_outputs[3468] = ~(layer4_outputs[2601]);
    assign layer5_outputs[3469] = (layer4_outputs[3847]) & ~(layer4_outputs[1561]);
    assign layer5_outputs[3470] = ~(layer4_outputs[4553]) | (layer4_outputs[3466]);
    assign layer5_outputs[3471] = (layer4_outputs[1742]) & (layer4_outputs[623]);
    assign layer5_outputs[3472] = ~(layer4_outputs[652]) | (layer4_outputs[1343]);
    assign layer5_outputs[3473] = ~((layer4_outputs[2613]) & (layer4_outputs[1642]));
    assign layer5_outputs[3474] = ~(layer4_outputs[3276]);
    assign layer5_outputs[3475] = ~(layer4_outputs[4798]);
    assign layer5_outputs[3476] = ~(layer4_outputs[1247]);
    assign layer5_outputs[3477] = (layer4_outputs[3077]) & (layer4_outputs[252]);
    assign layer5_outputs[3478] = ~((layer4_outputs[2588]) ^ (layer4_outputs[1578]));
    assign layer5_outputs[3479] = (layer4_outputs[4333]) & ~(layer4_outputs[4404]);
    assign layer5_outputs[3480] = (layer4_outputs[3468]) & (layer4_outputs[4699]);
    assign layer5_outputs[3481] = layer4_outputs[2283];
    assign layer5_outputs[3482] = ~((layer4_outputs[2527]) & (layer4_outputs[1618]));
    assign layer5_outputs[3483] = ~((layer4_outputs[367]) | (layer4_outputs[1197]));
    assign layer5_outputs[3484] = ~(layer4_outputs[274]);
    assign layer5_outputs[3485] = ~(layer4_outputs[1736]);
    assign layer5_outputs[3486] = (layer4_outputs[536]) & (layer4_outputs[2323]);
    assign layer5_outputs[3487] = ~(layer4_outputs[4697]);
    assign layer5_outputs[3488] = layer4_outputs[3603];
    assign layer5_outputs[3489] = (layer4_outputs[88]) & ~(layer4_outputs[2692]);
    assign layer5_outputs[3490] = ~(layer4_outputs[3260]);
    assign layer5_outputs[3491] = 1'b1;
    assign layer5_outputs[3492] = layer4_outputs[3893];
    assign layer5_outputs[3493] = ~((layer4_outputs[4634]) | (layer4_outputs[1225]));
    assign layer5_outputs[3494] = ~(layer4_outputs[2532]) | (layer4_outputs[502]);
    assign layer5_outputs[3495] = ~((layer4_outputs[4714]) & (layer4_outputs[3382]));
    assign layer5_outputs[3496] = layer4_outputs[5109];
    assign layer5_outputs[3497] = layer4_outputs[2809];
    assign layer5_outputs[3498] = (layer4_outputs[198]) & (layer4_outputs[1694]);
    assign layer5_outputs[3499] = layer4_outputs[1441];
    assign layer5_outputs[3500] = (layer4_outputs[2598]) & ~(layer4_outputs[4300]);
    assign layer5_outputs[3501] = (layer4_outputs[4901]) & (layer4_outputs[1495]);
    assign layer5_outputs[3502] = (layer4_outputs[3077]) ^ (layer4_outputs[1668]);
    assign layer5_outputs[3503] = layer4_outputs[3443];
    assign layer5_outputs[3504] = layer4_outputs[2559];
    assign layer5_outputs[3505] = (layer4_outputs[1368]) & (layer4_outputs[4481]);
    assign layer5_outputs[3506] = (layer4_outputs[915]) | (layer4_outputs[2110]);
    assign layer5_outputs[3507] = ~((layer4_outputs[4353]) & (layer4_outputs[605]));
    assign layer5_outputs[3508] = layer4_outputs[3145];
    assign layer5_outputs[3509] = ~(layer4_outputs[4343]) | (layer4_outputs[4337]);
    assign layer5_outputs[3510] = layer4_outputs[3652];
    assign layer5_outputs[3511] = ~((layer4_outputs[4987]) & (layer4_outputs[2011]));
    assign layer5_outputs[3512] = ~((layer4_outputs[389]) ^ (layer4_outputs[2320]));
    assign layer5_outputs[3513] = ~(layer4_outputs[4548]) | (layer4_outputs[2058]);
    assign layer5_outputs[3514] = ~(layer4_outputs[910]);
    assign layer5_outputs[3515] = layer4_outputs[3525];
    assign layer5_outputs[3516] = 1'b1;
    assign layer5_outputs[3517] = layer4_outputs[5011];
    assign layer5_outputs[3518] = ~(layer4_outputs[5031]) | (layer4_outputs[657]);
    assign layer5_outputs[3519] = ~((layer4_outputs[2766]) | (layer4_outputs[560]));
    assign layer5_outputs[3520] = ~(layer4_outputs[2918]) | (layer4_outputs[1831]);
    assign layer5_outputs[3521] = ~(layer4_outputs[1558]);
    assign layer5_outputs[3522] = layer4_outputs[2374];
    assign layer5_outputs[3523] = ~((layer4_outputs[952]) ^ (layer4_outputs[4858]));
    assign layer5_outputs[3524] = layer4_outputs[663];
    assign layer5_outputs[3525] = ~((layer4_outputs[2498]) & (layer4_outputs[3329]));
    assign layer5_outputs[3526] = ~((layer4_outputs[2233]) | (layer4_outputs[3327]));
    assign layer5_outputs[3527] = (layer4_outputs[2517]) & ~(layer4_outputs[1962]);
    assign layer5_outputs[3528] = ~(layer4_outputs[3682]);
    assign layer5_outputs[3529] = ~(layer4_outputs[1386]) | (layer4_outputs[3602]);
    assign layer5_outputs[3530] = (layer4_outputs[3560]) ^ (layer4_outputs[860]);
    assign layer5_outputs[3531] = layer4_outputs[93];
    assign layer5_outputs[3532] = (layer4_outputs[3688]) ^ (layer4_outputs[20]);
    assign layer5_outputs[3533] = 1'b0;
    assign layer5_outputs[3534] = ~(layer4_outputs[720]);
    assign layer5_outputs[3535] = ~(layer4_outputs[2563]);
    assign layer5_outputs[3536] = ~(layer4_outputs[2530]);
    assign layer5_outputs[3537] = ~(layer4_outputs[1932]);
    assign layer5_outputs[3538] = layer4_outputs[3771];
    assign layer5_outputs[3539] = ~((layer4_outputs[3050]) ^ (layer4_outputs[4813]));
    assign layer5_outputs[3540] = ~(layer4_outputs[1016]) | (layer4_outputs[3912]);
    assign layer5_outputs[3541] = ~(layer4_outputs[771]);
    assign layer5_outputs[3542] = ~(layer4_outputs[1712]);
    assign layer5_outputs[3543] = layer4_outputs[4633];
    assign layer5_outputs[3544] = ~(layer4_outputs[4102]);
    assign layer5_outputs[3545] = ~(layer4_outputs[4936]);
    assign layer5_outputs[3546] = ~(layer4_outputs[5035]);
    assign layer5_outputs[3547] = ~((layer4_outputs[832]) & (layer4_outputs[4490]));
    assign layer5_outputs[3548] = layer4_outputs[4250];
    assign layer5_outputs[3549] = layer4_outputs[3403];
    assign layer5_outputs[3550] = ~(layer4_outputs[2039]);
    assign layer5_outputs[3551] = ~((layer4_outputs[1759]) ^ (layer4_outputs[624]));
    assign layer5_outputs[3552] = ~(layer4_outputs[1755]);
    assign layer5_outputs[3553] = (layer4_outputs[1429]) & ~(layer4_outputs[2841]);
    assign layer5_outputs[3554] = ~((layer4_outputs[1217]) ^ (layer4_outputs[1406]));
    assign layer5_outputs[3555] = ~(layer4_outputs[4373]);
    assign layer5_outputs[3556] = ~(layer4_outputs[3530]);
    assign layer5_outputs[3557] = 1'b1;
    assign layer5_outputs[3558] = ~(layer4_outputs[3477]);
    assign layer5_outputs[3559] = ~(layer4_outputs[4727]);
    assign layer5_outputs[3560] = (layer4_outputs[3344]) & ~(layer4_outputs[2050]);
    assign layer5_outputs[3561] = layer4_outputs[859];
    assign layer5_outputs[3562] = layer4_outputs[2840];
    assign layer5_outputs[3563] = ~((layer4_outputs[3129]) | (layer4_outputs[3628]));
    assign layer5_outputs[3564] = ~((layer4_outputs[370]) | (layer4_outputs[2470]));
    assign layer5_outputs[3565] = (layer4_outputs[4860]) ^ (layer4_outputs[4355]);
    assign layer5_outputs[3566] = ~(layer4_outputs[4943]);
    assign layer5_outputs[3567] = ~((layer4_outputs[2651]) ^ (layer4_outputs[2362]));
    assign layer5_outputs[3568] = ~(layer4_outputs[3339]);
    assign layer5_outputs[3569] = (layer4_outputs[900]) | (layer4_outputs[2180]);
    assign layer5_outputs[3570] = ~(layer4_outputs[4469]) | (layer4_outputs[2286]);
    assign layer5_outputs[3571] = ~(layer4_outputs[1561]);
    assign layer5_outputs[3572] = ~(layer4_outputs[1706]) | (layer4_outputs[4629]);
    assign layer5_outputs[3573] = (layer4_outputs[861]) | (layer4_outputs[319]);
    assign layer5_outputs[3574] = ~((layer4_outputs[3350]) | (layer4_outputs[3017]));
    assign layer5_outputs[3575] = ~(layer4_outputs[2795]) | (layer4_outputs[2354]);
    assign layer5_outputs[3576] = 1'b0;
    assign layer5_outputs[3577] = 1'b1;
    assign layer5_outputs[3578] = (layer4_outputs[2313]) & ~(layer4_outputs[2394]);
    assign layer5_outputs[3579] = ~((layer4_outputs[2206]) | (layer4_outputs[4685]));
    assign layer5_outputs[3580] = layer4_outputs[2381];
    assign layer5_outputs[3581] = layer4_outputs[83];
    assign layer5_outputs[3582] = (layer4_outputs[4932]) ^ (layer4_outputs[1209]);
    assign layer5_outputs[3583] = (layer4_outputs[3014]) & ~(layer4_outputs[2224]);
    assign layer5_outputs[3584] = ~(layer4_outputs[5091]);
    assign layer5_outputs[3585] = layer4_outputs[2540];
    assign layer5_outputs[3586] = 1'b0;
    assign layer5_outputs[3587] = ~(layer4_outputs[2605]) | (layer4_outputs[4894]);
    assign layer5_outputs[3588] = ~(layer4_outputs[2876]);
    assign layer5_outputs[3589] = layer4_outputs[1145];
    assign layer5_outputs[3590] = layer4_outputs[4876];
    assign layer5_outputs[3591] = ~((layer4_outputs[3753]) | (layer4_outputs[4372]));
    assign layer5_outputs[3592] = layer4_outputs[2233];
    assign layer5_outputs[3593] = ~(layer4_outputs[3141]);
    assign layer5_outputs[3594] = layer4_outputs[4887];
    assign layer5_outputs[3595] = layer4_outputs[929];
    assign layer5_outputs[3596] = layer4_outputs[3172];
    assign layer5_outputs[3597] = layer4_outputs[747];
    assign layer5_outputs[3598] = ~((layer4_outputs[512]) & (layer4_outputs[4451]));
    assign layer5_outputs[3599] = ~((layer4_outputs[3182]) ^ (layer4_outputs[4620]));
    assign layer5_outputs[3600] = ~((layer4_outputs[4599]) ^ (layer4_outputs[2019]));
    assign layer5_outputs[3601] = (layer4_outputs[3272]) | (layer4_outputs[777]);
    assign layer5_outputs[3602] = 1'b1;
    assign layer5_outputs[3603] = ~((layer4_outputs[4710]) | (layer4_outputs[2907]));
    assign layer5_outputs[3604] = (layer4_outputs[4196]) & (layer4_outputs[2688]);
    assign layer5_outputs[3605] = (layer4_outputs[4168]) ^ (layer4_outputs[615]);
    assign layer5_outputs[3606] = ~(layer4_outputs[1792]);
    assign layer5_outputs[3607] = ~(layer4_outputs[4767]) | (layer4_outputs[2634]);
    assign layer5_outputs[3608] = ~(layer4_outputs[4185]);
    assign layer5_outputs[3609] = (layer4_outputs[4322]) ^ (layer4_outputs[1032]);
    assign layer5_outputs[3610] = (layer4_outputs[3778]) & ~(layer4_outputs[2606]);
    assign layer5_outputs[3611] = layer4_outputs[3196];
    assign layer5_outputs[3612] = ~(layer4_outputs[495]);
    assign layer5_outputs[3613] = ~(layer4_outputs[4548]);
    assign layer5_outputs[3614] = ~(layer4_outputs[3952]);
    assign layer5_outputs[3615] = (layer4_outputs[2048]) ^ (layer4_outputs[1741]);
    assign layer5_outputs[3616] = ~((layer4_outputs[1039]) | (layer4_outputs[4574]));
    assign layer5_outputs[3617] = layer4_outputs[353];
    assign layer5_outputs[3618] = ~(layer4_outputs[2987]) | (layer4_outputs[1774]);
    assign layer5_outputs[3619] = layer4_outputs[3435];
    assign layer5_outputs[3620] = ~(layer4_outputs[4188]);
    assign layer5_outputs[3621] = ~((layer4_outputs[5102]) | (layer4_outputs[200]));
    assign layer5_outputs[3622] = ~(layer4_outputs[4616]);
    assign layer5_outputs[3623] = 1'b0;
    assign layer5_outputs[3624] = (layer4_outputs[544]) | (layer4_outputs[1982]);
    assign layer5_outputs[3625] = ~(layer4_outputs[1531]);
    assign layer5_outputs[3626] = (layer4_outputs[63]) & (layer4_outputs[4753]);
    assign layer5_outputs[3627] = ~(layer4_outputs[1168]);
    assign layer5_outputs[3628] = (layer4_outputs[500]) & (layer4_outputs[4580]);
    assign layer5_outputs[3629] = (layer4_outputs[1077]) & ~(layer4_outputs[1853]);
    assign layer5_outputs[3630] = ~(layer4_outputs[2653]);
    assign layer5_outputs[3631] = layer4_outputs[2280];
    assign layer5_outputs[3632] = (layer4_outputs[1667]) ^ (layer4_outputs[525]);
    assign layer5_outputs[3633] = ~((layer4_outputs[2979]) | (layer4_outputs[130]));
    assign layer5_outputs[3634] = ~(layer4_outputs[3219]) | (layer4_outputs[4354]);
    assign layer5_outputs[3635] = layer4_outputs[458];
    assign layer5_outputs[3636] = (layer4_outputs[3474]) | (layer4_outputs[4438]);
    assign layer5_outputs[3637] = layer4_outputs[1101];
    assign layer5_outputs[3638] = layer4_outputs[2436];
    assign layer5_outputs[3639] = (layer4_outputs[4915]) & ~(layer4_outputs[3533]);
    assign layer5_outputs[3640] = layer4_outputs[2798];
    assign layer5_outputs[3641] = layer4_outputs[1044];
    assign layer5_outputs[3642] = ~(layer4_outputs[4054]);
    assign layer5_outputs[3643] = ~(layer4_outputs[341]) | (layer4_outputs[1361]);
    assign layer5_outputs[3644] = 1'b1;
    assign layer5_outputs[3645] = ~(layer4_outputs[2307]) | (layer4_outputs[255]);
    assign layer5_outputs[3646] = ~(layer4_outputs[1321]);
    assign layer5_outputs[3647] = layer4_outputs[649];
    assign layer5_outputs[3648] = (layer4_outputs[4150]) & ~(layer4_outputs[1939]);
    assign layer5_outputs[3649] = ~((layer4_outputs[1734]) | (layer4_outputs[4492]));
    assign layer5_outputs[3650] = (layer4_outputs[137]) ^ (layer4_outputs[4608]);
    assign layer5_outputs[3651] = ~(layer4_outputs[2597]);
    assign layer5_outputs[3652] = layer4_outputs[211];
    assign layer5_outputs[3653] = layer4_outputs[2431];
    assign layer5_outputs[3654] = (layer4_outputs[4698]) & (layer4_outputs[3455]);
    assign layer5_outputs[3655] = (layer4_outputs[4979]) & (layer4_outputs[3703]);
    assign layer5_outputs[3656] = ~(layer4_outputs[236]);
    assign layer5_outputs[3657] = ~(layer4_outputs[2462]);
    assign layer5_outputs[3658] = ~(layer4_outputs[4274]);
    assign layer5_outputs[3659] = ~(layer4_outputs[4824]) | (layer4_outputs[4090]);
    assign layer5_outputs[3660] = 1'b0;
    assign layer5_outputs[3661] = layer4_outputs[3931];
    assign layer5_outputs[3662] = (layer4_outputs[3516]) | (layer4_outputs[2460]);
    assign layer5_outputs[3663] = (layer4_outputs[836]) & (layer4_outputs[3449]);
    assign layer5_outputs[3664] = layer4_outputs[2301];
    assign layer5_outputs[3665] = ~(layer4_outputs[2277]);
    assign layer5_outputs[3666] = (layer4_outputs[1095]) ^ (layer4_outputs[1911]);
    assign layer5_outputs[3667] = ~(layer4_outputs[4695]);
    assign layer5_outputs[3668] = (layer4_outputs[1631]) & ~(layer4_outputs[2418]);
    assign layer5_outputs[3669] = ~(layer4_outputs[1119]);
    assign layer5_outputs[3670] = ~(layer4_outputs[2518]) | (layer4_outputs[3602]);
    assign layer5_outputs[3671] = ~(layer4_outputs[4721]);
    assign layer5_outputs[3672] = ~(layer4_outputs[4597]);
    assign layer5_outputs[3673] = layer4_outputs[2346];
    assign layer5_outputs[3674] = ~(layer4_outputs[4494]);
    assign layer5_outputs[3675] = (layer4_outputs[1597]) & ~(layer4_outputs[3836]);
    assign layer5_outputs[3676] = (layer4_outputs[2540]) | (layer4_outputs[1368]);
    assign layer5_outputs[3677] = layer4_outputs[660];
    assign layer5_outputs[3678] = (layer4_outputs[1468]) & (layer4_outputs[4214]);
    assign layer5_outputs[3679] = ~((layer4_outputs[380]) ^ (layer4_outputs[2310]));
    assign layer5_outputs[3680] = ~((layer4_outputs[87]) & (layer4_outputs[4299]));
    assign layer5_outputs[3681] = layer4_outputs[1678];
    assign layer5_outputs[3682] = ~(layer4_outputs[188]);
    assign layer5_outputs[3683] = ~(layer4_outputs[4036]);
    assign layer5_outputs[3684] = (layer4_outputs[3853]) & (layer4_outputs[4062]);
    assign layer5_outputs[3685] = ~((layer4_outputs[2281]) & (layer4_outputs[2489]));
    assign layer5_outputs[3686] = ~(layer4_outputs[25]);
    assign layer5_outputs[3687] = (layer4_outputs[4884]) | (layer4_outputs[3933]);
    assign layer5_outputs[3688] = layer4_outputs[3288];
    assign layer5_outputs[3689] = (layer4_outputs[818]) & (layer4_outputs[4043]);
    assign layer5_outputs[3690] = layer4_outputs[4325];
    assign layer5_outputs[3691] = ~((layer4_outputs[2216]) & (layer4_outputs[4375]));
    assign layer5_outputs[3692] = (layer4_outputs[5107]) | (layer4_outputs[2086]);
    assign layer5_outputs[3693] = layer4_outputs[264];
    assign layer5_outputs[3694] = (layer4_outputs[3848]) & ~(layer4_outputs[4628]);
    assign layer5_outputs[3695] = ~(layer4_outputs[55]);
    assign layer5_outputs[3696] = layer4_outputs[2099];
    assign layer5_outputs[3697] = ~((layer4_outputs[3858]) ^ (layer4_outputs[1502]));
    assign layer5_outputs[3698] = (layer4_outputs[4134]) & ~(layer4_outputs[4781]);
    assign layer5_outputs[3699] = ~(layer4_outputs[4427]) | (layer4_outputs[621]);
    assign layer5_outputs[3700] = layer4_outputs[342];
    assign layer5_outputs[3701] = ~(layer4_outputs[854]);
    assign layer5_outputs[3702] = ~(layer4_outputs[3637]);
    assign layer5_outputs[3703] = layer4_outputs[3980];
    assign layer5_outputs[3704] = layer4_outputs[2214];
    assign layer5_outputs[3705] = ~(layer4_outputs[489]) | (layer4_outputs[3544]);
    assign layer5_outputs[3706] = (layer4_outputs[4579]) & (layer4_outputs[4437]);
    assign layer5_outputs[3707] = layer4_outputs[4642];
    assign layer5_outputs[3708] = (layer4_outputs[292]) ^ (layer4_outputs[122]);
    assign layer5_outputs[3709] = ~(layer4_outputs[1136]) | (layer4_outputs[3112]);
    assign layer5_outputs[3710] = (layer4_outputs[1601]) & (layer4_outputs[4370]);
    assign layer5_outputs[3711] = layer4_outputs[3136];
    assign layer5_outputs[3712] = ~((layer4_outputs[4503]) & (layer4_outputs[4388]));
    assign layer5_outputs[3713] = 1'b0;
    assign layer5_outputs[3714] = ~(layer4_outputs[3306]) | (layer4_outputs[2973]);
    assign layer5_outputs[3715] = layer4_outputs[27];
    assign layer5_outputs[3716] = (layer4_outputs[2351]) & ~(layer4_outputs[2327]);
    assign layer5_outputs[3717] = ~(layer4_outputs[2416]);
    assign layer5_outputs[3718] = layer4_outputs[970];
    assign layer5_outputs[3719] = (layer4_outputs[2458]) & ~(layer4_outputs[4706]);
    assign layer5_outputs[3720] = ~(layer4_outputs[3889]);
    assign layer5_outputs[3721] = layer4_outputs[1258];
    assign layer5_outputs[3722] = (layer4_outputs[1053]) & (layer4_outputs[606]);
    assign layer5_outputs[3723] = ~(layer4_outputs[4788]);
    assign layer5_outputs[3724] = ~(layer4_outputs[4252]);
    assign layer5_outputs[3725] = ~(layer4_outputs[906]);
    assign layer5_outputs[3726] = layer4_outputs[1869];
    assign layer5_outputs[3727] = ~(layer4_outputs[4958]);
    assign layer5_outputs[3728] = ~((layer4_outputs[4441]) & (layer4_outputs[1953]));
    assign layer5_outputs[3729] = ~(layer4_outputs[275]);
    assign layer5_outputs[3730] = (layer4_outputs[3767]) ^ (layer4_outputs[3330]);
    assign layer5_outputs[3731] = ~(layer4_outputs[4701]);
    assign layer5_outputs[3732] = layer4_outputs[1479];
    assign layer5_outputs[3733] = layer4_outputs[4846];
    assign layer5_outputs[3734] = layer4_outputs[2991];
    assign layer5_outputs[3735] = (layer4_outputs[562]) ^ (layer4_outputs[1451]);
    assign layer5_outputs[3736] = layer4_outputs[1449];
    assign layer5_outputs[3737] = layer4_outputs[1779];
    assign layer5_outputs[3738] = (layer4_outputs[1709]) & (layer4_outputs[3929]);
    assign layer5_outputs[3739] = ~(layer4_outputs[2869]) | (layer4_outputs[1051]);
    assign layer5_outputs[3740] = layer4_outputs[733];
    assign layer5_outputs[3741] = ~((layer4_outputs[4198]) & (layer4_outputs[436]));
    assign layer5_outputs[3742] = layer4_outputs[314];
    assign layer5_outputs[3743] = ~(layer4_outputs[683]) | (layer4_outputs[4456]);
    assign layer5_outputs[3744] = layer4_outputs[1934];
    assign layer5_outputs[3745] = (layer4_outputs[3022]) & ~(layer4_outputs[4001]);
    assign layer5_outputs[3746] = layer4_outputs[4463];
    assign layer5_outputs[3747] = ~((layer4_outputs[801]) & (layer4_outputs[3592]));
    assign layer5_outputs[3748] = layer4_outputs[4560];
    assign layer5_outputs[3749] = layer4_outputs[4441];
    assign layer5_outputs[3750] = ~((layer4_outputs[3851]) ^ (layer4_outputs[4290]));
    assign layer5_outputs[3751] = (layer4_outputs[3777]) & (layer4_outputs[2811]);
    assign layer5_outputs[3752] = (layer4_outputs[2345]) & ~(layer4_outputs[426]);
    assign layer5_outputs[3753] = (layer4_outputs[1448]) ^ (layer4_outputs[4896]);
    assign layer5_outputs[3754] = ~(layer4_outputs[3336]) | (layer4_outputs[4199]);
    assign layer5_outputs[3755] = ~(layer4_outputs[2631]) | (layer4_outputs[272]);
    assign layer5_outputs[3756] = ~(layer4_outputs[1015]);
    assign layer5_outputs[3757] = ~((layer4_outputs[3643]) & (layer4_outputs[4300]));
    assign layer5_outputs[3758] = 1'b1;
    assign layer5_outputs[3759] = (layer4_outputs[4513]) & (layer4_outputs[3151]);
    assign layer5_outputs[3760] = layer4_outputs[4685];
    assign layer5_outputs[3761] = ~((layer4_outputs[2290]) | (layer4_outputs[1629]));
    assign layer5_outputs[3762] = ~(layer4_outputs[3553]);
    assign layer5_outputs[3763] = (layer4_outputs[4702]) ^ (layer4_outputs[2577]);
    assign layer5_outputs[3764] = (layer4_outputs[41]) & (layer4_outputs[3666]);
    assign layer5_outputs[3765] = layer4_outputs[821];
    assign layer5_outputs[3766] = ~(layer4_outputs[667]);
    assign layer5_outputs[3767] = ~((layer4_outputs[1006]) ^ (layer4_outputs[558]));
    assign layer5_outputs[3768] = ~(layer4_outputs[1228]);
    assign layer5_outputs[3769] = ~(layer4_outputs[1995]);
    assign layer5_outputs[3770] = ~(layer4_outputs[3954]);
    assign layer5_outputs[3771] = 1'b1;
    assign layer5_outputs[3772] = 1'b1;
    assign layer5_outputs[3773] = ~(layer4_outputs[234]) | (layer4_outputs[102]);
    assign layer5_outputs[3774] = layer4_outputs[3998];
    assign layer5_outputs[3775] = layer4_outputs[3532];
    assign layer5_outputs[3776] = (layer4_outputs[201]) ^ (layer4_outputs[1131]);
    assign layer5_outputs[3777] = (layer4_outputs[1677]) & ~(layer4_outputs[3619]);
    assign layer5_outputs[3778] = layer4_outputs[2330];
    assign layer5_outputs[3779] = ~((layer4_outputs[4292]) ^ (layer4_outputs[3601]));
    assign layer5_outputs[3780] = layer4_outputs[1467];
    assign layer5_outputs[3781] = ~((layer4_outputs[2497]) ^ (layer4_outputs[1582]));
    assign layer5_outputs[3782] = ~(layer4_outputs[808]);
    assign layer5_outputs[3783] = layer4_outputs[746];
    assign layer5_outputs[3784] = ~(layer4_outputs[4211]);
    assign layer5_outputs[3785] = (layer4_outputs[1740]) & ~(layer4_outputs[50]);
    assign layer5_outputs[3786] = layer4_outputs[1998];
    assign layer5_outputs[3787] = (layer4_outputs[3010]) | (layer4_outputs[3819]);
    assign layer5_outputs[3788] = (layer4_outputs[707]) & (layer4_outputs[418]);
    assign layer5_outputs[3789] = ~((layer4_outputs[3481]) & (layer4_outputs[1758]));
    assign layer5_outputs[3790] = ~(layer4_outputs[2144]) | (layer4_outputs[1301]);
    assign layer5_outputs[3791] = layer4_outputs[1555];
    assign layer5_outputs[3792] = ~((layer4_outputs[2819]) ^ (layer4_outputs[3209]));
    assign layer5_outputs[3793] = (layer4_outputs[1334]) ^ (layer4_outputs[4607]);
    assign layer5_outputs[3794] = ~(layer4_outputs[4893]);
    assign layer5_outputs[3795] = layer4_outputs[4057];
    assign layer5_outputs[3796] = (layer4_outputs[4342]) ^ (layer4_outputs[3143]);
    assign layer5_outputs[3797] = ~((layer4_outputs[2602]) ^ (layer4_outputs[1841]));
    assign layer5_outputs[3798] = (layer4_outputs[1333]) ^ (layer4_outputs[4351]);
    assign layer5_outputs[3799] = layer4_outputs[493];
    assign layer5_outputs[3800] = 1'b1;
    assign layer5_outputs[3801] = (layer4_outputs[5095]) & (layer4_outputs[2343]);
    assign layer5_outputs[3802] = layer4_outputs[257];
    assign layer5_outputs[3803] = (layer4_outputs[2849]) & ~(layer4_outputs[2906]);
    assign layer5_outputs[3804] = ~((layer4_outputs[314]) ^ (layer4_outputs[4920]));
    assign layer5_outputs[3805] = layer4_outputs[1931];
    assign layer5_outputs[3806] = ~((layer4_outputs[4002]) ^ (layer4_outputs[3856]));
    assign layer5_outputs[3807] = ~((layer4_outputs[1563]) | (layer4_outputs[4079]));
    assign layer5_outputs[3808] = ~(layer4_outputs[4511]);
    assign layer5_outputs[3809] = ~(layer4_outputs[2882]);
    assign layer5_outputs[3810] = ~(layer4_outputs[3058]);
    assign layer5_outputs[3811] = (layer4_outputs[3527]) & (layer4_outputs[2724]);
    assign layer5_outputs[3812] = layer4_outputs[3331];
    assign layer5_outputs[3813] = ~((layer4_outputs[4575]) ^ (layer4_outputs[2509]));
    assign layer5_outputs[3814] = layer4_outputs[752];
    assign layer5_outputs[3815] = 1'b1;
    assign layer5_outputs[3816] = (layer4_outputs[5092]) | (layer4_outputs[448]);
    assign layer5_outputs[3817] = (layer4_outputs[3270]) ^ (layer4_outputs[2648]);
    assign layer5_outputs[3818] = ~(layer4_outputs[518]);
    assign layer5_outputs[3819] = layer4_outputs[120];
    assign layer5_outputs[3820] = layer4_outputs[343];
    assign layer5_outputs[3821] = ~(layer4_outputs[3841]);
    assign layer5_outputs[3822] = layer4_outputs[3691];
    assign layer5_outputs[3823] = ~((layer4_outputs[2361]) ^ (layer4_outputs[4363]));
    assign layer5_outputs[3824] = (layer4_outputs[3258]) & ~(layer4_outputs[1884]);
    assign layer5_outputs[3825] = ~(layer4_outputs[4195]) | (layer4_outputs[4970]);
    assign layer5_outputs[3826] = ~(layer4_outputs[2469]);
    assign layer5_outputs[3827] = 1'b0;
    assign layer5_outputs[3828] = ~((layer4_outputs[1167]) | (layer4_outputs[847]));
    assign layer5_outputs[3829] = 1'b0;
    assign layer5_outputs[3830] = ~(layer4_outputs[395]);
    assign layer5_outputs[3831] = layer4_outputs[4951];
    assign layer5_outputs[3832] = ~(layer4_outputs[2725]);
    assign layer5_outputs[3833] = ~(layer4_outputs[4618]) | (layer4_outputs[3852]);
    assign layer5_outputs[3834] = 1'b0;
    assign layer5_outputs[3835] = ~(layer4_outputs[2210]) | (layer4_outputs[3015]);
    assign layer5_outputs[3836] = ~(layer4_outputs[4473]);
    assign layer5_outputs[3837] = ~(layer4_outputs[2706]);
    assign layer5_outputs[3838] = layer4_outputs[644];
    assign layer5_outputs[3839] = ~((layer4_outputs[1186]) ^ (layer4_outputs[4339]));
    assign layer5_outputs[3840] = ~((layer4_outputs[2269]) & (layer4_outputs[2551]));
    assign layer5_outputs[3841] = (layer4_outputs[131]) ^ (layer4_outputs[4389]);
    assign layer5_outputs[3842] = (layer4_outputs[2175]) & ~(layer4_outputs[2850]);
    assign layer5_outputs[3843] = (layer4_outputs[2833]) ^ (layer4_outputs[3315]);
    assign layer5_outputs[3844] = ~((layer4_outputs[973]) | (layer4_outputs[4801]));
    assign layer5_outputs[3845] = ~((layer4_outputs[275]) & (layer4_outputs[4072]));
    assign layer5_outputs[3846] = ~(layer4_outputs[93]);
    assign layer5_outputs[3847] = ~(layer4_outputs[2512]);
    assign layer5_outputs[3848] = ~((layer4_outputs[1446]) ^ (layer4_outputs[1566]));
    assign layer5_outputs[3849] = layer4_outputs[1174];
    assign layer5_outputs[3850] = ~(layer4_outputs[3640]);
    assign layer5_outputs[3851] = layer4_outputs[509];
    assign layer5_outputs[3852] = ~(layer4_outputs[2990]);
    assign layer5_outputs[3853] = ~(layer4_outputs[2445]) | (layer4_outputs[1500]);
    assign layer5_outputs[3854] = layer4_outputs[3861];
    assign layer5_outputs[3855] = ~(layer4_outputs[689]) | (layer4_outputs[3516]);
    assign layer5_outputs[3856] = ~((layer4_outputs[1606]) | (layer4_outputs[1433]));
    assign layer5_outputs[3857] = ~(layer4_outputs[2163]);
    assign layer5_outputs[3858] = ~(layer4_outputs[2728]) | (layer4_outputs[5060]);
    assign layer5_outputs[3859] = layer4_outputs[4177];
    assign layer5_outputs[3860] = layer4_outputs[4450];
    assign layer5_outputs[3861] = ~((layer4_outputs[3104]) & (layer4_outputs[1794]));
    assign layer5_outputs[3862] = layer4_outputs[351];
    assign layer5_outputs[3863] = ~(layer4_outputs[3955]) | (layer4_outputs[2187]);
    assign layer5_outputs[3864] = (layer4_outputs[608]) & ~(layer4_outputs[1360]);
    assign layer5_outputs[3865] = ~(layer4_outputs[626]);
    assign layer5_outputs[3866] = layer4_outputs[2364];
    assign layer5_outputs[3867] = (layer4_outputs[2983]) ^ (layer4_outputs[1134]);
    assign layer5_outputs[3868] = 1'b0;
    assign layer5_outputs[3869] = layer4_outputs[1230];
    assign layer5_outputs[3870] = layer4_outputs[1522];
    assign layer5_outputs[3871] = layer4_outputs[1135];
    assign layer5_outputs[3872] = layer4_outputs[738];
    assign layer5_outputs[3873] = (layer4_outputs[1528]) & (layer4_outputs[4474]);
    assign layer5_outputs[3874] = layer4_outputs[2484];
    assign layer5_outputs[3875] = ~(layer4_outputs[947]);
    assign layer5_outputs[3876] = (layer4_outputs[4916]) & ~(layer4_outputs[645]);
    assign layer5_outputs[3877] = ~(layer4_outputs[2295]);
    assign layer5_outputs[3878] = layer4_outputs[3707];
    assign layer5_outputs[3879] = ~(layer4_outputs[1049]);
    assign layer5_outputs[3880] = ~((layer4_outputs[4238]) | (layer4_outputs[2220]));
    assign layer5_outputs[3881] = (layer4_outputs[1148]) | (layer4_outputs[3907]);
    assign layer5_outputs[3882] = (layer4_outputs[1097]) & ~(layer4_outputs[1404]);
    assign layer5_outputs[3883] = ~(layer4_outputs[12]) | (layer4_outputs[390]);
    assign layer5_outputs[3884] = layer4_outputs[3978];
    assign layer5_outputs[3885] = ~((layer4_outputs[1970]) | (layer4_outputs[4769]));
    assign layer5_outputs[3886] = (layer4_outputs[2741]) & (layer4_outputs[2912]);
    assign layer5_outputs[3887] = ~((layer4_outputs[1797]) ^ (layer4_outputs[2087]));
    assign layer5_outputs[3888] = layer4_outputs[4128];
    assign layer5_outputs[3889] = ~(layer4_outputs[404]);
    assign layer5_outputs[3890] = (layer4_outputs[1669]) & ~(layer4_outputs[2917]);
    assign layer5_outputs[3891] = layer4_outputs[3631];
    assign layer5_outputs[3892] = (layer4_outputs[4083]) | (layer4_outputs[3]);
    assign layer5_outputs[3893] = layer4_outputs[159];
    assign layer5_outputs[3894] = ~((layer4_outputs[377]) | (layer4_outputs[3529]));
    assign layer5_outputs[3895] = (layer4_outputs[3704]) | (layer4_outputs[714]);
    assign layer5_outputs[3896] = ~((layer4_outputs[3360]) ^ (layer4_outputs[1157]));
    assign layer5_outputs[3897] = 1'b1;
    assign layer5_outputs[3898] = ~(layer4_outputs[503]);
    assign layer5_outputs[3899] = ~(layer4_outputs[4081]);
    assign layer5_outputs[3900] = ~(layer4_outputs[3947]);
    assign layer5_outputs[3901] = layer4_outputs[111];
    assign layer5_outputs[3902] = ~(layer4_outputs[4392]) | (layer4_outputs[3525]);
    assign layer5_outputs[3903] = layer4_outputs[797];
    assign layer5_outputs[3904] = ~(layer4_outputs[3093]);
    assign layer5_outputs[3905] = ~(layer4_outputs[4455]);
    assign layer5_outputs[3906] = ~(layer4_outputs[3080]);
    assign layer5_outputs[3907] = layer4_outputs[2764];
    assign layer5_outputs[3908] = (layer4_outputs[1670]) ^ (layer4_outputs[2532]);
    assign layer5_outputs[3909] = 1'b1;
    assign layer5_outputs[3910] = ~(layer4_outputs[4892]);
    assign layer5_outputs[3911] = layer4_outputs[2755];
    assign layer5_outputs[3912] = ~(layer4_outputs[146]) | (layer4_outputs[4957]);
    assign layer5_outputs[3913] = ~(layer4_outputs[1549]);
    assign layer5_outputs[3914] = ~(layer4_outputs[4776]);
    assign layer5_outputs[3915] = layer4_outputs[2712];
    assign layer5_outputs[3916] = (layer4_outputs[3015]) & (layer4_outputs[4487]);
    assign layer5_outputs[3917] = ~((layer4_outputs[2604]) ^ (layer4_outputs[2918]));
    assign layer5_outputs[3918] = ~(layer4_outputs[1957]) | (layer4_outputs[3366]);
    assign layer5_outputs[3919] = ~(layer4_outputs[2231]);
    assign layer5_outputs[3920] = layer4_outputs[3683];
    assign layer5_outputs[3921] = ~((layer4_outputs[702]) & (layer4_outputs[3928]));
    assign layer5_outputs[3922] = ~(layer4_outputs[4724]);
    assign layer5_outputs[3923] = ~((layer4_outputs[2478]) ^ (layer4_outputs[429]));
    assign layer5_outputs[3924] = (layer4_outputs[2171]) ^ (layer4_outputs[4233]);
    assign layer5_outputs[3925] = (layer4_outputs[3890]) ^ (layer4_outputs[2218]);
    assign layer5_outputs[3926] = ~((layer4_outputs[748]) | (layer4_outputs[396]));
    assign layer5_outputs[3927] = ~(layer4_outputs[3495]);
    assign layer5_outputs[3928] = ~(layer4_outputs[3856]);
    assign layer5_outputs[3929] = ~(layer4_outputs[3734]);
    assign layer5_outputs[3930] = (layer4_outputs[4387]) & ~(layer4_outputs[4690]);
    assign layer5_outputs[3931] = layer4_outputs[1588];
    assign layer5_outputs[3932] = layer4_outputs[1341];
    assign layer5_outputs[3933] = (layer4_outputs[1080]) & (layer4_outputs[3641]);
    assign layer5_outputs[3934] = ~((layer4_outputs[1647]) & (layer4_outputs[2090]));
    assign layer5_outputs[3935] = layer4_outputs[3484];
    assign layer5_outputs[3936] = ~(layer4_outputs[4087]) | (layer4_outputs[1459]);
    assign layer5_outputs[3937] = 1'b1;
    assign layer5_outputs[3938] = ~(layer4_outputs[770]);
    assign layer5_outputs[3939] = layer4_outputs[677];
    assign layer5_outputs[3940] = layer4_outputs[3819];
    assign layer5_outputs[3941] = (layer4_outputs[431]) | (layer4_outputs[2479]);
    assign layer5_outputs[3942] = layer4_outputs[309];
    assign layer5_outputs[3943] = 1'b1;
    assign layer5_outputs[3944] = ~(layer4_outputs[3774]);
    assign layer5_outputs[3945] = (layer4_outputs[1019]) ^ (layer4_outputs[1744]);
    assign layer5_outputs[3946] = 1'b0;
    assign layer5_outputs[3947] = ~(layer4_outputs[271]) | (layer4_outputs[2063]);
    assign layer5_outputs[3948] = layer4_outputs[3532];
    assign layer5_outputs[3949] = ~(layer4_outputs[235]) | (layer4_outputs[4707]);
    assign layer5_outputs[3950] = layer4_outputs[2208];
    assign layer5_outputs[3951] = (layer4_outputs[1457]) | (layer4_outputs[4282]);
    assign layer5_outputs[3952] = ~(layer4_outputs[1415]) | (layer4_outputs[4701]);
    assign layer5_outputs[3953] = layer4_outputs[163];
    assign layer5_outputs[3954] = (layer4_outputs[2256]) & ~(layer4_outputs[1545]);
    assign layer5_outputs[3955] = (layer4_outputs[1671]) ^ (layer4_outputs[2229]);
    assign layer5_outputs[3956] = layer4_outputs[999];
    assign layer5_outputs[3957] = (layer4_outputs[734]) & ~(layer4_outputs[2398]);
    assign layer5_outputs[3958] = layer4_outputs[698];
    assign layer5_outputs[3959] = 1'b0;
    assign layer5_outputs[3960] = ~(layer4_outputs[3701]) | (layer4_outputs[597]);
    assign layer5_outputs[3961] = (layer4_outputs[525]) ^ (layer4_outputs[3210]);
    assign layer5_outputs[3962] = (layer4_outputs[3949]) & (layer4_outputs[4282]);
    assign layer5_outputs[3963] = layer4_outputs[1723];
    assign layer5_outputs[3964] = (layer4_outputs[4053]) & (layer4_outputs[1313]);
    assign layer5_outputs[3965] = ~(layer4_outputs[5097]) | (layer4_outputs[4946]);
    assign layer5_outputs[3966] = layer4_outputs[2132];
    assign layer5_outputs[3967] = ~(layer4_outputs[179]);
    assign layer5_outputs[3968] = (layer4_outputs[2260]) ^ (layer4_outputs[3160]);
    assign layer5_outputs[3969] = ~((layer4_outputs[609]) ^ (layer4_outputs[383]));
    assign layer5_outputs[3970] = (layer4_outputs[3482]) ^ (layer4_outputs[4366]);
    assign layer5_outputs[3971] = 1'b1;
    assign layer5_outputs[3972] = ~((layer4_outputs[3099]) & (layer4_outputs[1892]));
    assign layer5_outputs[3973] = (layer4_outputs[2035]) ^ (layer4_outputs[142]);
    assign layer5_outputs[3974] = ~(layer4_outputs[2244]);
    assign layer5_outputs[3975] = 1'b0;
    assign layer5_outputs[3976] = ~((layer4_outputs[2462]) | (layer4_outputs[2995]));
    assign layer5_outputs[3977] = ~((layer4_outputs[559]) | (layer4_outputs[3536]));
    assign layer5_outputs[3978] = ~(layer4_outputs[4265]);
    assign layer5_outputs[3979] = ~(layer4_outputs[4070]);
    assign layer5_outputs[3980] = ~(layer4_outputs[3513]);
    assign layer5_outputs[3981] = ~(layer4_outputs[5041]);
    assign layer5_outputs[3982] = 1'b0;
    assign layer5_outputs[3983] = ~(layer4_outputs[666]);
    assign layer5_outputs[3984] = layer4_outputs[1513];
    assign layer5_outputs[3985] = 1'b0;
    assign layer5_outputs[3986] = ~(layer4_outputs[1192]);
    assign layer5_outputs[3987] = ~(layer4_outputs[497]);
    assign layer5_outputs[3988] = (layer4_outputs[2006]) & (layer4_outputs[3942]);
    assign layer5_outputs[3989] = ~(layer4_outputs[679]);
    assign layer5_outputs[3990] = layer4_outputs[592];
    assign layer5_outputs[3991] = (layer4_outputs[1151]) & ~(layer4_outputs[1706]);
    assign layer5_outputs[3992] = ~(layer4_outputs[2312]);
    assign layer5_outputs[3993] = layer4_outputs[2870];
    assign layer5_outputs[3994] = layer4_outputs[730];
    assign layer5_outputs[3995] = layer4_outputs[3924];
    assign layer5_outputs[3996] = ~((layer4_outputs[566]) & (layer4_outputs[1719]));
    assign layer5_outputs[3997] = (layer4_outputs[1281]) & ~(layer4_outputs[2098]);
    assign layer5_outputs[3998] = ~(layer4_outputs[772]);
    assign layer5_outputs[3999] = layer4_outputs[2417];
    assign layer5_outputs[4000] = layer4_outputs[3699];
    assign layer5_outputs[4001] = ~(layer4_outputs[4516]) | (layer4_outputs[2953]);
    assign layer5_outputs[4002] = ~((layer4_outputs[1435]) ^ (layer4_outputs[456]));
    assign layer5_outputs[4003] = ~(layer4_outputs[3472]);
    assign layer5_outputs[4004] = ~((layer4_outputs[1104]) & (layer4_outputs[150]));
    assign layer5_outputs[4005] = layer4_outputs[1689];
    assign layer5_outputs[4006] = ~(layer4_outputs[3408]);
    assign layer5_outputs[4007] = 1'b1;
    assign layer5_outputs[4008] = layer4_outputs[1445];
    assign layer5_outputs[4009] = ~((layer4_outputs[2999]) | (layer4_outputs[4234]));
    assign layer5_outputs[4010] = ~(layer4_outputs[4014]);
    assign layer5_outputs[4011] = (layer4_outputs[1035]) & ~(layer4_outputs[2807]);
    assign layer5_outputs[4012] = ~(layer4_outputs[4507]) | (layer4_outputs[704]);
    assign layer5_outputs[4013] = ~((layer4_outputs[1520]) | (layer4_outputs[4830]));
    assign layer5_outputs[4014] = ~((layer4_outputs[115]) ^ (layer4_outputs[3237]));
    assign layer5_outputs[4015] = (layer4_outputs[1438]) | (layer4_outputs[2002]);
    assign layer5_outputs[4016] = (layer4_outputs[1290]) & (layer4_outputs[3745]);
    assign layer5_outputs[4017] = layer4_outputs[1679];
    assign layer5_outputs[4018] = ~((layer4_outputs[4881]) & (layer4_outputs[3812]));
    assign layer5_outputs[4019] = ~(layer4_outputs[2804]);
    assign layer5_outputs[4020] = ~((layer4_outputs[998]) | (layer4_outputs[4416]));
    assign layer5_outputs[4021] = ~(layer4_outputs[3268]);
    assign layer5_outputs[4022] = ~((layer4_outputs[205]) ^ (layer4_outputs[2821]));
    assign layer5_outputs[4023] = layer4_outputs[838];
    assign layer5_outputs[4024] = layer4_outputs[4765];
    assign layer5_outputs[4025] = ~((layer4_outputs[3769]) | (layer4_outputs[1857]));
    assign layer5_outputs[4026] = layer4_outputs[2991];
    assign layer5_outputs[4027] = ~(layer4_outputs[4436]);
    assign layer5_outputs[4028] = layer4_outputs[4615];
    assign layer5_outputs[4029] = (layer4_outputs[2017]) ^ (layer4_outputs[3591]);
    assign layer5_outputs[4030] = ~((layer4_outputs[5044]) & (layer4_outputs[3445]));
    assign layer5_outputs[4031] = (layer4_outputs[511]) | (layer4_outputs[3044]);
    assign layer5_outputs[4032] = ~(layer4_outputs[1855]);
    assign layer5_outputs[4033] = (layer4_outputs[975]) & ~(layer4_outputs[3888]);
    assign layer5_outputs[4034] = layer4_outputs[3483];
    assign layer5_outputs[4035] = (layer4_outputs[706]) | (layer4_outputs[1462]);
    assign layer5_outputs[4036] = (layer4_outputs[2319]) | (layer4_outputs[1412]);
    assign layer5_outputs[4037] = layer4_outputs[2910];
    assign layer5_outputs[4038] = (layer4_outputs[1285]) & (layer4_outputs[2078]);
    assign layer5_outputs[4039] = (layer4_outputs[2812]) ^ (layer4_outputs[2229]);
    assign layer5_outputs[4040] = layer4_outputs[3378];
    assign layer5_outputs[4041] = (layer4_outputs[2552]) | (layer4_outputs[887]);
    assign layer5_outputs[4042] = ~(layer4_outputs[3530]);
    assign layer5_outputs[4043] = ~(layer4_outputs[233]);
    assign layer5_outputs[4044] = layer4_outputs[409];
    assign layer5_outputs[4045] = ~((layer4_outputs[4684]) ^ (layer4_outputs[4248]));
    assign layer5_outputs[4046] = ~((layer4_outputs[3790]) & (layer4_outputs[3231]));
    assign layer5_outputs[4047] = layer4_outputs[1141];
    assign layer5_outputs[4048] = ~(layer4_outputs[4515]);
    assign layer5_outputs[4049] = ~(layer4_outputs[4340]);
    assign layer5_outputs[4050] = layer4_outputs[4246];
    assign layer5_outputs[4051] = (layer4_outputs[1112]) & ~(layer4_outputs[3032]);
    assign layer5_outputs[4052] = (layer4_outputs[2170]) | (layer4_outputs[2449]);
    assign layer5_outputs[4053] = ~(layer4_outputs[1604]) | (layer4_outputs[2562]);
    assign layer5_outputs[4054] = 1'b0;
    assign layer5_outputs[4055] = ~((layer4_outputs[3543]) ^ (layer4_outputs[546]));
    assign layer5_outputs[4056] = layer4_outputs[718];
    assign layer5_outputs[4057] = (layer4_outputs[3163]) | (layer4_outputs[2829]);
    assign layer5_outputs[4058] = (layer4_outputs[677]) & (layer4_outputs[4789]);
    assign layer5_outputs[4059] = ~(layer4_outputs[3198]);
    assign layer5_outputs[4060] = (layer4_outputs[4063]) ^ (layer4_outputs[71]);
    assign layer5_outputs[4061] = (layer4_outputs[4048]) & ~(layer4_outputs[3085]);
    assign layer5_outputs[4062] = ~(layer4_outputs[945]);
    assign layer5_outputs[4063] = ~((layer4_outputs[4201]) & (layer4_outputs[4528]));
    assign layer5_outputs[4064] = ~(layer4_outputs[1376]);
    assign layer5_outputs[4065] = layer4_outputs[4059];
    assign layer5_outputs[4066] = ~(layer4_outputs[1964]);
    assign layer5_outputs[4067] = (layer4_outputs[708]) & ~(layer4_outputs[4953]);
    assign layer5_outputs[4068] = ~(layer4_outputs[918]);
    assign layer5_outputs[4069] = layer4_outputs[2707];
    assign layer5_outputs[4070] = (layer4_outputs[3774]) & ~(layer4_outputs[925]);
    assign layer5_outputs[4071] = (layer4_outputs[3404]) | (layer4_outputs[2790]);
    assign layer5_outputs[4072] = (layer4_outputs[504]) ^ (layer4_outputs[190]);
    assign layer5_outputs[4073] = ~(layer4_outputs[4133]);
    assign layer5_outputs[4074] = (layer4_outputs[4330]) & ~(layer4_outputs[4051]);
    assign layer5_outputs[4075] = ~(layer4_outputs[2485]);
    assign layer5_outputs[4076] = ~((layer4_outputs[1959]) & (layer4_outputs[2537]));
    assign layer5_outputs[4077] = layer4_outputs[4316];
    assign layer5_outputs[4078] = ~(layer4_outputs[1639]);
    assign layer5_outputs[4079] = layer4_outputs[3217];
    assign layer5_outputs[4080] = layer4_outputs[2199];
    assign layer5_outputs[4081] = ~(layer4_outputs[4565]) | (layer4_outputs[3576]);
    assign layer5_outputs[4082] = layer4_outputs[2859];
    assign layer5_outputs[4083] = ~((layer4_outputs[1201]) | (layer4_outputs[3939]));
    assign layer5_outputs[4084] = ~(layer4_outputs[3382]);
    assign layer5_outputs[4085] = ~(layer4_outputs[2067]);
    assign layer5_outputs[4086] = layer4_outputs[3158];
    assign layer5_outputs[4087] = ~(layer4_outputs[3340]);
    assign layer5_outputs[4088] = ~((layer4_outputs[3544]) | (layer4_outputs[5102]));
    assign layer5_outputs[4089] = ~((layer4_outputs[4918]) | (layer4_outputs[3041]));
    assign layer5_outputs[4090] = ~(layer4_outputs[4970]);
    assign layer5_outputs[4091] = (layer4_outputs[3949]) | (layer4_outputs[3965]);
    assign layer5_outputs[4092] = (layer4_outputs[2018]) ^ (layer4_outputs[3552]);
    assign layer5_outputs[4093] = layer4_outputs[2476];
    assign layer5_outputs[4094] = layer4_outputs[258];
    assign layer5_outputs[4095] = (layer4_outputs[2487]) | (layer4_outputs[4165]);
    assign layer5_outputs[4096] = (layer4_outputs[3740]) & ~(layer4_outputs[4641]);
    assign layer5_outputs[4097] = layer4_outputs[2992];
    assign layer5_outputs[4098] = ~(layer4_outputs[4204]);
    assign layer5_outputs[4099] = (layer4_outputs[4556]) & ~(layer4_outputs[5070]);
    assign layer5_outputs[4100] = (layer4_outputs[240]) & ~(layer4_outputs[972]);
    assign layer5_outputs[4101] = (layer4_outputs[3286]) & (layer4_outputs[1800]);
    assign layer5_outputs[4102] = (layer4_outputs[4550]) ^ (layer4_outputs[2222]);
    assign layer5_outputs[4103] = 1'b0;
    assign layer5_outputs[4104] = 1'b0;
    assign layer5_outputs[4105] = (layer4_outputs[2824]) ^ (layer4_outputs[2372]);
    assign layer5_outputs[4106] = ~((layer4_outputs[3187]) ^ (layer4_outputs[3467]));
    assign layer5_outputs[4107] = layer4_outputs[2810];
    assign layer5_outputs[4108] = ~((layer4_outputs[1377]) ^ (layer4_outputs[738]));
    assign layer5_outputs[4109] = ~((layer4_outputs[3974]) ^ (layer4_outputs[428]));
    assign layer5_outputs[4110] = ~(layer4_outputs[2055]);
    assign layer5_outputs[4111] = (layer4_outputs[4187]) & ~(layer4_outputs[1570]);
    assign layer5_outputs[4112] = ~(layer4_outputs[640]) | (layer4_outputs[3367]);
    assign layer5_outputs[4113] = layer4_outputs[4615];
    assign layer5_outputs[4114] = (layer4_outputs[2866]) ^ (layer4_outputs[1491]);
    assign layer5_outputs[4115] = ~(layer4_outputs[4046]) | (layer4_outputs[616]);
    assign layer5_outputs[4116] = (layer4_outputs[1239]) | (layer4_outputs[3751]);
    assign layer5_outputs[4117] = layer4_outputs[4429];
    assign layer5_outputs[4118] = layer4_outputs[472];
    assign layer5_outputs[4119] = ~((layer4_outputs[2695]) ^ (layer4_outputs[1204]));
    assign layer5_outputs[4120] = layer4_outputs[4347];
    assign layer5_outputs[4121] = (layer4_outputs[4378]) ^ (layer4_outputs[1267]);
    assign layer5_outputs[4122] = layer4_outputs[2528];
    assign layer5_outputs[4123] = (layer4_outputs[4804]) & ~(layer4_outputs[4757]);
    assign layer5_outputs[4124] = ~((layer4_outputs[451]) | (layer4_outputs[4949]));
    assign layer5_outputs[4125] = layer4_outputs[4394];
    assign layer5_outputs[4126] = ~((layer4_outputs[2650]) & (layer4_outputs[4745]));
    assign layer5_outputs[4127] = (layer4_outputs[4793]) ^ (layer4_outputs[521]);
    assign layer5_outputs[4128] = (layer4_outputs[1816]) & ~(layer4_outputs[209]);
    assign layer5_outputs[4129] = layer4_outputs[802];
    assign layer5_outputs[4130] = ~(layer4_outputs[135]);
    assign layer5_outputs[4131] = ~(layer4_outputs[1717]);
    assign layer5_outputs[4132] = ~((layer4_outputs[876]) ^ (layer4_outputs[782]));
    assign layer5_outputs[4133] = layer4_outputs[2685];
    assign layer5_outputs[4134] = (layer4_outputs[3576]) ^ (layer4_outputs[1074]);
    assign layer5_outputs[4135] = ~(layer4_outputs[2102]) | (layer4_outputs[3204]);
    assign layer5_outputs[4136] = 1'b1;
    assign layer5_outputs[4137] = ~((layer4_outputs[1973]) ^ (layer4_outputs[786]));
    assign layer5_outputs[4138] = layer4_outputs[1538];
    assign layer5_outputs[4139] = layer4_outputs[4808];
    assign layer5_outputs[4140] = ~(layer4_outputs[2295]);
    assign layer5_outputs[4141] = layer4_outputs[583];
    assign layer5_outputs[4142] = layer4_outputs[1265];
    assign layer5_outputs[4143] = layer4_outputs[1768];
    assign layer5_outputs[4144] = ~((layer4_outputs[483]) & (layer4_outputs[106]));
    assign layer5_outputs[4145] = ~(layer4_outputs[1992]);
    assign layer5_outputs[4146] = ~(layer4_outputs[3223]);
    assign layer5_outputs[4147] = ~(layer4_outputs[3217]);
    assign layer5_outputs[4148] = layer4_outputs[991];
    assign layer5_outputs[4149] = 1'b1;
    assign layer5_outputs[4150] = ~(layer4_outputs[3845]) | (layer4_outputs[840]);
    assign layer5_outputs[4151] = (layer4_outputs[498]) | (layer4_outputs[1097]);
    assign layer5_outputs[4152] = ~(layer4_outputs[2139]);
    assign layer5_outputs[4153] = ~(layer4_outputs[1699]);
    assign layer5_outputs[4154] = ~((layer4_outputs[2898]) ^ (layer4_outputs[3655]));
    assign layer5_outputs[4155] = ~((layer4_outputs[1531]) & (layer4_outputs[614]));
    assign layer5_outputs[4156] = ~(layer4_outputs[4656]) | (layer4_outputs[2590]);
    assign layer5_outputs[4157] = ~((layer4_outputs[2197]) & (layer4_outputs[141]));
    assign layer5_outputs[4158] = layer4_outputs[4943];
    assign layer5_outputs[4159] = layer4_outputs[618];
    assign layer5_outputs[4160] = ~(layer4_outputs[2247]);
    assign layer5_outputs[4161] = (layer4_outputs[1888]) ^ (layer4_outputs[191]);
    assign layer5_outputs[4162] = ~(layer4_outputs[708]);
    assign layer5_outputs[4163] = 1'b0;
    assign layer5_outputs[4164] = ~(layer4_outputs[4253]);
    assign layer5_outputs[4165] = (layer4_outputs[2093]) ^ (layer4_outputs[1548]);
    assign layer5_outputs[4166] = ~(layer4_outputs[2535]);
    assign layer5_outputs[4167] = layer4_outputs[615];
    assign layer5_outputs[4168] = ~(layer4_outputs[3188]);
    assign layer5_outputs[4169] = ~((layer4_outputs[3393]) & (layer4_outputs[1362]));
    assign layer5_outputs[4170] = 1'b0;
    assign layer5_outputs[4171] = (layer4_outputs[2149]) & (layer4_outputs[2089]);
    assign layer5_outputs[4172] = ~(layer4_outputs[2624]);
    assign layer5_outputs[4173] = ~(layer4_outputs[1117]) | (layer4_outputs[3114]);
    assign layer5_outputs[4174] = (layer4_outputs[3155]) | (layer4_outputs[811]);
    assign layer5_outputs[4175] = ~(layer4_outputs[1359]) | (layer4_outputs[4073]);
    assign layer5_outputs[4176] = (layer4_outputs[4665]) & ~(layer4_outputs[2519]);
    assign layer5_outputs[4177] = layer4_outputs[3283];
    assign layer5_outputs[4178] = (layer4_outputs[2572]) & (layer4_outputs[892]);
    assign layer5_outputs[4179] = (layer4_outputs[1092]) & ~(layer4_outputs[508]);
    assign layer5_outputs[4180] = ~(layer4_outputs[1203]);
    assign layer5_outputs[4181] = layer4_outputs[4079];
    assign layer5_outputs[4182] = 1'b1;
    assign layer5_outputs[4183] = ~(layer4_outputs[1625]);
    assign layer5_outputs[4184] = ~(layer4_outputs[1445]);
    assign layer5_outputs[4185] = layer4_outputs[4220];
    assign layer5_outputs[4186] = layer4_outputs[3867];
    assign layer5_outputs[4187] = layer4_outputs[2467];
    assign layer5_outputs[4188] = layer4_outputs[933];
    assign layer5_outputs[4189] = (layer4_outputs[1496]) ^ (layer4_outputs[522]);
    assign layer5_outputs[4190] = ~((layer4_outputs[3175]) & (layer4_outputs[2461]));
    assign layer5_outputs[4191] = (layer4_outputs[1054]) | (layer4_outputs[4737]);
    assign layer5_outputs[4192] = ~(layer4_outputs[817]);
    assign layer5_outputs[4193] = ~(layer4_outputs[4495]);
    assign layer5_outputs[4194] = layer4_outputs[2018];
    assign layer5_outputs[4195] = ~(layer4_outputs[4525]);
    assign layer5_outputs[4196] = layer4_outputs[1509];
    assign layer5_outputs[4197] = ~((layer4_outputs[4833]) ^ (layer4_outputs[4546]));
    assign layer5_outputs[4198] = layer4_outputs[1072];
    assign layer5_outputs[4199] = ~((layer4_outputs[590]) | (layer4_outputs[4205]));
    assign layer5_outputs[4200] = ~((layer4_outputs[3713]) & (layer4_outputs[3009]));
    assign layer5_outputs[4201] = layer4_outputs[363];
    assign layer5_outputs[4202] = ~(layer4_outputs[4147]);
    assign layer5_outputs[4203] = ~((layer4_outputs[337]) | (layer4_outputs[596]));
    assign layer5_outputs[4204] = ~((layer4_outputs[90]) & (layer4_outputs[2860]));
    assign layer5_outputs[4205] = ~(layer4_outputs[3454]);
    assign layer5_outputs[4206] = layer4_outputs[1567];
    assign layer5_outputs[4207] = ~(layer4_outputs[1456]);
    assign layer5_outputs[4208] = ~(layer4_outputs[107]);
    assign layer5_outputs[4209] = (layer4_outputs[3485]) ^ (layer4_outputs[2867]);
    assign layer5_outputs[4210] = layer4_outputs[2962];
    assign layer5_outputs[4211] = (layer4_outputs[3974]) & ~(layer4_outputs[4538]);
    assign layer5_outputs[4212] = layer4_outputs[3250];
    assign layer5_outputs[4213] = layer4_outputs[5016];
    assign layer5_outputs[4214] = ~((layer4_outputs[1752]) & (layer4_outputs[4568]));
    assign layer5_outputs[4215] = ~(layer4_outputs[495]);
    assign layer5_outputs[4216] = ~(layer4_outputs[2904]);
    assign layer5_outputs[4217] = layer4_outputs[1846];
    assign layer5_outputs[4218] = ~(layer4_outputs[3029]);
    assign layer5_outputs[4219] = ~(layer4_outputs[2797]) | (layer4_outputs[454]);
    assign layer5_outputs[4220] = ~(layer4_outputs[1757]);
    assign layer5_outputs[4221] = layer4_outputs[4128];
    assign layer5_outputs[4222] = ~(layer4_outputs[33]);
    assign layer5_outputs[4223] = layer4_outputs[4246];
    assign layer5_outputs[4224] = (layer4_outputs[809]) ^ (layer4_outputs[625]);
    assign layer5_outputs[4225] = (layer4_outputs[4106]) ^ (layer4_outputs[1984]);
    assign layer5_outputs[4226] = layer4_outputs[2912];
    assign layer5_outputs[4227] = ~(layer4_outputs[1323]) | (layer4_outputs[4652]);
    assign layer5_outputs[4228] = ~(layer4_outputs[3526]) | (layer4_outputs[123]);
    assign layer5_outputs[4229] = (layer4_outputs[1]) & (layer4_outputs[4160]);
    assign layer5_outputs[4230] = ~((layer4_outputs[2423]) ^ (layer4_outputs[2818]));
    assign layer5_outputs[4231] = ~((layer4_outputs[1607]) ^ (layer4_outputs[4249]));
    assign layer5_outputs[4232] = layer4_outputs[2434];
    assign layer5_outputs[4233] = ~(layer4_outputs[2055]);
    assign layer5_outputs[4234] = (layer4_outputs[3500]) & ~(layer4_outputs[3183]);
    assign layer5_outputs[4235] = layer4_outputs[3649];
    assign layer5_outputs[4236] = layer4_outputs[2960];
    assign layer5_outputs[4237] = ~(layer4_outputs[2732]);
    assign layer5_outputs[4238] = ~(layer4_outputs[1516]);
    assign layer5_outputs[4239] = 1'b0;
    assign layer5_outputs[4240] = (layer4_outputs[520]) & ~(layer4_outputs[1001]);
    assign layer5_outputs[4241] = layer4_outputs[107];
    assign layer5_outputs[4242] = ~(layer4_outputs[1413]);
    assign layer5_outputs[4243] = ~(layer4_outputs[4793]);
    assign layer5_outputs[4244] = (layer4_outputs[2307]) & (layer4_outputs[4511]);
    assign layer5_outputs[4245] = layer4_outputs[4786];
    assign layer5_outputs[4246] = ~((layer4_outputs[27]) | (layer4_outputs[948]));
    assign layer5_outputs[4247] = ~(layer4_outputs[1600]);
    assign layer5_outputs[4248] = layer4_outputs[2678];
    assign layer5_outputs[4249] = (layer4_outputs[3873]) | (layer4_outputs[2274]);
    assign layer5_outputs[4250] = ~(layer4_outputs[2645]);
    assign layer5_outputs[4251] = ~(layer4_outputs[1850]);
    assign layer5_outputs[4252] = ~((layer4_outputs[769]) & (layer4_outputs[1910]));
    assign layer5_outputs[4253] = layer4_outputs[1443];
    assign layer5_outputs[4254] = layer4_outputs[3426];
    assign layer5_outputs[4255] = layer4_outputs[1796];
    assign layer5_outputs[4256] = ~((layer4_outputs[2505]) ^ (layer4_outputs[3528]));
    assign layer5_outputs[4257] = ~(layer4_outputs[3432]);
    assign layer5_outputs[4258] = layer4_outputs[2942];
    assign layer5_outputs[4259] = ~(layer4_outputs[1896]);
    assign layer5_outputs[4260] = (layer4_outputs[328]) ^ (layer4_outputs[1682]);
    assign layer5_outputs[4261] = layer4_outputs[3710];
    assign layer5_outputs[4262] = 1'b1;
    assign layer5_outputs[4263] = ~(layer4_outputs[3040]) | (layer4_outputs[4108]);
    assign layer5_outputs[4264] = ~((layer4_outputs[2370]) | (layer4_outputs[101]));
    assign layer5_outputs[4265] = (layer4_outputs[4127]) | (layer4_outputs[1836]);
    assign layer5_outputs[4266] = (layer4_outputs[278]) ^ (layer4_outputs[4596]);
    assign layer5_outputs[4267] = ~(layer4_outputs[298]);
    assign layer5_outputs[4268] = layer4_outputs[3257];
    assign layer5_outputs[4269] = (layer4_outputs[3024]) & ~(layer4_outputs[1294]);
    assign layer5_outputs[4270] = 1'b1;
    assign layer5_outputs[4271] = layer4_outputs[342];
    assign layer5_outputs[4272] = layer4_outputs[3609];
    assign layer5_outputs[4273] = (layer4_outputs[3733]) & ~(layer4_outputs[2996]);
    assign layer5_outputs[4274] = 1'b1;
    assign layer5_outputs[4275] = (layer4_outputs[3754]) & ~(layer4_outputs[4326]);
    assign layer5_outputs[4276] = ~((layer4_outputs[3681]) & (layer4_outputs[4207]));
    assign layer5_outputs[4277] = ~((layer4_outputs[4160]) & (layer4_outputs[2305]));
    assign layer5_outputs[4278] = ~((layer4_outputs[4667]) & (layer4_outputs[1739]));
    assign layer5_outputs[4279] = ~(layer4_outputs[631]);
    assign layer5_outputs[4280] = (layer4_outputs[368]) & ~(layer4_outputs[1678]);
    assign layer5_outputs[4281] = (layer4_outputs[4135]) & ~(layer4_outputs[438]);
    assign layer5_outputs[4282] = layer4_outputs[2117];
    assign layer5_outputs[4283] = ~(layer4_outputs[3522]) | (layer4_outputs[3794]);
    assign layer5_outputs[4284] = ~((layer4_outputs[4043]) & (layer4_outputs[1260]));
    assign layer5_outputs[4285] = ~(layer4_outputs[1566]);
    assign layer5_outputs[4286] = ~(layer4_outputs[2630]) | (layer4_outputs[4301]);
    assign layer5_outputs[4287] = (layer4_outputs[3447]) ^ (layer4_outputs[4231]);
    assign layer5_outputs[4288] = 1'b1;
    assign layer5_outputs[4289] = (layer4_outputs[4132]) ^ (layer4_outputs[4422]);
    assign layer5_outputs[4290] = layer4_outputs[581];
    assign layer5_outputs[4291] = ~(layer4_outputs[514]);
    assign layer5_outputs[4292] = ~(layer4_outputs[2005]) | (layer4_outputs[2062]);
    assign layer5_outputs[4293] = ~(layer4_outputs[3957]) | (layer4_outputs[918]);
    assign layer5_outputs[4294] = (layer4_outputs[1844]) | (layer4_outputs[2521]);
    assign layer5_outputs[4295] = 1'b1;
    assign layer5_outputs[4296] = 1'b1;
    assign layer5_outputs[4297] = (layer4_outputs[5036]) | (layer4_outputs[4982]);
    assign layer5_outputs[4298] = layer4_outputs[3498];
    assign layer5_outputs[4299] = layer4_outputs[636];
    assign layer5_outputs[4300] = ~(layer4_outputs[3531]);
    assign layer5_outputs[4301] = ~(layer4_outputs[3042]) | (layer4_outputs[1323]);
    assign layer5_outputs[4302] = layer4_outputs[857];
    assign layer5_outputs[4303] = (layer4_outputs[399]) & ~(layer4_outputs[4981]);
    assign layer5_outputs[4304] = (layer4_outputs[2649]) ^ (layer4_outputs[139]);
    assign layer5_outputs[4305] = layer4_outputs[701];
    assign layer5_outputs[4306] = ~(layer4_outputs[31]);
    assign layer5_outputs[4307] = ~(layer4_outputs[3709]);
    assign layer5_outputs[4308] = (layer4_outputs[1124]) | (layer4_outputs[1685]);
    assign layer5_outputs[4309] = ~(layer4_outputs[5034]);
    assign layer5_outputs[4310] = ~((layer4_outputs[3828]) ^ (layer4_outputs[537]));
    assign layer5_outputs[4311] = (layer4_outputs[726]) & ~(layer4_outputs[4905]);
    assign layer5_outputs[4312] = (layer4_outputs[3870]) | (layer4_outputs[2730]);
    assign layer5_outputs[4313] = layer4_outputs[3395];
    assign layer5_outputs[4314] = (layer4_outputs[3680]) ^ (layer4_outputs[863]);
    assign layer5_outputs[4315] = ~(layer4_outputs[2947]);
    assign layer5_outputs[4316] = layer4_outputs[3255];
    assign layer5_outputs[4317] = ~(layer4_outputs[2356]) | (layer4_outputs[4803]);
    assign layer5_outputs[4318] = layer4_outputs[1809];
    assign layer5_outputs[4319] = ~((layer4_outputs[2725]) ^ (layer4_outputs[4563]));
    assign layer5_outputs[4320] = ~((layer4_outputs[2053]) | (layer4_outputs[2332]));
    assign layer5_outputs[4321] = ~((layer4_outputs[4733]) & (layer4_outputs[4875]));
    assign layer5_outputs[4322] = 1'b1;
    assign layer5_outputs[4323] = layer4_outputs[3784];
    assign layer5_outputs[4324] = ~(layer4_outputs[588]);
    assign layer5_outputs[4325] = ~((layer4_outputs[659]) ^ (layer4_outputs[5100]));
    assign layer5_outputs[4326] = ~(layer4_outputs[1473]);
    assign layer5_outputs[4327] = ~(layer4_outputs[4791]) | (layer4_outputs[5051]);
    assign layer5_outputs[4328] = layer4_outputs[4813];
    assign layer5_outputs[4329] = ~((layer4_outputs[657]) & (layer4_outputs[4854]));
    assign layer5_outputs[4330] = (layer4_outputs[2865]) & ~(layer4_outputs[4775]);
    assign layer5_outputs[4331] = layer4_outputs[2651];
    assign layer5_outputs[4332] = ~((layer4_outputs[1510]) | (layer4_outputs[4561]));
    assign layer5_outputs[4333] = ~((layer4_outputs[2499]) | (layer4_outputs[2021]));
    assign layer5_outputs[4334] = ~(layer4_outputs[4254]) | (layer4_outputs[1120]);
    assign layer5_outputs[4335] = (layer4_outputs[3898]) ^ (layer4_outputs[2914]);
    assign layer5_outputs[4336] = ~(layer4_outputs[1135]);
    assign layer5_outputs[4337] = ~((layer4_outputs[1790]) & (layer4_outputs[4809]));
    assign layer5_outputs[4338] = ~(layer4_outputs[2087]) | (layer4_outputs[1830]);
    assign layer5_outputs[4339] = ~(layer4_outputs[1871]) | (layer4_outputs[2506]);
    assign layer5_outputs[4340] = ~(layer4_outputs[4542]);
    assign layer5_outputs[4341] = ~((layer4_outputs[1707]) | (layer4_outputs[3055]));
    assign layer5_outputs[4342] = ~(layer4_outputs[3739]) | (layer4_outputs[4219]);
    assign layer5_outputs[4343] = (layer4_outputs[4907]) ^ (layer4_outputs[3548]);
    assign layer5_outputs[4344] = ~((layer4_outputs[443]) | (layer4_outputs[827]));
    assign layer5_outputs[4345] = (layer4_outputs[510]) & ~(layer4_outputs[120]);
    assign layer5_outputs[4346] = ~((layer4_outputs[4992]) ^ (layer4_outputs[116]));
    assign layer5_outputs[4347] = layer4_outputs[3846];
    assign layer5_outputs[4348] = layer4_outputs[4082];
    assign layer5_outputs[4349] = ~((layer4_outputs[4259]) ^ (layer4_outputs[3189]));
    assign layer5_outputs[4350] = layer4_outputs[2451];
    assign layer5_outputs[4351] = ~(layer4_outputs[3550]) | (layer4_outputs[60]);
    assign layer5_outputs[4352] = 1'b0;
    assign layer5_outputs[4353] = ~(layer4_outputs[949]);
    assign layer5_outputs[4354] = (layer4_outputs[1887]) | (layer4_outputs[1272]);
    assign layer5_outputs[4355] = (layer4_outputs[5006]) & (layer4_outputs[4137]);
    assign layer5_outputs[4356] = ~((layer4_outputs[2955]) | (layer4_outputs[2851]));
    assign layer5_outputs[4357] = ~(layer4_outputs[1896]) | (layer4_outputs[292]);
    assign layer5_outputs[4358] = layer4_outputs[1023];
    assign layer5_outputs[4359] = (layer4_outputs[920]) ^ (layer4_outputs[2643]);
    assign layer5_outputs[4360] = layer4_outputs[3923];
    assign layer5_outputs[4361] = (layer4_outputs[3125]) | (layer4_outputs[5092]);
    assign layer5_outputs[4362] = ~((layer4_outputs[773]) | (layer4_outputs[2392]));
    assign layer5_outputs[4363] = (layer4_outputs[1902]) | (layer4_outputs[3440]);
    assign layer5_outputs[4364] = layer4_outputs[198];
    assign layer5_outputs[4365] = (layer4_outputs[3236]) ^ (layer4_outputs[3440]);
    assign layer5_outputs[4366] = ~(layer4_outputs[742]) | (layer4_outputs[43]);
    assign layer5_outputs[4367] = layer4_outputs[3992];
    assign layer5_outputs[4368] = layer4_outputs[4674];
    assign layer5_outputs[4369] = ~(layer4_outputs[1140]);
    assign layer5_outputs[4370] = layer4_outputs[4197];
    assign layer5_outputs[4371] = (layer4_outputs[2304]) & ~(layer4_outputs[2017]);
    assign layer5_outputs[4372] = (layer4_outputs[4477]) & (layer4_outputs[1573]);
    assign layer5_outputs[4373] = layer4_outputs[5059];
    assign layer5_outputs[4374] = 1'b1;
    assign layer5_outputs[4375] = ~(layer4_outputs[1079]);
    assign layer5_outputs[4376] = ~((layer4_outputs[829]) & (layer4_outputs[4599]));
    assign layer5_outputs[4377] = ~(layer4_outputs[3952]);
    assign layer5_outputs[4378] = ~(layer4_outputs[679]) | (layer4_outputs[1610]);
    assign layer5_outputs[4379] = ~(layer4_outputs[2552]);
    assign layer5_outputs[4380] = ~((layer4_outputs[4442]) ^ (layer4_outputs[1526]));
    assign layer5_outputs[4381] = 1'b1;
    assign layer5_outputs[4382] = layer4_outputs[2261];
    assign layer5_outputs[4383] = ~(layer4_outputs[464]);
    assign layer5_outputs[4384] = layer4_outputs[678];
    assign layer5_outputs[4385] = (layer4_outputs[4110]) & (layer4_outputs[2292]);
    assign layer5_outputs[4386] = ~(layer4_outputs[698]);
    assign layer5_outputs[4387] = 1'b1;
    assign layer5_outputs[4388] = ~(layer4_outputs[3887]);
    assign layer5_outputs[4389] = layer4_outputs[4167];
    assign layer5_outputs[4390] = layer4_outputs[1990];
    assign layer5_outputs[4391] = (layer4_outputs[4714]) & (layer4_outputs[2900]);
    assign layer5_outputs[4392] = layer4_outputs[3858];
    assign layer5_outputs[4393] = (layer4_outputs[213]) | (layer4_outputs[65]);
    assign layer5_outputs[4394] = (layer4_outputs[3461]) & (layer4_outputs[4051]);
    assign layer5_outputs[4395] = ~(layer4_outputs[3031]);
    assign layer5_outputs[4396] = ~((layer4_outputs[654]) ^ (layer4_outputs[2054]));
    assign layer5_outputs[4397] = ~(layer4_outputs[4914]);
    assign layer5_outputs[4398] = 1'b1;
    assign layer5_outputs[4399] = (layer4_outputs[2374]) & (layer4_outputs[1981]);
    assign layer5_outputs[4400] = ~(layer4_outputs[4913]) | (layer4_outputs[3981]);
    assign layer5_outputs[4401] = ~(layer4_outputs[4961]);
    assign layer5_outputs[4402] = ~((layer4_outputs[2033]) & (layer4_outputs[4649]));
    assign layer5_outputs[4403] = layer4_outputs[1901];
    assign layer5_outputs[4404] = ~(layer4_outputs[4111]) | (layer4_outputs[3607]);
    assign layer5_outputs[4405] = ~(layer4_outputs[3345]);
    assign layer5_outputs[4406] = ~(layer4_outputs[3583]) | (layer4_outputs[1947]);
    assign layer5_outputs[4407] = layer4_outputs[1369];
    assign layer5_outputs[4408] = (layer4_outputs[1862]) & ~(layer4_outputs[2271]);
    assign layer5_outputs[4409] = ~(layer4_outputs[2584]);
    assign layer5_outputs[4410] = (layer4_outputs[2919]) & ~(layer4_outputs[3851]);
    assign layer5_outputs[4411] = layer4_outputs[4835];
    assign layer5_outputs[4412] = ~((layer4_outputs[3463]) ^ (layer4_outputs[1945]));
    assign layer5_outputs[4413] = (layer4_outputs[2842]) & ~(layer4_outputs[2184]);
    assign layer5_outputs[4414] = 1'b0;
    assign layer5_outputs[4415] = (layer4_outputs[2941]) & ~(layer4_outputs[2001]);
    assign layer5_outputs[4416] = layer4_outputs[1090];
    assign layer5_outputs[4417] = ~((layer4_outputs[3622]) & (layer4_outputs[5053]));
    assign layer5_outputs[4418] = (layer4_outputs[2334]) & ~(layer4_outputs[3547]);
    assign layer5_outputs[4419] = ~(layer4_outputs[2274]);
    assign layer5_outputs[4420] = layer4_outputs[3620];
    assign layer5_outputs[4421] = 1'b0;
    assign layer5_outputs[4422] = layer4_outputs[4089];
    assign layer5_outputs[4423] = (layer4_outputs[4481]) & ~(layer4_outputs[4105]);
    assign layer5_outputs[4424] = (layer4_outputs[723]) & ~(layer4_outputs[2608]);
    assign layer5_outputs[4425] = ~(layer4_outputs[1286]);
    assign layer5_outputs[4426] = (layer4_outputs[1223]) | (layer4_outputs[1829]);
    assign layer5_outputs[4427] = ~((layer4_outputs[466]) & (layer4_outputs[2042]));
    assign layer5_outputs[4428] = (layer4_outputs[267]) | (layer4_outputs[277]);
    assign layer5_outputs[4429] = ~(layer4_outputs[4694]) | (layer4_outputs[3915]);
    assign layer5_outputs[4430] = layer4_outputs[256];
    assign layer5_outputs[4431] = ~(layer4_outputs[2216]) | (layer4_outputs[32]);
    assign layer5_outputs[4432] = ~((layer4_outputs[4831]) & (layer4_outputs[3748]));
    assign layer5_outputs[4433] = layer4_outputs[1111];
    assign layer5_outputs[4434] = ~((layer4_outputs[338]) | (layer4_outputs[2689]));
    assign layer5_outputs[4435] = ~(layer4_outputs[3238]);
    assign layer5_outputs[4436] = ~((layer4_outputs[896]) ^ (layer4_outputs[798]));
    assign layer5_outputs[4437] = (layer4_outputs[3324]) | (layer4_outputs[255]);
    assign layer5_outputs[4438] = ~(layer4_outputs[3233]);
    assign layer5_outputs[4439] = ~(layer4_outputs[2603]);
    assign layer5_outputs[4440] = ~(layer4_outputs[792]);
    assign layer5_outputs[4441] = (layer4_outputs[2972]) & ~(layer4_outputs[817]);
    assign layer5_outputs[4442] = layer4_outputs[4792];
    assign layer5_outputs[4443] = 1'b1;
    assign layer5_outputs[4444] = ~((layer4_outputs[4535]) | (layer4_outputs[2750]));
    assign layer5_outputs[4445] = ~(layer4_outputs[3416]);
    assign layer5_outputs[4446] = ~(layer4_outputs[3897]);
    assign layer5_outputs[4447] = (layer4_outputs[2456]) & (layer4_outputs[773]);
    assign layer5_outputs[4448] = ~((layer4_outputs[304]) ^ (layer4_outputs[293]));
    assign layer5_outputs[4449] = ~((layer4_outputs[2245]) & (layer4_outputs[4434]));
    assign layer5_outputs[4450] = layer4_outputs[3307];
    assign layer5_outputs[4451] = ~(layer4_outputs[3728]);
    assign layer5_outputs[4452] = (layer4_outputs[2261]) & (layer4_outputs[1530]);
    assign layer5_outputs[4453] = ~(layer4_outputs[3114]) | (layer4_outputs[3073]);
    assign layer5_outputs[4454] = ~(layer4_outputs[779]) | (layer4_outputs[575]);
    assign layer5_outputs[4455] = ~((layer4_outputs[4108]) ^ (layer4_outputs[3607]));
    assign layer5_outputs[4456] = (layer4_outputs[3967]) & (layer4_outputs[4863]);
    assign layer5_outputs[4457] = ~(layer4_outputs[3556]);
    assign layer5_outputs[4458] = ~(layer4_outputs[2152]) | (layer4_outputs[2370]);
    assign layer5_outputs[4459] = ~(layer4_outputs[15]);
    assign layer5_outputs[4460] = ~((layer4_outputs[4241]) | (layer4_outputs[1432]));
    assign layer5_outputs[4461] = 1'b1;
    assign layer5_outputs[4462] = ~((layer4_outputs[1320]) | (layer4_outputs[1985]));
    assign layer5_outputs[4463] = layer4_outputs[3672];
    assign layer5_outputs[4464] = ~((layer4_outputs[3207]) | (layer4_outputs[4148]));
    assign layer5_outputs[4465] = ~(layer4_outputs[2546]) | (layer4_outputs[4547]);
    assign layer5_outputs[4466] = ~(layer4_outputs[3308]);
    assign layer5_outputs[4467] = ~(layer4_outputs[1216]);
    assign layer5_outputs[4468] = ~(layer4_outputs[4157]);
    assign layer5_outputs[4469] = (layer4_outputs[4595]) & (layer4_outputs[4015]);
    assign layer5_outputs[4470] = layer4_outputs[1542];
    assign layer5_outputs[4471] = layer4_outputs[4335];
    assign layer5_outputs[4472] = (layer4_outputs[4050]) & ~(layer4_outputs[3359]);
    assign layer5_outputs[4473] = layer4_outputs[2569];
    assign layer5_outputs[4474] = (layer4_outputs[4876]) & ~(layer4_outputs[964]);
    assign layer5_outputs[4475] = ~((layer4_outputs[785]) & (layer4_outputs[2085]));
    assign layer5_outputs[4476] = 1'b1;
    assign layer5_outputs[4477] = ~((layer4_outputs[4178]) ^ (layer4_outputs[4133]));
    assign layer5_outputs[4478] = ~((layer4_outputs[4120]) & (layer4_outputs[1054]));
    assign layer5_outputs[4479] = ~(layer4_outputs[3818]) | (layer4_outputs[1569]);
    assign layer5_outputs[4480] = ~(layer4_outputs[3076]);
    assign layer5_outputs[4481] = layer4_outputs[1704];
    assign layer5_outputs[4482] = ~((layer4_outputs[2772]) ^ (layer4_outputs[2040]));
    assign layer5_outputs[4483] = ~((layer4_outputs[296]) ^ (layer4_outputs[3268]));
    assign layer5_outputs[4484] = ~(layer4_outputs[251]);
    assign layer5_outputs[4485] = (layer4_outputs[1303]) | (layer4_outputs[4610]);
    assign layer5_outputs[4486] = layer4_outputs[3465];
    assign layer5_outputs[4487] = (layer4_outputs[2285]) & ~(layer4_outputs[109]);
    assign layer5_outputs[4488] = layer4_outputs[4728];
    assign layer5_outputs[4489] = (layer4_outputs[4302]) ^ (layer4_outputs[3975]);
    assign layer5_outputs[4490] = ~(layer4_outputs[4690]) | (layer4_outputs[1848]);
    assign layer5_outputs[4491] = ~((layer4_outputs[4237]) ^ (layer4_outputs[2748]));
    assign layer5_outputs[4492] = (layer4_outputs[3840]) & ~(layer4_outputs[2174]);
    assign layer5_outputs[4493] = ~(layer4_outputs[4039]);
    assign layer5_outputs[4494] = ~(layer4_outputs[2976]);
    assign layer5_outputs[4495] = ~(layer4_outputs[1180]);
    assign layer5_outputs[4496] = (layer4_outputs[4023]) & (layer4_outputs[2147]);
    assign layer5_outputs[4497] = layer4_outputs[2757];
    assign layer5_outputs[4498] = ~((layer4_outputs[4725]) & (layer4_outputs[3429]));
    assign layer5_outputs[4499] = layer4_outputs[2493];
    assign layer5_outputs[4500] = 1'b0;
    assign layer5_outputs[4501] = ~(layer4_outputs[2427]);
    assign layer5_outputs[4502] = layer4_outputs[810];
    assign layer5_outputs[4503] = (layer4_outputs[4289]) & (layer4_outputs[4726]);
    assign layer5_outputs[4504] = ~((layer4_outputs[3026]) | (layer4_outputs[1586]));
    assign layer5_outputs[4505] = ~(layer4_outputs[1738]);
    assign layer5_outputs[4506] = ~(layer4_outputs[3251]);
    assign layer5_outputs[4507] = ~(layer4_outputs[896]);
    assign layer5_outputs[4508] = layer4_outputs[2455];
    assign layer5_outputs[4509] = (layer4_outputs[3458]) & (layer4_outputs[46]);
    assign layer5_outputs[4510] = ~(layer4_outputs[2354]);
    assign layer5_outputs[4511] = ~(layer4_outputs[2204]) | (layer4_outputs[1346]);
    assign layer5_outputs[4512] = ~((layer4_outputs[2961]) | (layer4_outputs[3439]));
    assign layer5_outputs[4513] = (layer4_outputs[2397]) & ~(layer4_outputs[2138]);
    assign layer5_outputs[4514] = ~(layer4_outputs[860]) | (layer4_outputs[574]);
    assign layer5_outputs[4515] = layer4_outputs[3519];
    assign layer5_outputs[4516] = ~(layer4_outputs[4502]);
    assign layer5_outputs[4517] = layer4_outputs[2687];
    assign layer5_outputs[4518] = layer4_outputs[4020];
    assign layer5_outputs[4519] = (layer4_outputs[2506]) & ~(layer4_outputs[4935]);
    assign layer5_outputs[4520] = ~(layer4_outputs[5026]) | (layer4_outputs[557]);
    assign layer5_outputs[4521] = layer4_outputs[1300];
    assign layer5_outputs[4522] = (layer4_outputs[2970]) & (layer4_outputs[2315]);
    assign layer5_outputs[4523] = layer4_outputs[3226];
    assign layer5_outputs[4524] = layer4_outputs[4816];
    assign layer5_outputs[4525] = ~(layer4_outputs[4161]);
    assign layer5_outputs[4526] = (layer4_outputs[2736]) | (layer4_outputs[5018]);
    assign layer5_outputs[4527] = layer4_outputs[4262];
    assign layer5_outputs[4528] = layer4_outputs[1826];
    assign layer5_outputs[4529] = layer4_outputs[1832];
    assign layer5_outputs[4530] = 1'b0;
    assign layer5_outputs[4531] = ~((layer4_outputs[0]) ^ (layer4_outputs[1870]));
    assign layer5_outputs[4532] = ~(layer4_outputs[2516]);
    assign layer5_outputs[4533] = 1'b1;
    assign layer5_outputs[4534] = ~(layer4_outputs[2384]);
    assign layer5_outputs[4535] = ~(layer4_outputs[1702]);
    assign layer5_outputs[4536] = ~(layer4_outputs[1218]) | (layer4_outputs[4029]);
    assign layer5_outputs[4537] = ~(layer4_outputs[4165]);
    assign layer5_outputs[4538] = ~((layer4_outputs[4954]) & (layer4_outputs[1946]));
    assign layer5_outputs[4539] = ~(layer4_outputs[1150]) | (layer4_outputs[4453]);
    assign layer5_outputs[4540] = layer4_outputs[4867];
    assign layer5_outputs[4541] = ~((layer4_outputs[1867]) ^ (layer4_outputs[2719]));
    assign layer5_outputs[4542] = layer4_outputs[494];
    assign layer5_outputs[4543] = layer4_outputs[2028];
    assign layer5_outputs[4544] = layer4_outputs[5081];
    assign layer5_outputs[4545] = layer4_outputs[2483];
    assign layer5_outputs[4546] = layer4_outputs[1985];
    assign layer5_outputs[4547] = layer4_outputs[4142];
    assign layer5_outputs[4548] = ~(layer4_outputs[2136]);
    assign layer5_outputs[4549] = layer4_outputs[3482];
    assign layer5_outputs[4550] = ~(layer4_outputs[865]);
    assign layer5_outputs[4551] = layer4_outputs[2598];
    assign layer5_outputs[4552] = ~((layer4_outputs[755]) & (layer4_outputs[2077]));
    assign layer5_outputs[4553] = layer4_outputs[28];
    assign layer5_outputs[4554] = ~((layer4_outputs[1334]) ^ (layer4_outputs[2097]));
    assign layer5_outputs[4555] = layer4_outputs[486];
    assign layer5_outputs[4556] = ~((layer4_outputs[534]) ^ (layer4_outputs[3861]));
    assign layer5_outputs[4557] = layer4_outputs[763];
    assign layer5_outputs[4558] = ~(layer4_outputs[2739]);
    assign layer5_outputs[4559] = ~(layer4_outputs[3322]) | (layer4_outputs[3320]);
    assign layer5_outputs[4560] = ~(layer4_outputs[3051]);
    assign layer5_outputs[4561] = (layer4_outputs[1498]) & ~(layer4_outputs[573]);
    assign layer5_outputs[4562] = (layer4_outputs[2439]) | (layer4_outputs[2697]);
    assign layer5_outputs[4563] = layer4_outputs[3206];
    assign layer5_outputs[4564] = ~(layer4_outputs[4988]);
    assign layer5_outputs[4565] = layer4_outputs[4993];
    assign layer5_outputs[4566] = ~(layer4_outputs[1604]) | (layer4_outputs[655]);
    assign layer5_outputs[4567] = ~(layer4_outputs[793]);
    assign layer5_outputs[4568] = (layer4_outputs[688]) | (layer4_outputs[741]);
    assign layer5_outputs[4569] = (layer4_outputs[4241]) & (layer4_outputs[3224]);
    assign layer5_outputs[4570] = (layer4_outputs[2049]) & (layer4_outputs[1071]);
    assign layer5_outputs[4571] = ~(layer4_outputs[2135]);
    assign layer5_outputs[4572] = ~(layer4_outputs[3372]);
    assign layer5_outputs[4573] = (layer4_outputs[4630]) & ~(layer4_outputs[2482]);
    assign layer5_outputs[4574] = ~(layer4_outputs[3664]);
    assign layer5_outputs[4575] = ~(layer4_outputs[94]);
    assign layer5_outputs[4576] = ~(layer4_outputs[1842]);
    assign layer5_outputs[4577] = (layer4_outputs[4738]) & (layer4_outputs[3334]);
    assign layer5_outputs[4578] = layer4_outputs[114];
    assign layer5_outputs[4579] = (layer4_outputs[954]) & ~(layer4_outputs[2724]);
    assign layer5_outputs[4580] = 1'b1;
    assign layer5_outputs[4581] = (layer4_outputs[3164]) | (layer4_outputs[2527]);
    assign layer5_outputs[4582] = ~(layer4_outputs[4803]);
    assign layer5_outputs[4583] = ~(layer4_outputs[5045]);
    assign layer5_outputs[4584] = ~(layer4_outputs[831]) | (layer4_outputs[1074]);
    assign layer5_outputs[4585] = layer4_outputs[4465];
    assign layer5_outputs[4586] = ~(layer4_outputs[4853]);
    assign layer5_outputs[4587] = layer4_outputs[2291];
    assign layer5_outputs[4588] = ~((layer4_outputs[2959]) ^ (layer4_outputs[2047]));
    assign layer5_outputs[4589] = (layer4_outputs[764]) & ~(layer4_outputs[3090]);
    assign layer5_outputs[4590] = 1'b0;
    assign layer5_outputs[4591] = (layer4_outputs[3690]) & ~(layer4_outputs[343]);
    assign layer5_outputs[4592] = (layer4_outputs[599]) & ~(layer4_outputs[1139]);
    assign layer5_outputs[4593] = (layer4_outputs[3776]) & ~(layer4_outputs[1426]);
    assign layer5_outputs[4594] = ~(layer4_outputs[4325]);
    assign layer5_outputs[4595] = ~((layer4_outputs[498]) & (layer4_outputs[3393]));
    assign layer5_outputs[4596] = ~(layer4_outputs[3651]);
    assign layer5_outputs[4597] = (layer4_outputs[1971]) & ~(layer4_outputs[3132]);
    assign layer5_outputs[4598] = ~((layer4_outputs[1220]) ^ (layer4_outputs[2447]));
    assign layer5_outputs[4599] = (layer4_outputs[2711]) | (layer4_outputs[2463]);
    assign layer5_outputs[4600] = ~(layer4_outputs[197]);
    assign layer5_outputs[4601] = ~(layer4_outputs[3248]);
    assign layer5_outputs[4602] = (layer4_outputs[2201]) & ~(layer4_outputs[780]);
    assign layer5_outputs[4603] = ~(layer4_outputs[445]);
    assign layer5_outputs[4604] = ~(layer4_outputs[4665]) | (layer4_outputs[344]);
    assign layer5_outputs[4605] = ~((layer4_outputs[4616]) | (layer4_outputs[2179]));
    assign layer5_outputs[4606] = (layer4_outputs[4607]) & (layer4_outputs[1699]);
    assign layer5_outputs[4607] = ~((layer4_outputs[449]) | (layer4_outputs[4722]));
    assign layer5_outputs[4608] = layer4_outputs[995];
    assign layer5_outputs[4609] = layer4_outputs[3935];
    assign layer5_outputs[4610] = ~(layer4_outputs[2526]);
    assign layer5_outputs[4611] = (layer4_outputs[3271]) & (layer4_outputs[1629]);
    assign layer5_outputs[4612] = ~(layer4_outputs[2986]);
    assign layer5_outputs[4613] = layer4_outputs[3988];
    assign layer5_outputs[4614] = (layer4_outputs[4281]) & ~(layer4_outputs[682]);
    assign layer5_outputs[4615] = (layer4_outputs[3656]) ^ (layer4_outputs[1387]);
    assign layer5_outputs[4616] = ~(layer4_outputs[4668]);
    assign layer5_outputs[4617] = (layer4_outputs[1397]) & ~(layer4_outputs[4471]);
    assign layer5_outputs[4618] = ~((layer4_outputs[1013]) & (layer4_outputs[639]));
    assign layer5_outputs[4619] = ~(layer4_outputs[2732]);
    assign layer5_outputs[4620] = 1'b0;
    assign layer5_outputs[4621] = layer4_outputs[1849];
    assign layer5_outputs[4622] = ~(layer4_outputs[3771]);
    assign layer5_outputs[4623] = layer4_outputs[2582];
    assign layer5_outputs[4624] = (layer4_outputs[4569]) & (layer4_outputs[1663]);
    assign layer5_outputs[4625] = ~(layer4_outputs[152]);
    assign layer5_outputs[4626] = (layer4_outputs[1693]) & ~(layer4_outputs[3667]);
    assign layer5_outputs[4627] = (layer4_outputs[1162]) ^ (layer4_outputs[5027]);
    assign layer5_outputs[4628] = (layer4_outputs[4407]) & ~(layer4_outputs[3784]);
    assign layer5_outputs[4629] = ~(layer4_outputs[1343]);
    assign layer5_outputs[4630] = ~(layer4_outputs[2842]);
    assign layer5_outputs[4631] = ~(layer4_outputs[24]);
    assign layer5_outputs[4632] = ~((layer4_outputs[1153]) ^ (layer4_outputs[3033]));
    assign layer5_outputs[4633] = (layer4_outputs[4645]) ^ (layer4_outputs[1795]);
    assign layer5_outputs[4634] = ~(layer4_outputs[3638]) | (layer4_outputs[1425]);
    assign layer5_outputs[4635] = ~((layer4_outputs[1641]) | (layer4_outputs[945]));
    assign layer5_outputs[4636] = ~(layer4_outputs[4218]);
    assign layer5_outputs[4637] = (layer4_outputs[1018]) & ~(layer4_outputs[4605]);
    assign layer5_outputs[4638] = layer4_outputs[4957];
    assign layer5_outputs[4639] = (layer4_outputs[2241]) ^ (layer4_outputs[3668]);
    assign layer5_outputs[4640] = ~(layer4_outputs[1857]) | (layer4_outputs[3859]);
    assign layer5_outputs[4641] = ~(layer4_outputs[890]);
    assign layer5_outputs[4642] = ~(layer4_outputs[527]) | (layer4_outputs[3125]);
    assign layer5_outputs[4643] = ~(layer4_outputs[3052]);
    assign layer5_outputs[4644] = ~(layer4_outputs[4563]) | (layer4_outputs[4993]);
    assign layer5_outputs[4645] = ~((layer4_outputs[239]) ^ (layer4_outputs[4508]));
    assign layer5_outputs[4646] = ~(layer4_outputs[193]);
    assign layer5_outputs[4647] = ~(layer4_outputs[3367]);
    assign layer5_outputs[4648] = layer4_outputs[1156];
    assign layer5_outputs[4649] = ~(layer4_outputs[1838]);
    assign layer5_outputs[4650] = (layer4_outputs[400]) ^ (layer4_outputs[2921]);
    assign layer5_outputs[4651] = ~((layer4_outputs[2696]) & (layer4_outputs[4895]));
    assign layer5_outputs[4652] = (layer4_outputs[4419]) | (layer4_outputs[827]);
    assign layer5_outputs[4653] = (layer4_outputs[2316]) & ~(layer4_outputs[1999]);
    assign layer5_outputs[4654] = layer4_outputs[1855];
    assign layer5_outputs[4655] = ~(layer4_outputs[1808]) | (layer4_outputs[4416]);
    assign layer5_outputs[4656] = ~(layer4_outputs[430]);
    assign layer5_outputs[4657] = layer4_outputs[3803];
    assign layer5_outputs[4658] = 1'b0;
    assign layer5_outputs[4659] = layer4_outputs[3385];
    assign layer5_outputs[4660] = (layer4_outputs[3327]) ^ (layer4_outputs[2014]);
    assign layer5_outputs[4661] = ~((layer4_outputs[87]) | (layer4_outputs[1060]));
    assign layer5_outputs[4662] = 1'b0;
    assign layer5_outputs[4663] = ~(layer4_outputs[4502]);
    assign layer5_outputs[4664] = ~(layer4_outputs[2208]);
    assign layer5_outputs[4665] = (layer4_outputs[2927]) & (layer4_outputs[2746]);
    assign layer5_outputs[4666] = (layer4_outputs[1116]) & ~(layer4_outputs[2627]);
    assign layer5_outputs[4667] = ~(layer4_outputs[4293]);
    assign layer5_outputs[4668] = ~(layer4_outputs[4762]);
    assign layer5_outputs[4669] = ~(layer4_outputs[4848]);
    assign layer5_outputs[4670] = ~(layer4_outputs[1103]);
    assign layer5_outputs[4671] = ~(layer4_outputs[5117]) | (layer4_outputs[4293]);
    assign layer5_outputs[4672] = (layer4_outputs[3871]) & ~(layer4_outputs[2911]);
    assign layer5_outputs[4673] = ~((layer4_outputs[57]) | (layer4_outputs[4383]));
    assign layer5_outputs[4674] = (layer4_outputs[2289]) & (layer4_outputs[3392]);
    assign layer5_outputs[4675] = ~(layer4_outputs[642]) | (layer4_outputs[963]);
    assign layer5_outputs[4676] = ~(layer4_outputs[3193]);
    assign layer5_outputs[4677] = ~(layer4_outputs[3521]);
    assign layer5_outputs[4678] = (layer4_outputs[547]) & (layer4_outputs[5097]);
    assign layer5_outputs[4679] = ~(layer4_outputs[2142]);
    assign layer5_outputs[4680] = ~((layer4_outputs[4558]) ^ (layer4_outputs[1783]));
    assign layer5_outputs[4681] = ~(layer4_outputs[2789]);
    assign layer5_outputs[4682] = layer4_outputs[706];
    assign layer5_outputs[4683] = (layer4_outputs[1118]) | (layer4_outputs[3035]);
    assign layer5_outputs[4684] = (layer4_outputs[5066]) & ~(layer4_outputs[4216]);
    assign layer5_outputs[4685] = ~((layer4_outputs[1636]) ^ (layer4_outputs[4677]));
    assign layer5_outputs[4686] = ~(layer4_outputs[1025]);
    assign layer5_outputs[4687] = layer4_outputs[629];
    assign layer5_outputs[4688] = layer4_outputs[3823];
    assign layer5_outputs[4689] = ~(layer4_outputs[3593]);
    assign layer5_outputs[4690] = ~((layer4_outputs[2211]) & (layer4_outputs[3666]));
    assign layer5_outputs[4691] = ~((layer4_outputs[1233]) | (layer4_outputs[2099]));
    assign layer5_outputs[4692] = layer4_outputs[3980];
    assign layer5_outputs[4693] = ~(layer4_outputs[4324]);
    assign layer5_outputs[4694] = ~((layer4_outputs[2024]) | (layer4_outputs[2472]));
    assign layer5_outputs[4695] = ~(layer4_outputs[1773]);
    assign layer5_outputs[4696] = ~((layer4_outputs[143]) & (layer4_outputs[2063]));
    assign layer5_outputs[4697] = ~((layer4_outputs[2691]) & (layer4_outputs[3108]));
    assign layer5_outputs[4698] = (layer4_outputs[2183]) & ~(layer4_outputs[2907]);
    assign layer5_outputs[4699] = (layer4_outputs[4643]) & ~(layer4_outputs[3941]);
    assign layer5_outputs[4700] = ~(layer4_outputs[1107]) | (layer4_outputs[4650]);
    assign layer5_outputs[4701] = layer4_outputs[1993];
    assign layer5_outputs[4702] = (layer4_outputs[4295]) & ~(layer4_outputs[1303]);
    assign layer5_outputs[4703] = layer4_outputs[4272];
    assign layer5_outputs[4704] = layer4_outputs[2097];
    assign layer5_outputs[4705] = ~(layer4_outputs[2072]);
    assign layer5_outputs[4706] = layer4_outputs[3747];
    assign layer5_outputs[4707] = (layer4_outputs[168]) | (layer4_outputs[3419]);
    assign layer5_outputs[4708] = (layer4_outputs[1525]) | (layer4_outputs[2640]);
    assign layer5_outputs[4709] = 1'b0;
    assign layer5_outputs[4710] = 1'b0;
    assign layer5_outputs[4711] = ~(layer4_outputs[2744]) | (layer4_outputs[4181]);
    assign layer5_outputs[4712] = 1'b0;
    assign layer5_outputs[4713] = ~(layer4_outputs[4692]) | (layer4_outputs[2966]);
    assign layer5_outputs[4714] = ~(layer4_outputs[1465]);
    assign layer5_outputs[4715] = (layer4_outputs[2094]) & ~(layer4_outputs[3991]);
    assign layer5_outputs[4716] = (layer4_outputs[4431]) & (layer4_outputs[1751]);
    assign layer5_outputs[4717] = 1'b0;
    assign layer5_outputs[4718] = ~((layer4_outputs[3042]) ^ (layer4_outputs[1219]));
    assign layer5_outputs[4719] = layer4_outputs[3318];
    assign layer5_outputs[4720] = (layer4_outputs[4371]) ^ (layer4_outputs[381]);
    assign layer5_outputs[4721] = ~(layer4_outputs[3822]);
    assign layer5_outputs[4722] = ~(layer4_outputs[3256]);
    assign layer5_outputs[4723] = (layer4_outputs[882]) | (layer4_outputs[3227]);
    assign layer5_outputs[4724] = ~((layer4_outputs[2344]) & (layer4_outputs[2620]));
    assign layer5_outputs[4725] = (layer4_outputs[8]) | (layer4_outputs[868]);
    assign layer5_outputs[4726] = layer4_outputs[4085];
    assign layer5_outputs[4727] = ~((layer4_outputs[2250]) | (layer4_outputs[4117]));
    assign layer5_outputs[4728] = ~((layer4_outputs[4159]) & (layer4_outputs[1612]));
    assign layer5_outputs[4729] = layer4_outputs[4930];
    assign layer5_outputs[4730] = 1'b1;
    assign layer5_outputs[4731] = ~(layer4_outputs[2773]);
    assign layer5_outputs[4732] = (layer4_outputs[1585]) | (layer4_outputs[4368]);
    assign layer5_outputs[4733] = ~(layer4_outputs[1222]) | (layer4_outputs[3436]);
    assign layer5_outputs[4734] = 1'b0;
    assign layer5_outputs[4735] = (layer4_outputs[946]) ^ (layer4_outputs[1050]);
    assign layer5_outputs[4736] = (layer4_outputs[609]) & ~(layer4_outputs[4214]);
    assign layer5_outputs[4737] = ~(layer4_outputs[4978]) | (layer4_outputs[2792]);
    assign layer5_outputs[4738] = ~((layer4_outputs[4587]) | (layer4_outputs[4342]));
    assign layer5_outputs[4739] = ~(layer4_outputs[2647]) | (layer4_outputs[364]);
    assign layer5_outputs[4740] = ~((layer4_outputs[4349]) | (layer4_outputs[3665]));
    assign layer5_outputs[4741] = 1'b1;
    assign layer5_outputs[4742] = layer4_outputs[3683];
    assign layer5_outputs[4743] = (layer4_outputs[2190]) ^ (layer4_outputs[3449]);
    assign layer5_outputs[4744] = layer4_outputs[4780];
    assign layer5_outputs[4745] = ~(layer4_outputs[1599]);
    assign layer5_outputs[4746] = ~(layer4_outputs[3815]);
    assign layer5_outputs[4747] = ~((layer4_outputs[610]) ^ (layer4_outputs[1937]));
    assign layer5_outputs[4748] = layer4_outputs[4821];
    assign layer5_outputs[4749] = ~((layer4_outputs[1691]) ^ (layer4_outputs[1257]));
    assign layer5_outputs[4750] = (layer4_outputs[394]) | (layer4_outputs[4801]);
    assign layer5_outputs[4751] = layer4_outputs[2038];
    assign layer5_outputs[4752] = layer4_outputs[3429];
    assign layer5_outputs[4753] = (layer4_outputs[4379]) & ~(layer4_outputs[1821]);
    assign layer5_outputs[4754] = ~(layer4_outputs[3328]);
    assign layer5_outputs[4755] = ~((layer4_outputs[454]) ^ (layer4_outputs[1688]));
    assign layer5_outputs[4756] = layer4_outputs[2175];
    assign layer5_outputs[4757] = ~(layer4_outputs[290]);
    assign layer5_outputs[4758] = ~(layer4_outputs[2015]);
    assign layer5_outputs[4759] = (layer4_outputs[3633]) ^ (layer4_outputs[2150]);
    assign layer5_outputs[4760] = layer4_outputs[2633];
    assign layer5_outputs[4761] = ~((layer4_outputs[2739]) & (layer4_outputs[632]));
    assign layer5_outputs[4762] = ~(layer4_outputs[5054]);
    assign layer5_outputs[4763] = layer4_outputs[3053];
    assign layer5_outputs[4764] = layer4_outputs[148];
    assign layer5_outputs[4765] = layer4_outputs[371];
    assign layer5_outputs[4766] = layer4_outputs[1255];
    assign layer5_outputs[4767] = (layer4_outputs[1466]) & ~(layer4_outputs[994]);
    assign layer5_outputs[4768] = (layer4_outputs[457]) & ~(layer4_outputs[1881]);
    assign layer5_outputs[4769] = (layer4_outputs[1596]) & (layer4_outputs[2514]);
    assign layer5_outputs[4770] = ~(layer4_outputs[1093]) | (layer4_outputs[3720]);
    assign layer5_outputs[4771] = ~((layer4_outputs[4103]) | (layer4_outputs[94]));
    assign layer5_outputs[4772] = ~(layer4_outputs[3537]);
    assign layer5_outputs[4773] = layer4_outputs[3737];
    assign layer5_outputs[4774] = ~(layer4_outputs[1045]);
    assign layer5_outputs[4775] = ~(layer4_outputs[1293]) | (layer4_outputs[3824]);
    assign layer5_outputs[4776] = (layer4_outputs[4962]) | (layer4_outputs[381]);
    assign layer5_outputs[4777] = 1'b0;
    assign layer5_outputs[4778] = 1'b0;
    assign layer5_outputs[4779] = ~(layer4_outputs[2708]);
    assign layer5_outputs[4780] = (layer4_outputs[354]) & (layer4_outputs[4086]);
    assign layer5_outputs[4781] = (layer4_outputs[1297]) ^ (layer4_outputs[3660]);
    assign layer5_outputs[4782] = layer4_outputs[1990];
    assign layer5_outputs[4783] = ~(layer4_outputs[3475]);
    assign layer5_outputs[4784] = ~(layer4_outputs[3008]);
    assign layer5_outputs[4785] = ~(layer4_outputs[2252]) | (layer4_outputs[2052]);
    assign layer5_outputs[4786] = (layer4_outputs[2705]) | (layer4_outputs[3778]);
    assign layer5_outputs[4787] = 1'b0;
    assign layer5_outputs[4788] = (layer4_outputs[1331]) & ~(layer4_outputs[450]);
    assign layer5_outputs[4789] = layer4_outputs[2264];
    assign layer5_outputs[4790] = layer4_outputs[2357];
    assign layer5_outputs[4791] = ~(layer4_outputs[4177]);
    assign layer5_outputs[4792] = (layer4_outputs[3299]) & ~(layer4_outputs[1154]);
    assign layer5_outputs[4793] = layer4_outputs[2200];
    assign layer5_outputs[4794] = layer4_outputs[772];
    assign layer5_outputs[4795] = layer4_outputs[5068];
    assign layer5_outputs[4796] = ~(layer4_outputs[790]);
    assign layer5_outputs[4797] = layer4_outputs[3006];
    assign layer5_outputs[4798] = ~(layer4_outputs[3692]);
    assign layer5_outputs[4799] = ~(layer4_outputs[3126]);
    assign layer5_outputs[4800] = ~(layer4_outputs[2303]);
    assign layer5_outputs[4801] = ~(layer4_outputs[48]);
    assign layer5_outputs[4802] = (layer4_outputs[2560]) | (layer4_outputs[3418]);
    assign layer5_outputs[4803] = ~((layer4_outputs[1976]) & (layer4_outputs[3483]));
    assign layer5_outputs[4804] = (layer4_outputs[2684]) & ~(layer4_outputs[2336]);
    assign layer5_outputs[4805] = (layer4_outputs[610]) & ~(layer4_outputs[2075]);
    assign layer5_outputs[4806] = 1'b0;
    assign layer5_outputs[4807] = ~(layer4_outputs[4024]);
    assign layer5_outputs[4808] = ~(layer4_outputs[21]);
    assign layer5_outputs[4809] = ~(layer4_outputs[707]) | (layer4_outputs[2642]);
    assign layer5_outputs[4810] = (layer4_outputs[768]) | (layer4_outputs[2474]);
    assign layer5_outputs[4811] = ~(layer4_outputs[552]);
    assign layer5_outputs[4812] = ~(layer4_outputs[4988]);
    assign layer5_outputs[4813] = ~(layer4_outputs[2765]) | (layer4_outputs[1870]);
    assign layer5_outputs[4814] = layer4_outputs[2360];
    assign layer5_outputs[4815] = layer4_outputs[4848];
    assign layer5_outputs[4816] = ~(layer4_outputs[3916]);
    assign layer5_outputs[4817] = (layer4_outputs[4963]) & ~(layer4_outputs[2709]);
    assign layer5_outputs[4818] = 1'b0;
    assign layer5_outputs[4819] = ~(layer4_outputs[254]);
    assign layer5_outputs[4820] = ~(layer4_outputs[4648]);
    assign layer5_outputs[4821] = (layer4_outputs[3935]) | (layer4_outputs[2938]);
    assign layer5_outputs[4822] = ~((layer4_outputs[420]) | (layer4_outputs[2378]));
    assign layer5_outputs[4823] = 1'b0;
    assign layer5_outputs[4824] = layer4_outputs[4240];
    assign layer5_outputs[4825] = ~(layer4_outputs[3905]);
    assign layer5_outputs[4826] = ~(layer4_outputs[1170]);
    assign layer5_outputs[4827] = layer4_outputs[4843];
    assign layer5_outputs[4828] = ~((layer4_outputs[2210]) ^ (layer4_outputs[2122]));
    assign layer5_outputs[4829] = ~(layer4_outputs[2756]) | (layer4_outputs[2401]);
    assign layer5_outputs[4830] = ~(layer4_outputs[2202]);
    assign layer5_outputs[4831] = (layer4_outputs[619]) & ~(layer4_outputs[4671]);
    assign layer5_outputs[4832] = ~(layer4_outputs[2654]) | (layer4_outputs[3128]);
    assign layer5_outputs[4833] = ~(layer4_outputs[3674]);
    assign layer5_outputs[4834] = (layer4_outputs[2804]) & ~(layer4_outputs[1711]);
    assign layer5_outputs[4835] = layer4_outputs[2521];
    assign layer5_outputs[4836] = (layer4_outputs[3514]) & ~(layer4_outputs[5094]);
    assign layer5_outputs[4837] = ~((layer4_outputs[1056]) | (layer4_outputs[4104]));
    assign layer5_outputs[4838] = layer4_outputs[3148];
    assign layer5_outputs[4839] = layer4_outputs[4352];
    assign layer5_outputs[4840] = (layer4_outputs[3596]) & (layer4_outputs[388]);
    assign layer5_outputs[4841] = ~(layer4_outputs[2298]) | (layer4_outputs[5046]);
    assign layer5_outputs[4842] = (layer4_outputs[3932]) ^ (layer4_outputs[4186]);
    assign layer5_outputs[4843] = ~(layer4_outputs[4683]) | (layer4_outputs[1751]);
    assign layer5_outputs[4844] = ~(layer4_outputs[4539]);
    assign layer5_outputs[4845] = layer4_outputs[2673];
    assign layer5_outputs[4846] = layer4_outputs[2590];
    assign layer5_outputs[4847] = ~(layer4_outputs[1934]);
    assign layer5_outputs[4848] = ~(layer4_outputs[4980]);
    assign layer5_outputs[4849] = (layer4_outputs[4967]) & ~(layer4_outputs[2886]);
    assign layer5_outputs[4850] = ~(layer4_outputs[4158]) | (layer4_outputs[4396]);
    assign layer5_outputs[4851] = ~(layer4_outputs[2868]);
    assign layer5_outputs[4852] = ~(layer4_outputs[3025]);
    assign layer5_outputs[4853] = ~(layer4_outputs[4309]) | (layer4_outputs[4590]);
    assign layer5_outputs[4854] = ~(layer4_outputs[2074]);
    assign layer5_outputs[4855] = ~(layer4_outputs[270]);
    assign layer5_outputs[4856] = ~(layer4_outputs[1709]);
    assign layer5_outputs[4857] = layer4_outputs[358];
    assign layer5_outputs[4858] = ~(layer4_outputs[3969]);
    assign layer5_outputs[4859] = ~(layer4_outputs[2448]) | (layer4_outputs[3876]);
    assign layer5_outputs[4860] = layer4_outputs[2782];
    assign layer5_outputs[4861] = ~((layer4_outputs[1125]) & (layer4_outputs[4626]));
    assign layer5_outputs[4862] = ~(layer4_outputs[3433]) | (layer4_outputs[3930]);
    assign layer5_outputs[4863] = ~((layer4_outputs[4357]) | (layer4_outputs[4977]));
    assign layer5_outputs[4864] = ~(layer4_outputs[729]) | (layer4_outputs[1048]);
    assign layer5_outputs[4865] = ~(layer4_outputs[3896]);
    assign layer5_outputs[4866] = (layer4_outputs[3597]) ^ (layer4_outputs[2738]);
    assign layer5_outputs[4867] = ~(layer4_outputs[4586]);
    assign layer5_outputs[4868] = layer4_outputs[3885];
    assign layer5_outputs[4869] = (layer4_outputs[1536]) & (layer4_outputs[270]);
    assign layer5_outputs[4870] = (layer4_outputs[244]) | (layer4_outputs[244]);
    assign layer5_outputs[4871] = (layer4_outputs[3906]) & ~(layer4_outputs[1169]);
    assign layer5_outputs[4872] = ~(layer4_outputs[2877]);
    assign layer5_outputs[4873] = (layer4_outputs[5048]) | (layer4_outputs[3249]);
    assign layer5_outputs[4874] = ~(layer4_outputs[3968]);
    assign layer5_outputs[4875] = layer4_outputs[3726];
    assign layer5_outputs[4876] = layer4_outputs[2184];
    assign layer5_outputs[4877] = ~(layer4_outputs[1764]);
    assign layer5_outputs[4878] = (layer4_outputs[202]) & ~(layer4_outputs[2446]);
    assign layer5_outputs[4879] = ~(layer4_outputs[3694]);
    assign layer5_outputs[4880] = layer4_outputs[2069];
    assign layer5_outputs[4881] = (layer4_outputs[2838]) & ~(layer4_outputs[3572]);
    assign layer5_outputs[4882] = ~((layer4_outputs[1391]) | (layer4_outputs[3384]));
    assign layer5_outputs[4883] = ~((layer4_outputs[350]) & (layer4_outputs[4426]));
    assign layer5_outputs[4884] = layer4_outputs[845];
    assign layer5_outputs[4885] = layer4_outputs[2897];
    assign layer5_outputs[4886] = ~((layer4_outputs[1275]) & (layer4_outputs[2318]));
    assign layer5_outputs[4887] = ~(layer4_outputs[627]) | (layer4_outputs[4682]);
    assign layer5_outputs[4888] = layer4_outputs[410];
    assign layer5_outputs[4889] = ~((layer4_outputs[5111]) ^ (layer4_outputs[526]));
    assign layer5_outputs[4890] = ~(layer4_outputs[986]) | (layer4_outputs[4009]);
    assign layer5_outputs[4891] = ~((layer4_outputs[3462]) & (layer4_outputs[481]));
    assign layer5_outputs[4892] = (layer4_outputs[346]) | (layer4_outputs[4391]);
    assign layer5_outputs[4893] = ~(layer4_outputs[1819]);
    assign layer5_outputs[4894] = (layer4_outputs[4671]) & (layer4_outputs[686]);
    assign layer5_outputs[4895] = ~((layer4_outputs[330]) | (layer4_outputs[1352]));
    assign layer5_outputs[4896] = layer4_outputs[2743];
    assign layer5_outputs[4897] = ~((layer4_outputs[1344]) & (layer4_outputs[3464]));
    assign layer5_outputs[4898] = ~(layer4_outputs[4261]) | (layer4_outputs[1843]);
    assign layer5_outputs[4899] = ~(layer4_outputs[3816]);
    assign layer5_outputs[4900] = 1'b0;
    assign layer5_outputs[4901] = (layer4_outputs[2653]) ^ (layer4_outputs[3203]);
    assign layer5_outputs[4902] = ~(layer4_outputs[3434]);
    assign layer5_outputs[4903] = ~(layer4_outputs[1316]);
    assign layer5_outputs[4904] = ~(layer4_outputs[1311]);
    assign layer5_outputs[4905] = layer4_outputs[1265];
    assign layer5_outputs[4906] = layer4_outputs[134];
    assign layer5_outputs[4907] = ~(layer4_outputs[1634]);
    assign layer5_outputs[4908] = ~((layer4_outputs[1550]) | (layer4_outputs[3627]));
    assign layer5_outputs[4909] = layer4_outputs[1616];
    assign layer5_outputs[4910] = (layer4_outputs[267]) & ~(layer4_outputs[1123]);
    assign layer5_outputs[4911] = ~(layer4_outputs[4069]);
    assign layer5_outputs[4912] = ~((layer4_outputs[3788]) ^ (layer4_outputs[1861]));
    assign layer5_outputs[4913] = layer4_outputs[3166];
    assign layer5_outputs[4914] = (layer4_outputs[3341]) | (layer4_outputs[4100]);
    assign layer5_outputs[4915] = (layer4_outputs[2933]) ^ (layer4_outputs[2140]);
    assign layer5_outputs[4916] = (layer4_outputs[4524]) & (layer4_outputs[4791]);
    assign layer5_outputs[4917] = ~(layer4_outputs[4610]);
    assign layer5_outputs[4918] = (layer4_outputs[2575]) | (layer4_outputs[1676]);
    assign layer5_outputs[4919] = ~((layer4_outputs[5017]) & (layer4_outputs[3816]));
    assign layer5_outputs[4920] = (layer4_outputs[2667]) & (layer4_outputs[154]);
    assign layer5_outputs[4921] = ~(layer4_outputs[4770]);
    assign layer5_outputs[4922] = layer4_outputs[2495];
    assign layer5_outputs[4923] = ~((layer4_outputs[2825]) ^ (layer4_outputs[462]));
    assign layer5_outputs[4924] = layer4_outputs[3905];
    assign layer5_outputs[4925] = ~(layer4_outputs[512]) | (layer4_outputs[3153]);
    assign layer5_outputs[4926] = layer4_outputs[2713];
    assign layer5_outputs[4927] = layer4_outputs[916];
    assign layer5_outputs[4928] = (layer4_outputs[176]) ^ (layer4_outputs[2731]);
    assign layer5_outputs[4929] = layer4_outputs[2181];
    assign layer5_outputs[4930] = 1'b0;
    assign layer5_outputs[4931] = ~(layer4_outputs[4096]);
    assign layer5_outputs[4932] = (layer4_outputs[3612]) & ~(layer4_outputs[4663]);
    assign layer5_outputs[4933] = ~(layer4_outputs[3276]) | (layer4_outputs[3659]);
    assign layer5_outputs[4934] = ~(layer4_outputs[4229]) | (layer4_outputs[1786]);
    assign layer5_outputs[4935] = ~(layer4_outputs[888]) | (layer4_outputs[4617]);
    assign layer5_outputs[4936] = (layer4_outputs[3297]) & ~(layer4_outputs[4402]);
    assign layer5_outputs[4937] = ~(layer4_outputs[1529]);
    assign layer5_outputs[4938] = (layer4_outputs[4275]) ^ (layer4_outputs[3383]);
    assign layer5_outputs[4939] = ~((layer4_outputs[472]) | (layer4_outputs[3109]));
    assign layer5_outputs[4940] = ~(layer4_outputs[250]);
    assign layer5_outputs[4941] = layer4_outputs[823];
    assign layer5_outputs[4942] = layer4_outputs[2937];
    assign layer5_outputs[4943] = layer4_outputs[1588];
    assign layer5_outputs[4944] = ~(layer4_outputs[3581]);
    assign layer5_outputs[4945] = layer4_outputs[4162];
    assign layer5_outputs[4946] = (layer4_outputs[4842]) & (layer4_outputs[201]);
    assign layer5_outputs[4947] = (layer4_outputs[3214]) ^ (layer4_outputs[1772]);
    assign layer5_outputs[4948] = ~(layer4_outputs[2565]);
    assign layer5_outputs[4949] = ~(layer4_outputs[1879]) | (layer4_outputs[3606]);
    assign layer5_outputs[4950] = (layer4_outputs[1830]) & ~(layer4_outputs[3535]);
    assign layer5_outputs[4951] = ~((layer4_outputs[2618]) | (layer4_outputs[651]));
    assign layer5_outputs[4952] = layer4_outputs[4024];
    assign layer5_outputs[4953] = ~(layer4_outputs[1286]) | (layer4_outputs[3454]);
    assign layer5_outputs[4954] = (layer4_outputs[4879]) ^ (layer4_outputs[3746]);
    assign layer5_outputs[4955] = layer4_outputs[3459];
    assign layer5_outputs[4956] = ~(layer4_outputs[1098]) | (layer4_outputs[2754]);
    assign layer5_outputs[4957] = (layer4_outputs[1034]) | (layer4_outputs[2302]);
    assign layer5_outputs[4958] = layer4_outputs[4493];
    assign layer5_outputs[4959] = (layer4_outputs[1993]) & ~(layer4_outputs[4818]);
    assign layer5_outputs[4960] = ~((layer4_outputs[2803]) | (layer4_outputs[35]));
    assign layer5_outputs[4961] = (layer4_outputs[4622]) | (layer4_outputs[2663]);
    assign layer5_outputs[4962] = layer4_outputs[1288];
    assign layer5_outputs[4963] = layer4_outputs[4962];
    assign layer5_outputs[4964] = ~((layer4_outputs[235]) | (layer4_outputs[3439]));
    assign layer5_outputs[4965] = (layer4_outputs[4708]) & (layer4_outputs[3934]);
    assign layer5_outputs[4966] = layer4_outputs[1467];
    assign layer5_outputs[4967] = ~(layer4_outputs[630]);
    assign layer5_outputs[4968] = ~(layer4_outputs[1183]);
    assign layer5_outputs[4969] = (layer4_outputs[1933]) | (layer4_outputs[3635]);
    assign layer5_outputs[4970] = ~((layer4_outputs[3939]) ^ (layer4_outputs[4841]));
    assign layer5_outputs[4971] = ~((layer4_outputs[4433]) | (layer4_outputs[2126]));
    assign layer5_outputs[4972] = layer4_outputs[2265];
    assign layer5_outputs[4973] = ~(layer4_outputs[889]) | (layer4_outputs[2738]);
    assign layer5_outputs[4974] = ~((layer4_outputs[2939]) & (layer4_outputs[1757]));
    assign layer5_outputs[4975] = ~(layer4_outputs[5108]);
    assign layer5_outputs[4976] = ~((layer4_outputs[3756]) & (layer4_outputs[1986]));
    assign layer5_outputs[4977] = ~((layer4_outputs[2188]) ^ (layer4_outputs[2176]));
    assign layer5_outputs[4978] = (layer4_outputs[30]) ^ (layer4_outputs[628]);
    assign layer5_outputs[4979] = layer4_outputs[1735];
    assign layer5_outputs[4980] = layer4_outputs[467];
    assign layer5_outputs[4981] = ~(layer4_outputs[736]) | (layer4_outputs[2530]);
    assign layer5_outputs[4982] = ~(layer4_outputs[712]);
    assign layer5_outputs[4983] = layer4_outputs[4562];
    assign layer5_outputs[4984] = layer4_outputs[4916];
    assign layer5_outputs[4985] = 1'b1;
    assign layer5_outputs[4986] = ~((layer4_outputs[2464]) ^ (layer4_outputs[1381]));
    assign layer5_outputs[4987] = ~(layer4_outputs[2545]) | (layer4_outputs[2021]);
    assign layer5_outputs[4988] = layer4_outputs[2314];
    assign layer5_outputs[4989] = layer4_outputs[1672];
    assign layer5_outputs[4990] = layer4_outputs[3639];
    assign layer5_outputs[4991] = ~((layer4_outputs[4888]) & (layer4_outputs[20]));
    assign layer5_outputs[4992] = (layer4_outputs[488]) ^ (layer4_outputs[1841]);
    assign layer5_outputs[4993] = ~((layer4_outputs[2899]) & (layer4_outputs[874]));
    assign layer5_outputs[4994] = (layer4_outputs[4360]) & (layer4_outputs[1460]);
    assign layer5_outputs[4995] = layer4_outputs[1770];
    assign layer5_outputs[4996] = ~(layer4_outputs[2611]);
    assign layer5_outputs[4997] = ~(layer4_outputs[40]) | (layer4_outputs[569]);
    assign layer5_outputs[4998] = (layer4_outputs[161]) ^ (layer4_outputs[4965]);
    assign layer5_outputs[4999] = (layer4_outputs[2432]) | (layer4_outputs[967]);
    assign layer5_outputs[5000] = (layer4_outputs[1394]) | (layer4_outputs[1643]);
    assign layer5_outputs[5001] = ~(layer4_outputs[2615]) | (layer4_outputs[4845]);
    assign layer5_outputs[5002] = ~(layer4_outputs[12]) | (layer4_outputs[2125]);
    assign layer5_outputs[5003] = (layer4_outputs[167]) & ~(layer4_outputs[1384]);
    assign layer5_outputs[5004] = layer4_outputs[1784];
    assign layer5_outputs[5005] = layer4_outputs[3640];
    assign layer5_outputs[5006] = (layer4_outputs[703]) ^ (layer4_outputs[4230]);
    assign layer5_outputs[5007] = layer4_outputs[5078];
    assign layer5_outputs[5008] = ~(layer4_outputs[4496]);
    assign layer5_outputs[5009] = (layer4_outputs[4700]) & ~(layer4_outputs[2299]);
    assign layer5_outputs[5010] = ~(layer4_outputs[2861]);
    assign layer5_outputs[5011] = ~((layer4_outputs[3503]) ^ (layer4_outputs[1807]));
    assign layer5_outputs[5012] = ~(layer4_outputs[2337]) | (layer4_outputs[4386]);
    assign layer5_outputs[5013] = 1'b0;
    assign layer5_outputs[5014] = 1'b0;
    assign layer5_outputs[5015] = layer4_outputs[921];
    assign layer5_outputs[5016] = ~(layer4_outputs[697]);
    assign layer5_outputs[5017] = layer4_outputs[2685];
    assign layer5_outputs[5018] = layer4_outputs[2964];
    assign layer5_outputs[5019] = ~((layer4_outputs[3300]) | (layer4_outputs[814]));
    assign layer5_outputs[5020] = (layer4_outputs[1856]) | (layer4_outputs[3039]);
    assign layer5_outputs[5021] = ~(layer4_outputs[2794]);
    assign layer5_outputs[5022] = ~((layer4_outputs[1926]) ^ (layer4_outputs[3414]));
    assign layer5_outputs[5023] = (layer4_outputs[1871]) & ~(layer4_outputs[2825]);
    assign layer5_outputs[5024] = ~(layer4_outputs[884]);
    assign layer5_outputs[5025] = ~(layer4_outputs[671]);
    assign layer5_outputs[5026] = (layer4_outputs[1189]) | (layer4_outputs[912]);
    assign layer5_outputs[5027] = ~(layer4_outputs[4031]) | (layer4_outputs[1839]);
    assign layer5_outputs[5028] = (layer4_outputs[684]) & ~(layer4_outputs[2951]);
    assign layer5_outputs[5029] = layer4_outputs[3344];
    assign layer5_outputs[5030] = (layer4_outputs[2550]) & (layer4_outputs[88]);
    assign layer5_outputs[5031] = ~(layer4_outputs[1852]);
    assign layer5_outputs[5032] = 1'b0;
    assign layer5_outputs[5033] = layer4_outputs[4653];
    assign layer5_outputs[5034] = (layer4_outputs[3373]) & ~(layer4_outputs[3586]);
    assign layer5_outputs[5035] = ~((layer4_outputs[1939]) | (layer4_outputs[438]));
    assign layer5_outputs[5036] = ~(layer4_outputs[1923]);
    assign layer5_outputs[5037] = (layer4_outputs[2747]) & ~(layer4_outputs[1598]);
    assign layer5_outputs[5038] = 1'b1;
    assign layer5_outputs[5039] = 1'b0;
    assign layer5_outputs[5040] = ~((layer4_outputs[828]) & (layer4_outputs[5043]));
    assign layer5_outputs[5041] = layer4_outputs[3074];
    assign layer5_outputs[5042] = ~((layer4_outputs[901]) | (layer4_outputs[2982]));
    assign layer5_outputs[5043] = ~(layer4_outputs[3901]);
    assign layer5_outputs[5044] = ~(layer4_outputs[2698]) | (layer4_outputs[2276]);
    assign layer5_outputs[5045] = ~(layer4_outputs[1412]) | (layer4_outputs[1251]);
    assign layer5_outputs[5046] = layer4_outputs[4716];
    assign layer5_outputs[5047] = ~(layer4_outputs[4354]) | (layer4_outputs[4544]);
    assign layer5_outputs[5048] = ~(layer4_outputs[3117]);
    assign layer5_outputs[5049] = 1'b0;
    assign layer5_outputs[5050] = 1'b1;
    assign layer5_outputs[5051] = ~(layer4_outputs[2064]) | (layer4_outputs[4096]);
    assign layer5_outputs[5052] = (layer4_outputs[4999]) & (layer4_outputs[181]);
    assign layer5_outputs[5053] = layer4_outputs[318];
    assign layer5_outputs[5054] = (layer4_outputs[3143]) | (layer4_outputs[879]);
    assign layer5_outputs[5055] = (layer4_outputs[1278]) & ~(layer4_outputs[1890]);
    assign layer5_outputs[5056] = layer4_outputs[4480];
    assign layer5_outputs[5057] = (layer4_outputs[3020]) | (layer4_outputs[210]);
    assign layer5_outputs[5058] = ~((layer4_outputs[2246]) ^ (layer4_outputs[993]));
    assign layer5_outputs[5059] = (layer4_outputs[4050]) & ~(layer4_outputs[163]);
    assign layer5_outputs[5060] = layer4_outputs[2588];
    assign layer5_outputs[5061] = layer4_outputs[3914];
    assign layer5_outputs[5062] = ~(layer4_outputs[2092]);
    assign layer5_outputs[5063] = layer4_outputs[952];
    assign layer5_outputs[5064] = 1'b0;
    assign layer5_outputs[5065] = ~((layer4_outputs[405]) ^ (layer4_outputs[2477]));
    assign layer5_outputs[5066] = (layer4_outputs[3919]) & (layer4_outputs[1989]);
    assign layer5_outputs[5067] = layer4_outputs[3412];
    assign layer5_outputs[5068] = (layer4_outputs[3194]) & ~(layer4_outputs[3337]);
    assign layer5_outputs[5069] = ~(layer4_outputs[914]);
    assign layer5_outputs[5070] = ~(layer4_outputs[2329]);
    assign layer5_outputs[5071] = (layer4_outputs[3190]) ^ (layer4_outputs[2969]);
    assign layer5_outputs[5072] = ~(layer4_outputs[2775]);
    assign layer5_outputs[5073] = (layer4_outputs[924]) | (layer4_outputs[1296]);
    assign layer5_outputs[5074] = layer4_outputs[4206];
    assign layer5_outputs[5075] = layer4_outputs[1590];
    assign layer5_outputs[5076] = ~(layer4_outputs[1507]);
    assign layer5_outputs[5077] = layer4_outputs[64];
    assign layer5_outputs[5078] = (layer4_outputs[841]) ^ (layer4_outputs[3946]);
    assign layer5_outputs[5079] = ~(layer4_outputs[727]);
    assign layer5_outputs[5080] = layer4_outputs[3507];
    assign layer5_outputs[5081] = ~((layer4_outputs[4129]) | (layer4_outputs[4412]));
    assign layer5_outputs[5082] = (layer4_outputs[3236]) & ~(layer4_outputs[1450]);
    assign layer5_outputs[5083] = 1'b1;
    assign layer5_outputs[5084] = layer4_outputs[725];
    assign layer5_outputs[5085] = 1'b0;
    assign layer5_outputs[5086] = (layer4_outputs[4620]) & ~(layer4_outputs[4058]);
    assign layer5_outputs[5087] = layer4_outputs[1847];
    assign layer5_outputs[5088] = (layer4_outputs[856]) & (layer4_outputs[1089]);
    assign layer5_outputs[5089] = ~((layer4_outputs[136]) & (layer4_outputs[182]));
    assign layer5_outputs[5090] = ~(layer4_outputs[2561]);
    assign layer5_outputs[5091] = ~(layer4_outputs[1065]);
    assign layer5_outputs[5092] = ~(layer4_outputs[3383]) | (layer4_outputs[1498]);
    assign layer5_outputs[5093] = ~(layer4_outputs[23]);
    assign layer5_outputs[5094] = 1'b1;
    assign layer5_outputs[5095] = ~(layer4_outputs[3130]);
    assign layer5_outputs[5096] = ~(layer4_outputs[1391]) | (layer4_outputs[4658]);
    assign layer5_outputs[5097] = (layer4_outputs[1187]) & (layer4_outputs[877]);
    assign layer5_outputs[5098] = ~((layer4_outputs[1428]) | (layer4_outputs[3803]));
    assign layer5_outputs[5099] = ~(layer4_outputs[1610]);
    assign layer5_outputs[5100] = layer4_outputs[1032];
    assign layer5_outputs[5101] = ~(layer4_outputs[1714]);
    assign layer5_outputs[5102] = ~((layer4_outputs[3111]) & (layer4_outputs[3524]));
    assign layer5_outputs[5103] = (layer4_outputs[1268]) ^ (layer4_outputs[2007]);
    assign layer5_outputs[5104] = 1'b1;
    assign layer5_outputs[5105] = (layer4_outputs[3474]) ^ (layer4_outputs[4037]);
    assign layer5_outputs[5106] = layer4_outputs[4468];
    assign layer5_outputs[5107] = ~(layer4_outputs[1977]);
    assign layer5_outputs[5108] = ~(layer4_outputs[3005]);
    assign layer5_outputs[5109] = layer4_outputs[3476];
    assign layer5_outputs[5110] = ~(layer4_outputs[4125]) | (layer4_outputs[2550]);
    assign layer5_outputs[5111] = (layer4_outputs[3808]) & ~(layer4_outputs[983]);
    assign layer5_outputs[5112] = ~(layer4_outputs[105]);
    assign layer5_outputs[5113] = ~((layer4_outputs[384]) & (layer4_outputs[1918]));
    assign layer5_outputs[5114] = layer4_outputs[1434];
    assign layer5_outputs[5115] = (layer4_outputs[1532]) | (layer4_outputs[1951]);
    assign layer5_outputs[5116] = layer4_outputs[4533];
    assign layer5_outputs[5117] = layer4_outputs[1697];
    assign layer5_outputs[5118] = (layer4_outputs[2615]) ^ (layer4_outputs[803]);
    assign layer5_outputs[5119] = (layer4_outputs[415]) ^ (layer4_outputs[1207]);
    assign layer6_outputs[0] = layer5_outputs[1456];
    assign layer6_outputs[1] = ~((layer5_outputs[57]) ^ (layer5_outputs[2363]));
    assign layer6_outputs[2] = layer5_outputs[2162];
    assign layer6_outputs[3] = ~((layer5_outputs[4109]) ^ (layer5_outputs[801]));
    assign layer6_outputs[4] = ~((layer5_outputs[3029]) & (layer5_outputs[2548]));
    assign layer6_outputs[5] = (layer5_outputs[954]) & (layer5_outputs[4473]);
    assign layer6_outputs[6] = layer5_outputs[4499];
    assign layer6_outputs[7] = layer5_outputs[1830];
    assign layer6_outputs[8] = layer5_outputs[945];
    assign layer6_outputs[9] = ~((layer5_outputs[3064]) ^ (layer5_outputs[611]));
    assign layer6_outputs[10] = ~((layer5_outputs[4450]) ^ (layer5_outputs[563]));
    assign layer6_outputs[11] = ~((layer5_outputs[1375]) ^ (layer5_outputs[4241]));
    assign layer6_outputs[12] = ~(layer5_outputs[4142]);
    assign layer6_outputs[13] = layer5_outputs[1523];
    assign layer6_outputs[14] = ~((layer5_outputs[267]) ^ (layer5_outputs[1075]));
    assign layer6_outputs[15] = layer5_outputs[2585];
    assign layer6_outputs[16] = (layer5_outputs[1952]) | (layer5_outputs[3179]);
    assign layer6_outputs[17] = ~(layer5_outputs[853]);
    assign layer6_outputs[18] = (layer5_outputs[3166]) | (layer5_outputs[2241]);
    assign layer6_outputs[19] = (layer5_outputs[4257]) & (layer5_outputs[2942]);
    assign layer6_outputs[20] = ~(layer5_outputs[3130]);
    assign layer6_outputs[21] = ~(layer5_outputs[2558]) | (layer5_outputs[810]);
    assign layer6_outputs[22] = ~(layer5_outputs[940]);
    assign layer6_outputs[23] = (layer5_outputs[294]) & ~(layer5_outputs[850]);
    assign layer6_outputs[24] = layer5_outputs[3922];
    assign layer6_outputs[25] = ~((layer5_outputs[1720]) ^ (layer5_outputs[5100]));
    assign layer6_outputs[26] = layer5_outputs[4593];
    assign layer6_outputs[27] = ~((layer5_outputs[2432]) ^ (layer5_outputs[4900]));
    assign layer6_outputs[28] = ~(layer5_outputs[1329]);
    assign layer6_outputs[29] = layer5_outputs[3850];
    assign layer6_outputs[30] = (layer5_outputs[4377]) & (layer5_outputs[3164]);
    assign layer6_outputs[31] = layer5_outputs[5116];
    assign layer6_outputs[32] = layer5_outputs[651];
    assign layer6_outputs[33] = ~(layer5_outputs[1835]);
    assign layer6_outputs[34] = layer5_outputs[1457];
    assign layer6_outputs[35] = (layer5_outputs[3116]) | (layer5_outputs[2278]);
    assign layer6_outputs[36] = 1'b0;
    assign layer6_outputs[37] = ~((layer5_outputs[2518]) & (layer5_outputs[3301]));
    assign layer6_outputs[38] = ~(layer5_outputs[1147]);
    assign layer6_outputs[39] = ~(layer5_outputs[1421]);
    assign layer6_outputs[40] = (layer5_outputs[2869]) & ~(layer5_outputs[1247]);
    assign layer6_outputs[41] = layer5_outputs[107];
    assign layer6_outputs[42] = ~(layer5_outputs[798]) | (layer5_outputs[3219]);
    assign layer6_outputs[43] = layer5_outputs[4758];
    assign layer6_outputs[44] = ~(layer5_outputs[3362]);
    assign layer6_outputs[45] = ~((layer5_outputs[1719]) ^ (layer5_outputs[4496]));
    assign layer6_outputs[46] = (layer5_outputs[2569]) ^ (layer5_outputs[1484]);
    assign layer6_outputs[47] = (layer5_outputs[2037]) & ~(layer5_outputs[1179]);
    assign layer6_outputs[48] = ~(layer5_outputs[3690]);
    assign layer6_outputs[49] = ~(layer5_outputs[1178]);
    assign layer6_outputs[50] = layer5_outputs[4986];
    assign layer6_outputs[51] = ~(layer5_outputs[2488]) | (layer5_outputs[4897]);
    assign layer6_outputs[52] = 1'b1;
    assign layer6_outputs[53] = ~(layer5_outputs[2084]) | (layer5_outputs[1793]);
    assign layer6_outputs[54] = ~(layer5_outputs[4819]);
    assign layer6_outputs[55] = ~(layer5_outputs[1804]) | (layer5_outputs[5042]);
    assign layer6_outputs[56] = layer5_outputs[2044];
    assign layer6_outputs[57] = (layer5_outputs[182]) & (layer5_outputs[2774]);
    assign layer6_outputs[58] = ~((layer5_outputs[2448]) ^ (layer5_outputs[2023]));
    assign layer6_outputs[59] = 1'b1;
    assign layer6_outputs[60] = ~(layer5_outputs[2201]);
    assign layer6_outputs[61] = ~((layer5_outputs[3664]) & (layer5_outputs[3300]));
    assign layer6_outputs[62] = layer5_outputs[3465];
    assign layer6_outputs[63] = layer5_outputs[893];
    assign layer6_outputs[64] = (layer5_outputs[578]) ^ (layer5_outputs[2378]);
    assign layer6_outputs[65] = ~(layer5_outputs[4873]);
    assign layer6_outputs[66] = ~(layer5_outputs[1164]) | (layer5_outputs[3752]);
    assign layer6_outputs[67] = ~(layer5_outputs[934]);
    assign layer6_outputs[68] = layer5_outputs[4079];
    assign layer6_outputs[69] = ~(layer5_outputs[2029]);
    assign layer6_outputs[70] = ~(layer5_outputs[4979]);
    assign layer6_outputs[71] = (layer5_outputs[645]) & ~(layer5_outputs[5071]);
    assign layer6_outputs[72] = ~(layer5_outputs[3782]);
    assign layer6_outputs[73] = ~((layer5_outputs[3652]) ^ (layer5_outputs[4108]));
    assign layer6_outputs[74] = (layer5_outputs[2509]) | (layer5_outputs[4493]);
    assign layer6_outputs[75] = ~(layer5_outputs[5097]) | (layer5_outputs[1287]);
    assign layer6_outputs[76] = ~((layer5_outputs[4533]) & (layer5_outputs[2712]));
    assign layer6_outputs[77] = (layer5_outputs[890]) ^ (layer5_outputs[1660]);
    assign layer6_outputs[78] = layer5_outputs[15];
    assign layer6_outputs[79] = layer5_outputs[3493];
    assign layer6_outputs[80] = ~(layer5_outputs[3939]);
    assign layer6_outputs[81] = ~(layer5_outputs[4178]) | (layer5_outputs[708]);
    assign layer6_outputs[82] = ~(layer5_outputs[956]);
    assign layer6_outputs[83] = ~(layer5_outputs[3898]);
    assign layer6_outputs[84] = (layer5_outputs[1221]) ^ (layer5_outputs[2417]);
    assign layer6_outputs[85] = layer5_outputs[243];
    assign layer6_outputs[86] = ~((layer5_outputs[400]) ^ (layer5_outputs[3170]));
    assign layer6_outputs[87] = layer5_outputs[4065];
    assign layer6_outputs[88] = (layer5_outputs[889]) & (layer5_outputs[2985]);
    assign layer6_outputs[89] = ~(layer5_outputs[4124]);
    assign layer6_outputs[90] = (layer5_outputs[4727]) | (layer5_outputs[2672]);
    assign layer6_outputs[91] = (layer5_outputs[567]) & (layer5_outputs[1542]);
    assign layer6_outputs[92] = layer5_outputs[1091];
    assign layer6_outputs[93] = (layer5_outputs[3643]) & (layer5_outputs[1549]);
    assign layer6_outputs[94] = ~((layer5_outputs[622]) ^ (layer5_outputs[113]));
    assign layer6_outputs[95] = ~(layer5_outputs[4240]);
    assign layer6_outputs[96] = (layer5_outputs[4062]) ^ (layer5_outputs[4280]);
    assign layer6_outputs[97] = (layer5_outputs[2033]) ^ (layer5_outputs[912]);
    assign layer6_outputs[98] = ~(layer5_outputs[3072]);
    assign layer6_outputs[99] = (layer5_outputs[561]) ^ (layer5_outputs[263]);
    assign layer6_outputs[100] = layer5_outputs[3296];
    assign layer6_outputs[101] = layer5_outputs[2203];
    assign layer6_outputs[102] = (layer5_outputs[4926]) & (layer5_outputs[1280]);
    assign layer6_outputs[103] = ~(layer5_outputs[801]);
    assign layer6_outputs[104] = (layer5_outputs[1190]) | (layer5_outputs[3070]);
    assign layer6_outputs[105] = ~(layer5_outputs[2073]);
    assign layer6_outputs[106] = (layer5_outputs[2592]) | (layer5_outputs[1615]);
    assign layer6_outputs[107] = layer5_outputs[3284];
    assign layer6_outputs[108] = ~(layer5_outputs[666]);
    assign layer6_outputs[109] = ~(layer5_outputs[2280]);
    assign layer6_outputs[110] = ~(layer5_outputs[3804]) | (layer5_outputs[4867]);
    assign layer6_outputs[111] = ~(layer5_outputs[3232]) | (layer5_outputs[1551]);
    assign layer6_outputs[112] = (layer5_outputs[5114]) & ~(layer5_outputs[2554]);
    assign layer6_outputs[113] = ~(layer5_outputs[31]);
    assign layer6_outputs[114] = (layer5_outputs[4898]) & ~(layer5_outputs[1281]);
    assign layer6_outputs[115] = ~(layer5_outputs[4789]);
    assign layer6_outputs[116] = layer5_outputs[198];
    assign layer6_outputs[117] = ~(layer5_outputs[3220]);
    assign layer6_outputs[118] = layer5_outputs[2436];
    assign layer6_outputs[119] = (layer5_outputs[2331]) & ~(layer5_outputs[2889]);
    assign layer6_outputs[120] = layer5_outputs[3478];
    assign layer6_outputs[121] = ~(layer5_outputs[1246]);
    assign layer6_outputs[122] = ~(layer5_outputs[918]);
    assign layer6_outputs[123] = ~(layer5_outputs[1086]);
    assign layer6_outputs[124] = ~((layer5_outputs[2552]) | (layer5_outputs[4949]));
    assign layer6_outputs[125] = ~(layer5_outputs[1187]);
    assign layer6_outputs[126] = layer5_outputs[4857];
    assign layer6_outputs[127] = ~(layer5_outputs[4149]) | (layer5_outputs[4028]);
    assign layer6_outputs[128] = ~(layer5_outputs[1762]);
    assign layer6_outputs[129] = (layer5_outputs[2190]) ^ (layer5_outputs[485]);
    assign layer6_outputs[130] = (layer5_outputs[3383]) | (layer5_outputs[2105]);
    assign layer6_outputs[131] = ~(layer5_outputs[3675]);
    assign layer6_outputs[132] = ~((layer5_outputs[1369]) ^ (layer5_outputs[2693]));
    assign layer6_outputs[133] = 1'b1;
    assign layer6_outputs[134] = (layer5_outputs[2317]) & (layer5_outputs[4432]);
    assign layer6_outputs[135] = ~(layer5_outputs[30]);
    assign layer6_outputs[136] = ~(layer5_outputs[4112]);
    assign layer6_outputs[137] = (layer5_outputs[974]) & ~(layer5_outputs[4149]);
    assign layer6_outputs[138] = 1'b0;
    assign layer6_outputs[139] = ~(layer5_outputs[1858]);
    assign layer6_outputs[140] = ~(layer5_outputs[1448]) | (layer5_outputs[4213]);
    assign layer6_outputs[141] = (layer5_outputs[1101]) | (layer5_outputs[360]);
    assign layer6_outputs[142] = layer5_outputs[3136];
    assign layer6_outputs[143] = ~((layer5_outputs[698]) & (layer5_outputs[4551]));
    assign layer6_outputs[144] = ~(layer5_outputs[4708]);
    assign layer6_outputs[145] = (layer5_outputs[2401]) & ~(layer5_outputs[2409]);
    assign layer6_outputs[146] = ~(layer5_outputs[466]);
    assign layer6_outputs[147] = layer5_outputs[37];
    assign layer6_outputs[148] = ~(layer5_outputs[1781]);
    assign layer6_outputs[149] = (layer5_outputs[1891]) ^ (layer5_outputs[543]);
    assign layer6_outputs[150] = layer5_outputs[3182];
    assign layer6_outputs[151] = layer5_outputs[754];
    assign layer6_outputs[152] = 1'b0;
    assign layer6_outputs[153] = ~(layer5_outputs[1680]);
    assign layer6_outputs[154] = ~((layer5_outputs[2063]) ^ (layer5_outputs[441]));
    assign layer6_outputs[155] = ~(layer5_outputs[476]);
    assign layer6_outputs[156] = ~(layer5_outputs[2741]);
    assign layer6_outputs[157] = ~(layer5_outputs[150]);
    assign layer6_outputs[158] = ~(layer5_outputs[1117]);
    assign layer6_outputs[159] = ~(layer5_outputs[1043]);
    assign layer6_outputs[160] = layer5_outputs[5006];
    assign layer6_outputs[161] = ~(layer5_outputs[4484]);
    assign layer6_outputs[162] = ~(layer5_outputs[223]);
    assign layer6_outputs[163] = layer5_outputs[2724];
    assign layer6_outputs[164] = (layer5_outputs[1880]) | (layer5_outputs[971]);
    assign layer6_outputs[165] = layer5_outputs[4238];
    assign layer6_outputs[166] = layer5_outputs[2912];
    assign layer6_outputs[167] = ~(layer5_outputs[747]);
    assign layer6_outputs[168] = (layer5_outputs[97]) ^ (layer5_outputs[4083]);
    assign layer6_outputs[169] = layer5_outputs[1745];
    assign layer6_outputs[170] = ~((layer5_outputs[2584]) | (layer5_outputs[4642]));
    assign layer6_outputs[171] = ~(layer5_outputs[2030]);
    assign layer6_outputs[172] = ~((layer5_outputs[3847]) | (layer5_outputs[3177]));
    assign layer6_outputs[173] = 1'b1;
    assign layer6_outputs[174] = ~(layer5_outputs[2662]);
    assign layer6_outputs[175] = layer5_outputs[2982];
    assign layer6_outputs[176] = ~(layer5_outputs[2014]);
    assign layer6_outputs[177] = layer5_outputs[682];
    assign layer6_outputs[178] = layer5_outputs[3021];
    assign layer6_outputs[179] = (layer5_outputs[3304]) ^ (layer5_outputs[4205]);
    assign layer6_outputs[180] = layer5_outputs[2428];
    assign layer6_outputs[181] = (layer5_outputs[2537]) ^ (layer5_outputs[770]);
    assign layer6_outputs[182] = layer5_outputs[55];
    assign layer6_outputs[183] = layer5_outputs[756];
    assign layer6_outputs[184] = ~(layer5_outputs[781]);
    assign layer6_outputs[185] = (layer5_outputs[1608]) & (layer5_outputs[2707]);
    assign layer6_outputs[186] = layer5_outputs[3619];
    assign layer6_outputs[187] = (layer5_outputs[4078]) | (layer5_outputs[272]);
    assign layer6_outputs[188] = ~(layer5_outputs[4850]) | (layer5_outputs[1356]);
    assign layer6_outputs[189] = (layer5_outputs[3790]) & ~(layer5_outputs[3580]);
    assign layer6_outputs[190] = (layer5_outputs[884]) & ~(layer5_outputs[183]);
    assign layer6_outputs[191] = (layer5_outputs[4568]) & (layer5_outputs[4222]);
    assign layer6_outputs[192] = layer5_outputs[275];
    assign layer6_outputs[193] = layer5_outputs[1173];
    assign layer6_outputs[194] = layer5_outputs[3859];
    assign layer6_outputs[195] = layer5_outputs[2403];
    assign layer6_outputs[196] = (layer5_outputs[3262]) ^ (layer5_outputs[1475]);
    assign layer6_outputs[197] = ~((layer5_outputs[2410]) ^ (layer5_outputs[25]));
    assign layer6_outputs[198] = (layer5_outputs[3794]) | (layer5_outputs[3351]);
    assign layer6_outputs[199] = ~(layer5_outputs[3229]) | (layer5_outputs[2717]);
    assign layer6_outputs[200] = (layer5_outputs[4963]) ^ (layer5_outputs[845]);
    assign layer6_outputs[201] = layer5_outputs[2208];
    assign layer6_outputs[202] = ~(layer5_outputs[4718]);
    assign layer6_outputs[203] = 1'b1;
    assign layer6_outputs[204] = ~(layer5_outputs[1892]);
    assign layer6_outputs[205] = ~(layer5_outputs[1420]);
    assign layer6_outputs[206] = ~((layer5_outputs[4372]) & (layer5_outputs[2845]));
    assign layer6_outputs[207] = ~(layer5_outputs[4188]);
    assign layer6_outputs[208] = (layer5_outputs[2122]) ^ (layer5_outputs[5072]);
    assign layer6_outputs[209] = ~(layer5_outputs[1924]);
    assign layer6_outputs[210] = ~(layer5_outputs[4889]);
    assign layer6_outputs[211] = ~(layer5_outputs[1621]) | (layer5_outputs[4468]);
    assign layer6_outputs[212] = layer5_outputs[120];
    assign layer6_outputs[213] = (layer5_outputs[4666]) ^ (layer5_outputs[2476]);
    assign layer6_outputs[214] = layer5_outputs[1691];
    assign layer6_outputs[215] = ~(layer5_outputs[3842]);
    assign layer6_outputs[216] = ~(layer5_outputs[4908]);
    assign layer6_outputs[217] = (layer5_outputs[4347]) & (layer5_outputs[2366]);
    assign layer6_outputs[218] = ~(layer5_outputs[3561]);
    assign layer6_outputs[219] = (layer5_outputs[2371]) & ~(layer5_outputs[1167]);
    assign layer6_outputs[220] = ~(layer5_outputs[244]);
    assign layer6_outputs[221] = layer5_outputs[4723];
    assign layer6_outputs[222] = (layer5_outputs[3591]) ^ (layer5_outputs[333]);
    assign layer6_outputs[223] = layer5_outputs[3741];
    assign layer6_outputs[224] = ~(layer5_outputs[2755]) | (layer5_outputs[2105]);
    assign layer6_outputs[225] = 1'b0;
    assign layer6_outputs[226] = ~(layer5_outputs[676]);
    assign layer6_outputs[227] = ~(layer5_outputs[19]);
    assign layer6_outputs[228] = layer5_outputs[1928];
    assign layer6_outputs[229] = ~(layer5_outputs[4848]);
    assign layer6_outputs[230] = ~(layer5_outputs[2751]);
    assign layer6_outputs[231] = ~(layer5_outputs[4507]);
    assign layer6_outputs[232] = ~((layer5_outputs[5028]) | (layer5_outputs[1089]));
    assign layer6_outputs[233] = (layer5_outputs[2778]) & ~(layer5_outputs[2344]);
    assign layer6_outputs[234] = ~((layer5_outputs[3744]) ^ (layer5_outputs[5008]));
    assign layer6_outputs[235] = ~((layer5_outputs[4801]) ^ (layer5_outputs[2658]));
    assign layer6_outputs[236] = layer5_outputs[2438];
    assign layer6_outputs[237] = ~(layer5_outputs[4548]) | (layer5_outputs[4767]);
    assign layer6_outputs[238] = ~(layer5_outputs[2235]);
    assign layer6_outputs[239] = (layer5_outputs[609]) & (layer5_outputs[213]);
    assign layer6_outputs[240] = ~(layer5_outputs[3241]);
    assign layer6_outputs[241] = ~(layer5_outputs[2360]);
    assign layer6_outputs[242] = layer5_outputs[3379];
    assign layer6_outputs[243] = ~(layer5_outputs[2617]);
    assign layer6_outputs[244] = ~(layer5_outputs[4180]) | (layer5_outputs[1228]);
    assign layer6_outputs[245] = layer5_outputs[4231];
    assign layer6_outputs[246] = ~((layer5_outputs[2573]) ^ (layer5_outputs[4422]));
    assign layer6_outputs[247] = ~(layer5_outputs[3549]);
    assign layer6_outputs[248] = ~((layer5_outputs[1944]) ^ (layer5_outputs[3930]));
    assign layer6_outputs[249] = (layer5_outputs[2486]) ^ (layer5_outputs[3466]);
    assign layer6_outputs[250] = ~(layer5_outputs[4426]);
    assign layer6_outputs[251] = ~(layer5_outputs[1]);
    assign layer6_outputs[252] = (layer5_outputs[3353]) & (layer5_outputs[751]);
    assign layer6_outputs[253] = layer5_outputs[4835];
    assign layer6_outputs[254] = 1'b1;
    assign layer6_outputs[255] = (layer5_outputs[3303]) ^ (layer5_outputs[706]);
    assign layer6_outputs[256] = layer5_outputs[541];
    assign layer6_outputs[257] = (layer5_outputs[5075]) & ~(layer5_outputs[5070]);
    assign layer6_outputs[258] = layer5_outputs[1039];
    assign layer6_outputs[259] = ~(layer5_outputs[2243]);
    assign layer6_outputs[260] = ~((layer5_outputs[3319]) ^ (layer5_outputs[702]));
    assign layer6_outputs[261] = ~((layer5_outputs[2893]) & (layer5_outputs[3042]));
    assign layer6_outputs[262] = (layer5_outputs[832]) | (layer5_outputs[2828]);
    assign layer6_outputs[263] = ~(layer5_outputs[3569]);
    assign layer6_outputs[264] = layer5_outputs[2579];
    assign layer6_outputs[265] = ~(layer5_outputs[1735]);
    assign layer6_outputs[266] = layer5_outputs[3005];
    assign layer6_outputs[267] = layer5_outputs[1762];
    assign layer6_outputs[268] = ~(layer5_outputs[3325]);
    assign layer6_outputs[269] = layer5_outputs[2689];
    assign layer6_outputs[270] = ~(layer5_outputs[3932]);
    assign layer6_outputs[271] = ~(layer5_outputs[4048]);
    assign layer6_outputs[272] = 1'b1;
    assign layer6_outputs[273] = layer5_outputs[1523];
    assign layer6_outputs[274] = ~(layer5_outputs[501]);
    assign layer6_outputs[275] = ~((layer5_outputs[508]) & (layer5_outputs[2331]));
    assign layer6_outputs[276] = ~(layer5_outputs[3740]);
    assign layer6_outputs[277] = ~(layer5_outputs[755]);
    assign layer6_outputs[278] = layer5_outputs[3764];
    assign layer6_outputs[279] = layer5_outputs[3175];
    assign layer6_outputs[280] = ~(layer5_outputs[888]);
    assign layer6_outputs[281] = layer5_outputs[1784];
    assign layer6_outputs[282] = ~(layer5_outputs[4813]);
    assign layer6_outputs[283] = layer5_outputs[4062];
    assign layer6_outputs[284] = ~(layer5_outputs[3852]);
    assign layer6_outputs[285] = ~((layer5_outputs[3985]) | (layer5_outputs[5012]));
    assign layer6_outputs[286] = layer5_outputs[2795];
    assign layer6_outputs[287] = ~(layer5_outputs[4582]);
    assign layer6_outputs[288] = ~(layer5_outputs[2295]);
    assign layer6_outputs[289] = (layer5_outputs[2783]) | (layer5_outputs[1224]);
    assign layer6_outputs[290] = layer5_outputs[2673];
    assign layer6_outputs[291] = ~(layer5_outputs[1082]) | (layer5_outputs[3778]);
    assign layer6_outputs[292] = ~(layer5_outputs[2807]);
    assign layer6_outputs[293] = (layer5_outputs[2605]) | (layer5_outputs[1339]);
    assign layer6_outputs[294] = (layer5_outputs[46]) ^ (layer5_outputs[1887]);
    assign layer6_outputs[295] = layer5_outputs[170];
    assign layer6_outputs[296] = layer5_outputs[2429];
    assign layer6_outputs[297] = ~(layer5_outputs[2834]);
    assign layer6_outputs[298] = layer5_outputs[2451];
    assign layer6_outputs[299] = ~(layer5_outputs[1378]) | (layer5_outputs[3390]);
    assign layer6_outputs[300] = ~((layer5_outputs[335]) ^ (layer5_outputs[1953]));
    assign layer6_outputs[301] = layer5_outputs[4619];
    assign layer6_outputs[302] = layer5_outputs[1229];
    assign layer6_outputs[303] = layer5_outputs[4693];
    assign layer6_outputs[304] = ~((layer5_outputs[3381]) ^ (layer5_outputs[3435]));
    assign layer6_outputs[305] = (layer5_outputs[1794]) & ~(layer5_outputs[4960]);
    assign layer6_outputs[306] = ~(layer5_outputs[4179]);
    assign layer6_outputs[307] = layer5_outputs[2038];
    assign layer6_outputs[308] = layer5_outputs[1229];
    assign layer6_outputs[309] = ~(layer5_outputs[4950]);
    assign layer6_outputs[310] = ~(layer5_outputs[4008]);
    assign layer6_outputs[311] = ~((layer5_outputs[3070]) ^ (layer5_outputs[402]));
    assign layer6_outputs[312] = ~(layer5_outputs[2094]);
    assign layer6_outputs[313] = layer5_outputs[218];
    assign layer6_outputs[314] = layer5_outputs[321];
    assign layer6_outputs[315] = ~(layer5_outputs[1729]);
    assign layer6_outputs[316] = ~(layer5_outputs[2022]);
    assign layer6_outputs[317] = layer5_outputs[4624];
    assign layer6_outputs[318] = ~((layer5_outputs[2948]) | (layer5_outputs[886]));
    assign layer6_outputs[319] = layer5_outputs[3984];
    assign layer6_outputs[320] = (layer5_outputs[1608]) & (layer5_outputs[2541]);
    assign layer6_outputs[321] = ~(layer5_outputs[3184]);
    assign layer6_outputs[322] = layer5_outputs[980];
    assign layer6_outputs[323] = ~(layer5_outputs[1034]) | (layer5_outputs[2065]);
    assign layer6_outputs[324] = layer5_outputs[4689];
    assign layer6_outputs[325] = ~((layer5_outputs[4799]) & (layer5_outputs[4953]));
    assign layer6_outputs[326] = ~(layer5_outputs[4914]);
    assign layer6_outputs[327] = ~(layer5_outputs[1167]);
    assign layer6_outputs[328] = layer5_outputs[3271];
    assign layer6_outputs[329] = layer5_outputs[3454];
    assign layer6_outputs[330] = layer5_outputs[4475];
    assign layer6_outputs[331] = ~((layer5_outputs[3395]) ^ (layer5_outputs[2854]));
    assign layer6_outputs[332] = ~(layer5_outputs[859]);
    assign layer6_outputs[333] = (layer5_outputs[2226]) & ~(layer5_outputs[3869]);
    assign layer6_outputs[334] = (layer5_outputs[2094]) ^ (layer5_outputs[289]);
    assign layer6_outputs[335] = ~(layer5_outputs[1783]);
    assign layer6_outputs[336] = ~(layer5_outputs[1157]);
    assign layer6_outputs[337] = layer5_outputs[4041];
    assign layer6_outputs[338] = (layer5_outputs[3750]) | (layer5_outputs[4919]);
    assign layer6_outputs[339] = ~((layer5_outputs[1078]) ^ (layer5_outputs[2906]));
    assign layer6_outputs[340] = ~(layer5_outputs[2639]);
    assign layer6_outputs[341] = ~((layer5_outputs[1188]) ^ (layer5_outputs[2988]));
    assign layer6_outputs[342] = ~(layer5_outputs[2648]) | (layer5_outputs[2034]);
    assign layer6_outputs[343] = ~(layer5_outputs[4432]);
    assign layer6_outputs[344] = ~((layer5_outputs[2683]) & (layer5_outputs[1700]));
    assign layer6_outputs[345] = 1'b1;
    assign layer6_outputs[346] = layer5_outputs[3273];
    assign layer6_outputs[347] = ~(layer5_outputs[253]);
    assign layer6_outputs[348] = (layer5_outputs[2883]) & ~(layer5_outputs[4549]);
    assign layer6_outputs[349] = ~((layer5_outputs[574]) ^ (layer5_outputs[206]));
    assign layer6_outputs[350] = ~(layer5_outputs[1809]);
    assign layer6_outputs[351] = ~(layer5_outputs[1641]);
    assign layer6_outputs[352] = (layer5_outputs[4182]) & (layer5_outputs[1279]);
    assign layer6_outputs[353] = ~(layer5_outputs[3058]);
    assign layer6_outputs[354] = layer5_outputs[2588];
    assign layer6_outputs[355] = (layer5_outputs[3429]) ^ (layer5_outputs[4854]);
    assign layer6_outputs[356] = (layer5_outputs[1238]) & (layer5_outputs[4770]);
    assign layer6_outputs[357] = (layer5_outputs[3691]) | (layer5_outputs[4305]);
    assign layer6_outputs[358] = ~(layer5_outputs[1959]);
    assign layer6_outputs[359] = (layer5_outputs[3648]) | (layer5_outputs[4061]);
    assign layer6_outputs[360] = 1'b1;
    assign layer6_outputs[361] = (layer5_outputs[3629]) & ~(layer5_outputs[898]);
    assign layer6_outputs[362] = ~(layer5_outputs[3885]);
    assign layer6_outputs[363] = layer5_outputs[2780];
    assign layer6_outputs[364] = ~(layer5_outputs[696]);
    assign layer6_outputs[365] = layer5_outputs[3286];
    assign layer6_outputs[366] = ~(layer5_outputs[1107]);
    assign layer6_outputs[367] = layer5_outputs[253];
    assign layer6_outputs[368] = (layer5_outputs[1345]) & ~(layer5_outputs[4622]);
    assign layer6_outputs[369] = ~(layer5_outputs[2692]);
    assign layer6_outputs[370] = (layer5_outputs[2079]) | (layer5_outputs[4306]);
    assign layer6_outputs[371] = layer5_outputs[2612];
    assign layer6_outputs[372] = (layer5_outputs[2924]) ^ (layer5_outputs[216]);
    assign layer6_outputs[373] = 1'b1;
    assign layer6_outputs[374] = layer5_outputs[446];
    assign layer6_outputs[375] = ~(layer5_outputs[2555]);
    assign layer6_outputs[376] = layer5_outputs[4327];
    assign layer6_outputs[377] = ~(layer5_outputs[452]) | (layer5_outputs[2143]);
    assign layer6_outputs[378] = ~(layer5_outputs[551]);
    assign layer6_outputs[379] = ~(layer5_outputs[1719]);
    assign layer6_outputs[380] = layer5_outputs[4523];
    assign layer6_outputs[381] = layer5_outputs[2490];
    assign layer6_outputs[382] = ~(layer5_outputs[614]) | (layer5_outputs[2508]);
    assign layer6_outputs[383] = ~((layer5_outputs[4451]) ^ (layer5_outputs[2864]));
    assign layer6_outputs[384] = ~((layer5_outputs[3236]) ^ (layer5_outputs[1736]));
    assign layer6_outputs[385] = ~(layer5_outputs[2365]);
    assign layer6_outputs[386] = ~(layer5_outputs[4173]);
    assign layer6_outputs[387] = ~((layer5_outputs[4326]) | (layer5_outputs[4480]));
    assign layer6_outputs[388] = (layer5_outputs[1245]) & (layer5_outputs[3304]);
    assign layer6_outputs[389] = (layer5_outputs[3885]) ^ (layer5_outputs[4672]);
    assign layer6_outputs[390] = ~((layer5_outputs[3997]) & (layer5_outputs[2642]));
    assign layer6_outputs[391] = layer5_outputs[4192];
    assign layer6_outputs[392] = ~(layer5_outputs[4526]) | (layer5_outputs[2572]);
    assign layer6_outputs[393] = layer5_outputs[4137];
    assign layer6_outputs[394] = layer5_outputs[1707];
    assign layer6_outputs[395] = (layer5_outputs[4711]) & (layer5_outputs[4666]);
    assign layer6_outputs[396] = layer5_outputs[1225];
    assign layer6_outputs[397] = ~(layer5_outputs[2703]);
    assign layer6_outputs[398] = layer5_outputs[1547];
    assign layer6_outputs[399] = ~(layer5_outputs[3839]);
    assign layer6_outputs[400] = layer5_outputs[1440];
    assign layer6_outputs[401] = ~((layer5_outputs[1322]) ^ (layer5_outputs[4832]));
    assign layer6_outputs[402] = (layer5_outputs[716]) & ~(layer5_outputs[3832]);
    assign layer6_outputs[403] = (layer5_outputs[868]) ^ (layer5_outputs[2419]);
    assign layer6_outputs[404] = layer5_outputs[1900];
    assign layer6_outputs[405] = layer5_outputs[2910];
    assign layer6_outputs[406] = (layer5_outputs[227]) & (layer5_outputs[3963]);
    assign layer6_outputs[407] = ~((layer5_outputs[2449]) & (layer5_outputs[2857]));
    assign layer6_outputs[408] = ~(layer5_outputs[4996]);
    assign layer6_outputs[409] = 1'b0;
    assign layer6_outputs[410] = ~(layer5_outputs[1852]);
    assign layer6_outputs[411] = (layer5_outputs[1559]) & (layer5_outputs[4197]);
    assign layer6_outputs[412] = ~(layer5_outputs[2807]);
    assign layer6_outputs[413] = (layer5_outputs[1529]) & ~(layer5_outputs[909]);
    assign layer6_outputs[414] = (layer5_outputs[1181]) & ~(layer5_outputs[3356]);
    assign layer6_outputs[415] = ~(layer5_outputs[4305]);
    assign layer6_outputs[416] = ~((layer5_outputs[1038]) ^ (layer5_outputs[492]));
    assign layer6_outputs[417] = 1'b0;
    assign layer6_outputs[418] = layer5_outputs[276];
    assign layer6_outputs[419] = ~(layer5_outputs[3218]);
    assign layer6_outputs[420] = layer5_outputs[1863];
    assign layer6_outputs[421] = ~((layer5_outputs[4709]) ^ (layer5_outputs[1891]));
    assign layer6_outputs[422] = ~((layer5_outputs[4126]) & (layer5_outputs[1322]));
    assign layer6_outputs[423] = layer5_outputs[290];
    assign layer6_outputs[424] = ~(layer5_outputs[4106]) | (layer5_outputs[4099]);
    assign layer6_outputs[425] = ~(layer5_outputs[4792]);
    assign layer6_outputs[426] = (layer5_outputs[1696]) ^ (layer5_outputs[1320]);
    assign layer6_outputs[427] = (layer5_outputs[4675]) | (layer5_outputs[5014]);
    assign layer6_outputs[428] = layer5_outputs[4029];
    assign layer6_outputs[429] = ~((layer5_outputs[4052]) ^ (layer5_outputs[318]));
    assign layer6_outputs[430] = (layer5_outputs[719]) & ~(layer5_outputs[4303]);
    assign layer6_outputs[431] = (layer5_outputs[4095]) & (layer5_outputs[4414]);
    assign layer6_outputs[432] = ~((layer5_outputs[5001]) & (layer5_outputs[4987]));
    assign layer6_outputs[433] = ~((layer5_outputs[4782]) & (layer5_outputs[2975]));
    assign layer6_outputs[434] = layer5_outputs[4052];
    assign layer6_outputs[435] = (layer5_outputs[1232]) & ~(layer5_outputs[946]);
    assign layer6_outputs[436] = ~(layer5_outputs[246]);
    assign layer6_outputs[437] = layer5_outputs[100];
    assign layer6_outputs[438] = layer5_outputs[2347];
    assign layer6_outputs[439] = ~(layer5_outputs[652]) | (layer5_outputs[4391]);
    assign layer6_outputs[440] = (layer5_outputs[4820]) & (layer5_outputs[4585]);
    assign layer6_outputs[441] = (layer5_outputs[972]) & ~(layer5_outputs[5117]);
    assign layer6_outputs[442] = layer5_outputs[4461];
    assign layer6_outputs[443] = layer5_outputs[2330];
    assign layer6_outputs[444] = ~(layer5_outputs[234]);
    assign layer6_outputs[445] = (layer5_outputs[3609]) & ~(layer5_outputs[2604]);
    assign layer6_outputs[446] = layer5_outputs[4161];
    assign layer6_outputs[447] = layer5_outputs[4143];
    assign layer6_outputs[448] = layer5_outputs[3409];
    assign layer6_outputs[449] = (layer5_outputs[2993]) & ~(layer5_outputs[2317]);
    assign layer6_outputs[450] = layer5_outputs[4429];
    assign layer6_outputs[451] = layer5_outputs[2929];
    assign layer6_outputs[452] = layer5_outputs[4832];
    assign layer6_outputs[453] = layer5_outputs[2867];
    assign layer6_outputs[454] = ~(layer5_outputs[2967]);
    assign layer6_outputs[455] = ~(layer5_outputs[4812]);
    assign layer6_outputs[456] = ~((layer5_outputs[2006]) ^ (layer5_outputs[2580]));
    assign layer6_outputs[457] = (layer5_outputs[4878]) & ~(layer5_outputs[839]);
    assign layer6_outputs[458] = (layer5_outputs[102]) ^ (layer5_outputs[3875]);
    assign layer6_outputs[459] = ~(layer5_outputs[1070]);
    assign layer6_outputs[460] = layer5_outputs[3043];
    assign layer6_outputs[461] = ~(layer5_outputs[868]);
    assign layer6_outputs[462] = (layer5_outputs[530]) ^ (layer5_outputs[4987]);
    assign layer6_outputs[463] = ~(layer5_outputs[990]) | (layer5_outputs[604]);
    assign layer6_outputs[464] = layer5_outputs[3361];
    assign layer6_outputs[465] = layer5_outputs[2137];
    assign layer6_outputs[466] = ~(layer5_outputs[3907]);
    assign layer6_outputs[467] = ~(layer5_outputs[1008]);
    assign layer6_outputs[468] = layer5_outputs[2576];
    assign layer6_outputs[469] = layer5_outputs[3697];
    assign layer6_outputs[470] = ~(layer5_outputs[613]);
    assign layer6_outputs[471] = ~(layer5_outputs[3195]);
    assign layer6_outputs[472] = ~(layer5_outputs[1873]);
    assign layer6_outputs[473] = layer5_outputs[1226];
    assign layer6_outputs[474] = (layer5_outputs[3897]) & ~(layer5_outputs[5055]);
    assign layer6_outputs[475] = layer5_outputs[1284];
    assign layer6_outputs[476] = layer5_outputs[803];
    assign layer6_outputs[477] = ~(layer5_outputs[2763]) | (layer5_outputs[332]);
    assign layer6_outputs[478] = ~(layer5_outputs[877]);
    assign layer6_outputs[479] = ~(layer5_outputs[3138]);
    assign layer6_outputs[480] = ~(layer5_outputs[1663]);
    assign layer6_outputs[481] = ~(layer5_outputs[681]) | (layer5_outputs[4674]);
    assign layer6_outputs[482] = ~(layer5_outputs[3934]) | (layer5_outputs[590]);
    assign layer6_outputs[483] = layer5_outputs[4314];
    assign layer6_outputs[484] = layer5_outputs[4873];
    assign layer6_outputs[485] = (layer5_outputs[4782]) ^ (layer5_outputs[5101]);
    assign layer6_outputs[486] = (layer5_outputs[827]) | (layer5_outputs[3028]);
    assign layer6_outputs[487] = layer5_outputs[42];
    assign layer6_outputs[488] = layer5_outputs[671];
    assign layer6_outputs[489] = ~(layer5_outputs[1163]) | (layer5_outputs[2122]);
    assign layer6_outputs[490] = ~((layer5_outputs[2366]) ^ (layer5_outputs[1648]));
    assign layer6_outputs[491] = layer5_outputs[129];
    assign layer6_outputs[492] = layer5_outputs[4517];
    assign layer6_outputs[493] = layer5_outputs[4872];
    assign layer6_outputs[494] = layer5_outputs[3331];
    assign layer6_outputs[495] = (layer5_outputs[1623]) | (layer5_outputs[3719]);
    assign layer6_outputs[496] = layer5_outputs[3522];
    assign layer6_outputs[497] = ~((layer5_outputs[4731]) | (layer5_outputs[2947]));
    assign layer6_outputs[498] = layer5_outputs[3238];
    assign layer6_outputs[499] = ~(layer5_outputs[4619]) | (layer5_outputs[4716]);
    assign layer6_outputs[500] = (layer5_outputs[1620]) | (layer5_outputs[2385]);
    assign layer6_outputs[501] = ~(layer5_outputs[736]) | (layer5_outputs[931]);
    assign layer6_outputs[502] = ~(layer5_outputs[4691]);
    assign layer6_outputs[503] = ~((layer5_outputs[2714]) & (layer5_outputs[423]));
    assign layer6_outputs[504] = (layer5_outputs[1025]) ^ (layer5_outputs[3019]);
    assign layer6_outputs[505] = layer5_outputs[5097];
    assign layer6_outputs[506] = ~(layer5_outputs[4632]);
    assign layer6_outputs[507] = layer5_outputs[3253];
    assign layer6_outputs[508] = ~((layer5_outputs[334]) ^ (layer5_outputs[2217]));
    assign layer6_outputs[509] = ~(layer5_outputs[1213]);
    assign layer6_outputs[510] = layer5_outputs[4593];
    assign layer6_outputs[511] = ~(layer5_outputs[3542]);
    assign layer6_outputs[512] = (layer5_outputs[1211]) ^ (layer5_outputs[2737]);
    assign layer6_outputs[513] = (layer5_outputs[3930]) & (layer5_outputs[2768]);
    assign layer6_outputs[514] = ~(layer5_outputs[757]);
    assign layer6_outputs[515] = ~((layer5_outputs[474]) & (layer5_outputs[3189]));
    assign layer6_outputs[516] = ~(layer5_outputs[1911]);
    assign layer6_outputs[517] = (layer5_outputs[1904]) & ~(layer5_outputs[781]);
    assign layer6_outputs[518] = (layer5_outputs[4755]) & (layer5_outputs[9]);
    assign layer6_outputs[519] = ~(layer5_outputs[1760]);
    assign layer6_outputs[520] = ~(layer5_outputs[4670]) | (layer5_outputs[4888]);
    assign layer6_outputs[521] = ~(layer5_outputs[428]);
    assign layer6_outputs[522] = layer5_outputs[1909];
    assign layer6_outputs[523] = (layer5_outputs[2493]) ^ (layer5_outputs[3188]);
    assign layer6_outputs[524] = layer5_outputs[1806];
    assign layer6_outputs[525] = ~(layer5_outputs[1982]) | (layer5_outputs[3004]);
    assign layer6_outputs[526] = ~((layer5_outputs[4830]) ^ (layer5_outputs[2941]));
    assign layer6_outputs[527] = ~((layer5_outputs[4129]) ^ (layer5_outputs[2296]));
    assign layer6_outputs[528] = layer5_outputs[4983];
    assign layer6_outputs[529] = ~(layer5_outputs[3365]);
    assign layer6_outputs[530] = ~(layer5_outputs[4605]);
    assign layer6_outputs[531] = ~((layer5_outputs[1974]) | (layer5_outputs[1059]));
    assign layer6_outputs[532] = ~(layer5_outputs[2297]) | (layer5_outputs[4427]);
    assign layer6_outputs[533] = (layer5_outputs[284]) ^ (layer5_outputs[3299]);
    assign layer6_outputs[534] = ~(layer5_outputs[3873]);
    assign layer6_outputs[535] = ~(layer5_outputs[4695]);
    assign layer6_outputs[536] = layer5_outputs[4201];
    assign layer6_outputs[537] = layer5_outputs[5098];
    assign layer6_outputs[538] = (layer5_outputs[4150]) & ~(layer5_outputs[2691]);
    assign layer6_outputs[539] = ~(layer5_outputs[4166]) | (layer5_outputs[270]);
    assign layer6_outputs[540] = ~(layer5_outputs[327]) | (layer5_outputs[5088]);
    assign layer6_outputs[541] = ~(layer5_outputs[2322]);
    assign layer6_outputs[542] = layer5_outputs[510];
    assign layer6_outputs[543] = ~(layer5_outputs[968]);
    assign layer6_outputs[544] = ~(layer5_outputs[5043]);
    assign layer6_outputs[545] = layer5_outputs[2809];
    assign layer6_outputs[546] = layer5_outputs[878];
    assign layer6_outputs[547] = (layer5_outputs[1626]) & ~(layer5_outputs[722]);
    assign layer6_outputs[548] = ~((layer5_outputs[1539]) ^ (layer5_outputs[3658]));
    assign layer6_outputs[549] = ~(layer5_outputs[4600]);
    assign layer6_outputs[550] = ~((layer5_outputs[3628]) ^ (layer5_outputs[1705]));
    assign layer6_outputs[551] = (layer5_outputs[1713]) & (layer5_outputs[4564]);
    assign layer6_outputs[552] = (layer5_outputs[3423]) & (layer5_outputs[1895]);
    assign layer6_outputs[553] = layer5_outputs[3674];
    assign layer6_outputs[554] = ~(layer5_outputs[876]);
    assign layer6_outputs[555] = layer5_outputs[3874];
    assign layer6_outputs[556] = ~(layer5_outputs[1632]);
    assign layer6_outputs[557] = layer5_outputs[3671];
    assign layer6_outputs[558] = ~((layer5_outputs[4394]) ^ (layer5_outputs[3777]));
    assign layer6_outputs[559] = ~((layer5_outputs[644]) ^ (layer5_outputs[2526]));
    assign layer6_outputs[560] = ~(layer5_outputs[1564]) | (layer5_outputs[1240]);
    assign layer6_outputs[561] = layer5_outputs[3124];
    assign layer6_outputs[562] = layer5_outputs[4606];
    assign layer6_outputs[563] = ~((layer5_outputs[2539]) ^ (layer5_outputs[3549]));
    assign layer6_outputs[564] = ~((layer5_outputs[3474]) ^ (layer5_outputs[2048]));
    assign layer6_outputs[565] = layer5_outputs[3342];
    assign layer6_outputs[566] = ~(layer5_outputs[4037]);
    assign layer6_outputs[567] = ~(layer5_outputs[2923]);
    assign layer6_outputs[568] = ~(layer5_outputs[2855]) | (layer5_outputs[835]);
    assign layer6_outputs[569] = ~(layer5_outputs[3117]) | (layer5_outputs[3798]);
    assign layer6_outputs[570] = ~(layer5_outputs[1834]);
    assign layer6_outputs[571] = ~(layer5_outputs[3290]);
    assign layer6_outputs[572] = ~(layer5_outputs[4910]);
    assign layer6_outputs[573] = layer5_outputs[3517];
    assign layer6_outputs[574] = ~(layer5_outputs[40]) | (layer5_outputs[1757]);
    assign layer6_outputs[575] = ~(layer5_outputs[968]) | (layer5_outputs[4594]);
    assign layer6_outputs[576] = layer5_outputs[2128];
    assign layer6_outputs[577] = (layer5_outputs[3606]) ^ (layer5_outputs[3529]);
    assign layer6_outputs[578] = ~((layer5_outputs[6]) | (layer5_outputs[3518]));
    assign layer6_outputs[579] = ~(layer5_outputs[3186]) | (layer5_outputs[3181]);
    assign layer6_outputs[580] = layer5_outputs[4228];
    assign layer6_outputs[581] = layer5_outputs[4825];
    assign layer6_outputs[582] = ~((layer5_outputs[4393]) | (layer5_outputs[3057]));
    assign layer6_outputs[583] = ~((layer5_outputs[2054]) | (layer5_outputs[3039]));
    assign layer6_outputs[584] = (layer5_outputs[4415]) | (layer5_outputs[2381]);
    assign layer6_outputs[585] = ~(layer5_outputs[1290]) | (layer5_outputs[4250]);
    assign layer6_outputs[586] = layer5_outputs[3288];
    assign layer6_outputs[587] = (layer5_outputs[3104]) | (layer5_outputs[716]);
    assign layer6_outputs[588] = ~(layer5_outputs[3151]);
    assign layer6_outputs[589] = layer5_outputs[3661];
    assign layer6_outputs[590] = (layer5_outputs[3823]) & ~(layer5_outputs[2408]);
    assign layer6_outputs[591] = ~(layer5_outputs[1032]);
    assign layer6_outputs[592] = ~(layer5_outputs[3874]);
    assign layer6_outputs[593] = ~((layer5_outputs[850]) ^ (layer5_outputs[4975]));
    assign layer6_outputs[594] = ~(layer5_outputs[3982]);
    assign layer6_outputs[595] = ~(layer5_outputs[4303]) | (layer5_outputs[1900]);
    assign layer6_outputs[596] = layer5_outputs[258];
    assign layer6_outputs[597] = layer5_outputs[4609];
    assign layer6_outputs[598] = (layer5_outputs[5050]) | (layer5_outputs[176]);
    assign layer6_outputs[599] = layer5_outputs[4800];
    assign layer6_outputs[600] = ~(layer5_outputs[2664]);
    assign layer6_outputs[601] = ~(layer5_outputs[3634]);
    assign layer6_outputs[602] = layer5_outputs[4413];
    assign layer6_outputs[603] = layer5_outputs[4410];
    assign layer6_outputs[604] = ~(layer5_outputs[1833]);
    assign layer6_outputs[605] = layer5_outputs[3085];
    assign layer6_outputs[606] = ~(layer5_outputs[1842]);
    assign layer6_outputs[607] = (layer5_outputs[2578]) ^ (layer5_outputs[4861]);
    assign layer6_outputs[608] = layer5_outputs[421];
    assign layer6_outputs[609] = (layer5_outputs[1346]) & ~(layer5_outputs[1720]);
    assign layer6_outputs[610] = ~(layer5_outputs[4431]);
    assign layer6_outputs[611] = layer5_outputs[4641];
    assign layer6_outputs[612] = (layer5_outputs[1666]) ^ (layer5_outputs[1591]);
    assign layer6_outputs[613] = ~(layer5_outputs[1852]);
    assign layer6_outputs[614] = ~((layer5_outputs[4080]) ^ (layer5_outputs[4074]));
    assign layer6_outputs[615] = layer5_outputs[249];
    assign layer6_outputs[616] = (layer5_outputs[1662]) ^ (layer5_outputs[4404]);
    assign layer6_outputs[617] = ~(layer5_outputs[1926]) | (layer5_outputs[2568]);
    assign layer6_outputs[618] = layer5_outputs[2067];
    assign layer6_outputs[619] = ~(layer5_outputs[5]) | (layer5_outputs[4039]);
    assign layer6_outputs[620] = layer5_outputs[2863];
    assign layer6_outputs[621] = layer5_outputs[4417];
    assign layer6_outputs[622] = ~((layer5_outputs[77]) & (layer5_outputs[3905]));
    assign layer6_outputs[623] = ~(layer5_outputs[4824]);
    assign layer6_outputs[624] = ~(layer5_outputs[4808]);
    assign layer6_outputs[625] = ~(layer5_outputs[3788]);
    assign layer6_outputs[626] = ~(layer5_outputs[548]) | (layer5_outputs[2777]);
    assign layer6_outputs[627] = layer5_outputs[3644];
    assign layer6_outputs[628] = ~(layer5_outputs[760]) | (layer5_outputs[3682]);
    assign layer6_outputs[629] = (layer5_outputs[1190]) & (layer5_outputs[3388]);
    assign layer6_outputs[630] = (layer5_outputs[2903]) & ~(layer5_outputs[4431]);
    assign layer6_outputs[631] = ~((layer5_outputs[3494]) | (layer5_outputs[3401]));
    assign layer6_outputs[632] = ~(layer5_outputs[2161]);
    assign layer6_outputs[633] = ~(layer5_outputs[4176]);
    assign layer6_outputs[634] = layer5_outputs[3137];
    assign layer6_outputs[635] = (layer5_outputs[1458]) & (layer5_outputs[3038]);
    assign layer6_outputs[636] = layer5_outputs[4459];
    assign layer6_outputs[637] = layer5_outputs[3654];
    assign layer6_outputs[638] = (layer5_outputs[2865]) & (layer5_outputs[2399]);
    assign layer6_outputs[639] = (layer5_outputs[2667]) & ~(layer5_outputs[3123]);
    assign layer6_outputs[640] = (layer5_outputs[4736]) | (layer5_outputs[1678]);
    assign layer6_outputs[641] = ~(layer5_outputs[2979]);
    assign layer6_outputs[642] = layer5_outputs[4535];
    assign layer6_outputs[643] = ~(layer5_outputs[4862]);
    assign layer6_outputs[644] = ~((layer5_outputs[2093]) | (layer5_outputs[2497]));
    assign layer6_outputs[645] = ~(layer5_outputs[1435]);
    assign layer6_outputs[646] = ~(layer5_outputs[592]);
    assign layer6_outputs[647] = ~(layer5_outputs[1966]);
    assign layer6_outputs[648] = ~(layer5_outputs[1319]) | (layer5_outputs[525]);
    assign layer6_outputs[649] = 1'b0;
    assign layer6_outputs[650] = ~(layer5_outputs[3734]);
    assign layer6_outputs[651] = ~((layer5_outputs[307]) | (layer5_outputs[883]));
    assign layer6_outputs[652] = ~((layer5_outputs[2050]) ^ (layer5_outputs[1928]));
    assign layer6_outputs[653] = layer5_outputs[2051];
    assign layer6_outputs[654] = ~(layer5_outputs[2038]);
    assign layer6_outputs[655] = ~(layer5_outputs[1932]);
    assign layer6_outputs[656] = layer5_outputs[108];
    assign layer6_outputs[657] = ~(layer5_outputs[459]);
    assign layer6_outputs[658] = layer5_outputs[3999];
    assign layer6_outputs[659] = layer5_outputs[1695];
    assign layer6_outputs[660] = (layer5_outputs[3582]) & ~(layer5_outputs[345]);
    assign layer6_outputs[661] = 1'b1;
    assign layer6_outputs[662] = ~(layer5_outputs[4504]);
    assign layer6_outputs[663] = ~(layer5_outputs[3942]) | (layer5_outputs[2091]);
    assign layer6_outputs[664] = (layer5_outputs[685]) ^ (layer5_outputs[1738]);
    assign layer6_outputs[665] = layer5_outputs[3737];
    assign layer6_outputs[666] = layer5_outputs[2814];
    assign layer6_outputs[667] = (layer5_outputs[2799]) ^ (layer5_outputs[1836]);
    assign layer6_outputs[668] = layer5_outputs[142];
    assign layer6_outputs[669] = ~((layer5_outputs[4005]) ^ (layer5_outputs[3742]));
    assign layer6_outputs[670] = (layer5_outputs[3853]) ^ (layer5_outputs[169]);
    assign layer6_outputs[671] = ~((layer5_outputs[4256]) | (layer5_outputs[936]));
    assign layer6_outputs[672] = (layer5_outputs[3597]) & ~(layer5_outputs[3190]);
    assign layer6_outputs[673] = layer5_outputs[2764];
    assign layer6_outputs[674] = ~((layer5_outputs[3078]) & (layer5_outputs[737]));
    assign layer6_outputs[675] = layer5_outputs[4216];
    assign layer6_outputs[676] = ~(layer5_outputs[529]);
    assign layer6_outputs[677] = (layer5_outputs[729]) & (layer5_outputs[2181]);
    assign layer6_outputs[678] = ~((layer5_outputs[3388]) | (layer5_outputs[4367]));
    assign layer6_outputs[679] = ~(layer5_outputs[4141]);
    assign layer6_outputs[680] = layer5_outputs[5094];
    assign layer6_outputs[681] = ~((layer5_outputs[4218]) ^ (layer5_outputs[1509]));
    assign layer6_outputs[682] = (layer5_outputs[2109]) & ~(layer5_outputs[281]);
    assign layer6_outputs[683] = 1'b0;
    assign layer6_outputs[684] = ~(layer5_outputs[4681]);
    assign layer6_outputs[685] = (layer5_outputs[2266]) & ~(layer5_outputs[2542]);
    assign layer6_outputs[686] = layer5_outputs[457];
    assign layer6_outputs[687] = ~(layer5_outputs[4719]) | (layer5_outputs[3364]);
    assign layer6_outputs[688] = ~(layer5_outputs[2472]) | (layer5_outputs[1370]);
    assign layer6_outputs[689] = (layer5_outputs[283]) & ~(layer5_outputs[3695]);
    assign layer6_outputs[690] = ~((layer5_outputs[3767]) ^ (layer5_outputs[3911]));
    assign layer6_outputs[691] = ~(layer5_outputs[3894]);
    assign layer6_outputs[692] = ~((layer5_outputs[4389]) | (layer5_outputs[1744]));
    assign layer6_outputs[693] = ~(layer5_outputs[1935]) | (layer5_outputs[5117]);
    assign layer6_outputs[694] = ~(layer5_outputs[636]);
    assign layer6_outputs[695] = layer5_outputs[4498];
    assign layer6_outputs[696] = 1'b1;
    assign layer6_outputs[697] = ~(layer5_outputs[1607]) | (layer5_outputs[843]);
    assign layer6_outputs[698] = ~(layer5_outputs[2111]) | (layer5_outputs[2142]);
    assign layer6_outputs[699] = ~(layer5_outputs[3970]);
    assign layer6_outputs[700] = ~((layer5_outputs[411]) | (layer5_outputs[982]));
    assign layer6_outputs[701] = ~(layer5_outputs[366]);
    assign layer6_outputs[702] = ~(layer5_outputs[3245]);
    assign layer6_outputs[703] = (layer5_outputs[1282]) | (layer5_outputs[5044]);
    assign layer6_outputs[704] = ~(layer5_outputs[749]);
    assign layer6_outputs[705] = (layer5_outputs[3676]) ^ (layer5_outputs[4556]);
    assign layer6_outputs[706] = layer5_outputs[3405];
    assign layer6_outputs[707] = (layer5_outputs[4323]) | (layer5_outputs[1398]);
    assign layer6_outputs[708] = layer5_outputs[3725];
    assign layer6_outputs[709] = layer5_outputs[4917];
    assign layer6_outputs[710] = ~(layer5_outputs[145]);
    assign layer6_outputs[711] = layer5_outputs[4328];
    assign layer6_outputs[712] = ~(layer5_outputs[4648]) | (layer5_outputs[3614]);
    assign layer6_outputs[713] = (layer5_outputs[3297]) ^ (layer5_outputs[2314]);
    assign layer6_outputs[714] = (layer5_outputs[1535]) & ~(layer5_outputs[2219]);
    assign layer6_outputs[715] = layer5_outputs[100];
    assign layer6_outputs[716] = ~(layer5_outputs[1032]);
    assign layer6_outputs[717] = layer5_outputs[4094];
    assign layer6_outputs[718] = layer5_outputs[1803];
    assign layer6_outputs[719] = (layer5_outputs[2400]) | (layer5_outputs[3616]);
    assign layer6_outputs[720] = ~(layer5_outputs[3948]);
    assign layer6_outputs[721] = layer5_outputs[1126];
    assign layer6_outputs[722] = ~(layer5_outputs[3573]);
    assign layer6_outputs[723] = ~((layer5_outputs[3326]) ^ (layer5_outputs[4588]));
    assign layer6_outputs[724] = ~((layer5_outputs[818]) ^ (layer5_outputs[4267]));
    assign layer6_outputs[725] = ~(layer5_outputs[2957]);
    assign layer6_outputs[726] = ~((layer5_outputs[2527]) ^ (layer5_outputs[1581]));
    assign layer6_outputs[727] = ~(layer5_outputs[3489]) | (layer5_outputs[3592]);
    assign layer6_outputs[728] = ~(layer5_outputs[3653]);
    assign layer6_outputs[729] = layer5_outputs[3988];
    assign layer6_outputs[730] = (layer5_outputs[3964]) | (layer5_outputs[3849]);
    assign layer6_outputs[731] = ~(layer5_outputs[1115]);
    assign layer6_outputs[732] = ~(layer5_outputs[3935]);
    assign layer6_outputs[733] = layer5_outputs[709];
    assign layer6_outputs[734] = ~(layer5_outputs[439]);
    assign layer6_outputs[735] = (layer5_outputs[1494]) & ~(layer5_outputs[2968]);
    assign layer6_outputs[736] = layer5_outputs[2090];
    assign layer6_outputs[737] = 1'b1;
    assign layer6_outputs[738] = layer5_outputs[578];
    assign layer6_outputs[739] = ~((layer5_outputs[1463]) & (layer5_outputs[3625]));
    assign layer6_outputs[740] = ~(layer5_outputs[2276]) | (layer5_outputs[2237]);
    assign layer6_outputs[741] = ~((layer5_outputs[2275]) | (layer5_outputs[2125]));
    assign layer6_outputs[742] = ~(layer5_outputs[2141]);
    assign layer6_outputs[743] = layer5_outputs[3578];
    assign layer6_outputs[744] = ~(layer5_outputs[854]);
    assign layer6_outputs[745] = ~(layer5_outputs[1516]) | (layer5_outputs[3131]);
    assign layer6_outputs[746] = (layer5_outputs[1905]) | (layer5_outputs[3979]);
    assign layer6_outputs[747] = ~((layer5_outputs[1432]) | (layer5_outputs[2432]));
    assign layer6_outputs[748] = (layer5_outputs[3419]) ^ (layer5_outputs[3773]);
    assign layer6_outputs[749] = ~(layer5_outputs[674]);
    assign layer6_outputs[750] = ~(layer5_outputs[3118]);
    assign layer6_outputs[751] = 1'b0;
    assign layer6_outputs[752] = (layer5_outputs[2447]) & (layer5_outputs[4222]);
    assign layer6_outputs[753] = ~((layer5_outputs[1299]) | (layer5_outputs[2666]));
    assign layer6_outputs[754] = layer5_outputs[4091];
    assign layer6_outputs[755] = 1'b1;
    assign layer6_outputs[756] = ~(layer5_outputs[4209]) | (layer5_outputs[3632]);
    assign layer6_outputs[757] = layer5_outputs[2478];
    assign layer6_outputs[758] = ~(layer5_outputs[2483]);
    assign layer6_outputs[759] = ~(layer5_outputs[1646]);
    assign layer6_outputs[760] = ~(layer5_outputs[3528]);
    assign layer6_outputs[761] = ~((layer5_outputs[87]) | (layer5_outputs[4737]));
    assign layer6_outputs[762] = ~((layer5_outputs[4504]) & (layer5_outputs[187]));
    assign layer6_outputs[763] = layer5_outputs[1645];
    assign layer6_outputs[764] = layer5_outputs[5021];
    assign layer6_outputs[765] = ~((layer5_outputs[955]) ^ (layer5_outputs[483]));
    assign layer6_outputs[766] = layer5_outputs[4252];
    assign layer6_outputs[767] = ~(layer5_outputs[2816]);
    assign layer6_outputs[768] = ~(layer5_outputs[1332]);
    assign layer6_outputs[769] = (layer5_outputs[755]) & (layer5_outputs[3551]);
    assign layer6_outputs[770] = layer5_outputs[4278];
    assign layer6_outputs[771] = (layer5_outputs[28]) ^ (layer5_outputs[1020]);
    assign layer6_outputs[772] = ~(layer5_outputs[2899]);
    assign layer6_outputs[773] = (layer5_outputs[5044]) | (layer5_outputs[659]);
    assign layer6_outputs[774] = ~((layer5_outputs[2725]) & (layer5_outputs[4829]));
    assign layer6_outputs[775] = (layer5_outputs[4180]) | (layer5_outputs[5047]);
    assign layer6_outputs[776] = ~(layer5_outputs[191]) | (layer5_outputs[1018]);
    assign layer6_outputs[777] = ~(layer5_outputs[1400]);
    assign layer6_outputs[778] = ~(layer5_outputs[3428]);
    assign layer6_outputs[779] = ~(layer5_outputs[2952]);
    assign layer6_outputs[780] = (layer5_outputs[3274]) & ~(layer5_outputs[1352]);
    assign layer6_outputs[781] = layer5_outputs[4392];
    assign layer6_outputs[782] = (layer5_outputs[3565]) ^ (layer5_outputs[1452]);
    assign layer6_outputs[783] = ~(layer5_outputs[915]);
    assign layer6_outputs[784] = ~(layer5_outputs[2822]) | (layer5_outputs[471]);
    assign layer6_outputs[785] = ~(layer5_outputs[2337]);
    assign layer6_outputs[786] = layer5_outputs[2003];
    assign layer6_outputs[787] = layer5_outputs[2322];
    assign layer6_outputs[788] = ~(layer5_outputs[75]) | (layer5_outputs[4960]);
    assign layer6_outputs[789] = layer5_outputs[1463];
    assign layer6_outputs[790] = layer5_outputs[4877];
    assign layer6_outputs[791] = ~(layer5_outputs[2910]);
    assign layer6_outputs[792] = (layer5_outputs[2566]) ^ (layer5_outputs[3467]);
    assign layer6_outputs[793] = ~(layer5_outputs[48]);
    assign layer6_outputs[794] = ~(layer5_outputs[1568]) | (layer5_outputs[2308]);
    assign layer6_outputs[795] = ~(layer5_outputs[836]);
    assign layer6_outputs[796] = ~((layer5_outputs[3804]) ^ (layer5_outputs[1575]));
    assign layer6_outputs[797] = ~(layer5_outputs[4466]);
    assign layer6_outputs[798] = layer5_outputs[4990];
    assign layer6_outputs[799] = ~(layer5_outputs[2794]);
    assign layer6_outputs[800] = ~(layer5_outputs[875]) | (layer5_outputs[4779]);
    assign layer6_outputs[801] = (layer5_outputs[4932]) | (layer5_outputs[4405]);
    assign layer6_outputs[802] = (layer5_outputs[4144]) & ~(layer5_outputs[733]);
    assign layer6_outputs[803] = ~((layer5_outputs[0]) | (layer5_outputs[2077]));
    assign layer6_outputs[804] = layer5_outputs[1013];
    assign layer6_outputs[805] = ~(layer5_outputs[3594]);
    assign layer6_outputs[806] = ~(layer5_outputs[4797]);
    assign layer6_outputs[807] = ~((layer5_outputs[2576]) & (layer5_outputs[2711]));
    assign layer6_outputs[808] = ~(layer5_outputs[2156]);
    assign layer6_outputs[809] = ~(layer5_outputs[4340]);
    assign layer6_outputs[810] = (layer5_outputs[3872]) & ~(layer5_outputs[3367]);
    assign layer6_outputs[811] = ~(layer5_outputs[4831]);
    assign layer6_outputs[812] = (layer5_outputs[1429]) ^ (layer5_outputs[413]);
    assign layer6_outputs[813] = ~(layer5_outputs[2194]);
    assign layer6_outputs[814] = ~((layer5_outputs[4893]) & (layer5_outputs[4647]));
    assign layer6_outputs[815] = ~(layer5_outputs[137]);
    assign layer6_outputs[816] = ~(layer5_outputs[5035]);
    assign layer6_outputs[817] = ~(layer5_outputs[4630]);
    assign layer6_outputs[818] = ~(layer5_outputs[3321]) | (layer5_outputs[2394]);
    assign layer6_outputs[819] = ~(layer5_outputs[4520]);
    assign layer6_outputs[820] = layer5_outputs[467];
    assign layer6_outputs[821] = ~((layer5_outputs[4074]) & (layer5_outputs[1291]));
    assign layer6_outputs[822] = (layer5_outputs[2191]) & ~(layer5_outputs[1413]);
    assign layer6_outputs[823] = ~(layer5_outputs[3294]) | (layer5_outputs[1028]);
    assign layer6_outputs[824] = (layer5_outputs[3543]) & ~(layer5_outputs[2949]);
    assign layer6_outputs[825] = (layer5_outputs[2099]) | (layer5_outputs[2097]);
    assign layer6_outputs[826] = layer5_outputs[1847];
    assign layer6_outputs[827] = ~(layer5_outputs[2168]);
    assign layer6_outputs[828] = ~((layer5_outputs[2698]) ^ (layer5_outputs[2756]));
    assign layer6_outputs[829] = layer5_outputs[3998];
    assign layer6_outputs[830] = ~((layer5_outputs[369]) & (layer5_outputs[1917]));
    assign layer6_outputs[831] = layer5_outputs[1818];
    assign layer6_outputs[832] = ~(layer5_outputs[4034]);
    assign layer6_outputs[833] = (layer5_outputs[349]) & ~(layer5_outputs[31]);
    assign layer6_outputs[834] = ~((layer5_outputs[4273]) ^ (layer5_outputs[140]));
    assign layer6_outputs[835] = ~(layer5_outputs[1697]);
    assign layer6_outputs[836] = ~(layer5_outputs[4130]) | (layer5_outputs[1570]);
    assign layer6_outputs[837] = ~(layer5_outputs[1746]) | (layer5_outputs[2974]);
    assign layer6_outputs[838] = layer5_outputs[1525];
    assign layer6_outputs[839] = (layer5_outputs[4037]) ^ (layer5_outputs[437]);
    assign layer6_outputs[840] = ~(layer5_outputs[4495]);
    assign layer6_outputs[841] = ~(layer5_outputs[3366]);
    assign layer6_outputs[842] = ~(layer5_outputs[2555]);
    assign layer6_outputs[843] = (layer5_outputs[2741]) ^ (layer5_outputs[1088]);
    assign layer6_outputs[844] = (layer5_outputs[3259]) | (layer5_outputs[2595]);
    assign layer6_outputs[845] = (layer5_outputs[3877]) ^ (layer5_outputs[2149]);
    assign layer6_outputs[846] = ~(layer5_outputs[1431]);
    assign layer6_outputs[847] = ~(layer5_outputs[800]);
    assign layer6_outputs[848] = (layer5_outputs[3169]) ^ (layer5_outputs[4364]);
    assign layer6_outputs[849] = (layer5_outputs[3232]) | (layer5_outputs[2751]);
    assign layer6_outputs[850] = ~((layer5_outputs[3370]) | (layer5_outputs[2026]));
    assign layer6_outputs[851] = ~(layer5_outputs[762]) | (layer5_outputs[82]);
    assign layer6_outputs[852] = (layer5_outputs[4974]) & ~(layer5_outputs[3798]);
    assign layer6_outputs[853] = ~(layer5_outputs[3330]) | (layer5_outputs[977]);
    assign layer6_outputs[854] = ~(layer5_outputs[2024]) | (layer5_outputs[461]);
    assign layer6_outputs[855] = ~(layer5_outputs[4563]);
    assign layer6_outputs[856] = layer5_outputs[2986];
    assign layer6_outputs[857] = ~(layer5_outputs[3588]) | (layer5_outputs[4576]);
    assign layer6_outputs[858] = layer5_outputs[418];
    assign layer6_outputs[859] = ~((layer5_outputs[1694]) ^ (layer5_outputs[751]));
    assign layer6_outputs[860] = (layer5_outputs[292]) ^ (layer5_outputs[3248]);
    assign layer6_outputs[861] = ~(layer5_outputs[4598]);
    assign layer6_outputs[862] = layer5_outputs[2519];
    assign layer6_outputs[863] = 1'b0;
    assign layer6_outputs[864] = (layer5_outputs[2075]) & (layer5_outputs[817]);
    assign layer6_outputs[865] = ~(layer5_outputs[2479]);
    assign layer6_outputs[866] = (layer5_outputs[3115]) ^ (layer5_outputs[2375]);
    assign layer6_outputs[867] = ~(layer5_outputs[3309]) | (layer5_outputs[1667]);
    assign layer6_outputs[868] = (layer5_outputs[2405]) | (layer5_outputs[3617]);
    assign layer6_outputs[869] = ~(layer5_outputs[4000]);
    assign layer6_outputs[870] = ~(layer5_outputs[4435]);
    assign layer6_outputs[871] = (layer5_outputs[2653]) & (layer5_outputs[2759]);
    assign layer6_outputs[872] = ~(layer5_outputs[3010]);
    assign layer6_outputs[873] = ~((layer5_outputs[3807]) | (layer5_outputs[2341]));
    assign layer6_outputs[874] = 1'b1;
    assign layer6_outputs[875] = ~(layer5_outputs[2301]);
    assign layer6_outputs[876] = layer5_outputs[2466];
    assign layer6_outputs[877] = layer5_outputs[4600];
    assign layer6_outputs[878] = layer5_outputs[4312];
    assign layer6_outputs[879] = ~(layer5_outputs[3275]);
    assign layer6_outputs[880] = (layer5_outputs[2670]) ^ (layer5_outputs[1601]);
    assign layer6_outputs[881] = ~(layer5_outputs[2958]);
    assign layer6_outputs[882] = ~(layer5_outputs[1194]) | (layer5_outputs[4118]);
    assign layer6_outputs[883] = layer5_outputs[4460];
    assign layer6_outputs[884] = layer5_outputs[3878];
    assign layer6_outputs[885] = ~(layer5_outputs[1266]) | (layer5_outputs[4029]);
    assign layer6_outputs[886] = layer5_outputs[2115];
    assign layer6_outputs[887] = (layer5_outputs[576]) ^ (layer5_outputs[3183]);
    assign layer6_outputs[888] = ~(layer5_outputs[852]) | (layer5_outputs[4268]);
    assign layer6_outputs[889] = layer5_outputs[1790];
    assign layer6_outputs[890] = (layer5_outputs[4941]) & ~(layer5_outputs[4234]);
    assign layer6_outputs[891] = layer5_outputs[3067];
    assign layer6_outputs[892] = ~(layer5_outputs[3700]) | (layer5_outputs[3197]);
    assign layer6_outputs[893] = (layer5_outputs[1596]) & ~(layer5_outputs[2199]);
    assign layer6_outputs[894] = (layer5_outputs[1964]) ^ (layer5_outputs[1384]);
    assign layer6_outputs[895] = layer5_outputs[4682];
    assign layer6_outputs[896] = (layer5_outputs[1172]) ^ (layer5_outputs[254]);
    assign layer6_outputs[897] = ~(layer5_outputs[3692]);
    assign layer6_outputs[898] = (layer5_outputs[1156]) | (layer5_outputs[3475]);
    assign layer6_outputs[899] = 1'b1;
    assign layer6_outputs[900] = layer5_outputs[658];
    assign layer6_outputs[901] = ~(layer5_outputs[2615]);
    assign layer6_outputs[902] = ~((layer5_outputs[1317]) | (layer5_outputs[1625]));
    assign layer6_outputs[903] = (layer5_outputs[4533]) & ~(layer5_outputs[1347]);
    assign layer6_outputs[904] = (layer5_outputs[830]) & ~(layer5_outputs[1083]);
    assign layer6_outputs[905] = layer5_outputs[5001];
    assign layer6_outputs[906] = layer5_outputs[1467];
    assign layer6_outputs[907] = 1'b0;
    assign layer6_outputs[908] = ~(layer5_outputs[1710]) | (layer5_outputs[4847]);
    assign layer6_outputs[909] = ~(layer5_outputs[4462]) | (layer5_outputs[670]);
    assign layer6_outputs[910] = ~(layer5_outputs[1654]) | (layer5_outputs[2841]);
    assign layer6_outputs[911] = (layer5_outputs[2174]) ^ (layer5_outputs[3956]);
    assign layer6_outputs[912] = layer5_outputs[3960];
    assign layer6_outputs[913] = 1'b1;
    assign layer6_outputs[914] = (layer5_outputs[2609]) | (layer5_outputs[4194]);
    assign layer6_outputs[915] = ~(layer5_outputs[1791]);
    assign layer6_outputs[916] = layer5_outputs[4169];
    assign layer6_outputs[917] = ~((layer5_outputs[1878]) ^ (layer5_outputs[734]));
    assign layer6_outputs[918] = (layer5_outputs[2891]) ^ (layer5_outputs[3553]);
    assign layer6_outputs[919] = (layer5_outputs[4143]) & (layer5_outputs[3241]);
    assign layer6_outputs[920] = (layer5_outputs[1649]) & (layer5_outputs[3247]);
    assign layer6_outputs[921] = ~(layer5_outputs[2403]);
    assign layer6_outputs[922] = ~((layer5_outputs[97]) ^ (layer5_outputs[1656]));
    assign layer6_outputs[923] = layer5_outputs[1866];
    assign layer6_outputs[924] = ~((layer5_outputs[3218]) ^ (layer5_outputs[1112]));
    assign layer6_outputs[925] = ~(layer5_outputs[3826]) | (layer5_outputs[2895]);
    assign layer6_outputs[926] = ~((layer5_outputs[408]) ^ (layer5_outputs[1971]));
    assign layer6_outputs[927] = ~(layer5_outputs[925]);
    assign layer6_outputs[928] = (layer5_outputs[4119]) ^ (layer5_outputs[3383]);
    assign layer6_outputs[929] = ~(layer5_outputs[4172]);
    assign layer6_outputs[930] = (layer5_outputs[3510]) ^ (layer5_outputs[3615]);
    assign layer6_outputs[931] = layer5_outputs[236];
    assign layer6_outputs[932] = (layer5_outputs[3906]) & (layer5_outputs[2393]);
    assign layer6_outputs[933] = ~((layer5_outputs[139]) | (layer5_outputs[1252]));
    assign layer6_outputs[934] = layer5_outputs[1232];
    assign layer6_outputs[935] = ~(layer5_outputs[3697]);
    assign layer6_outputs[936] = ~(layer5_outputs[1681]);
    assign layer6_outputs[937] = (layer5_outputs[1686]) & (layer5_outputs[1983]);
    assign layer6_outputs[938] = (layer5_outputs[4390]) | (layer5_outputs[2920]);
    assign layer6_outputs[939] = ~(layer5_outputs[3961]) | (layer5_outputs[4673]);
    assign layer6_outputs[940] = (layer5_outputs[2945]) ^ (layer5_outputs[306]);
    assign layer6_outputs[941] = ~(layer5_outputs[2161]);
    assign layer6_outputs[942] = ~(layer5_outputs[1553]) | (layer5_outputs[3110]);
    assign layer6_outputs[943] = ~(layer5_outputs[1984]) | (layer5_outputs[5083]);
    assign layer6_outputs[944] = layer5_outputs[5023];
    assign layer6_outputs[945] = ~(layer5_outputs[921]);
    assign layer6_outputs[946] = ~((layer5_outputs[3238]) ^ (layer5_outputs[736]));
    assign layer6_outputs[947] = ~(layer5_outputs[3550]);
    assign layer6_outputs[948] = (layer5_outputs[3991]) & ~(layer5_outputs[4662]);
    assign layer6_outputs[949] = layer5_outputs[1801];
    assign layer6_outputs[950] = ~(layer5_outputs[562]);
    assign layer6_outputs[951] = ~((layer5_outputs[2793]) ^ (layer5_outputs[2854]));
    assign layer6_outputs[952] = ~(layer5_outputs[4261]) | (layer5_outputs[569]);
    assign layer6_outputs[953] = ~(layer5_outputs[1822]);
    assign layer6_outputs[954] = ~(layer5_outputs[2292]) | (layer5_outputs[3695]);
    assign layer6_outputs[955] = layer5_outputs[2930];
    assign layer6_outputs[956] = ~(layer5_outputs[2185]) | (layer5_outputs[939]);
    assign layer6_outputs[957] = ~(layer5_outputs[765]);
    assign layer6_outputs[958] = ~(layer5_outputs[4085]) | (layer5_outputs[4738]);
    assign layer6_outputs[959] = (layer5_outputs[1437]) & (layer5_outputs[1710]);
    assign layer6_outputs[960] = ~((layer5_outputs[4696]) | (layer5_outputs[3359]));
    assign layer6_outputs[961] = layer5_outputs[1207];
    assign layer6_outputs[962] = ~(layer5_outputs[5022]);
    assign layer6_outputs[963] = ~(layer5_outputs[192]) | (layer5_outputs[189]);
    assign layer6_outputs[964] = ~(layer5_outputs[4055]);
    assign layer6_outputs[965] = (layer5_outputs[4225]) ^ (layer5_outputs[4059]);
    assign layer6_outputs[966] = ~(layer5_outputs[4924]);
    assign layer6_outputs[967] = ~(layer5_outputs[3547]) | (layer5_outputs[1246]);
    assign layer6_outputs[968] = (layer5_outputs[1001]) & (layer5_outputs[604]);
    assign layer6_outputs[969] = ~((layer5_outputs[3190]) ^ (layer5_outputs[1616]));
    assign layer6_outputs[970] = layer5_outputs[1752];
    assign layer6_outputs[971] = ~(layer5_outputs[931]) | (layer5_outputs[1272]);
    assign layer6_outputs[972] = layer5_outputs[4880];
    assign layer6_outputs[973] = layer5_outputs[4627];
    assign layer6_outputs[974] = ~(layer5_outputs[1519]);
    assign layer6_outputs[975] = layer5_outputs[1312];
    assign layer6_outputs[976] = ~(layer5_outputs[3613]);
    assign layer6_outputs[977] = ~(layer5_outputs[3125]) | (layer5_outputs[2982]);
    assign layer6_outputs[978] = ~(layer5_outputs[830]);
    assign layer6_outputs[979] = ~(layer5_outputs[3598]);
    assign layer6_outputs[980] = ~(layer5_outputs[2108]) | (layer5_outputs[79]);
    assign layer6_outputs[981] = ~((layer5_outputs[2312]) & (layer5_outputs[3040]));
    assign layer6_outputs[982] = ~(layer5_outputs[454]) | (layer5_outputs[981]);
    assign layer6_outputs[983] = (layer5_outputs[1791]) & ~(layer5_outputs[1745]);
    assign layer6_outputs[984] = ~(layer5_outputs[303]);
    assign layer6_outputs[985] = ~(layer5_outputs[3650]);
    assign layer6_outputs[986] = ~(layer5_outputs[4860]) | (layer5_outputs[795]);
    assign layer6_outputs[987] = (layer5_outputs[4730]) | (layer5_outputs[864]);
    assign layer6_outputs[988] = ~((layer5_outputs[2997]) ^ (layer5_outputs[392]));
    assign layer6_outputs[989] = (layer5_outputs[3964]) | (layer5_outputs[2113]);
    assign layer6_outputs[990] = layer5_outputs[2202];
    assign layer6_outputs[991] = ~(layer5_outputs[1678]);
    assign layer6_outputs[992] = layer5_outputs[1688];
    assign layer6_outputs[993] = ~(layer5_outputs[4907]);
    assign layer6_outputs[994] = ~(layer5_outputs[1595]) | (layer5_outputs[2900]);
    assign layer6_outputs[995] = layer5_outputs[2829];
    assign layer6_outputs[996] = (layer5_outputs[2963]) | (layer5_outputs[3937]);
    assign layer6_outputs[997] = ~((layer5_outputs[632]) | (layer5_outputs[4088]));
    assign layer6_outputs[998] = ~(layer5_outputs[3577]) | (layer5_outputs[2135]);
    assign layer6_outputs[999] = layer5_outputs[4995];
    assign layer6_outputs[1000] = ~(layer5_outputs[1308]) | (layer5_outputs[91]);
    assign layer6_outputs[1001] = ~(layer5_outputs[328]);
    assign layer6_outputs[1002] = ~(layer5_outputs[237]);
    assign layer6_outputs[1003] = layer5_outputs[2483];
    assign layer6_outputs[1004] = ~(layer5_outputs[4438]);
    assign layer6_outputs[1005] = ~(layer5_outputs[1164]);
    assign layer6_outputs[1006] = ~(layer5_outputs[2806]);
    assign layer6_outputs[1007] = ~(layer5_outputs[3017]) | (layer5_outputs[2934]);
    assign layer6_outputs[1008] = (layer5_outputs[4477]) & (layer5_outputs[933]);
    assign layer6_outputs[1009] = 1'b1;
    assign layer6_outputs[1010] = layer5_outputs[1782];
    assign layer6_outputs[1011] = layer5_outputs[5069];
    assign layer6_outputs[1012] = layer5_outputs[4870];
    assign layer6_outputs[1013] = ~((layer5_outputs[916]) & (layer5_outputs[348]));
    assign layer6_outputs[1014] = (layer5_outputs[477]) | (layer5_outputs[2510]);
    assign layer6_outputs[1015] = (layer5_outputs[1275]) ^ (layer5_outputs[2345]);
    assign layer6_outputs[1016] = layer5_outputs[4014];
    assign layer6_outputs[1017] = ~(layer5_outputs[4424]) | (layer5_outputs[278]);
    assign layer6_outputs[1018] = ~(layer5_outputs[1502]) | (layer5_outputs[5107]);
    assign layer6_outputs[1019] = ~(layer5_outputs[4594]);
    assign layer6_outputs[1020] = (layer5_outputs[1711]) & ~(layer5_outputs[2886]);
    assign layer6_outputs[1021] = (layer5_outputs[589]) & ~(layer5_outputs[1902]);
    assign layer6_outputs[1022] = ~(layer5_outputs[2370]);
    assign layer6_outputs[1023] = (layer5_outputs[86]) & ~(layer5_outputs[32]);
    assign layer6_outputs[1024] = ~(layer5_outputs[405]);
    assign layer6_outputs[1025] = layer5_outputs[4728];
    assign layer6_outputs[1026] = ~(layer5_outputs[3141]);
    assign layer6_outputs[1027] = (layer5_outputs[3739]) | (layer5_outputs[2804]);
    assign layer6_outputs[1028] = layer5_outputs[4127];
    assign layer6_outputs[1029] = (layer5_outputs[3519]) & (layer5_outputs[3466]);
    assign layer6_outputs[1030] = ~(layer5_outputs[2265]);
    assign layer6_outputs[1031] = (layer5_outputs[2078]) ^ (layer5_outputs[1781]);
    assign layer6_outputs[1032] = layer5_outputs[4974];
    assign layer6_outputs[1033] = layer5_outputs[1966];
    assign layer6_outputs[1034] = layer5_outputs[2389];
    assign layer6_outputs[1035] = ~(layer5_outputs[4444]);
    assign layer6_outputs[1036] = layer5_outputs[1860];
    assign layer6_outputs[1037] = 1'b0;
    assign layer6_outputs[1038] = ~((layer5_outputs[3501]) ^ (layer5_outputs[2953]));
    assign layer6_outputs[1039] = ~((layer5_outputs[1636]) & (layer5_outputs[2131]));
    assign layer6_outputs[1040] = layer5_outputs[3396];
    assign layer6_outputs[1041] = ~(layer5_outputs[1036]);
    assign layer6_outputs[1042] = layer5_outputs[438];
    assign layer6_outputs[1043] = layer5_outputs[4845];
    assign layer6_outputs[1044] = layer5_outputs[4812];
    assign layer6_outputs[1045] = ~(layer5_outputs[2744]);
    assign layer6_outputs[1046] = ~(layer5_outputs[2983]);
    assign layer6_outputs[1047] = layer5_outputs[1987];
    assign layer6_outputs[1048] = ~((layer5_outputs[2504]) ^ (layer5_outputs[3959]));
    assign layer6_outputs[1049] = ~(layer5_outputs[3148]);
    assign layer6_outputs[1050] = (layer5_outputs[4778]) ^ (layer5_outputs[4572]);
    assign layer6_outputs[1051] = ~(layer5_outputs[2304]);
    assign layer6_outputs[1052] = ~((layer5_outputs[3295]) ^ (layer5_outputs[2508]));
    assign layer6_outputs[1053] = ~(layer5_outputs[440]) | (layer5_outputs[4225]);
    assign layer6_outputs[1054] = layer5_outputs[1623];
    assign layer6_outputs[1055] = (layer5_outputs[4170]) ^ (layer5_outputs[4998]);
    assign layer6_outputs[1056] = ~(layer5_outputs[3327]);
    assign layer6_outputs[1057] = (layer5_outputs[3063]) ^ (layer5_outputs[4016]);
    assign layer6_outputs[1058] = ~(layer5_outputs[1125]);
    assign layer6_outputs[1059] = ~((layer5_outputs[2775]) | (layer5_outputs[4791]));
    assign layer6_outputs[1060] = ~(layer5_outputs[3503]) | (layer5_outputs[621]);
    assign layer6_outputs[1061] = layer5_outputs[1145];
    assign layer6_outputs[1062] = layer5_outputs[3360];
    assign layer6_outputs[1063] = (layer5_outputs[2254]) & ~(layer5_outputs[3627]);
    assign layer6_outputs[1064] = layer5_outputs[1358];
    assign layer6_outputs[1065] = (layer5_outputs[3884]) ^ (layer5_outputs[891]);
    assign layer6_outputs[1066] = ~(layer5_outputs[2443]);
    assign layer6_outputs[1067] = ~((layer5_outputs[600]) ^ (layer5_outputs[3532]));
    assign layer6_outputs[1068] = layer5_outputs[2299];
    assign layer6_outputs[1069] = ~((layer5_outputs[156]) | (layer5_outputs[4610]));
    assign layer6_outputs[1070] = ~((layer5_outputs[705]) & (layer5_outputs[3224]));
    assign layer6_outputs[1071] = ~(layer5_outputs[999]);
    assign layer6_outputs[1072] = ~(layer5_outputs[4045]);
    assign layer6_outputs[1073] = ~(layer5_outputs[3646]);
    assign layer6_outputs[1074] = layer5_outputs[4701];
    assign layer6_outputs[1075] = layer5_outputs[2018];
    assign layer6_outputs[1076] = 1'b0;
    assign layer6_outputs[1077] = ~((layer5_outputs[4626]) | (layer5_outputs[326]));
    assign layer6_outputs[1078] = layer5_outputs[4724];
    assign layer6_outputs[1079] = ~((layer5_outputs[4603]) & (layer5_outputs[4311]));
    assign layer6_outputs[1080] = ~(layer5_outputs[4909]);
    assign layer6_outputs[1081] = ~(layer5_outputs[2439]) | (layer5_outputs[2196]);
    assign layer6_outputs[1082] = ~(layer5_outputs[2922]);
    assign layer6_outputs[1083] = ~((layer5_outputs[3441]) | (layer5_outputs[1629]));
    assign layer6_outputs[1084] = ~(layer5_outputs[1260]) | (layer5_outputs[2478]);
    assign layer6_outputs[1085] = ~(layer5_outputs[811]);
    assign layer6_outputs[1086] = ~((layer5_outputs[3996]) ^ (layer5_outputs[2041]));
    assign layer6_outputs[1087] = ~(layer5_outputs[1730]);
    assign layer6_outputs[1088] = layer5_outputs[2324];
    assign layer6_outputs[1089] = layer5_outputs[1468];
    assign layer6_outputs[1090] = ~((layer5_outputs[1557]) & (layer5_outputs[4558]));
    assign layer6_outputs[1091] = layer5_outputs[545];
    assign layer6_outputs[1092] = ~((layer5_outputs[4657]) ^ (layer5_outputs[4200]));
    assign layer6_outputs[1093] = ~((layer5_outputs[1026]) & (layer5_outputs[1485]));
    assign layer6_outputs[1094] = (layer5_outputs[5002]) & ~(layer5_outputs[1567]);
    assign layer6_outputs[1095] = ~((layer5_outputs[4076]) ^ (layer5_outputs[846]));
    assign layer6_outputs[1096] = ~((layer5_outputs[2708]) ^ (layer5_outputs[4279]));
    assign layer6_outputs[1097] = (layer5_outputs[3730]) ^ (layer5_outputs[5037]);
    assign layer6_outputs[1098] = (layer5_outputs[1449]) & ~(layer5_outputs[2818]);
    assign layer6_outputs[1099] = ~(layer5_outputs[4809]);
    assign layer6_outputs[1100] = ~((layer5_outputs[1208]) & (layer5_outputs[1361]));
    assign layer6_outputs[1101] = ~(layer5_outputs[2381]);
    assign layer6_outputs[1102] = layer5_outputs[3469];
    assign layer6_outputs[1103] = ~(layer5_outputs[4469]);
    assign layer6_outputs[1104] = layer5_outputs[270];
    assign layer6_outputs[1105] = (layer5_outputs[2682]) | (layer5_outputs[1007]);
    assign layer6_outputs[1106] = layer5_outputs[234];
    assign layer6_outputs[1107] = layer5_outputs[4963];
    assign layer6_outputs[1108] = (layer5_outputs[4875]) & ~(layer5_outputs[2571]);
    assign layer6_outputs[1109] = layer5_outputs[3760];
    assign layer6_outputs[1110] = layer5_outputs[4992];
    assign layer6_outputs[1111] = (layer5_outputs[3950]) & ~(layer5_outputs[2859]);
    assign layer6_outputs[1112] = layer5_outputs[2644];
    assign layer6_outputs[1113] = (layer5_outputs[1894]) & ~(layer5_outputs[983]);
    assign layer6_outputs[1114] = ~((layer5_outputs[209]) & (layer5_outputs[4916]));
    assign layer6_outputs[1115] = ~(layer5_outputs[314]);
    assign layer6_outputs[1116] = layer5_outputs[5100];
    assign layer6_outputs[1117] = (layer5_outputs[1231]) | (layer5_outputs[4765]);
    assign layer6_outputs[1118] = 1'b1;
    assign layer6_outputs[1119] = layer5_outputs[921];
    assign layer6_outputs[1120] = ~(layer5_outputs[2021]);
    assign layer6_outputs[1121] = (layer5_outputs[3120]) & (layer5_outputs[4032]);
    assign layer6_outputs[1122] = ~((layer5_outputs[2823]) | (layer5_outputs[1090]));
    assign layer6_outputs[1123] = layer5_outputs[3700];
    assign layer6_outputs[1124] = layer5_outputs[4444];
    assign layer6_outputs[1125] = ~((layer5_outputs[584]) | (layer5_outputs[1367]));
    assign layer6_outputs[1126] = (layer5_outputs[2677]) ^ (layer5_outputs[1597]);
    assign layer6_outputs[1127] = (layer5_outputs[2569]) ^ (layer5_outputs[2251]);
    assign layer6_outputs[1128] = layer5_outputs[3028];
    assign layer6_outputs[1129] = layer5_outputs[1570];
    assign layer6_outputs[1130] = ~((layer5_outputs[188]) | (layer5_outputs[1479]));
    assign layer6_outputs[1131] = ~(layer5_outputs[1089]);
    assign layer6_outputs[1132] = ~((layer5_outputs[81]) | (layer5_outputs[4072]));
    assign layer6_outputs[1133] = layer5_outputs[2496];
    assign layer6_outputs[1134] = ~((layer5_outputs[2046]) ^ (layer5_outputs[536]));
    assign layer6_outputs[1135] = (layer5_outputs[7]) & ~(layer5_outputs[861]);
    assign layer6_outputs[1136] = ~(layer5_outputs[2142]) | (layer5_outputs[4505]);
    assign layer6_outputs[1137] = layer5_outputs[812];
    assign layer6_outputs[1138] = layer5_outputs[3633];
    assign layer6_outputs[1139] = ~(layer5_outputs[3124]);
    assign layer6_outputs[1140] = ~(layer5_outputs[2901]);
    assign layer6_outputs[1141] = ~(layer5_outputs[1242]);
    assign layer6_outputs[1142] = ~(layer5_outputs[3647]) | (layer5_outputs[3470]);
    assign layer6_outputs[1143] = ~(layer5_outputs[4379]) | (layer5_outputs[4434]);
    assign layer6_outputs[1144] = ~(layer5_outputs[5093]);
    assign layer6_outputs[1145] = ~((layer5_outputs[1945]) ^ (layer5_outputs[562]));
    assign layer6_outputs[1146] = layer5_outputs[3351];
    assign layer6_outputs[1147] = (layer5_outputs[892]) ^ (layer5_outputs[3101]);
    assign layer6_outputs[1148] = ~(layer5_outputs[1940]);
    assign layer6_outputs[1149] = ~(layer5_outputs[4895]);
    assign layer6_outputs[1150] = ~(layer5_outputs[1961]);
    assign layer6_outputs[1151] = ~(layer5_outputs[529]);
    assign layer6_outputs[1152] = ~((layer5_outputs[1926]) & (layer5_outputs[994]));
    assign layer6_outputs[1153] = layer5_outputs[964];
    assign layer6_outputs[1154] = ~((layer5_outputs[2056]) ^ (layer5_outputs[2006]));
    assign layer6_outputs[1155] = (layer5_outputs[1777]) & ~(layer5_outputs[3683]);
    assign layer6_outputs[1156] = ~(layer5_outputs[68]);
    assign layer6_outputs[1157] = ~(layer5_outputs[1787]);
    assign layer6_outputs[1158] = (layer5_outputs[4160]) | (layer5_outputs[3065]);
    assign layer6_outputs[1159] = layer5_outputs[122];
    assign layer6_outputs[1160] = ~(layer5_outputs[2481]) | (layer5_outputs[3774]);
    assign layer6_outputs[1161] = 1'b0;
    assign layer6_outputs[1162] = ~(layer5_outputs[1576]);
    assign layer6_outputs[1163] = ~((layer5_outputs[779]) ^ (layer5_outputs[963]));
    assign layer6_outputs[1164] = ~(layer5_outputs[4581]) | (layer5_outputs[2976]);
    assign layer6_outputs[1165] = (layer5_outputs[1015]) ^ (layer5_outputs[3269]);
    assign layer6_outputs[1166] = ~((layer5_outputs[3984]) | (layer5_outputs[3650]));
    assign layer6_outputs[1167] = ~((layer5_outputs[1829]) & (layer5_outputs[2029]));
    assign layer6_outputs[1168] = ~((layer5_outputs[2463]) & (layer5_outputs[2218]));
    assign layer6_outputs[1169] = ~(layer5_outputs[4843]);
    assign layer6_outputs[1170] = ~(layer5_outputs[3683]);
    assign layer6_outputs[1171] = ~((layer5_outputs[2099]) & (layer5_outputs[1912]));
    assign layer6_outputs[1172] = (layer5_outputs[598]) | (layer5_outputs[1061]);
    assign layer6_outputs[1173] = layer5_outputs[3626];
    assign layer6_outputs[1174] = ~(layer5_outputs[3628]) | (layer5_outputs[767]);
    assign layer6_outputs[1175] = layer5_outputs[2231];
    assign layer6_outputs[1176] = ~(layer5_outputs[2130]);
    assign layer6_outputs[1177] = ~(layer5_outputs[3994]);
    assign layer6_outputs[1178] = (layer5_outputs[614]) | (layer5_outputs[1892]);
    assign layer6_outputs[1179] = layer5_outputs[4341];
    assign layer6_outputs[1180] = ~(layer5_outputs[435]);
    assign layer6_outputs[1181] = (layer5_outputs[4292]) & ~(layer5_outputs[3464]);
    assign layer6_outputs[1182] = ~(layer5_outputs[2901]);
    assign layer6_outputs[1183] = ~(layer5_outputs[3569]);
    assign layer6_outputs[1184] = ~(layer5_outputs[3850]);
    assign layer6_outputs[1185] = ~(layer5_outputs[3006]);
    assign layer6_outputs[1186] = layer5_outputs[1717];
    assign layer6_outputs[1187] = ~(layer5_outputs[29]);
    assign layer6_outputs[1188] = layer5_outputs[2768];
    assign layer6_outputs[1189] = ~((layer5_outputs[2026]) ^ (layer5_outputs[1546]));
    assign layer6_outputs[1190] = ~((layer5_outputs[3037]) & (layer5_outputs[1806]));
    assign layer6_outputs[1191] = (layer5_outputs[3888]) & ~(layer5_outputs[948]);
    assign layer6_outputs[1192] = (layer5_outputs[4532]) & ~(layer5_outputs[1474]);
    assign layer6_outputs[1193] = (layer5_outputs[3856]) & ~(layer5_outputs[3784]);
    assign layer6_outputs[1194] = ~((layer5_outputs[4334]) ^ (layer5_outputs[1571]));
    assign layer6_outputs[1195] = ~(layer5_outputs[438]);
    assign layer6_outputs[1196] = layer5_outputs[4];
    assign layer6_outputs[1197] = ~(layer5_outputs[4051]);
    assign layer6_outputs[1198] = layer5_outputs[418];
    assign layer6_outputs[1199] = ~(layer5_outputs[3067]);
    assign layer6_outputs[1200] = (layer5_outputs[2873]) & (layer5_outputs[1404]);
    assign layer6_outputs[1201] = ~((layer5_outputs[3220]) | (layer5_outputs[2085]));
    assign layer6_outputs[1202] = layer5_outputs[4727];
    assign layer6_outputs[1203] = (layer5_outputs[1915]) | (layer5_outputs[3194]);
    assign layer6_outputs[1204] = layer5_outputs[3830];
    assign layer6_outputs[1205] = layer5_outputs[1783];
    assign layer6_outputs[1206] = ~(layer5_outputs[1150]);
    assign layer6_outputs[1207] = ~((layer5_outputs[2267]) | (layer5_outputs[2153]));
    assign layer6_outputs[1208] = (layer5_outputs[2131]) & ~(layer5_outputs[4063]);
    assign layer6_outputs[1209] = ~(layer5_outputs[3851]) | (layer5_outputs[117]);
    assign layer6_outputs[1210] = ~(layer5_outputs[3872]);
    assign layer6_outputs[1211] = (layer5_outputs[2391]) & ~(layer5_outputs[1643]);
    assign layer6_outputs[1212] = ~((layer5_outputs[4394]) | (layer5_outputs[3338]));
    assign layer6_outputs[1213] = layer5_outputs[4282];
    assign layer6_outputs[1214] = ~((layer5_outputs[1810]) & (layer5_outputs[4331]));
    assign layer6_outputs[1215] = (layer5_outputs[763]) | (layer5_outputs[1818]);
    assign layer6_outputs[1216] = ~((layer5_outputs[41]) ^ (layer5_outputs[645]));
    assign layer6_outputs[1217] = ~(layer5_outputs[3479]) | (layer5_outputs[3372]);
    assign layer6_outputs[1218] = (layer5_outputs[4257]) & ~(layer5_outputs[1076]);
    assign layer6_outputs[1219] = ~(layer5_outputs[1217]);
    assign layer6_outputs[1220] = ~(layer5_outputs[2077]);
    assign layer6_outputs[1221] = layer5_outputs[5087];
    assign layer6_outputs[1222] = ~(layer5_outputs[4066]);
    assign layer6_outputs[1223] = ~(layer5_outputs[588]);
    assign layer6_outputs[1224] = (layer5_outputs[4580]) ^ (layer5_outputs[3575]);
    assign layer6_outputs[1225] = (layer5_outputs[1123]) ^ (layer5_outputs[151]);
    assign layer6_outputs[1226] = ~(layer5_outputs[5111]);
    assign layer6_outputs[1227] = ~(layer5_outputs[914]) | (layer5_outputs[4800]);
    assign layer6_outputs[1228] = ~(layer5_outputs[3142]) | (layer5_outputs[4752]);
    assign layer6_outputs[1229] = layer5_outputs[846];
    assign layer6_outputs[1230] = ~(layer5_outputs[1362]);
    assign layer6_outputs[1231] = ~(layer5_outputs[263]);
    assign layer6_outputs[1232] = layer5_outputs[950];
    assign layer6_outputs[1233] = ~(layer5_outputs[1995]) | (layer5_outputs[799]);
    assign layer6_outputs[1234] = ~(layer5_outputs[3564]);
    assign layer6_outputs[1235] = layer5_outputs[2238];
    assign layer6_outputs[1236] = (layer5_outputs[4237]) & (layer5_outputs[1634]);
    assign layer6_outputs[1237] = (layer5_outputs[4316]) & (layer5_outputs[3937]);
    assign layer6_outputs[1238] = (layer5_outputs[1467]) & ~(layer5_outputs[5084]);
    assign layer6_outputs[1239] = layer5_outputs[177];
    assign layer6_outputs[1240] = ~(layer5_outputs[3564]) | (layer5_outputs[3268]);
    assign layer6_outputs[1241] = ~((layer5_outputs[2675]) ^ (layer5_outputs[3041]));
    assign layer6_outputs[1242] = ~(layer5_outputs[2556]);
    assign layer6_outputs[1243] = layer5_outputs[1417];
    assign layer6_outputs[1244] = layer5_outputs[3981];
    assign layer6_outputs[1245] = layer5_outputs[3777];
    assign layer6_outputs[1246] = ~((layer5_outputs[883]) & (layer5_outputs[1171]));
    assign layer6_outputs[1247] = ~(layer5_outputs[76]);
    assign layer6_outputs[1248] = layer5_outputs[1515];
    assign layer6_outputs[1249] = 1'b0;
    assign layer6_outputs[1250] = ~((layer5_outputs[2973]) ^ (layer5_outputs[3963]));
    assign layer6_outputs[1251] = ~((layer5_outputs[168]) & (layer5_outputs[2960]));
    assign layer6_outputs[1252] = ~(layer5_outputs[2025]);
    assign layer6_outputs[1253] = ~((layer5_outputs[5079]) & (layer5_outputs[2411]));
    assign layer6_outputs[1254] = ~(layer5_outputs[3827]);
    assign layer6_outputs[1255] = (layer5_outputs[141]) ^ (layer5_outputs[1158]);
    assign layer6_outputs[1256] = ~(layer5_outputs[2468]) | (layer5_outputs[1572]);
    assign layer6_outputs[1257] = layer5_outputs[439];
    assign layer6_outputs[1258] = layer5_outputs[5005];
    assign layer6_outputs[1259] = layer5_outputs[1701];
    assign layer6_outputs[1260] = ~(layer5_outputs[3990]);
    assign layer6_outputs[1261] = ~(layer5_outputs[987]) | (layer5_outputs[3394]);
    assign layer6_outputs[1262] = (layer5_outputs[624]) & ~(layer5_outputs[217]);
    assign layer6_outputs[1263] = layer5_outputs[2446];
    assign layer6_outputs[1264] = layer5_outputs[2382];
    assign layer6_outputs[1265] = ~(layer5_outputs[2307]);
    assign layer6_outputs[1266] = (layer5_outputs[2475]) ^ (layer5_outputs[2178]);
    assign layer6_outputs[1267] = 1'b1;
    assign layer6_outputs[1268] = layer5_outputs[64];
    assign layer6_outputs[1269] = ~(layer5_outputs[4613]);
    assign layer6_outputs[1270] = layer5_outputs[4833];
    assign layer6_outputs[1271] = ~(layer5_outputs[1910]);
    assign layer6_outputs[1272] = ~(layer5_outputs[3502]);
    assign layer6_outputs[1273] = layer5_outputs[4720];
    assign layer6_outputs[1274] = ~(layer5_outputs[251]);
    assign layer6_outputs[1275] = layer5_outputs[5068];
    assign layer6_outputs[1276] = layer5_outputs[384];
    assign layer6_outputs[1277] = ~((layer5_outputs[4488]) ^ (layer5_outputs[2707]));
    assign layer6_outputs[1278] = ~(layer5_outputs[224]);
    assign layer6_outputs[1279] = ~(layer5_outputs[4233]);
    assign layer6_outputs[1280] = ~(layer5_outputs[4685]);
    assign layer6_outputs[1281] = (layer5_outputs[4684]) ^ (layer5_outputs[157]);
    assign layer6_outputs[1282] = ~(layer5_outputs[2997]) | (layer5_outputs[4709]);
    assign layer6_outputs[1283] = layer5_outputs[835];
    assign layer6_outputs[1284] = layer5_outputs[2562];
    assign layer6_outputs[1285] = ~(layer5_outputs[3625]);
    assign layer6_outputs[1286] = (layer5_outputs[395]) & (layer5_outputs[2626]);
    assign layer6_outputs[1287] = layer5_outputs[3202];
    assign layer6_outputs[1288] = layer5_outputs[102];
    assign layer6_outputs[1289] = ~(layer5_outputs[4058]);
    assign layer6_outputs[1290] = ~((layer5_outputs[4038]) ^ (layer5_outputs[2925]));
    assign layer6_outputs[1291] = layer5_outputs[2469];
    assign layer6_outputs[1292] = layer5_outputs[1281];
    assign layer6_outputs[1293] = layer5_outputs[2881];
    assign layer6_outputs[1294] = ~(layer5_outputs[3594]);
    assign layer6_outputs[1295] = ~((layer5_outputs[4163]) | (layer5_outputs[2600]));
    assign layer6_outputs[1296] = (layer5_outputs[4486]) & (layer5_outputs[1760]);
    assign layer6_outputs[1297] = layer5_outputs[4941];
    assign layer6_outputs[1298] = layer5_outputs[3813];
    assign layer6_outputs[1299] = ~(layer5_outputs[2353]) | (layer5_outputs[3585]);
    assign layer6_outputs[1300] = ~(layer5_outputs[510]);
    assign layer6_outputs[1301] = ~((layer5_outputs[826]) | (layer5_outputs[225]));
    assign layer6_outputs[1302] = (layer5_outputs[192]) ^ (layer5_outputs[1030]);
    assign layer6_outputs[1303] = ~(layer5_outputs[3406]);
    assign layer6_outputs[1304] = layer5_outputs[352];
    assign layer6_outputs[1305] = ~((layer5_outputs[618]) ^ (layer5_outputs[2284]));
    assign layer6_outputs[1306] = ~((layer5_outputs[2975]) ^ (layer5_outputs[1670]));
    assign layer6_outputs[1307] = (layer5_outputs[2661]) ^ (layer5_outputs[1054]);
    assign layer6_outputs[1308] = layer5_outputs[1295];
    assign layer6_outputs[1309] = (layer5_outputs[2892]) & (layer5_outputs[1092]);
    assign layer6_outputs[1310] = (layer5_outputs[2547]) & ~(layer5_outputs[2429]);
    assign layer6_outputs[1311] = ~(layer5_outputs[1055]);
    assign layer6_outputs[1312] = ~(layer5_outputs[3809]) | (layer5_outputs[1001]);
    assign layer6_outputs[1313] = layer5_outputs[2669];
    assign layer6_outputs[1314] = layer5_outputs[4676];
    assign layer6_outputs[1315] = ~(layer5_outputs[387]);
    assign layer6_outputs[1316] = ~((layer5_outputs[2383]) ^ (layer5_outputs[3486]));
    assign layer6_outputs[1317] = ~(layer5_outputs[2148]);
    assign layer6_outputs[1318] = ~(layer5_outputs[3469]);
    assign layer6_outputs[1319] = ~((layer5_outputs[2814]) ^ (layer5_outputs[4161]));
    assign layer6_outputs[1320] = layer5_outputs[3189];
    assign layer6_outputs[1321] = ~(layer5_outputs[1937]);
    assign layer6_outputs[1322] = ~(layer5_outputs[2]);
    assign layer6_outputs[1323] = ~((layer5_outputs[4950]) & (layer5_outputs[1017]));
    assign layer6_outputs[1324] = ~((layer5_outputs[3415]) ^ (layer5_outputs[2148]));
    assign layer6_outputs[1325] = layer5_outputs[2395];
    assign layer6_outputs[1326] = (layer5_outputs[3751]) ^ (layer5_outputs[1122]);
    assign layer6_outputs[1327] = ~(layer5_outputs[101]) | (layer5_outputs[5026]);
    assign layer6_outputs[1328] = (layer5_outputs[2359]) & (layer5_outputs[2888]);
    assign layer6_outputs[1329] = layer5_outputs[4866];
    assign layer6_outputs[1330] = ~(layer5_outputs[4030]);
    assign layer6_outputs[1331] = layer5_outputs[4063];
    assign layer6_outputs[1332] = ~(layer5_outputs[1311]);
    assign layer6_outputs[1333] = ~((layer5_outputs[2243]) ^ (layer5_outputs[3533]));
    assign layer6_outputs[1334] = ~(layer5_outputs[1380]);
    assign layer6_outputs[1335] = (layer5_outputs[3215]) & ~(layer5_outputs[1997]);
    assign layer6_outputs[1336] = (layer5_outputs[1782]) & ~(layer5_outputs[1611]);
    assign layer6_outputs[1337] = layer5_outputs[988];
    assign layer6_outputs[1338] = (layer5_outputs[1448]) ^ (layer5_outputs[4060]);
    assign layer6_outputs[1339] = ~(layer5_outputs[1769]);
    assign layer6_outputs[1340] = ~((layer5_outputs[1920]) | (layer5_outputs[1854]));
    assign layer6_outputs[1341] = ~(layer5_outputs[5003]);
    assign layer6_outputs[1342] = layer5_outputs[2098];
    assign layer6_outputs[1343] = ~(layer5_outputs[1692]) | (layer5_outputs[757]);
    assign layer6_outputs[1344] = (layer5_outputs[2622]) & (layer5_outputs[215]);
    assign layer6_outputs[1345] = (layer5_outputs[4336]) ^ (layer5_outputs[3312]);
    assign layer6_outputs[1346] = (layer5_outputs[2994]) & ~(layer5_outputs[3149]);
    assign layer6_outputs[1347] = ~(layer5_outputs[2355]);
    assign layer6_outputs[1348] = ~((layer5_outputs[3641]) & (layer5_outputs[2072]));
    assign layer6_outputs[1349] = layer5_outputs[4791];
    assign layer6_outputs[1350] = layer5_outputs[1454];
    assign layer6_outputs[1351] = ~((layer5_outputs[2577]) | (layer5_outputs[4320]));
    assign layer6_outputs[1352] = layer5_outputs[3252];
    assign layer6_outputs[1353] = layer5_outputs[1992];
    assign layer6_outputs[1354] = ~((layer5_outputs[5065]) ^ (layer5_outputs[3544]));
    assign layer6_outputs[1355] = layer5_outputs[795];
    assign layer6_outputs[1356] = layer5_outputs[1453];
    assign layer6_outputs[1357] = layer5_outputs[2955];
    assign layer6_outputs[1358] = ~(layer5_outputs[1162]);
    assign layer6_outputs[1359] = layer5_outputs[2836];
    assign layer6_outputs[1360] = ~((layer5_outputs[3754]) & (layer5_outputs[1470]));
    assign layer6_outputs[1361] = (layer5_outputs[4314]) ^ (layer5_outputs[390]);
    assign layer6_outputs[1362] = ~(layer5_outputs[3799]) | (layer5_outputs[2856]);
    assign layer6_outputs[1363] = (layer5_outputs[5110]) ^ (layer5_outputs[3156]);
    assign layer6_outputs[1364] = ~(layer5_outputs[3281]);
    assign layer6_outputs[1365] = (layer5_outputs[1409]) & ~(layer5_outputs[331]);
    assign layer6_outputs[1366] = ~(layer5_outputs[265]);
    assign layer6_outputs[1367] = (layer5_outputs[3893]) & (layer5_outputs[4688]);
    assign layer6_outputs[1368] = ~(layer5_outputs[903]);
    assign layer6_outputs[1369] = ~(layer5_outputs[3405]);
    assign layer6_outputs[1370] = layer5_outputs[4022];
    assign layer6_outputs[1371] = layer5_outputs[4507];
    assign layer6_outputs[1372] = ~(layer5_outputs[4211]);
    assign layer6_outputs[1373] = (layer5_outputs[175]) ^ (layer5_outputs[1685]);
    assign layer6_outputs[1374] = layer5_outputs[703];
    assign layer6_outputs[1375] = ~(layer5_outputs[3541]);
    assign layer6_outputs[1376] = (layer5_outputs[1619]) & ~(layer5_outputs[4720]);
    assign layer6_outputs[1377] = (layer5_outputs[1722]) | (layer5_outputs[1236]);
    assign layer6_outputs[1378] = ~((layer5_outputs[36]) ^ (layer5_outputs[808]));
    assign layer6_outputs[1379] = ~(layer5_outputs[656]);
    assign layer6_outputs[1380] = (layer5_outputs[4107]) & (layer5_outputs[3952]);
    assign layer6_outputs[1381] = layer5_outputs[118];
    assign layer6_outputs[1382] = layer5_outputs[33];
    assign layer6_outputs[1383] = (layer5_outputs[3077]) ^ (layer5_outputs[1492]);
    assign layer6_outputs[1384] = ~(layer5_outputs[3416]);
    assign layer6_outputs[1385] = layer5_outputs[4116];
    assign layer6_outputs[1386] = ~(layer5_outputs[412]);
    assign layer6_outputs[1387] = layer5_outputs[4220];
    assign layer6_outputs[1388] = ~(layer5_outputs[4939]);
    assign layer6_outputs[1389] = layer5_outputs[3040];
    assign layer6_outputs[1390] = (layer5_outputs[4418]) ^ (layer5_outputs[2614]);
    assign layer6_outputs[1391] = ~(layer5_outputs[1921]);
    assign layer6_outputs[1392] = layer5_outputs[3875];
    assign layer6_outputs[1393] = ~(layer5_outputs[3210]);
    assign layer6_outputs[1394] = (layer5_outputs[1214]) ^ (layer5_outputs[3720]);
    assign layer6_outputs[1395] = ~(layer5_outputs[3750]);
    assign layer6_outputs[1396] = ~(layer5_outputs[2986]);
    assign layer6_outputs[1397] = (layer5_outputs[2040]) & ~(layer5_outputs[978]);
    assign layer6_outputs[1398] = layer5_outputs[166];
    assign layer6_outputs[1399] = ~(layer5_outputs[2106]);
    assign layer6_outputs[1400] = (layer5_outputs[273]) ^ (layer5_outputs[1110]);
    assign layer6_outputs[1401] = (layer5_outputs[3266]) ^ (layer5_outputs[486]);
    assign layer6_outputs[1402] = ~(layer5_outputs[1482]);
    assign layer6_outputs[1403] = ~((layer5_outputs[1261]) ^ (layer5_outputs[1537]));
    assign layer6_outputs[1404] = layer5_outputs[5024];
    assign layer6_outputs[1405] = 1'b0;
    assign layer6_outputs[1406] = ~(layer5_outputs[2246]);
    assign layer6_outputs[1407] = layer5_outputs[2991];
    assign layer6_outputs[1408] = ~((layer5_outputs[3631]) ^ (layer5_outputs[3105]));
    assign layer6_outputs[1409] = ~((layer5_outputs[2134]) | (layer5_outputs[1159]));
    assign layer6_outputs[1410] = ~(layer5_outputs[1785]) | (layer5_outputs[3535]);
    assign layer6_outputs[1411] = ~(layer5_outputs[3759]);
    assign layer6_outputs[1412] = ~(layer5_outputs[2942]);
    assign layer6_outputs[1413] = (layer5_outputs[4430]) ^ (layer5_outputs[3490]);
    assign layer6_outputs[1414] = ~(layer5_outputs[2783]);
    assign layer6_outputs[1415] = ~(layer5_outputs[874]);
    assign layer6_outputs[1416] = layer5_outputs[3818];
    assign layer6_outputs[1417] = ~(layer5_outputs[4686]) | (layer5_outputs[3687]);
    assign layer6_outputs[1418] = (layer5_outputs[2373]) | (layer5_outputs[1455]);
    assign layer6_outputs[1419] = ~(layer5_outputs[3235]);
    assign layer6_outputs[1420] = (layer5_outputs[3961]) & (layer5_outputs[4665]);
    assign layer6_outputs[1421] = (layer5_outputs[4973]) ^ (layer5_outputs[53]);
    assign layer6_outputs[1422] = layer5_outputs[4330];
    assign layer6_outputs[1423] = layer5_outputs[3187];
    assign layer6_outputs[1424] = ~((layer5_outputs[2290]) ^ (layer5_outputs[343]));
    assign layer6_outputs[1425] = ~(layer5_outputs[2902]) | (layer5_outputs[581]);
    assign layer6_outputs[1426] = (layer5_outputs[320]) | (layer5_outputs[1102]);
    assign layer6_outputs[1427] = (layer5_outputs[1712]) ^ (layer5_outputs[516]);
    assign layer6_outputs[1428] = layer5_outputs[1045];
    assign layer6_outputs[1429] = (layer5_outputs[2342]) & ~(layer5_outputs[1408]);
    assign layer6_outputs[1430] = 1'b1;
    assign layer6_outputs[1431] = ~(layer5_outputs[3912]);
    assign layer6_outputs[1432] = layer5_outputs[3392];
    assign layer6_outputs[1433] = ~(layer5_outputs[3448]);
    assign layer6_outputs[1434] = ~(layer5_outputs[3657]) | (layer5_outputs[2140]);
    assign layer6_outputs[1435] = layer5_outputs[3844];
    assign layer6_outputs[1436] = ~(layer5_outputs[1573]) | (layer5_outputs[1948]);
    assign layer6_outputs[1437] = layer5_outputs[3690];
    assign layer6_outputs[1438] = ~(layer5_outputs[3356]) | (layer5_outputs[4472]);
    assign layer6_outputs[1439] = ~(layer5_outputs[3704]);
    assign layer6_outputs[1440] = ~(layer5_outputs[3947]);
    assign layer6_outputs[1441] = layer5_outputs[3162];
    assign layer6_outputs[1442] = (layer5_outputs[1550]) | (layer5_outputs[2880]);
    assign layer6_outputs[1443] = (layer5_outputs[2607]) ^ (layer5_outputs[3462]);
    assign layer6_outputs[1444] = (layer5_outputs[4505]) & (layer5_outputs[3596]);
    assign layer6_outputs[1445] = ~(layer5_outputs[3249]) | (layer5_outputs[2596]);
    assign layer6_outputs[1446] = (layer5_outputs[264]) & (layer5_outputs[2788]);
    assign layer6_outputs[1447] = ~(layer5_outputs[4512]);
    assign layer6_outputs[1448] = layer5_outputs[1038];
    assign layer6_outputs[1449] = (layer5_outputs[2844]) & (layer5_outputs[3761]);
    assign layer6_outputs[1450] = layer5_outputs[3671];
    assign layer6_outputs[1451] = 1'b1;
    assign layer6_outputs[1452] = (layer5_outputs[3152]) & ~(layer5_outputs[2803]);
    assign layer6_outputs[1453] = ~(layer5_outputs[5030]);
    assign layer6_outputs[1454] = layer5_outputs[1405];
    assign layer6_outputs[1455] = ~((layer5_outputs[5083]) & (layer5_outputs[1655]));
    assign layer6_outputs[1456] = ~(layer5_outputs[1080]);
    assign layer6_outputs[1457] = ~(layer5_outputs[1739]);
    assign layer6_outputs[1458] = 1'b0;
    assign layer6_outputs[1459] = layer5_outputs[334];
    assign layer6_outputs[1460] = (layer5_outputs[4283]) | (layer5_outputs[3978]);
    assign layer6_outputs[1461] = layer5_outputs[2334];
    assign layer6_outputs[1462] = ~((layer5_outputs[3814]) ^ (layer5_outputs[4302]));
    assign layer6_outputs[1463] = ~((layer5_outputs[414]) | (layer5_outputs[5086]));
    assign layer6_outputs[1464] = (layer5_outputs[1019]) & (layer5_outputs[5106]);
    assign layer6_outputs[1465] = (layer5_outputs[92]) | (layer5_outputs[5074]);
    assign layer6_outputs[1466] = (layer5_outputs[4751]) & ~(layer5_outputs[1439]);
    assign layer6_outputs[1467] = ~((layer5_outputs[4470]) ^ (layer5_outputs[3133]));
    assign layer6_outputs[1468] = 1'b0;
    assign layer6_outputs[1469] = ~(layer5_outputs[3976]);
    assign layer6_outputs[1470] = (layer5_outputs[507]) & ~(layer5_outputs[1731]);
    assign layer6_outputs[1471] = layer5_outputs[1677];
    assign layer6_outputs[1472] = ~(layer5_outputs[1302]);
    assign layer6_outputs[1473] = layer5_outputs[3051];
    assign layer6_outputs[1474] = ~(layer5_outputs[4095]);
    assign layer6_outputs[1475] = ~((layer5_outputs[4461]) ^ (layer5_outputs[2126]));
    assign layer6_outputs[1476] = ~((layer5_outputs[196]) & (layer5_outputs[3575]));
    assign layer6_outputs[1477] = ~((layer5_outputs[3503]) & (layer5_outputs[1043]));
    assign layer6_outputs[1478] = ~(layer5_outputs[5051]);
    assign layer6_outputs[1479] = layer5_outputs[1588];
    assign layer6_outputs[1480] = (layer5_outputs[1626]) & (layer5_outputs[4230]);
    assign layer6_outputs[1481] = ~(layer5_outputs[4288]) | (layer5_outputs[385]);
    assign layer6_outputs[1482] = ~((layer5_outputs[224]) & (layer5_outputs[3860]));
    assign layer6_outputs[1483] = ~((layer5_outputs[1807]) | (layer5_outputs[1097]));
    assign layer6_outputs[1484] = ~(layer5_outputs[3085]);
    assign layer6_outputs[1485] = ~((layer5_outputs[1599]) ^ (layer5_outputs[2529]));
    assign layer6_outputs[1486] = layer5_outputs[766];
    assign layer6_outputs[1487] = ~((layer5_outputs[962]) ^ (layer5_outputs[1921]));
    assign layer6_outputs[1488] = ~(layer5_outputs[3559]);
    assign layer6_outputs[1489] = layer5_outputs[1925];
    assign layer6_outputs[1490] = (layer5_outputs[3769]) ^ (layer5_outputs[1675]);
    assign layer6_outputs[1491] = layer5_outputs[4750];
    assign layer6_outputs[1492] = ~((layer5_outputs[3147]) | (layer5_outputs[4671]));
    assign layer6_outputs[1493] = layer5_outputs[1016];
    assign layer6_outputs[1494] = ~(layer5_outputs[2619]);
    assign layer6_outputs[1495] = ~((layer5_outputs[4354]) ^ (layer5_outputs[3518]));
    assign layer6_outputs[1496] = ~((layer5_outputs[4921]) ^ (layer5_outputs[4004]));
    assign layer6_outputs[1497] = ~(layer5_outputs[2261]);
    assign layer6_outputs[1498] = ~(layer5_outputs[5062]);
    assign layer6_outputs[1499] = layer5_outputs[2374];
    assign layer6_outputs[1500] = ~(layer5_outputs[2843]) | (layer5_outputs[1958]);
    assign layer6_outputs[1501] = ~(layer5_outputs[237]);
    assign layer6_outputs[1502] = layer5_outputs[2059];
    assign layer6_outputs[1503] = (layer5_outputs[4637]) ^ (layer5_outputs[1759]);
    assign layer6_outputs[1504] = layer5_outputs[1104];
    assign layer6_outputs[1505] = ~(layer5_outputs[4377]) | (layer5_outputs[1329]);
    assign layer6_outputs[1506] = ~((layer5_outputs[4408]) ^ (layer5_outputs[4937]));
    assign layer6_outputs[1507] = layer5_outputs[4213];
    assign layer6_outputs[1508] = ~((layer5_outputs[1430]) & (layer5_outputs[3668]));
    assign layer6_outputs[1509] = 1'b0;
    assign layer6_outputs[1510] = ~(layer5_outputs[111]) | (layer5_outputs[3216]);
    assign layer6_outputs[1511] = (layer5_outputs[2903]) | (layer5_outputs[4761]);
    assign layer6_outputs[1512] = (layer5_outputs[889]) ^ (layer5_outputs[3531]);
    assign layer6_outputs[1513] = (layer5_outputs[2233]) ^ (layer5_outputs[1936]);
    assign layer6_outputs[1514] = ~(layer5_outputs[152]);
    assign layer6_outputs[1515] = (layer5_outputs[1962]) & ~(layer5_outputs[1325]);
    assign layer6_outputs[1516] = ~(layer5_outputs[4032]);
    assign layer6_outputs[1517] = (layer5_outputs[4815]) & ~(layer5_outputs[3370]);
    assign layer6_outputs[1518] = ~(layer5_outputs[3355]) | (layer5_outputs[528]);
    assign layer6_outputs[1519] = (layer5_outputs[1698]) ^ (layer5_outputs[1403]);
    assign layer6_outputs[1520] = ~((layer5_outputs[504]) ^ (layer5_outputs[4421]));
    assign layer6_outputs[1521] = ~((layer5_outputs[3805]) | (layer5_outputs[4804]));
    assign layer6_outputs[1522] = (layer5_outputs[4850]) & (layer5_outputs[3]);
    assign layer6_outputs[1523] = layer5_outputs[3114];
    assign layer6_outputs[1524] = (layer5_outputs[2316]) | (layer5_outputs[1949]);
    assign layer6_outputs[1525] = layer5_outputs[2230];
    assign layer6_outputs[1526] = ~(layer5_outputs[4906]) | (layer5_outputs[1707]);
    assign layer6_outputs[1527] = ~(layer5_outputs[2945]);
    assign layer6_outputs[1528] = layer5_outputs[3836];
    assign layer6_outputs[1529] = ~(layer5_outputs[4524]);
    assign layer6_outputs[1530] = ~(layer5_outputs[3580]);
    assign layer6_outputs[1531] = ~(layer5_outputs[3097]);
    assign layer6_outputs[1532] = ~(layer5_outputs[3698]);
    assign layer6_outputs[1533] = (layer5_outputs[4263]) & (layer5_outputs[3560]);
    assign layer6_outputs[1534] = (layer5_outputs[1761]) & (layer5_outputs[4152]);
    assign layer6_outputs[1535] = ~((layer5_outputs[1973]) ^ (layer5_outputs[4321]));
    assign layer6_outputs[1536] = (layer5_outputs[1750]) ^ (layer5_outputs[369]);
    assign layer6_outputs[1537] = layer5_outputs[47];
    assign layer6_outputs[1538] = layer5_outputs[4920];
    assign layer6_outputs[1539] = layer5_outputs[2946];
    assign layer6_outputs[1540] = layer5_outputs[4547];
    assign layer6_outputs[1541] = layer5_outputs[2951];
    assign layer6_outputs[1542] = ~((layer5_outputs[3574]) ^ (layer5_outputs[70]));
    assign layer6_outputs[1543] = ~(layer5_outputs[2544]);
    assign layer6_outputs[1544] = layer5_outputs[2813];
    assign layer6_outputs[1545] = layer5_outputs[2169];
    assign layer6_outputs[1546] = ~(layer5_outputs[4251]);
    assign layer6_outputs[1547] = (layer5_outputs[4102]) ^ (layer5_outputs[3211]);
    assign layer6_outputs[1548] = ~(layer5_outputs[4744]);
    assign layer6_outputs[1549] = ~(layer5_outputs[2684]);
    assign layer6_outputs[1550] = ~(layer5_outputs[873]) | (layer5_outputs[1091]);
    assign layer6_outputs[1551] = layer5_outputs[2952];
    assign layer6_outputs[1552] = (layer5_outputs[4275]) | (layer5_outputs[4026]);
    assign layer6_outputs[1553] = layer5_outputs[3536];
    assign layer6_outputs[1554] = (layer5_outputs[239]) ^ (layer5_outputs[782]);
    assign layer6_outputs[1555] = ~((layer5_outputs[4570]) ^ (layer5_outputs[2457]));
    assign layer6_outputs[1556] = layer5_outputs[4092];
    assign layer6_outputs[1557] = layer5_outputs[4119];
    assign layer6_outputs[1558] = ~((layer5_outputs[2356]) & (layer5_outputs[543]));
    assign layer6_outputs[1559] = 1'b1;
    assign layer6_outputs[1560] = layer5_outputs[4405];
    assign layer6_outputs[1561] = 1'b1;
    assign layer6_outputs[1562] = (layer5_outputs[3546]) & ~(layer5_outputs[5096]);
    assign layer6_outputs[1563] = (layer5_outputs[3153]) & ~(layer5_outputs[1050]);
    assign layer6_outputs[1564] = layer5_outputs[4361];
    assign layer6_outputs[1565] = ~(layer5_outputs[427]);
    assign layer6_outputs[1566] = layer5_outputs[3640];
    assign layer6_outputs[1567] = ~((layer5_outputs[3670]) & (layer5_outputs[75]));
    assign layer6_outputs[1568] = 1'b0;
    assign layer6_outputs[1569] = layer5_outputs[4905];
    assign layer6_outputs[1570] = ~(layer5_outputs[279]);
    assign layer6_outputs[1571] = ~(layer5_outputs[2833]);
    assign layer6_outputs[1572] = ~(layer5_outputs[869]);
    assign layer6_outputs[1573] = (layer5_outputs[3091]) & (layer5_outputs[319]);
    assign layer6_outputs[1574] = ~(layer5_outputs[1728]);
    assign layer6_outputs[1575] = ~(layer5_outputs[225]);
    assign layer6_outputs[1576] = ~((layer5_outputs[3283]) & (layer5_outputs[2145]));
    assign layer6_outputs[1577] = ~(layer5_outputs[494]);
    assign layer6_outputs[1578] = layer5_outputs[1554];
    assign layer6_outputs[1579] = layer5_outputs[3159];
    assign layer6_outputs[1580] = (layer5_outputs[2998]) ^ (layer5_outputs[5038]);
    assign layer6_outputs[1581] = layer5_outputs[970];
    assign layer6_outputs[1582] = layer5_outputs[871];
    assign layer6_outputs[1583] = (layer5_outputs[4172]) & ~(layer5_outputs[1426]);
    assign layer6_outputs[1584] = layer5_outputs[3334];
    assign layer6_outputs[1585] = (layer5_outputs[2320]) & (layer5_outputs[4788]);
    assign layer6_outputs[1586] = ~((layer5_outputs[1227]) | (layer5_outputs[1047]));
    assign layer6_outputs[1587] = layer5_outputs[4179];
    assign layer6_outputs[1588] = layer5_outputs[4078];
    assign layer6_outputs[1589] = layer5_outputs[2458];
    assign layer6_outputs[1590] = 1'b0;
    assign layer6_outputs[1591] = ~(layer5_outputs[1271]);
    assign layer6_outputs[1592] = (layer5_outputs[4097]) & ~(layer5_outputs[3626]);
    assign layer6_outputs[1593] = ~(layer5_outputs[1396]);
    assign layer6_outputs[1594] = layer5_outputs[1767];
    assign layer6_outputs[1595] = ~(layer5_outputs[4616]);
    assign layer6_outputs[1596] = layer5_outputs[3199];
    assign layer6_outputs[1597] = ~((layer5_outputs[4253]) ^ (layer5_outputs[885]));
    assign layer6_outputs[1598] = ~(layer5_outputs[2813]);
    assign layer6_outputs[1599] = (layer5_outputs[5027]) ^ (layer5_outputs[2010]);
    assign layer6_outputs[1600] = ~(layer5_outputs[2116]);
    assign layer6_outputs[1601] = layer5_outputs[1473];
    assign layer6_outputs[1602] = ~((layer5_outputs[4255]) ^ (layer5_outputs[3706]));
    assign layer6_outputs[1603] = layer5_outputs[1824];
    assign layer6_outputs[1604] = ~(layer5_outputs[3889]) | (layer5_outputs[1155]);
    assign layer6_outputs[1605] = ~((layer5_outputs[882]) ^ (layer5_outputs[282]));
    assign layer6_outputs[1606] = layer5_outputs[3965];
    assign layer6_outputs[1607] = layer5_outputs[2282];
    assign layer6_outputs[1608] = ~(layer5_outputs[1976]);
    assign layer6_outputs[1609] = (layer5_outputs[1789]) | (layer5_outputs[874]);
    assign layer6_outputs[1610] = ~((layer5_outputs[4668]) ^ (layer5_outputs[4577]));
    assign layer6_outputs[1611] = ~(layer5_outputs[4502]);
    assign layer6_outputs[1612] = 1'b1;
    assign layer6_outputs[1613] = ~(layer5_outputs[1799]);
    assign layer6_outputs[1614] = layer5_outputs[1220];
    assign layer6_outputs[1615] = ~(layer5_outputs[1133]);
    assign layer6_outputs[1616] = (layer5_outputs[1267]) ^ (layer5_outputs[226]);
    assign layer6_outputs[1617] = ~(layer5_outputs[4122]);
    assign layer6_outputs[1618] = ~((layer5_outputs[1906]) ^ (layer5_outputs[101]));
    assign layer6_outputs[1619] = ~(layer5_outputs[3803]) | (layer5_outputs[2676]);
    assign layer6_outputs[1620] = ~(layer5_outputs[1446]) | (layer5_outputs[1770]);
    assign layer6_outputs[1621] = layer5_outputs[78];
    assign layer6_outputs[1622] = (layer5_outputs[119]) & ~(layer5_outputs[4947]);
    assign layer6_outputs[1623] = (layer5_outputs[2187]) & ~(layer5_outputs[2875]);
    assign layer6_outputs[1624] = layer5_outputs[1160];
    assign layer6_outputs[1625] = ~(layer5_outputs[1846]);
    assign layer6_outputs[1626] = layer5_outputs[3472];
    assign layer6_outputs[1627] = ~(layer5_outputs[4237]);
    assign layer6_outputs[1628] = (layer5_outputs[4656]) & ~(layer5_outputs[4979]);
    assign layer6_outputs[1629] = layer5_outputs[1365];
    assign layer6_outputs[1630] = layer5_outputs[3472];
    assign layer6_outputs[1631] = layer5_outputs[1663];
    assign layer6_outputs[1632] = ~(layer5_outputs[1337]) | (layer5_outputs[2442]);
    assign layer6_outputs[1633] = ~(layer5_outputs[4051]);
    assign layer6_outputs[1634] = ~(layer5_outputs[2404]);
    assign layer6_outputs[1635] = ~(layer5_outputs[2721]);
    assign layer6_outputs[1636] = ~(layer5_outputs[0]);
    assign layer6_outputs[1637] = (layer5_outputs[2218]) & ~(layer5_outputs[4198]);
    assign layer6_outputs[1638] = ~(layer5_outputs[464]);
    assign layer6_outputs[1639] = ~((layer5_outputs[626]) ^ (layer5_outputs[704]));
    assign layer6_outputs[1640] = ~((layer5_outputs[3221]) ^ (layer5_outputs[4821]));
    assign layer6_outputs[1641] = ~((layer5_outputs[4576]) ^ (layer5_outputs[3103]));
    assign layer6_outputs[1642] = ~(layer5_outputs[1805]) | (layer5_outputs[2894]);
    assign layer6_outputs[1643] = ~(layer5_outputs[4955]);
    assign layer6_outputs[1644] = ~((layer5_outputs[2057]) | (layer5_outputs[708]));
    assign layer6_outputs[1645] = ~(layer5_outputs[4214]);
    assign layer6_outputs[1646] = ~((layer5_outputs[4356]) ^ (layer5_outputs[5024]));
    assign layer6_outputs[1647] = (layer5_outputs[3359]) | (layer5_outputs[857]);
    assign layer6_outputs[1648] = layer5_outputs[72];
    assign layer6_outputs[1649] = (layer5_outputs[2368]) & ~(layer5_outputs[2930]);
    assign layer6_outputs[1650] = ~(layer5_outputs[2246]) | (layer5_outputs[4457]);
    assign layer6_outputs[1651] = ~((layer5_outputs[1827]) ^ (layer5_outputs[60]));
    assign layer6_outputs[1652] = ~((layer5_outputs[1901]) & (layer5_outputs[1010]));
    assign layer6_outputs[1653] = layer5_outputs[735];
    assign layer6_outputs[1654] = ~(layer5_outputs[3707]);
    assign layer6_outputs[1655] = (layer5_outputs[832]) | (layer5_outputs[3558]);
    assign layer6_outputs[1656] = layer5_outputs[2928];
    assign layer6_outputs[1657] = ~(layer5_outputs[917]) | (layer5_outputs[964]);
    assign layer6_outputs[1658] = ~((layer5_outputs[3882]) | (layer5_outputs[3838]));
    assign layer6_outputs[1659] = (layer5_outputs[3064]) & ~(layer5_outputs[3908]);
    assign layer6_outputs[1660] = (layer5_outputs[1630]) & (layer5_outputs[2532]);
    assign layer6_outputs[1661] = layer5_outputs[4707];
    assign layer6_outputs[1662] = (layer5_outputs[2837]) ^ (layer5_outputs[3340]);
    assign layer6_outputs[1663] = (layer5_outputs[4740]) & (layer5_outputs[2971]);
    assign layer6_outputs[1664] = (layer5_outputs[4768]) & ~(layer5_outputs[1090]);
    assign layer6_outputs[1665] = ~(layer5_outputs[2625]);
    assign layer6_outputs[1666] = ~(layer5_outputs[63]);
    assign layer6_outputs[1667] = ~(layer5_outputs[547]);
    assign layer6_outputs[1668] = ~(layer5_outputs[3251]);
    assign layer6_outputs[1669] = (layer5_outputs[887]) & ~(layer5_outputs[471]);
    assign layer6_outputs[1670] = layer5_outputs[4637];
    assign layer6_outputs[1671] = 1'b1;
    assign layer6_outputs[1672] = (layer5_outputs[2421]) & (layer5_outputs[901]);
    assign layer6_outputs[1673] = ~(layer5_outputs[3825]);
    assign layer6_outputs[1674] = (layer5_outputs[1196]) ^ (layer5_outputs[3845]);
    assign layer6_outputs[1675] = ~(layer5_outputs[22]);
    assign layer6_outputs[1676] = layer5_outputs[2683];
    assign layer6_outputs[1677] = ~((layer5_outputs[2147]) ^ (layer5_outputs[2847]));
    assign layer6_outputs[1678] = ~(layer5_outputs[1510]);
    assign layer6_outputs[1679] = ~((layer5_outputs[978]) & (layer5_outputs[3119]));
    assign layer6_outputs[1680] = (layer5_outputs[3680]) ^ (layer5_outputs[3113]);
    assign layer6_outputs[1681] = ~(layer5_outputs[3109]);
    assign layer6_outputs[1682] = layer5_outputs[2898];
    assign layer6_outputs[1683] = layer5_outputs[4878];
    assign layer6_outputs[1684] = ~(layer5_outputs[2042]);
    assign layer6_outputs[1685] = ~(layer5_outputs[1287]);
    assign layer6_outputs[1686] = (layer5_outputs[2758]) & (layer5_outputs[2740]);
    assign layer6_outputs[1687] = ~(layer5_outputs[3582]);
    assign layer6_outputs[1688] = ~((layer5_outputs[1136]) ^ (layer5_outputs[3840]));
    assign layer6_outputs[1689] = (layer5_outputs[5056]) | (layer5_outputs[2754]);
    assign layer6_outputs[1690] = (layer5_outputs[1422]) | (layer5_outputs[3193]);
    assign layer6_outputs[1691] = ~(layer5_outputs[3465]);
    assign layer6_outputs[1692] = ~(layer5_outputs[1354]);
    assign layer6_outputs[1693] = layer5_outputs[2376];
    assign layer6_outputs[1694] = ~((layer5_outputs[4500]) ^ (layer5_outputs[4706]));
    assign layer6_outputs[1695] = ~(layer5_outputs[140]);
    assign layer6_outputs[1696] = ~(layer5_outputs[3368]) | (layer5_outputs[1436]);
    assign layer6_outputs[1697] = ~(layer5_outputs[2835]);
    assign layer6_outputs[1698] = ~((layer5_outputs[2558]) ^ (layer5_outputs[1936]));
    assign layer6_outputs[1699] = ~(layer5_outputs[2675]) | (layer5_outputs[4933]);
    assign layer6_outputs[1700] = layer5_outputs[4841];
    assign layer6_outputs[1701] = layer5_outputs[4258];
    assign layer6_outputs[1702] = layer5_outputs[4744];
    assign layer6_outputs[1703] = layer5_outputs[1885];
    assign layer6_outputs[1704] = layer5_outputs[3391];
    assign layer6_outputs[1705] = layer5_outputs[4174];
    assign layer6_outputs[1706] = (layer5_outputs[1853]) ^ (layer5_outputs[317]);
    assign layer6_outputs[1707] = (layer5_outputs[442]) & ~(layer5_outputs[4317]);
    assign layer6_outputs[1708] = ~((layer5_outputs[4525]) & (layer5_outputs[2877]));
    assign layer6_outputs[1709] = layer5_outputs[180];
    assign layer6_outputs[1710] = (layer5_outputs[3455]) ^ (layer5_outputs[455]);
    assign layer6_outputs[1711] = layer5_outputs[2535];
    assign layer6_outputs[1712] = ~(layer5_outputs[4195]);
    assign layer6_outputs[1713] = ~(layer5_outputs[2150]) | (layer5_outputs[1625]);
    assign layer6_outputs[1714] = ~(layer5_outputs[1062]);
    assign layer6_outputs[1715] = layer5_outputs[4360];
    assign layer6_outputs[1716] = ~((layer5_outputs[3045]) & (layer5_outputs[1545]));
    assign layer6_outputs[1717] = ~(layer5_outputs[2215]);
    assign layer6_outputs[1718] = (layer5_outputs[4376]) & ~(layer5_outputs[1694]);
    assign layer6_outputs[1719] = layer5_outputs[989];
    assign layer6_outputs[1720] = (layer5_outputs[3324]) | (layer5_outputs[1053]);
    assign layer6_outputs[1721] = ~(layer5_outputs[4286]) | (layer5_outputs[3716]);
    assign layer6_outputs[1722] = ~((layer5_outputs[4004]) | (layer5_outputs[2885]));
    assign layer6_outputs[1723] = (layer5_outputs[2816]) ^ (layer5_outputs[515]);
    assign layer6_outputs[1724] = 1'b0;
    assign layer6_outputs[1725] = ~(layer5_outputs[4750]);
    assign layer6_outputs[1726] = (layer5_outputs[1824]) | (layer5_outputs[5069]);
    assign layer6_outputs[1727] = (layer5_outputs[4226]) & ~(layer5_outputs[1176]);
    assign layer6_outputs[1728] = ~(layer5_outputs[4046]) | (layer5_outputs[2361]);
    assign layer6_outputs[1729] = ~(layer5_outputs[3688]);
    assign layer6_outputs[1730] = layer5_outputs[800];
    assign layer6_outputs[1731] = ~(layer5_outputs[3126]);
    assign layer6_outputs[1732] = ~(layer5_outputs[4206]);
    assign layer6_outputs[1733] = ~(layer5_outputs[1929]) | (layer5_outputs[1464]);
    assign layer6_outputs[1734] = (layer5_outputs[256]) & ~(layer5_outputs[300]);
    assign layer6_outputs[1735] = ~(layer5_outputs[909]);
    assign layer6_outputs[1736] = ~(layer5_outputs[1621]);
    assign layer6_outputs[1737] = (layer5_outputs[1068]) ^ (layer5_outputs[3732]);
    assign layer6_outputs[1738] = (layer5_outputs[1185]) & ~(layer5_outputs[2133]);
    assign layer6_outputs[1739] = ~(layer5_outputs[341]);
    assign layer6_outputs[1740] = layer5_outputs[2267];
    assign layer6_outputs[1741] = (layer5_outputs[1464]) | (layer5_outputs[4640]);
    assign layer6_outputs[1742] = layer5_outputs[3724];
    assign layer6_outputs[1743] = ~(layer5_outputs[460]) | (layer5_outputs[2968]);
    assign layer6_outputs[1744] = (layer5_outputs[4376]) ^ (layer5_outputs[4573]);
    assign layer6_outputs[1745] = ~((layer5_outputs[2817]) ^ (layer5_outputs[4911]));
    assign layer6_outputs[1746] = (layer5_outputs[3484]) & ~(layer5_outputs[1179]);
    assign layer6_outputs[1747] = (layer5_outputs[2349]) & (layer5_outputs[2547]);
    assign layer6_outputs[1748] = layer5_outputs[2867];
    assign layer6_outputs[1749] = ~((layer5_outputs[161]) & (layer5_outputs[1795]));
    assign layer6_outputs[1750] = ~(layer5_outputs[1945]);
    assign layer6_outputs[1751] = ~((layer5_outputs[5025]) ^ (layer5_outputs[2885]));
    assign layer6_outputs[1752] = layer5_outputs[2506];
    assign layer6_outputs[1753] = ~(layer5_outputs[2001]);
    assign layer6_outputs[1754] = ~((layer5_outputs[936]) | (layer5_outputs[1687]));
    assign layer6_outputs[1755] = 1'b1;
    assign layer6_outputs[1756] = (layer5_outputs[4259]) & ~(layer5_outputs[3439]);
    assign layer6_outputs[1757] = ~((layer5_outputs[5095]) ^ (layer5_outputs[105]));
    assign layer6_outputs[1758] = 1'b0;
    assign layer6_outputs[1759] = ~((layer5_outputs[3744]) & (layer5_outputs[4463]));
    assign layer6_outputs[1760] = (layer5_outputs[664]) & ~(layer5_outputs[3630]);
    assign layer6_outputs[1761] = (layer5_outputs[2430]) ^ (layer5_outputs[231]);
    assign layer6_outputs[1762] = ~(layer5_outputs[1256]);
    assign layer6_outputs[1763] = (layer5_outputs[1902]) & (layer5_outputs[3365]);
    assign layer6_outputs[1764] = ~(layer5_outputs[4462]);
    assign layer6_outputs[1765] = ~(layer5_outputs[1568]);
    assign layer6_outputs[1766] = ~((layer5_outputs[2495]) ^ (layer5_outputs[423]));
    assign layer6_outputs[1767] = (layer5_outputs[667]) ^ (layer5_outputs[872]);
    assign layer6_outputs[1768] = (layer5_outputs[2269]) ^ (layer5_outputs[1404]);
    assign layer6_outputs[1769] = layer5_outputs[4440];
    assign layer6_outputs[1770] = (layer5_outputs[3270]) ^ (layer5_outputs[3267]);
    assign layer6_outputs[1771] = (layer5_outputs[2389]) & (layer5_outputs[4570]);
    assign layer6_outputs[1772] = (layer5_outputs[4530]) & (layer5_outputs[51]);
    assign layer6_outputs[1773] = ~((layer5_outputs[1981]) ^ (layer5_outputs[3482]));
    assign layer6_outputs[1774] = ~(layer5_outputs[3000]);
    assign layer6_outputs[1775] = ~(layer5_outputs[3278]) | (layer5_outputs[2716]);
    assign layer6_outputs[1776] = ~(layer5_outputs[754]);
    assign layer6_outputs[1777] = ~((layer5_outputs[760]) | (layer5_outputs[3181]));
    assign layer6_outputs[1778] = layer5_outputs[133];
    assign layer6_outputs[1779] = layer5_outputs[4713];
    assign layer6_outputs[1780] = ~(layer5_outputs[3337]);
    assign layer6_outputs[1781] = layer5_outputs[583];
    assign layer6_outputs[1782] = ~(layer5_outputs[3440]);
    assign layer6_outputs[1783] = (layer5_outputs[2726]) & ~(layer5_outputs[3699]);
    assign layer6_outputs[1784] = ~((layer5_outputs[4904]) | (layer5_outputs[786]));
    assign layer6_outputs[1785] = ~((layer5_outputs[992]) ^ (layer5_outputs[1449]));
    assign layer6_outputs[1786] = layer5_outputs[4554];
    assign layer6_outputs[1787] = ~((layer5_outputs[3895]) & (layer5_outputs[2091]));
    assign layer6_outputs[1788] = ~((layer5_outputs[3829]) ^ (layer5_outputs[4608]));
    assign layer6_outputs[1789] = layer5_outputs[4546];
    assign layer6_outputs[1790] = (layer5_outputs[3285]) & (layer5_outputs[4970]);
    assign layer6_outputs[1791] = layer5_outputs[2613];
    assign layer6_outputs[1792] = layer5_outputs[3506];
    assign layer6_outputs[1793] = ~(layer5_outputs[3812]);
    assign layer6_outputs[1794] = layer5_outputs[656];
    assign layer6_outputs[1795] = ~((layer5_outputs[2937]) | (layer5_outputs[296]));
    assign layer6_outputs[1796] = ~((layer5_outputs[2355]) ^ (layer5_outputs[3357]));
    assign layer6_outputs[1797] = layer5_outputs[1244];
    assign layer6_outputs[1798] = 1'b1;
    assign layer6_outputs[1799] = ~(layer5_outputs[1763]);
    assign layer6_outputs[1800] = ~(layer5_outputs[1544]);
    assign layer6_outputs[1801] = ~(layer5_outputs[789]);
    assign layer6_outputs[1802] = (layer5_outputs[416]) ^ (layer5_outputs[304]);
    assign layer6_outputs[1803] = (layer5_outputs[3882]) & ~(layer5_outputs[553]);
    assign layer6_outputs[1804] = (layer5_outputs[4520]) & ~(layer5_outputs[718]);
    assign layer6_outputs[1805] = ~(layer5_outputs[4609]) | (layer5_outputs[397]);
    assign layer6_outputs[1806] = ~((layer5_outputs[612]) & (layer5_outputs[2820]));
    assign layer6_outputs[1807] = ~((layer5_outputs[5068]) ^ (layer5_outputs[2658]));
    assign layer6_outputs[1808] = ~(layer5_outputs[1859]) | (layer5_outputs[667]);
    assign layer6_outputs[1809] = ~((layer5_outputs[4381]) ^ (layer5_outputs[761]));
    assign layer6_outputs[1810] = (layer5_outputs[4966]) ^ (layer5_outputs[1066]);
    assign layer6_outputs[1811] = layer5_outputs[1873];
    assign layer6_outputs[1812] = ~(layer5_outputs[4043]);
    assign layer6_outputs[1813] = layer5_outputs[1572];
    assign layer6_outputs[1814] = ~((layer5_outputs[3721]) | (layer5_outputs[4245]));
    assign layer6_outputs[1815] = layer5_outputs[1134];
    assign layer6_outputs[1816] = ~(layer5_outputs[4534]);
    assign layer6_outputs[1817] = layer5_outputs[919];
    assign layer6_outputs[1818] = layer5_outputs[4817];
    assign layer6_outputs[1819] = layer5_outputs[4243];
    assign layer6_outputs[1820] = ~(layer5_outputs[3087]);
    assign layer6_outputs[1821] = layer5_outputs[3334];
    assign layer6_outputs[1822] = layer5_outputs[340];
    assign layer6_outputs[1823] = layer5_outputs[1704];
    assign layer6_outputs[1824] = layer5_outputs[1601];
    assign layer6_outputs[1825] = ~(layer5_outputs[4724]) | (layer5_outputs[2743]);
    assign layer6_outputs[1826] = layer5_outputs[4437];
    assign layer6_outputs[1827] = ~((layer5_outputs[3320]) & (layer5_outputs[3668]));
    assign layer6_outputs[1828] = ~(layer5_outputs[4687]);
    assign layer6_outputs[1829] = (layer5_outputs[4938]) & (layer5_outputs[887]);
    assign layer6_outputs[1830] = ~(layer5_outputs[2470]) | (layer5_outputs[3587]);
    assign layer6_outputs[1831] = (layer5_outputs[2184]) & (layer5_outputs[2115]);
    assign layer6_outputs[1832] = layer5_outputs[1084];
    assign layer6_outputs[1833] = ~((layer5_outputs[3407]) ^ (layer5_outputs[2960]));
    assign layer6_outputs[1834] = (layer5_outputs[4929]) | (layer5_outputs[2456]);
    assign layer6_outputs[1835] = (layer5_outputs[603]) ^ (layer5_outputs[3880]);
    assign layer6_outputs[1836] = ~(layer5_outputs[577]);
    assign layer6_outputs[1837] = layer5_outputs[2004];
    assign layer6_outputs[1838] = 1'b0;
    assign layer6_outputs[1839] = (layer5_outputs[3529]) | (layer5_outputs[4075]);
    assign layer6_outputs[1840] = ~((layer5_outputs[1664]) ^ (layer5_outputs[879]));
    assign layer6_outputs[1841] = layer5_outputs[184];
    assign layer6_outputs[1842] = layer5_outputs[1561];
    assign layer6_outputs[1843] = (layer5_outputs[794]) & ~(layer5_outputs[4901]);
    assign layer6_outputs[1844] = ~((layer5_outputs[2177]) ^ (layer5_outputs[3508]));
    assign layer6_outputs[1845] = (layer5_outputs[181]) & ~(layer5_outputs[4281]);
    assign layer6_outputs[1846] = ~(layer5_outputs[912]);
    assign layer6_outputs[1847] = 1'b1;
    assign layer6_outputs[1848] = layer5_outputs[1304];
    assign layer6_outputs[1849] = ~(layer5_outputs[4412]);
    assign layer6_outputs[1850] = layer5_outputs[3781];
    assign layer6_outputs[1851] = ~(layer5_outputs[4289]);
    assign layer6_outputs[1852] = (layer5_outputs[2480]) ^ (layer5_outputs[1826]);
    assign layer6_outputs[1853] = (layer5_outputs[1821]) ^ (layer5_outputs[3135]);
    assign layer6_outputs[1854] = ~((layer5_outputs[1024]) ^ (layer5_outputs[4729]));
    assign layer6_outputs[1855] = layer5_outputs[1373];
    assign layer6_outputs[1856] = ~(layer5_outputs[4068]);
    assign layer6_outputs[1857] = (layer5_outputs[287]) ^ (layer5_outputs[248]);
    assign layer6_outputs[1858] = layer5_outputs[3406];
    assign layer6_outputs[1859] = ~(layer5_outputs[924]) | (layer5_outputs[1577]);
    assign layer6_outputs[1860] = layer5_outputs[4043];
    assign layer6_outputs[1861] = (layer5_outputs[2592]) ^ (layer5_outputs[4187]);
    assign layer6_outputs[1862] = (layer5_outputs[5029]) & ~(layer5_outputs[2611]);
    assign layer6_outputs[1863] = (layer5_outputs[511]) & (layer5_outputs[3724]);
    assign layer6_outputs[1864] = layer5_outputs[1751];
    assign layer6_outputs[1865] = layer5_outputs[1292];
    assign layer6_outputs[1866] = ~(layer5_outputs[1131]);
    assign layer6_outputs[1867] = ~((layer5_outputs[819]) ^ (layer5_outputs[4497]));
    assign layer6_outputs[1868] = layer5_outputs[739];
    assign layer6_outputs[1869] = (layer5_outputs[2155]) & ~(layer5_outputs[1896]);
    assign layer6_outputs[1870] = ~((layer5_outputs[2696]) ^ (layer5_outputs[4474]));
    assign layer6_outputs[1871] = layer5_outputs[794];
    assign layer6_outputs[1872] = layer5_outputs[2129];
    assign layer6_outputs[1873] = 1'b0;
    assign layer6_outputs[1874] = ~(layer5_outputs[1]);
    assign layer6_outputs[1875] = ~(layer5_outputs[831]);
    assign layer6_outputs[1876] = ~((layer5_outputs[4519]) ^ (layer5_outputs[1993]));
    assign layer6_outputs[1877] = ~((layer5_outputs[1288]) | (layer5_outputs[2358]));
    assign layer6_outputs[1878] = ~(layer5_outputs[1893]) | (layer5_outputs[1916]);
    assign layer6_outputs[1879] = ~(layer5_outputs[3151]);
    assign layer6_outputs[1880] = (layer5_outputs[627]) ^ (layer5_outputs[1521]);
    assign layer6_outputs[1881] = (layer5_outputs[3814]) & (layer5_outputs[1658]);
    assign layer6_outputs[1882] = ~(layer5_outputs[1018]) | (layer5_outputs[3036]);
    assign layer6_outputs[1883] = layer5_outputs[1275];
    assign layer6_outputs[1884] = layer5_outputs[4794];
    assign layer6_outputs[1885] = ~((layer5_outputs[4590]) ^ (layer5_outputs[222]));
    assign layer6_outputs[1886] = ~((layer5_outputs[361]) | (layer5_outputs[2259]));
    assign layer6_outputs[1887] = ~(layer5_outputs[4382]);
    assign layer6_outputs[1888] = layer5_outputs[1724];
    assign layer6_outputs[1889] = ~(layer5_outputs[5118]);
    assign layer6_outputs[1890] = layer5_outputs[201];
    assign layer6_outputs[1891] = 1'b0;
    assign layer6_outputs[1892] = (layer5_outputs[575]) & ~(layer5_outputs[470]);
    assign layer6_outputs[1893] = ~(layer5_outputs[333]) | (layer5_outputs[4384]);
    assign layer6_outputs[1894] = ~((layer5_outputs[880]) & (layer5_outputs[2193]));
    assign layer6_outputs[1895] = layer5_outputs[2261];
    assign layer6_outputs[1896] = ~(layer5_outputs[2811]) | (layer5_outputs[4757]);
    assign layer6_outputs[1897] = ~(layer5_outputs[1847]);
    assign layer6_outputs[1898] = layer5_outputs[4056];
    assign layer6_outputs[1899] = (layer5_outputs[4168]) ^ (layer5_outputs[717]);
    assign layer6_outputs[1900] = layer5_outputs[4489];
    assign layer6_outputs[1901] = ~((layer5_outputs[643]) | (layer5_outputs[1639]));
    assign layer6_outputs[1902] = ~(layer5_outputs[844]);
    assign layer6_outputs[1903] = layer5_outputs[1062];
    assign layer6_outputs[1904] = 1'b1;
    assign layer6_outputs[1905] = ~(layer5_outputs[5025]);
    assign layer6_outputs[1906] = ~(layer5_outputs[3818]);
    assign layer6_outputs[1907] = (layer5_outputs[3431]) ^ (layer5_outputs[4066]);
    assign layer6_outputs[1908] = ~(layer5_outputs[2222]);
    assign layer6_outputs[1909] = layer5_outputs[4318];
    assign layer6_outputs[1910] = ~(layer5_outputs[3978]);
    assign layer6_outputs[1911] = ~(layer5_outputs[1831]);
    assign layer6_outputs[1912] = layer5_outputs[4265];
    assign layer6_outputs[1913] = ~(layer5_outputs[3645]) | (layer5_outputs[3506]);
    assign layer6_outputs[1914] = layer5_outputs[377];
    assign layer6_outputs[1915] = layer5_outputs[575];
    assign layer6_outputs[1916] = layer5_outputs[460];
    assign layer6_outputs[1917] = (layer5_outputs[1233]) & (layer5_outputs[4406]);
    assign layer6_outputs[1918] = 1'b1;
    assign layer6_outputs[1919] = layer5_outputs[3228];
    assign layer6_outputs[1920] = ~((layer5_outputs[1069]) & (layer5_outputs[2926]));
    assign layer6_outputs[1921] = ~(layer5_outputs[3253]);
    assign layer6_outputs[1922] = ~((layer5_outputs[4628]) | (layer5_outputs[3720]));
    assign layer6_outputs[1923] = ~(layer5_outputs[805]);
    assign layer6_outputs[1924] = layer5_outputs[2897];
    assign layer6_outputs[1925] = ~(layer5_outputs[454]);
    assign layer6_outputs[1926] = (layer5_outputs[2346]) & ~(layer5_outputs[1771]);
    assign layer6_outputs[1927] = layer5_outputs[2794];
    assign layer6_outputs[1928] = ~(layer5_outputs[3641]);
    assign layer6_outputs[1929] = ~(layer5_outputs[1412]);
    assign layer6_outputs[1930] = ~(layer5_outputs[4586]);
    assign layer6_outputs[1931] = ~((layer5_outputs[2339]) ^ (layer5_outputs[3098]));
    assign layer6_outputs[1932] = (layer5_outputs[1606]) | (layer5_outputs[3386]);
    assign layer6_outputs[1933] = ~(layer5_outputs[4496]);
    assign layer6_outputs[1934] = ~(layer5_outputs[1292]);
    assign layer6_outputs[1935] = ~(layer5_outputs[482]) | (layer5_outputs[3311]);
    assign layer6_outputs[1936] = ~(layer5_outputs[593]);
    assign layer6_outputs[1937] = ~(layer5_outputs[4450]) | (layer5_outputs[4293]);
    assign layer6_outputs[1938] = ~(layer5_outputs[2287]) | (layer5_outputs[1603]);
    assign layer6_outputs[1939] = ~(layer5_outputs[2511]) | (layer5_outputs[1505]);
    assign layer6_outputs[1940] = ~(layer5_outputs[2175]);
    assign layer6_outputs[1941] = (layer5_outputs[3660]) ^ (layer5_outputs[2575]);
    assign layer6_outputs[1942] = (layer5_outputs[4406]) & ~(layer5_outputs[556]);
    assign layer6_outputs[1943] = ~(layer5_outputs[3679]);
    assign layer6_outputs[1944] = (layer5_outputs[3802]) & ~(layer5_outputs[2550]);
    assign layer6_outputs[1945] = (layer5_outputs[5115]) & (layer5_outputs[2037]);
    assign layer6_outputs[1946] = layer5_outputs[350];
    assign layer6_outputs[1947] = layer5_outputs[3061];
    assign layer6_outputs[1948] = ~(layer5_outputs[987]);
    assign layer6_outputs[1949] = (layer5_outputs[4734]) & ~(layer5_outputs[1166]);
    assign layer6_outputs[1950] = (layer5_outputs[2985]) ^ (layer5_outputs[3226]);
    assign layer6_outputs[1951] = layer5_outputs[4046];
    assign layer6_outputs[1952] = ~((layer5_outputs[3705]) ^ (layer5_outputs[927]));
    assign layer6_outputs[1953] = ~(layer5_outputs[698]) | (layer5_outputs[4442]);
    assign layer6_outputs[1954] = layer5_outputs[1653];
    assign layer6_outputs[1955] = ~(layer5_outputs[2520]);
    assign layer6_outputs[1956] = ~(layer5_outputs[1008]);
    assign layer6_outputs[1957] = layer5_outputs[4704];
    assign layer6_outputs[1958] = ~(layer5_outputs[4702]);
    assign layer6_outputs[1959] = layer5_outputs[4088];
    assign layer6_outputs[1960] = ~(layer5_outputs[4931]);
    assign layer6_outputs[1961] = ~(layer5_outputs[286]);
    assign layer6_outputs[1962] = (layer5_outputs[2728]) ^ (layer5_outputs[3713]);
    assign layer6_outputs[1963] = layer5_outputs[1778];
    assign layer6_outputs[1964] = (layer5_outputs[3692]) & ~(layer5_outputs[3603]);
    assign layer6_outputs[1965] = layer5_outputs[4704];
    assign layer6_outputs[1966] = ~(layer5_outputs[2114]) | (layer5_outputs[727]);
    assign layer6_outputs[1967] = ~(layer5_outputs[2861]);
    assign layer6_outputs[1968] = layer5_outputs[2710];
    assign layer6_outputs[1969] = (layer5_outputs[4940]) ^ (layer5_outputs[3229]);
    assign layer6_outputs[1970] = layer5_outputs[198];
    assign layer6_outputs[1971] = layer5_outputs[4547];
    assign layer6_outputs[1972] = ~((layer5_outputs[4290]) ^ (layer5_outputs[2514]));
    assign layer6_outputs[1973] = (layer5_outputs[2324]) & ~(layer5_outputs[5103]);
    assign layer6_outputs[1974] = layer5_outputs[996];
    assign layer6_outputs[1975] = ~((layer5_outputs[684]) ^ (layer5_outputs[1076]));
    assign layer6_outputs[1976] = layer5_outputs[5000];
    assign layer6_outputs[1977] = (layer5_outputs[2616]) | (layer5_outputs[3128]);
    assign layer6_outputs[1978] = layer5_outputs[2277];
    assign layer6_outputs[1979] = layer5_outputs[1474];
    assign layer6_outputs[1980] = layer5_outputs[2606];
    assign layer6_outputs[1981] = (layer5_outputs[3705]) & ~(layer5_outputs[2431]);
    assign layer6_outputs[1982] = (layer5_outputs[4407]) & ~(layer5_outputs[4109]);
    assign layer6_outputs[1983] = 1'b0;
    assign layer6_outputs[1984] = (layer5_outputs[4141]) & ~(layer5_outputs[2682]);
    assign layer6_outputs[1985] = layer5_outputs[1946];
    assign layer6_outputs[1986] = ~(layer5_outputs[753]);
    assign layer6_outputs[1987] = ~(layer5_outputs[3473]);
    assign layer6_outputs[1988] = layer5_outputs[2908];
    assign layer6_outputs[1989] = ~(layer5_outputs[2852]);
    assign layer6_outputs[1990] = ~(layer5_outputs[4996]);
    assign layer6_outputs[1991] = layer5_outputs[672];
    assign layer6_outputs[1992] = ~((layer5_outputs[2450]) | (layer5_outputs[1045]));
    assign layer6_outputs[1993] = ~(layer5_outputs[380]) | (layer5_outputs[2915]);
    assign layer6_outputs[1994] = ~(layer5_outputs[375]);
    assign layer6_outputs[1995] = ~(layer5_outputs[3239]);
    assign layer6_outputs[1996] = layer5_outputs[4147];
    assign layer6_outputs[1997] = (layer5_outputs[1495]) ^ (layer5_outputs[2868]);
    assign layer6_outputs[1998] = (layer5_outputs[2762]) ^ (layer5_outputs[4559]);
    assign layer6_outputs[1999] = (layer5_outputs[2036]) ^ (layer5_outputs[109]);
    assign layer6_outputs[2000] = ~((layer5_outputs[1575]) & (layer5_outputs[2151]));
    assign layer6_outputs[2001] = layer5_outputs[2939];
    assign layer6_outputs[2002] = layer5_outputs[4221];
    assign layer6_outputs[2003] = ~((layer5_outputs[4890]) ^ (layer5_outputs[3516]));
    assign layer6_outputs[2004] = layer5_outputs[4050];
    assign layer6_outputs[2005] = ~((layer5_outputs[3384]) ^ (layer5_outputs[2866]));
    assign layer6_outputs[2006] = ~(layer5_outputs[1583]);
    assign layer6_outputs[2007] = ~((layer5_outputs[3480]) | (layer5_outputs[3074]));
    assign layer6_outputs[2008] = layer5_outputs[2012];
    assign layer6_outputs[2009] = ~((layer5_outputs[1374]) | (layer5_outputs[4555]));
    assign layer6_outputs[2010] = ~(layer5_outputs[1552]);
    assign layer6_outputs[2011] = layer5_outputs[4879];
    assign layer6_outputs[2012] = layer5_outputs[3496];
    assign layer6_outputs[2013] = ~(layer5_outputs[4928]);
    assign layer6_outputs[2014] = layer5_outputs[5005];
    assign layer6_outputs[2015] = ~(layer5_outputs[4044]);
    assign layer6_outputs[2016] = 1'b1;
    assign layer6_outputs[2017] = (layer5_outputs[3762]) & (layer5_outputs[788]);
    assign layer6_outputs[2018] = ~((layer5_outputs[2459]) ^ (layer5_outputs[2634]));
    assign layer6_outputs[2019] = ~((layer5_outputs[610]) ^ (layer5_outputs[2649]));
    assign layer6_outputs[2020] = (layer5_outputs[2736]) | (layer5_outputs[2519]);
    assign layer6_outputs[2021] = ~((layer5_outputs[3471]) & (layer5_outputs[2390]));
    assign layer6_outputs[2022] = ~((layer5_outputs[1341]) ^ (layer5_outputs[1934]));
    assign layer6_outputs[2023] = ~(layer5_outputs[3116]);
    assign layer6_outputs[2024] = layer5_outputs[768];
    assign layer6_outputs[2025] = 1'b0;
    assign layer6_outputs[2026] = layer5_outputs[1815];
    assign layer6_outputs[2027] = layer5_outputs[3849];
    assign layer6_outputs[2028] = layer5_outputs[4411];
    assign layer6_outputs[2029] = ~((layer5_outputs[2134]) ^ (layer5_outputs[3642]));
    assign layer6_outputs[2030] = layer5_outputs[1268];
    assign layer6_outputs[2031] = ~(layer5_outputs[2314]);
    assign layer6_outputs[2032] = ~(layer5_outputs[3215]);
    assign layer6_outputs[2033] = ~(layer5_outputs[1165]);
    assign layer6_outputs[2034] = (layer5_outputs[3958]) & (layer5_outputs[3958]);
    assign layer6_outputs[2035] = layer5_outputs[50];
    assign layer6_outputs[2036] = layer5_outputs[462];
    assign layer6_outputs[2037] = layer5_outputs[4212];
    assign layer6_outputs[2038] = ~(layer5_outputs[2027]);
    assign layer6_outputs[2039] = (layer5_outputs[125]) & ~(layer5_outputs[486]);
    assign layer6_outputs[2040] = ~(layer5_outputs[466]);
    assign layer6_outputs[2041] = (layer5_outputs[1751]) ^ (layer5_outputs[1051]);
    assign layer6_outputs[2042] = ~(layer5_outputs[3595]);
    assign layer6_outputs[2043] = ~(layer5_outputs[3266]) | (layer5_outputs[1504]);
    assign layer6_outputs[2044] = ~((layer5_outputs[633]) & (layer5_outputs[2225]));
    assign layer6_outputs[2045] = ~((layer5_outputs[3205]) ^ (layer5_outputs[3789]));
    assign layer6_outputs[2046] = ~(layer5_outputs[3102]);
    assign layer6_outputs[2047] = layer5_outputs[4943];
    assign layer6_outputs[2048] = ~(layer5_outputs[4177]);
    assign layer6_outputs[2049] = ~(layer5_outputs[2049]);
    assign layer6_outputs[2050] = 1'b0;
    assign layer6_outputs[2051] = ~(layer5_outputs[2173]);
    assign layer6_outputs[2052] = ~((layer5_outputs[580]) ^ (layer5_outputs[3259]));
    assign layer6_outputs[2053] = ~(layer5_outputs[585]) | (layer5_outputs[5007]);
    assign layer6_outputs[2054] = (layer5_outputs[4618]) & ~(layer5_outputs[2745]);
    assign layer6_outputs[2055] = (layer5_outputs[4349]) ^ (layer5_outputs[1895]);
    assign layer6_outputs[2056] = layer5_outputs[4742];
    assign layer6_outputs[2057] = (layer5_outputs[4401]) ^ (layer5_outputs[1108]);
    assign layer6_outputs[2058] = ~(layer5_outputs[2466]);
    assign layer6_outputs[2059] = layer5_outputs[2680];
    assign layer6_outputs[2060] = ~(layer5_outputs[5018]);
    assign layer6_outputs[2061] = layer5_outputs[4107];
    assign layer6_outputs[2062] = ~(layer5_outputs[404]);
    assign layer6_outputs[2063] = ~(layer5_outputs[2943]);
    assign layer6_outputs[2064] = (layer5_outputs[4531]) & ~(layer5_outputs[3309]);
    assign layer6_outputs[2065] = ~(layer5_outputs[2673]) | (layer5_outputs[969]);
    assign layer6_outputs[2066] = ~(layer5_outputs[1371]);
    assign layer6_outputs[2067] = layer5_outputs[4104];
    assign layer6_outputs[2068] = (layer5_outputs[1356]) ^ (layer5_outputs[217]);
    assign layer6_outputs[2069] = (layer5_outputs[4795]) & (layer5_outputs[2700]);
    assign layer6_outputs[2070] = (layer5_outputs[1177]) ^ (layer5_outputs[4629]);
    assign layer6_outputs[2071] = ~((layer5_outputs[2963]) ^ (layer5_outputs[1415]));
    assign layer6_outputs[2072] = ~(layer5_outputs[3454]);
    assign layer6_outputs[2073] = ~((layer5_outputs[2660]) ^ (layer5_outputs[2065]));
    assign layer6_outputs[2074] = ~(layer5_outputs[3856]);
    assign layer6_outputs[2075] = (layer5_outputs[2476]) & (layer5_outputs[4922]);
    assign layer6_outputs[2076] = ~(layer5_outputs[4223]);
    assign layer6_outputs[2077] = (layer5_outputs[2740]) ^ (layer5_outputs[3177]);
    assign layer6_outputs[2078] = ~(layer5_outputs[3089]);
    assign layer6_outputs[2079] = (layer5_outputs[4545]) ^ (layer5_outputs[1833]);
    assign layer6_outputs[2080] = ~(layer5_outputs[2384]);
    assign layer6_outputs[2081] = ~((layer5_outputs[3621]) ^ (layer5_outputs[1579]));
    assign layer6_outputs[2082] = ~((layer5_outputs[2338]) ^ (layer5_outputs[2524]));
    assign layer6_outputs[2083] = (layer5_outputs[3462]) ^ (layer5_outputs[484]);
    assign layer6_outputs[2084] = (layer5_outputs[211]) ^ (layer5_outputs[1979]);
    assign layer6_outputs[2085] = ~(layer5_outputs[722]);
    assign layer6_outputs[2086] = layer5_outputs[4404];
    assign layer6_outputs[2087] = ~((layer5_outputs[4045]) & (layer5_outputs[3636]));
    assign layer6_outputs[2088] = ~(layer5_outputs[1470]);
    assign layer6_outputs[2089] = ~(layer5_outputs[3155]);
    assign layer6_outputs[2090] = (layer5_outputs[3263]) ^ (layer5_outputs[3020]);
    assign layer6_outputs[2091] = layer5_outputs[2979];
    assign layer6_outputs[2092] = ~(layer5_outputs[2792]) | (layer5_outputs[4980]);
    assign layer6_outputs[2093] = layer5_outputs[2163];
    assign layer6_outputs[2094] = (layer5_outputs[943]) & (layer5_outputs[4678]);
    assign layer6_outputs[2095] = (layer5_outputs[2518]) & ~(layer5_outputs[3323]);
    assign layer6_outputs[2096] = ~(layer5_outputs[4552]);
    assign layer6_outputs[2097] = layer5_outputs[2413];
    assign layer6_outputs[2098] = ~(layer5_outputs[2195]);
    assign layer6_outputs[2099] = (layer5_outputs[503]) ^ (layer5_outputs[2872]);
    assign layer6_outputs[2100] = ~((layer5_outputs[1546]) & (layer5_outputs[991]));
    assign layer6_outputs[2101] = ~(layer5_outputs[4617]);
    assign layer6_outputs[2102] = (layer5_outputs[200]) & (layer5_outputs[1867]);
    assign layer6_outputs[2103] = ~(layer5_outputs[1991]);
    assign layer6_outputs[2104] = ~(layer5_outputs[4391]) | (layer5_outputs[1911]);
    assign layer6_outputs[2105] = (layer5_outputs[3224]) ^ (layer5_outputs[1857]);
    assign layer6_outputs[2106] = ~((layer5_outputs[4676]) ^ (layer5_outputs[2660]));
    assign layer6_outputs[2107] = (layer5_outputs[973]) ^ (layer5_outputs[2343]);
    assign layer6_outputs[2108] = ~(layer5_outputs[838]);
    assign layer6_outputs[2109] = 1'b1;
    assign layer6_outputs[2110] = ~(layer5_outputs[4309]);
    assign layer6_outputs[2111] = layer5_outputs[3138];
    assign layer6_outputs[2112] = ~((layer5_outputs[3929]) ^ (layer5_outputs[4123]));
    assign layer6_outputs[2113] = layer5_outputs[2962];
    assign layer6_outputs[2114] = layer5_outputs[3143];
    assign layer6_outputs[2115] = layer5_outputs[4069];
    assign layer6_outputs[2116] = layer5_outputs[3786];
    assign layer6_outputs[2117] = 1'b1;
    assign layer6_outputs[2118] = layer5_outputs[4805];
    assign layer6_outputs[2119] = (layer5_outputs[943]) ^ (layer5_outputs[2749]);
    assign layer6_outputs[2120] = layer5_outputs[905];
    assign layer6_outputs[2121] = ~((layer5_outputs[4925]) ^ (layer5_outputs[3140]));
    assign layer6_outputs[2122] = layer5_outputs[1273];
    assign layer6_outputs[2123] = 1'b1;
    assign layer6_outputs[2124] = (layer5_outputs[660]) | (layer5_outputs[4101]);
    assign layer6_outputs[2125] = ~((layer5_outputs[4138]) & (layer5_outputs[3050]));
    assign layer6_outputs[2126] = ~(layer5_outputs[4518]) | (layer5_outputs[3281]);
    assign layer6_outputs[2127] = layer5_outputs[3021];
    assign layer6_outputs[2128] = layer5_outputs[506];
    assign layer6_outputs[2129] = ~(layer5_outputs[5016]);
    assign layer6_outputs[2130] = ~(layer5_outputs[2080]);
    assign layer6_outputs[2131] = layer5_outputs[2479];
    assign layer6_outputs[2132] = layer5_outputs[271];
    assign layer6_outputs[2133] = ~(layer5_outputs[3206]);
    assign layer6_outputs[2134] = ~(layer5_outputs[3313]) | (layer5_outputs[3305]);
    assign layer6_outputs[2135] = (layer5_outputs[1666]) & ~(layer5_outputs[3062]);
    assign layer6_outputs[2136] = ~(layer5_outputs[4362]) | (layer5_outputs[4425]);
    assign layer6_outputs[2137] = layer5_outputs[2438];
    assign layer6_outputs[2138] = layer5_outputs[552];
    assign layer6_outputs[2139] = ~(layer5_outputs[110]) | (layer5_outputs[3277]);
    assign layer6_outputs[2140] = ~(layer5_outputs[1274]) | (layer5_outputs[2560]);
    assign layer6_outputs[2141] = ~(layer5_outputs[2397]);
    assign layer6_outputs[2142] = ~(layer5_outputs[2563]);
    assign layer6_outputs[2143] = layer5_outputs[1123];
    assign layer6_outputs[2144] = ~((layer5_outputs[796]) ^ (layer5_outputs[3891]));
    assign layer6_outputs[2145] = ~(layer5_outputs[5021]) | (layer5_outputs[3223]);
    assign layer6_outputs[2146] = ~((layer5_outputs[1594]) ^ (layer5_outputs[3417]));
    assign layer6_outputs[2147] = (layer5_outputs[3066]) & ~(layer5_outputs[3389]);
    assign layer6_outputs[2148] = ~((layer5_outputs[2422]) ^ (layer5_outputs[123]));
    assign layer6_outputs[2149] = (layer5_outputs[396]) & ~(layer5_outputs[3773]);
    assign layer6_outputs[2150] = layer5_outputs[643];
    assign layer6_outputs[2151] = layer5_outputs[3245];
    assign layer6_outputs[2152] = layer5_outputs[2922];
    assign layer6_outputs[2153] = ~(layer5_outputs[4564]);
    assign layer6_outputs[2154] = ~(layer5_outputs[4339]);
    assign layer6_outputs[2155] = layer5_outputs[3240];
    assign layer6_outputs[2156] = ~(layer5_outputs[777]) | (layer5_outputs[635]);
    assign layer6_outputs[2157] = ~(layer5_outputs[905]);
    assign layer6_outputs[2158] = ~(layer5_outputs[4796]);
    assign layer6_outputs[2159] = layer5_outputs[3748];
    assign layer6_outputs[2160] = ~(layer5_outputs[4901]) | (layer5_outputs[2884]);
    assign layer6_outputs[2161] = (layer5_outputs[4400]) & ~(layer5_outputs[4844]);
    assign layer6_outputs[2162] = ~(layer5_outputs[3306]);
    assign layer6_outputs[2163] = ~(layer5_outputs[1766]);
    assign layer6_outputs[2164] = layer5_outputs[4021];
    assign layer6_outputs[2165] = 1'b1;
    assign layer6_outputs[2166] = (layer5_outputs[355]) & ~(layer5_outputs[2713]);
    assign layer6_outputs[2167] = layer5_outputs[2687];
    assign layer6_outputs[2168] = ~(layer5_outputs[2914]);
    assign layer6_outputs[2169] = layer5_outputs[302];
    assign layer6_outputs[2170] = ~(layer5_outputs[3460]) | (layer5_outputs[3546]);
    assign layer6_outputs[2171] = ~(layer5_outputs[847]);
    assign layer6_outputs[2172] = ~((layer5_outputs[3049]) | (layer5_outputs[4545]));
    assign layer6_outputs[2173] = layer5_outputs[2590];
    assign layer6_outputs[2174] = layer5_outputs[1633];
    assign layer6_outputs[2175] = (layer5_outputs[3434]) | (layer5_outputs[117]);
    assign layer6_outputs[2176] = ~(layer5_outputs[3137]);
    assign layer6_outputs[2177] = layer5_outputs[284];
    assign layer6_outputs[2178] = ~((layer5_outputs[1946]) & (layer5_outputs[366]));
    assign layer6_outputs[2179] = ~((layer5_outputs[450]) & (layer5_outputs[332]));
    assign layer6_outputs[2180] = layer5_outputs[3046];
    assign layer6_outputs[2181] = layer5_outputs[4814];
    assign layer6_outputs[2182] = ~(layer5_outputs[4994]);
    assign layer6_outputs[2183] = layer5_outputs[4638];
    assign layer6_outputs[2184] = layer5_outputs[2530];
    assign layer6_outputs[2185] = layer5_outputs[4342];
    assign layer6_outputs[2186] = layer5_outputs[1914];
    assign layer6_outputs[2187] = layer5_outputs[4255];
    assign layer6_outputs[2188] = ~((layer5_outputs[4886]) | (layer5_outputs[1201]));
    assign layer6_outputs[2189] = (layer5_outputs[2236]) & ~(layer5_outputs[2877]);
    assign layer6_outputs[2190] = (layer5_outputs[1508]) | (layer5_outputs[1701]);
    assign layer6_outputs[2191] = layer5_outputs[405];
    assign layer6_outputs[2192] = layer5_outputs[2705];
    assign layer6_outputs[2193] = ~(layer5_outputs[365]);
    assign layer6_outputs[2194] = (layer5_outputs[323]) & (layer5_outputs[1285]);
    assign layer6_outputs[2195] = layer5_outputs[1199];
    assign layer6_outputs[2196] = ~(layer5_outputs[3708]);
    assign layer6_outputs[2197] = ~((layer5_outputs[2164]) & (layer5_outputs[617]));
    assign layer6_outputs[2198] = layer5_outputs[4575];
    assign layer6_outputs[2199] = layer5_outputs[3538];
    assign layer6_outputs[2200] = ~(layer5_outputs[4235]);
    assign layer6_outputs[2201] = (layer5_outputs[370]) ^ (layer5_outputs[4889]);
    assign layer6_outputs[2202] = layer5_outputs[3155];
    assign layer6_outputs[2203] = layer5_outputs[5058];
    assign layer6_outputs[2204] = layer5_outputs[4568];
    assign layer6_outputs[2205] = layer5_outputs[1152];
    assign layer6_outputs[2206] = ~((layer5_outputs[836]) ^ (layer5_outputs[4592]));
    assign layer6_outputs[2207] = ~((layer5_outputs[3030]) & (layer5_outputs[4021]));
    assign layer6_outputs[2208] = ~(layer5_outputs[2893]);
    assign layer6_outputs[2209] = (layer5_outputs[3667]) ^ (layer5_outputs[3642]);
    assign layer6_outputs[2210] = layer5_outputs[5109];
    assign layer6_outputs[2211] = (layer5_outputs[3185]) & ~(layer5_outputs[447]);
    assign layer6_outputs[2212] = 1'b0;
    assign layer6_outputs[2213] = (layer5_outputs[4338]) ^ (layer5_outputs[888]);
    assign layer6_outputs[2214] = (layer5_outputs[5088]) & ~(layer5_outputs[2133]);
    assign layer6_outputs[2215] = (layer5_outputs[191]) | (layer5_outputs[135]);
    assign layer6_outputs[2216] = ~(layer5_outputs[371]) | (layer5_outputs[1160]);
    assign layer6_outputs[2217] = ~((layer5_outputs[4402]) ^ (layer5_outputs[3117]));
    assign layer6_outputs[2218] = layer5_outputs[4962];
    assign layer6_outputs[2219] = layer5_outputs[90];
    assign layer6_outputs[2220] = (layer5_outputs[2858]) ^ (layer5_outputs[1765]);
    assign layer6_outputs[2221] = ~(layer5_outputs[2723]);
    assign layer6_outputs[2222] = ~(layer5_outputs[1802]) | (layer5_outputs[3134]);
    assign layer6_outputs[2223] = ~((layer5_outputs[1139]) ^ (layer5_outputs[3368]));
    assign layer6_outputs[2224] = layer5_outputs[3494];
    assign layer6_outputs[2225] = (layer5_outputs[848]) ^ (layer5_outputs[4034]);
    assign layer6_outputs[2226] = ~((layer5_outputs[1382]) ^ (layer5_outputs[713]));
    assign layer6_outputs[2227] = (layer5_outputs[4903]) & (layer5_outputs[5054]);
    assign layer6_outputs[2228] = (layer5_outputs[988]) ^ (layer5_outputs[4930]);
    assign layer6_outputs[2229] = ~(layer5_outputs[5074]);
    assign layer6_outputs[2230] = ~((layer5_outputs[5043]) | (layer5_outputs[493]));
    assign layer6_outputs[2231] = (layer5_outputs[1797]) & ~(layer5_outputs[3096]);
    assign layer6_outputs[2232] = (layer5_outputs[1598]) ^ (layer5_outputs[17]);
    assign layer6_outputs[2233] = (layer5_outputs[3352]) ^ (layer5_outputs[608]);
    assign layer6_outputs[2234] = ~((layer5_outputs[2123]) ^ (layer5_outputs[4706]));
    assign layer6_outputs[2235] = ~((layer5_outputs[2177]) ^ (layer5_outputs[2000]));
    assign layer6_outputs[2236] = ~(layer5_outputs[2305]) | (layer5_outputs[1733]);
    assign layer6_outputs[2237] = (layer5_outputs[3278]) ^ (layer5_outputs[693]);
    assign layer6_outputs[2238] = ~((layer5_outputs[783]) | (layer5_outputs[2328]));
    assign layer6_outputs[2239] = layer5_outputs[4922];
    assign layer6_outputs[2240] = ~(layer5_outputs[1564]);
    assign layer6_outputs[2241] = layer5_outputs[88];
    assign layer6_outputs[2242] = layer5_outputs[2391];
    assign layer6_outputs[2243] = ~(layer5_outputs[3317]);
    assign layer6_outputs[2244] = ~((layer5_outputs[3154]) & (layer5_outputs[342]));
    assign layer6_outputs[2245] = ~(layer5_outputs[5098]);
    assign layer6_outputs[2246] = ~((layer5_outputs[2638]) | (layer5_outputs[1704]));
    assign layer6_outputs[2247] = layer5_outputs[1333];
    assign layer6_outputs[2248] = layer5_outputs[1661];
    assign layer6_outputs[2249] = 1'b1;
    assign layer6_outputs[2250] = ~(layer5_outputs[135]);
    assign layer6_outputs[2251] = layer5_outputs[4116];
    assign layer6_outputs[2252] = ~(layer5_outputs[4134]);
    assign layer6_outputs[2253] = (layer5_outputs[1756]) ^ (layer5_outputs[3353]);
    assign layer6_outputs[2254] = (layer5_outputs[496]) ^ (layer5_outputs[3346]);
    assign layer6_outputs[2255] = layer5_outputs[4758];
    assign layer6_outputs[2256] = ~(layer5_outputs[2959]);
    assign layer6_outputs[2257] = ~(layer5_outputs[1481]);
    assign layer6_outputs[2258] = layer5_outputs[1273];
    assign layer6_outputs[2259] = layer5_outputs[1922];
    assign layer6_outputs[2260] = ~(layer5_outputs[1034]);
    assign layer6_outputs[2261] = layer5_outputs[3012];
    assign layer6_outputs[2262] = (layer5_outputs[2821]) & ~(layer5_outputs[3507]);
    assign layer6_outputs[2263] = layer5_outputs[4792];
    assign layer6_outputs[2264] = ~(layer5_outputs[1057]);
    assign layer6_outputs[2265] = layer5_outputs[3419];
    assign layer6_outputs[2266] = layer5_outputs[4773];
    assign layer6_outputs[2267] = layer5_outputs[278];
    assign layer6_outputs[2268] = ~(layer5_outputs[1350]);
    assign layer6_outputs[2269] = (layer5_outputs[1869]) ^ (layer5_outputs[4663]);
    assign layer6_outputs[2270] = ~((layer5_outputs[1487]) ^ (layer5_outputs[185]));
    assign layer6_outputs[2271] = layer5_outputs[1017];
    assign layer6_outputs[2272] = layer5_outputs[2577];
    assign layer6_outputs[2273] = ~(layer5_outputs[1003]);
    assign layer6_outputs[2274] = ~(layer5_outputs[661]);
    assign layer6_outputs[2275] = ~(layer5_outputs[3945]) | (layer5_outputs[4784]);
    assign layer6_outputs[2276] = layer5_outputs[122];
    assign layer6_outputs[2277] = layer5_outputs[648];
    assign layer6_outputs[2278] = (layer5_outputs[73]) & (layer5_outputs[2780]);
    assign layer6_outputs[2279] = (layer5_outputs[3022]) ^ (layer5_outputs[1598]);
    assign layer6_outputs[2280] = ~((layer5_outputs[3205]) ^ (layer5_outputs[2671]));
    assign layer6_outputs[2281] = ~(layer5_outputs[853]);
    assign layer6_outputs[2282] = (layer5_outputs[1031]) ^ (layer5_outputs[4258]);
    assign layer6_outputs[2283] = ~(layer5_outputs[252]);
    assign layer6_outputs[2284] = 1'b0;
    assign layer6_outputs[2285] = ~((layer5_outputs[1959]) ^ (layer5_outputs[4434]));
    assign layer6_outputs[2286] = ~(layer5_outputs[1670]);
    assign layer6_outputs[2287] = ~(layer5_outputs[451]);
    assign layer6_outputs[2288] = ~(layer5_outputs[2415]) | (layer5_outputs[1571]);
    assign layer6_outputs[2289] = (layer5_outputs[4599]) | (layer5_outputs[2439]);
    assign layer6_outputs[2290] = layer5_outputs[632];
    assign layer6_outputs[2291] = layer5_outputs[204];
    assign layer6_outputs[2292] = ~(layer5_outputs[1988]);
    assign layer6_outputs[2293] = ~(layer5_outputs[2767]);
    assign layer6_outputs[2294] = ~(layer5_outputs[2158]) | (layer5_outputs[4626]);
    assign layer6_outputs[2295] = ~(layer5_outputs[4493]) | (layer5_outputs[594]);
    assign layer6_outputs[2296] = (layer5_outputs[779]) & ~(layer5_outputs[3983]);
    assign layer6_outputs[2297] = (layer5_outputs[387]) | (layer5_outputs[4584]);
    assign layer6_outputs[2298] = (layer5_outputs[4281]) & ~(layer5_outputs[2298]);
    assign layer6_outputs[2299] = layer5_outputs[350];
    assign layer6_outputs[2300] = ~(layer5_outputs[4526]);
    assign layer6_outputs[2301] = (layer5_outputs[3429]) | (layer5_outputs[392]);
    assign layer6_outputs[2302] = 1'b1;
    assign layer6_outputs[2303] = ~(layer5_outputs[427]);
    assign layer6_outputs[2304] = layer5_outputs[329];
    assign layer6_outputs[2305] = ~(layer5_outputs[2406]);
    assign layer6_outputs[2306] = (layer5_outputs[4632]) & ~(layer5_outputs[2937]);
    assign layer6_outputs[2307] = layer5_outputs[3223];
    assign layer6_outputs[2308] = ~(layer5_outputs[2339]);
    assign layer6_outputs[2309] = (layer5_outputs[1912]) ^ (layer5_outputs[2265]);
    assign layer6_outputs[2310] = ~(layer5_outputs[1584]);
    assign layer6_outputs[2311] = ~(layer5_outputs[957]);
    assign layer6_outputs[2312] = ~((layer5_outputs[3607]) | (layer5_outputs[4202]));
    assign layer6_outputs[2313] = ~((layer5_outputs[2543]) ^ (layer5_outputs[1156]));
    assign layer6_outputs[2314] = ~(layer5_outputs[4747]);
    assign layer6_outputs[2315] = layer5_outputs[3521];
    assign layer6_outputs[2316] = layer5_outputs[4096];
    assign layer6_outputs[2317] = ~(layer5_outputs[4190]) | (layer5_outputs[4315]);
    assign layer6_outputs[2318] = (layer5_outputs[1459]) | (layer5_outputs[4636]);
    assign layer6_outputs[2319] = ~(layer5_outputs[1205]);
    assign layer6_outputs[2320] = ~(layer5_outputs[721]);
    assign layer6_outputs[2321] = ~(layer5_outputs[3473]) | (layer5_outputs[4478]);
    assign layer6_outputs[2322] = (layer5_outputs[677]) & ~(layer5_outputs[4712]);
    assign layer6_outputs[2323] = ~(layer5_outputs[2082]);
    assign layer6_outputs[2324] = layer5_outputs[654];
    assign layer6_outputs[2325] = (layer5_outputs[1552]) ^ (layer5_outputs[1855]);
    assign layer6_outputs[2326] = ~(layer5_outputs[4597]);
    assign layer6_outputs[2327] = ~((layer5_outputs[1612]) & (layer5_outputs[4]));
    assign layer6_outputs[2328] = layer5_outputs[1058];
    assign layer6_outputs[2329] = ~(layer5_outputs[1674]);
    assign layer6_outputs[2330] = layer5_outputs[3001];
    assign layer6_outputs[2331] = ~(layer5_outputs[2782]);
    assign layer6_outputs[2332] = (layer5_outputs[3547]) & (layer5_outputs[158]);
    assign layer6_outputs[2333] = 1'b1;
    assign layer6_outputs[2334] = (layer5_outputs[3057]) ^ (layer5_outputs[3864]);
    assign layer6_outputs[2335] = ~((layer5_outputs[3402]) ^ (layer5_outputs[4010]));
    assign layer6_outputs[2336] = (layer5_outputs[1986]) & ~(layer5_outputs[29]);
    assign layer6_outputs[2337] = ~((layer5_outputs[3794]) & (layer5_outputs[3468]));
    assign layer6_outputs[2338] = ~(layer5_outputs[469]);
    assign layer6_outputs[2339] = ~(layer5_outputs[1293]) | (layer5_outputs[1393]);
    assign layer6_outputs[2340] = layer5_outputs[1856];
    assign layer6_outputs[2341] = ~(layer5_outputs[3411]);
    assign layer6_outputs[2342] = layer5_outputs[2076];
    assign layer6_outputs[2343] = layer5_outputs[4195];
    assign layer6_outputs[2344] = ~(layer5_outputs[2333]);
    assign layer6_outputs[2345] = layer5_outputs[4698];
    assign layer6_outputs[2346] = layer5_outputs[401];
    assign layer6_outputs[2347] = layer5_outputs[4068];
    assign layer6_outputs[2348] = ~(layer5_outputs[2599]);
    assign layer6_outputs[2349] = ~(layer5_outputs[5016]);
    assign layer6_outputs[2350] = (layer5_outputs[2352]) ^ (layer5_outputs[4771]);
    assign layer6_outputs[2351] = layer5_outputs[712];
    assign layer6_outputs[2352] = ~(layer5_outputs[2991]);
    assign layer6_outputs[2353] = ~((layer5_outputs[4869]) ^ (layer5_outputs[1130]));
    assign layer6_outputs[2354] = layer5_outputs[2920];
    assign layer6_outputs[2355] = layer5_outputs[2069];
    assign layer6_outputs[2356] = ~(layer5_outputs[3206]);
    assign layer6_outputs[2357] = ~((layer5_outputs[4940]) | (layer5_outputs[1614]));
    assign layer6_outputs[2358] = ~((layer5_outputs[3670]) ^ (layer5_outputs[4855]));
    assign layer6_outputs[2359] = layer5_outputs[625];
    assign layer6_outputs[2360] = ~((layer5_outputs[1489]) ^ (layer5_outputs[3648]));
    assign layer6_outputs[2361] = ~((layer5_outputs[1817]) | (layer5_outputs[498]));
    assign layer6_outputs[2362] = ~(layer5_outputs[619]);
    assign layer6_outputs[2363] = ~(layer5_outputs[2457]);
    assign layer6_outputs[2364] = (layer5_outputs[65]) ^ (layer5_outputs[4426]);
    assign layer6_outputs[2365] = ~((layer5_outputs[5102]) & (layer5_outputs[1175]));
    assign layer6_outputs[2366] = (layer5_outputs[2443]) | (layer5_outputs[3925]);
    assign layer6_outputs[2367] = ~(layer5_outputs[1430]);
    assign layer6_outputs[2368] = ~((layer5_outputs[4892]) ^ (layer5_outputs[630]));
    assign layer6_outputs[2369] = ~(layer5_outputs[3633]) | (layer5_outputs[2358]);
    assign layer6_outputs[2370] = layer5_outputs[2117];
    assign layer6_outputs[2371] = ~(layer5_outputs[1749]) | (layer5_outputs[1775]);
    assign layer6_outputs[2372] = layer5_outputs[3061];
    assign layer6_outputs[2373] = layer5_outputs[2904];
    assign layer6_outputs[2374] = ~((layer5_outputs[1359]) ^ (layer5_outputs[3270]));
    assign layer6_outputs[2375] = layer5_outputs[4824];
    assign layer6_outputs[2376] = layer5_outputs[3399];
    assign layer6_outputs[2377] = ~(layer5_outputs[2383]);
    assign layer6_outputs[2378] = ~(layer5_outputs[4951]) | (layer5_outputs[3523]);
    assign layer6_outputs[2379] = (layer5_outputs[2801]) & ~(layer5_outputs[2455]);
    assign layer6_outputs[2380] = ~(layer5_outputs[1659]);
    assign layer6_outputs[2381] = ~((layer5_outputs[517]) ^ (layer5_outputs[4828]));
    assign layer6_outputs[2382] = (layer5_outputs[4554]) & (layer5_outputs[4707]);
    assign layer6_outputs[2383] = ~((layer5_outputs[1682]) & (layer5_outputs[2124]));
    assign layer6_outputs[2384] = ~(layer5_outputs[1595]) | (layer5_outputs[1811]);
    assign layer6_outputs[2385] = (layer5_outputs[4333]) ^ (layer5_outputs[4114]);
    assign layer6_outputs[2386] = layer5_outputs[1500];
    assign layer6_outputs[2387] = (layer5_outputs[571]) ^ (layer5_outputs[1510]);
    assign layer6_outputs[2388] = (layer5_outputs[4259]) & (layer5_outputs[631]);
    assign layer6_outputs[2389] = ~(layer5_outputs[90]) | (layer5_outputs[3285]);
    assign layer6_outputs[2390] = ~(layer5_outputs[249]) | (layer5_outputs[3709]);
    assign layer6_outputs[2391] = ~((layer5_outputs[3976]) | (layer5_outputs[4111]));
    assign layer6_outputs[2392] = (layer5_outputs[2323]) & (layer5_outputs[1447]);
    assign layer6_outputs[2393] = layer5_outputs[3097];
    assign layer6_outputs[2394] = ~(layer5_outputs[2839]);
    assign layer6_outputs[2395] = layer5_outputs[3175];
    assign layer6_outputs[2396] = (layer5_outputs[3447]) | (layer5_outputs[3340]);
    assign layer6_outputs[2397] = ~((layer5_outputs[1622]) ^ (layer5_outputs[1974]));
    assign layer6_outputs[2398] = (layer5_outputs[3910]) & ~(layer5_outputs[1200]);
    assign layer6_outputs[2399] = layer5_outputs[561];
    assign layer6_outputs[2400] = ~(layer5_outputs[1407]) | (layer5_outputs[1828]);
    assign layer6_outputs[2401] = layer5_outputs[4092];
    assign layer6_outputs[2402] = ~(layer5_outputs[555]) | (layer5_outputs[115]);
    assign layer6_outputs[2403] = layer5_outputs[4959];
    assign layer6_outputs[2404] = layer5_outputs[1898];
    assign layer6_outputs[2405] = layer5_outputs[3890];
    assign layer6_outputs[2406] = ~(layer5_outputs[4741]);
    assign layer6_outputs[2407] = (layer5_outputs[3554]) ^ (layer5_outputs[3276]);
    assign layer6_outputs[2408] = ~(layer5_outputs[3292]);
    assign layer6_outputs[2409] = layer5_outputs[4216];
    assign layer6_outputs[2410] = ~(layer5_outputs[2060]);
    assign layer6_outputs[2411] = layer5_outputs[672];
    assign layer6_outputs[2412] = ~((layer5_outputs[300]) | (layer5_outputs[1633]));
    assign layer6_outputs[2413] = ~(layer5_outputs[3201]) | (layer5_outputs[1668]);
    assign layer6_outputs[2414] = (layer5_outputs[164]) & ~(layer5_outputs[2015]);
    assign layer6_outputs[2415] = 1'b1;
    assign layer6_outputs[2416] = layer5_outputs[3222];
    assign layer6_outputs[2417] = (layer5_outputs[505]) & (layer5_outputs[5067]);
    assign layer6_outputs[2418] = (layer5_outputs[4668]) ^ (layer5_outputs[3599]);
    assign layer6_outputs[2419] = layer5_outputs[4773];
    assign layer6_outputs[2420] = (layer5_outputs[2641]) & ~(layer5_outputs[4414]);
    assign layer6_outputs[2421] = ~((layer5_outputs[2882]) ^ (layer5_outputs[3661]));
    assign layer6_outputs[2422] = ~((layer5_outputs[3735]) | (layer5_outputs[18]));
    assign layer6_outputs[2423] = ~((layer5_outputs[1320]) | (layer5_outputs[3525]));
    assign layer6_outputs[2424] = ~(layer5_outputs[4437]) | (layer5_outputs[4031]);
    assign layer6_outputs[2425] = 1'b1;
    assign layer6_outputs[2426] = ~(layer5_outputs[1676]) | (layer5_outputs[516]);
    assign layer6_outputs[2427] = (layer5_outputs[1836]) & ~(layer5_outputs[502]);
    assign layer6_outputs[2428] = (layer5_outputs[4942]) & (layer5_outputs[3815]);
    assign layer6_outputs[2429] = ~((layer5_outputs[159]) | (layer5_outputs[4424]));
    assign layer6_outputs[2430] = ~(layer5_outputs[2523]);
    assign layer6_outputs[2431] = ~(layer5_outputs[3974]);
    assign layer6_outputs[2432] = 1'b1;
    assign layer6_outputs[2433] = ~((layer5_outputs[1191]) ^ (layer5_outputs[1867]));
    assign layer6_outputs[2434] = (layer5_outputs[4060]) & ~(layer5_outputs[1002]);
    assign layer6_outputs[2435] = ~(layer5_outputs[2321]);
    assign layer6_outputs[2436] = ~(layer5_outputs[1177]);
    assign layer6_outputs[2437] = (layer5_outputs[1277]) | (layer5_outputs[1868]);
    assign layer6_outputs[2438] = ~(layer5_outputs[3428]);
    assign layer6_outputs[2439] = (layer5_outputs[3537]) | (layer5_outputs[4726]);
    assign layer6_outputs[2440] = ~(layer5_outputs[2140]);
    assign layer6_outputs[2441] = ~(layer5_outputs[5028]);
    assign layer6_outputs[2442] = ~(layer5_outputs[4118]);
    assign layer6_outputs[2443] = ~(layer5_outputs[4749]);
    assign layer6_outputs[2444] = (layer5_outputs[5057]) & (layer5_outputs[1331]);
    assign layer6_outputs[2445] = (layer5_outputs[1061]) | (layer5_outputs[1505]);
    assign layer6_outputs[2446] = (layer5_outputs[4905]) ^ (layer5_outputs[2278]);
    assign layer6_outputs[2447] = layer5_outputs[3980];
    assign layer6_outputs[2448] = ~(layer5_outputs[2831]);
    assign layer6_outputs[2449] = (layer5_outputs[1705]) & (layer5_outputs[76]);
    assign layer6_outputs[2450] = layer5_outputs[3543];
    assign layer6_outputs[2451] = ~((layer5_outputs[1889]) | (layer5_outputs[5051]));
    assign layer6_outputs[2452] = layer5_outputs[2777];
    assign layer6_outputs[2453] = layer5_outputs[3821];
    assign layer6_outputs[2454] = (layer5_outputs[3203]) & ~(layer5_outputs[1445]);
    assign layer6_outputs[2455] = layer5_outputs[2621];
    assign layer6_outputs[2456] = ~(layer5_outputs[1662]);
    assign layer6_outputs[2457] = ~(layer5_outputs[4283]);
    assign layer6_outputs[2458] = layer5_outputs[2761];
    assign layer6_outputs[2459] = layer5_outputs[3745];
    assign layer6_outputs[2460] = layer5_outputs[993];
    assign layer6_outputs[2461] = layer5_outputs[4932];
    assign layer6_outputs[2462] = layer5_outputs[2856];
    assign layer6_outputs[2463] = layer5_outputs[1012];
    assign layer6_outputs[2464] = ~(layer5_outputs[3842]);
    assign layer6_outputs[2465] = layer5_outputs[2205];
    assign layer6_outputs[2466] = ~(layer5_outputs[2631]);
    assign layer6_outputs[2467] = layer5_outputs[3727];
    assign layer6_outputs[2468] = ~((layer5_outputs[4683]) ^ (layer5_outputs[2234]));
    assign layer6_outputs[2469] = layer5_outputs[3318];
    assign layer6_outputs[2470] = (layer5_outputs[1691]) & (layer5_outputs[2536]);
    assign layer6_outputs[2471] = layer5_outputs[4097];
    assign layer6_outputs[2472] = (layer5_outputs[4586]) & ~(layer5_outputs[2533]);
    assign layer6_outputs[2473] = (layer5_outputs[3348]) ^ (layer5_outputs[2407]);
    assign layer6_outputs[2474] = ~(layer5_outputs[1618]);
    assign layer6_outputs[2475] = (layer5_outputs[4667]) ^ (layer5_outputs[26]);
    assign layer6_outputs[2476] = (layer5_outputs[2608]) & (layer5_outputs[804]);
    assign layer6_outputs[2477] = layer5_outputs[1334];
    assign layer6_outputs[2478] = (layer5_outputs[4538]) & ~(layer5_outputs[3846]);
    assign layer6_outputs[2479] = (layer5_outputs[184]) | (layer5_outputs[1703]);
    assign layer6_outputs[2480] = layer5_outputs[1244];
    assign layer6_outputs[2481] = (layer5_outputs[4551]) & (layer5_outputs[2189]);
    assign layer6_outputs[2482] = ~(layer5_outputs[2656]);
    assign layer6_outputs[2483] = ~((layer5_outputs[1789]) | (layer5_outputs[1922]));
    assign layer6_outputs[2484] = ~(layer5_outputs[3664]);
    assign layer6_outputs[2485] = (layer5_outputs[4697]) & ~(layer5_outputs[5081]);
    assign layer6_outputs[2486] = layer5_outputs[3609];
    assign layer6_outputs[2487] = ~(layer5_outputs[3723]) | (layer5_outputs[2798]);
    assign layer6_outputs[2488] = (layer5_outputs[1483]) & ~(layer5_outputs[3025]);
    assign layer6_outputs[2489] = ~((layer5_outputs[615]) & (layer5_outputs[2655]));
    assign layer6_outputs[2490] = ~(layer5_outputs[4804]) | (layer5_outputs[4658]);
    assign layer6_outputs[2491] = 1'b0;
    assign layer6_outputs[2492] = layer5_outputs[1753];
    assign layer6_outputs[2493] = ~(layer5_outputs[1296]);
    assign layer6_outputs[2494] = ~(layer5_outputs[2688]);
    assign layer6_outputs[2495] = ~((layer5_outputs[4144]) & (layer5_outputs[3991]));
    assign layer6_outputs[2496] = ~(layer5_outputs[3071]);
    assign layer6_outputs[2497] = layer5_outputs[2587];
    assign layer6_outputs[2498] = (layer5_outputs[4464]) ^ (layer5_outputs[3047]);
    assign layer6_outputs[2499] = (layer5_outputs[3583]) & ~(layer5_outputs[654]);
    assign layer6_outputs[2500] = ~(layer5_outputs[1028]);
    assign layer6_outputs[2501] = ~(layer5_outputs[4044]) | (layer5_outputs[5034]);
    assign layer6_outputs[2502] = layer5_outputs[4039];
    assign layer6_outputs[2503] = ~(layer5_outputs[2126]);
    assign layer6_outputs[2504] = ~((layer5_outputs[2610]) | (layer5_outputs[220]));
    assign layer6_outputs[2505] = 1'b1;
    assign layer6_outputs[2506] = layer5_outputs[746];
    assign layer6_outputs[2507] = ~(layer5_outputs[2733]);
    assign layer6_outputs[2508] = ~((layer5_outputs[2319]) ^ (layer5_outputs[3483]));
    assign layer6_outputs[2509] = (layer5_outputs[4565]) | (layer5_outputs[72]);
    assign layer6_outputs[2510] = (layer5_outputs[3924]) & ~(layer5_outputs[4977]);
    assign layer6_outputs[2511] = ~(layer5_outputs[1350]);
    assign layer6_outputs[2512] = ~(layer5_outputs[4669]);
    assign layer6_outputs[2513] = ~((layer5_outputs[4532]) ^ (layer5_outputs[1869]));
    assign layer6_outputs[2514] = ~(layer5_outputs[3119]);
    assign layer6_outputs[2515] = layer5_outputs[4515];
    assign layer6_outputs[2516] = ~(layer5_outputs[2528]) | (layer5_outputs[4454]);
    assign layer6_outputs[2517] = ~(layer5_outputs[4981]);
    assign layer6_outputs[2518] = ~(layer5_outputs[3440]) | (layer5_outputs[3282]);
    assign layer6_outputs[2519] = layer5_outputs[1444];
    assign layer6_outputs[2520] = ~(layer5_outputs[4606]);
    assign layer6_outputs[2521] = (layer5_outputs[828]) & (layer5_outputs[4171]);
    assign layer6_outputs[2522] = ~(layer5_outputs[4284]);
    assign layer6_outputs[2523] = layer5_outputs[274];
    assign layer6_outputs[2524] = ~(layer5_outputs[4208]) | (layer5_outputs[4548]);
    assign layer6_outputs[2525] = ~(layer5_outputs[1628]);
    assign layer6_outputs[2526] = layer5_outputs[4135];
    assign layer6_outputs[2527] = ~((layer5_outputs[3446]) | (layer5_outputs[523]));
    assign layer6_outputs[2528] = ~(layer5_outputs[3192]);
    assign layer6_outputs[2529] = layer5_outputs[1000];
    assign layer6_outputs[2530] = (layer5_outputs[3592]) ^ (layer5_outputs[2896]);
    assign layer6_outputs[2531] = layer5_outputs[2912];
    assign layer6_outputs[2532] = ~(layer5_outputs[4899]) | (layer5_outputs[2035]);
    assign layer6_outputs[2533] = layer5_outputs[4613];
    assign layer6_outputs[2534] = layer5_outputs[4164];
    assign layer6_outputs[2535] = layer5_outputs[4839];
    assign layer6_outputs[2536] = layer5_outputs[106];
    assign layer6_outputs[2537] = (layer5_outputs[2448]) ^ (layer5_outputs[2632]);
    assign layer6_outputs[2538] = (layer5_outputs[923]) & (layer5_outputs[2255]);
    assign layer6_outputs[2539] = ~(layer5_outputs[847]);
    assign layer6_outputs[2540] = (layer5_outputs[3745]) | (layer5_outputs[4453]);
    assign layer6_outputs[2541] = ~(layer5_outputs[3904]);
    assign layer6_outputs[2542] = ~(layer5_outputs[3555]);
    assign layer6_outputs[2543] = ~(layer5_outputs[2290]);
    assign layer6_outputs[2544] = layer5_outputs[4909];
    assign layer6_outputs[2545] = ~((layer5_outputs[1611]) ^ (layer5_outputs[4209]));
    assign layer6_outputs[2546] = layer5_outputs[3537];
    assign layer6_outputs[2547] = ~(layer5_outputs[2003]) | (layer5_outputs[104]);
    assign layer6_outputs[2548] = 1'b0;
    assign layer6_outputs[2549] = ~(layer5_outputs[2132]);
    assign layer6_outputs[2550] = (layer5_outputs[3056]) ^ (layer5_outputs[2550]);
    assign layer6_outputs[2551] = layer5_outputs[1539];
    assign layer6_outputs[2552] = layer5_outputs[855];
    assign layer6_outputs[2553] = ~((layer5_outputs[1634]) ^ (layer5_outputs[1065]));
    assign layer6_outputs[2554] = layer5_outputs[2776];
    assign layer6_outputs[2555] = ~(layer5_outputs[11]) | (layer5_outputs[3240]);
    assign layer6_outputs[2556] = layer5_outputs[4113];
    assign layer6_outputs[2557] = (layer5_outputs[5080]) & ~(layer5_outputs[568]);
    assign layer6_outputs[2558] = ~(layer5_outputs[1908]) | (layer5_outputs[1642]);
    assign layer6_outputs[2559] = ~(layer5_outputs[1128]);
    assign layer6_outputs[2560] = (layer5_outputs[3969]) & (layer5_outputs[1391]);
    assign layer6_outputs[2561] = (layer5_outputs[1357]) & (layer5_outputs[2233]);
    assign layer6_outputs[2562] = layer5_outputs[4236];
    assign layer6_outputs[2563] = ~(layer5_outputs[343]) | (layer5_outputs[1029]);
    assign layer6_outputs[2564] = (layer5_outputs[1140]) | (layer5_outputs[3965]);
    assign layer6_outputs[2565] = (layer5_outputs[3451]) ^ (layer5_outputs[2169]);
    assign layer6_outputs[2566] = ~(layer5_outputs[559]);
    assign layer6_outputs[2567] = layer5_outputs[3712];
    assign layer6_outputs[2568] = (layer5_outputs[1392]) ^ (layer5_outputs[2206]);
    assign layer6_outputs[2569] = layer5_outputs[1210];
    assign layer6_outputs[2570] = layer5_outputs[2510];
    assign layer6_outputs[2571] = ~(layer5_outputs[2109]);
    assign layer6_outputs[2572] = (layer5_outputs[3486]) ^ (layer5_outputs[2597]);
    assign layer6_outputs[2573] = ~(layer5_outputs[2996]) | (layer5_outputs[4690]);
    assign layer6_outputs[2574] = layer5_outputs[858];
    assign layer6_outputs[2575] = ~(layer5_outputs[412]);
    assign layer6_outputs[2576] = ~((layer5_outputs[3862]) ^ (layer5_outputs[1711]));
    assign layer6_outputs[2577] = layer5_outputs[2538];
    assign layer6_outputs[2578] = layer5_outputs[4220];
    assign layer6_outputs[2579] = ~(layer5_outputs[4694]) | (layer5_outputs[2760]);
    assign layer6_outputs[2580] = ~(layer5_outputs[3135]);
    assign layer6_outputs[2581] = ~(layer5_outputs[652]);
    assign layer6_outputs[2582] = ~((layer5_outputs[5045]) ^ (layer5_outputs[5090]));
    assign layer6_outputs[2583] = ~((layer5_outputs[767]) | (layer5_outputs[2594]));
    assign layer6_outputs[2584] = (layer5_outputs[3362]) & ~(layer5_outputs[899]);
    assign layer6_outputs[2585] = ~(layer5_outputs[2745]);
    assign layer6_outputs[2586] = (layer5_outputs[1149]) & ~(layer5_outputs[1102]);
    assign layer6_outputs[2587] = ~(layer5_outputs[1631]);
    assign layer6_outputs[2588] = ~(layer5_outputs[4866]);
    assign layer6_outputs[2589] = ~(layer5_outputs[2030]);
    assign layer6_outputs[2590] = (layer5_outputs[3824]) & ~(layer5_outputs[3612]);
    assign layer6_outputs[2591] = ~(layer5_outputs[298]);
    assign layer6_outputs[2592] = layer5_outputs[2052];
    assign layer6_outputs[2593] = ~(layer5_outputs[3049]);
    assign layer6_outputs[2594] = ~((layer5_outputs[1532]) ^ (layer5_outputs[4639]));
    assign layer6_outputs[2595] = layer5_outputs[4447];
    assign layer6_outputs[2596] = (layer5_outputs[3225]) & ~(layer5_outputs[823]);
    assign layer6_outputs[2597] = (layer5_outputs[2686]) ^ (layer5_outputs[2929]);
    assign layer6_outputs[2598] = (layer5_outputs[3210]) ^ (layer5_outputs[3888]);
    assign layer6_outputs[2599] = (layer5_outputs[829]) ^ (layer5_outputs[2273]);
    assign layer6_outputs[2600] = layer5_outputs[752];
    assign layer6_outputs[2601] = (layer5_outputs[3498]) & ~(layer5_outputs[3055]);
    assign layer6_outputs[2602] = layer5_outputs[2957];
    assign layer6_outputs[2603] = ~((layer5_outputs[1560]) | (layer5_outputs[1077]));
    assign layer6_outputs[2604] = ~((layer5_outputs[1455]) ^ (layer5_outputs[296]));
    assign layer6_outputs[2605] = layer5_outputs[1170];
    assign layer6_outputs[2606] = ~((layer5_outputs[5013]) ^ (layer5_outputs[2851]));
    assign layer6_outputs[2607] = ~(layer5_outputs[1655]);
    assign layer6_outputs[2608] = 1'b1;
    assign layer6_outputs[2609] = (layer5_outputs[388]) & ~(layer5_outputs[422]);
    assign layer6_outputs[2610] = layer5_outputs[3979];
    assign layer6_outputs[2611] = ~(layer5_outputs[4523]);
    assign layer6_outputs[2612] = ~(layer5_outputs[384]);
    assign layer6_outputs[2613] = layer5_outputs[1579];
    assign layer6_outputs[2614] = layer5_outputs[3035];
    assign layer6_outputs[2615] = 1'b0;
    assign layer6_outputs[2616] = layer5_outputs[906];
    assign layer6_outputs[2617] = layer5_outputs[5011];
    assign layer6_outputs[2618] = (layer5_outputs[3434]) & ~(layer5_outputs[4145]);
    assign layer6_outputs[2619] = layer5_outputs[4299];
    assign layer6_outputs[2620] = layer5_outputs[4024];
    assign layer6_outputs[2621] = (layer5_outputs[728]) & ~(layer5_outputs[4276]);
    assign layer6_outputs[2622] = 1'b1;
    assign layer6_outputs[2623] = ~(layer5_outputs[499]);
    assign layer6_outputs[2624] = ~(layer5_outputs[1069]);
    assign layer6_outputs[2625] = ~((layer5_outputs[4475]) & (layer5_outputs[4396]));
    assign layer6_outputs[2626] = ~((layer5_outputs[1618]) ^ (layer5_outputs[2653]));
    assign layer6_outputs[2627] = layer5_outputs[4891];
    assign layer6_outputs[2628] = layer5_outputs[250];
    assign layer6_outputs[2629] = (layer5_outputs[3227]) | (layer5_outputs[4033]);
    assign layer6_outputs[2630] = ~(layer5_outputs[3269]) | (layer5_outputs[4379]);
    assign layer6_outputs[2631] = (layer5_outputs[3758]) ^ (layer5_outputs[4651]);
    assign layer6_outputs[2632] = (layer5_outputs[4350]) | (layer5_outputs[4684]);
    assign layer6_outputs[2633] = layer5_outputs[1202];
    assign layer6_outputs[2634] = ~(layer5_outputs[3808]);
    assign layer6_outputs[2635] = layer5_outputs[52];
    assign layer6_outputs[2636] = (layer5_outputs[1478]) & ~(layer5_outputs[3741]);
    assign layer6_outputs[2637] = (layer5_outputs[2013]) & (layer5_outputs[2329]);
    assign layer6_outputs[2638] = ~(layer5_outputs[1175]);
    assign layer6_outputs[2639] = ~(layer5_outputs[4298]);
    assign layer6_outputs[2640] = (layer5_outputs[143]) & ~(layer5_outputs[3292]);
    assign layer6_outputs[2641] = ~(layer5_outputs[3678]);
    assign layer6_outputs[2642] = ~(layer5_outputs[1969]) | (layer5_outputs[3562]);
    assign layer6_outputs[2643] = ~(layer5_outputs[2289]);
    assign layer6_outputs[2644] = ~(layer5_outputs[3584]);
    assign layer6_outputs[2645] = layer5_outputs[4956];
    assign layer6_outputs[2646] = ~((layer5_outputs[3337]) & (layer5_outputs[4403]));
    assign layer6_outputs[2647] = ~(layer5_outputs[2520]);
    assign layer6_outputs[2648] = ~(layer5_outputs[3759]);
    assign layer6_outputs[2649] = ~(layer5_outputs[146]);
    assign layer6_outputs[2650] = (layer5_outputs[3685]) & ~(layer5_outputs[4567]);
    assign layer6_outputs[2651] = (layer5_outputs[802]) ^ (layer5_outputs[854]);
    assign layer6_outputs[2652] = layer5_outputs[5056];
    assign layer6_outputs[2653] = ~(layer5_outputs[2047]);
    assign layer6_outputs[2654] = ~(layer5_outputs[3159]);
    assign layer6_outputs[2655] = ~(layer5_outputs[2292]);
    assign layer6_outputs[2656] = layer5_outputs[1004];
    assign layer6_outputs[2657] = ~(layer5_outputs[1848]);
    assign layer6_outputs[2658] = ~((layer5_outputs[4309]) ^ (layer5_outputs[3234]));
    assign layer6_outputs[2659] = 1'b0;
    assign layer6_outputs[2660] = ~(layer5_outputs[993]);
    assign layer6_outputs[2661] = layer5_outputs[3267];
    assign layer6_outputs[2662] = ~(layer5_outputs[4251]) | (layer5_outputs[3390]);
    assign layer6_outputs[2663] = layer5_outputs[3316];
    assign layer6_outputs[2664] = ~((layer5_outputs[1541]) ^ (layer5_outputs[3100]));
    assign layer6_outputs[2665] = (layer5_outputs[2238]) & ~(layer5_outputs[997]);
    assign layer6_outputs[2666] = (layer5_outputs[2567]) & (layer5_outputs[4335]);
    assign layer6_outputs[2667] = ~(layer5_outputs[3920]) | (layer5_outputs[3837]);
    assign layer6_outputs[2668] = (layer5_outputs[2637]) & ~(layer5_outputs[3034]);
    assign layer6_outputs[2669] = ~(layer5_outputs[2818]);
    assign layer6_outputs[2670] = ~(layer5_outputs[4610]) | (layer5_outputs[1041]);
    assign layer6_outputs[2671] = layer5_outputs[4053];
    assign layer6_outputs[2672] = (layer5_outputs[582]) ^ (layer5_outputs[5082]);
    assign layer6_outputs[2673] = (layer5_outputs[1235]) ^ (layer5_outputs[4083]);
    assign layer6_outputs[2674] = (layer5_outputs[1424]) & ~(layer5_outputs[3031]);
    assign layer6_outputs[2675] = ~((layer5_outputs[2726]) ^ (layer5_outputs[235]));
    assign layer6_outputs[2676] = ~(layer5_outputs[4479]) | (layer5_outputs[3314]);
    assign layer6_outputs[2677] = ~(layer5_outputs[3167]);
    assign layer6_outputs[2678] = (layer5_outputs[409]) ^ (layer5_outputs[4612]);
    assign layer6_outputs[2679] = ~(layer5_outputs[877]);
    assign layer6_outputs[2680] = ~(layer5_outputs[4946]);
    assign layer6_outputs[2681] = ~(layer5_outputs[2183]);
    assign layer6_outputs[2682] = (layer5_outputs[2453]) & ~(layer5_outputs[4687]);
    assign layer6_outputs[2683] = layer5_outputs[4890];
    assign layer6_outputs[2684] = ~(layer5_outputs[189]);
    assign layer6_outputs[2685] = (layer5_outputs[324]) & (layer5_outputs[2087]);
    assign layer6_outputs[2686] = ~((layer5_outputs[4193]) ^ (layer5_outputs[732]));
    assign layer6_outputs[2687] = layer5_outputs[3087];
    assign layer6_outputs[2688] = ~(layer5_outputs[1416]);
    assign layer6_outputs[2689] = ~(layer5_outputs[266]);
    assign layer6_outputs[2690] = ~(layer5_outputs[2229]);
    assign layer6_outputs[2691] = layer5_outputs[4535];
    assign layer6_outputs[2692] = ~(layer5_outputs[1735]);
    assign layer6_outputs[2693] = ~((layer5_outputs[89]) ^ (layer5_outputs[3170]));
    assign layer6_outputs[2694] = (layer5_outputs[1658]) & ~(layer5_outputs[3144]);
    assign layer6_outputs[2695] = ~(layer5_outputs[3768]);
    assign layer6_outputs[2696] = (layer5_outputs[4717]) ^ (layer5_outputs[3757]);
    assign layer6_outputs[2697] = ~(layer5_outputs[1935]);
    assign layer6_outputs[2698] = ~((layer5_outputs[2718]) ^ (layer5_outputs[1301]));
    assign layer6_outputs[2699] = (layer5_outputs[3590]) & ~(layer5_outputs[345]);
    assign layer6_outputs[2700] = layer5_outputs[3279];
    assign layer6_outputs[2701] = ~((layer5_outputs[5026]) & (layer5_outputs[1656]));
    assign layer6_outputs[2702] = (layer5_outputs[132]) & ~(layer5_outputs[2482]);
    assign layer6_outputs[2703] = (layer5_outputs[1559]) & ~(layer5_outputs[3701]);
    assign layer6_outputs[2704] = ~(layer5_outputs[4142]);
    assign layer6_outputs[2705] = ~(layer5_outputs[4887]);
    assign layer6_outputs[2706] = ~(layer5_outputs[878]) | (layer5_outputs[38]);
    assign layer6_outputs[2707] = ~((layer5_outputs[1257]) ^ (layer5_outputs[4592]));
    assign layer6_outputs[2708] = layer5_outputs[3526];
    assign layer6_outputs[2709] = ~((layer5_outputs[202]) | (layer5_outputs[146]));
    assign layer6_outputs[2710] = ~(layer5_outputs[2222]);
    assign layer6_outputs[2711] = ~(layer5_outputs[27]);
    assign layer6_outputs[2712] = layer5_outputs[4077];
    assign layer6_outputs[2713] = ~(layer5_outputs[505]);
    assign layer6_outputs[2714] = ~(layer5_outputs[897]);
    assign layer6_outputs[2715] = ~((layer5_outputs[4759]) ^ (layer5_outputs[2204]));
    assign layer6_outputs[2716] = layer5_outputs[1197];
    assign layer6_outputs[2717] = ~((layer5_outputs[4945]) & (layer5_outputs[4770]));
    assign layer6_outputs[2718] = ~(layer5_outputs[4951]);
    assign layer6_outputs[2719] = layer5_outputs[1923];
    assign layer6_outputs[2720] = ~(layer5_outputs[241]) | (layer5_outputs[4679]);
    assign layer6_outputs[2721] = (layer5_outputs[4175]) ^ (layer5_outputs[3400]);
    assign layer6_outputs[2722] = layer5_outputs[1636];
    assign layer6_outputs[2723] = ~(layer5_outputs[862]) | (layer5_outputs[2679]);
    assign layer6_outputs[2724] = layer5_outputs[1885];
    assign layer6_outputs[2725] = (layer5_outputs[3617]) | (layer5_outputs[2521]);
    assign layer6_outputs[2726] = (layer5_outputs[2819]) & (layer5_outputs[4602]);
    assign layer6_outputs[2727] = layer5_outputs[3068];
    assign layer6_outputs[2728] = layer5_outputs[2217];
    assign layer6_outputs[2729] = ~(layer5_outputs[4942]);
    assign layer6_outputs[2730] = ~((layer5_outputs[3432]) ^ (layer5_outputs[2086]));
    assign layer6_outputs[2731] = (layer5_outputs[3658]) | (layer5_outputs[3163]);
    assign layer6_outputs[2732] = ~(layer5_outputs[1957]);
    assign layer6_outputs[2733] = ~(layer5_outputs[2200]);
    assign layer6_outputs[2734] = ~(layer5_outputs[3498]);
    assign layer6_outputs[2735] = ~(layer5_outputs[3532]);
    assign layer6_outputs[2736] = ~(layer5_outputs[956]) | (layer5_outputs[4601]);
    assign layer6_outputs[2737] = layer5_outputs[1052];
    assign layer6_outputs[2738] = (layer5_outputs[408]) ^ (layer5_outputs[4364]);
    assign layer6_outputs[2739] = (layer5_outputs[4923]) & (layer5_outputs[3727]);
    assign layer6_outputs[2740] = ~(layer5_outputs[1709]);
    assign layer6_outputs[2741] = layer5_outputs[1466];
    assign layer6_outputs[2742] = ~(layer5_outputs[3866]);
    assign layer6_outputs[2743] = ~(layer5_outputs[4176]);
    assign layer6_outputs[2744] = ~((layer5_outputs[5009]) | (layer5_outputs[4842]));
    assign layer6_outputs[2745] = (layer5_outputs[182]) & ~(layer5_outputs[4147]);
    assign layer6_outputs[2746] = layer5_outputs[1478];
    assign layer6_outputs[2747] = ~((layer5_outputs[5036]) ^ (layer5_outputs[4984]));
    assign layer6_outputs[2748] = (layer5_outputs[566]) & ~(layer5_outputs[1880]);
    assign layer6_outputs[2749] = (layer5_outputs[1729]) ^ (layer5_outputs[913]);
    assign layer6_outputs[2750] = layer5_outputs[821];
    assign layer6_outputs[2751] = layer5_outputs[976];
    assign layer6_outputs[2752] = ~(layer5_outputs[1446]);
    assign layer6_outputs[2753] = (layer5_outputs[1325]) ^ (layer5_outputs[3193]);
    assign layer6_outputs[2754] = ~(layer5_outputs[4327]);
    assign layer6_outputs[2755] = ~((layer5_outputs[3208]) & (layer5_outputs[3435]));
    assign layer6_outputs[2756] = layer5_outputs[3812];
    assign layer6_outputs[2757] = (layer5_outputs[2272]) & (layer5_outputs[2784]);
    assign layer6_outputs[2758] = ~(layer5_outputs[1217]) | (layer5_outputs[4285]);
    assign layer6_outputs[2759] = layer5_outputs[1602];
    assign layer6_outputs[2760] = ~(layer5_outputs[1615]) | (layer5_outputs[2497]);
    assign layer6_outputs[2761] = ~((layer5_outputs[1668]) ^ (layer5_outputs[982]));
    assign layer6_outputs[2762] = ~((layer5_outputs[2491]) ^ (layer5_outputs[4944]));
    assign layer6_outputs[2763] = (layer5_outputs[3198]) & ~(layer5_outputs[3780]);
    assign layer6_outputs[2764] = layer5_outputs[4587];
    assign layer6_outputs[2765] = layer5_outputs[1216];
    assign layer6_outputs[2766] = layer5_outputs[1078];
    assign layer6_outputs[2767] = layer5_outputs[513];
    assign layer6_outputs[2768] = ~((layer5_outputs[1971]) ^ (layer5_outputs[3902]));
    assign layer6_outputs[2769] = ~(layer5_outputs[3835]);
    assign layer6_outputs[2770] = layer5_outputs[1941];
    assign layer6_outputs[2771] = layer5_outputs[4819];
    assign layer6_outputs[2772] = ~((layer5_outputs[1787]) | (layer5_outputs[390]));
    assign layer6_outputs[2773] = ~((layer5_outputs[190]) & (layer5_outputs[2987]));
    assign layer6_outputs[2774] = layer5_outputs[4957];
    assign layer6_outputs[2775] = ~((layer5_outputs[595]) ^ (layer5_outputs[1518]));
    assign layer6_outputs[2776] = (layer5_outputs[105]) ^ (layer5_outputs[1022]);
    assign layer6_outputs[2777] = ~(layer5_outputs[2311]);
    assign layer6_outputs[2778] = layer5_outputs[3645];
    assign layer6_outputs[2779] = ~(layer5_outputs[3540]) | (layer5_outputs[4228]);
    assign layer6_outputs[2780] = ~((layer5_outputs[3381]) ^ (layer5_outputs[200]));
    assign layer6_outputs[2781] = ~((layer5_outputs[1962]) & (layer5_outputs[3157]));
    assign layer6_outputs[2782] = layer5_outputs[4343];
    assign layer6_outputs[2783] = ~(layer5_outputs[2549]) | (layer5_outputs[2307]);
    assign layer6_outputs[2784] = ~(layer5_outputs[1569]);
    assign layer6_outputs[2785] = ~((layer5_outputs[4561]) & (layer5_outputs[2153]));
    assign layer6_outputs[2786] = ~(layer5_outputs[1341]);
    assign layer6_outputs[2787] = ~(layer5_outputs[4989]);
    assign layer6_outputs[2788] = (layer5_outputs[531]) & ~(layer5_outputs[3719]);
    assign layer6_outputs[2789] = ~(layer5_outputs[4263]);
    assign layer6_outputs[2790] = (layer5_outputs[1932]) & (layer5_outputs[2923]);
    assign layer6_outputs[2791] = layer5_outputs[3260];
    assign layer6_outputs[2792] = (layer5_outputs[3501]) ^ (layer5_outputs[548]);
    assign layer6_outputs[2793] = (layer5_outputs[8]) | (layer5_outputs[2260]);
    assign layer6_outputs[2794] = layer5_outputs[703];
    assign layer6_outputs[2795] = ~((layer5_outputs[546]) ^ (layer5_outputs[2500]));
    assign layer6_outputs[2796] = 1'b1;
    assign layer6_outputs[2797] = (layer5_outputs[3284]) & ~(layer5_outputs[4920]);
    assign layer6_outputs[2798] = ~(layer5_outputs[4411]);
    assign layer6_outputs[2799] = (layer5_outputs[3079]) & (layer5_outputs[1888]);
    assign layer6_outputs[2800] = layer5_outputs[3200];
    assign layer6_outputs[2801] = 1'b0;
    assign layer6_outputs[2802] = ~((layer5_outputs[2649]) ^ (layer5_outputs[2139]));
    assign layer6_outputs[2803] = layer5_outputs[749];
    assign layer6_outputs[2804] = (layer5_outputs[2561]) & ~(layer5_outputs[1937]);
    assign layer6_outputs[2805] = ~(layer5_outputs[4557]) | (layer5_outputs[2853]);
    assign layer6_outputs[2806] = ~(layer5_outputs[1050]) | (layer5_outputs[2266]);
    assign layer6_outputs[2807] = ~(layer5_outputs[1262]);
    assign layer6_outputs[2808] = layer5_outputs[552];
    assign layer6_outputs[2809] = layer5_outputs[3973];
    assign layer6_outputs[2810] = layer5_outputs[4924];
    assign layer6_outputs[2811] = layer5_outputs[4837];
    assign layer6_outputs[2812] = (layer5_outputs[1146]) & ~(layer5_outputs[2980]);
    assign layer6_outputs[2813] = layer5_outputs[3793];
    assign layer6_outputs[2814] = ~((layer5_outputs[1421]) & (layer5_outputs[2141]));
    assign layer6_outputs[2815] = ~(layer5_outputs[1340]);
    assign layer6_outputs[2816] = ~(layer5_outputs[5082]);
    assign layer6_outputs[2817] = layer5_outputs[3715];
    assign layer6_outputs[2818] = (layer5_outputs[3624]) & ~(layer5_outputs[4183]);
    assign layer6_outputs[2819] = layer5_outputs[837];
    assign layer6_outputs[2820] = 1'b0;
    assign layer6_outputs[2821] = (layer5_outputs[786]) & (layer5_outputs[1387]);
    assign layer6_outputs[2822] = (layer5_outputs[2977]) | (layer5_outputs[1072]);
    assign layer6_outputs[2823] = 1'b1;
    assign layer6_outputs[2824] = ~(layer5_outputs[2360]);
    assign layer6_outputs[2825] = ~((layer5_outputs[3693]) | (layer5_outputs[2624]));
    assign layer6_outputs[2826] = layer5_outputs[4611];
    assign layer6_outputs[2827] = ~(layer5_outputs[3514]);
    assign layer6_outputs[2828] = (layer5_outputs[2186]) ^ (layer5_outputs[3807]);
    assign layer6_outputs[2829] = (layer5_outputs[1044]) | (layer5_outputs[4776]);
    assign layer6_outputs[2830] = layer5_outputs[4002];
    assign layer6_outputs[2831] = ~((layer5_outputs[1115]) | (layer5_outputs[3100]));
    assign layer6_outputs[2832] = (layer5_outputs[1237]) & (layer5_outputs[824]);
    assign layer6_outputs[2833] = (layer5_outputs[3883]) | (layer5_outputs[4771]);
    assign layer6_outputs[2834] = (layer5_outputs[4332]) ^ (layer5_outputs[4057]);
    assign layer6_outputs[2835] = ~(layer5_outputs[5046]);
    assign layer6_outputs[2836] = ~(layer5_outputs[4383]);
    assign layer6_outputs[2837] = (layer5_outputs[441]) & (layer5_outputs[357]);
    assign layer6_outputs[2838] = 1'b0;
    assign layer6_outputs[2839] = ~(layer5_outputs[4261]);
    assign layer6_outputs[2840] = ~((layer5_outputs[1517]) ^ (layer5_outputs[2918]));
    assign layer6_outputs[2841] = ~(layer5_outputs[2454]);
    assign layer6_outputs[2842] = ~((layer5_outputs[2411]) | (layer5_outputs[478]));
    assign layer6_outputs[2843] = ~(layer5_outputs[2127]);
    assign layer6_outputs[2844] = layer5_outputs[3185];
    assign layer6_outputs[2845] = layer5_outputs[1706];
    assign layer6_outputs[2846] = layer5_outputs[2704];
    assign layer6_outputs[2847] = 1'b0;
    assign layer6_outputs[2848] = ~((layer5_outputs[763]) ^ (layer5_outputs[16]));
    assign layer6_outputs[2849] = (layer5_outputs[922]) & ~(layer5_outputs[3235]);
    assign layer6_outputs[2850] = ~(layer5_outputs[1639]) | (layer5_outputs[2212]);
    assign layer6_outputs[2851] = layer5_outputs[4207];
    assign layer6_outputs[2852] = ~(layer5_outputs[2652]);
    assign layer6_outputs[2853] = ~((layer5_outputs[981]) ^ (layer5_outputs[1426]));
    assign layer6_outputs[2854] = ~(layer5_outputs[1755]) | (layer5_outputs[1360]);
    assign layer6_outputs[2855] = layer5_outputs[1300];
    assign layer6_outputs[2856] = (layer5_outputs[2171]) ^ (layer5_outputs[4521]);
    assign layer6_outputs[2857] = (layer5_outputs[1247]) & ~(layer5_outputs[3305]);
    assign layer6_outputs[2858] = layer5_outputs[4971];
    assign layer6_outputs[2859] = (layer5_outputs[3343]) ^ (layer5_outputs[3374]);
    assign layer6_outputs[2860] = layer5_outputs[3231];
    assign layer6_outputs[2861] = layer5_outputs[4826];
    assign layer6_outputs[2862] = ~((layer5_outputs[4196]) ^ (layer5_outputs[2101]));
    assign layer6_outputs[2863] = ~(layer5_outputs[3360]);
    assign layer6_outputs[2864] = ~(layer5_outputs[4718]);
    assign layer6_outputs[2865] = ~(layer5_outputs[5034]);
    assign layer6_outputs[2866] = ~(layer5_outputs[3786]);
    assign layer6_outputs[2867] = ~(layer5_outputs[4667]) | (layer5_outputs[1543]);
    assign layer6_outputs[2868] = layer5_outputs[4999];
    assign layer6_outputs[2869] = (layer5_outputs[2566]) ^ (layer5_outputs[3826]);
    assign layer6_outputs[2870] = layer5_outputs[4433];
    assign layer6_outputs[2871] = (layer5_outputs[4852]) & (layer5_outputs[3781]);
    assign layer6_outputs[2872] = layer5_outputs[4382];
    assign layer6_outputs[2873] = (layer5_outputs[2207]) & (layer5_outputs[2098]);
    assign layer6_outputs[2874] = layer5_outputs[22];
    assign layer6_outputs[2875] = layer5_outputs[3619];
    assign layer6_outputs[2876] = ~(layer5_outputs[2013]) | (layer5_outputs[1438]);
    assign layer6_outputs[2877] = layer5_outputs[2152];
    assign layer6_outputs[2878] = ~(layer5_outputs[3595]);
    assign layer6_outputs[2879] = (layer5_outputs[3115]) | (layer5_outputs[1263]);
    assign layer6_outputs[2880] = ~(layer5_outputs[2321]);
    assign layer6_outputs[2881] = (layer5_outputs[3845]) & ~(layer5_outputs[2063]);
    assign layer6_outputs[2882] = ~(layer5_outputs[1965]);
    assign layer6_outputs[2883] = ~(layer5_outputs[4699]) | (layer5_outputs[2423]);
    assign layer6_outputs[2884] = layer5_outputs[1444];
    assign layer6_outputs[2885] = (layer5_outputs[1687]) | (layer5_outputs[3327]);
    assign layer6_outputs[2886] = ~(layer5_outputs[540]);
    assign layer6_outputs[2887] = ~(layer5_outputs[3636]);
    assign layer6_outputs[2888] = layer5_outputs[3527];
    assign layer6_outputs[2889] = (layer5_outputs[4338]) & ~(layer5_outputs[951]);
    assign layer6_outputs[2890] = layer5_outputs[1650];
    assign layer6_outputs[2891] = ~(layer5_outputs[2715]);
    assign layer6_outputs[2892] = ~((layer5_outputs[149]) | (layer5_outputs[3892]));
    assign layer6_outputs[2893] = ~((layer5_outputs[1004]) & (layer5_outputs[904]));
    assign layer6_outputs[2894] = (layer5_outputs[170]) & ~(layer5_outputs[2641]);
    assign layer6_outputs[2895] = layer5_outputs[306];
    assign layer6_outputs[2896] = ~(layer5_outputs[2075]);
    assign layer6_outputs[2897] = (layer5_outputs[4335]) & ~(layer5_outputs[3476]);
    assign layer6_outputs[2898] = ~(layer5_outputs[4793]);
    assign layer6_outputs[2899] = ~(layer5_outputs[5019]) | (layer5_outputs[5076]);
    assign layer6_outputs[2900] = ~(layer5_outputs[1286]);
    assign layer6_outputs[2901] = layer5_outputs[4153];
    assign layer6_outputs[2902] = (layer5_outputs[4388]) & (layer5_outputs[1193]);
    assign layer6_outputs[2903] = ~((layer5_outputs[844]) & (layer5_outputs[4686]));
    assign layer6_outputs[2904] = ~(layer5_outputs[126]);
    assign layer6_outputs[2905] = ~(layer5_outputs[3792]);
    assign layer6_outputs[2906] = ~((layer5_outputs[1442]) ^ (layer5_outputs[4645]));
    assign layer6_outputs[2907] = ~((layer5_outputs[712]) & (layer5_outputs[1942]));
    assign layer6_outputs[2908] = layer5_outputs[1307];
    assign layer6_outputs[2909] = ~(layer5_outputs[1073]);
    assign layer6_outputs[2910] = ~((layer5_outputs[4991]) & (layer5_outputs[4761]));
    assign layer6_outputs[2911] = ~(layer5_outputs[1221]) | (layer5_outputs[626]);
    assign layer6_outputs[2912] = layer5_outputs[3012];
    assign layer6_outputs[2913] = layer5_outputs[2865];
    assign layer6_outputs[2914] = layer5_outputs[1209];
    assign layer6_outputs[2915] = layer5_outputs[4420];
    assign layer6_outputs[2916] = layer5_outputs[2244];
    assign layer6_outputs[2917] = ~(layer5_outputs[3442]);
    assign layer6_outputs[2918] = (layer5_outputs[1776]) ^ (layer5_outputs[2860]);
    assign layer6_outputs[2919] = ~((layer5_outputs[2571]) | (layer5_outputs[696]));
    assign layer6_outputs[2920] = layer5_outputs[5114];
    assign layer6_outputs[2921] = ~((layer5_outputs[186]) ^ (layer5_outputs[1007]));
    assign layer6_outputs[2922] = layer5_outputs[4301];
    assign layer6_outputs[2923] = (layer5_outputs[2162]) & (layer5_outputs[2495]);
    assign layer6_outputs[2924] = ~(layer5_outputs[1149]);
    assign layer6_outputs[2925] = ~((layer5_outputs[4786]) ^ (layer5_outputs[2456]));
    assign layer6_outputs[2926] = layer5_outputs[52];
    assign layer6_outputs[2927] = ~(layer5_outputs[3938]);
    assign layer6_outputs[2928] = ~(layer5_outputs[2271]);
    assign layer6_outputs[2929] = layer5_outputs[4856];
    assign layer6_outputs[2930] = ~(layer5_outputs[1881]);
    assign layer6_outputs[2931] = ~(layer5_outputs[3060]);
    assign layer6_outputs[2932] = layer5_outputs[3393];
    assign layer6_outputs[2933] = layer5_outputs[959];
    assign layer6_outputs[2934] = ~(layer5_outputs[4868]);
    assign layer6_outputs[2935] = layer5_outputs[3074];
    assign layer6_outputs[2936] = (layer5_outputs[2274]) & ~(layer5_outputs[3840]);
    assign layer6_outputs[2937] = ~(layer5_outputs[2674]);
    assign layer6_outputs[2938] = layer5_outputs[957];
    assign layer6_outputs[2939] = (layer5_outputs[1985]) & ~(layer5_outputs[2422]);
    assign layer6_outputs[2940] = (layer5_outputs[1617]) & (layer5_outputs[639]);
    assign layer6_outputs[2941] = ~((layer5_outputs[1250]) ^ (layer5_outputs[428]));
    assign layer6_outputs[2942] = layer5_outputs[2080];
    assign layer6_outputs[2943] = ~(layer5_outputs[287]);
    assign layer6_outputs[2944] = ~(layer5_outputs[3214]) | (layer5_outputs[1799]);
    assign layer6_outputs[2945] = ~(layer5_outputs[2897]) | (layer5_outputs[4883]);
    assign layer6_outputs[2946] = (layer5_outputs[3384]) ^ (layer5_outputs[920]);
    assign layer6_outputs[2947] = ~(layer5_outputs[269]);
    assign layer6_outputs[2948] = layer5_outputs[4385];
    assign layer6_outputs[2949] = ~((layer5_outputs[951]) | (layer5_outputs[4527]));
    assign layer6_outputs[2950] = (layer5_outputs[724]) ^ (layer5_outputs[3846]);
    assign layer6_outputs[2951] = ~(layer5_outputs[624]);
    assign layer6_outputs[2952] = ~(layer5_outputs[1276]) | (layer5_outputs[4348]);
    assign layer6_outputs[2953] = ~(layer5_outputs[2305]);
    assign layer6_outputs[2954] = ~((layer5_outputs[3920]) & (layer5_outputs[3011]));
    assign layer6_outputs[2955] = ~((layer5_outputs[483]) ^ (layer5_outputs[4206]));
    assign layer6_outputs[2956] = (layer5_outputs[2014]) & (layer5_outputs[902]);
    assign layer6_outputs[2957] = ~(layer5_outputs[4663]);
    assign layer6_outputs[2958] = (layer5_outputs[3274]) & ~(layer5_outputs[4857]);
    assign layer6_outputs[2959] = ~(layer5_outputs[3157]);
    assign layer6_outputs[2960] = (layer5_outputs[1144]) ^ (layer5_outputs[3308]);
    assign layer6_outputs[2961] = layer5_outputs[1779];
    assign layer6_outputs[2962] = ~((layer5_outputs[646]) ^ (layer5_outputs[4899]));
    assign layer6_outputs[2963] = ~(layer5_outputs[1285]);
    assign layer6_outputs[2964] = layer5_outputs[1832];
    assign layer6_outputs[2965] = (layer5_outputs[2112]) ^ (layer5_outputs[4601]);
    assign layer6_outputs[2966] = ~((layer5_outputs[1368]) ^ (layer5_outputs[710]));
    assign layer6_outputs[2967] = ~(layer5_outputs[180]);
    assign layer6_outputs[2968] = ~(layer5_outputs[701]);
    assign layer6_outputs[2969] = ~(layer5_outputs[2458]);
    assign layer6_outputs[2970] = ~(layer5_outputs[4689]);
    assign layer6_outputs[2971] = layer5_outputs[3998];
    assign layer6_outputs[2972] = ~(layer5_outputs[4158]);
    assign layer6_outputs[2973] = ~(layer5_outputs[3431]);
    assign layer6_outputs[2974] = layer5_outputs[737];
    assign layer6_outputs[2975] = ~(layer5_outputs[3275]);
    assign layer6_outputs[2976] = layer5_outputs[822];
    assign layer6_outputs[2977] = ~(layer5_outputs[4925]);
    assign layer6_outputs[2978] = ~(layer5_outputs[3716]);
    assign layer6_outputs[2979] = (layer5_outputs[3032]) | (layer5_outputs[4166]);
    assign layer6_outputs[2980] = layer5_outputs[2638];
    assign layer6_outputs[2981] = ~(layer5_outputs[1916]);
    assign layer6_outputs[2982] = (layer5_outputs[4820]) ^ (layer5_outputs[4543]);
    assign layer6_outputs[2983] = layer5_outputs[2076];
    assign layer6_outputs[2984] = layer5_outputs[2620];
    assign layer6_outputs[2985] = layer5_outputs[4760];
    assign layer6_outputs[2986] = layer5_outputs[3746];
    assign layer6_outputs[2987] = (layer5_outputs[2990]) & ~(layer5_outputs[2052]);
    assign layer6_outputs[2988] = ~(layer5_outputs[4654]);
    assign layer6_outputs[2989] = (layer5_outputs[2241]) ^ (layer5_outputs[4067]);
    assign layer6_outputs[2990] = layer5_outputs[1685];
    assign layer6_outputs[2991] = ~((layer5_outputs[4148]) ^ (layer5_outputs[372]));
    assign layer6_outputs[2992] = ~(layer5_outputs[1410]);
    assign layer6_outputs[2993] = (layer5_outputs[175]) | (layer5_outputs[663]);
    assign layer6_outputs[2994] = (layer5_outputs[1777]) ^ (layer5_outputs[2384]);
    assign layer6_outputs[2995] = layer5_outputs[4760];
    assign layer6_outputs[2996] = ~(layer5_outputs[1589]) | (layer5_outputs[2059]);
    assign layer6_outputs[2997] = ~(layer5_outputs[2454]);
    assign layer6_outputs[2998] = layer5_outputs[1871];
    assign layer6_outputs[2999] = (layer5_outputs[1020]) & ~(layer5_outputs[4425]);
    assign layer6_outputs[3000] = layer5_outputs[2832];
    assign layer6_outputs[3001] = (layer5_outputs[3212]) & ~(layer5_outputs[3254]);
    assign layer6_outputs[3002] = (layer5_outputs[2790]) & (layer5_outputs[2757]);
    assign layer6_outputs[3003] = ~((layer5_outputs[4449]) ^ (layer5_outputs[3349]));
    assign layer6_outputs[3004] = layer5_outputs[4775];
    assign layer6_outputs[3005] = ~(layer5_outputs[3698]);
    assign layer6_outputs[3006] = ~(layer5_outputs[3562]) | (layer5_outputs[5078]);
    assign layer6_outputs[3007] = ~((layer5_outputs[2249]) & (layer5_outputs[2822]));
    assign layer6_outputs[3008] = ~(layer5_outputs[984]);
    assign layer6_outputs[3009] = (layer5_outputs[925]) ^ (layer5_outputs[5075]);
    assign layer6_outputs[3010] = ~(layer5_outputs[3694]);
    assign layer6_outputs[3011] = ~(layer5_outputs[1163]);
    assign layer6_outputs[3012] = ~((layer5_outputs[3968]) | (layer5_outputs[1465]));
    assign layer6_outputs[3013] = (layer5_outputs[3442]) ^ (layer5_outputs[1355]);
    assign layer6_outputs[3014] = ~(layer5_outputs[3379]);
    assign layer6_outputs[3015] = layer5_outputs[3302];
    assign layer6_outputs[3016] = (layer5_outputs[3164]) & ~(layer5_outputs[4859]);
    assign layer6_outputs[3017] = (layer5_outputs[16]) & ~(layer5_outputs[2107]);
    assign layer6_outputs[3018] = ~((layer5_outputs[3299]) ^ (layer5_outputs[1409]));
    assign layer6_outputs[3019] = layer5_outputs[3147];
    assign layer6_outputs[3020] = ~(layer5_outputs[5062]);
    assign layer6_outputs[3021] = ~(layer5_outputs[1586]);
    assign layer6_outputs[3022] = ~(layer5_outputs[3865]) | (layer5_outputs[3500]);
    assign layer6_outputs[3023] = layer5_outputs[1081];
    assign layer6_outputs[3024] = ~((layer5_outputs[1385]) | (layer5_outputs[3314]));
    assign layer6_outputs[3025] = layer5_outputs[1128];
    assign layer6_outputs[3026] = ~(layer5_outputs[4231]);
    assign layer6_outputs[3027] = (layer5_outputs[4537]) & (layer5_outputs[218]);
    assign layer6_outputs[3028] = layer5_outputs[241];
    assign layer6_outputs[3029] = ~(layer5_outputs[761]);
    assign layer6_outputs[3030] = layer5_outputs[5078];
    assign layer6_outputs[3031] = (layer5_outputs[4802]) & ~(layer5_outputs[1537]);
    assign layer6_outputs[3032] = (layer5_outputs[607]) & ~(layer5_outputs[3414]);
    assign layer6_outputs[3033] = ~(layer5_outputs[5059]);
    assign layer6_outputs[3034] = ~(layer5_outputs[4913]) | (layer5_outputs[3828]);
    assign layer6_outputs[3035] = (layer5_outputs[1223]) & ~(layer5_outputs[3385]);
    assign layer6_outputs[3036] = ~((layer5_outputs[3654]) & (layer5_outputs[3718]));
    assign layer6_outputs[3037] = ~(layer5_outputs[1079]);
    assign layer6_outputs[3038] = layer5_outputs[557];
    assign layer6_outputs[3039] = ~(layer5_outputs[2081]);
    assign layer6_outputs[3040] = layer5_outputs[282];
    assign layer6_outputs[3041] = layer5_outputs[1348];
    assign layer6_outputs[3042] = layer5_outputs[424];
    assign layer6_outputs[3043] = ~(layer5_outputs[2778]);
    assign layer6_outputs[3044] = layer5_outputs[3302];
    assign layer6_outputs[3045] = (layer5_outputs[3747]) ^ (layer5_outputs[2697]);
    assign layer6_outputs[3046] = (layer5_outputs[4186]) & ~(layer5_outputs[4633]);
    assign layer6_outputs[3047] = layer5_outputs[4802];
    assign layer6_outputs[3048] = ~(layer5_outputs[873]);
    assign layer6_outputs[3049] = layer5_outputs[1307];
    assign layer6_outputs[3050] = ~((layer5_outputs[2587]) & (layer5_outputs[415]));
    assign layer6_outputs[3051] = ~(layer5_outputs[4571]);
    assign layer6_outputs[3052] = ~((layer5_outputs[4958]) ^ (layer5_outputs[3928]));
    assign layer6_outputs[3053] = layer5_outputs[3298];
    assign layer6_outputs[3054] = (layer5_outputs[1138]) | (layer5_outputs[2138]);
    assign layer6_outputs[3055] = ~(layer5_outputs[5018]);
    assign layer6_outputs[3056] = ~(layer5_outputs[787]);
    assign layer6_outputs[3057] = layer5_outputs[3150];
    assign layer6_outputs[3058] = layer5_outputs[1766];
    assign layer6_outputs[3059] = ~(layer5_outputs[4301]);
    assign layer6_outputs[3060] = ~((layer5_outputs[2372]) | (layer5_outputs[4344]));
    assign layer6_outputs[3061] = ~(layer5_outputs[195]);
    assign layer6_outputs[3062] = (layer5_outputs[3916]) ^ (layer5_outputs[4672]);
    assign layer6_outputs[3063] = ~(layer5_outputs[4790]);
    assign layer6_outputs[3064] = ~((layer5_outputs[601]) ^ (layer5_outputs[1191]));
    assign layer6_outputs[3065] = ~(layer5_outputs[1294]);
    assign layer6_outputs[3066] = ~((layer5_outputs[4089]) ^ (layer5_outputs[3163]));
    assign layer6_outputs[3067] = ~(layer5_outputs[4967]);
    assign layer6_outputs[3068] = ~(layer5_outputs[4378]);
    assign layer6_outputs[3069] = layer5_outputs[1490];
    assign layer6_outputs[3070] = ~((layer5_outputs[325]) ^ (layer5_outputs[3749]));
    assign layer6_outputs[3071] = 1'b1;
    assign layer6_outputs[3072] = ~((layer5_outputs[3450]) | (layer5_outputs[4138]));
    assign layer6_outputs[3073] = ~(layer5_outputs[3907]);
    assign layer6_outputs[3074] = ~(layer5_outputs[1122]) | (layer5_outputs[1264]);
    assign layer6_outputs[3075] = ~(layer5_outputs[842]);
    assign layer6_outputs[3076] = ~(layer5_outputs[3871]);
    assign layer6_outputs[3077] = layer5_outputs[2390];
    assign layer6_outputs[3078] = (layer5_outputs[1956]) & ~(layer5_outputs[2911]);
    assign layer6_outputs[3079] = ~(layer5_outputs[2788]);
    assign layer6_outputs[3080] = ~((layer5_outputs[2954]) | (layer5_outputs[2409]));
    assign layer6_outputs[3081] = ~(layer5_outputs[1084]);
    assign layer6_outputs[3082] = layer5_outputs[3412];
    assign layer6_outputs[3083] = ~(layer5_outputs[3389]);
    assign layer6_outputs[3084] = 1'b1;
    assign layer6_outputs[3085] = (layer5_outputs[3830]) ^ (layer5_outputs[741]);
    assign layer6_outputs[3086] = (layer5_outputs[316]) ^ (layer5_outputs[2665]);
    assign layer6_outputs[3087] = layer5_outputs[2467];
    assign layer6_outputs[3088] = layer5_outputs[2304];
    assign layer6_outputs[3089] = layer5_outputs[3078];
    assign layer6_outputs[3090] = ~(layer5_outputs[2310]);
    assign layer6_outputs[3091] = (layer5_outputs[3942]) ^ (layer5_outputs[2677]);
    assign layer6_outputs[3092] = (layer5_outputs[488]) ^ (layer5_outputs[3328]);
    assign layer6_outputs[3093] = ~((layer5_outputs[4733]) ^ (layer5_outputs[804]));
    assign layer6_outputs[3094] = ~(layer5_outputs[911]);
    assign layer6_outputs[3095] = (layer5_outputs[1993]) ^ (layer5_outputs[838]);
    assign layer6_outputs[3096] = layer5_outputs[231];
    assign layer6_outputs[3097] = ~((layer5_outputs[2112]) | (layer5_outputs[2965]));
    assign layer6_outputs[3098] = ~(layer5_outputs[4438]);
    assign layer6_outputs[3099] = layer5_outputs[1348];
    assign layer6_outputs[3100] = layer5_outputs[4271];
    assign layer6_outputs[3101] = (layer5_outputs[3373]) & ~(layer5_outputs[367]);
    assign layer6_outputs[3102] = ~(layer5_outputs[2066]) | (layer5_outputs[1734]);
    assign layer6_outputs[3103] = ~(layer5_outputs[4359]);
    assign layer6_outputs[3104] = 1'b0;
    assign layer6_outputs[3105] = layer5_outputs[2859];
    assign layer6_outputs[3106] = (layer5_outputs[2285]) ^ (layer5_outputs[1714]);
    assign layer6_outputs[3107] = (layer5_outputs[2911]) | (layer5_outputs[126]);
    assign layer6_outputs[3108] = layer5_outputs[3130];
    assign layer6_outputs[3109] = layer5_outputs[4682];
    assign layer6_outputs[3110] = ~((layer5_outputs[383]) & (layer5_outputs[410]));
    assign layer6_outputs[3111] = 1'b0;
    assign layer6_outputs[3112] = layer5_outputs[4849];
    assign layer6_outputs[3113] = ~(layer5_outputs[3250]);
    assign layer6_outputs[3114] = 1'b0;
    assign layer6_outputs[3115] = ~((layer5_outputs[341]) ^ (layer5_outputs[1813]));
    assign layer6_outputs[3116] = layer5_outputs[2123];
    assign layer6_outputs[3117] = ~(layer5_outputs[1527]) | (layer5_outputs[4500]);
    assign layer6_outputs[3118] = ~((layer5_outputs[816]) | (layer5_outputs[2367]));
    assign layer6_outputs[3119] = layer5_outputs[3600];
    assign layer6_outputs[3120] = layer5_outputs[2900];
    assign layer6_outputs[3121] = ~((layer5_outputs[3867]) | (layer5_outputs[2034]));
    assign layer6_outputs[3122] = ~(layer5_outputs[2832]) | (layer5_outputs[2623]);
    assign layer6_outputs[3123] = layer5_outputs[99];
    assign layer6_outputs[3124] = ~(layer5_outputs[1924]);
    assign layer6_outputs[3125] = ~(layer5_outputs[1544]) | (layer5_outputs[3251]);
    assign layer6_outputs[3126] = ~(layer5_outputs[81]);
    assign layer6_outputs[3127] = ~(layer5_outputs[3433]);
    assign layer6_outputs[3128] = ~(layer5_outputs[772]);
    assign layer6_outputs[3129] = (layer5_outputs[1085]) ^ (layer5_outputs[2593]);
    assign layer6_outputs[3130] = ~(layer5_outputs[1578]);
    assign layer6_outputs[3131] = ~((layer5_outputs[2760]) & (layer5_outputs[4241]));
    assign layer6_outputs[3132] = (layer5_outputs[3891]) ^ (layer5_outputs[4846]);
    assign layer6_outputs[3133] = (layer5_outputs[4452]) ^ (layer5_outputs[1199]);
    assign layer6_outputs[3134] = layer5_outputs[792];
    assign layer6_outputs[3135] = (layer5_outputs[648]) & ~(layer5_outputs[4290]);
    assign layer6_outputs[3136] = ~(layer5_outputs[1197]);
    assign layer6_outputs[3137] = ~((layer5_outputs[719]) & (layer5_outputs[1159]));
    assign layer6_outputs[3138] = ~(layer5_outputs[4081]);
    assign layer6_outputs[3139] = (layer5_outputs[3524]) & ~(layer5_outputs[1923]);
    assign layer6_outputs[3140] = (layer5_outputs[2549]) & (layer5_outputs[4935]);
    assign layer6_outputs[3141] = ~(layer5_outputs[960]) | (layer5_outputs[4459]);
    assign layer6_outputs[3142] = ~((layer5_outputs[2382]) | (layer5_outputs[2288]));
    assign layer6_outputs[3143] = ~(layer5_outputs[1481]);
    assign layer6_outputs[3144] = (layer5_outputs[4747]) ^ (layer5_outputs[4018]);
    assign layer6_outputs[3145] = ~(layer5_outputs[45]);
    assign layer6_outputs[3146] = ~((layer5_outputs[3410]) ^ (layer5_outputs[2820]));
    assign layer6_outputs[3147] = (layer5_outputs[2631]) ^ (layer5_outputs[613]);
    assign layer6_outputs[3148] = (layer5_outputs[2987]) & ~(layer5_outputs[3179]);
    assign layer6_outputs[3149] = (layer5_outputs[3675]) & (layer5_outputs[521]);
    assign layer6_outputs[3150] = (layer5_outputs[2008]) & ~(layer5_outputs[447]);
    assign layer6_outputs[3151] = (layer5_outputs[681]) & ~(layer5_outputs[1920]);
    assign layer6_outputs[3152] = ~(layer5_outputs[2347]) | (layer5_outputs[2981]);
    assign layer6_outputs[3153] = layer5_outputs[3987];
    assign layer6_outputs[3154] = ~((layer5_outputs[1222]) | (layer5_outputs[4731]));
    assign layer6_outputs[3155] = ~(layer5_outputs[1148]);
    assign layer6_outputs[3156] = (layer5_outputs[3513]) ^ (layer5_outputs[4277]);
    assign layer6_outputs[3157] = ~((layer5_outputs[23]) ^ (layer5_outputs[3977]));
    assign layer6_outputs[3158] = layer5_outputs[3613];
    assign layer6_outputs[3159] = ~(layer5_outputs[692]);
    assign layer6_outputs[3160] = ~(layer5_outputs[368]);
    assign layer6_outputs[3161] = ~(layer5_outputs[4780]);
    assign layer6_outputs[3162] = ~(layer5_outputs[518]) | (layer5_outputs[962]);
    assign layer6_outputs[3163] = layer5_outputs[3132];
    assign layer6_outputs[3164] = 1'b0;
    assign layer6_outputs[3165] = layer5_outputs[3363];
    assign layer6_outputs[3166] = layer5_outputs[1005];
    assign layer6_outputs[3167] = layer5_outputs[493];
    assign layer6_outputs[3168] = layer5_outputs[4476];
    assign layer6_outputs[3169] = (layer5_outputs[1486]) ^ (layer5_outputs[3590]);
    assign layer6_outputs[3170] = layer5_outputs[4976];
    assign layer6_outputs[3171] = (layer5_outputs[3505]) | (layer5_outputs[1255]);
    assign layer6_outputs[3172] = layer5_outputs[2564];
    assign layer6_outputs[3173] = (layer5_outputs[4977]) & ~(layer5_outputs[260]);
    assign layer6_outputs[3174] = (layer5_outputs[4304]) & ~(layer5_outputs[391]);
    assign layer6_outputs[3175] = ~(layer5_outputs[1178]);
    assign layer6_outputs[3176] = ~((layer5_outputs[4783]) | (layer5_outputs[1938]));
    assign layer6_outputs[3177] = ~(layer5_outputs[4615]);
    assign layer6_outputs[3178] = ~(layer5_outputs[2513]);
    assign layer6_outputs[3179] = ~(layer5_outputs[1465]) | (layer5_outputs[381]);
    assign layer6_outputs[3180] = layer5_outputs[1419];
    assign layer6_outputs[3181] = ~(layer5_outputs[3173]);
    assign layer6_outputs[3182] = ~(layer5_outputs[3775]) | (layer5_outputs[4939]);
    assign layer6_outputs[3183] = layer5_outputs[2913];
    assign layer6_outputs[3184] = (layer5_outputs[1391]) & ~(layer5_outputs[1858]);
    assign layer6_outputs[3185] = ~((layer5_outputs[4542]) ^ (layer5_outputs[3593]));
    assign layer6_outputs[3186] = layer5_outputs[1411];
    assign layer6_outputs[3187] = layer5_outputs[489];
    assign layer6_outputs[3188] = (layer5_outputs[1841]) & ~(layer5_outputs[4728]);
    assign layer6_outputs[3189] = ~(layer5_outputs[2871]) | (layer5_outputs[4562]);
    assign layer6_outputs[3190] = layer5_outputs[2664];
    assign layer6_outputs[3191] = layer5_outputs[1527];
    assign layer6_outputs[3192] = ~(layer5_outputs[1605]);
    assign layer6_outputs[3193] = (layer5_outputs[1402]) & ~(layer5_outputs[4012]);
    assign layer6_outputs[3194] = (layer5_outputs[521]) & ~(layer5_outputs[431]);
    assign layer6_outputs[3195] = (layer5_outputs[1503]) & ~(layer5_outputs[2990]);
    assign layer6_outputs[3196] = ~(layer5_outputs[1862]);
    assign layer6_outputs[3197] = ~((layer5_outputs[576]) | (layer5_outputs[1131]));
    assign layer6_outputs[3198] = (layer5_outputs[2964]) | (layer5_outputs[314]);
    assign layer6_outputs[3199] = layer5_outputs[380];
    assign layer6_outputs[3200] = layer5_outputs[3345];
    assign layer6_outputs[3201] = (layer5_outputs[932]) & ~(layer5_outputs[4121]);
    assign layer6_outputs[3202] = layer5_outputs[2127];
    assign layer6_outputs[3203] = layer5_outputs[1397];
    assign layer6_outputs[3204] = (layer5_outputs[2763]) ^ (layer5_outputs[2564]);
    assign layer6_outputs[3205] = ~(layer5_outputs[927]) | (layer5_outputs[891]);
    assign layer6_outputs[3206] = layer5_outputs[3805];
    assign layer6_outputs[3207] = (layer5_outputs[154]) & ~(layer5_outputs[3161]);
    assign layer6_outputs[3208] = ~((layer5_outputs[2387]) ^ (layer5_outputs[3131]));
    assign layer6_outputs[3209] = ~((layer5_outputs[1686]) | (layer5_outputs[3560]));
    assign layer6_outputs[3210] = (layer5_outputs[1100]) ^ (layer5_outputs[2055]);
    assign layer6_outputs[3211] = (layer5_outputs[2024]) & ~(layer5_outputs[1030]);
    assign layer6_outputs[3212] = ~(layer5_outputs[2913]) | (layer5_outputs[3587]);
    assign layer6_outputs[3213] = ~(layer5_outputs[3306]);
    assign layer6_outputs[3214] = (layer5_outputs[4968]) & ~(layer5_outputs[393]);
    assign layer6_outputs[3215] = layer5_outputs[1702];
    assign layer6_outputs[3216] = (layer5_outputs[633]) ^ (layer5_outputs[4990]);
    assign layer6_outputs[3217] = ~(layer5_outputs[1563]);
    assign layer6_outputs[3218] = layer5_outputs[822];
    assign layer6_outputs[3219] = layer5_outputs[3792];
    assign layer6_outputs[3220] = (layer5_outputs[1897]) ^ (layer5_outputs[2825]);
    assign layer6_outputs[3221] = layer5_outputs[1985];
    assign layer6_outputs[3222] = ~(layer5_outputs[3321]) | (layer5_outputs[1741]);
    assign layer6_outputs[3223] = ~((layer5_outputs[4409]) & (layer5_outputs[2734]));
    assign layer6_outputs[3224] = layer5_outputs[3656];
    assign layer6_outputs[3225] = ~(layer5_outputs[1612]) | (layer5_outputs[2188]);
    assign layer6_outputs[3226] = ~(layer5_outputs[1124]);
    assign layer6_outputs[3227] = layer5_outputs[3433];
    assign layer6_outputs[3228] = ~(layer5_outputs[881]);
    assign layer6_outputs[3229] = ~((layer5_outputs[2031]) | (layer5_outputs[2242]));
    assign layer6_outputs[3230] = layer5_outputs[3286];
    assign layer6_outputs[3231] = layer5_outputs[2451];
    assign layer6_outputs[3232] = (layer5_outputs[2486]) ^ (layer5_outputs[446]);
    assign layer6_outputs[3233] = ~(layer5_outputs[1052]) | (layer5_outputs[1702]);
    assign layer6_outputs[3234] = layer5_outputs[1056];
    assign layer6_outputs[3235] = layer5_outputs[1909];
    assign layer6_outputs[3236] = (layer5_outputs[4834]) | (layer5_outputs[3507]);
    assign layer6_outputs[3237] = ~(layer5_outputs[4739]) | (layer5_outputs[3869]);
    assign layer6_outputs[3238] = layer5_outputs[4885];
    assign layer6_outputs[3239] = ~(layer5_outputs[194]);
    assign layer6_outputs[3240] = ~(layer5_outputs[2239]);
    assign layer6_outputs[3241] = layer5_outputs[2801];
    assign layer6_outputs[3242] = ~(layer5_outputs[1109]);
    assign layer6_outputs[3243] = ~(layer5_outputs[1889]);
    assign layer6_outputs[3244] = ~(layer5_outputs[989]);
    assign layer6_outputs[3245] = ~(layer5_outputs[4772]);
    assign layer6_outputs[3246] = ~(layer5_outputs[2460]);
    assign layer6_outputs[3247] = ~(layer5_outputs[451]);
    assign layer6_outputs[3248] = layer5_outputs[1215];
    assign layer6_outputs[3249] = ~(layer5_outputs[295]);
    assign layer6_outputs[3250] = layer5_outputs[1830];
    assign layer6_outputs[3251] = ~(layer5_outputs[1182]);
    assign layer6_outputs[3252] = ~(layer5_outputs[1757]);
    assign layer6_outputs[3253] = layer5_outputs[5029];
    assign layer6_outputs[3254] = ~(layer5_outputs[3066]);
    assign layer6_outputs[3255] = layer5_outputs[1023];
    assign layer6_outputs[3256] = ~(layer5_outputs[3332]) | (layer5_outputs[2291]);
    assign layer6_outputs[3257] = ~(layer5_outputs[4680]) | (layer5_outputs[4446]);
    assign layer6_outputs[3258] = ~(layer5_outputs[2286]) | (layer5_outputs[518]);
    assign layer6_outputs[3259] = layer5_outputs[4916];
    assign layer6_outputs[3260] = (layer5_outputs[4346]) & (layer5_outputs[1493]);
    assign layer6_outputs[3261] = ~(layer5_outputs[929]) | (layer5_outputs[1844]);
    assign layer6_outputs[3262] = ~(layer5_outputs[4191]);
    assign layer6_outputs[3263] = ~((layer5_outputs[785]) ^ (layer5_outputs[1141]));
    assign layer6_outputs[3264] = ~(layer5_outputs[3854]);
    assign layer6_outputs[3265] = layer5_outputs[538];
    assign layer6_outputs[3266] = layer5_outputs[771];
    assign layer6_outputs[3267] = ~(layer5_outputs[2230]);
    assign layer6_outputs[3268] = layer5_outputs[3919];
    assign layer6_outputs[3269] = (layer5_outputs[4700]) & ~(layer5_outputs[3992]);
    assign layer6_outputs[3270] = ~(layer5_outputs[2301]) | (layer5_outputs[4769]);
    assign layer6_outputs[3271] = ~((layer5_outputs[726]) & (layer5_outputs[2433]));
    assign layer6_outputs[3272] = ~((layer5_outputs[1265]) | (layer5_outputs[346]));
    assign layer6_outputs[3273] = layer5_outputs[2812];
    assign layer6_outputs[3274] = layer5_outputs[1105];
    assign layer6_outputs[3275] = ~((layer5_outputs[4861]) ^ (layer5_outputs[3659]));
    assign layer6_outputs[3276] = (layer5_outputs[1585]) ^ (layer5_outputs[1676]);
    assign layer6_outputs[3277] = layer5_outputs[4853];
    assign layer6_outputs[3278] = (layer5_outputs[4082]) ^ (layer5_outputs[2663]);
    assign layer6_outputs[3279] = (layer5_outputs[57]) ^ (layer5_outputs[4754]);
    assign layer6_outputs[3280] = layer5_outputs[972];
    assign layer6_outputs[3281] = (layer5_outputs[5115]) & (layer5_outputs[1406]);
    assign layer6_outputs[3282] = ~(layer5_outputs[3242]);
    assign layer6_outputs[3283] = ~(layer5_outputs[1451]);
    assign layer6_outputs[3284] = ~(layer5_outputs[4677]);
    assign layer6_outputs[3285] = ~(layer5_outputs[2074]);
    assign layer6_outputs[3286] = layer5_outputs[2285];
    assign layer6_outputs[3287] = layer5_outputs[1162];
    assign layer6_outputs[3288] = ~(layer5_outputs[3490]) | (layer5_outputs[3746]);
    assign layer6_outputs[3289] = layer5_outputs[937];
    assign layer6_outputs[3290] = (layer5_outputs[725]) & (layer5_outputs[2849]);
    assign layer6_outputs[3291] = ~((layer5_outputs[3310]) & (layer5_outputs[3848]));
    assign layer6_outputs[3292] = ~((layer5_outputs[4329]) ^ (layer5_outputs[1475]));
    assign layer6_outputs[3293] = layer5_outputs[4774];
    assign layer6_outputs[3294] = layer5_outputs[4572];
    assign layer6_outputs[3295] = ~((layer5_outputs[2506]) ^ (layer5_outputs[4181]));
    assign layer6_outputs[3296] = ~(layer5_outputs[742]);
    assign layer6_outputs[3297] = (layer5_outputs[2058]) & ~(layer5_outputs[4537]);
    assign layer6_outputs[3298] = ~(layer5_outputs[906]);
    assign layer6_outputs[3299] = (layer5_outputs[4588]) | (layer5_outputs[4390]);
    assign layer6_outputs[3300] = ~((layer5_outputs[3461]) ^ (layer5_outputs[2779]));
    assign layer6_outputs[3301] = ~((layer5_outputs[4659]) ^ (layer5_outputs[1029]));
    assign layer6_outputs[3302] = layer5_outputs[2250];
    assign layer6_outputs[3303] = layer5_outputs[4466];
    assign layer6_outputs[3304] = ~((layer5_outputs[3332]) ^ (layer5_outputs[5000]));
    assign layer6_outputs[3305] = ~((layer5_outputs[616]) ^ (layer5_outputs[3534]));
    assign layer6_outputs[3306] = (layer5_outputs[4093]) & ~(layer5_outputs[5103]);
    assign layer6_outputs[3307] = ~((layer5_outputs[1286]) ^ (layer5_outputs[1094]));
    assign layer6_outputs[3308] = layer5_outputs[938];
    assign layer6_outputs[3309] = ~(layer5_outputs[4840]);
    assign layer6_outputs[3310] = 1'b1;
    assign layer6_outputs[3311] = ~((layer5_outputs[1399]) ^ (layer5_outputs[966]));
    assign layer6_outputs[3312] = ~(layer5_outputs[4665]);
    assign layer6_outputs[3313] = ~(layer5_outputs[2594]) | (layer5_outputs[4270]);
    assign layer6_outputs[3314] = layer5_outputs[1983];
    assign layer6_outputs[3315] = layer5_outputs[1990];
    assign layer6_outputs[3316] = layer5_outputs[445];
    assign layer6_outputs[3317] = (layer5_outputs[859]) | (layer5_outputs[4070]);
    assign layer6_outputs[3318] = ~((layer5_outputs[436]) ^ (layer5_outputs[4300]));
    assign layer6_outputs[3319] = layer5_outputs[3756];
    assign layer6_outputs[3320] = layer5_outputs[3071];
    assign layer6_outputs[3321] = layer5_outputs[3187];
    assign layer6_outputs[3322] = ~(layer5_outputs[148]) | (layer5_outputs[4248]);
    assign layer6_outputs[3323] = (layer5_outputs[1508]) | (layer5_outputs[2485]);
    assign layer6_outputs[3324] = ~(layer5_outputs[4117]);
    assign layer6_outputs[3325] = (layer5_outputs[5112]) & (layer5_outputs[3542]);
    assign layer6_outputs[3326] = ~((layer5_outputs[245]) & (layer5_outputs[680]));
    assign layer6_outputs[3327] = layer5_outputs[2293];
    assign layer6_outputs[3328] = layer5_outputs[3152];
    assign layer6_outputs[3329] = (layer5_outputs[3335]) & (layer5_outputs[4178]);
    assign layer6_outputs[3330] = layer5_outputs[2855];
    assign layer6_outputs[3331] = ~(layer5_outputs[4997]);
    assign layer6_outputs[3332] = (layer5_outputs[2019]) & ~(layer5_outputs[1171]);
    assign layer6_outputs[3333] = (layer5_outputs[2425]) & (layer5_outputs[2491]);
    assign layer6_outputs[3334] = (layer5_outputs[2595]) & (layer5_outputs[1577]);
    assign layer6_outputs[3335] = (layer5_outputs[1466]) & ~(layer5_outputs[1309]);
    assign layer6_outputs[3336] = ~((layer5_outputs[49]) & (layer5_outputs[3098]));
    assign layer6_outputs[3337] = ~(layer5_outputs[2224]);
    assign layer6_outputs[3338] = layer5_outputs[480];
    assign layer6_outputs[3339] = (layer5_outputs[1186]) & ~(layer5_outputs[934]);
    assign layer6_outputs[3340] = layer5_outputs[3072];
    assign layer6_outputs[3341] = ~(layer5_outputs[787]);
    assign layer6_outputs[3342] = (layer5_outputs[4982]) ^ (layer5_outputs[3914]);
    assign layer6_outputs[3343] = ~((layer5_outputs[82]) | (layer5_outputs[3896]));
    assign layer6_outputs[3344] = ~(layer5_outputs[4927]);
    assign layer6_outputs[3345] = ~((layer5_outputs[4481]) ^ (layer5_outputs[2237]));
    assign layer6_outputs[3346] = ~(layer5_outputs[374]);
    assign layer6_outputs[3347] = layer5_outputs[904];
    assign layer6_outputs[3348] = ~(layer5_outputs[407]);
    assign layer6_outputs[3349] = layer5_outputs[142];
    assign layer6_outputs[3350] = 1'b0;
    assign layer6_outputs[3351] = layer5_outputs[2811];
    assign layer6_outputs[3352] = layer5_outputs[4984];
    assign layer6_outputs[3353] = layer5_outputs[2402];
    assign layer6_outputs[3354] = layer5_outputs[4618];
    assign layer6_outputs[3355] = layer5_outputs[3396];
    assign layer6_outputs[3356] = ~(layer5_outputs[2603]);
    assign layer6_outputs[3357] = ~(layer5_outputs[2340]);
    assign layer6_outputs[3358] = layer5_outputs[491];
    assign layer6_outputs[3359] = ~((layer5_outputs[3372]) & (layer5_outputs[3775]));
    assign layer6_outputs[3360] = layer5_outputs[710];
    assign layer6_outputs[3361] = layer5_outputs[111];
    assign layer6_outputs[3362] = ~((layer5_outputs[4014]) ^ (layer5_outputs[961]));
    assign layer6_outputs[3363] = ~(layer5_outputs[623]);
    assign layer6_outputs[3364] = (layer5_outputs[3674]) & ~(layer5_outputs[2724]);
    assign layer6_outputs[3365] = layer5_outputs[1461];
    assign layer6_outputs[3366] = (layer5_outputs[851]) & ~(layer5_outputs[3487]);
    assign layer6_outputs[3367] = layer5_outputs[3033];
    assign layer6_outputs[3368] = layer5_outputs[1874];
    assign layer6_outputs[3369] = ~(layer5_outputs[1846]) | (layer5_outputs[2523]);
    assign layer6_outputs[3370] = layer5_outputs[1342];
    assign layer6_outputs[3371] = ~((layer5_outputs[1006]) | (layer5_outputs[5033]));
    assign layer6_outputs[3372] = (layer5_outputs[2375]) | (layer5_outputs[777]);
    assign layer6_outputs[3373] = ~(layer5_outputs[4328]);
    assign layer6_outputs[3374] = layer5_outputs[433];
    assign layer6_outputs[3375] = ~(layer5_outputs[527]) | (layer5_outputs[2362]);
    assign layer6_outputs[3376] = ~((layer5_outputs[1290]) & (layer5_outputs[129]));
    assign layer6_outputs[3377] = ~((layer5_outputs[1647]) ^ (layer5_outputs[2356]));
    assign layer6_outputs[3378] = ~(layer5_outputs[2717]);
    assign layer6_outputs[3379] = layer5_outputs[4360];
    assign layer6_outputs[3380] = ~((layer5_outputs[1793]) ^ (layer5_outputs[4652]));
    assign layer6_outputs[3381] = ~((layer5_outputs[4798]) & (layer5_outputs[3696]));
    assign layer6_outputs[3382] = ~((layer5_outputs[5096]) | (layer5_outputs[994]));
    assign layer6_outputs[3383] = layer5_outputs[2502];
    assign layer6_outputs[3384] = ~(layer5_outputs[1706]);
    assign layer6_outputs[3385] = ~(layer5_outputs[311]);
    assign layer6_outputs[3386] = ~(layer5_outputs[640]);
    assign layer6_outputs[3387] = (layer5_outputs[1829]) & (layer5_outputs[2970]);
    assign layer6_outputs[3388] = layer5_outputs[208];
    assign layer6_outputs[3389] = ~(layer5_outputs[1507]);
    assign layer6_outputs[3390] = ~((layer5_outputs[715]) ^ (layer5_outputs[3713]));
    assign layer6_outputs[3391] = layer5_outputs[1715];
    assign layer6_outputs[3392] = (layer5_outputs[1999]) & ~(layer5_outputs[2644]);
    assign layer6_outputs[3393] = layer5_outputs[3974];
    assign layer6_outputs[3394] = ~(layer5_outputs[4086]);
    assign layer6_outputs[3395] = (layer5_outputs[1216]) & ~(layer5_outputs[2446]);
    assign layer6_outputs[3396] = ~(layer5_outputs[290]);
    assign layer6_outputs[3397] = layer5_outputs[559];
    assign layer6_outputs[3398] = (layer5_outputs[1640]) | (layer5_outputs[66]);
    assign layer6_outputs[3399] = ~(layer5_outputs[163]);
    assign layer6_outputs[3400] = (layer5_outputs[5070]) | (layer5_outputs[2522]);
    assign layer6_outputs[3401] = (layer5_outputs[3168]) & ~(layer5_outputs[96]);
    assign layer6_outputs[3402] = ~(layer5_outputs[4965]);
    assign layer6_outputs[3403] = ~(layer5_outputs[941]);
    assign layer6_outputs[3404] = ~(layer5_outputs[2919]);
    assign layer6_outputs[3405] = ~(layer5_outputs[3481]);
    assign layer6_outputs[3406] = (layer5_outputs[4003]) ^ (layer5_outputs[2473]);
    assign layer6_outputs[3407] = ~(layer5_outputs[4912]);
    assign layer6_outputs[3408] = (layer5_outputs[321]) | (layer5_outputs[1752]);
    assign layer6_outputs[3409] = (layer5_outputs[1132]) ^ (layer5_outputs[406]);
    assign layer6_outputs[3410] = ~(layer5_outputs[4035]);
    assign layer6_outputs[3411] = ~(layer5_outputs[945]);
    assign layer6_outputs[3412] = ~((layer5_outputs[792]) | (layer5_outputs[4441]));
    assign layer6_outputs[3413] = ~((layer5_outputs[4958]) & (layer5_outputs[434]));
    assign layer6_outputs[3414] = ~((layer5_outputs[3243]) | (layer5_outputs[5110]));
    assign layer6_outputs[3415] = layer5_outputs[855];
    assign layer6_outputs[3416] = ~((layer5_outputs[2753]) ^ (layer5_outputs[2176]));
    assign layer6_outputs[3417] = layer5_outputs[2738];
    assign layer6_outputs[3418] = ~(layer5_outputs[537]);
    assign layer6_outputs[3419] = ~(layer5_outputs[4373]);
    assign layer6_outputs[3420] = ~(layer5_outputs[2809]);
    assign layer6_outputs[3421] = ~(layer5_outputs[2568]);
    assign layer6_outputs[3422] = ~((layer5_outputs[2296]) & (layer5_outputs[2668]));
    assign layer6_outputs[3423] = (layer5_outputs[1918]) & ~(layer5_outputs[4334]);
    assign layer6_outputs[3424] = ~(layer5_outputs[59]) | (layer5_outputs[2588]);
    assign layer6_outputs[3425] = ~(layer5_outputs[2941]) | (layer5_outputs[605]);
    assign layer6_outputs[3426] = (layer5_outputs[2888]) & ~(layer5_outputs[4949]);
    assign layer6_outputs[3427] = 1'b1;
    assign layer6_outputs[3428] = ~((layer5_outputs[4844]) | (layer5_outputs[166]));
    assign layer6_outputs[3429] = layer5_outputs[4025];
    assign layer6_outputs[3430] = layer5_outputs[1119];
    assign layer6_outputs[3431] = (layer5_outputs[1066]) & ~(layer5_outputs[1840]);
    assign layer6_outputs[3432] = layer5_outputs[42];
    assign layer6_outputs[3433] = ~(layer5_outputs[1082]) | (layer5_outputs[1488]);
    assign layer6_outputs[3434] = ~((layer5_outputs[28]) ^ (layer5_outputs[1979]));
    assign layer6_outputs[3435] = layer5_outputs[4784];
    assign layer6_outputs[3436] = ~(layer5_outputs[2280]);
    assign layer6_outputs[3437] = layer5_outputs[5031];
    assign layer6_outputs[3438] = ~(layer5_outputs[96]);
    assign layer6_outputs[3439] = (layer5_outputs[490]) & ~(layer5_outputs[3345]);
    assign layer6_outputs[3440] = layer5_outputs[398];
    assign layer6_outputs[3441] = layer5_outputs[4906];
    assign layer6_outputs[3442] = (layer5_outputs[4696]) & (layer5_outputs[2352]);
    assign layer6_outputs[3443] = ~((layer5_outputs[174]) & (layer5_outputs[5011]));
    assign layer6_outputs[3444] = (layer5_outputs[545]) & ~(layer5_outputs[4614]);
    assign layer6_outputs[3445] = layer5_outputs[3307];
    assign layer6_outputs[3446] = layer5_outputs[3715];
    assign layer6_outputs[3447] = layer5_outputs[3610];
    assign layer6_outputs[3448] = ~((layer5_outputs[2898]) ^ (layer5_outputs[2657]));
    assign layer6_outputs[3449] = ~((layer5_outputs[3921]) ^ (layer5_outputs[974]));
    assign layer6_outputs[3450] = layer5_outputs[2907];
    assign layer6_outputs[3451] = layer5_outputs[255];
    assign layer6_outputs[3452] = ~(layer5_outputs[2152]);
    assign layer6_outputs[3453] = ~(layer5_outputs[4427]);
    assign layer6_outputs[3454] = ~(layer5_outputs[4439]);
    assign layer6_outputs[3455] = ~(layer5_outputs[902]);
    assign layer6_outputs[3456] = layer5_outputs[1174];
    assign layer6_outputs[3457] = (layer5_outputs[4371]) ^ (layer5_outputs[1344]);
    assign layer6_outputs[3458] = layer5_outputs[4723];
    assign layer6_outputs[3459] = layer5_outputs[1037];
    assign layer6_outputs[3460] = ~((layer5_outputs[1388]) ^ (layer5_outputs[2011]));
    assign layer6_outputs[3461] = ~(layer5_outputs[312]);
    assign layer6_outputs[3462] = layer5_outputs[1127];
    assign layer6_outputs[3463] = (layer5_outputs[4692]) & (layer5_outputs[1605]);
    assign layer6_outputs[3464] = (layer5_outputs[4540]) & ~(layer5_outputs[464]);
    assign layer6_outputs[3465] = layer5_outputs[3566];
    assign layer6_outputs[3466] = ~(layer5_outputs[2761]);
    assign layer6_outputs[3467] = ~(layer5_outputs[2556]) | (layer5_outputs[2565]);
    assign layer6_outputs[3468] = ~(layer5_outputs[655]);
    assign layer6_outputs[3469] = (layer5_outputs[285]) & ~(layer5_outputs[3165]);
    assign layer6_outputs[3470] = ~(layer5_outputs[3250]);
    assign layer6_outputs[3471] = 1'b1;
    assign layer6_outputs[3472] = (layer5_outputs[522]) ^ (layer5_outputs[497]);
    assign layer6_outputs[3473] = ~((layer5_outputs[2032]) ^ (layer5_outputs[4192]));
    assign layer6_outputs[3474] = (layer5_outputs[4756]) & ~(layer5_outputs[2460]);
    assign layer6_outputs[3475] = layer5_outputs[69];
    assign layer6_outputs[3476] = ~(layer5_outputs[2424]);
    assign layer6_outputs[3477] = (layer5_outputs[4099]) & ~(layer5_outputs[4087]);
    assign layer6_outputs[3478] = layer5_outputs[699];
    assign layer6_outputs[3479] = layer5_outputs[4344];
    assign layer6_outputs[3480] = ~((layer5_outputs[1967]) ^ (layer5_outputs[4558]));
    assign layer6_outputs[3481] = 1'b0;
    assign layer6_outputs[3482] = ~(layer5_outputs[2157]) | (layer5_outputs[2194]);
    assign layer6_outputs[3483] = ~((layer5_outputs[1573]) ^ (layer5_outputs[2950]));
    assign layer6_outputs[3484] = ~(layer5_outputs[1096]);
    assign layer6_outputs[3485] = ~((layer5_outputs[5048]) ^ (layer5_outputs[2102]));
    assign layer6_outputs[3486] = ~(layer5_outputs[78]);
    assign layer6_outputs[3487] = 1'b1;
    assign layer6_outputs[3488] = layer5_outputs[472];
    assign layer6_outputs[3489] = ~(layer5_outputs[2058]);
    assign layer6_outputs[3490] = ~(layer5_outputs[1492]) | (layer5_outputs[2404]);
    assign layer6_outputs[3491] = ~(layer5_outputs[1316]);
    assign layer6_outputs[3492] = (layer5_outputs[5031]) ^ (layer5_outputs[3414]);
    assign layer6_outputs[3493] = layer5_outputs[2946];
    assign layer6_outputs[3494] = ~((layer5_outputs[315]) | (layer5_outputs[780]));
    assign layer6_outputs[3495] = ~(layer5_outputs[1451]);
    assign layer6_outputs[3496] = ~(layer5_outputs[1773]);
    assign layer6_outputs[3497] = layer5_outputs[1980];
    assign layer6_outputs[3498] = ~(layer5_outputs[2471]);
    assign layer6_outputs[3499] = ~(layer5_outputs[3783]);
    assign layer6_outputs[3500] = (layer5_outputs[467]) & ~(layer5_outputs[2700]);
    assign layer6_outputs[3501] = (layer5_outputs[772]) & (layer5_outputs[167]);
    assign layer6_outputs[3502] = ~(layer5_outputs[998]);
    assign layer6_outputs[3503] = (layer5_outputs[765]) | (layer5_outputs[71]);
    assign layer6_outputs[3504] = (layer5_outputs[4011]) & ~(layer5_outputs[3176]);
    assign layer6_outputs[3505] = 1'b1;
    assign layer6_outputs[3506] = (layer5_outputs[4653]) & ~(layer5_outputs[666]);
    assign layer6_outputs[3507] = (layer5_outputs[455]) | (layer5_outputs[858]);
    assign layer6_outputs[3508] = (layer5_outputs[3191]) ^ (layer5_outputs[2905]);
    assign layer6_outputs[3509] = layer5_outputs[764];
    assign layer6_outputs[3510] = layer5_outputs[707];
    assign layer6_outputs[3511] = (layer5_outputs[3947]) | (layer5_outputs[2926]);
    assign layer6_outputs[3512] = layer5_outputs[494];
    assign layer6_outputs[3513] = ~((layer5_outputs[1016]) ^ (layer5_outputs[3737]));
    assign layer6_outputs[3514] = layer5_outputs[448];
    assign layer6_outputs[3515] = ~(layer5_outputs[114]) | (layer5_outputs[771]);
    assign layer6_outputs[3516] = (layer5_outputs[669]) & ~(layer5_outputs[2754]);
    assign layer6_outputs[3517] = layer5_outputs[3612];
    assign layer6_outputs[3518] = (layer5_outputs[2332]) ^ (layer5_outputs[399]);
    assign layer6_outputs[3519] = ~((layer5_outputs[4182]) | (layer5_outputs[599]));
    assign layer6_outputs[3520] = ~((layer5_outputs[4743]) ^ (layer5_outputs[1252]));
    assign layer6_outputs[3521] = (layer5_outputs[3770]) & ~(layer5_outputs[3194]);
    assign layer6_outputs[3522] = ~(layer5_outputs[766]);
    assign layer6_outputs[3523] = layer5_outputs[46];
    assign layer6_outputs[3524] = (layer5_outputs[3721]) & ~(layer5_outputs[261]);
    assign layer6_outputs[3525] = ~(layer5_outputs[4084]);
    assign layer6_outputs[3526] = ~((layer5_outputs[2706]) ^ (layer5_outputs[2781]));
    assign layer6_outputs[3527] = ~(layer5_outputs[2998]);
    assign layer6_outputs[3528] = layer5_outputs[2545];
    assign layer6_outputs[3529] = layer5_outputs[2750];
    assign layer6_outputs[3530] = (layer5_outputs[3016]) ^ (layer5_outputs[819]);
    assign layer6_outputs[3531] = layer5_outputs[1965];
    assign layer6_outputs[3532] = (layer5_outputs[2407]) ^ (layer5_outputs[4199]);
    assign layer6_outputs[3533] = ~(layer5_outputs[4122]) | (layer5_outputs[1574]);
    assign layer6_outputs[3534] = layer5_outputs[3568];
    assign layer6_outputs[3535] = layer5_outputs[3793];
    assign layer6_outputs[3536] = ~(layer5_outputs[2444]);
    assign layer6_outputs[3537] = ~(layer5_outputs[2117]);
    assign layer6_outputs[3538] = ~(layer5_outputs[1893]);
    assign layer6_outputs[3539] = ~((layer5_outputs[1335]) ^ (layer5_outputs[1214]));
    assign layer6_outputs[3540] = layer5_outputs[35];
    assign layer6_outputs[3541] = ~((layer5_outputs[155]) ^ (layer5_outputs[3921]));
    assign layer6_outputs[3542] = (layer5_outputs[4858]) ^ (layer5_outputs[966]);
    assign layer6_outputs[3543] = 1'b0;
    assign layer6_outputs[3544] = layer5_outputs[4934];
    assign layer6_outputs[3545] = ~(layer5_outputs[2871]);
    assign layer6_outputs[3546] = layer5_outputs[3126];
    assign layer6_outputs[3547] = layer5_outputs[4876];
    assign layer6_outputs[3548] = layer5_outputs[676];
    assign layer6_outputs[3549] = layer5_outputs[2303];
    assign layer6_outputs[3550] = ~(layer5_outputs[4026]);
    assign layer6_outputs[3551] = (layer5_outputs[3196]) & ~(layer5_outputs[3940]);
    assign layer6_outputs[3552] = ~(layer5_outputs[1699]);
    assign layer6_outputs[3553] = ~((layer5_outputs[120]) | (layer5_outputs[473]));
    assign layer6_outputs[3554] = 1'b0;
    assign layer6_outputs[3555] = layer5_outputs[3730];
    assign layer6_outputs[3556] = ~((layer5_outputs[20]) & (layer5_outputs[2766]));
    assign layer6_outputs[3557] = ~((layer5_outputs[714]) ^ (layer5_outputs[1650]));
    assign layer6_outputs[3558] = ~((layer5_outputs[1717]) ^ (layer5_outputs[4352]));
    assign layer6_outputs[3559] = layer5_outputs[2753];
    assign layer6_outputs[3560] = ~(layer5_outputs[3495]);
    assign layer6_outputs[3561] = ~((layer5_outputs[1323]) | (layer5_outputs[4156]));
    assign layer6_outputs[3562] = layer5_outputs[1730];
    assign layer6_outputs[3563] = ~(layer5_outputs[2062]);
    assign layer6_outputs[3564] = ~(layer5_outputs[3288]);
    assign layer6_outputs[3565] = layer5_outputs[79];
    assign layer6_outputs[3566] = (layer5_outputs[610]) ^ (layer5_outputs[839]);
    assign layer6_outputs[3567] = ~(layer5_outputs[1725]);
    assign layer6_outputs[3568] = layer5_outputs[3653];
    assign layer6_outputs[3569] = ~(layer5_outputs[1006]);
    assign layer6_outputs[3570] = ~(layer5_outputs[3819]);
    assign layer6_outputs[3571] = (layer5_outputs[2887]) & (layer5_outputs[1253]);
    assign layer6_outputs[3572] = layer5_outputs[4419];
    assign layer6_outputs[3573] = ~(layer5_outputs[1435]);
    assign layer6_outputs[3574] = ~((layer5_outputs[1526]) & (layer5_outputs[664]));
    assign layer6_outputs[3575] = layer5_outputs[509];
    assign layer6_outputs[3576] = (layer5_outputs[4886]) ^ (layer5_outputs[3458]);
    assign layer6_outputs[3577] = layer5_outputs[3246];
    assign layer6_outputs[3578] = (layer5_outputs[4823]) ^ (layer5_outputs[3387]);
    assign layer6_outputs[3579] = ~(layer5_outputs[3378]);
    assign layer6_outputs[3580] = layer5_outputs[1944];
    assign layer6_outputs[3581] = ~(layer5_outputs[1913]) | (layer5_outputs[4366]);
    assign layer6_outputs[3582] = (layer5_outputs[2647]) | (layer5_outputs[162]);
    assign layer6_outputs[3583] = ~(layer5_outputs[2260]);
    assign layer6_outputs[3584] = ~(layer5_outputs[1610]) | (layer5_outputs[2007]);
    assign layer6_outputs[3585] = (layer5_outputs[939]) & ~(layer5_outputs[4670]);
    assign layer6_outputs[3586] = layer5_outputs[3094];
    assign layer6_outputs[3587] = layer5_outputs[4781];
    assign layer6_outputs[3588] = layer5_outputs[1954];
    assign layer6_outputs[3589] = ~(layer5_outputs[2316]);
    assign layer6_outputs[3590] = (layer5_outputs[1497]) & ~(layer5_outputs[3254]);
    assign layer6_outputs[3591] = layer5_outputs[2018];
    assign layer6_outputs[3592] = layer5_outputs[2943];
    assign layer6_outputs[3593] = ~((layer5_outputs[3082]) & (layer5_outputs[1305]));
    assign layer6_outputs[3594] = layer5_outputs[4072];
    assign layer6_outputs[3595] = ~(layer5_outputs[1941]);
    assign layer6_outputs[3596] = layer5_outputs[4036];
    assign layer6_outputs[3597] = layer5_outputs[2999];
    assign layer6_outputs[3598] = ~(layer5_outputs[519]);
    assign layer6_outputs[3599] = 1'b0;
    assign layer6_outputs[3600] = (layer5_outputs[3584]) & ~(layer5_outputs[93]);
    assign layer6_outputs[3601] = (layer5_outputs[2045]) | (layer5_outputs[4085]);
    assign layer6_outputs[3602] = ~(layer5_outputs[1228]);
    assign layer6_outputs[3603] = ~((layer5_outputs[5037]) | (layer5_outputs[863]));
    assign layer6_outputs[3604] = ~(layer5_outputs[678]);
    assign layer6_outputs[3605] = ~(layer5_outputs[2728]);
    assign layer6_outputs[3606] = ~(layer5_outputs[983]) | (layer5_outputs[649]);
    assign layer6_outputs[3607] = ~((layer5_outputs[2799]) ^ (layer5_outputs[4098]));
    assign layer6_outputs[3608] = ~((layer5_outputs[1340]) ^ (layer5_outputs[322]));
    assign layer6_outputs[3609] = (layer5_outputs[2191]) & ~(layer5_outputs[1933]);
    assign layer6_outputs[3610] = layer5_outputs[2200];
    assign layer6_outputs[3611] = ~((layer5_outputs[1142]) & (layer5_outputs[591]));
    assign layer6_outputs[3612] = ~((layer5_outputs[1074]) | (layer5_outputs[3538]));
    assign layer6_outputs[3613] = ~(layer5_outputs[3669]);
    assign layer6_outputs[3614] = layer5_outputs[3420];
    assign layer6_outputs[3615] = layer5_outputs[3458];
    assign layer6_outputs[3616] = ~(layer5_outputs[396]);
    assign layer6_outputs[3617] = ~((layer5_outputs[2543]) & (layer5_outputs[2178]));
    assign layer6_outputs[3618] = ~((layer5_outputs[2769]) ^ (layer5_outputs[1074]));
    assign layer6_outputs[3619] = (layer5_outputs[3776]) & (layer5_outputs[4715]);
    assign layer6_outputs[3620] = ~((layer5_outputs[1914]) & (layer5_outputs[3445]));
    assign layer6_outputs[3621] = (layer5_outputs[212]) & (layer5_outputs[1958]);
    assign layer6_outputs[3622] = (layer5_outputs[3800]) & (layer5_outputs[4486]);
    assign layer6_outputs[3623] = ~(layer5_outputs[2766]) | (layer5_outputs[4299]);
    assign layer6_outputs[3624] = (layer5_outputs[2951]) & (layer5_outputs[2028]);
    assign layer6_outputs[3625] = ~(layer5_outputs[4553]);
    assign layer6_outputs[3626] = ~(layer5_outputs[208]) | (layer5_outputs[1258]);
    assign layer6_outputs[3627] = (layer5_outputs[849]) ^ (layer5_outputs[1296]);
    assign layer6_outputs[3628] = ~(layer5_outputs[3707]);
    assign layer6_outputs[3629] = ~(layer5_outputs[1372]);
    assign layer6_outputs[3630] = ~(layer5_outputs[3795]);
    assign layer6_outputs[3631] = ~(layer5_outputs[4683]) | (layer5_outputs[1854]);
    assign layer6_outputs[3632] = (layer5_outputs[442]) & ~(layer5_outputs[2263]);
    assign layer6_outputs[3633] = layer5_outputs[2757];
    assign layer6_outputs[3634] = layer5_outputs[1631];
    assign layer6_outputs[3635] = (layer5_outputs[2966]) ^ (layer5_outputs[551]);
    assign layer6_outputs[3636] = (layer5_outputs[1433]) | (layer5_outputs[1896]);
    assign layer6_outputs[3637] = ~((layer5_outputs[923]) & (layer5_outputs[2081]));
    assign layer6_outputs[3638] = ~(layer5_outputs[2043]);
    assign layer6_outputs[3639] = ~(layer5_outputs[3851]);
    assign layer6_outputs[3640] = ~(layer5_outputs[4170]) | (layer5_outputs[587]);
    assign layer6_outputs[3641] = ~((layer5_outputs[3191]) ^ (layer5_outputs[4073]));
    assign layer6_outputs[3642] = ~(layer5_outputs[3647]);
    assign layer6_outputs[3643] = layer5_outputs[3870];
    assign layer6_outputs[3644] = layer5_outputs[1786];
    assign layer6_outputs[3645] = (layer5_outputs[1025]) & (layer5_outputs[2716]);
    assign layer6_outputs[3646] = ~(layer5_outputs[1955]) | (layer5_outputs[3394]);
    assign layer6_outputs[3647] = ~(layer5_outputs[1477]);
    assign layer6_outputs[3648] = ~(layer5_outputs[3734]) | (layer5_outputs[65]);
    assign layer6_outputs[3649] = ~((layer5_outputs[4746]) & (layer5_outputs[5020]));
    assign layer6_outputs[3650] = ~(layer5_outputs[1125]) | (layer5_outputs[5105]);
    assign layer6_outputs[3651] = layer5_outputs[3514];
    assign layer6_outputs[3652] = (layer5_outputs[2639]) & ~(layer5_outputs[1638]);
    assign layer6_outputs[3653] = ~((layer5_outputs[856]) ^ (layer5_outputs[4513]));
    assign layer6_outputs[3654] = ~(layer5_outputs[368]);
    assign layer6_outputs[3655] = 1'b1;
    assign layer6_outputs[3656] = layer5_outputs[4033];
    assign layer6_outputs[3657] = layer5_outputs[4035];
    assign layer6_outputs[3658] = ~((layer5_outputs[373]) & (layer5_outputs[462]));
    assign layer6_outputs[3659] = (layer5_outputs[273]) ^ (layer5_outputs[1825]);
    assign layer6_outputs[3660] = (layer5_outputs[3485]) | (layer5_outputs[1734]);
    assign layer6_outputs[3661] = (layer5_outputs[2654]) & (layer5_outputs[2202]);
    assign layer6_outputs[3662] = ~(layer5_outputs[3225]);
    assign layer6_outputs[3663] = ~(layer5_outputs[4789]);
    assign layer6_outputs[3664] = ~((layer5_outputs[39]) & (layer5_outputs[4642]));
    assign layer6_outputs[3665] = (layer5_outputs[4795]) ^ (layer5_outputs[4194]);
    assign layer6_outputs[3666] = layer5_outputs[1872];
    assign layer6_outputs[3667] = ~(layer5_outputs[3662]);
    assign layer6_outputs[3668] = (layer5_outputs[1071]) & ~(layer5_outputs[214]);
    assign layer6_outputs[3669] = ~(layer5_outputs[2650]);
    assign layer6_outputs[3670] = (layer5_outputs[4501]) & ~(layer5_outputs[4635]);
    assign layer6_outputs[3671] = layer5_outputs[3669];
    assign layer6_outputs[3672] = ~((layer5_outputs[4319]) & (layer5_outputs[3197]));
    assign layer6_outputs[3673] = (layer5_outputs[1808]) & (layer5_outputs[690]);
    assign layer6_outputs[3674] = layer5_outputs[3009];
    assign layer6_outputs[3675] = (layer5_outputs[124]) & ~(layer5_outputs[1337]);
    assign layer6_outputs[3676] = ~(layer5_outputs[1352]) | (layer5_outputs[4120]);
    assign layer6_outputs[3677] = layer5_outputs[1534];
    assign layer6_outputs[3678] = ~(layer5_outputs[2089]);
    assign layer6_outputs[3679] = ~((layer5_outputs[2300]) ^ (layer5_outputs[45]));
    assign layer6_outputs[3680] = layer5_outputs[2];
    assign layer6_outputs[3681] = ~(layer5_outputs[924]);
    assign layer6_outputs[3682] = (layer5_outputs[4133]) & ~(layer5_outputs[2343]);
    assign layer6_outputs[3683] = layer5_outputs[739];
    assign layer6_outputs[3684] = ~(layer5_outputs[1206]) | (layer5_outputs[2353]);
    assign layer6_outputs[3685] = (layer5_outputs[2878]) ^ (layer5_outputs[5015]);
    assign layer6_outputs[3686] = ~(layer5_outputs[3148]);
    assign layer6_outputs[3687] = 1'b0;
    assign layer6_outputs[3688] = layer5_outputs[165];
    assign layer6_outputs[3689] = layer5_outputs[1170];
    assign layer6_outputs[3690] = (layer5_outputs[3027]) & (layer5_outputs[1453]);
    assign layer6_outputs[3691] = layer5_outputs[3403];
    assign layer6_outputs[3692] = layer5_outputs[3556];
    assign layer6_outputs[3693] = layer5_outputs[4641];
    assign layer6_outputs[3694] = (layer5_outputs[1336]) & ~(layer5_outputs[2693]);
    assign layer6_outputs[3695] = ~(layer5_outputs[2144]);
    assign layer6_outputs[3696] = ~(layer5_outputs[3630]);
    assign layer6_outputs[3697] = ~(layer5_outputs[2723]) | (layer5_outputs[233]);
    assign layer6_outputs[3698] = (layer5_outputs[2089]) & ~(layer5_outputs[3517]);
    assign layer6_outputs[3699] = ~(layer5_outputs[1747]);
    assign layer6_outputs[3700] = (layer5_outputs[4169]) & (layer5_outputs[823]);
    assign layer6_outputs[3701] = (layer5_outputs[821]) & ~(layer5_outputs[4794]);
    assign layer6_outputs[3702] = ~((layer5_outputs[1555]) ^ (layer5_outputs[1165]));
    assign layer6_outputs[3703] = ~((layer5_outputs[3325]) | (layer5_outputs[2948]));
    assign layer6_outputs[3704] = ~(layer5_outputs[4463]) | (layer5_outputs[4602]);
    assign layer6_outputs[3705] = ~((layer5_outputs[2597]) | (layer5_outputs[1511]));
    assign layer6_outputs[3706] = ~(layer5_outputs[1450]);
    assign layer6_outputs[3707] = ~(layer5_outputs[1804]);
    assign layer6_outputs[3708] = ~(layer5_outputs[3002]) | (layer5_outputs[4725]);
    assign layer6_outputs[3709] = layer5_outputs[1773];
    assign layer6_outputs[3710] = (layer5_outputs[2507]) & ~(layer5_outputs[2399]);
    assign layer6_outputs[3711] = ~(layer5_outputs[398]);
    assign layer6_outputs[3712] = ~(layer5_outputs[337]);
    assign layer6_outputs[3713] = layer5_outputs[1968];
    assign layer6_outputs[3714] = ~(layer5_outputs[721]);
    assign layer6_outputs[3715] = ~((layer5_outputs[4139]) & (layer5_outputs[2630]));
    assign layer6_outputs[3716] = (layer5_outputs[4308]) & ~(layer5_outputs[277]);
    assign layer6_outputs[3717] = ~(layer5_outputs[586]) | (layer5_outputs[305]);
    assign layer6_outputs[3718] = ~((layer5_outputs[3900]) ^ (layer5_outputs[675]));
    assign layer6_outputs[3719] = ~(layer5_outputs[2079]) | (layer5_outputs[4503]);
    assign layer6_outputs[3720] = layer5_outputs[3714];
    assign layer6_outputs[3721] = layer5_outputs[1877];
    assign layer6_outputs[3722] = ~(layer5_outputs[1343]);
    assign layer6_outputs[3723] = ~(layer5_outputs[1472]);
    assign layer6_outputs[3724] = (layer5_outputs[1279]) & ~(layer5_outputs[3611]);
    assign layer6_outputs[3725] = (layer5_outputs[2350]) & (layer5_outputs[4219]);
    assign layer6_outputs[3726] = ~((layer5_outputs[2609]) | (layer5_outputs[3371]));
    assign layer6_outputs[3727] = ~((layer5_outputs[3864]) ^ (layer5_outputs[4308]));
    assign layer6_outputs[3728] = ~((layer5_outputs[4751]) ^ (layer5_outputs[3540]));
    assign layer6_outputs[3729] = (layer5_outputs[66]) | (layer5_outputs[621]);
    assign layer6_outputs[3730] = (layer5_outputs[227]) & (layer5_outputs[4114]);
    assign layer6_outputs[3731] = layer5_outputs[3672];
    assign layer6_outputs[3732] = 1'b0;
    assign layer6_outputs[3733] = layer5_outputs[2396];
    assign layer6_outputs[3734] = ~(layer5_outputs[4541]) | (layer5_outputs[2096]);
    assign layer6_outputs[3735] = layer5_outputs[758];
    assign layer6_outputs[3736] = ~(layer5_outputs[1780]);
    assign layer6_outputs[3737] = (layer5_outputs[3711]) & ~(layer5_outputs[3453]);
    assign layer6_outputs[3738] = ~(layer5_outputs[3180]);
    assign layer6_outputs[3739] = ~((layer5_outputs[1427]) | (layer5_outputs[5030]));
    assign layer6_outputs[3740] = (layer5_outputs[1114]) & ~(layer5_outputs[4105]);
    assign layer6_outputs[3741] = layer5_outputs[4552];
    assign layer6_outputs[3742] = ~(layer5_outputs[4467]);
    assign layer6_outputs[3743] = ~(layer5_outputs[348]);
    assign layer6_outputs[3744] = layer5_outputs[2870];
    assign layer6_outputs[3745] = ~(layer5_outputs[513]);
    assign layer6_outputs[3746] = layer5_outputs[4372];
    assign layer6_outputs[3747] = ~(layer5_outputs[1593]);
    assign layer6_outputs[3748] = ~(layer5_outputs[2905]);
    assign layer6_outputs[3749] = ~(layer5_outputs[3567]);
    assign layer6_outputs[3750] = ~(layer5_outputs[1529]);
    assign layer6_outputs[3751] = ~((layer5_outputs[3324]) | (layer5_outputs[2297]));
    assign layer6_outputs[3752] = ~(layer5_outputs[5091]);
    assign layer6_outputs[3753] = ~(layer5_outputs[2537]) | (layer5_outputs[3056]);
    assign layer6_outputs[3754] = ~(layer5_outputs[3493]);
    assign layer6_outputs[3755] = ~((layer5_outputs[47]) | (layer5_outputs[3566]));
    assign layer6_outputs[3756] = layer5_outputs[2121];
    assign layer6_outputs[3757] = layer5_outputs[1980];
    assign layer6_outputs[3758] = layer5_outputs[3879];
    assign layer6_outputs[3759] = layer5_outputs[3459];
    assign layer6_outputs[3760] = ~((layer5_outputs[1405]) ^ (layer5_outputs[3203]));
    assign layer6_outputs[3761] = ~((layer5_outputs[688]) & (layer5_outputs[1456]));
    assign layer6_outputs[3762] = ~((layer5_outputs[3955]) ^ (layer5_outputs[3862]));
    assign layer6_outputs[3763] = layer5_outputs[2197];
    assign layer6_outputs[3764] = ~(layer5_outputs[4297]) | (layer5_outputs[1371]);
    assign layer6_outputs[3765] = ~((layer5_outputs[1898]) & (layer5_outputs[2834]));
    assign layer6_outputs[3766] = (layer5_outputs[539]) ^ (layer5_outputs[4397]);
    assign layer6_outputs[3767] = layer5_outputs[4877];
    assign layer6_outputs[3768] = (layer5_outputs[815]) | (layer5_outputs[4243]);
    assign layer6_outputs[3769] = ~((layer5_outputs[915]) ^ (layer5_outputs[1148]));
    assign layer6_outputs[3770] = ~((layer5_outputs[4778]) ^ (layer5_outputs[1145]));
    assign layer6_outputs[3771] = layer5_outputs[769];
    assign layer6_outputs[3772] = layer5_outputs[2436];
    assign layer6_outputs[3773] = layer5_outputs[3425];
    assign layer6_outputs[3774] = layer5_outputs[98];
    assign layer6_outputs[3775] = ~((layer5_outputs[2715]) | (layer5_outputs[4528]));
    assign layer6_outputs[3776] = ~(layer5_outputs[2939]);
    assign layer6_outputs[3777] = ~(layer5_outputs[4266]);
    assign layer6_outputs[3778] = layer5_outputs[4595];
    assign layer6_outputs[3779] = ~((layer5_outputs[1841]) & (layer5_outputs[2464]));
    assign layer6_outputs[3780] = ~(layer5_outputs[2005]);
    assign layer6_outputs[3781] = ~(layer5_outputs[4183]);
    assign layer6_outputs[3782] = layer5_outputs[373];
    assign layer6_outputs[3783] = ~(layer5_outputs[4030]);
    assign layer6_outputs[3784] = layer5_outputs[240];
    assign layer6_outputs[3785] = (layer5_outputs[456]) | (layer5_outputs[172]);
    assign layer6_outputs[3786] = layer5_outputs[3242];
    assign layer6_outputs[3787] = ~(layer5_outputs[3949]) | (layer5_outputs[3075]);
    assign layer6_outputs[3788] = layer5_outputs[429];
    assign layer6_outputs[3789] = layer5_outputs[3144];
    assign layer6_outputs[3790] = ~(layer5_outputs[3180]);
    assign layer6_outputs[3791] = (layer5_outputs[539]) ^ (layer5_outputs[357]);
    assign layer6_outputs[3792] = ~(layer5_outputs[970]);
    assign layer6_outputs[3793] = ~(layer5_outputs[316]);
    assign layer6_outputs[3794] = 1'b1;
    assign layer6_outputs[3795] = ~(layer5_outputs[3369]);
    assign layer6_outputs[3796] = (layer5_outputs[740]) & ~(layer5_outputs[1501]);
    assign layer6_outputs[3797] = layer5_outputs[3375];
    assign layer6_outputs[3798] = layer5_outputs[2173];
    assign layer6_outputs[3799] = 1'b0;
    assign layer6_outputs[3800] = ~(layer5_outputs[4381]) | (layer5_outputs[4774]);
    assign layer6_outputs[3801] = ~((layer5_outputs[2632]) | (layer5_outputs[1907]));
    assign layer6_outputs[3802] = layer5_outputs[2287];
    assign layer6_outputs[3803] = ~(layer5_outputs[1349]);
    assign layer6_outputs[3804] = ~(layer5_outputs[176]);
    assign layer6_outputs[3805] = ~((layer5_outputs[4244]) ^ (layer5_outputs[4596]));
    assign layer6_outputs[3806] = (layer5_outputs[1372]) ^ (layer5_outputs[3401]);
    assign layer6_outputs[3807] = 1'b1;
    assign layer6_outputs[3808] = layer5_outputs[1584];
    assign layer6_outputs[3809] = (layer5_outputs[706]) & ~(layer5_outputs[2183]);
    assign layer6_outputs[3810] = ~(layer5_outputs[4015]);
    assign layer6_outputs[3811] = ~(layer5_outputs[549]);
    assign layer6_outputs[3812] = (layer5_outputs[649]) ^ (layer5_outputs[1169]);
    assign layer6_outputs[3813] = ~(layer5_outputs[1560]);
    assign layer6_outputs[3814] = ~(layer5_outputs[2357]) | (layer5_outputs[2419]);
    assign layer6_outputs[3815] = (layer5_outputs[1056]) ^ (layer5_outputs[2732]);
    assign layer6_outputs[3816] = (layer5_outputs[4272]) & (layer5_outputs[4185]);
    assign layer6_outputs[3817] = layer5_outputs[4636];
    assign layer6_outputs[3818] = layer5_outputs[895];
    assign layer6_outputs[3819] = ~(layer5_outputs[688]) | (layer5_outputs[1198]);
    assign layer6_outputs[3820] = ~((layer5_outputs[4137]) | (layer5_outputs[3610]));
    assign layer6_outputs[3821] = layer5_outputs[4597];
    assign layer6_outputs[3822] = layer5_outputs[80];
    assign layer6_outputs[3823] = layer5_outputs[3967];
    assign layer6_outputs[3824] = layer5_outputs[3168];
    assign layer6_outputs[3825] = ~(layer5_outputs[3408]);
    assign layer6_outputs[3826] = ~((layer5_outputs[663]) & (layer5_outputs[2651]));
    assign layer6_outputs[3827] = ~((layer5_outputs[3515]) ^ (layer5_outputs[121]));
    assign layer6_outputs[3828] = layer5_outputs[547];
    assign layer6_outputs[3829] = (layer5_outputs[4185]) & ~(layer5_outputs[1040]);
    assign layer6_outputs[3830] = ~((layer5_outputs[504]) & (layer5_outputs[2369]));
    assign layer6_outputs[3831] = ~(layer5_outputs[2071]);
    assign layer6_outputs[3832] = (layer5_outputs[4839]) | (layer5_outputs[2949]);
    assign layer6_outputs[3833] = ~(layer5_outputs[530]);
    assign layer6_outputs[3834] = ~((layer5_outputs[4173]) ^ (layer5_outputs[376]));
    assign layer6_outputs[3835] = layer5_outputs[4943];
    assign layer6_outputs[3836] = layer5_outputs[1727];
    assign layer6_outputs[3837] = layer5_outputs[424];
    assign layer6_outputs[3838] = ~(layer5_outputs[4702]);
    assign layer6_outputs[3839] = ~((layer5_outputs[3977]) ^ (layer5_outputs[711]));
    assign layer6_outputs[3840] = ~(layer5_outputs[1033]);
    assign layer6_outputs[3841] = layer5_outputs[2535];
    assign layer6_outputs[3842] = ~(layer5_outputs[788]) | (layer5_outputs[309]);
    assign layer6_outputs[3843] = ~((layer5_outputs[319]) ^ (layer5_outputs[3316]));
    assign layer6_outputs[3844] = ~(layer5_outputs[2936]);
    assign layer6_outputs[3845] = (layer5_outputs[4218]) | (layer5_outputs[3600]);
    assign layer6_outputs[3846] = ~((layer5_outputs[4478]) ^ (layer5_outputs[1521]));
    assign layer6_outputs[3847] = layer5_outputs[60];
    assign layer6_outputs[3848] = (layer5_outputs[4651]) & ~(layer5_outputs[4022]);
    assign layer6_outputs[3849] = ~(layer5_outputs[123]);
    assign layer6_outputs[3850] = ~(layer5_outputs[3204]);
    assign layer6_outputs[3851] = (layer5_outputs[1919]) ^ (layer5_outputs[4810]);
    assign layer6_outputs[3852] = layer5_outputs[39];
    assign layer6_outputs[3853] = layer5_outputs[728];
    assign layer6_outputs[3854] = ~((layer5_outputs[2765]) | (layer5_outputs[2019]));
    assign layer6_outputs[3855] = 1'b1;
    assign layer6_outputs[3856] = layer5_outputs[3788];
    assign layer6_outputs[3857] = layer5_outputs[4270];
    assign layer6_outputs[3858] = ~(layer5_outputs[1925]);
    assign layer6_outputs[3859] = layer5_outputs[2531];
    assign layer6_outputs[3860] = 1'b0;
    assign layer6_outputs[3861] = ~((layer5_outputs[4871]) ^ (layer5_outputs[4203]));
    assign layer6_outputs[3862] = ~(layer5_outputs[2199]);
    assign layer6_outputs[3863] = ~(layer5_outputs[865]);
    assign layer6_outputs[3864] = ~((layer5_outputs[173]) & (layer5_outputs[2608]));
    assign layer6_outputs[3865] = ~((layer5_outputs[5066]) | (layer5_outputs[527]));
    assign layer6_outputs[3866] = ~(layer5_outputs[509]);
    assign layer6_outputs[3867] = layer5_outputs[695];
    assign layer6_outputs[3868] = (layer5_outputs[4625]) | (layer5_outputs[3656]);
    assign layer6_outputs[3869] = layer5_outputs[4090];
    assign layer6_outputs[3870] = ~(layer5_outputs[818]) | (layer5_outputs[1335]);
    assign layer6_outputs[3871] = 1'b0;
    assign layer6_outputs[3872] = (layer5_outputs[2515]) & ~(layer5_outputs[4408]);
    assign layer6_outputs[3873] = ~(layer5_outputs[2121]);
    assign layer6_outputs[3874] = layer5_outputs[1933];
    assign layer6_outputs[3875] = ~((layer5_outputs[4634]) & (layer5_outputs[3571]));
    assign layer6_outputs[3876] = ~((layer5_outputs[1120]) ^ (layer5_outputs[1153]));
    assign layer6_outputs[3877] = ~(layer5_outputs[2424]);
    assign layer6_outputs[3878] = ~((layer5_outputs[4304]) | (layer5_outputs[946]));
    assign layer6_outputs[3879] = ~(layer5_outputs[2782]);
    assign layer6_outputs[3880] = (layer5_outputs[443]) | (layer5_outputs[826]);
    assign layer6_outputs[3881] = (layer5_outputs[1100]) ^ (layer5_outputs[1714]);
    assign layer6_outputs[3882] = layer5_outputs[1788];
    assign layer6_outputs[3883] = (layer5_outputs[4549]) & ~(layer5_outputs[3871]);
    assign layer6_outputs[3884] = ~((layer5_outputs[5061]) & (layer5_outputs[2512]));
    assign layer6_outputs[3885] = layer5_outputs[150];
    assign layer6_outputs[3886] = ~(layer5_outputs[1882]);
    assign layer6_outputs[3887] = layer5_outputs[297];
    assign layer6_outputs[3888] = layer5_outputs[1271];
    assign layer6_outputs[3889] = ~(layer5_outputs[711]);
    assign layer6_outputs[3890] = layer5_outputs[4151];
    assign layer6_outputs[3891] = 1'b0;
    assign layer6_outputs[3892] = ~(layer5_outputs[2185]);
    assign layer6_outputs[3893] = ~((layer5_outputs[2488]) ^ (layer5_outputs[756]));
    assign layer6_outputs[3894] = layer5_outputs[3456];
    assign layer6_outputs[3895] = (layer5_outputs[4017]) ^ (layer5_outputs[313]);
    assign layer6_outputs[3896] = ~(layer5_outputs[692]) | (layer5_outputs[2110]);
    assign layer6_outputs[3897] = layer5_outputs[1262];
    assign layer6_outputs[3898] = (layer5_outputs[3025]) ^ (layer5_outputs[1548]);
    assign layer6_outputs[3899] = (layer5_outputs[1283]) ^ (layer5_outputs[1499]);
    assign layer6_outputs[3900] = ~(layer5_outputs[4541]);
    assign layer6_outputs[3901] = layer5_outputs[3966];
    assign layer6_outputs[3902] = ~(layer5_outputs[3387]);
    assign layer6_outputs[3903] = (layer5_outputs[3684]) ^ (layer5_outputs[3461]);
    assign layer6_outputs[3904] = ~((layer5_outputs[2729]) & (layer5_outputs[119]));
    assign layer6_outputs[3905] = ~((layer5_outputs[2239]) | (layer5_outputs[3110]));
    assign layer6_outputs[3906] = ~(layer5_outputs[4300]);
    assign layer6_outputs[3907] = layer5_outputs[1943];
    assign layer6_outputs[3908] = ~((layer5_outputs[1310]) & (layer5_outputs[353]));
    assign layer6_outputs[3909] = (layer5_outputs[3579]) ^ (layer5_outputs[4417]);
    assign layer6_outputs[3910] = (layer5_outputs[5017]) | (layer5_outputs[603]);
    assign layer6_outputs[3911] = ~(layer5_outputs[691]) | (layer5_outputs[615]);
    assign layer6_outputs[3912] = ~(layer5_outputs[1289]);
    assign layer6_outputs[3913] = ~(layer5_outputs[4386]);
    assign layer6_outputs[3914] = layer5_outputs[3421];
    assign layer6_outputs[3915] = ~(layer5_outputs[3748]);
    assign layer6_outputs[3916] = layer5_outputs[2300];
    assign layer6_outputs[3917] = layer5_outputs[4019];
    assign layer6_outputs[3918] = (layer5_outputs[1161]) & ~(layer5_outputs[4705]);
    assign layer6_outputs[3919] = ~(layer5_outputs[1530]);
    assign layer6_outputs[3920] = (layer5_outputs[4645]) ^ (layer5_outputs[2481]);
    assign layer6_outputs[3921] = ~(layer5_outputs[2964]);
    assign layer6_outputs[3922] = ~(layer5_outputs[3449]);
    assign layer6_outputs[3923] = (layer5_outputs[104]) ^ (layer5_outputs[867]);
    assign layer6_outputs[3924] = ~(layer5_outputs[2270]);
    assign layer6_outputs[3925] = (layer5_outputs[2771]) | (layer5_outputs[2574]);
    assign layer6_outputs[3926] = layer5_outputs[4560];
    assign layer6_outputs[3927] = (layer5_outputs[4508]) & (layer5_outputs[4310]);
    assign layer6_outputs[3928] = layer5_outputs[674];
    assign layer6_outputs[3929] = ~((layer5_outputs[898]) ^ (layer5_outputs[389]));
    assign layer6_outputs[3930] = layer5_outputs[2863];
    assign layer6_outputs[3931] = layer5_outputs[1142];
    assign layer6_outputs[3932] = (layer5_outputs[3160]) ^ (layer5_outputs[3932]);
    assign layer6_outputs[3933] = ~(layer5_outputs[2570]);
    assign layer6_outputs[3934] = (layer5_outputs[1934]) | (layer5_outputs[1215]);
    assign layer6_outputs[3935] = ~((layer5_outputs[3408]) ^ (layer5_outputs[1314]));
    assign layer6_outputs[3936] = layer5_outputs[1151];
    assign layer6_outputs[3937] = layer5_outputs[1578];
    assign layer6_outputs[3938] = layer5_outputs[3222];
    assign layer6_outputs[3939] = ~(layer5_outputs[1939]) | (layer5_outputs[1738]);
    assign layer6_outputs[3940] = layer5_outputs[1779];
    assign layer6_outputs[3941] = ~(layer5_outputs[2132]);
    assign layer6_outputs[3942] = (layer5_outputs[3635]) ^ (layer5_outputs[1202]);
    assign layer6_outputs[3943] = (layer5_outputs[1862]) | (layer5_outputs[1715]);
    assign layer6_outputs[3944] = layer5_outputs[4947];
    assign layer6_outputs[3945] = (layer5_outputs[340]) ^ (layer5_outputs[4275]);
    assign layer6_outputs[3946] = (layer5_outputs[2579]) & (layer5_outputs[1237]);
    assign layer6_outputs[3947] = (layer5_outputs[2678]) ^ (layer5_outputs[522]);
    assign layer6_outputs[3948] = (layer5_outputs[304]) | (layer5_outputs[4625]);
    assign layer6_outputs[3949] = ~(layer5_outputs[4027]);
    assign layer6_outputs[3950] = ~(layer5_outputs[971]);
    assign layer6_outputs[3951] = ~((layer5_outputs[4510]) & (layer5_outputs[776]));
    assign layer6_outputs[3952] = (layer5_outputs[1297]) ^ (layer5_outputs[1587]);
    assign layer6_outputs[3953] = ~(layer5_outputs[1079]);
    assign layer6_outputs[3954] = (layer5_outputs[2915]) & ~(layer5_outputs[1569]);
    assign layer6_outputs[3955] = layer5_outputs[5099];
    assign layer6_outputs[3956] = ~(layer5_outputs[18]);
    assign layer6_outputs[3957] = (layer5_outputs[1680]) & ~(layer5_outputs[2170]);
    assign layer6_outputs[3958] = ~((layer5_outputs[3816]) ^ (layer5_outputs[3451]));
    assign layer6_outputs[3959] = (layer5_outputs[24]) ^ (layer5_outputs[1879]);
    assign layer6_outputs[3960] = ~(layer5_outputs[335]) | (layer5_outputs[4199]);
    assign layer6_outputs[3961] = ~(layer5_outputs[2800]);
    assign layer6_outputs[3962] = layer5_outputs[2209];
    assign layer6_outputs[3963] = (layer5_outputs[4757]) & ~(layer5_outputs[141]);
    assign layer6_outputs[3964] = layer5_outputs[3338];
    assign layer6_outputs[3965] = (layer5_outputs[785]) & ~(layer5_outputs[4797]);
    assign layer6_outputs[3966] = (layer5_outputs[478]) | (layer5_outputs[2061]);
    assign layer6_outputs[3967] = (layer5_outputs[665]) & (layer5_outputs[4081]);
    assign layer6_outputs[3968] = (layer5_outputs[623]) | (layer5_outputs[1042]);
    assign layer6_outputs[3969] = ~((layer5_outputs[3769]) ^ (layer5_outputs[1808]));
    assign layer6_outputs[3970] = layer5_outputs[139];
    assign layer6_outputs[3971] = layer5_outputs[3509];
    assign layer6_outputs[3972] = layer5_outputs[1643];
    assign layer6_outputs[3973] = (layer5_outputs[185]) | (layer5_outputs[4098]);
    assign layer6_outputs[3974] = ~(layer5_outputs[2047]);
    assign layer6_outputs[3975] = ~(layer5_outputs[3122]);
    assign layer6_outputs[3976] = ~(layer5_outputs[106]) | (layer5_outputs[3092]);
    assign layer6_outputs[3977] = ~(layer5_outputs[4484]);
    assign layer6_outputs[3978] = ~(layer5_outputs[389]);
    assign layer6_outputs[3979] = ~(layer5_outputs[2559]);
    assign layer6_outputs[3980] = ~(layer5_outputs[2873]) | (layer5_outputs[5108]);
    assign layer6_outputs[3981] = ~(layer5_outputs[1695]);
    assign layer6_outputs[3982] = ~((layer5_outputs[4324]) & (layer5_outputs[299]));
    assign layer6_outputs[3983] = ~(layer5_outputs[4705]);
    assign layer6_outputs[3984] = ~((layer5_outputs[1407]) ^ (layer5_outputs[1582]));
    assign layer6_outputs[3985] = (layer5_outputs[3001]) & ~(layer5_outputs[5039]);
    assign layer6_outputs[3986] = ~(layer5_outputs[2279]);
    assign layer6_outputs[3987] = layer5_outputs[4810];
    assign layer6_outputs[3988] = ~(layer5_outputs[138]);
    assign layer6_outputs[3989] = ~((layer5_outputs[5014]) ^ (layer5_outputs[2846]));
    assign layer6_outputs[3990] = ~((layer5_outputs[730]) & (layer5_outputs[2214]));
    assign layer6_outputs[3991] = ~((layer5_outputs[4071]) ^ (layer5_outputs[163]));
    assign layer6_outputs[3992] = ~(layer5_outputs[83]);
    assign layer6_outputs[3993] = (layer5_outputs[1844]) & ~(layer5_outputs[4106]);
    assign layer6_outputs[3994] = (layer5_outputs[668]) ^ (layer5_outputs[1672]);
    assign layer6_outputs[3995] = layer5_outputs[5053];
    assign layer6_outputs[3996] = layer5_outputs[2434];
    assign layer6_outputs[3997] = ~(layer5_outputs[1147]);
    assign layer6_outputs[3998] = ~(layer5_outputs[2282]);
    assign layer6_outputs[3999] = (layer5_outputs[4374]) ^ (layer5_outputs[2351]);
    assign layer6_outputs[4000] = ~(layer5_outputs[1712]) | (layer5_outputs[3941]);
    assign layer6_outputs[4001] = layer5_outputs[3213];
    assign layer6_outputs[4002] = ~((layer5_outputs[1204]) ^ (layer5_outputs[1110]));
    assign layer6_outputs[4003] = layer5_outputs[1180];
    assign layer6_outputs[4004] = (layer5_outputs[658]) & ~(layer5_outputs[1723]);
    assign layer6_outputs[4005] = (layer5_outputs[1243]) & ~(layer5_outputs[3933]);
    assign layer6_outputs[4006] = ~(layer5_outputs[4762]);
    assign layer6_outputs[4007] = ~(layer5_outputs[3931]);
    assign layer6_outputs[4008] = ~((layer5_outputs[2654]) | (layer5_outputs[1313]));
    assign layer6_outputs[4009] = ~(layer5_outputs[3699]) | (layer5_outputs[1557]);
    assign layer6_outputs[4010] = layer5_outputs[2119];
    assign layer6_outputs[4011] = ~(layer5_outputs[3033]) | (layer5_outputs[4903]);
    assign layer6_outputs[4012] = ~((layer5_outputs[2503]) ^ (layer5_outputs[4440]));
    assign layer6_outputs[4013] = ~(layer5_outputs[4821]);
    assign layer6_outputs[4014] = layer5_outputs[2271];
    assign layer6_outputs[4015] = layer5_outputs[4089];
    assign layer6_outputs[4016] = ~(layer5_outputs[556]);
    assign layer6_outputs[4017] = ~((layer5_outputs[933]) ^ (layer5_outputs[1200]));
    assign layer6_outputs[4018] = (layer5_outputs[1058]) & (layer5_outputs[540]);
    assign layer6_outputs[4019] = (layer5_outputs[2102]) ^ (layer5_outputs[535]);
    assign layer6_outputs[4020] = ~(layer5_outputs[2590]);
    assign layer6_outputs[4021] = ~(layer5_outputs[453]);
    assign layer6_outputs[4022] = ~(layer5_outputs[3209]) | (layer5_outputs[1051]);
    assign layer6_outputs[4023] = ~(layer5_outputs[2043]);
    assign layer6_outputs[4024] = ~(layer5_outputs[3838]) | (layer5_outputs[3757]);
    assign layer6_outputs[4025] = ~(layer5_outputs[813]);
    assign layer6_outputs[4026] = (layer5_outputs[3143]) & ~(layer5_outputs[554]);
    assign layer6_outputs[4027] = layer5_outputs[4972];
    assign layer6_outputs[4028] = ~((layer5_outputs[2113]) ^ (layer5_outputs[3361]));
    assign layer6_outputs[4029] = ~(layer5_outputs[1561]) | (layer5_outputs[358]);
    assign layer6_outputs[4030] = (layer5_outputs[2179]) ^ (layer5_outputs[1754]);
    assign layer6_outputs[4031] = (layer5_outputs[507]) ^ (layer5_outputs[1094]);
    assign layer6_outputs[4032] = (layer5_outputs[630]) & (layer5_outputs[489]);
    assign layer6_outputs[4033] = ~((layer5_outputs[3810]) & (layer5_outputs[51]));
    assign layer6_outputs[4034] = ~((layer5_outputs[1955]) & (layer5_outputs[896]));
    assign layer6_outputs[4035] = layer5_outputs[407];
    assign layer6_outputs[4036] = ~(layer5_outputs[1740]);
    assign layer6_outputs[4037] = layer5_outputs[4048];
    assign layer6_outputs[4038] = ~(layer5_outputs[2270]) | (layer5_outputs[5104]);
    assign layer6_outputs[4039] = 1'b1;
    assign layer6_outputs[4040] = layer5_outputs[2795];
    assign layer6_outputs[4041] = ~((layer5_outputs[3300]) ^ (layer5_outputs[3604]));
    assign layer6_outputs[4042] = ~((layer5_outputs[193]) | (layer5_outputs[1362]));
    assign layer6_outputs[4043] = ~(layer5_outputs[2211]);
    assign layer6_outputs[4044] = (layer5_outputs[2892]) & ~(layer5_outputs[5049]);
    assign layer6_outputs[4045] = (layer5_outputs[3616]) ^ (layer5_outputs[3161]);
    assign layer6_outputs[4046] = ~(layer5_outputs[3444]);
    assign layer6_outputs[4047] = ~(layer5_outputs[3421]) | (layer5_outputs[354]);
    assign layer6_outputs[4048] = ~(layer5_outputs[2268]);
    assign layer6_outputs[4049] = (layer5_outputs[1312]) & (layer5_outputs[733]);
    assign layer6_outputs[4050] = ~(layer5_outputs[572]);
    assign layer6_outputs[4051] = ~(layer5_outputs[4827]) | (layer5_outputs[187]);
    assign layer6_outputs[4052] = ~(layer5_outputs[918]) | (layer5_outputs[2784]);
    assign layer6_outputs[4053] = layer5_outputs[1826];
    assign layer6_outputs[4054] = ~(layer5_outputs[3107]);
    assign layer6_outputs[4055] = ~(layer5_outputs[4938]);
    assign layer6_outputs[4056] = ~((layer5_outputs[450]) & (layer5_outputs[4204]));
    assign layer6_outputs[4057] = layer5_outputs[3088];
    assign layer6_outputs[4058] = ~((layer5_outputs[2743]) ^ (layer5_outputs[3090]));
    assign layer6_outputs[4059] = layer5_outputs[1434];
    assign layer6_outputs[4060] = ~((layer5_outputs[2124]) ^ (layer5_outputs[3870]));
    assign layer6_outputs[4061] = (layer5_outputs[1977]) | (layer5_outputs[669]);
    assign layer6_outputs[4062] = ~(layer5_outputs[2294]);
    assign layer6_outputs[4063] = layer5_outputs[1684];
    assign layer6_outputs[4064] = ~(layer5_outputs[3992]);
    assign layer6_outputs[4065] = ~(layer5_outputs[2044]);
    assign layer6_outputs[4066] = ~(layer5_outputs[1461]);
    assign layer6_outputs[4067] = ~(layer5_outputs[3216]);
    assign layer6_outputs[4068] = ~(layer5_outputs[701]);
    assign layer6_outputs[4069] = ~(layer5_outputs[1866]);
    assign layer6_outputs[4070] = ~((layer5_outputs[2612]) | (layer5_outputs[3747]));
    assign layer6_outputs[4071] = layer5_outputs[3568];
    assign layer6_outputs[4072] = (layer5_outputs[1978]) ^ (layer5_outputs[2522]);
    assign layer6_outputs[4073] = ~((layer5_outputs[3908]) ^ (layer5_outputs[3946]));
    assign layer6_outputs[4074] = ~(layer5_outputs[2539]);
    assign layer6_outputs[4075] = (layer5_outputs[2921]) | (layer5_outputs[149]);
    assign layer6_outputs[4076] = (layer5_outputs[453]) & ~(layer5_outputs[186]);
    assign layer6_outputs[4077] = (layer5_outputs[2156]) & ~(layer5_outputs[43]);
    assign layer6_outputs[4078] = ~(layer5_outputs[3492]);
    assign layer6_outputs[4079] = ~((layer5_outputs[115]) | (layer5_outputs[5052]));
    assign layer6_outputs[4080] = ~(layer5_outputs[232]);
    assign layer6_outputs[4081] = ~(layer5_outputs[3348]);
    assign layer6_outputs[4082] = ~((layer5_outputs[3014]) ^ (layer5_outputs[3861]));
    assign layer6_outputs[4083] = layer5_outputs[4786];
    assign layer6_outputs[4084] = (layer5_outputs[903]) ^ (layer5_outputs[4983]);
    assign layer6_outputs[4085] = (layer5_outputs[2289]) & (layer5_outputs[4827]);
    assign layer6_outputs[4086] = ~(layer5_outputs[816]);
    assign layer6_outputs[4087] = (layer5_outputs[1021]) | (layer5_outputs[4446]);
    assign layer6_outputs[4088] = ~(layer5_outputs[355]);
    assign layer6_outputs[4089] = layer5_outputs[1304];
    assign layer6_outputs[4090] = ~(layer5_outputs[3395]);
    assign layer6_outputs[4091] = (layer5_outputs[2572]) | (layer5_outputs[3424]);
    assign layer6_outputs[4092] = ~(layer5_outputs[2365]);
    assign layer6_outputs[4093] = ~(layer5_outputs[4935]) | (layer5_outputs[318]);
    assign layer6_outputs[4094] = ~(layer5_outputs[1743]);
    assign layer6_outputs[4095] = layer5_outputs[3009];
    assign layer6_outputs[4096] = 1'b0;
    assign layer6_outputs[4097] = ~(layer5_outputs[315]);
    assign layer6_outputs[4098] = (layer5_outputs[2272]) & ~(layer5_outputs[3430]);
    assign layer6_outputs[4099] = ~((layer5_outputs[330]) ^ (layer5_outputs[3174]));
    assign layer6_outputs[4100] = layer5_outputs[2528];
    assign layer6_outputs[4101] = ~(layer5_outputs[2819]);
    assign layer6_outputs[4102] = layer5_outputs[2739];
    assign layer6_outputs[4103] = layer5_outputs[3182];
    assign layer6_outputs[4104] = ~((layer5_outputs[4240]) | (layer5_outputs[2540]));
    assign layer6_outputs[4105] = (layer5_outputs[2235]) & ~(layer5_outputs[222]);
    assign layer6_outputs[4106] = ~(layer5_outputs[3268]);
    assign layer6_outputs[4107] = ~(layer5_outputs[4620]);
    assign layer6_outputs[4108] = layer5_outputs[4198];
    assign layer6_outputs[4109] = (layer5_outputs[1737]) | (layer5_outputs[3298]);
    assign layer6_outputs[4110] = layer5_outputs[1682];
    assign layer6_outputs[4111] = (layer5_outputs[4550]) | (layer5_outputs[752]);
    assign layer6_outputs[4112] = ~((layer5_outputs[1718]) ^ (layer5_outputs[1736]));
    assign layer6_outputs[4113] = layer5_outputs[4157];
    assign layer6_outputs[4114] = ~(layer5_outputs[2731]);
    assign layer6_outputs[4115] = (layer5_outputs[153]) ^ (layer5_outputs[975]);
    assign layer6_outputs[4116] = 1'b1;
    assign layer6_outputs[4117] = ~(layer5_outputs[3884]);
    assign layer6_outputs[4118] = layer5_outputs[2286];
    assign layer6_outputs[4119] = layer5_outputs[4858];
    assign layer6_outputs[4120] = ~((layer5_outputs[2166]) & (layer5_outputs[420]));
    assign layer6_outputs[4121] = layer5_outputs[2441];
    assign layer6_outputs[4122] = layer5_outputs[4621];
    assign layer6_outputs[4123] = ~(layer5_outputs[2767]);
    assign layer6_outputs[4124] = layer5_outputs[1741];
    assign layer6_outputs[4125] = (layer5_outputs[4345]) | (layer5_outputs[4777]);
    assign layer6_outputs[4126] = layer5_outputs[1870];
    assign layer6_outputs[4127] = layer5_outputs[948];
    assign layer6_outputs[4128] = (layer5_outputs[1379]) & ~(layer5_outputs[2827]);
    assign layer6_outputs[4129] = layer5_outputs[4212];
    assign layer6_outputs[4130] = (layer5_outputs[2068]) & ~(layer5_outputs[4822]);
    assign layer6_outputs[4131] = layer5_outputs[3557];
    assign layer6_outputs[4132] = (layer5_outputs[503]) & ~(layer5_outputs[3496]);
    assign layer6_outputs[4133] = layer5_outputs[3892];
    assign layer6_outputs[4134] = layer5_outputs[1576];
    assign layer6_outputs[4135] = layer5_outputs[1098];
    assign layer6_outputs[4136] = layer5_outputs[4716];
    assign layer6_outputs[4137] = (layer5_outputs[2440]) ^ (layer5_outputs[173]);
    assign layer6_outputs[4138] = layer5_outputs[3231];
    assign layer6_outputs[4139] = 1'b0;
    assign layer6_outputs[4140] = ~((layer5_outputs[4661]) ^ (layer5_outputs[3488]));
    assign layer6_outputs[4141] = ~(layer5_outputs[1590]);
    assign layer6_outputs[4142] = (layer5_outputs[1208]) ^ (layer5_outputs[1483]);
    assign layer6_outputs[4143] = layer5_outputs[937];
    assign layer6_outputs[4144] = ~(layer5_outputs[5009]);
    assign layer6_outputs[4145] = (layer5_outputs[4491]) | (layer5_outputs[2167]);
    assign layer6_outputs[4146] = ~(layer5_outputs[3994]);
    assign layer6_outputs[4147] = (layer5_outputs[4442]) | (layer5_outputs[3764]);
    assign layer6_outputs[4148] = layer5_outputs[2430];
    assign layer6_outputs[4149] = (layer5_outputs[1890]) & ~(layer5_outputs[4511]);
    assign layer6_outputs[4150] = (layer5_outputs[2247]) ^ (layer5_outputs[2281]);
    assign layer6_outputs[4151] = 1'b0;
    assign layer6_outputs[4152] = ~((layer5_outputs[4393]) ^ (layer5_outputs[3258]));
    assign layer6_outputs[4153] = ~(layer5_outputs[1616]) | (layer5_outputs[3732]);
    assign layer6_outputs[4154] = ~(layer5_outputs[4001]);
    assign layer6_outputs[4155] = layer5_outputs[1420];
    assign layer6_outputs[4156] = layer5_outputs[644];
    assign layer6_outputs[4157] = layer5_outputs[3073];
    assign layer6_outputs[4158] = ~((layer5_outputs[6]) & (layer5_outputs[3572]));
    assign layer6_outputs[4159] = (layer5_outputs[3728]) ^ (layer5_outputs[1048]);
    assign layer6_outputs[4160] = (layer5_outputs[4249]) & ~(layer5_outputs[3865]);
    assign layer6_outputs[4161] = ~(layer5_outputs[3894]);
    assign layer6_outputs[4162] = layer5_outputs[4917];
    assign layer6_outputs[4163] = ~((layer5_outputs[2414]) & (layer5_outputs[238]));
    assign layer6_outputs[4164] = ~(layer5_outputs[3330]) | (layer5_outputs[914]);
    assign layer6_outputs[4165] = ~(layer5_outputs[564]) | (layer5_outputs[1495]);
    assign layer6_outputs[4166] = ~(layer5_outputs[1951]) | (layer5_outputs[2376]);
    assign layer6_outputs[4167] = layer5_outputs[1382];
    assign layer6_outputs[4168] = ~(layer5_outputs[1013]) | (layer5_outputs[292]);
    assign layer6_outputs[4169] = (layer5_outputs[3342]) & ~(layer5_outputs[4361]);
    assign layer6_outputs[4170] = ~((layer5_outputs[2251]) ^ (layer5_outputs[3015]));
    assign layer6_outputs[4171] = ~(layer5_outputs[194]);
    assign layer6_outputs[4172] = layer5_outputs[3123];
    assign layer6_outputs[4173] = 1'b0;
    assign layer6_outputs[4174] = layer5_outputs[4752];
    assign layer6_outputs[4175] = ~(layer5_outputs[3890]) | (layer5_outputs[896]);
    assign layer6_outputs[4176] = ~(layer5_outputs[4713]);
    assign layer6_outputs[4177] = (layer5_outputs[374]) | (layer5_outputs[93]);
    assign layer6_outputs[4178] = layer5_outputs[3178];
    assign layer6_outputs[4179] = layer5_outputs[4289];
    assign layer6_outputs[4180] = layer5_outputs[4323];
    assign layer6_outputs[4181] = layer5_outputs[1835];
    assign layer6_outputs[4182] = ~((layer5_outputs[1210]) | (layer5_outputs[2711]));
    assign layer6_outputs[4183] = layer5_outputs[2620];
    assign layer6_outputs[4184] = layer5_outputs[4369];
    assign layer6_outputs[4185] = ~(layer5_outputs[5086]);
    assign layer6_outputs[4186] = layer5_outputs[926];
    assign layer6_outputs[4187] = layer5_outputs[179];
    assign layer6_outputs[4188] = layer5_outputs[1939];
    assign layer6_outputs[4189] = ~((layer5_outputs[14]) ^ (layer5_outputs[238]));
    assign layer6_outputs[4190] = ~((layer5_outputs[1080]) ^ (layer5_outputs[4700]));
    assign layer6_outputs[4191] = layer5_outputs[2426];
    assign layer6_outputs[4192] = ~((layer5_outputs[3702]) & (layer5_outputs[84]));
    assign layer6_outputs[4193] = layer5_outputs[5063];
    assign layer6_outputs[4194] = ~((layer5_outputs[1264]) | (layer5_outputs[3706]));
    assign layer6_outputs[4195] = ~((layer5_outputs[2172]) ^ (layer5_outputs[1117]));
    assign layer6_outputs[4196] = (layer5_outputs[3738]) & ~(layer5_outputs[4355]);
    assign layer6_outputs[4197] = ~((layer5_outputs[4561]) ^ (layer5_outputs[2225]));
    assign layer6_outputs[4198] = ~(layer5_outputs[911]) | (layer5_outputs[351]);
    assign layer6_outputs[4199] = layer5_outputs[3258];
    assign layer6_outputs[4200] = layer5_outputs[2049];
    assign layer6_outputs[4201] = ~((layer5_outputs[269]) & (layer5_outputs[1306]));
    assign layer6_outputs[4202] = ~(layer5_outputs[3505]) | (layer5_outputs[668]);
    assign layer6_outputs[4203] = ~(layer5_outputs[3060]);
    assign layer6_outputs[4204] = 1'b0;
    assign layer6_outputs[4205] = layer5_outputs[1471];
    assign layer6_outputs[4206] = (layer5_outputs[4973]) ^ (layer5_outputs[5080]);
    assign layer6_outputs[4207] = ~(layer5_outputs[4690]);
    assign layer6_outputs[4208] = 1'b0;
    assign layer6_outputs[4209] = layer5_outputs[1610];
    assign layer6_outputs[4210] = (layer5_outputs[2427]) & (layer5_outputs[134]);
    assign layer6_outputs[4211] = (layer5_outputs[4644]) & (layer5_outputs[1377]);
    assign layer6_outputs[4212] = ~(layer5_outputs[3968]);
    assign layer6_outputs[4213] = (layer5_outputs[4317]) | (layer5_outputs[1011]);
    assign layer6_outputs[4214] = ~(layer5_outputs[3953]);
    assign layer6_outputs[4215] = ~((layer5_outputs[3896]) ^ (layer5_outputs[252]));
    assign layer6_outputs[4216] = (layer5_outputs[3354]) & ~(layer5_outputs[4350]);
    assign layer6_outputs[4217] = ~(layer5_outputs[4473]) | (layer5_outputs[3358]);
    assign layer6_outputs[4218] = layer5_outputs[2988];
    assign layer6_outputs[4219] = ~(layer5_outputs[3971]);
    assign layer6_outputs[4220] = (layer5_outputs[4380]) & ~(layer5_outputs[4557]);
    assign layer6_outputs[4221] = (layer5_outputs[2095]) ^ (layer5_outputs[1541]);
    assign layer6_outputs[4222] = layer5_outputs[3289];
    assign layer6_outputs[4223] = layer5_outputs[425];
    assign layer6_outputs[4224] = ~((layer5_outputs[3910]) & (layer5_outputs[5040]));
    assign layer6_outputs[4225] = ~(layer5_outputs[197]);
    assign layer6_outputs[4226] = (layer5_outputs[4224]) | (layer5_outputs[3606]);
    assign layer6_outputs[4227] = (layer5_outputs[588]) ^ (layer5_outputs[1848]);
    assign layer6_outputs[4228] = (layer5_outputs[2001]) & ~(layer5_outputs[1500]);
    assign layer6_outputs[4229] = layer5_outputs[5092];
    assign layer6_outputs[4230] = layer5_outputs[3132];
    assign layer6_outputs[4231] = ~(layer5_outputs[3449]);
    assign layer6_outputs[4232] = ~(layer5_outputs[4780]);
    assign layer6_outputs[4233] = ~(layer5_outputs[928]) | (layer5_outputs[2924]);
    assign layer6_outputs[4234] = ~(layer5_outputs[5048]);
    assign layer6_outputs[4235] = layer5_outputs[480];
    assign layer6_outputs[4236] = layer5_outputs[601];
    assign layer6_outputs[4237] = ~(layer5_outputs[1677]) | (layer5_outputs[4691]);
    assign layer6_outputs[4238] = ~((layer5_outputs[1241]) | (layer5_outputs[4944]));
    assign layer6_outputs[4239] = layer5_outputs[4145];
    assign layer6_outputs[4240] = ~(layer5_outputs[3837]) | (layer5_outputs[653]);
    assign layer6_outputs[4241] = ~((layer5_outputs[112]) | (layer5_outputs[88]));
    assign layer6_outputs[4242] = layer5_outputs[4358];
    assign layer6_outputs[4243] = ~(layer5_outputs[2370]);
    assign layer6_outputs[4244] = ~(layer5_outputs[1877]);
    assign layer6_outputs[4245] = ~(layer5_outputs[4456]);
    assign layer6_outputs[4246] = ~(layer5_outputs[992]);
    assign layer6_outputs[4247] = (layer5_outputs[1950]) & ~(layer5_outputs[474]);
    assign layer6_outputs[4248] = layer5_outputs[4413];
    assign layer6_outputs[4249] = ~((layer5_outputs[2604]) | (layer5_outputs[1969]));
    assign layer6_outputs[4250] = 1'b0;
    assign layer6_outputs[4251] = layer5_outputs[726];
    assign layer6_outputs[4252] = layer5_outputs[3418];
    assign layer6_outputs[4253] = ~(layer5_outputs[143]);
    assign layer6_outputs[4254] = (layer5_outputs[3477]) & ~(layer5_outputs[3796]);
    assign layer6_outputs[4255] = ~((layer5_outputs[3062]) ^ (layer5_outputs[1460]));
    assign layer6_outputs[4256] = (layer5_outputs[409]) ^ (layer5_outputs[1860]);
    assign layer6_outputs[4257] = ~(layer5_outputs[3352]) | (layer5_outputs[2684]);
    assign layer6_outputs[4258] = ~((layer5_outputs[2363]) & (layer5_outputs[286]));
    assign layer6_outputs[4259] = ~((layer5_outputs[2248]) ^ (layer5_outputs[2277]));
    assign layer6_outputs[4260] = (layer5_outputs[1319]) | (layer5_outputs[1395]);
    assign layer6_outputs[4261] = ~(layer5_outputs[2695]) | (layer5_outputs[74]);
    assign layer6_outputs[4262] = (layer5_outputs[1377]) & (layer5_outputs[1250]);
    assign layer6_outputs[4263] = ~(layer5_outputs[860]);
    assign layer6_outputs[4264] = layer5_outputs[4697];
    assign layer6_outputs[4265] = ~((layer5_outputs[411]) ^ (layer5_outputs[590]));
    assign layer6_outputs[4266] = layer5_outputs[4064];
    assign layer6_outputs[4267] = layer5_outputs[1551];
    assign layer6_outputs[4268] = layer5_outputs[1358];
    assign layer6_outputs[4269] = (layer5_outputs[431]) & ~(layer5_outputs[4154]);
    assign layer6_outputs[4270] = ~(layer5_outputs[358]);
    assign layer6_outputs[4271] = layer5_outputs[4648];
    assign layer6_outputs[4272] = layer5_outputs[2601];
    assign layer6_outputs[4273] = ~((layer5_outputs[130]) | (layer5_outputs[3427]));
    assign layer6_outputs[4274] = (layer5_outputs[4604]) ^ (layer5_outputs[221]);
    assign layer6_outputs[4275] = ~((layer5_outputs[3731]) | (layer5_outputs[1905]));
    assign layer6_outputs[4276] = ~(layer5_outputs[1976]);
    assign layer6_outputs[4277] = layer5_outputs[2529];
    assign layer6_outputs[4278] = 1'b1;
    assign layer6_outputs[4279] = ~((layer5_outputs[4615]) ^ (layer5_outputs[3423]));
    assign layer6_outputs[4280] = ~(layer5_outputs[4307]);
    assign layer6_outputs[4281] = layer5_outputs[3172];
    assign layer6_outputs[4282] = ~(layer5_outputs[258]);
    assign layer6_outputs[4283] = ~((layer5_outputs[2838]) ^ (layer5_outputs[2017]));
    assign layer6_outputs[4284] = ~(layer5_outputs[463]);
    assign layer6_outputs[4285] = layer5_outputs[2750];
    assign layer6_outputs[4286] = ~(layer5_outputs[3809]) | (layer5_outputs[2862]);
    assign layer6_outputs[4287] = ~(layer5_outputs[2203]) | (layer5_outputs[421]);
    assign layer6_outputs[4288] = ~(layer5_outputs[3914]);
    assign layer6_outputs[4289] = ~((layer5_outputs[2462]) & (layer5_outputs[1388]));
    assign layer6_outputs[4290] = layer5_outputs[2254];
    assign layer6_outputs[4291] = (layer5_outputs[4930]) & ~(layer5_outputs[1324]);
    assign layer6_outputs[4292] = ~((layer5_outputs[1169]) | (layer5_outputs[2341]));
    assign layer6_outputs[4293] = ~(layer5_outputs[2619]) | (layer5_outputs[1876]);
    assign layer6_outputs[4294] = ~(layer5_outputs[2719]);
    assign layer6_outputs[4295] = ~(layer5_outputs[2849]) | (layer5_outputs[2971]);
    assign layer6_outputs[4296] = layer5_outputs[165];
    assign layer6_outputs[4297] = layer5_outputs[3621];
    assign layer6_outputs[4298] = ~((layer5_outputs[4528]) ^ (layer5_outputs[2895]));
    assign layer6_outputs[4299] = layer5_outputs[2536];
    assign layer6_outputs[4300] = ~(layer5_outputs[4879]) | (layer5_outputs[1913]);
    assign layer6_outputs[4301] = (layer5_outputs[4445]) & ~(layer5_outputs[364]);
    assign layer6_outputs[4302] = layer5_outputs[4492];
    assign layer6_outputs[4303] = 1'b0;
    assign layer6_outputs[4304] = 1'b0;
    assign layer6_outputs[4305] = ~((layer5_outputs[4732]) & (layer5_outputs[71]));
    assign layer6_outputs[4306] = ~(layer5_outputs[636]);
    assign layer6_outputs[4307] = ~(layer5_outputs[4976]) | (layer5_outputs[3957]);
    assign layer6_outputs[4308] = ~(layer5_outputs[1831]);
    assign layer6_outputs[4309] = ~((layer5_outputs[2252]) & (layer5_outputs[1355]));
    assign layer6_outputs[4310] = 1'b0;
    assign layer6_outputs[4311] = ~((layer5_outputs[2108]) ^ (layer5_outputs[4279]));
    assign layer6_outputs[4312] = layer5_outputs[4457];
    assign layer6_outputs[4313] = layer5_outputs[4467];
    assign layer6_outputs[4314] = ~(layer5_outputs[5002]);
    assign layer6_outputs[4315] = layer5_outputs[3404];
    assign layer6_outputs[4316] = layer5_outputs[2447];
    assign layer6_outputs[4317] = layer5_outputs[3779];
    assign layer6_outputs[4318] = (layer5_outputs[212]) | (layer5_outputs[1328]);
    assign layer6_outputs[4319] = ~(layer5_outputs[3766]);
    assign layer6_outputs[4320] = ~((layer5_outputs[5094]) | (layer5_outputs[378]));
    assign layer6_outputs[4321] = layer5_outputs[4838];
    assign layer6_outputs[4322] = layer5_outputs[2214];
    assign layer6_outputs[4323] = ~(layer5_outputs[3703]);
    assign layer6_outputs[4324] = layer5_outputs[3570];
    assign layer6_outputs[4325] = layer5_outputs[2195];
    assign layer6_outputs[4326] = ~(layer5_outputs[919]);
    assign layer6_outputs[4327] = layer5_outputs[2586];
    assign layer6_outputs[4328] = ~((layer5_outputs[650]) ^ (layer5_outputs[2346]));
    assign layer6_outputs[4329] = layer5_outputs[3039];
    assign layer6_outputs[4330] = ~(layer5_outputs[2965]);
    assign layer6_outputs[4331] = ~(layer5_outputs[3426]);
    assign layer6_outputs[4332] = ~((layer5_outputs[651]) & (layer5_outputs[1749]));
    assign layer6_outputs[4333] = layer5_outputs[1927];
    assign layer6_outputs[4334] = (layer5_outputs[4714]) & ~(layer5_outputs[2662]);
    assign layer6_outputs[4335] = ~(layer5_outputs[4380]);
    assign layer6_outputs[4336] = ~(layer5_outputs[1907]);
    assign layer6_outputs[4337] = ~(layer5_outputs[3084]);
    assign layer6_outputs[4338] = ~((layer5_outputs[4785]) | (layer5_outputs[4798]));
    assign layer6_outputs[4339] = layer5_outputs[2736];
    assign layer6_outputs[4340] = layer5_outputs[11];
    assign layer6_outputs[4341] = ~(layer5_outputs[2392]);
    assign layer6_outputs[4342] = (layer5_outputs[758]) & (layer5_outputs[965]);
    assign layer6_outputs[4343] = ~(layer5_outputs[1207]);
    assign layer6_outputs[4344] = (layer5_outputs[627]) | (layer5_outputs[74]);
    assign layer6_outputs[4345] = ~(layer5_outputs[2838]) | (layer5_outputs[2648]);
    assign layer6_outputs[4346] = layer5_outputs[961];
    assign layer6_outputs[4347] = ~(layer5_outputs[700]) | (layer5_outputs[4834]);
    assign layer6_outputs[4348] = layer5_outputs[1346];
    assign layer6_outputs[4349] = (layer5_outputs[62]) & (layer5_outputs[4421]);
    assign layer6_outputs[4350] = ~(layer5_outputs[3667]) | (layer5_outputs[3037]);
    assign layer6_outputs[4351] = ~(layer5_outputs[4808]);
    assign layer6_outputs[4352] = layer5_outputs[1460];
    assign layer6_outputs[4353] = (layer5_outputs[4215]) & (layer5_outputs[294]);
    assign layer6_outputs[4354] = 1'b1;
    assign layer6_outputs[4355] = layer5_outputs[1439];
    assign layer6_outputs[4356] = ~(layer5_outputs[1542]);
    assign layer6_outputs[4357] = ~(layer5_outputs[363]);
    assign layer6_outputs[4358] = ~(layer5_outputs[570]) | (layer5_outputs[3524]);
    assign layer6_outputs[4359] = (layer5_outputs[354]) & (layer5_outputs[2739]);
    assign layer6_outputs[4360] = ~(layer5_outputs[4959]);
    assign layer6_outputs[4361] = (layer5_outputs[3103]) & ~(layer5_outputs[1047]);
    assign layer6_outputs[4362] = ~((layer5_outputs[262]) ^ (layer5_outputs[1814]));
    assign layer6_outputs[4363] = ~(layer5_outputs[3053]) | (layer5_outputs[977]);
    assign layer6_outputs[4364] = ~(layer5_outputs[484]) | (layer5_outputs[308]);
    assign layer6_outputs[4365] = ~(layer5_outputs[1842]) | (layer5_outputs[2416]);
    assign layer6_outputs[4366] = layer5_outputs[4140];
    assign layer6_outputs[4367] = (layer5_outputs[4669]) | (layer5_outputs[3689]);
    assign layer6_outputs[4368] = layer5_outputs[4685];
    assign layer6_outputs[4369] = layer5_outputs[1792];
    assign layer6_outputs[4370] = layer5_outputs[2354];
    assign layer6_outputs[4371] = layer5_outputs[4491];
    assign layer6_outputs[4372] = ~((layer5_outputs[339]) ^ (layer5_outputs[2821]));
    assign layer6_outputs[4373] = ~(layer5_outputs[2601]) | (layer5_outputs[2593]);
    assign layer6_outputs[4374] = ~(layer5_outputs[3125]) | (layer5_outputs[4418]);
    assign layer6_outputs[4375] = (layer5_outputs[3900]) ^ (layer5_outputs[1035]);
    assign layer6_outputs[4376] = ~(layer5_outputs[2129]) | (layer5_outputs[4159]);
    assign layer6_outputs[4377] = ~(layer5_outputs[3273]);
    assign layer6_outputs[4378] = (layer5_outputs[2465]) & ~(layer5_outputs[1876]);
    assign layer6_outputs[4379] = ~((layer5_outputs[1381]) & (layer5_outputs[1929]));
    assign layer6_outputs[4380] = (layer5_outputs[2364]) & ~(layer5_outputs[2493]);
    assign layer6_outputs[4381] = layer5_outputs[2636];
    assign layer6_outputs[4382] = ~(layer5_outputs[2283]) | (layer5_outputs[2487]);
    assign layer6_outputs[4383] = (layer5_outputs[582]) ^ (layer5_outputs[3820]);
    assign layer6_outputs[4384] = (layer5_outputs[534]) ^ (layer5_outputs[2408]);
    assign layer6_outputs[4385] = layer5_outputs[1257];
    assign layer6_outputs[4386] = (layer5_outputs[365]) | (layer5_outputs[4596]);
    assign layer6_outputs[4387] = layer5_outputs[4015];
    assign layer6_outputs[4388] = ~((layer5_outputs[4128]) | (layer5_outputs[2907]));
    assign layer6_outputs[4389] = (layer5_outputs[4002]) & ~(layer5_outputs[3059]);
    assign layer6_outputs[4390] = ~(layer5_outputs[322]) | (layer5_outputs[1203]);
    assign layer6_outputs[4391] = layer5_outputs[2216];
    assign layer6_outputs[4392] = (layer5_outputs[807]) & (layer5_outputs[1613]);
    assign layer6_outputs[4393] = (layer5_outputs[4205]) | (layer5_outputs[1820]);
    assign layer6_outputs[4394] = (layer5_outputs[1871]) | (layer5_outputs[85]);
    assign layer6_outputs[4395] = layer5_outputs[963];
    assign layer6_outputs[4396] = layer5_outputs[381];
    assign layer6_outputs[4397] = ~((layer5_outputs[3565]) ^ (layer5_outputs[5004]));
    assign layer6_outputs[4398] = layer5_outputs[4049];
    assign layer6_outputs[4399] = layer5_outputs[2372];
    assign layer6_outputs[4400] = (layer5_outputs[4481]) ^ (layer5_outputs[735]);
    assign layer6_outputs[4401] = layer5_outputs[3296];
    assign layer6_outputs[4402] = ~((layer5_outputs[3883]) & (layer5_outputs[2332]));
    assign layer6_outputs[4403] = ~(layer5_outputs[2635]);
    assign layer6_outputs[4404] = ~(layer5_outputs[1763]) | (layer5_outputs[3313]);
    assign layer6_outputs[4405] = layer5_outputs[4501];
    assign layer6_outputs[4406] = (layer5_outputs[3339]) | (layer5_outputs[3069]);
    assign layer6_outputs[4407] = layer5_outputs[910];
    assign layer6_outputs[4408] = layer5_outputs[2492];
    assign layer6_outputs[4409] = 1'b1;
    assign layer6_outputs[4410] = layer5_outputs[2470];
    assign layer6_outputs[4411] = layer5_outputs[4566];
    assign layer6_outputs[4412] = ~((layer5_outputs[1368]) ^ (layer5_outputs[637]));
    assign layer6_outputs[4413] = ~(layer5_outputs[3766]);
    assign layer6_outputs[4414] = layer5_outputs[2242];
    assign layer6_outputs[4415] = (layer5_outputs[1755]) ^ (layer5_outputs[3271]);
    assign layer6_outputs[4416] = layer5_outputs[4569];
    assign layer6_outputs[4417] = layer5_outputs[1086];
    assign layer6_outputs[4418] = ~((layer5_outputs[1999]) | (layer5_outputs[3867]));
    assign layer6_outputs[4419] = ~(layer5_outputs[4238]);
    assign layer6_outputs[4420] = ~(layer5_outputs[3776]) | (layer5_outputs[3608]);
    assign layer6_outputs[4421] = ~((layer5_outputs[4902]) & (layer5_outputs[1992]));
    assign layer6_outputs[4422] = layer5_outputs[3797];
    assign layer6_outputs[4423] = 1'b0;
    assign layer6_outputs[4424] = (layer5_outputs[4006]) & (layer5_outputs[3638]);
    assign layer6_outputs[4425] = layer5_outputs[4266];
    assign layer6_outputs[4426] = ~(layer5_outputs[2410]);
    assign layer6_outputs[4427] = ~(layer5_outputs[1975]) | (layer5_outputs[4337]);
    assign layer6_outputs[4428] = (layer5_outputs[4936]) & ~(layer5_outputs[197]);
    assign layer6_outputs[4429] = (layer5_outputs[2909]) & ~(layer5_outputs[837]);
    assign layer6_outputs[4430] = ~(layer5_outputs[351]);
    assign layer6_outputs[4431] = ~(layer5_outputs[4232]) | (layer5_outputs[256]);
    assign layer6_outputs[4432] = ~(layer5_outputs[3150]);
    assign layer6_outputs[4433] = (layer5_outputs[3954]) & ~(layer5_outputs[3843]);
    assign layer6_outputs[4434] = (layer5_outputs[1111]) & ~(layer5_outputs[4803]);
    assign layer6_outputs[4435] = ~(layer5_outputs[1205]);
    assign layer6_outputs[4436] = (layer5_outputs[5095]) | (layer5_outputs[986]);
    assign layer6_outputs[4437] = ~(layer5_outputs[1821]);
    assign layer6_outputs[4438] = ~(layer5_outputs[3016]) | (layer5_outputs[1071]);
    assign layer6_outputs[4439] = ~((layer5_outputs[5108]) | (layer5_outputs[679]));
    assign layer6_outputs[4440] = ~((layer5_outputs[3139]) ^ (layer5_outputs[1732]));
    assign layer6_outputs[4441] = ~((layer5_outputs[1637]) ^ (layer5_outputs[1679]));
    assign layer6_outputs[4442] = ~(layer5_outputs[2262]);
    assign layer6_outputs[4443] = ~(layer5_outputs[2315]);
    assign layer6_outputs[4444] = layer5_outputs[2042];
    assign layer6_outputs[4445] = layer5_outputs[3024];
    assign layer6_outputs[4446] = layer5_outputs[3048];
    assign layer6_outputs[4447] = (layer5_outputs[517]) | (layer5_outputs[3108]);
    assign layer6_outputs[4448] = layer5_outputs[34];
    assign layer6_outputs[4449] = ~(layer5_outputs[49]);
    assign layer6_outputs[4450] = (layer5_outputs[1225]) | (layer5_outputs[4710]);
    assign layer6_outputs[4451] = ~(layer5_outputs[487]);
    assign layer6_outputs[4452] = (layer5_outputs[2944]) | (layer5_outputs[2955]);
    assign layer6_outputs[4453] = layer5_outputs[2377];
    assign layer6_outputs[4454] = ~(layer5_outputs[4489]);
    assign layer6_outputs[4455] = ~((layer5_outputs[3940]) & (layer5_outputs[616]));
    assign layer6_outputs[4456] = layer5_outputs[1443];
    assign layer6_outputs[4457] = (layer5_outputs[183]) ^ (layer5_outputs[4649]);
    assign layer6_outputs[4458] = (layer5_outputs[347]) | (layer5_outputs[456]);
    assign layer6_outputs[4459] = ~(layer5_outputs[1987]);
    assign layer6_outputs[4460] = ~(layer5_outputs[293]);
    assign layer6_outputs[4461] = (layer5_outputs[2455]) & ~(layer5_outputs[3145]);
    assign layer6_outputs[4462] = ~(layer5_outputs[2765]);
    assign layer6_outputs[4463] = ~((layer5_outputs[4041]) ^ (layer5_outputs[3044]));
    assign layer6_outputs[4464] = layer5_outputs[1600];
    assign layer6_outputs[4465] = layer5_outputs[2020];
    assign layer6_outputs[4466] = layer5_outputs[673];
    assign layer6_outputs[4467] = layer5_outputs[4907];
    assign layer6_outputs[4468] = ~(layer5_outputs[85]);
    assign layer6_outputs[4469] = ~(layer5_outputs[4336]);
    assign layer6_outputs[4470] = layer5_outputs[2210];
    assign layer6_outputs[4471] = (layer5_outputs[171]) & ~(layer5_outputs[5093]);
    assign layer6_outputs[4472] = ~(layer5_outputs[3953]) | (layer5_outputs[2306]);
    assign layer6_outputs[4473] = ~((layer5_outputs[4204]) ^ (layer5_outputs[3756]));
    assign layer6_outputs[4474] = layer5_outputs[4714];
    assign layer6_outputs[4475] = (layer5_outputs[3679]) ^ (layer5_outputs[3188]);
    assign layer6_outputs[4476] = ~(layer5_outputs[3347]);
    assign layer6_outputs[4477] = ~(layer5_outputs[501]);
    assign layer6_outputs[4478] = (layer5_outputs[3861]) & ~(layer5_outputs[2719]);
    assign layer6_outputs[4479] = ~(layer5_outputs[4197]);
    assign layer6_outputs[4480] = ~(layer5_outputs[4207]);
    assign layer6_outputs[4481] = layer5_outputs[3398];
    assign layer6_outputs[4482] = (layer5_outputs[3413]) & ~(layer5_outputs[638]);
    assign layer6_outputs[4483] = ~((layer5_outputs[1774]) & (layer5_outputs[1135]));
    assign layer6_outputs[4484] = ~(layer5_outputs[58]) | (layer5_outputs[1192]);
    assign layer6_outputs[4485] = layer5_outputs[3836];
    assign layer6_outputs[4486] = ~(layer5_outputs[2083]) | (layer5_outputs[3504]);
    assign layer6_outputs[4487] = ~(layer5_outputs[4016]) | (layer5_outputs[10]);
    assign layer6_outputs[4488] = ~((layer5_outputs[3289]) ^ (layer5_outputs[3903]));
    assign layer6_outputs[4489] = layer5_outputs[3901];
    assign layer6_outputs[4490] = ~(layer5_outputs[3936]);
    assign layer6_outputs[4491] = layer5_outputs[5118];
    assign layer6_outputs[4492] = (layer5_outputs[4584]) & (layer5_outputs[1360]);
    assign layer6_outputs[4493] = ~(layer5_outputs[3694]);
    assign layer6_outputs[4494] = ~(layer5_outputs[2505]);
    assign layer6_outputs[4495] = layer5_outputs[4285];
    assign layer6_outputs[4496] = ~(layer5_outputs[4946]);
    assign layer6_outputs[4497] = ~(layer5_outputs[2610]);
    assign layer6_outputs[4498] = ~(layer5_outputs[3385]);
    assign layer6_outputs[4499] = (layer5_outputs[4494]) & ~(layer5_outputs[959]);
    assign layer6_outputs[4500] = ~(layer5_outputs[4151]);
    assign layer6_outputs[4501] = layer5_outputs[3868];
    assign layer6_outputs[4502] = ~(layer5_outputs[3923]);
    assign layer6_outputs[4503] = ~(layer5_outputs[3261]);
    assign layer6_outputs[4504] = ~(layer5_outputs[1949]);
    assign layer6_outputs[4505] = (layer5_outputs[4136]) & ~(layer5_outputs[715]);
    assign layer6_outputs[4506] = (layer5_outputs[4392]) & (layer5_outputs[1592]);
    assign layer6_outputs[4507] = ~((layer5_outputs[1816]) ^ (layer5_outputs[2932]));
    assign layer6_outputs[4508] = ~(layer5_outputs[2643]);
    assign layer6_outputs[4509] = ~((layer5_outputs[4739]) ^ (layer5_outputs[229]));
    assign layer6_outputs[4510] = layer5_outputs[4854];
    assign layer6_outputs[4511] = ~((layer5_outputs[4429]) | (layer5_outputs[4955]));
    assign layer6_outputs[4512] = layer5_outputs[3172];
    assign layer6_outputs[4513] = ~(layer5_outputs[203]);
    assign layer6_outputs[4514] = (layer5_outputs[2640]) & ~(layer5_outputs[3303]);
    assign layer6_outputs[4515] = ~((layer5_outputs[1689]) ^ (layer5_outputs[4269]));
    assign layer6_outputs[4516] = ~(layer5_outputs[2858]);
    assign layer6_outputs[4517] = ~(layer5_outputs[3876]);
    assign layer6_outputs[4518] = ~(layer5_outputs[4785]) | (layer5_outputs[4399]);
    assign layer6_outputs[4519] = ~(layer5_outputs[1364]);
    assign layer6_outputs[4520] = ~(layer5_outputs[2513]);
    assign layer6_outputs[4521] = ~(layer5_outputs[4497]);
    assign layer6_outputs[4522] = ~(layer5_outputs[1394]);
    assign layer6_outputs[4523] = (layer5_outputs[511]) & ~(layer5_outputs[4247]);
    assign layer6_outputs[4524] = layer5_outputs[705];
    assign layer6_outputs[4525] = ~(layer5_outputs[4764]) | (layer5_outputs[2008]);
    assign layer6_outputs[4526] = layer5_outputs[4351];
    assign layer6_outputs[4527] = layer5_outputs[2841];
    assign layer6_outputs[4528] = layer5_outputs[3255];
    assign layer6_outputs[4529] = (layer5_outputs[958]) & ~(layer5_outputs[4621]);
    assign layer6_outputs[4530] = ~(layer5_outputs[3403]);
    assign layer6_outputs[4531] = layer5_outputs[593];
    assign layer6_outputs[4532] = ~(layer5_outputs[3765]) | (layer5_outputs[4357]);
    assign layer6_outputs[4533] = ~(layer5_outputs[3640]) | (layer5_outputs[3558]);
    assign layer6_outputs[4534] = ~(layer5_outputs[2646]) | (layer5_outputs[3525]);
    assign layer6_outputs[4535] = (layer5_outputs[640]) ^ (layer5_outputs[618]);
    assign layer6_outputs[4536] = ~(layer5_outputs[1105]);
    assign layer6_outputs[4537] = ~((layer5_outputs[1402]) | (layer5_outputs[4993]));
    assign layer6_outputs[4538] = (layer5_outputs[458]) ^ (layer5_outputs[213]);
    assign layer6_outputs[4539] = ~(layer5_outputs[4898]);
    assign layer6_outputs[4540] = (layer5_outputs[984]) & ~(layer5_outputs[4025]);
    assign layer6_outputs[4541] = ~((layer5_outputs[1184]) ^ (layer5_outputs[861]));
    assign layer6_outputs[4542] = (layer5_outputs[4560]) & (layer5_outputs[3944]);
    assign layer6_outputs[4543] = (layer5_outputs[1127]) & (layer5_outputs[1758]);
    assign layer6_outputs[4544] = ~(layer5_outputs[2802]);
    assign layer6_outputs[4545] = layer5_outputs[1357];
    assign layer6_outputs[4546] = ~(layer5_outputs[3767]);
    assign layer6_outputs[4547] = (layer5_outputs[2504]) ^ (layer5_outputs[1665]);
    assign layer6_outputs[4548] = ~(layer5_outputs[2166]);
    assign layer6_outputs[4549] = (layer5_outputs[2312]) ^ (layer5_outputs[1284]);
    assign layer6_outputs[4550] = ~((layer5_outputs[3129]) & (layer5_outputs[4911]));
    assign layer6_outputs[4551] = (layer5_outputs[4653]) | (layer5_outputs[4833]);
    assign layer6_outputs[4552] = ~(layer5_outputs[5036]);
    assign layer6_outputs[4553] = (layer5_outputs[3457]) ^ (layer5_outputs[330]);
    assign layer6_outputs[4554] = layer5_outputs[5099];
    assign layer6_outputs[4555] = layer5_outputs[1302];
    assign layer6_outputs[4556] = ~(layer5_outputs[2737]) | (layer5_outputs[3430]);
    assign layer6_outputs[4557] = ~(layer5_outputs[1298]);
    assign layer6_outputs[4558] = (layer5_outputs[281]) | (layer5_outputs[1130]);
    assign layer6_outputs[4559] = 1'b0;
    assign layer6_outputs[4560] = ~(layer5_outputs[3995]) | (layer5_outputs[3217]);
    assign layer6_outputs[4561] = (layer5_outputs[1853]) ^ (layer5_outputs[2016]);
    assign layer6_outputs[4562] = (layer5_outputs[2908]) & ~(layer5_outputs[942]);
    assign layer6_outputs[4563] = ~((layer5_outputs[4894]) & (layer5_outputs[1764]));
    assign layer6_outputs[4564] = layer5_outputs[293];
    assign layer6_outputs[4565] = ~((layer5_outputs[1434]) | (layer5_outputs[461]));
    assign layer6_outputs[4566] = layer5_outputs[3996];
    assign layer6_outputs[4567] = ~((layer5_outputs[4108]) ^ (layer5_outputs[3023]));
    assign layer6_outputs[4568] = layer5_outputs[3294];
    assign layer6_outputs[4569] = ~(layer5_outputs[94]);
    assign layer6_outputs[4570] = ~((layer5_outputs[564]) & (layer5_outputs[4069]));
    assign layer6_outputs[4571] = ~(layer5_outputs[356]);
    assign layer6_outputs[4572] = (layer5_outputs[3859]) & ~(layer5_outputs[2396]);
    assign layer6_outputs[4573] = layer5_outputs[403];
    assign layer6_outputs[4574] = (layer5_outputs[2542]) ^ (layer5_outputs[4607]);
    assign layer6_outputs[4575] = ~(layer5_outputs[3948]);
    assign layer6_outputs[4576] = layer5_outputs[3585];
    assign layer6_outputs[4577] = layer5_outputs[2263];
    assign layer6_outputs[4578] = ~((layer5_outputs[1887]) | (layer5_outputs[1915]));
    assign layer6_outputs[4579] = layer5_outputs[2007];
    assign layer6_outputs[4580] = ~(layer5_outputs[1602]);
    assign layer6_outputs[4581] = layer5_outputs[1201];
    assign layer6_outputs[4582] = (layer5_outputs[56]) & (layer5_outputs[759]);
    assign layer6_outputs[4583] = ~(layer5_outputs[4617]);
    assign layer6_outputs[4584] = layer5_outputs[2618];
    assign layer6_outputs[4585] = ~((layer5_outputs[3412]) & (layer5_outputs[1211]));
    assign layer6_outputs[4586] = ~(layer5_outputs[3366]);
    assign layer6_outputs[4587] = layer5_outputs[2831];
    assign layer6_outputs[4588] = layer5_outputs[831];
    assign layer6_outputs[4589] = (layer5_outputs[1157]) & (layer5_outputs[4595]);
    assign layer6_outputs[4590] = (layer5_outputs[1501]) & ~(layer5_outputs[4915]);
    assign layer6_outputs[4591] = layer5_outputs[1220];
    assign layer6_outputs[4592] = ~(layer5_outputs[1023]);
    assign layer6_outputs[4593] = ~(layer5_outputs[2917]) | (layer5_outputs[4127]);
    assign layer6_outputs[4594] = layer5_outputs[3962];
    assign layer6_outputs[4595] = (layer5_outputs[3925]) & ~(layer5_outputs[2309]);
    assign layer6_outputs[4596] = ~((layer5_outputs[910]) ^ (layer5_outputs[2993]));
    assign layer6_outputs[4597] = ~(layer5_outputs[1046]);
    assign layer6_outputs[4598] = (layer5_outputs[3510]) ^ (layer5_outputs[687]);
    assign layer6_outputs[4599] = ~(layer5_outputs[2138]);
    assign layer6_outputs[4600] = ~(layer5_outputs[814]);
    assign layer6_outputs[4601] = ~(layer5_outputs[4293]);
    assign layer6_outputs[4602] = layer5_outputs[26];
    assign layer6_outputs[4603] = ~((layer5_outputs[1254]) ^ (layer5_outputs[103]));
    assign layer6_outputs[4604] = layer5_outputs[2627];
    assign layer6_outputs[4605] = layer5_outputs[2104];
    assign layer6_outputs[4606] = layer5_outputs[1308];
    assign layer6_outputs[4607] = ~(layer5_outputs[1386]);
    assign layer6_outputs[4608] = (layer5_outputs[2919]) & ~(layer5_outputs[4735]);
    assign layer6_outputs[4609] = ~(layer5_outputs[2676]);
    assign layer6_outputs[4610] = layer5_outputs[3649];
    assign layer6_outputs[4611] = ~(layer5_outputs[1443]);
    assign layer6_outputs[4612] = layer5_outputs[415];
    assign layer6_outputs[4613] = ~((layer5_outputs[147]) ^ (layer5_outputs[2629]));
    assign layer6_outputs[4614] = layer5_outputs[2220];
    assign layer6_outputs[4615] = (layer5_outputs[3255]) ^ (layer5_outputs[744]);
    assign layer6_outputs[4616] = ~(layer5_outputs[69]);
    assign layer6_outputs[4617] = ~(layer5_outputs[3927]);
    assign layer6_outputs[4618] = ~(layer5_outputs[3043]);
    assign layer6_outputs[4619] = (layer5_outputs[3160]) & ~(layer5_outputs[4538]);
    assign layer6_outputs[4620] = ~(layer5_outputs[3096]);
    assign layer6_outputs[4621] = ~(layer5_outputs[4276]);
    assign layer6_outputs[4622] = (layer5_outputs[4876]) ^ (layer5_outputs[2894]);
    assign layer6_outputs[4623] = layer5_outputs[3371];
    assign layer6_outputs[4624] = (layer5_outputs[534]) & (layer5_outputs[1748]);
    assign layer6_outputs[4625] = ~((layer5_outputs[1947]) ^ (layer5_outputs[5119]));
    assign layer6_outputs[4626] = layer5_outputs[2561];
    assign layer6_outputs[4627] = ~(layer5_outputs[4252]) | (layer5_outputs[2879]);
    assign layer6_outputs[4628] = ~(layer5_outputs[1530]);
    assign layer6_outputs[4629] = ~(layer5_outputs[1236]);
    assign layer6_outputs[4630] = ~(layer5_outputs[1044]);
    assign layer6_outputs[4631] = ~(layer5_outputs[1641]);
    assign layer6_outputs[4632] = ~((layer5_outputs[4246]) ^ (layer5_outputs[1651]));
    assign layer6_outputs[4633] = (layer5_outputs[1981]) ^ (layer5_outputs[2521]);
    assign layer6_outputs[4634] = ~((layer5_outputs[2749]) ^ (layer5_outputs[2967]));
    assign layer6_outputs[4635] = layer5_outputs[3411];
    assign layer6_outputs[4636] = ~(layer5_outputs[1550]);
    assign layer6_outputs[4637] = ~(layer5_outputs[40]);
    assign layer6_outputs[4638] = ~(layer5_outputs[913]);
    assign layer6_outputs[4639] = (layer5_outputs[2917]) & (layer5_outputs[4807]);
    assign layer6_outputs[4640] = ~((layer5_outputs[1496]) & (layer5_outputs[2554]));
    assign layer6_outputs[4641] = ~(layer5_outputs[520]);
    assign layer6_outputs[4642] = layer5_outputs[3539];
    assign layer6_outputs[4643] = ~((layer5_outputs[4368]) & (layer5_outputs[372]));
    assign layer6_outputs[4644] = ~((layer5_outputs[841]) & (layer5_outputs[3436]));
    assign layer6_outputs[4645] = layer5_outputs[2434];
    assign layer6_outputs[4646] = ~(layer5_outputs[4165]) | (layer5_outputs[414]);
    assign layer6_outputs[4647] = ~(layer5_outputs[4875]) | (layer5_outputs[1733]);
    assign layer6_outputs[4648] = ~(layer5_outputs[4654]);
    assign layer6_outputs[4649] = ~(layer5_outputs[3726]);
    assign layer6_outputs[4650] = (layer5_outputs[4644]) ^ (layer5_outputs[419]);
    assign layer6_outputs[4651] = (layer5_outputs[2040]) ^ (layer5_outputs[3982]);
    assign layer6_outputs[4652] = (layer5_outputs[1886]) | (layer5_outputs[2039]);
    assign layer6_outputs[4653] = (layer5_outputs[3857]) ^ (layer5_outputs[4027]);
    assign layer6_outputs[4654] = ~((layer5_outputs[3854]) ^ (layer5_outputs[2928]));
    assign layer6_outputs[4655] = ~((layer5_outputs[2840]) ^ (layer5_outputs[5102]));
    assign layer6_outputs[4656] = ~((layer5_outputs[3684]) ^ (layer5_outputs[1139]));
    assign layer6_outputs[4657] = ~(layer5_outputs[1259]);
    assign layer6_outputs[4658] = ~(layer5_outputs[1099]);
    assign layer6_outputs[4659] = ~(layer5_outputs[1390]) | (layer5_outputs[4156]);
    assign layer6_outputs[4660] = ~(layer5_outputs[3006]);
    assign layer6_outputs[4661] = (layer5_outputs[1784]) | (layer5_outputs[3024]);
    assign layer6_outputs[4662] = ~(layer5_outputs[2534]);
    assign layer6_outputs[4663] = ~(layer5_outputs[1240]);
    assign layer6_outputs[4664] = layer5_outputs[1607];
    assign layer6_outputs[4665] = 1'b0;
    assign layer6_outputs[4666] = ~(layer5_outputs[2752]);
    assign layer6_outputs[4667] = ~((layer5_outputs[3446]) ^ (layer5_outputs[2186]));
    assign layer6_outputs[4668] = ~(layer5_outputs[2976]);
    assign layer6_outputs[4669] = (layer5_outputs[110]) & (layer5_outputs[4635]);
    assign layer6_outputs[4670] = layer5_outputs[1864];
    assign layer6_outputs[4671] = ~((layer5_outputs[4124]) ^ (layer5_outputs[4287]));
    assign layer6_outputs[4672] = ~((layer5_outputs[1630]) & (layer5_outputs[4616]));
    assign layer6_outputs[4673] = ~(layer5_outputs[3945]);
    assign layer6_outputs[4674] = ~(layer5_outputs[3031]);
    assign layer6_outputs[4675] = (layer5_outputs[1310]) & ~(layer5_outputs[584]);
    assign layer6_outputs[4676] = layer5_outputs[3058];
    assign layer6_outputs[4677] = ~(layer5_outputs[1300]);
    assign layer6_outputs[4678] = layer5_outputs[1754];
    assign layer6_outputs[4679] = ~(layer5_outputs[2544]) | (layer5_outputs[3083]);
    assign layer6_outputs[4680] = ~(layer5_outputs[4534]);
    assign layer6_outputs[4681] = ~((layer5_outputs[3753]) ^ (layer5_outputs[3655]));
    assign layer6_outputs[4682] = ~(layer5_outputs[2420]);
    assign layer6_outputs[4683] = ~(layer5_outputs[177]);
    assign layer6_outputs[4684] = (layer5_outputs[2934]) ^ (layer5_outputs[1097]);
    assign layer6_outputs[4685] = ~(layer5_outputs[691]);
    assign layer6_outputs[4686] = (layer5_outputs[1917]) & ~(layer5_outputs[1796]);
    assign layer6_outputs[4687] = ~(layer5_outputs[2469]);
    assign layer6_outputs[4688] = ~(layer5_outputs[2580]) | (layer5_outputs[4811]);
    assign layer6_outputs[4689] = layer5_outputs[2748];
    assign layer6_outputs[4690] = (layer5_outputs[2729]) & (layer5_outputs[158]);
    assign layer6_outputs[4691] = layer5_outputs[2445];
    assign layer6_outputs[4692] = layer5_outputs[2925];
    assign layer6_outputs[4693] = layer5_outputs[2009];
    assign layer6_outputs[4694] = (layer5_outputs[2427]) & ~(layer5_outputs[1948]);
    assign layer6_outputs[4695] = (layer5_outputs[3415]) ^ (layer5_outputs[3315]);
    assign layer6_outputs[4696] = ~((layer5_outputs[3672]) ^ (layer5_outputs[265]));
    assign layer6_outputs[4697] = ~((layer5_outputs[27]) | (layer5_outputs[3331]));
    assign layer6_outputs[4698] = 1'b1;
    assign layer6_outputs[4699] = ~(layer5_outputs[1851]);
    assign layer6_outputs[4700] = layer5_outputs[4896];
    assign layer6_outputs[4701] = layer5_outputs[1168];
    assign layer6_outputs[4702] = (layer5_outputs[3833]) ^ (layer5_outputs[221]);
    assign layer6_outputs[4703] = (layer5_outputs[1471]) ^ (layer5_outputs[2070]);
    assign layer6_outputs[4704] = layer5_outputs[1261];
    assign layer6_outputs[4705] = ~(layer5_outputs[3755]);
    assign layer6_outputs[4706] = layer5_outputs[4842];
    assign layer6_outputs[4707] = ~(layer5_outputs[1283]) | (layer5_outputs[3092]);
    assign layer6_outputs[4708] = ~(layer5_outputs[2402]);
    assign layer6_outputs[4709] = ~(layer5_outputs[3886]);
    assign layer6_outputs[4710] = (layer5_outputs[4546]) ^ (layer5_outputs[3589]);
    assign layer6_outputs[4711] = (layer5_outputs[219]) & ~(layer5_outputs[3614]);
    assign layer6_outputs[4712] = (layer5_outputs[2340]) ^ (layer5_outputs[3265]);
    assign layer6_outputs[4713] = ~((layer5_outputs[2170]) | (layer5_outputs[2681]));
    assign layer6_outputs[4714] = ~((layer5_outputs[2201]) & (layer5_outputs[4235]));
    assign layer6_outputs[4715] = layer5_outputs[881];
    assign layer6_outputs[4716] = layer5_outputs[1800];
    assign layer6_outputs[4717] = layer5_outputs[3686];
    assign layer6_outputs[4718] = ~((layer5_outputs[4302]) ^ (layer5_outputs[1609]));
    assign layer6_outputs[4719] = ~((layer5_outputs[4952]) & (layer5_outputs[3080]));
    assign layer6_outputs[4720] = layer5_outputs[1146];
    assign layer6_outputs[4721] = ~(layer5_outputs[3731]);
    assign layer6_outputs[4722] = layer5_outputs[5073];
    assign layer6_outputs[4723] = ~(layer5_outputs[172]);
    assign layer6_outputs[4724] = (layer5_outputs[1878]) & ~(layer5_outputs[1235]);
    assign layer6_outputs[4725] = 1'b1;
    assign layer6_outputs[4726] = ~((layer5_outputs[1294]) & (layer5_outputs[327]));
    assign layer6_outputs[4727] = (layer5_outputs[2215]) & ~(layer5_outputs[2589]);
    assign layer6_outputs[4728] = ~((layer5_outputs[3291]) ^ (layer5_outputs[4292]));
    assign layer6_outputs[4729] = layer5_outputs[1828];
    assign layer6_outputs[4730] = ~((layer5_outputs[4038]) | (layer5_outputs[2426]));
    assign layer6_outputs[4731] = ~((layer5_outputs[2022]) | (layer5_outputs[3832]));
    assign layer6_outputs[4732] = layer5_outputs[3236];
    assign layer6_outputs[4733] = ~(layer5_outputs[4249]);
    assign layer6_outputs[4734] = ~((layer5_outputs[4957]) ^ (layer5_outputs[359]));
    assign layer6_outputs[4735] = layer5_outputs[138];
    assign layer6_outputs[4736] = layer5_outputs[1314];
    assign layer6_outputs[4737] = ~((layer5_outputs[2829]) | (layer5_outputs[1547]));
    assign layer6_outputs[4738] = layer5_outputs[4090];
    assign layer6_outputs[4739] = ~(layer5_outputs[980]);
    assign layer6_outputs[4740] = layer5_outputs[4502];
    assign layer6_outputs[4741] = ~(layer5_outputs[353]) | (layer5_outputs[199]);
    assign layer6_outputs[4742] = ~(layer5_outputs[2530]);
    assign layer6_outputs[4743] = (layer5_outputs[2977]) | (layer5_outputs[4882]);
    assign layer6_outputs[4744] = layer5_outputs[3444];
    assign layer6_outputs[4745] = ~(layer5_outputs[4053]);
    assign layer6_outputs[4746] = layer5_outputs[3902];
    assign layer6_outputs[4747] = ~((layer5_outputs[1859]) & (layer5_outputs[894]));
    assign layer6_outputs[4748] = ~((layer5_outputs[4298]) & (layer5_outputs[1906]));
    assign layer6_outputs[4749] = ~((layer5_outputs[3986]) | (layer5_outputs[4659]));
    assign layer6_outputs[4750] = layer5_outputs[1800];
    assign layer6_outputs[4751] = (layer5_outputs[160]) | (layer5_outputs[1053]);
    assign layer6_outputs[4752] = (layer5_outputs[4851]) | (layer5_outputs[2418]);
    assign layer6_outputs[4753] = ~(layer5_outputs[162]);
    assign layer6_outputs[4754] = ~(layer5_outputs[2655]);
    assign layer6_outputs[4755] = layer5_outputs[686];
    assign layer6_outputs[4756] = ~(layer5_outputs[370]);
    assign layer6_outputs[4757] = layer5_outputs[4410];
    assign layer6_outputs[4758] = ~(layer5_outputs[4813]);
    assign layer6_outputs[4759] = (layer5_outputs[2056]) | (layer5_outputs[4542]);
    assign layer6_outputs[4760] = layer5_outputs[2093];
    assign layer6_outputs[4761] = layer5_outputs[2671];
    assign layer6_outputs[4762] = layer5_outputs[4849];
    assign layer6_outputs[4763] = (layer5_outputs[2250]) | (layer5_outputs[4177]);
    assign layer6_outputs[4764] = (layer5_outputs[3391]) | (layer5_outputs[1617]);
    assign layer6_outputs[4765] = ~((layer5_outputs[1504]) ^ (layer5_outputs[764]));
    assign layer6_outputs[4766] = ~(layer5_outputs[3280]);
    assign layer6_outputs[4767] = ~(layer5_outputs[1459]);
    assign layer6_outputs[4768] = layer5_outputs[4125];
    assign layer6_outputs[4769] = (layer5_outputs[1073]) ^ (layer5_outputs[867]);
    assign layer6_outputs[4770] = ~((layer5_outputs[680]) & (layer5_outputs[1795]));
    assign layer6_outputs[4771] = (layer5_outputs[3404]) | (layer5_outputs[870]);
    assign layer6_outputs[4772] = ~(layer5_outputs[2070]);
    assign layer6_outputs[4773] = layer5_outputs[195];
    assign layer6_outputs[4774] = (layer5_outputs[3322]) | (layer5_outputs[4407]);
    assign layer6_outputs[4775] = (layer5_outputs[3114]) | (layer5_outputs[3184]);
    assign layer6_outputs[4776] = (layer5_outputs[2712]) ^ (layer5_outputs[2054]);
    assign layer6_outputs[4777] = ~(layer5_outputs[2659]);
    assign layer6_outputs[4778] = layer5_outputs[289];
    assign layer6_outputs[4779] = ~(layer5_outputs[2730]) | (layer5_outputs[4499]);
    assign layer6_outputs[4780] = ~((layer5_outputs[2053]) & (layer5_outputs[3548]));
    assign layer6_outputs[4781] = (layer5_outputs[2258]) | (layer5_outputs[3099]);
    assign layer6_outputs[4782] = layer5_outputs[4776];
    assign layer6_outputs[4783] = layer5_outputs[2319];
    assign layer6_outputs[4784] = ~(layer5_outputs[3425]);
    assign layer6_outputs[4785] = ~(layer5_outputs[2802]);
    assign layer6_outputs[4786] = 1'b1;
    assign layer6_outputs[4787] = ~(layer5_outputs[2294]) | (layer5_outputs[4215]);
    assign layer6_outputs[4788] = ~(layer5_outputs[1927]);
    assign layer6_outputs[4789] = layer5_outputs[1774];
    assign layer6_outputs[4790] = ~(layer5_outputs[995]);
    assign layer6_outputs[4791] = layer5_outputs[1884];
    assign layer6_outputs[4792] = layer5_outputs[4485];
    assign layer6_outputs[4793] = ~(layer5_outputs[2146]);
    assign layer6_outputs[4794] = ~((layer5_outputs[2958]) ^ (layer5_outputs[1855]));
    assign layer6_outputs[4795] = layer5_outputs[3733];
    assign layer6_outputs[4796] = ~(layer5_outputs[1251]);
    assign layer6_outputs[4797] = (layer5_outputs[2705]) | (layer5_outputs[1450]);
    assign layer6_outputs[4798] = ~(layer5_outputs[397]);
    assign layer6_outputs[4799] = layer5_outputs[3848];
    assign layer6_outputs[4800] = ~(layer5_outputs[4174]);
    assign layer6_outputs[4801] = ~(layer5_outputs[557]);
    assign layer6_outputs[4802] = layer5_outputs[1135];
    assign layer6_outputs[4803] = ~(layer5_outputs[2490]);
    assign layer6_outputs[4804] = ~((layer5_outputs[1673]) | (layer5_outputs[1503]));
    assign layer6_outputs[4805] = 1'b0;
    assign layer6_outputs[4806] = ~(layer5_outputs[463]);
    assign layer6_outputs[4807] = ~(layer5_outputs[520]);
    assign layer6_outputs[4808] = (layer5_outputs[1027]) & ~(layer5_outputs[1251]);
    assign layer6_outputs[4809] = (layer5_outputs[1385]) | (layer5_outputs[264]);
    assign layer6_outputs[4810] = (layer5_outputs[4286]) ^ (layer5_outputs[1863]);
    assign layer6_outputs[4811] = ~(layer5_outputs[4157]) | (layer5_outputs[950]);
    assign layer6_outputs[4812] = ~((layer5_outputs[775]) ^ (layer5_outputs[3531]));
    assign layer6_outputs[4813] = ~(layer5_outputs[3008]);
    assign layer6_outputs[4814] = (layer5_outputs[570]) & ~(layer5_outputs[2524]);
    assign layer6_outputs[4815] = (layer5_outputs[4622]) & (layer5_outputs[3643]);
    assign layer6_outputs[4816] = ~(layer5_outputs[4763]);
    assign layer6_outputs[4817] = layer5_outputs[4972];
    assign layer6_outputs[4818] = ~(layer5_outputs[3634]);
    assign layer6_outputs[4819] = ~(layer5_outputs[4447]);
    assign layer6_outputs[4820] = (layer5_outputs[3881]) ^ (layer5_outputs[3796]);
    assign layer6_outputs[4821] = ~((layer5_outputs[2362]) | (layer5_outputs[3003]));
    assign layer6_outputs[4822] = ~((layer5_outputs[899]) ^ (layer5_outputs[2796]));
    assign layer6_outputs[4823] = ~(layer5_outputs[3556]);
    assign layer6_outputs[4824] = ~(layer5_outputs[942]);
    assign layer6_outputs[4825] = layer5_outputs[3521];
    assign layer6_outputs[4826] = ~(layer5_outputs[901]);
    assign layer6_outputs[4827] = layer5_outputs[4837];
    assign layer6_outputs[4828] = ~(layer5_outputs[3559]);
    assign layer6_outputs[4829] = ~(layer5_outputs[2228]);
    assign layer6_outputs[4830] = layer5_outputs[2878];
    assign layer6_outputs[4831] = 1'b1;
    assign layer6_outputs[4832] = ~(layer5_outputs[4008]);
    assign layer6_outputs[4833] = ~((layer5_outputs[2546]) & (layer5_outputs[1059]));
    assign layer6_outputs[4834] = ~(layer5_outputs[3153]) | (layer5_outputs[935]);
    assign layer6_outputs[4835] = ~(layer5_outputs[2904]);
    assign layer6_outputs[4836] = ~((layer5_outputs[401]) & (layer5_outputs[3234]));
    assign layer6_outputs[4837] = layer5_outputs[4681];
    assign layer6_outputs[4838] = layer5_outputs[4337];
    assign layer6_outputs[4839] = layer5_outputs[1672];
    assign layer6_outputs[4840] = layer5_outputs[825];
    assign layer6_outputs[4841] = layer5_outputs[4403];
    assign layer6_outputs[4842] = layer5_outputs[2302];
    assign layer6_outputs[4843] = layer5_outputs[246];
    assign layer6_outputs[4844] = layer5_outputs[2440];
    assign layer6_outputs[4845] = (layer5_outputs[338]) ^ (layer5_outputs[2603]);
    assign layer6_outputs[4846] = ~((layer5_outputs[2950]) ^ (layer5_outputs[4084]));
    assign layer6_outputs[4847] = ~((layer5_outputs[3897]) ^ (layer5_outputs[3196]));
    assign layer6_outputs[4848] = ~(layer5_outputs[4680]);
    assign layer6_outputs[4849] = ~(layer5_outputs[3007]) | (layer5_outputs[1654]);
    assign layer6_outputs[4850] = (layer5_outputs[4395]) & (layer5_outputs[3112]);
    assign layer6_outputs[4851] = layer5_outputs[617];
    assign layer6_outputs[4852] = (layer5_outputs[2938]) ^ (layer5_outputs[3491]);
    assign layer6_outputs[4853] = 1'b0;
    assign layer6_outputs[4854] = (layer5_outputs[1942]) & ~(layer5_outputs[2069]);
    assign layer6_outputs[4855] = layer5_outputs[2586];
    assign layer6_outputs[4856] = ~(layer5_outputs[1690]);
    assign layer6_outputs[4857] = ~(layer5_outputs[884]) | (layer5_outputs[4189]);
    assign layer6_outputs[4858] = ~((layer5_outputs[935]) & (layer5_outputs[1780]));
    assign layer6_outputs[4859] = ~(layer5_outputs[3726]);
    assign layer6_outputs[4860] = (layer5_outputs[2002]) & (layer5_outputs[3597]);
    assign layer6_outputs[4861] = layer5_outputs[179];
    assign layer6_outputs[4862] = ~(layer5_outputs[3386]);
    assign layer6_outputs[4863] = (layer5_outputs[2806]) & (layer5_outputs[2916]);
    assign layer6_outputs[4864] = layer5_outputs[3311];
    assign layer6_outputs[4865] = ~(layer5_outputs[3183]);
    assign layer6_outputs[4866] = ~(layer5_outputs[3283]);
    assign layer6_outputs[4867] = layer5_outputs[2064];
    assign layer6_outputs[4868] = ~(layer5_outputs[1525]);
    assign layer6_outputs[4869] = (layer5_outputs[611]) & ~(layer5_outputs[3801]);
    assign layer6_outputs[4870] = layer5_outputs[4908];
    assign layer6_outputs[4871] = layer5_outputs[3711];
    assign layer6_outputs[4872] = layer5_outputs[2167];
    assign layer6_outputs[4873] = ~((layer5_outputs[2253]) ^ (layer5_outputs[1827]));
    assign layer6_outputs[4874] = ~(layer5_outputs[193]);
    assign layer6_outputs[4875] = ~(layer5_outputs[4017]) | (layer5_outputs[4384]);
    assign layer6_outputs[4876] = ~(layer5_outputs[870]);
    assign layer6_outputs[4877] = (layer5_outputs[2401]) & ~(layer5_outputs[4736]);
    assign layer6_outputs[4878] = (layer5_outputs[3014]) | (layer5_outputs[1317]);
    assign layer6_outputs[4879] = ~(layer5_outputs[3519]) | (layer5_outputs[2327]);
    assign layer6_outputs[4880] = layer5_outputs[2151];
    assign layer6_outputs[4881] = layer5_outputs[1864];
    assign layer6_outputs[4882] = layer5_outputs[8];
    assign layer6_outputs[4883] = ~(layer5_outputs[2380]);
    assign layer6_outputs[4884] = (layer5_outputs[232]) | (layer5_outputs[3962]);
    assign layer6_outputs[4885] = ~(layer5_outputs[3439]);
    assign layer6_outputs[4886] = ~(layer5_outputs[4544]);
    assign layer6_outputs[4887] = ~((layer5_outputs[3347]) ^ (layer5_outputs[3913]));
    assign layer6_outputs[4888] = ~((layer5_outputs[3823]) ^ (layer5_outputs[190]));
    assign layer6_outputs[4889] = layer5_outputs[3111];
    assign layer6_outputs[4890] = (layer5_outputs[5008]) & (layer5_outputs[2582]);
    assign layer6_outputs[4891] = (layer5_outputs[3341]) | (layer5_outputs[748]);
    assign layer6_outputs[4892] = ~((layer5_outputs[1657]) | (layer5_outputs[1418]));
    assign layer6_outputs[4893] = layer5_outputs[4047];
    assign layer6_outputs[4894] = layer5_outputs[178];
    assign layer6_outputs[4895] = layer5_outputs[3813];
    assign layer6_outputs[4896] = (layer5_outputs[4514]) ^ (layer5_outputs[3526]);
    assign layer6_outputs[4897] = layer5_outputs[3939];
    assign layer6_outputs[4898] = layer5_outputs[2548];
    assign layer6_outputs[4899] = layer5_outputs[3987];
    assign layer6_outputs[4900] = layer5_outputs[1347];
    assign layer6_outputs[4901] = (layer5_outputs[4767]) & ~(layer5_outputs[329]);
    assign layer6_outputs[4902] = (layer5_outputs[5107]) & ~(layer5_outputs[3717]);
    assign layer6_outputs[4903] = ~(layer5_outputs[2328]);
    assign layer6_outputs[4904] = ~(layer5_outputs[738]);
    assign layer6_outputs[4905] = ~(layer5_outputs[4516]);
    assign layer6_outputs[4906] = 1'b1;
    assign layer6_outputs[4907] = ~(layer5_outputs[470]) | (layer5_outputs[2062]);
    assign layer6_outputs[4908] = layer5_outputs[828];
    assign layer6_outputs[4909] = ~((layer5_outputs[2333]) ^ (layer5_outputs[295]));
    assign layer6_outputs[4910] = ~((layer5_outputs[4840]) | (layer5_outputs[2659]));
    assign layer6_outputs[4911] = (layer5_outputs[55]) & ~(layer5_outputs[809]);
    assign layer6_outputs[4912] = layer5_outputs[361];
    assign layer6_outputs[4913] = ~(layer5_outputs[204]);
    assign layer6_outputs[4914] = layer5_outputs[4521];
    assign layer6_outputs[4915] = ~(layer5_outputs[2559]);
    assign layer6_outputs[4916] = ~(layer5_outputs[1837]) | (layer5_outputs[388]);
    assign layer6_outputs[4917] = layer5_outputs[168];
    assign layer6_outputs[4918] = ~(layer5_outputs[3763]);
    assign layer6_outputs[4919] = layer5_outputs[1422];
    assign layer6_outputs[4920] = 1'b0;
    assign layer6_outputs[4921] = 1'b0;
    assign layer6_outputs[4922] = ~(layer5_outputs[586]);
    assign layer6_outputs[4923] = (layer5_outputs[4891]) & ~(layer5_outputs[2525]);
    assign layer6_outputs[4924] = (layer5_outputs[4494]) ^ (layer5_outputs[2735]);
    assign layer6_outputs[4925] = (layer5_outputs[3156]) & ~(layer5_outputs[5063]);
    assign layer6_outputs[4926] = ~(layer5_outputs[4633]);
    assign layer6_outputs[4927] = ~(layer5_outputs[2974]);
    assign layer6_outputs[4928] = (layer5_outputs[2231]) & ~(layer5_outputs[3926]);
    assign layer6_outputs[4929] = ~(layer5_outputs[1874]);
    assign layer6_outputs[4930] = ~(layer5_outputs[1778]);
    assign layer6_outputs[4931] = (layer5_outputs[3301]) & ~(layer5_outputs[4783]);
    assign layer6_outputs[4932] = layer5_outputs[2674];
    assign layer6_outputs[4933] = ~((layer5_outputs[4660]) ^ (layer5_outputs[2245]));
    assign layer6_outputs[4934] = layer5_outputs[2804];
    assign layer6_outputs[4935] = ~(layer5_outputs[1543]);
    assign layer6_outputs[4936] = ~(layer5_outputs[2565]);
    assign layer6_outputs[4937] = ~(layer5_outputs[144]);
    assign layer6_outputs[4938] = layer5_outputs[1339];
    assign layer6_outputs[4939] = ~(layer5_outputs[3154]);
    assign layer6_outputs[4940] = ~((layer5_outputs[2011]) ^ (layer5_outputs[2627]));
    assign layer6_outputs[4941] = ~(layer5_outputs[1740]);
    assign layer6_outputs[4942] = (layer5_outputs[4386]) ^ (layer5_outputs[4902]);
    assign layer6_outputs[4943] = ~(layer5_outputs[3134]);
    assign layer6_outputs[4944] = ~((layer5_outputs[3437]) ^ (layer5_outputs[3376]));
    assign layer6_outputs[4945] = layer5_outputs[2120];
    assign layer6_outputs[4946] = ~(layer5_outputs[2507]);
    assign layer6_outputs[4947] = layer5_outputs[2605];
    assign layer6_outputs[4948] = ~((layer5_outputs[1342]) & (layer5_outputs[4864]));
    assign layer6_outputs[4949] = layer5_outputs[769];
    assign layer6_outputs[4950] = ~((layer5_outputs[1967]) & (layer5_outputs[1599]));
    assign layer6_outputs[4951] = ~((layer5_outputs[325]) | (layer5_outputs[4643]));
    assign layer6_outputs[4952] = ~(layer5_outputs[2212]);
    assign layer6_outputs[4953] = layer5_outputs[3013];
    assign layer6_outputs[4954] = layer5_outputs[682];
    assign layer6_outputs[4955] = layer5_outputs[3703];
    assign layer6_outputs[4956] = ~(layer5_outputs[3980]);
    assign layer6_outputs[4957] = layer5_outputs[2692];
    assign layer6_outputs[4958] = ~((layer5_outputs[4310]) & (layer5_outputs[1624]));
    assign layer6_outputs[4959] = (layer5_outputs[3586]) ^ (layer5_outputs[3931]);
    assign layer6_outputs[4960] = ~(layer5_outputs[4852]);
    assign layer6_outputs[4961] = layer5_outputs[2120];
    assign layer6_outputs[4962] = ~(layer5_outputs[2198]);
    assign layer6_outputs[4963] = (layer5_outputs[2701]) & (layer5_outputs[5081]);
    assign layer6_outputs[4964] = ~((layer5_outputs[417]) ^ (layer5_outputs[1327]));
    assign layer6_outputs[4965] = layer5_outputs[469];
    assign layer6_outputs[4966] = (layer5_outputs[4433]) & ~(layer5_outputs[4262]);
    assign layer6_outputs[4967] = layer5_outputs[3567];
    assign layer6_outputs[4968] = layer5_outputs[3828];
    assign layer6_outputs[4969] = ~(layer5_outputs[612]);
    assign layer6_outputs[4970] = ~(layer5_outputs[3993]) | (layer5_outputs[4611]);
    assign layer6_outputs[4971] = (layer5_outputs[2386]) & ~(layer5_outputs[21]);
    assign layer6_outputs[4972] = (layer5_outputs[4460]) & ~(layer5_outputs[2160]);
    assign layer6_outputs[4973] = ~(layer5_outputs[566]);
    assign layer6_outputs[4974] = ~(layer5_outputs[4995]);
    assign layer6_outputs[4975] = ~((layer5_outputs[1212]) & (layer5_outputs[1490]));
    assign layer6_outputs[4976] = (layer5_outputs[1797]) | (layer5_outputs[3754]);
    assign layer6_outputs[4977] = layer5_outputs[908];
    assign layer6_outputs[4978] = (layer5_outputs[4765]) & ~(layer5_outputs[1400]);
    assign layer6_outputs[4979] = ~(layer5_outputs[2931]);
    assign layer6_outputs[4980] = layer5_outputs[167];
    assign layer6_outputs[4981] = ~(layer5_outputs[3954]);
    assign layer6_outputs[4982] = (layer5_outputs[53]) ^ (layer5_outputs[4756]);
    assign layer6_outputs[4983] = ~(layer5_outputs[259]);
    assign layer6_outputs[4984] = ~(layer5_outputs[2668]);
    assign layer6_outputs[4985] = layer5_outputs[2431];
    assign layer6_outputs[4986] = ~((layer5_outputs[4969]) ^ (layer5_outputs[1282]));
    assign layer6_outputs[4987] = ~(layer5_outputs[3899]) | (layer5_outputs[1374]);
    assign layer6_outputs[4988] = (layer5_outputs[4362]) & ~(layer5_outputs[3858]);
    assign layer6_outputs[4989] = (layer5_outputs[1961]) ^ (layer5_outputs[1376]);
    assign layer6_outputs[4990] = (layer5_outputs[1472]) & (layer5_outputs[1681]);
    assign layer6_outputs[4991] = (layer5_outputs[573]) & ~(layer5_outputs[2159]);
    assign layer6_outputs[4992] = layer5_outputs[2302];
    assign layer6_outputs[4993] = 1'b1;
    assign layer6_outputs[4994] = (layer5_outputs[3729]) ^ (layer5_outputs[3899]);
    assign layer6_outputs[4995] = ~((layer5_outputs[3109]) | (layer5_outputs[496]));
    assign layer6_outputs[4996] = 1'b1;
    assign layer6_outputs[4997] = ~(layer5_outputs[243]);
    assign layer6_outputs[4998] = layer5_outputs[598];
    assign layer6_outputs[4999] = ~(layer5_outputs[3677]);
    assign layer6_outputs[5000] = ~(layer5_outputs[768]);
    assign layer6_outputs[5001] = (layer5_outputs[1140]) | (layer5_outputs[3635]);
    assign layer6_outputs[5002] = ~((layer5_outputs[2067]) | (layer5_outputs[3799]));
    assign layer6_outputs[5003] = ~(layer5_outputs[2703]);
    assign layer6_outputs[5004] = ~(layer5_outputs[4825]);
    assign layer6_outputs[5005] = layer5_outputs[2853];
    assign layer6_outputs[5006] = ~((layer5_outputs[2973]) ^ (layer5_outputs[2933]));
    assign layer6_outputs[5007] = layer5_outputs[2970];
    assign layer6_outputs[5008] = ~(layer5_outputs[4064]);
    assign layer6_outputs[5009] = ~(layer5_outputs[2656]);
    assign layer6_outputs[5010] = layer5_outputs[4703];
    assign layer6_outputs[5011] = ~(layer5_outputs[1351]);
    assign layer6_outputs[5012] = ~(layer5_outputs[508]);
    assign layer6_outputs[5013] = 1'b1;
    assign layer6_outputs[5014] = (layer5_outputs[2163]) ^ (layer5_outputs[3397]);
    assign layer6_outputs[5015] = (layer5_outputs[4233]) ^ (layer5_outputs[3563]);
    assign layer6_outputs[5016] = ~(layer5_outputs[1233]);
    assign layer6_outputs[5017] = layer5_outputs[4347];
    assign layer6_outputs[5018] = layer5_outputs[3933];
    assign layer6_outputs[5019] = layer5_outputs[2721];
    assign layer6_outputs[5020] = ~(layer5_outputs[3382]);
    assign layer6_outputs[5021] = ~((layer5_outputs[2823]) | (layer5_outputs[3551]));
    assign layer6_outputs[5022] = ~(layer5_outputs[1039]);
    assign layer6_outputs[5023] = layer5_outputs[33];
    assign layer6_outputs[5024] = ~(layer5_outputs[796]);
    assign layer6_outputs[5025] = layer5_outputs[876];
    assign layer6_outputs[5026] = ~(layer5_outputs[5050]);
    assign layer6_outputs[5027] = ~((layer5_outputs[4399]) ^ (layer5_outputs[2787]));
    assign layer6_outputs[5028] = (layer5_outputs[4341]) & ~(layer5_outputs[3886]);
    assign layer6_outputs[5029] = ~(layer5_outputs[64]) | (layer5_outputs[3599]);
    assign layer6_outputs[5030] = ~((layer5_outputs[5065]) ^ (layer5_outputs[2525]));
    assign layer6_outputs[5031] = ~(layer5_outputs[3410]);
    assign layer6_outputs[5032] = ~(layer5_outputs[695]);
    assign layer6_outputs[5033] = layer5_outputs[3108];
    assign layer6_outputs[5034] = ~(layer5_outputs[2101]);
    assign layer6_outputs[5035] = ~((layer5_outputs[4831]) ^ (layer5_outputs[4226]));
    assign layer6_outputs[5036] = (layer5_outputs[4397]) | (layer5_outputs[3280]);
    assign layer6_outputs[5037] = ~(layer5_outputs[2602]);
    assign layer6_outputs[5038] = layer5_outputs[2474];
    assign layer6_outputs[5039] = ~(layer5_outputs[3701]);
    assign layer6_outputs[5040] = ~(layer5_outputs[560]);
    assign layer6_outputs[5041] = ~(layer5_outputs[2687]);
    assign layer6_outputs[5042] = (layer5_outputs[3122]) ^ (layer5_outputs[2747]);
    assign layer6_outputs[5043] = ~(layer5_outputs[2635]);
    assign layer6_outputs[5044] = ~((layer5_outputs[12]) ^ (layer5_outputs[362]));
    assign layer6_outputs[5045] = layer5_outputs[2437];
    assign layer6_outputs[5046] = ~(layer5_outputs[4159]);
    assign layer6_outputs[5047] = ~(layer5_outputs[5027]) | (layer5_outputs[1203]);
    assign layer6_outputs[5048] = layer5_outputs[2405];
    assign layer6_outputs[5049] = ~((layer5_outputs[1295]) ^ (layer5_outputs[13]));
    assign layer6_outputs[5050] = ~(layer5_outputs[1137]);
    assign layer6_outputs[5051] = layer5_outputs[485];
    assign layer6_outputs[5052] = ~(layer5_outputs[4435]);
    assign layer6_outputs[5053] = layer5_outputs[3045];
    assign layer6_outputs[5054] = layer5_outputs[1101];
    assign layer6_outputs[5055] = (layer5_outputs[825]) & ~(layer5_outputs[3765]);
    assign layer6_outputs[5056] = ~((layer5_outputs[699]) | (layer5_outputs[1555]));
    assign layer6_outputs[5057] = ~((layer5_outputs[3173]) ^ (layer5_outputs[2936]));
    assign layer6_outputs[5058] = ~(layer5_outputs[1613]);
    assign layer6_outputs[5059] = layer5_outputs[1840];
    assign layer6_outputs[5060] = ~(layer5_outputs[1129]);
    assign layer6_outputs[5061] = ~((layer5_outputs[4042]) ^ (layer5_outputs[2291]));
    assign layer6_outputs[5062] = (layer5_outputs[3520]) & ~(layer5_outputs[3935]);
    assign layer6_outputs[5063] = ~((layer5_outputs[1747]) | (layer5_outputs[4247]));
    assign layer6_outputs[5064] = ~((layer5_outputs[500]) ^ (layer5_outputs[3026]));
    assign layer6_outputs[5065] = ~(layer5_outputs[4614]);
    assign layer6_outputs[5066] = ~((layer5_outputs[1249]) ^ (layer5_outputs[2313]));
    assign layer6_outputs[5067] = ~(layer5_outputs[2489]);
    assign layer6_outputs[5068] = layer5_outputs[4028];
    assign layer6_outputs[5069] = layer5_outputs[1642];
    assign layer6_outputs[5070] = (layer5_outputs[73]) ^ (layer5_outputs[514]);
    assign layer6_outputs[5071] = layer5_outputs[871];
    assign layer6_outputs[5072] = layer5_outputs[3105];
    assign layer6_outputs[5073] = layer5_outputs[4799];
    assign layer6_outputs[5074] = (layer5_outputs[1121]) & ~(layer5_outputs[3753]);
    assign layer6_outputs[5075] = layer5_outputs[4605];
    assign layer6_outputs[5076] = ~(layer5_outputs[2318]) | (layer5_outputs[2196]);
    assign layer6_outputs[5077] = (layer5_outputs[3121]) & ~(layer5_outputs[3233]);
    assign layer6_outputs[5078] = ~((layer5_outputs[2465]) & (layer5_outputs[3441]));
    assign layer6_outputs[5079] = ~(layer5_outputs[4184]);
    assign layer6_outputs[5080] = ~(layer5_outputs[2310]);
    assign layer6_outputs[5081] = (layer5_outputs[2735]) ^ (layer5_outputs[1881]);
    assign layer6_outputs[5082] = ~(layer5_outputs[145]) | (layer5_outputs[1333]);
    assign layer6_outputs[5083] = ~(layer5_outputs[3013]);
    assign layer6_outputs[5084] = ~(layer5_outputs[2074]) | (layer5_outputs[3952]);
    assign layer6_outputs[5085] = ~(layer5_outputs[4895]);
    assign layer6_outputs[5086] = ~((layer5_outputs[799]) | (layer5_outputs[207]));
    assign layer6_outputs[5087] = ~(layer5_outputs[4608]) | (layer5_outputs[261]);
    assign layer6_outputs[5088] = layer5_outputs[4049];
    assign layer6_outputs[5089] = ~(layer5_outputs[4725]);
    assign layer6_outputs[5090] = ~((layer5_outputs[399]) & (layer5_outputs[2793]));
    assign layer6_outputs[5091] = ~((layer5_outputs[2899]) | (layer5_outputs[2645]));
    assign layer6_outputs[5092] = (layer5_outputs[4865]) & (layer5_outputs[1077]);
    assign layer6_outputs[5093] = ~(layer5_outputs[1756]);
    assign layer6_outputs[5094] = layer5_outputs[3003];
    assign layer6_outputs[5095] = ~(layer5_outputs[2755]);
    assign layer6_outputs[5096] = (layer5_outputs[4065]) & (layer5_outputs[4091]);
    assign layer6_outputs[5097] = ~(layer5_outputs[4566]) | (layer5_outputs[3926]);
    assign layer6_outputs[5098] = layer5_outputs[3929];
    assign layer6_outputs[5099] = (layer5_outputs[3555]) & ~(layer5_outputs[4647]);
    assign layer6_outputs[5100] = ~((layer5_outputs[2337]) & (layer5_outputs[4719]));
    assign layer6_outputs[5101] = ~(layer5_outputs[3657]);
    assign layer6_outputs[5102] = layer5_outputs[3535];
    assign layer6_outputs[5103] = layer5_outputs[2090];
    assign layer6_outputs[5104] = ~(layer5_outputs[4031]);
    assign layer6_outputs[5105] = ~((layer5_outputs[2257]) | (layer5_outputs[94]));
    assign layer6_outputs[5106] = ~((layer5_outputs[4146]) ^ (layer5_outputs[2293]));
    assign layer6_outputs[5107] = ~(layer5_outputs[3951]);
    assign layer6_outputs[5108] = layer5_outputs[2096];
    assign layer6_outputs[5109] = layer5_outputs[2031];
    assign layer6_outputs[5110] = ~((layer5_outputs[3201]) & (layer5_outputs[4125]));
    assign layer6_outputs[5111] = ~(layer5_outputs[2257]);
    assign layer6_outputs[5112] = ~(layer5_outputs[236]);
    assign layer6_outputs[5113] = layer5_outputs[4646];
    assign layer6_outputs[5114] = (layer5_outputs[1218]) ^ (layer5_outputs[4111]);
    assign layer6_outputs[5115] = layer5_outputs[720];
    assign layer6_outputs[5116] = ~(layer5_outputs[3816]) | (layer5_outputs[679]);
    assign layer6_outputs[5117] = ~(layer5_outputs[2371]);
    assign layer6_outputs[5118] = layer5_outputs[4999];
    assign layer6_outputs[5119] = ~(layer5_outputs[4769]);
    assign outputs[0] = ~(layer6_outputs[1064]);
    assign outputs[1] = ~(layer6_outputs[3992]);
    assign outputs[2] = (layer6_outputs[1046]) ^ (layer6_outputs[3290]);
    assign outputs[3] = ~(layer6_outputs[4324]);
    assign outputs[4] = ~(layer6_outputs[1616]);
    assign outputs[5] = ~(layer6_outputs[4135]);
    assign outputs[6] = ~(layer6_outputs[1921]);
    assign outputs[7] = ~(layer6_outputs[2578]);
    assign outputs[8] = layer6_outputs[2309];
    assign outputs[9] = layer6_outputs[2733];
    assign outputs[10] = layer6_outputs[103];
    assign outputs[11] = layer6_outputs[1292];
    assign outputs[12] = ~(layer6_outputs[4221]);
    assign outputs[13] = ~(layer6_outputs[4097]);
    assign outputs[14] = layer6_outputs[2815];
    assign outputs[15] = layer6_outputs[567];
    assign outputs[16] = layer6_outputs[2068];
    assign outputs[17] = ~(layer6_outputs[18]);
    assign outputs[18] = layer6_outputs[4333];
    assign outputs[19] = layer6_outputs[1792];
    assign outputs[20] = layer6_outputs[815];
    assign outputs[21] = (layer6_outputs[3863]) ^ (layer6_outputs[4488]);
    assign outputs[22] = ~(layer6_outputs[41]);
    assign outputs[23] = layer6_outputs[5024];
    assign outputs[24] = ~((layer6_outputs[885]) ^ (layer6_outputs[3844]));
    assign outputs[25] = ~(layer6_outputs[2956]);
    assign outputs[26] = layer6_outputs[1341];
    assign outputs[27] = layer6_outputs[4944];
    assign outputs[28] = (layer6_outputs[2712]) & ~(layer6_outputs[1170]);
    assign outputs[29] = layer6_outputs[4883];
    assign outputs[30] = ~((layer6_outputs[4796]) & (layer6_outputs[707]));
    assign outputs[31] = ~(layer6_outputs[1289]);
    assign outputs[32] = ~((layer6_outputs[509]) | (layer6_outputs[4995]));
    assign outputs[33] = ~(layer6_outputs[2765]);
    assign outputs[34] = layer6_outputs[1848];
    assign outputs[35] = ~((layer6_outputs[4627]) ^ (layer6_outputs[4672]));
    assign outputs[36] = (layer6_outputs[4635]) ^ (layer6_outputs[1835]);
    assign outputs[37] = ~(layer6_outputs[2108]);
    assign outputs[38] = ~(layer6_outputs[619]) | (layer6_outputs[870]);
    assign outputs[39] = layer6_outputs[2529];
    assign outputs[40] = ~(layer6_outputs[3373]);
    assign outputs[41] = ~(layer6_outputs[2752]);
    assign outputs[42] = ~(layer6_outputs[2959]);
    assign outputs[43] = (layer6_outputs[718]) ^ (layer6_outputs[2062]);
    assign outputs[44] = ~(layer6_outputs[1698]);
    assign outputs[45] = (layer6_outputs[1720]) ^ (layer6_outputs[1409]);
    assign outputs[46] = ~((layer6_outputs[4465]) ^ (layer6_outputs[4326]));
    assign outputs[47] = ~((layer6_outputs[4351]) ^ (layer6_outputs[2027]));
    assign outputs[48] = ~(layer6_outputs[3377]);
    assign outputs[49] = ~(layer6_outputs[3384]);
    assign outputs[50] = layer6_outputs[645];
    assign outputs[51] = layer6_outputs[4390];
    assign outputs[52] = ~(layer6_outputs[2581]);
    assign outputs[53] = ~((layer6_outputs[643]) | (layer6_outputs[3351]));
    assign outputs[54] = ~(layer6_outputs[1859]);
    assign outputs[55] = layer6_outputs[5000];
    assign outputs[56] = layer6_outputs[3194];
    assign outputs[57] = layer6_outputs[3999];
    assign outputs[58] = ~((layer6_outputs[1787]) & (layer6_outputs[1323]));
    assign outputs[59] = layer6_outputs[949];
    assign outputs[60] = ~(layer6_outputs[3584]);
    assign outputs[61] = ~(layer6_outputs[3416]);
    assign outputs[62] = (layer6_outputs[2350]) & ~(layer6_outputs[1723]);
    assign outputs[63] = ~(layer6_outputs[3617]);
    assign outputs[64] = layer6_outputs[2077];
    assign outputs[65] = ~(layer6_outputs[2667]);
    assign outputs[66] = layer6_outputs[1345];
    assign outputs[67] = ~((layer6_outputs[3152]) ^ (layer6_outputs[2998]));
    assign outputs[68] = ~(layer6_outputs[236]);
    assign outputs[69] = ~((layer6_outputs[1877]) ^ (layer6_outputs[2771]));
    assign outputs[70] = ~(layer6_outputs[4927]) | (layer6_outputs[3502]);
    assign outputs[71] = (layer6_outputs[1015]) ^ (layer6_outputs[2004]);
    assign outputs[72] = layer6_outputs[4415];
    assign outputs[73] = ~(layer6_outputs[4523]);
    assign outputs[74] = ~(layer6_outputs[4885]);
    assign outputs[75] = ~(layer6_outputs[3648]);
    assign outputs[76] = layer6_outputs[263];
    assign outputs[77] = layer6_outputs[1800];
    assign outputs[78] = layer6_outputs[5111];
    assign outputs[79] = ~(layer6_outputs[4328]) | (layer6_outputs[4050]);
    assign outputs[80] = (layer6_outputs[3374]) ^ (layer6_outputs[1102]);
    assign outputs[81] = ~(layer6_outputs[3675]);
    assign outputs[82] = layer6_outputs[3539];
    assign outputs[83] = ~((layer6_outputs[4695]) ^ (layer6_outputs[3712]));
    assign outputs[84] = ~(layer6_outputs[665]);
    assign outputs[85] = ~(layer6_outputs[2616]);
    assign outputs[86] = ~(layer6_outputs[2776]);
    assign outputs[87] = ~((layer6_outputs[817]) ^ (layer6_outputs[4304]));
    assign outputs[88] = layer6_outputs[2164];
    assign outputs[89] = ~(layer6_outputs[3191]);
    assign outputs[90] = ~(layer6_outputs[602]);
    assign outputs[91] = ~(layer6_outputs[1953]);
    assign outputs[92] = ~(layer6_outputs[703]);
    assign outputs[93] = layer6_outputs[726];
    assign outputs[94] = layer6_outputs[2346];
    assign outputs[95] = ~((layer6_outputs[1150]) ^ (layer6_outputs[4344]));
    assign outputs[96] = ~(layer6_outputs[3738]);
    assign outputs[97] = (layer6_outputs[2579]) & ~(layer6_outputs[4388]);
    assign outputs[98] = ~(layer6_outputs[2022]);
    assign outputs[99] = ~(layer6_outputs[1299]);
    assign outputs[100] = layer6_outputs[2422];
    assign outputs[101] = layer6_outputs[476];
    assign outputs[102] = layer6_outputs[30];
    assign outputs[103] = layer6_outputs[1734];
    assign outputs[104] = layer6_outputs[1985];
    assign outputs[105] = ~(layer6_outputs[957]);
    assign outputs[106] = layer6_outputs[1725];
    assign outputs[107] = layer6_outputs[4869];
    assign outputs[108] = ~((layer6_outputs[1594]) ^ (layer6_outputs[4729]));
    assign outputs[109] = ~(layer6_outputs[1363]);
    assign outputs[110] = layer6_outputs[443];
    assign outputs[111] = ~(layer6_outputs[4719]);
    assign outputs[112] = layer6_outputs[4565];
    assign outputs[113] = layer6_outputs[4446];
    assign outputs[114] = ~(layer6_outputs[2106]);
    assign outputs[115] = layer6_outputs[4064];
    assign outputs[116] = layer6_outputs[3361];
    assign outputs[117] = ~(layer6_outputs[968]);
    assign outputs[118] = ~(layer6_outputs[4197]);
    assign outputs[119] = layer6_outputs[1718];
    assign outputs[120] = ~((layer6_outputs[4450]) ^ (layer6_outputs[4865]));
    assign outputs[121] = ~(layer6_outputs[1667]);
    assign outputs[122] = (layer6_outputs[996]) & ~(layer6_outputs[1024]);
    assign outputs[123] = layer6_outputs[2008];
    assign outputs[124] = ~((layer6_outputs[810]) | (layer6_outputs[961]));
    assign outputs[125] = ~((layer6_outputs[2610]) | (layer6_outputs[1600]));
    assign outputs[126] = (layer6_outputs[1842]) ^ (layer6_outputs[827]);
    assign outputs[127] = ~(layer6_outputs[4002]);
    assign outputs[128] = ~(layer6_outputs[2105]);
    assign outputs[129] = (layer6_outputs[2769]) & (layer6_outputs[4729]);
    assign outputs[130] = ~(layer6_outputs[4312]);
    assign outputs[131] = layer6_outputs[4222];
    assign outputs[132] = layer6_outputs[2293];
    assign outputs[133] = ~(layer6_outputs[668]);
    assign outputs[134] = ~(layer6_outputs[3608]);
    assign outputs[135] = layer6_outputs[1780];
    assign outputs[136] = ~(layer6_outputs[4025]);
    assign outputs[137] = layer6_outputs[4176];
    assign outputs[138] = layer6_outputs[2201];
    assign outputs[139] = ~(layer6_outputs[4739]);
    assign outputs[140] = ~(layer6_outputs[247]);
    assign outputs[141] = (layer6_outputs[1023]) ^ (layer6_outputs[3806]);
    assign outputs[142] = (layer6_outputs[1732]) & (layer6_outputs[5059]);
    assign outputs[143] = ~((layer6_outputs[3413]) ^ (layer6_outputs[4969]));
    assign outputs[144] = layer6_outputs[2026];
    assign outputs[145] = ~(layer6_outputs[1603]);
    assign outputs[146] = layer6_outputs[2263];
    assign outputs[147] = ~(layer6_outputs[4180]);
    assign outputs[148] = ~(layer6_outputs[1003]);
    assign outputs[149] = ~((layer6_outputs[853]) ^ (layer6_outputs[3038]));
    assign outputs[150] = layer6_outputs[3847];
    assign outputs[151] = layer6_outputs[2130];
    assign outputs[152] = ~((layer6_outputs[1640]) ^ (layer6_outputs[1845]));
    assign outputs[153] = ~(layer6_outputs[3370]);
    assign outputs[154] = ~(layer6_outputs[1830]);
    assign outputs[155] = (layer6_outputs[3054]) & (layer6_outputs[190]);
    assign outputs[156] = ~(layer6_outputs[3533]);
    assign outputs[157] = ~(layer6_outputs[4121]);
    assign outputs[158] = layer6_outputs[1734];
    assign outputs[159] = ~((layer6_outputs[4287]) | (layer6_outputs[2241]));
    assign outputs[160] = ~(layer6_outputs[2794]) | (layer6_outputs[3446]);
    assign outputs[161] = layer6_outputs[385];
    assign outputs[162] = (layer6_outputs[1589]) ^ (layer6_outputs[3104]);
    assign outputs[163] = layer6_outputs[1899];
    assign outputs[164] = layer6_outputs[188];
    assign outputs[165] = ~(layer6_outputs[342]);
    assign outputs[166] = ~((layer6_outputs[1454]) ^ (layer6_outputs[1302]));
    assign outputs[167] = ~(layer6_outputs[2070]);
    assign outputs[168] = layer6_outputs[118];
    assign outputs[169] = (layer6_outputs[2072]) | (layer6_outputs[4632]);
    assign outputs[170] = layer6_outputs[4561];
    assign outputs[171] = ~((layer6_outputs[743]) ^ (layer6_outputs[2662]));
    assign outputs[172] = (layer6_outputs[2407]) | (layer6_outputs[3821]);
    assign outputs[173] = layer6_outputs[211];
    assign outputs[174] = ~((layer6_outputs[686]) ^ (layer6_outputs[124]));
    assign outputs[175] = layer6_outputs[870];
    assign outputs[176] = ~(layer6_outputs[3763]);
    assign outputs[177] = layer6_outputs[3695];
    assign outputs[178] = layer6_outputs[4897];
    assign outputs[179] = layer6_outputs[405];
    assign outputs[180] = layer6_outputs[1773];
    assign outputs[181] = ~(layer6_outputs[3478]);
    assign outputs[182] = layer6_outputs[3663];
    assign outputs[183] = layer6_outputs[1972];
    assign outputs[184] = layer6_outputs[4108];
    assign outputs[185] = ~(layer6_outputs[3330]);
    assign outputs[186] = layer6_outputs[4884];
    assign outputs[187] = layer6_outputs[4649];
    assign outputs[188] = layer6_outputs[3321];
    assign outputs[189] = layer6_outputs[2399];
    assign outputs[190] = layer6_outputs[4844];
    assign outputs[191] = ~((layer6_outputs[4699]) | (layer6_outputs[3053]));
    assign outputs[192] = ~(layer6_outputs[4413]);
    assign outputs[193] = layer6_outputs[4083];
    assign outputs[194] = ~(layer6_outputs[97]);
    assign outputs[195] = ~(layer6_outputs[1351]);
    assign outputs[196] = layer6_outputs[1050];
    assign outputs[197] = ~(layer6_outputs[3897]);
    assign outputs[198] = ~(layer6_outputs[5011]);
    assign outputs[199] = ~(layer6_outputs[1898]);
    assign outputs[200] = ~(layer6_outputs[2001]);
    assign outputs[201] = ~(layer6_outputs[4572]);
    assign outputs[202] = layer6_outputs[3514];
    assign outputs[203] = ~(layer6_outputs[2934]);
    assign outputs[204] = layer6_outputs[3684];
    assign outputs[205] = ~(layer6_outputs[2059]);
    assign outputs[206] = ~(layer6_outputs[4401]);
    assign outputs[207] = layer6_outputs[897];
    assign outputs[208] = layer6_outputs[3955];
    assign outputs[209] = ~(layer6_outputs[716]);
    assign outputs[210] = (layer6_outputs[2697]) & (layer6_outputs[3333]);
    assign outputs[211] = (layer6_outputs[1812]) ^ (layer6_outputs[1468]);
    assign outputs[212] = layer6_outputs[4148];
    assign outputs[213] = layer6_outputs[1005];
    assign outputs[214] = layer6_outputs[1271];
    assign outputs[215] = ~(layer6_outputs[3513]);
    assign outputs[216] = ~(layer6_outputs[2744]);
    assign outputs[217] = layer6_outputs[2239];
    assign outputs[218] = ~(layer6_outputs[487]);
    assign outputs[219] = layer6_outputs[1127];
    assign outputs[220] = ~(layer6_outputs[4012]);
    assign outputs[221] = (layer6_outputs[3852]) & ~(layer6_outputs[3521]);
    assign outputs[222] = layer6_outputs[4671];
    assign outputs[223] = ~(layer6_outputs[3007]);
    assign outputs[224] = ~(layer6_outputs[2834]);
    assign outputs[225] = (layer6_outputs[2546]) ^ (layer6_outputs[3931]);
    assign outputs[226] = layer6_outputs[2479];
    assign outputs[227] = (layer6_outputs[1065]) & ~(layer6_outputs[3012]);
    assign outputs[228] = ~(layer6_outputs[375]);
    assign outputs[229] = ~(layer6_outputs[1475]);
    assign outputs[230] = layer6_outputs[3025];
    assign outputs[231] = ~(layer6_outputs[1221]);
    assign outputs[232] = layer6_outputs[2330];
    assign outputs[233] = layer6_outputs[1398];
    assign outputs[234] = ~((layer6_outputs[1519]) & (layer6_outputs[472]));
    assign outputs[235] = ~((layer6_outputs[88]) | (layer6_outputs[588]));
    assign outputs[236] = layer6_outputs[1760];
    assign outputs[237] = ~((layer6_outputs[1362]) & (layer6_outputs[1204]));
    assign outputs[238] = ~(layer6_outputs[955]);
    assign outputs[239] = ~(layer6_outputs[1879]);
    assign outputs[240] = (layer6_outputs[1544]) & ~(layer6_outputs[768]);
    assign outputs[241] = ~((layer6_outputs[2338]) ^ (layer6_outputs[417]));
    assign outputs[242] = (layer6_outputs[4979]) & ~(layer6_outputs[1478]);
    assign outputs[243] = ~(layer6_outputs[2629]);
    assign outputs[244] = ~(layer6_outputs[3420]);
    assign outputs[245] = ~(layer6_outputs[3076]);
    assign outputs[246] = ~(layer6_outputs[786]);
    assign outputs[247] = layer6_outputs[3088];
    assign outputs[248] = ~((layer6_outputs[4592]) ^ (layer6_outputs[2424]));
    assign outputs[249] = ~((layer6_outputs[4908]) ^ (layer6_outputs[2791]));
    assign outputs[250] = (layer6_outputs[2047]) ^ (layer6_outputs[4163]);
    assign outputs[251] = layer6_outputs[103];
    assign outputs[252] = ~((layer6_outputs[326]) ^ (layer6_outputs[1569]));
    assign outputs[253] = ~(layer6_outputs[1629]);
    assign outputs[254] = layer6_outputs[3435];
    assign outputs[255] = layer6_outputs[3573];
    assign outputs[256] = (layer6_outputs[4103]) ^ (layer6_outputs[4063]);
    assign outputs[257] = ~(layer6_outputs[4442]);
    assign outputs[258] = layer6_outputs[324];
    assign outputs[259] = ~(layer6_outputs[334]);
    assign outputs[260] = layer6_outputs[3613];
    assign outputs[261] = ~(layer6_outputs[1298]);
    assign outputs[262] = ~(layer6_outputs[4885]);
    assign outputs[263] = (layer6_outputs[4843]) ^ (layer6_outputs[3038]);
    assign outputs[264] = ~(layer6_outputs[3510]);
    assign outputs[265] = ~(layer6_outputs[4591]);
    assign outputs[266] = layer6_outputs[2286];
    assign outputs[267] = (layer6_outputs[2544]) ^ (layer6_outputs[1106]);
    assign outputs[268] = ~((layer6_outputs[434]) ^ (layer6_outputs[2310]));
    assign outputs[269] = layer6_outputs[1173];
    assign outputs[270] = ~(layer6_outputs[371]);
    assign outputs[271] = ~(layer6_outputs[4694]);
    assign outputs[272] = ~(layer6_outputs[928]);
    assign outputs[273] = ~((layer6_outputs[3014]) ^ (layer6_outputs[4768]));
    assign outputs[274] = ~(layer6_outputs[143]);
    assign outputs[275] = layer6_outputs[815];
    assign outputs[276] = ~(layer6_outputs[4283]);
    assign outputs[277] = layer6_outputs[2501];
    assign outputs[278] = layer6_outputs[1043];
    assign outputs[279] = layer6_outputs[1199];
    assign outputs[280] = ~(layer6_outputs[72]);
    assign outputs[281] = layer6_outputs[3813];
    assign outputs[282] = ~((layer6_outputs[1944]) ^ (layer6_outputs[2265]));
    assign outputs[283] = layer6_outputs[704];
    assign outputs[284] = layer6_outputs[1915];
    assign outputs[285] = (layer6_outputs[2399]) | (layer6_outputs[2561]);
    assign outputs[286] = ~(layer6_outputs[44]);
    assign outputs[287] = ~(layer6_outputs[2178]);
    assign outputs[288] = ~((layer6_outputs[3440]) ^ (layer6_outputs[1877]));
    assign outputs[289] = layer6_outputs[3726];
    assign outputs[290] = layer6_outputs[1230];
    assign outputs[291] = ~(layer6_outputs[2690]);
    assign outputs[292] = layer6_outputs[3646];
    assign outputs[293] = layer6_outputs[4049];
    assign outputs[294] = ~((layer6_outputs[5109]) ^ (layer6_outputs[1544]));
    assign outputs[295] = ~(layer6_outputs[2913]);
    assign outputs[296] = layer6_outputs[62];
    assign outputs[297] = ~(layer6_outputs[4866]);
    assign outputs[298] = layer6_outputs[1416];
    assign outputs[299] = ~(layer6_outputs[1924]);
    assign outputs[300] = ~(layer6_outputs[4289]);
    assign outputs[301] = ~(layer6_outputs[4102]);
    assign outputs[302] = layer6_outputs[4481];
    assign outputs[303] = ~((layer6_outputs[1954]) ^ (layer6_outputs[2414]));
    assign outputs[304] = layer6_outputs[4870];
    assign outputs[305] = ~(layer6_outputs[611]);
    assign outputs[306] = layer6_outputs[1473];
    assign outputs[307] = ~((layer6_outputs[438]) ^ (layer6_outputs[1599]));
    assign outputs[308] = (layer6_outputs[2425]) & ~(layer6_outputs[1223]);
    assign outputs[309] = ~((layer6_outputs[3457]) ^ (layer6_outputs[3412]));
    assign outputs[310] = layer6_outputs[3472];
    assign outputs[311] = ~(layer6_outputs[1787]);
    assign outputs[312] = ~(layer6_outputs[3495]);
    assign outputs[313] = ~(layer6_outputs[2353]);
    assign outputs[314] = (layer6_outputs[3260]) ^ (layer6_outputs[1368]);
    assign outputs[315] = ~(layer6_outputs[21]);
    assign outputs[316] = layer6_outputs[4867];
    assign outputs[317] = ~(layer6_outputs[2156]) | (layer6_outputs[3218]);
    assign outputs[318] = ~(layer6_outputs[1358]);
    assign outputs[319] = (layer6_outputs[609]) ^ (layer6_outputs[4955]);
    assign outputs[320] = ~(layer6_outputs[1438]);
    assign outputs[321] = ~((layer6_outputs[4854]) | (layer6_outputs[192]));
    assign outputs[322] = ~(layer6_outputs[970]);
    assign outputs[323] = layer6_outputs[410];
    assign outputs[324] = layer6_outputs[3674];
    assign outputs[325] = ~(layer6_outputs[3850]);
    assign outputs[326] = layer6_outputs[3450];
    assign outputs[327] = (layer6_outputs[1945]) | (layer6_outputs[2492]);
    assign outputs[328] = ~(layer6_outputs[2544]);
    assign outputs[329] = ~(layer6_outputs[1220]);
    assign outputs[330] = layer6_outputs[1067];
    assign outputs[331] = layer6_outputs[3021];
    assign outputs[332] = layer6_outputs[1160];
    assign outputs[333] = layer6_outputs[1647];
    assign outputs[334] = layer6_outputs[2364];
    assign outputs[335] = ~(layer6_outputs[242]);
    assign outputs[336] = layer6_outputs[3867];
    assign outputs[337] = layer6_outputs[2937];
    assign outputs[338] = ~(layer6_outputs[1580]);
    assign outputs[339] = ~((layer6_outputs[947]) ^ (layer6_outputs[2376]));
    assign outputs[340] = ~(layer6_outputs[4085]);
    assign outputs[341] = layer6_outputs[257];
    assign outputs[342] = ~(layer6_outputs[1178]);
    assign outputs[343] = (layer6_outputs[83]) ^ (layer6_outputs[2633]);
    assign outputs[344] = ~(layer6_outputs[3061]);
    assign outputs[345] = layer6_outputs[4915];
    assign outputs[346] = ~(layer6_outputs[5017]);
    assign outputs[347] = (layer6_outputs[834]) ^ (layer6_outputs[4479]);
    assign outputs[348] = ~(layer6_outputs[804]);
    assign outputs[349] = ~(layer6_outputs[3982]);
    assign outputs[350] = (layer6_outputs[4265]) ^ (layer6_outputs[4660]);
    assign outputs[351] = layer6_outputs[4270];
    assign outputs[352] = layer6_outputs[4372];
    assign outputs[353] = ~((layer6_outputs[1334]) & (layer6_outputs[2065]));
    assign outputs[354] = layer6_outputs[343];
    assign outputs[355] = ~(layer6_outputs[3546]);
    assign outputs[356] = (layer6_outputs[1339]) ^ (layer6_outputs[4682]);
    assign outputs[357] = ~(layer6_outputs[3704]);
    assign outputs[358] = ~((layer6_outputs[556]) ^ (layer6_outputs[2092]));
    assign outputs[359] = ~(layer6_outputs[4814]);
    assign outputs[360] = layer6_outputs[4055];
    assign outputs[361] = ~((layer6_outputs[4962]) ^ (layer6_outputs[152]));
    assign outputs[362] = ~(layer6_outputs[2851]);
    assign outputs[363] = ~(layer6_outputs[4524]);
    assign outputs[364] = layer6_outputs[1188];
    assign outputs[365] = layer6_outputs[2246];
    assign outputs[366] = ~((layer6_outputs[1265]) | (layer6_outputs[2262]));
    assign outputs[367] = ~((layer6_outputs[1029]) ^ (layer6_outputs[4689]));
    assign outputs[368] = layer6_outputs[1654];
    assign outputs[369] = ~(layer6_outputs[2249]) | (layer6_outputs[234]);
    assign outputs[370] = ~(layer6_outputs[1997]);
    assign outputs[371] = ~(layer6_outputs[1999]);
    assign outputs[372] = layer6_outputs[1494];
    assign outputs[373] = ~((layer6_outputs[2922]) ^ (layer6_outputs[3469]));
    assign outputs[374] = ~((layer6_outputs[1379]) ^ (layer6_outputs[739]));
    assign outputs[375] = ~(layer6_outputs[4629]);
    assign outputs[376] = layer6_outputs[4512];
    assign outputs[377] = ~(layer6_outputs[4878]) | (layer6_outputs[748]);
    assign outputs[378] = (layer6_outputs[3552]) ^ (layer6_outputs[1727]);
    assign outputs[379] = ~(layer6_outputs[210]);
    assign outputs[380] = layer6_outputs[4476];
    assign outputs[381] = ~(layer6_outputs[4463]);
    assign outputs[382] = layer6_outputs[3509];
    assign outputs[383] = ~(layer6_outputs[865]);
    assign outputs[384] = ~(layer6_outputs[1499]);
    assign outputs[385] = ~(layer6_outputs[3593]) | (layer6_outputs[975]);
    assign outputs[386] = layer6_outputs[1642];
    assign outputs[387] = layer6_outputs[3517];
    assign outputs[388] = layer6_outputs[1107];
    assign outputs[389] = ~(layer6_outputs[3982]);
    assign outputs[390] = (layer6_outputs[1327]) ^ (layer6_outputs[3693]);
    assign outputs[391] = (layer6_outputs[4585]) & ~(layer6_outputs[920]);
    assign outputs[392] = (layer6_outputs[4660]) ^ (layer6_outputs[2803]);
    assign outputs[393] = ~(layer6_outputs[2657]) | (layer6_outputs[1585]);
    assign outputs[394] = ~(layer6_outputs[4227]);
    assign outputs[395] = layer6_outputs[2446];
    assign outputs[396] = ~(layer6_outputs[4036]);
    assign outputs[397] = (layer6_outputs[2615]) ^ (layer6_outputs[4307]);
    assign outputs[398] = layer6_outputs[4773];
    assign outputs[399] = ~(layer6_outputs[4924]);
    assign outputs[400] = ~(layer6_outputs[87]);
    assign outputs[401] = ~((layer6_outputs[3032]) ^ (layer6_outputs[39]));
    assign outputs[402] = (layer6_outputs[3973]) ^ (layer6_outputs[2177]);
    assign outputs[403] = ~(layer6_outputs[1786]);
    assign outputs[404] = ~(layer6_outputs[3527]);
    assign outputs[405] = ~(layer6_outputs[1916]);
    assign outputs[406] = layer6_outputs[4232];
    assign outputs[407] = layer6_outputs[4428];
    assign outputs[408] = ~(layer6_outputs[3890]);
    assign outputs[409] = ~(layer6_outputs[1810]);
    assign outputs[410] = (layer6_outputs[2056]) ^ (layer6_outputs[50]);
    assign outputs[411] = ~(layer6_outputs[457]);
    assign outputs[412] = layer6_outputs[2418];
    assign outputs[413] = layer6_outputs[2194];
    assign outputs[414] = (layer6_outputs[427]) & ~(layer6_outputs[1635]);
    assign outputs[415] = layer6_outputs[2093];
    assign outputs[416] = layer6_outputs[4696];
    assign outputs[417] = (layer6_outputs[3900]) & ~(layer6_outputs[1906]);
    assign outputs[418] = ~(layer6_outputs[4419]);
    assign outputs[419] = ~(layer6_outputs[4489]) | (layer6_outputs[202]);
    assign outputs[420] = (layer6_outputs[2265]) ^ (layer6_outputs[1355]);
    assign outputs[421] = ~((layer6_outputs[3093]) ^ (layer6_outputs[1430]));
    assign outputs[422] = layer6_outputs[1762];
    assign outputs[423] = (layer6_outputs[3903]) & (layer6_outputs[679]);
    assign outputs[424] = layer6_outputs[1263];
    assign outputs[425] = ~(layer6_outputs[684]);
    assign outputs[426] = ~((layer6_outputs[534]) ^ (layer6_outputs[43]));
    assign outputs[427] = ~((layer6_outputs[4106]) ^ (layer6_outputs[2124]));
    assign outputs[428] = layer6_outputs[4207];
    assign outputs[429] = ~(layer6_outputs[5100]);
    assign outputs[430] = ~(layer6_outputs[3961]);
    assign outputs[431] = ~(layer6_outputs[4205]);
    assign outputs[432] = ~(layer6_outputs[936]);
    assign outputs[433] = layer6_outputs[3723];
    assign outputs[434] = layer6_outputs[4094];
    assign outputs[435] = ~(layer6_outputs[5035]);
    assign outputs[436] = layer6_outputs[4330];
    assign outputs[437] = ~(layer6_outputs[4547]);
    assign outputs[438] = layer6_outputs[1961];
    assign outputs[439] = ~(layer6_outputs[4532]) | (layer6_outputs[1101]);
    assign outputs[440] = layer6_outputs[4644];
    assign outputs[441] = ~(layer6_outputs[3618]);
    assign outputs[442] = layer6_outputs[508];
    assign outputs[443] = (layer6_outputs[2855]) & ~(layer6_outputs[1942]);
    assign outputs[444] = ~(layer6_outputs[2509]) | (layer6_outputs[393]);
    assign outputs[445] = (layer6_outputs[2357]) ^ (layer6_outputs[3537]);
    assign outputs[446] = ~(layer6_outputs[2329]);
    assign outputs[447] = layer6_outputs[3117];
    assign outputs[448] = ~(layer6_outputs[2311]);
    assign outputs[449] = layer6_outputs[4594];
    assign outputs[450] = ~(layer6_outputs[411]);
    assign outputs[451] = ~((layer6_outputs[809]) ^ (layer6_outputs[578]));
    assign outputs[452] = layer6_outputs[4706];
    assign outputs[453] = layer6_outputs[2496];
    assign outputs[454] = layer6_outputs[1457];
    assign outputs[455] = layer6_outputs[3934];
    assign outputs[456] = ~(layer6_outputs[1735]);
    assign outputs[457] = layer6_outputs[2122];
    assign outputs[458] = layer6_outputs[2194];
    assign outputs[459] = ~(layer6_outputs[549]) | (layer6_outputs[3215]);
    assign outputs[460] = ~(layer6_outputs[1456]);
    assign outputs[461] = (layer6_outputs[3967]) ^ (layer6_outputs[3096]);
    assign outputs[462] = layer6_outputs[2644];
    assign outputs[463] = layer6_outputs[3156];
    assign outputs[464] = ~((layer6_outputs[3483]) & (layer6_outputs[2785]));
    assign outputs[465] = layer6_outputs[3344];
    assign outputs[466] = layer6_outputs[2718];
    assign outputs[467] = ~(layer6_outputs[429]);
    assign outputs[468] = layer6_outputs[1090];
    assign outputs[469] = layer6_outputs[678];
    assign outputs[470] = layer6_outputs[4738];
    assign outputs[471] = layer6_outputs[4089];
    assign outputs[472] = ~(layer6_outputs[127]);
    assign outputs[473] = layer6_outputs[1320];
    assign outputs[474] = layer6_outputs[2285];
    assign outputs[475] = layer6_outputs[639];
    assign outputs[476] = ~((layer6_outputs[3687]) ^ (layer6_outputs[3788]));
    assign outputs[477] = ~(layer6_outputs[4288]);
    assign outputs[478] = (layer6_outputs[1825]) & ~(layer6_outputs[961]);
    assign outputs[479] = layer6_outputs[820];
    assign outputs[480] = layer6_outputs[1525];
    assign outputs[481] = layer6_outputs[115];
    assign outputs[482] = (layer6_outputs[2789]) ^ (layer6_outputs[5027]);
    assign outputs[483] = layer6_outputs[1332];
    assign outputs[484] = ~(layer6_outputs[2947]);
    assign outputs[485] = layer6_outputs[1577];
    assign outputs[486] = (layer6_outputs[2475]) ^ (layer6_outputs[1352]);
    assign outputs[487] = (layer6_outputs[2344]) & ~(layer6_outputs[4721]);
    assign outputs[488] = layer6_outputs[3900];
    assign outputs[489] = ~((layer6_outputs[1222]) ^ (layer6_outputs[4409]));
    assign outputs[490] = ~(layer6_outputs[228]) | (layer6_outputs[3188]);
    assign outputs[491] = layer6_outputs[2551];
    assign outputs[492] = layer6_outputs[3390];
    assign outputs[493] = ~(layer6_outputs[4506]);
    assign outputs[494] = ~(layer6_outputs[4214]);
    assign outputs[495] = (layer6_outputs[2428]) & (layer6_outputs[1743]);
    assign outputs[496] = layer6_outputs[2828];
    assign outputs[497] = layer6_outputs[749];
    assign outputs[498] = (layer6_outputs[4627]) & (layer6_outputs[1577]);
    assign outputs[499] = ~((layer6_outputs[3196]) ^ (layer6_outputs[3595]));
    assign outputs[500] = ~(layer6_outputs[4217]);
    assign outputs[501] = layer6_outputs[255];
    assign outputs[502] = ~((layer6_outputs[3131]) & (layer6_outputs[3006]));
    assign outputs[503] = (layer6_outputs[1236]) ^ (layer6_outputs[4966]);
    assign outputs[504] = (layer6_outputs[134]) ^ (layer6_outputs[500]);
    assign outputs[505] = ~(layer6_outputs[2879]);
    assign outputs[506] = ~(layer6_outputs[1025]);
    assign outputs[507] = ~(layer6_outputs[2922]);
    assign outputs[508] = layer6_outputs[4276];
    assign outputs[509] = layer6_outputs[2276];
    assign outputs[510] = (layer6_outputs[3824]) & ~(layer6_outputs[4608]);
    assign outputs[511] = ~(layer6_outputs[1916]) | (layer6_outputs[1063]);
    assign outputs[512] = ~(layer6_outputs[3654]);
    assign outputs[513] = (layer6_outputs[2379]) & ~(layer6_outputs[4969]);
    assign outputs[514] = (layer6_outputs[2905]) & ~(layer6_outputs[2206]);
    assign outputs[515] = ~(layer6_outputs[2755]) | (layer6_outputs[225]);
    assign outputs[516] = layer6_outputs[53];
    assign outputs[517] = layer6_outputs[1262];
    assign outputs[518] = layer6_outputs[1330];
    assign outputs[519] = ~(layer6_outputs[4421]);
    assign outputs[520] = layer6_outputs[3805];
    assign outputs[521] = (layer6_outputs[1184]) & ~(layer6_outputs[1017]);
    assign outputs[522] = ~(layer6_outputs[2456]);
    assign outputs[523] = ~(layer6_outputs[2930]);
    assign outputs[524] = layer6_outputs[3428];
    assign outputs[525] = ~(layer6_outputs[2245]);
    assign outputs[526] = ~(layer6_outputs[1055]);
    assign outputs[527] = ~(layer6_outputs[4671]);
    assign outputs[528] = layer6_outputs[3878];
    assign outputs[529] = ~(layer6_outputs[776]);
    assign outputs[530] = (layer6_outputs[2484]) ^ (layer6_outputs[176]);
    assign outputs[531] = ~(layer6_outputs[2978]);
    assign outputs[532] = 1'b0;
    assign outputs[533] = (layer6_outputs[1943]) & ~(layer6_outputs[4771]);
    assign outputs[534] = ~(layer6_outputs[1160]);
    assign outputs[535] = layer6_outputs[1223];
    assign outputs[536] = ~(layer6_outputs[1806]);
    assign outputs[537] = ~(layer6_outputs[851]);
    assign outputs[538] = ~((layer6_outputs[4664]) ^ (layer6_outputs[1675]));
    assign outputs[539] = (layer6_outputs[2311]) & ~(layer6_outputs[2427]);
    assign outputs[540] = ~(layer6_outputs[3768]);
    assign outputs[541] = (layer6_outputs[1423]) ^ (layer6_outputs[3252]);
    assign outputs[542] = ~(layer6_outputs[279]);
    assign outputs[543] = ~(layer6_outputs[1726]);
    assign outputs[544] = layer6_outputs[3325];
    assign outputs[545] = ~(layer6_outputs[4130]);
    assign outputs[546] = layer6_outputs[3302];
    assign outputs[547] = layer6_outputs[361];
    assign outputs[548] = ~(layer6_outputs[4257]);
    assign outputs[549] = layer6_outputs[4071];
    assign outputs[550] = ~(layer6_outputs[4584]);
    assign outputs[551] = ~(layer6_outputs[1009]);
    assign outputs[552] = layer6_outputs[4991];
    assign outputs[553] = ~(layer6_outputs[3326]);
    assign outputs[554] = ~(layer6_outputs[967]);
    assign outputs[555] = layer6_outputs[2253];
    assign outputs[556] = ~(layer6_outputs[3065]);
    assign outputs[557] = ~(layer6_outputs[4874]);
    assign outputs[558] = ~((layer6_outputs[439]) ^ (layer6_outputs[128]));
    assign outputs[559] = (layer6_outputs[4114]) & ~(layer6_outputs[1104]);
    assign outputs[560] = ~(layer6_outputs[3023]);
    assign outputs[561] = layer6_outputs[219];
    assign outputs[562] = ~(layer6_outputs[2415]) | (layer6_outputs[459]);
    assign outputs[563] = (layer6_outputs[4979]) & (layer6_outputs[2627]);
    assign outputs[564] = ~(layer6_outputs[4308]);
    assign outputs[565] = ~((layer6_outputs[1381]) ^ (layer6_outputs[1505]));
    assign outputs[566] = (layer6_outputs[3170]) ^ (layer6_outputs[3754]);
    assign outputs[567] = (layer6_outputs[238]) & ~(layer6_outputs[1756]);
    assign outputs[568] = ~(layer6_outputs[3616]);
    assign outputs[569] = (layer6_outputs[4435]) & (layer6_outputs[1930]);
    assign outputs[570] = ~((layer6_outputs[3149]) ^ (layer6_outputs[1731]));
    assign outputs[571] = ~(layer6_outputs[4432]);
    assign outputs[572] = (layer6_outputs[3354]) & ~(layer6_outputs[2699]);
    assign outputs[573] = ~(layer6_outputs[3699]);
    assign outputs[574] = (layer6_outputs[1293]) & (layer6_outputs[818]);
    assign outputs[575] = ~((layer6_outputs[204]) | (layer6_outputs[2978]));
    assign outputs[576] = ~(layer6_outputs[279]);
    assign outputs[577] = layer6_outputs[3571];
    assign outputs[578] = layer6_outputs[2250];
    assign outputs[579] = ~(layer6_outputs[4386]);
    assign outputs[580] = layer6_outputs[2448];
    assign outputs[581] = ~(layer6_outputs[3935]);
    assign outputs[582] = layer6_outputs[1117];
    assign outputs[583] = ~(layer6_outputs[1561]);
    assign outputs[584] = layer6_outputs[4321];
    assign outputs[585] = ~(layer6_outputs[246]);
    assign outputs[586] = ~((layer6_outputs[3627]) ^ (layer6_outputs[1130]));
    assign outputs[587] = ~(layer6_outputs[4420]) | (layer6_outputs[1409]);
    assign outputs[588] = ~((layer6_outputs[232]) ^ (layer6_outputs[2557]));
    assign outputs[589] = (layer6_outputs[5096]) & (layer6_outputs[487]);
    assign outputs[590] = ~((layer6_outputs[116]) | (layer6_outputs[1837]));
    assign outputs[591] = layer6_outputs[864];
    assign outputs[592] = ~(layer6_outputs[4186]);
    assign outputs[593] = ~(layer6_outputs[1112]);
    assign outputs[594] = (layer6_outputs[2238]) ^ (layer6_outputs[802]);
    assign outputs[595] = ~((layer6_outputs[153]) ^ (layer6_outputs[4698]));
    assign outputs[596] = (layer6_outputs[5008]) & ~(layer6_outputs[3002]);
    assign outputs[597] = layer6_outputs[3130];
    assign outputs[598] = ~((layer6_outputs[1276]) | (layer6_outputs[2821]));
    assign outputs[599] = ~(layer6_outputs[763]);
    assign outputs[600] = layer6_outputs[1719];
    assign outputs[601] = ~(layer6_outputs[1731]);
    assign outputs[602] = (layer6_outputs[111]) & ~(layer6_outputs[1144]);
    assign outputs[603] = ~((layer6_outputs[1867]) | (layer6_outputs[2910]));
    assign outputs[604] = layer6_outputs[4728];
    assign outputs[605] = ~(layer6_outputs[4976]);
    assign outputs[606] = (layer6_outputs[1974]) & ~(layer6_outputs[1532]);
    assign outputs[607] = ~(layer6_outputs[1277]);
    assign outputs[608] = layer6_outputs[576];
    assign outputs[609] = ~(layer6_outputs[1230]);
    assign outputs[610] = (layer6_outputs[2367]) & ~(layer6_outputs[4505]);
    assign outputs[611] = (layer6_outputs[5010]) ^ (layer6_outputs[2042]);
    assign outputs[612] = ~((layer6_outputs[4846]) | (layer6_outputs[3039]));
    assign outputs[613] = ~((layer6_outputs[2680]) ^ (layer6_outputs[2597]));
    assign outputs[614] = ~(layer6_outputs[4996]) | (layer6_outputs[3733]);
    assign outputs[615] = layer6_outputs[1670];
    assign outputs[616] = ~((layer6_outputs[3145]) ^ (layer6_outputs[213]));
    assign outputs[617] = ~(layer6_outputs[3304]);
    assign outputs[618] = layer6_outputs[1786];
    assign outputs[619] = (layer6_outputs[1105]) ^ (layer6_outputs[4987]);
    assign outputs[620] = layer6_outputs[3388];
    assign outputs[621] = layer6_outputs[4093];
    assign outputs[622] = ~((layer6_outputs[3687]) ^ (layer6_outputs[875]));
    assign outputs[623] = ~(layer6_outputs[2157]);
    assign outputs[624] = layer6_outputs[3454];
    assign outputs[625] = ~(layer6_outputs[3752]);
    assign outputs[626] = layer6_outputs[300];
    assign outputs[627] = (layer6_outputs[2091]) & (layer6_outputs[3159]);
    assign outputs[628] = layer6_outputs[2571];
    assign outputs[629] = ~(layer6_outputs[1394]);
    assign outputs[630] = (layer6_outputs[4850]) ^ (layer6_outputs[3470]);
    assign outputs[631] = layer6_outputs[1668];
    assign outputs[632] = layer6_outputs[2772];
    assign outputs[633] = ~(layer6_outputs[278]);
    assign outputs[634] = layer6_outputs[2902];
    assign outputs[635] = ~(layer6_outputs[3988]);
    assign outputs[636] = ~(layer6_outputs[2317]);
    assign outputs[637] = (layer6_outputs[2422]) ^ (layer6_outputs[3498]);
    assign outputs[638] = ~(layer6_outputs[4165]);
    assign outputs[639] = (layer6_outputs[4623]) ^ (layer6_outputs[3305]);
    assign outputs[640] = layer6_outputs[1470];
    assign outputs[641] = (layer6_outputs[1675]) ^ (layer6_outputs[254]);
    assign outputs[642] = (layer6_outputs[3347]) & ~(layer6_outputs[4858]);
    assign outputs[643] = ~(layer6_outputs[2057]);
    assign outputs[644] = ~((layer6_outputs[4867]) | (layer6_outputs[3019]));
    assign outputs[645] = ~(layer6_outputs[4693]);
    assign outputs[646] = ~((layer6_outputs[3246]) ^ (layer6_outputs[2790]));
    assign outputs[647] = ~(layer6_outputs[4358]);
    assign outputs[648] = ~((layer6_outputs[3778]) | (layer6_outputs[1270]));
    assign outputs[649] = ~((layer6_outputs[1860]) ^ (layer6_outputs[3305]));
    assign outputs[650] = layer6_outputs[4273];
    assign outputs[651] = layer6_outputs[2961];
    assign outputs[652] = ~(layer6_outputs[3233]);
    assign outputs[653] = ~(layer6_outputs[595]) | (layer6_outputs[1078]);
    assign outputs[654] = layer6_outputs[5118];
    assign outputs[655] = ~(layer6_outputs[832]);
    assign outputs[656] = ~(layer6_outputs[489]);
    assign outputs[657] = ~(layer6_outputs[165]);
    assign outputs[658] = (layer6_outputs[414]) & ~(layer6_outputs[1497]);
    assign outputs[659] = ~(layer6_outputs[1011]);
    assign outputs[660] = (layer6_outputs[3349]) ^ (layer6_outputs[3419]);
    assign outputs[661] = ~(layer6_outputs[2977]);
    assign outputs[662] = layer6_outputs[25];
    assign outputs[663] = (layer6_outputs[4583]) ^ (layer6_outputs[2871]);
    assign outputs[664] = layer6_outputs[3743];
    assign outputs[665] = layer6_outputs[1925];
    assign outputs[666] = (layer6_outputs[4613]) & (layer6_outputs[1142]);
    assign outputs[667] = layer6_outputs[1631];
    assign outputs[668] = layer6_outputs[3494];
    assign outputs[669] = layer6_outputs[3534];
    assign outputs[670] = ~((layer6_outputs[4708]) | (layer6_outputs[4023]));
    assign outputs[671] = layer6_outputs[2492];
    assign outputs[672] = (layer6_outputs[2330]) & ~(layer6_outputs[1635]);
    assign outputs[673] = (layer6_outputs[654]) & (layer6_outputs[4779]);
    assign outputs[674] = layer6_outputs[656];
    assign outputs[675] = (layer6_outputs[102]) & (layer6_outputs[4318]);
    assign outputs[676] = ~(layer6_outputs[2366]);
    assign outputs[677] = ~(layer6_outputs[258]);
    assign outputs[678] = (layer6_outputs[1624]) ^ (layer6_outputs[598]);
    assign outputs[679] = ~((layer6_outputs[1093]) | (layer6_outputs[4707]));
    assign outputs[680] = (layer6_outputs[5104]) & ~(layer6_outputs[3628]);
    assign outputs[681] = ~((layer6_outputs[1400]) ^ (layer6_outputs[139]));
    assign outputs[682] = layer6_outputs[988];
    assign outputs[683] = (layer6_outputs[3859]) ^ (layer6_outputs[3686]);
    assign outputs[684] = ~(layer6_outputs[1379]);
    assign outputs[685] = layer6_outputs[2266];
    assign outputs[686] = ~(layer6_outputs[4415]);
    assign outputs[687] = ~(layer6_outputs[2006]);
    assign outputs[688] = layer6_outputs[4826];
    assign outputs[689] = ~(layer6_outputs[3728]);
    assign outputs[690] = layer6_outputs[3836];
    assign outputs[691] = ~(layer6_outputs[4493]);
    assign outputs[692] = (layer6_outputs[844]) & ~(layer6_outputs[2020]);
    assign outputs[693] = ~(layer6_outputs[3076]) | (layer6_outputs[2444]);
    assign outputs[694] = layer6_outputs[610];
    assign outputs[695] = ~((layer6_outputs[4757]) | (layer6_outputs[438]));
    assign outputs[696] = ~((layer6_outputs[1477]) | (layer6_outputs[17]));
    assign outputs[697] = layer6_outputs[2184];
    assign outputs[698] = ~(layer6_outputs[1190]);
    assign outputs[699] = (layer6_outputs[1169]) ^ (layer6_outputs[2361]);
    assign outputs[700] = ~(layer6_outputs[3823]);
    assign outputs[701] = (layer6_outputs[2356]) ^ (layer6_outputs[2039]);
    assign outputs[702] = (layer6_outputs[1376]) & (layer6_outputs[1046]);
    assign outputs[703] = (layer6_outputs[15]) & ~(layer6_outputs[2381]);
    assign outputs[704] = layer6_outputs[4783];
    assign outputs[705] = ~((layer6_outputs[4976]) ^ (layer6_outputs[4734]));
    assign outputs[706] = layer6_outputs[4615];
    assign outputs[707] = layer6_outputs[1275];
    assign outputs[708] = layer6_outputs[3956];
    assign outputs[709] = (layer6_outputs[2785]) ^ (layer6_outputs[5047]);
    assign outputs[710] = (layer6_outputs[1501]) ^ (layer6_outputs[2009]);
    assign outputs[711] = (layer6_outputs[2909]) ^ (layer6_outputs[880]);
    assign outputs[712] = layer6_outputs[3089];
    assign outputs[713] = (layer6_outputs[601]) & ~(layer6_outputs[4605]);
    assign outputs[714] = ~(layer6_outputs[2359]) | (layer6_outputs[2147]);
    assign outputs[715] = layer6_outputs[2763];
    assign outputs[716] = ~(layer6_outputs[2620]);
    assign outputs[717] = ~(layer6_outputs[4497]);
    assign outputs[718] = ~((layer6_outputs[1648]) | (layer6_outputs[2336]));
    assign outputs[719] = (layer6_outputs[1333]) & (layer6_outputs[1430]);
    assign outputs[720] = ~(layer6_outputs[1418]) | (layer6_outputs[1020]);
    assign outputs[721] = (layer6_outputs[4758]) ^ (layer6_outputs[3783]);
    assign outputs[722] = ~(layer6_outputs[4035]);
    assign outputs[723] = (layer6_outputs[1910]) & (layer6_outputs[728]);
    assign outputs[724] = ~((layer6_outputs[945]) | (layer6_outputs[3031]));
    assign outputs[725] = ~(layer6_outputs[4066]);
    assign outputs[726] = layer6_outputs[811];
    assign outputs[727] = ~(layer6_outputs[4452]) | (layer6_outputs[2312]);
    assign outputs[728] = layer6_outputs[2935];
    assign outputs[729] = (layer6_outputs[150]) & ~(layer6_outputs[2609]);
    assign outputs[730] = layer6_outputs[4310];
    assign outputs[731] = ~((layer6_outputs[1863]) ^ (layer6_outputs[4467]));
    assign outputs[732] = ~((layer6_outputs[4558]) ^ (layer6_outputs[3426]));
    assign outputs[733] = layer6_outputs[3874];
    assign outputs[734] = layer6_outputs[3193];
    assign outputs[735] = ~(layer6_outputs[4453]);
    assign outputs[736] = ~((layer6_outputs[3487]) ^ (layer6_outputs[2895]));
    assign outputs[737] = (layer6_outputs[1386]) ^ (layer6_outputs[3236]);
    assign outputs[738] = ~(layer6_outputs[4564]);
    assign outputs[739] = ~((layer6_outputs[2911]) ^ (layer6_outputs[754]));
    assign outputs[740] = layer6_outputs[3751];
    assign outputs[741] = layer6_outputs[432];
    assign outputs[742] = ~(layer6_outputs[3851]);
    assign outputs[743] = ~((layer6_outputs[47]) ^ (layer6_outputs[4970]));
    assign outputs[744] = ~(layer6_outputs[3362]);
    assign outputs[745] = ~((layer6_outputs[1854]) | (layer6_outputs[1679]));
    assign outputs[746] = ~((layer6_outputs[3789]) | (layer6_outputs[6]));
    assign outputs[747] = (layer6_outputs[3688]) & (layer6_outputs[3003]);
    assign outputs[748] = ~(layer6_outputs[1436]);
    assign outputs[749] = ~((layer6_outputs[3333]) | (layer6_outputs[3198]));
    assign outputs[750] = ~((layer6_outputs[56]) | (layer6_outputs[4701]));
    assign outputs[751] = (layer6_outputs[4540]) & ~(layer6_outputs[3270]);
    assign outputs[752] = ~(layer6_outputs[1206]);
    assign outputs[753] = layer6_outputs[3172];
    assign outputs[754] = ~((layer6_outputs[3387]) | (layer6_outputs[2274]));
    assign outputs[755] = ~(layer6_outputs[1245]);
    assign outputs[756] = (layer6_outputs[3494]) & (layer6_outputs[3591]);
    assign outputs[757] = ~((layer6_outputs[4961]) & (layer6_outputs[900]));
    assign outputs[758] = layer6_outputs[2451];
    assign outputs[759] = ~((layer6_outputs[1559]) ^ (layer6_outputs[3087]));
    assign outputs[760] = layer6_outputs[1001];
    assign outputs[761] = ~(layer6_outputs[4083]);
    assign outputs[762] = ~((layer6_outputs[2505]) ^ (layer6_outputs[1986]));
    assign outputs[763] = ~(layer6_outputs[3911]);
    assign outputs[764] = ~(layer6_outputs[1883]);
    assign outputs[765] = layer6_outputs[4760];
    assign outputs[766] = ~(layer6_outputs[2485]);
    assign outputs[767] = (layer6_outputs[1451]) & (layer6_outputs[218]);
    assign outputs[768] = (layer6_outputs[2467]) & (layer6_outputs[3886]);
    assign outputs[769] = layer6_outputs[2266];
    assign outputs[770] = ~(layer6_outputs[1741]) | (layer6_outputs[2096]);
    assign outputs[771] = ~(layer6_outputs[4521]);
    assign outputs[772] = (layer6_outputs[1827]) & ~(layer6_outputs[1128]);
    assign outputs[773] = (layer6_outputs[3905]) & (layer6_outputs[4159]);
    assign outputs[774] = (layer6_outputs[4748]) ^ (layer6_outputs[3938]);
    assign outputs[775] = ~(layer6_outputs[243]);
    assign outputs[776] = ~((layer6_outputs[4703]) | (layer6_outputs[3453]));
    assign outputs[777] = (layer6_outputs[3060]) & (layer6_outputs[4654]);
    assign outputs[778] = ~(layer6_outputs[4379]);
    assign outputs[779] = (layer6_outputs[176]) ^ (layer6_outputs[1692]);
    assign outputs[780] = ~(layer6_outputs[3005]);
    assign outputs[781] = ~((layer6_outputs[4424]) ^ (layer6_outputs[3697]));
    assign outputs[782] = ~(layer6_outputs[2145]);
    assign outputs[783] = ~(layer6_outputs[541]);
    assign outputs[784] = ~(layer6_outputs[721]);
    assign outputs[785] = (layer6_outputs[4514]) ^ (layer6_outputs[2231]);
    assign outputs[786] = ~(layer6_outputs[2908]);
    assign outputs[787] = layer6_outputs[1610];
    assign outputs[788] = layer6_outputs[2064];
    assign outputs[789] = layer6_outputs[4077];
    assign outputs[790] = ~((layer6_outputs[3741]) ^ (layer6_outputs[3055]));
    assign outputs[791] = ~((layer6_outputs[4925]) ^ (layer6_outputs[1951]));
    assign outputs[792] = ~(layer6_outputs[3611]);
    assign outputs[793] = layer6_outputs[1665];
    assign outputs[794] = (layer6_outputs[900]) & ~(layer6_outputs[502]);
    assign outputs[795] = layer6_outputs[2562];
    assign outputs[796] = ~((layer6_outputs[1935]) | (layer6_outputs[4707]));
    assign outputs[797] = ~(layer6_outputs[3198]) | (layer6_outputs[1533]);
    assign outputs[798] = layer6_outputs[604];
    assign outputs[799] = ~(layer6_outputs[4796]);
    assign outputs[800] = ~(layer6_outputs[3073]);
    assign outputs[801] = (layer6_outputs[4305]) & (layer6_outputs[510]);
    assign outputs[802] = layer6_outputs[5114];
    assign outputs[803] = layer6_outputs[1472];
    assign outputs[804] = ~(layer6_outputs[3116]);
    assign outputs[805] = ~(layer6_outputs[347]);
    assign outputs[806] = ~((layer6_outputs[4286]) ^ (layer6_outputs[1329]));
    assign outputs[807] = (layer6_outputs[3297]) & ~(layer6_outputs[368]);
    assign outputs[808] = (layer6_outputs[3882]) & ~(layer6_outputs[1170]);
    assign outputs[809] = ~(layer6_outputs[4464]);
    assign outputs[810] = layer6_outputs[1895];
    assign outputs[811] = ~(layer6_outputs[5085]);
    assign outputs[812] = (layer6_outputs[1795]) & ~(layer6_outputs[4241]);
    assign outputs[813] = ~(layer6_outputs[1537]);
    assign outputs[814] = layer6_outputs[1259];
    assign outputs[815] = ~(layer6_outputs[3064]);
    assign outputs[816] = ~((layer6_outputs[4621]) | (layer6_outputs[2264]));
    assign outputs[817] = layer6_outputs[3462];
    assign outputs[818] = layer6_outputs[54];
    assign outputs[819] = layer6_outputs[4340];
    assign outputs[820] = (layer6_outputs[4253]) & ~(layer6_outputs[2758]);
    assign outputs[821] = (layer6_outputs[4938]) & (layer6_outputs[2247]);
    assign outputs[822] = ~(layer6_outputs[2148]);
    assign outputs[823] = ~(layer6_outputs[1893]);
    assign outputs[824] = ~(layer6_outputs[3312]);
    assign outputs[825] = ~(layer6_outputs[4454]);
    assign outputs[826] = ~(layer6_outputs[3023]);
    assign outputs[827] = layer6_outputs[2798];
    assign outputs[828] = ~((layer6_outputs[3509]) | (layer6_outputs[2428]));
    assign outputs[829] = ~(layer6_outputs[4732]);
    assign outputs[830] = ~((layer6_outputs[1006]) ^ (layer6_outputs[4129]));
    assign outputs[831] = (layer6_outputs[4946]) & (layer6_outputs[3225]);
    assign outputs[832] = (layer6_outputs[2120]) & ~(layer6_outputs[191]);
    assign outputs[833] = (layer6_outputs[2339]) ^ (layer6_outputs[1825]);
    assign outputs[834] = (layer6_outputs[436]) | (layer6_outputs[3210]);
    assign outputs[835] = layer6_outputs[3273];
    assign outputs[836] = layer6_outputs[2289];
    assign outputs[837] = (layer6_outputs[4552]) & ~(layer6_outputs[5041]);
    assign outputs[838] = layer6_outputs[591];
    assign outputs[839] = layer6_outputs[121];
    assign outputs[840] = ~(layer6_outputs[5047]);
    assign outputs[841] = (layer6_outputs[5002]) & ~(layer6_outputs[4422]);
    assign outputs[842] = ~(layer6_outputs[3312]);
    assign outputs[843] = layer6_outputs[3597];
    assign outputs[844] = ~(layer6_outputs[4810]);
    assign outputs[845] = ~(layer6_outputs[2890]);
    assign outputs[846] = layer6_outputs[1208];
    assign outputs[847] = ~(layer6_outputs[3652]);
    assign outputs[848] = ~(layer6_outputs[3337]);
    assign outputs[849] = (layer6_outputs[2668]) & ~(layer6_outputs[1149]);
    assign outputs[850] = ~((layer6_outputs[1022]) | (layer6_outputs[3418]));
    assign outputs[851] = (layer6_outputs[3662]) & ~(layer6_outputs[3525]);
    assign outputs[852] = (layer6_outputs[1803]) ^ (layer6_outputs[2147]);
    assign outputs[853] = ~(layer6_outputs[4417]);
    assign outputs[854] = ~(layer6_outputs[1761]);
    assign outputs[855] = layer6_outputs[1354];
    assign outputs[856] = ~(layer6_outputs[4509]);
    assign outputs[857] = ~(layer6_outputs[3284]);
    assign outputs[858] = layer6_outputs[123];
    assign outputs[859] = layer6_outputs[4460];
    assign outputs[860] = layer6_outputs[3334];
    assign outputs[861] = (layer6_outputs[4855]) & ~(layer6_outputs[3438]);
    assign outputs[862] = ~(layer6_outputs[3672]);
    assign outputs[863] = ~(layer6_outputs[602]);
    assign outputs[864] = ~((layer6_outputs[2980]) ^ (layer6_outputs[477]));
    assign outputs[865] = layer6_outputs[4478];
    assign outputs[866] = layer6_outputs[2784];
    assign outputs[867] = ~(layer6_outputs[330]);
    assign outputs[868] = (layer6_outputs[2971]) & (layer6_outputs[352]);
    assign outputs[869] = ~((layer6_outputs[719]) | (layer6_outputs[1567]));
    assign outputs[870] = ~((layer6_outputs[4624]) | (layer6_outputs[3033]));
    assign outputs[871] = (layer6_outputs[3692]) & ~(layer6_outputs[3697]);
    assign outputs[872] = ~(layer6_outputs[3679]);
    assign outputs[873] = (layer6_outputs[4445]) & ~(layer6_outputs[2555]);
    assign outputs[874] = ~(layer6_outputs[3166]);
    assign outputs[875] = (layer6_outputs[944]) ^ (layer6_outputs[1008]);
    assign outputs[876] = ~(layer6_outputs[3511]);
    assign outputs[877] = ~(layer6_outputs[2326]) | (layer6_outputs[2331]);
    assign outputs[878] = ~((layer6_outputs[2123]) ^ (layer6_outputs[4237]));
    assign outputs[879] = layer6_outputs[3000];
    assign outputs[880] = ~((layer6_outputs[1218]) ^ (layer6_outputs[2439]));
    assign outputs[881] = ~(layer6_outputs[310]);
    assign outputs[882] = ~(layer6_outputs[1733]);
    assign outputs[883] = layer6_outputs[4543];
    assign outputs[884] = ~(layer6_outputs[3711]);
    assign outputs[885] = ~(layer6_outputs[905]);
    assign outputs[886] = ~(layer6_outputs[302]);
    assign outputs[887] = (layer6_outputs[216]) & ~(layer6_outputs[2695]);
    assign outputs[888] = ~(layer6_outputs[2313]);
    assign outputs[889] = (layer6_outputs[3255]) & ~(layer6_outputs[1637]);
    assign outputs[890] = layer6_outputs[3085];
    assign outputs[891] = (layer6_outputs[3694]) & ~(layer6_outputs[616]);
    assign outputs[892] = ~(layer6_outputs[3731]);
    assign outputs[893] = ~(layer6_outputs[742]);
    assign outputs[894] = layer6_outputs[3879];
    assign outputs[895] = layer6_outputs[4065];
    assign outputs[896] = (layer6_outputs[2526]) & ~(layer6_outputs[2436]);
    assign outputs[897] = layer6_outputs[1351];
    assign outputs[898] = layer6_outputs[2527];
    assign outputs[899] = ~((layer6_outputs[2582]) ^ (layer6_outputs[5101]));
    assign outputs[900] = ~((layer6_outputs[3214]) ^ (layer6_outputs[3920]));
    assign outputs[901] = layer6_outputs[1888];
    assign outputs[902] = ~((layer6_outputs[873]) ^ (layer6_outputs[1137]));
    assign outputs[903] = layer6_outputs[1863];
    assign outputs[904] = ~(layer6_outputs[1836]);
    assign outputs[905] = (layer6_outputs[595]) & (layer6_outputs[1075]);
    assign outputs[906] = ~((layer6_outputs[5007]) ^ (layer6_outputs[3958]));
    assign outputs[907] = ~(layer6_outputs[3650]);
    assign outputs[908] = (layer6_outputs[4034]) & ~(layer6_outputs[4316]);
    assign outputs[909] = layer6_outputs[4974];
    assign outputs[910] = (layer6_outputs[895]) & (layer6_outputs[747]);
    assign outputs[911] = ~((layer6_outputs[3143]) | (layer6_outputs[4353]));
    assign outputs[912] = layer6_outputs[3370];
    assign outputs[913] = ~(layer6_outputs[80]);
    assign outputs[914] = layer6_outputs[1140];
    assign outputs[915] = (layer6_outputs[2761]) ^ (layer6_outputs[1280]);
    assign outputs[916] = ~(layer6_outputs[2268]);
    assign outputs[917] = (layer6_outputs[2801]) & ~(layer6_outputs[3997]);
    assign outputs[918] = ~(layer6_outputs[3314]);
    assign outputs[919] = ~(layer6_outputs[1450]);
    assign outputs[920] = (layer6_outputs[3009]) & ~(layer6_outputs[640]);
    assign outputs[921] = (layer6_outputs[2884]) ^ (layer6_outputs[5082]);
    assign outputs[922] = (layer6_outputs[4604]) & (layer6_outputs[4307]);
    assign outputs[923] = layer6_outputs[3755];
    assign outputs[924] = (layer6_outputs[2343]) & ~(layer6_outputs[776]);
    assign outputs[925] = layer6_outputs[3296];
    assign outputs[926] = ~(layer6_outputs[2725]);
    assign outputs[927] = ~(layer6_outputs[1503]);
    assign outputs[928] = ~((layer6_outputs[1861]) | (layer6_outputs[118]));
    assign outputs[929] = (layer6_outputs[4134]) & (layer6_outputs[1033]);
    assign outputs[930] = layer6_outputs[4482];
    assign outputs[931] = (layer6_outputs[427]) & ~(layer6_outputs[489]);
    assign outputs[932] = (layer6_outputs[3170]) ^ (layer6_outputs[1120]);
    assign outputs[933] = layer6_outputs[3949];
    assign outputs[934] = (layer6_outputs[436]) ^ (layer6_outputs[4531]);
    assign outputs[935] = ~(layer6_outputs[4343]);
    assign outputs[936] = layer6_outputs[393];
    assign outputs[937] = ~((layer6_outputs[2249]) ^ (layer6_outputs[4517]));
    assign outputs[938] = layer6_outputs[1119];
    assign outputs[939] = layer6_outputs[4761];
    assign outputs[940] = ~(layer6_outputs[502]) | (layer6_outputs[3612]);
    assign outputs[941] = ~(layer6_outputs[1228]);
    assign outputs[942] = layer6_outputs[4473];
    assign outputs[943] = layer6_outputs[4897];
    assign outputs[944] = ~(layer6_outputs[3531]);
    assign outputs[945] = (layer6_outputs[3179]) ^ (layer6_outputs[4556]);
    assign outputs[946] = layer6_outputs[3516];
    assign outputs[947] = (layer6_outputs[2689]) & ~(layer6_outputs[1386]);
    assign outputs[948] = ~(layer6_outputs[5094]);
    assign outputs[949] = layer6_outputs[2840];
    assign outputs[950] = ~(layer6_outputs[1710]);
    assign outputs[951] = ~((layer6_outputs[4902]) | (layer6_outputs[1521]));
    assign outputs[952] = layer6_outputs[1440];
    assign outputs[953] = ~(layer6_outputs[877]);
    assign outputs[954] = ~(layer6_outputs[291]) | (layer6_outputs[5089]);
    assign outputs[955] = layer6_outputs[5002];
    assign outputs[956] = layer6_outputs[864];
    assign outputs[957] = layer6_outputs[3340];
    assign outputs[958] = ~(layer6_outputs[3500]);
    assign outputs[959] = layer6_outputs[724];
    assign outputs[960] = (layer6_outputs[750]) ^ (layer6_outputs[2702]);
    assign outputs[961] = ~(layer6_outputs[412]);
    assign outputs[962] = ~(layer6_outputs[3668]);
    assign outputs[963] = layer6_outputs[1239];
    assign outputs[964] = (layer6_outputs[630]) & (layer6_outputs[311]);
    assign outputs[965] = (layer6_outputs[4982]) & ~(layer6_outputs[3543]);
    assign outputs[966] = (layer6_outputs[1769]) | (layer6_outputs[629]);
    assign outputs[967] = layer6_outputs[1262];
    assign outputs[968] = ~(layer6_outputs[2411]);
    assign outputs[969] = (layer6_outputs[1198]) & (layer6_outputs[2129]);
    assign outputs[970] = (layer6_outputs[2787]) & ~(layer6_outputs[1711]);
    assign outputs[971] = ~((layer6_outputs[1264]) | (layer6_outputs[910]));
    assign outputs[972] = layer6_outputs[4821];
    assign outputs[973] = layer6_outputs[3069];
    assign outputs[974] = layer6_outputs[2149];
    assign outputs[975] = ~(layer6_outputs[3205]) | (layer6_outputs[1898]);
    assign outputs[976] = layer6_outputs[1094];
    assign outputs[977] = ~(layer6_outputs[2736]);
    assign outputs[978] = (layer6_outputs[3556]) | (layer6_outputs[1520]);
    assign outputs[979] = (layer6_outputs[3604]) ^ (layer6_outputs[921]);
    assign outputs[980] = layer6_outputs[2536];
    assign outputs[981] = layer6_outputs[2848];
    assign outputs[982] = layer6_outputs[326];
    assign outputs[983] = (layer6_outputs[311]) & ~(layer6_outputs[3146]);
    assign outputs[984] = (layer6_outputs[1186]) ^ (layer6_outputs[4907]);
    assign outputs[985] = (layer6_outputs[2097]) & ~(layer6_outputs[2945]);
    assign outputs[986] = layer6_outputs[3283];
    assign outputs[987] = ~((layer6_outputs[2340]) | (layer6_outputs[1532]));
    assign outputs[988] = layer6_outputs[4425];
    assign outputs[989] = layer6_outputs[1831];
    assign outputs[990] = ~(layer6_outputs[2221]);
    assign outputs[991] = ~((layer6_outputs[3079]) & (layer6_outputs[3814]));
    assign outputs[992] = ~(layer6_outputs[4092]);
    assign outputs[993] = ~(layer6_outputs[2114]);
    assign outputs[994] = ~(layer6_outputs[1377]);
    assign outputs[995] = layer6_outputs[4733];
    assign outputs[996] = ~((layer6_outputs[2134]) ^ (layer6_outputs[3283]));
    assign outputs[997] = (layer6_outputs[4122]) & ~(layer6_outputs[3877]);
    assign outputs[998] = ~(layer6_outputs[1655]);
    assign outputs[999] = (layer6_outputs[769]) ^ (layer6_outputs[4275]);
    assign outputs[1000] = (layer6_outputs[3263]) & ~(layer6_outputs[4124]);
    assign outputs[1001] = ~(layer6_outputs[2016]);
    assign outputs[1002] = (layer6_outputs[3605]) & ~(layer6_outputs[3092]);
    assign outputs[1003] = layer6_outputs[5096];
    assign outputs[1004] = ~((layer6_outputs[3395]) | (layer6_outputs[4884]));
    assign outputs[1005] = (layer6_outputs[490]) & ~(layer6_outputs[5006]);
    assign outputs[1006] = ~(layer6_outputs[568]) | (layer6_outputs[3701]);
    assign outputs[1007] = (layer6_outputs[2495]) ^ (layer6_outputs[2608]);
    assign outputs[1008] = layer6_outputs[314];
    assign outputs[1009] = layer6_outputs[5022];
    assign outputs[1010] = ~((layer6_outputs[4564]) ^ (layer6_outputs[1048]));
    assign outputs[1011] = layer6_outputs[153];
    assign outputs[1012] = ~(layer6_outputs[4904]);
    assign outputs[1013] = layer6_outputs[4818];
    assign outputs[1014] = ~(layer6_outputs[4505]);
    assign outputs[1015] = (layer6_outputs[1514]) & (layer6_outputs[1549]);
    assign outputs[1016] = ~((layer6_outputs[3451]) ^ (layer6_outputs[3968]));
    assign outputs[1017] = layer6_outputs[779];
    assign outputs[1018] = (layer6_outputs[3515]) ^ (layer6_outputs[2716]);
    assign outputs[1019] = layer6_outputs[25];
    assign outputs[1020] = ~(layer6_outputs[1080]);
    assign outputs[1021] = ~((layer6_outputs[4725]) ^ (layer6_outputs[2849]));
    assign outputs[1022] = (layer6_outputs[1942]) & ~(layer6_outputs[2114]);
    assign outputs[1023] = ~((layer6_outputs[3796]) ^ (layer6_outputs[2371]));
    assign outputs[1024] = ~((layer6_outputs[631]) ^ (layer6_outputs[3765]));
    assign outputs[1025] = (layer6_outputs[3837]) ^ (layer6_outputs[3505]);
    assign outputs[1026] = layer6_outputs[49];
    assign outputs[1027] = ~(layer6_outputs[59]) | (layer6_outputs[3742]);
    assign outputs[1028] = layer6_outputs[310];
    assign outputs[1029] = layer6_outputs[638];
    assign outputs[1030] = ~((layer6_outputs[1302]) ^ (layer6_outputs[4942]));
    assign outputs[1031] = ~(layer6_outputs[4655]);
    assign outputs[1032] = ~(layer6_outputs[3399]);
    assign outputs[1033] = ~(layer6_outputs[1174]) | (layer6_outputs[252]);
    assign outputs[1034] = ~(layer6_outputs[3699]);
    assign outputs[1035] = (layer6_outputs[2478]) ^ (layer6_outputs[1746]);
    assign outputs[1036] = (layer6_outputs[1682]) ^ (layer6_outputs[4550]);
    assign outputs[1037] = layer6_outputs[3803];
    assign outputs[1038] = layer6_outputs[4322];
    assign outputs[1039] = ~((layer6_outputs[352]) ^ (layer6_outputs[3753]));
    assign outputs[1040] = (layer6_outputs[3236]) & ~(layer6_outputs[2538]);
    assign outputs[1041] = layer6_outputs[4576];
    assign outputs[1042] = ~((layer6_outputs[3531]) & (layer6_outputs[4661]));
    assign outputs[1043] = ~(layer6_outputs[2765]);
    assign outputs[1044] = ~(layer6_outputs[2671]);
    assign outputs[1045] = ~((layer6_outputs[1954]) ^ (layer6_outputs[4894]));
    assign outputs[1046] = ~(layer6_outputs[4380]);
    assign outputs[1047] = ~(layer6_outputs[4339]);
    assign outputs[1048] = ~(layer6_outputs[3451]);
    assign outputs[1049] = ~((layer6_outputs[1296]) ^ (layer6_outputs[4311]));
    assign outputs[1050] = ~(layer6_outputs[474]);
    assign outputs[1051] = ~(layer6_outputs[1687]);
    assign outputs[1052] = ~(layer6_outputs[4523]);
    assign outputs[1053] = (layer6_outputs[574]) ^ (layer6_outputs[1153]);
    assign outputs[1054] = ~((layer6_outputs[4009]) ^ (layer6_outputs[4840]));
    assign outputs[1055] = layer6_outputs[2882];
    assign outputs[1056] = (layer6_outputs[2496]) & (layer6_outputs[1281]);
    assign outputs[1057] = ~(layer6_outputs[2073]);
    assign outputs[1058] = layer6_outputs[542];
    assign outputs[1059] = ~((layer6_outputs[1326]) ^ (layer6_outputs[4736]));
    assign outputs[1060] = layer6_outputs[391];
    assign outputs[1061] = ~((layer6_outputs[4718]) & (layer6_outputs[275]));
    assign outputs[1062] = layer6_outputs[1144];
    assign outputs[1063] = layer6_outputs[215];
    assign outputs[1064] = ~(layer6_outputs[1317]);
    assign outputs[1065] = ~(layer6_outputs[681]);
    assign outputs[1066] = ~(layer6_outputs[5001]);
    assign outputs[1067] = (layer6_outputs[3855]) ^ (layer6_outputs[8]);
    assign outputs[1068] = ~(layer6_outputs[1019]);
    assign outputs[1069] = layer6_outputs[1242];
    assign outputs[1070] = layer6_outputs[1790];
    assign outputs[1071] = ~((layer6_outputs[4810]) ^ (layer6_outputs[4436]));
    assign outputs[1072] = layer6_outputs[161];
    assign outputs[1073] = ~(layer6_outputs[4518]);
    assign outputs[1074] = ~(layer6_outputs[852]);
    assign outputs[1075] = layer6_outputs[936];
    assign outputs[1076] = ~(layer6_outputs[4521]);
    assign outputs[1077] = layer6_outputs[2190];
    assign outputs[1078] = ~(layer6_outputs[239]);
    assign outputs[1079] = layer6_outputs[2286];
    assign outputs[1080] = layer6_outputs[2877];
    assign outputs[1081] = (layer6_outputs[3909]) ^ (layer6_outputs[1752]);
    assign outputs[1082] = layer6_outputs[2217];
    assign outputs[1083] = layer6_outputs[623];
    assign outputs[1084] = (layer6_outputs[720]) & ~(layer6_outputs[4037]);
    assign outputs[1085] = ~((layer6_outputs[3190]) ^ (layer6_outputs[3955]));
    assign outputs[1086] = (layer6_outputs[2024]) | (layer6_outputs[2167]);
    assign outputs[1087] = ~(layer6_outputs[4127]);
    assign outputs[1088] = (layer6_outputs[2756]) ^ (layer6_outputs[2630]);
    assign outputs[1089] = ~(layer6_outputs[906]);
    assign outputs[1090] = (layer6_outputs[1887]) ^ (layer6_outputs[4308]);
    assign outputs[1091] = layer6_outputs[4716];
    assign outputs[1092] = ~(layer6_outputs[3772]);
    assign outputs[1093] = (layer6_outputs[3848]) ^ (layer6_outputs[3011]);
    assign outputs[1094] = ~(layer6_outputs[653]);
    assign outputs[1095] = ~((layer6_outputs[192]) | (layer6_outputs[3662]));
    assign outputs[1096] = ~(layer6_outputs[1962]);
    assign outputs[1097] = ~((layer6_outputs[2142]) | (layer6_outputs[4330]));
    assign outputs[1098] = ~(layer6_outputs[2440]);
    assign outputs[1099] = ~(layer6_outputs[3618]);
    assign outputs[1100] = layer6_outputs[4323];
    assign outputs[1101] = ~(layer6_outputs[2128]);
    assign outputs[1102] = layer6_outputs[4503];
    assign outputs[1103] = ~(layer6_outputs[2972]);
    assign outputs[1104] = (layer6_outputs[3022]) & (layer6_outputs[4462]);
    assign outputs[1105] = layer6_outputs[2894];
    assign outputs[1106] = layer6_outputs[2497];
    assign outputs[1107] = layer6_outputs[1414];
    assign outputs[1108] = ~((layer6_outputs[4642]) ^ (layer6_outputs[503]));
    assign outputs[1109] = ~(layer6_outputs[17]);
    assign outputs[1110] = ~(layer6_outputs[3769]);
    assign outputs[1111] = ~((layer6_outputs[2246]) | (layer6_outputs[3157]));
    assign outputs[1112] = ~(layer6_outputs[2063]);
    assign outputs[1113] = ~(layer6_outputs[313]);
    assign outputs[1114] = ~(layer6_outputs[70]) | (layer6_outputs[2443]);
    assign outputs[1115] = ~(layer6_outputs[934]);
    assign outputs[1116] = ~((layer6_outputs[4930]) ^ (layer6_outputs[654]));
    assign outputs[1117] = layer6_outputs[5103];
    assign outputs[1118] = (layer6_outputs[3495]) & ~(layer6_outputs[4872]);
    assign outputs[1119] = ~((layer6_outputs[846]) & (layer6_outputs[4036]));
    assign outputs[1120] = ~(layer6_outputs[4378]);
    assign outputs[1121] = layer6_outputs[4282];
    assign outputs[1122] = layer6_outputs[4914];
    assign outputs[1123] = layer6_outputs[3270];
    assign outputs[1124] = layer6_outputs[4171];
    assign outputs[1125] = ~((layer6_outputs[808]) | (layer6_outputs[2964]));
    assign outputs[1126] = layer6_outputs[2891];
    assign outputs[1127] = (layer6_outputs[4466]) ^ (layer6_outputs[1037]);
    assign outputs[1128] = ~(layer6_outputs[3319]);
    assign outputs[1129] = ~(layer6_outputs[3712]);
    assign outputs[1130] = ~((layer6_outputs[4290]) ^ (layer6_outputs[2185]));
    assign outputs[1131] = ~(layer6_outputs[3761]);
    assign outputs[1132] = ~((layer6_outputs[2641]) ^ (layer6_outputs[3044]));
    assign outputs[1133] = layer6_outputs[55];
    assign outputs[1134] = layer6_outputs[4516];
    assign outputs[1135] = ~(layer6_outputs[3033]);
    assign outputs[1136] = layer6_outputs[2226];
    assign outputs[1137] = ~(layer6_outputs[3559]) | (layer6_outputs[1435]);
    assign outputs[1138] = (layer6_outputs[2232]) ^ (layer6_outputs[1929]);
    assign outputs[1139] = layer6_outputs[3707];
    assign outputs[1140] = (layer6_outputs[3717]) & (layer6_outputs[3825]);
    assign outputs[1141] = ~(layer6_outputs[1841]);
    assign outputs[1142] = ~(layer6_outputs[1627]);
    assign outputs[1143] = (layer6_outputs[463]) & (layer6_outputs[4079]);
    assign outputs[1144] = ~(layer6_outputs[4391]) | (layer6_outputs[2659]);
    assign outputs[1145] = (layer6_outputs[2725]) ^ (layer6_outputs[4853]);
    assign outputs[1146] = ~((layer6_outputs[2202]) ^ (layer6_outputs[1862]));
    assign outputs[1147] = layer6_outputs[4750];
    assign outputs[1148] = layer6_outputs[5034];
    assign outputs[1149] = (layer6_outputs[4769]) ^ (layer6_outputs[261]);
    assign outputs[1150] = ~((layer6_outputs[1541]) & (layer6_outputs[4877]));
    assign outputs[1151] = ~((layer6_outputs[1150]) ^ (layer6_outputs[1387]));
    assign outputs[1152] = layer6_outputs[3353];
    assign outputs[1153] = layer6_outputs[3153];
    assign outputs[1154] = layer6_outputs[207];
    assign outputs[1155] = layer6_outputs[2250];
    assign outputs[1156] = ~(layer6_outputs[3317]);
    assign outputs[1157] = layer6_outputs[979];
    assign outputs[1158] = layer6_outputs[2651];
    assign outputs[1159] = ~(layer6_outputs[2901]);
    assign outputs[1160] = layer6_outputs[1260];
    assign outputs[1161] = ~((layer6_outputs[667]) ^ (layer6_outputs[1001]));
    assign outputs[1162] = ~((layer6_outputs[1309]) ^ (layer6_outputs[2334]));
    assign outputs[1163] = layer6_outputs[3044];
    assign outputs[1164] = (layer6_outputs[534]) & (layer6_outputs[1576]);
    assign outputs[1165] = layer6_outputs[3015];
    assign outputs[1166] = (layer6_outputs[1107]) & ~(layer6_outputs[2375]);
    assign outputs[1167] = layer6_outputs[4557];
    assign outputs[1168] = layer6_outputs[2894];
    assign outputs[1169] = layer6_outputs[48];
    assign outputs[1170] = ~(layer6_outputs[4916]);
    assign outputs[1171] = ~(layer6_outputs[1188]);
    assign outputs[1172] = ~(layer6_outputs[3379]);
    assign outputs[1173] = layer6_outputs[123];
    assign outputs[1174] = ~(layer6_outputs[1802]);
    assign outputs[1175] = ~(layer6_outputs[3815]);
    assign outputs[1176] = ~(layer6_outputs[3026]);
    assign outputs[1177] = ~(layer6_outputs[4577]);
    assign outputs[1178] = ~((layer6_outputs[1266]) ^ (layer6_outputs[954]));
    assign outputs[1179] = (layer6_outputs[424]) & ~(layer6_outputs[1669]);
    assign outputs[1180] = layer6_outputs[32];
    assign outputs[1181] = ~(layer6_outputs[2442]);
    assign outputs[1182] = ~(layer6_outputs[3950]);
    assign outputs[1183] = layer6_outputs[5027];
    assign outputs[1184] = layer6_outputs[66];
    assign outputs[1185] = (layer6_outputs[1749]) ^ (layer6_outputs[566]);
    assign outputs[1186] = ~((layer6_outputs[894]) ^ (layer6_outputs[2850]));
    assign outputs[1187] = (layer6_outputs[1938]) ^ (layer6_outputs[3954]);
    assign outputs[1188] = layer6_outputs[4901];
    assign outputs[1189] = ~(layer6_outputs[28]);
    assign outputs[1190] = ~(layer6_outputs[1428]);
    assign outputs[1191] = layer6_outputs[2919];
    assign outputs[1192] = ~((layer6_outputs[2517]) ^ (layer6_outputs[2260]));
    assign outputs[1193] = layer6_outputs[4971];
    assign outputs[1194] = layer6_outputs[4340];
    assign outputs[1195] = ~(layer6_outputs[4363]);
    assign outputs[1196] = ~((layer6_outputs[3214]) ^ (layer6_outputs[2197]));
    assign outputs[1197] = layer6_outputs[271];
    assign outputs[1198] = ~(layer6_outputs[4910]);
    assign outputs[1199] = ~((layer6_outputs[1536]) ^ (layer6_outputs[2825]));
    assign outputs[1200] = ~((layer6_outputs[4891]) ^ (layer6_outputs[4144]));
    assign outputs[1201] = layer6_outputs[1947];
    assign outputs[1202] = (layer6_outputs[2280]) ^ (layer6_outputs[4978]);
    assign outputs[1203] = layer6_outputs[2419];
    assign outputs[1204] = layer6_outputs[2583];
    assign outputs[1205] = ~(layer6_outputs[4183]);
    assign outputs[1206] = ~(layer6_outputs[1420]);
    assign outputs[1207] = ~(layer6_outputs[3898]);
    assign outputs[1208] = ~(layer6_outputs[4488]);
    assign outputs[1209] = ~(layer6_outputs[734]);
    assign outputs[1210] = layer6_outputs[2213];
    assign outputs[1211] = ~((layer6_outputs[2857]) | (layer6_outputs[4188]));
    assign outputs[1212] = layer6_outputs[3849];
    assign outputs[1213] = layer6_outputs[539];
    assign outputs[1214] = ~((layer6_outputs[3959]) ^ (layer6_outputs[3798]));
    assign outputs[1215] = layer6_outputs[1956];
    assign outputs[1216] = layer6_outputs[2220];
    assign outputs[1217] = (layer6_outputs[3441]) ^ (layer6_outputs[4695]);
    assign outputs[1218] = ~((layer6_outputs[335]) ^ (layer6_outputs[4581]));
    assign outputs[1219] = ~((layer6_outputs[1290]) & (layer6_outputs[2204]));
    assign outputs[1220] = ~(layer6_outputs[2269]);
    assign outputs[1221] = (layer6_outputs[4405]) & ~(layer6_outputs[744]);
    assign outputs[1222] = ~(layer6_outputs[3178]);
    assign outputs[1223] = ~(layer6_outputs[2995]);
    assign outputs[1224] = ~((layer6_outputs[4046]) ^ (layer6_outputs[2727]));
    assign outputs[1225] = (layer6_outputs[3510]) & ~(layer6_outputs[4864]);
    assign outputs[1226] = layer6_outputs[4980];
    assign outputs[1227] = ~(layer6_outputs[1300]);
    assign outputs[1228] = ~(layer6_outputs[4191]);
    assign outputs[1229] = ~(layer6_outputs[3025]);
    assign outputs[1230] = ~(layer6_outputs[4977]) | (layer6_outputs[4699]);
    assign outputs[1231] = ~((layer6_outputs[1998]) ^ (layer6_outputs[511]));
    assign outputs[1232] = ~(layer6_outputs[501]);
    assign outputs[1233] = layer6_outputs[3017];
    assign outputs[1234] = ~(layer6_outputs[289]);
    assign outputs[1235] = ~((layer6_outputs[19]) ^ (layer6_outputs[2994]));
    assign outputs[1236] = (layer6_outputs[3872]) ^ (layer6_outputs[197]);
    assign outputs[1237] = layer6_outputs[3159];
    assign outputs[1238] = layer6_outputs[250];
    assign outputs[1239] = (layer6_outputs[984]) ^ (layer6_outputs[627]);
    assign outputs[1240] = (layer6_outputs[4272]) ^ (layer6_outputs[4722]);
    assign outputs[1241] = ~((layer6_outputs[4097]) | (layer6_outputs[3176]));
    assign outputs[1242] = layer6_outputs[1992];
    assign outputs[1243] = ~((layer6_outputs[531]) ^ (layer6_outputs[2869]));
    assign outputs[1244] = layer6_outputs[4051];
    assign outputs[1245] = layer6_outputs[2570];
    assign outputs[1246] = (layer6_outputs[525]) ^ (layer6_outputs[1079]);
    assign outputs[1247] = layer6_outputs[1087];
    assign outputs[1248] = layer6_outputs[4104];
    assign outputs[1249] = layer6_outputs[4327];
    assign outputs[1250] = ~((layer6_outputs[2801]) ^ (layer6_outputs[141]));
    assign outputs[1251] = ~((layer6_outputs[3833]) ^ (layer6_outputs[4751]));
    assign outputs[1252] = ~(layer6_outputs[1442]);
    assign outputs[1253] = ~(layer6_outputs[2870]);
    assign outputs[1254] = layer6_outputs[3396];
    assign outputs[1255] = ~(layer6_outputs[4200]);
    assign outputs[1256] = ~(layer6_outputs[3455]) | (layer6_outputs[4813]);
    assign outputs[1257] = (layer6_outputs[3615]) ^ (layer6_outputs[3795]);
    assign outputs[1258] = ~(layer6_outputs[4168]);
    assign outputs[1259] = layer6_outputs[1868];
    assign outputs[1260] = (layer6_outputs[1788]) ^ (layer6_outputs[3931]);
    assign outputs[1261] = ~(layer6_outputs[4556]);
    assign outputs[1262] = (layer6_outputs[3744]) ^ (layer6_outputs[4059]);
    assign outputs[1263] = ~((layer6_outputs[3556]) ^ (layer6_outputs[2883]));
    assign outputs[1264] = ~((layer6_outputs[635]) ^ (layer6_outputs[4443]));
    assign outputs[1265] = (layer6_outputs[2950]) ^ (layer6_outputs[2156]);
    assign outputs[1266] = layer6_outputs[709];
    assign outputs[1267] = (layer6_outputs[4622]) ^ (layer6_outputs[1286]);
    assign outputs[1268] = ~((layer6_outputs[5092]) ^ (layer6_outputs[861]));
    assign outputs[1269] = layer6_outputs[662];
    assign outputs[1270] = ~(layer6_outputs[87]);
    assign outputs[1271] = ~(layer6_outputs[2701]);
    assign outputs[1272] = ~(layer6_outputs[3587]);
    assign outputs[1273] = (layer6_outputs[266]) ^ (layer6_outputs[3735]);
    assign outputs[1274] = layer6_outputs[3058];
    assign outputs[1275] = ~(layer6_outputs[1943]);
    assign outputs[1276] = ~(layer6_outputs[1963]);
    assign outputs[1277] = ~(layer6_outputs[3221]);
    assign outputs[1278] = layer6_outputs[4485];
    assign outputs[1279] = layer6_outputs[140];
    assign outputs[1280] = ~((layer6_outputs[1892]) | (layer6_outputs[2435]));
    assign outputs[1281] = (layer6_outputs[1807]) ^ (layer6_outputs[874]);
    assign outputs[1282] = layer6_outputs[1197];
    assign outputs[1283] = ~(layer6_outputs[1146]);
    assign outputs[1284] = ~(layer6_outputs[2026]);
    assign outputs[1285] = layer6_outputs[3735];
    assign outputs[1286] = layer6_outputs[4095];
    assign outputs[1287] = ~(layer6_outputs[938]);
    assign outputs[1288] = ~((layer6_outputs[4471]) ^ (layer6_outputs[5075]));
    assign outputs[1289] = (layer6_outputs[4280]) ^ (layer6_outputs[3136]);
    assign outputs[1290] = ~(layer6_outputs[1364]);
    assign outputs[1291] = ~(layer6_outputs[3610]);
    assign outputs[1292] = ~(layer6_outputs[2017]);
    assign outputs[1293] = ~(layer6_outputs[3246]);
    assign outputs[1294] = ~(layer6_outputs[1514]);
    assign outputs[1295] = layer6_outputs[60];
    assign outputs[1296] = layer6_outputs[257];
    assign outputs[1297] = layer6_outputs[4616];
    assign outputs[1298] = (layer6_outputs[1021]) | (layer6_outputs[2482]);
    assign outputs[1299] = ~((layer6_outputs[874]) ^ (layer6_outputs[2414]));
    assign outputs[1300] = ~(layer6_outputs[532]);
    assign outputs[1301] = ~((layer6_outputs[2277]) ^ (layer6_outputs[197]));
    assign outputs[1302] = ~((layer6_outputs[2892]) ^ (layer6_outputs[3597]));
    assign outputs[1303] = layer6_outputs[2230];
    assign outputs[1304] = layer6_outputs[4855];
    assign outputs[1305] = (layer6_outputs[3421]) ^ (layer6_outputs[790]);
    assign outputs[1306] = ~((layer6_outputs[3905]) ^ (layer6_outputs[1847]));
    assign outputs[1307] = layer6_outputs[4903];
    assign outputs[1308] = ~(layer6_outputs[2039]) | (layer6_outputs[449]);
    assign outputs[1309] = ~(layer6_outputs[1715]);
    assign outputs[1310] = ~((layer6_outputs[346]) & (layer6_outputs[594]));
    assign outputs[1311] = layer6_outputs[2556];
    assign outputs[1312] = ~(layer6_outputs[3301]);
    assign outputs[1313] = layer6_outputs[3991];
    assign outputs[1314] = layer6_outputs[667];
    assign outputs[1315] = ~(layer6_outputs[399]);
    assign outputs[1316] = ~(layer6_outputs[1741]) | (layer6_outputs[4343]);
    assign outputs[1317] = ~(layer6_outputs[2498]);
    assign outputs[1318] = ~(layer6_outputs[5113]);
    assign outputs[1319] = ~((layer6_outputs[3753]) ^ (layer6_outputs[2843]));
    assign outputs[1320] = layer6_outputs[3731];
    assign outputs[1321] = layer6_outputs[3977];
    assign outputs[1322] = layer6_outputs[3431];
    assign outputs[1323] = ~(layer6_outputs[4332]);
    assign outputs[1324] = ~(layer6_outputs[122]);
    assign outputs[1325] = (layer6_outputs[3437]) ^ (layer6_outputs[4062]);
    assign outputs[1326] = layer6_outputs[1921];
    assign outputs[1327] = ~(layer6_outputs[4313]);
    assign outputs[1328] = layer6_outputs[2448];
    assign outputs[1329] = ~(layer6_outputs[4933]);
    assign outputs[1330] = ~(layer6_outputs[4957]);
    assign outputs[1331] = ~(layer6_outputs[3867]);
    assign outputs[1332] = ~(layer6_outputs[2693]) | (layer6_outputs[3660]);
    assign outputs[1333] = ~(layer6_outputs[4487]) | (layer6_outputs[669]);
    assign outputs[1334] = ~(layer6_outputs[218]) | (layer6_outputs[2751]);
    assign outputs[1335] = (layer6_outputs[482]) & ~(layer6_outputs[57]);
    assign outputs[1336] = ~(layer6_outputs[2455]);
    assign outputs[1337] = (layer6_outputs[400]) ^ (layer6_outputs[1476]);
    assign outputs[1338] = ~((layer6_outputs[3129]) ^ (layer6_outputs[2748]));
    assign outputs[1339] = layer6_outputs[2446];
    assign outputs[1340] = layer6_outputs[2643];
    assign outputs[1341] = ~(layer6_outputs[78]);
    assign outputs[1342] = layer6_outputs[797];
    assign outputs[1343] = ~(layer6_outputs[2270]);
    assign outputs[1344] = layer6_outputs[2301];
    assign outputs[1345] = ~(layer6_outputs[4573]);
    assign outputs[1346] = layer6_outputs[1108];
    assign outputs[1347] = layer6_outputs[4162];
    assign outputs[1348] = (layer6_outputs[2589]) & ~(layer6_outputs[387]);
    assign outputs[1349] = layer6_outputs[1289];
    assign outputs[1350] = layer6_outputs[4904];
    assign outputs[1351] = ~(layer6_outputs[807]);
    assign outputs[1352] = ~(layer6_outputs[3804]) | (layer6_outputs[4393]);
    assign outputs[1353] = (layer6_outputs[617]) | (layer6_outputs[4816]);
    assign outputs[1354] = layer6_outputs[29];
    assign outputs[1355] = (layer6_outputs[951]) & ~(layer6_outputs[2757]);
    assign outputs[1356] = ~((layer6_outputs[525]) ^ (layer6_outputs[269]));
    assign outputs[1357] = layer6_outputs[623];
    assign outputs[1358] = layer6_outputs[1604];
    assign outputs[1359] = ~(layer6_outputs[3133]);
    assign outputs[1360] = layer6_outputs[4029];
    assign outputs[1361] = layer6_outputs[3929];
    assign outputs[1362] = layer6_outputs[163];
    assign outputs[1363] = ~((layer6_outputs[3211]) ^ (layer6_outputs[1088]));
    assign outputs[1364] = layer6_outputs[1538];
    assign outputs[1365] = layer6_outputs[3304];
    assign outputs[1366] = ~(layer6_outputs[2555]);
    assign outputs[1367] = (layer6_outputs[649]) ^ (layer6_outputs[3251]);
    assign outputs[1368] = ~(layer6_outputs[4828]);
    assign outputs[1369] = layer6_outputs[726];
    assign outputs[1370] = layer6_outputs[4930];
    assign outputs[1371] = layer6_outputs[3589];
    assign outputs[1372] = ~(layer6_outputs[3999]);
    assign outputs[1373] = layer6_outputs[4425];
    assign outputs[1374] = (layer6_outputs[2657]) ^ (layer6_outputs[2731]);
    assign outputs[1375] = ~(layer6_outputs[652]);
    assign outputs[1376] = ~(layer6_outputs[214]);
    assign outputs[1377] = (layer6_outputs[4189]) ^ (layer6_outputs[4080]);
    assign outputs[1378] = ~((layer6_outputs[1251]) ^ (layer6_outputs[2534]));
    assign outputs[1379] = (layer6_outputs[3819]) ^ (layer6_outputs[2865]);
    assign outputs[1380] = layer6_outputs[4263];
    assign outputs[1381] = ~(layer6_outputs[2957]);
    assign outputs[1382] = ~(layer6_outputs[4548]);
    assign outputs[1383] = layer6_outputs[5053];
    assign outputs[1384] = ~((layer6_outputs[2811]) & (layer6_outputs[1500]));
    assign outputs[1385] = (layer6_outputs[18]) & (layer6_outputs[3757]);
    assign outputs[1386] = ~(layer6_outputs[4828]);
    assign outputs[1387] = ~((layer6_outputs[999]) ^ (layer6_outputs[1458]));
    assign outputs[1388] = layer6_outputs[4650];
    assign outputs[1389] = ~((layer6_outputs[2985]) & (layer6_outputs[3557]));
    assign outputs[1390] = (layer6_outputs[3808]) ^ (layer6_outputs[3422]);
    assign outputs[1391] = ~(layer6_outputs[3031]);
    assign outputs[1392] = layer6_outputs[412];
    assign outputs[1393] = layer6_outputs[2081];
    assign outputs[1394] = ~(layer6_outputs[533]);
    assign outputs[1395] = ~(layer6_outputs[3976]);
    assign outputs[1396] = layer6_outputs[4598];
    assign outputs[1397] = ~((layer6_outputs[2100]) ^ (layer6_outputs[2962]));
    assign outputs[1398] = layer6_outputs[4806];
    assign outputs[1399] = ~(layer6_outputs[71]);
    assign outputs[1400] = ~(layer6_outputs[3516]);
    assign outputs[1401] = ~(layer6_outputs[1010]);
    assign outputs[1402] = layer6_outputs[3775];
    assign outputs[1403] = ~(layer6_outputs[2588]);
    assign outputs[1404] = ~((layer6_outputs[3794]) & (layer6_outputs[3292]));
    assign outputs[1405] = (layer6_outputs[4217]) ^ (layer6_outputs[2784]);
    assign outputs[1406] = layer6_outputs[4999];
    assign outputs[1407] = (layer6_outputs[3637]) & ~(layer6_outputs[1572]);
    assign outputs[1408] = (layer6_outputs[3474]) ^ (layer6_outputs[1232]);
    assign outputs[1409] = layer6_outputs[4035];
    assign outputs[1410] = layer6_outputs[4331];
    assign outputs[1411] = layer6_outputs[4277];
    assign outputs[1412] = layer6_outputs[333];
    assign outputs[1413] = layer6_outputs[4060];
    assign outputs[1414] = ~(layer6_outputs[597]);
    assign outputs[1415] = ~((layer6_outputs[264]) & (layer6_outputs[409]));
    assign outputs[1416] = ~(layer6_outputs[3634]);
    assign outputs[1417] = layer6_outputs[1377];
    assign outputs[1418] = layer6_outputs[1216];
    assign outputs[1419] = ~((layer6_outputs[1200]) | (layer6_outputs[2684]));
    assign outputs[1420] = ~(layer6_outputs[1866]);
    assign outputs[1421] = layer6_outputs[4268];
    assign outputs[1422] = ~(layer6_outputs[3410]);
    assign outputs[1423] = layer6_outputs[3391];
    assign outputs[1424] = (layer6_outputs[4531]) ^ (layer6_outputs[2180]);
    assign outputs[1425] = layer6_outputs[3771];
    assign outputs[1426] = ~(layer6_outputs[1864]);
    assign outputs[1427] = (layer6_outputs[3182]) & ~(layer6_outputs[5016]);
    assign outputs[1428] = ~(layer6_outputs[31]);
    assign outputs[1429] = ~((layer6_outputs[3970]) ^ (layer6_outputs[1031]));
    assign outputs[1430] = ~(layer6_outputs[4352]);
    assign outputs[1431] = ~((layer6_outputs[4543]) ^ (layer6_outputs[974]));
    assign outputs[1432] = ~((layer6_outputs[625]) & (layer6_outputs[4596]));
    assign outputs[1433] = (layer6_outputs[3195]) ^ (layer6_outputs[1599]);
    assign outputs[1434] = ~((layer6_outputs[91]) ^ (layer6_outputs[3839]));
    assign outputs[1435] = ~(layer6_outputs[2191]);
    assign outputs[1436] = ~(layer6_outputs[3458]) | (layer6_outputs[742]);
    assign outputs[1437] = layer6_outputs[3275];
    assign outputs[1438] = ~(layer6_outputs[501]);
    assign outputs[1439] = ~(layer6_outputs[2665]);
    assign outputs[1440] = ~((layer6_outputs[3860]) ^ (layer6_outputs[4957]));
    assign outputs[1441] = layer6_outputs[875];
    assign outputs[1442] = ~((layer6_outputs[319]) ^ (layer6_outputs[5074]));
    assign outputs[1443] = layer6_outputs[1677];
    assign outputs[1444] = layer6_outputs[2975];
    assign outputs[1445] = ~(layer6_outputs[1060]);
    assign outputs[1446] = (layer6_outputs[1552]) & ~(layer6_outputs[2234]);
    assign outputs[1447] = ~((layer6_outputs[833]) & (layer6_outputs[3899]));
    assign outputs[1448] = ~(layer6_outputs[4329]);
    assign outputs[1449] = ~((layer6_outputs[483]) ^ (layer6_outputs[4813]));
    assign outputs[1450] = layer6_outputs[4609];
    assign outputs[1451] = layer6_outputs[3569];
    assign outputs[1452] = layer6_outputs[904];
    assign outputs[1453] = ~(layer6_outputs[994]) | (layer6_outputs[429]);
    assign outputs[1454] = ~(layer6_outputs[1662]);
    assign outputs[1455] = layer6_outputs[3866];
    assign outputs[1456] = ~((layer6_outputs[2571]) | (layer6_outputs[2503]));
    assign outputs[1457] = layer6_outputs[4132];
    assign outputs[1458] = layer6_outputs[4585];
    assign outputs[1459] = ~(layer6_outputs[3303]) | (layer6_outputs[979]);
    assign outputs[1460] = layer6_outputs[3525];
    assign outputs[1461] = ~((layer6_outputs[1255]) ^ (layer6_outputs[14]));
    assign outputs[1462] = layer6_outputs[2295];
    assign outputs[1463] = layer6_outputs[222];
    assign outputs[1464] = ~((layer6_outputs[1980]) & (layer6_outputs[1091]));
    assign outputs[1465] = ~(layer6_outputs[4374]) | (layer6_outputs[1681]);
    assign outputs[1466] = ~((layer6_outputs[3115]) ^ (layer6_outputs[4940]));
    assign outputs[1467] = ~(layer6_outputs[991]);
    assign outputs[1468] = (layer6_outputs[2575]) & ~(layer6_outputs[2393]);
    assign outputs[1469] = ~(layer6_outputs[1918]) | (layer6_outputs[2372]);
    assign outputs[1470] = layer6_outputs[467];
    assign outputs[1471] = ~(layer6_outputs[2520]);
    assign outputs[1472] = ~(layer6_outputs[3835]);
    assign outputs[1473] = layer6_outputs[1073];
    assign outputs[1474] = ~((layer6_outputs[1973]) | (layer6_outputs[1440]));
    assign outputs[1475] = layer6_outputs[3902];
    assign outputs[1476] = ~(layer6_outputs[3600]);
    assign outputs[1477] = (layer6_outputs[2152]) ^ (layer6_outputs[3400]);
    assign outputs[1478] = layer6_outputs[383];
    assign outputs[1479] = ~(layer6_outputs[1763]);
    assign outputs[1480] = ~(layer6_outputs[2395]);
    assign outputs[1481] = ~(layer6_outputs[4264]);
    assign outputs[1482] = layer6_outputs[4846];
    assign outputs[1483] = layer6_outputs[1739];
    assign outputs[1484] = layer6_outputs[1197];
    assign outputs[1485] = ~((layer6_outputs[4985]) ^ (layer6_outputs[3758]));
    assign outputs[1486] = (layer6_outputs[39]) | (layer6_outputs[3]);
    assign outputs[1487] = layer6_outputs[3849];
    assign outputs[1488] = layer6_outputs[4274];
    assign outputs[1489] = layer6_outputs[2980];
    assign outputs[1490] = ~(layer6_outputs[168]);
    assign outputs[1491] = layer6_outputs[646];
    assign outputs[1492] = ~(layer6_outputs[3710]);
    assign outputs[1493] = ~(layer6_outputs[90]);
    assign outputs[1494] = ~(layer6_outputs[2917]);
    assign outputs[1495] = ~(layer6_outputs[2965]);
    assign outputs[1496] = (layer6_outputs[3232]) ^ (layer6_outputs[2425]);
    assign outputs[1497] = ~((layer6_outputs[1740]) ^ (layer6_outputs[4000]));
    assign outputs[1498] = (layer6_outputs[1612]) ^ (layer6_outputs[930]);
    assign outputs[1499] = layer6_outputs[4258];
    assign outputs[1500] = (layer6_outputs[5086]) | (layer6_outputs[5050]);
    assign outputs[1501] = ~((layer6_outputs[3073]) ^ (layer6_outputs[1031]));
    assign outputs[1502] = (layer6_outputs[793]) ^ (layer6_outputs[1523]);
    assign outputs[1503] = ~((layer6_outputs[2252]) ^ (layer6_outputs[1785]));
    assign outputs[1504] = (layer6_outputs[2795]) ^ (layer6_outputs[2794]);
    assign outputs[1505] = ~(layer6_outputs[2875]);
    assign outputs[1506] = layer6_outputs[3002];
    assign outputs[1507] = ~((layer6_outputs[131]) ^ (layer6_outputs[1159]));
    assign outputs[1508] = ~(layer6_outputs[2063]);
    assign outputs[1509] = ~((layer6_outputs[2997]) & (layer6_outputs[4129]));
    assign outputs[1510] = ~((layer6_outputs[4701]) ^ (layer6_outputs[1803]));
    assign outputs[1511] = layer6_outputs[1824];
    assign outputs[1512] = (layer6_outputs[4750]) ^ (layer6_outputs[4249]);
    assign outputs[1513] = (layer6_outputs[3698]) & ~(layer6_outputs[3536]);
    assign outputs[1514] = ~((layer6_outputs[1298]) | (layer6_outputs[504]));
    assign outputs[1515] = ~(layer6_outputs[1826]);
    assign outputs[1516] = ~(layer6_outputs[2993]) | (layer6_outputs[1294]);
    assign outputs[1517] = ~(layer6_outputs[4378]);
    assign outputs[1518] = (layer6_outputs[1190]) & ~(layer6_outputs[2498]);
    assign outputs[1519] = ~((layer6_outputs[4831]) ^ (layer6_outputs[468]));
    assign outputs[1520] = layer6_outputs[3626];
    assign outputs[1521] = ~(layer6_outputs[3913]);
    assign outputs[1522] = (layer6_outputs[3490]) ^ (layer6_outputs[925]);
    assign outputs[1523] = ~(layer6_outputs[1682]);
    assign outputs[1524] = ~((layer6_outputs[152]) ^ (layer6_outputs[4325]));
    assign outputs[1525] = (layer6_outputs[2471]) ^ (layer6_outputs[2610]);
    assign outputs[1526] = ~((layer6_outputs[4382]) ^ (layer6_outputs[3795]));
    assign outputs[1527] = layer6_outputs[1583];
    assign outputs[1528] = ~(layer6_outputs[913]) | (layer6_outputs[3497]);
    assign outputs[1529] = layer6_outputs[2308];
    assign outputs[1530] = ~((layer6_outputs[600]) | (layer6_outputs[629]));
    assign outputs[1531] = ~(layer6_outputs[3452]);
    assign outputs[1532] = layer6_outputs[3996];
    assign outputs[1533] = layer6_outputs[3126];
    assign outputs[1534] = ~(layer6_outputs[3538]);
    assign outputs[1535] = layer6_outputs[963];
    assign outputs[1536] = layer6_outputs[3467];
    assign outputs[1537] = ~((layer6_outputs[3503]) | (layer6_outputs[1542]));
    assign outputs[1538] = layer6_outputs[86];
    assign outputs[1539] = (layer6_outputs[829]) ^ (layer6_outputs[4424]);
    assign outputs[1540] = ~(layer6_outputs[2906]);
    assign outputs[1541] = layer6_outputs[325];
    assign outputs[1542] = ~((layer6_outputs[3759]) | (layer6_outputs[1135]));
    assign outputs[1543] = ~(layer6_outputs[4992]);
    assign outputs[1544] = (layer6_outputs[857]) & ~(layer6_outputs[3450]);
    assign outputs[1545] = ~(layer6_outputs[4460]);
    assign outputs[1546] = ~(layer6_outputs[769]) | (layer6_outputs[1963]);
    assign outputs[1547] = (layer6_outputs[688]) ^ (layer6_outputs[2319]);
    assign outputs[1548] = (layer6_outputs[2470]) & ~(layer6_outputs[959]);
    assign outputs[1549] = (layer6_outputs[1896]) & (layer6_outputs[5050]);
    assign outputs[1550] = (layer6_outputs[3486]) ^ (layer6_outputs[5048]);
    assign outputs[1551] = ~(layer6_outputs[2698]);
    assign outputs[1552] = (layer6_outputs[246]) ^ (layer6_outputs[1312]);
    assign outputs[1553] = layer6_outputs[4082];
    assign outputs[1554] = ~(layer6_outputs[5087]);
    assign outputs[1555] = (layer6_outputs[4504]) & ~(layer6_outputs[3542]);
    assign outputs[1556] = ~(layer6_outputs[1123]);
    assign outputs[1557] = ~(layer6_outputs[3568]);
    assign outputs[1558] = (layer6_outputs[2567]) ^ (layer6_outputs[1578]);
    assign outputs[1559] = (layer6_outputs[2865]) ^ (layer6_outputs[237]);
    assign outputs[1560] = layer6_outputs[4917];
    assign outputs[1561] = layer6_outputs[2553];
    assign outputs[1562] = ~((layer6_outputs[1902]) | (layer6_outputs[1626]));
    assign outputs[1563] = ~((layer6_outputs[4148]) ^ (layer6_outputs[3364]));
    assign outputs[1564] = ~(layer6_outputs[2462]);
    assign outputs[1565] = ~((layer6_outputs[2215]) & (layer6_outputs[3890]));
    assign outputs[1566] = (layer6_outputs[1874]) & (layer6_outputs[1136]);
    assign outputs[1567] = ~(layer6_outputs[2013]);
    assign outputs[1568] = layer6_outputs[324];
    assign outputs[1569] = layer6_outputs[4524];
    assign outputs[1570] = ~(layer6_outputs[1684]);
    assign outputs[1571] = (layer6_outputs[4683]) ^ (layer6_outputs[4338]);
    assign outputs[1572] = (layer6_outputs[3838]) ^ (layer6_outputs[1923]);
    assign outputs[1573] = (layer6_outputs[2897]) | (layer6_outputs[1495]);
    assign outputs[1574] = layer6_outputs[3288];
    assign outputs[1575] = ~((layer6_outputs[4418]) | (layer6_outputs[3811]));
    assign outputs[1576] = (layer6_outputs[766]) & ~(layer6_outputs[983]);
    assign outputs[1577] = ~(layer6_outputs[5034]);
    assign outputs[1578] = layer6_outputs[2404];
    assign outputs[1579] = layer6_outputs[4348];
    assign outputs[1580] = layer6_outputs[1926];
    assign outputs[1581] = ~(layer6_outputs[4189]);
    assign outputs[1582] = layer6_outputs[3146];
    assign outputs[1583] = ~((layer6_outputs[3210]) ^ (layer6_outputs[3091]));
    assign outputs[1584] = ~(layer6_outputs[271]);
    assign outputs[1585] = (layer6_outputs[2333]) & (layer6_outputs[196]);
    assign outputs[1586] = ~(layer6_outputs[245]);
    assign outputs[1587] = layer6_outputs[3077];
    assign outputs[1588] = (layer6_outputs[4726]) ^ (layer6_outputs[111]);
    assign outputs[1589] = ~(layer6_outputs[2525]);
    assign outputs[1590] = layer6_outputs[3059];
    assign outputs[1591] = ~(layer6_outputs[712]);
    assign outputs[1592] = (layer6_outputs[2189]) ^ (layer6_outputs[3340]);
    assign outputs[1593] = (layer6_outputs[2899]) ^ (layer6_outputs[92]);
    assign outputs[1594] = layer6_outputs[1310];
    assign outputs[1595] = layer6_outputs[2273];
    assign outputs[1596] = ~(layer6_outputs[460]);
    assign outputs[1597] = layer6_outputs[3118];
    assign outputs[1598] = layer6_outputs[2196];
    assign outputs[1599] = layer6_outputs[1047];
    assign outputs[1600] = layer6_outputs[548];
    assign outputs[1601] = ~(layer6_outputs[4251]);
    assign outputs[1602] = ~((layer6_outputs[2390]) ^ (layer6_outputs[2724]));
    assign outputs[1603] = layer6_outputs[27];
    assign outputs[1604] = layer6_outputs[4443];
    assign outputs[1605] = layer6_outputs[933];
    assign outputs[1606] = layer6_outputs[543];
    assign outputs[1607] = ~((layer6_outputs[12]) ^ (layer6_outputs[1995]));
    assign outputs[1608] = layer6_outputs[2616];
    assign outputs[1609] = layer6_outputs[1906];
    assign outputs[1610] = ~(layer6_outputs[1839]) | (layer6_outputs[3080]);
    assign outputs[1611] = ~((layer6_outputs[4601]) ^ (layer6_outputs[1032]));
    assign outputs[1612] = ~((layer6_outputs[1502]) ^ (layer6_outputs[2463]));
    assign outputs[1613] = layer6_outputs[3748];
    assign outputs[1614] = layer6_outputs[1097];
    assign outputs[1615] = (layer6_outputs[1411]) & ~(layer6_outputs[3854]);
    assign outputs[1616] = (layer6_outputs[2049]) ^ (layer6_outputs[917]);
    assign outputs[1617] = (layer6_outputs[2833]) & ~(layer6_outputs[881]);
    assign outputs[1618] = layer6_outputs[3638];
    assign outputs[1619] = (layer6_outputs[1460]) ^ (layer6_outputs[924]);
    assign outputs[1620] = ~((layer6_outputs[2940]) ^ (layer6_outputs[739]));
    assign outputs[1621] = layer6_outputs[4359];
    assign outputs[1622] = (layer6_outputs[1567]) & ~(layer6_outputs[1404]);
    assign outputs[1623] = ~(layer6_outputs[3615]);
    assign outputs[1624] = ~(layer6_outputs[2948]);
    assign outputs[1625] = layer6_outputs[2308];
    assign outputs[1626] = ~((layer6_outputs[3298]) | (layer6_outputs[346]));
    assign outputs[1627] = ~(layer6_outputs[4429]);
    assign outputs[1628] = ~(layer6_outputs[4191]);
    assign outputs[1629] = ~((layer6_outputs[2032]) ^ (layer6_outputs[4269]));
    assign outputs[1630] = ~(layer6_outputs[486]);
    assign outputs[1631] = (layer6_outputs[2568]) & (layer6_outputs[1407]);
    assign outputs[1632] = layer6_outputs[1503];
    assign outputs[1633] = layer6_outputs[5080];
    assign outputs[1634] = (layer6_outputs[1857]) & ~(layer6_outputs[3150]);
    assign outputs[1635] = (layer6_outputs[2837]) ^ (layer6_outputs[8]);
    assign outputs[1636] = ~(layer6_outputs[973]);
    assign outputs[1637] = (layer6_outputs[3933]) & ~(layer6_outputs[3979]);
    assign outputs[1638] = layer6_outputs[396];
    assign outputs[1639] = layer6_outputs[5081];
    assign outputs[1640] = ~(layer6_outputs[2699]);
    assign outputs[1641] = layer6_outputs[4062];
    assign outputs[1642] = ~(layer6_outputs[4742]);
    assign outputs[1643] = layer6_outputs[1050];
    assign outputs[1644] = ~((layer6_outputs[803]) ^ (layer6_outputs[1434]));
    assign outputs[1645] = ~((layer6_outputs[741]) ^ (layer6_outputs[2518]));
    assign outputs[1646] = layer6_outputs[965];
    assign outputs[1647] = layer6_outputs[2199];
    assign outputs[1648] = layer6_outputs[3040];
    assign outputs[1649] = ~(layer6_outputs[3418]);
    assign outputs[1650] = layer6_outputs[4568];
    assign outputs[1651] = ~((layer6_outputs[3631]) ^ (layer6_outputs[2788]));
    assign outputs[1652] = ~(layer6_outputs[205]);
    assign outputs[1653] = ~(layer6_outputs[4153]);
    assign outputs[1654] = ~(layer6_outputs[869]);
    assign outputs[1655] = ~(layer6_outputs[973]);
    assign outputs[1656] = ~(layer6_outputs[4431]);
    assign outputs[1657] = ~(layer6_outputs[4202]);
    assign outputs[1658] = ~(layer6_outputs[1860]) | (layer6_outputs[1467]);
    assign outputs[1659] = ~((layer6_outputs[3876]) ^ (layer6_outputs[2360]));
    assign outputs[1660] = (layer6_outputs[2932]) ^ (layer6_outputs[1437]);
    assign outputs[1661] = ~((layer6_outputs[1213]) ^ (layer6_outputs[4675]));
    assign outputs[1662] = (layer6_outputs[1040]) & ~(layer6_outputs[4108]);
    assign outputs[1663] = ~(layer6_outputs[3046]);
    assign outputs[1664] = ~(layer6_outputs[3828]);
    assign outputs[1665] = ~(layer6_outputs[2061]) | (layer6_outputs[3619]);
    assign outputs[1666] = (layer6_outputs[3286]) & ~(layer6_outputs[4845]);
    assign outputs[1667] = layer6_outputs[3365];
    assign outputs[1668] = (layer6_outputs[513]) ^ (layer6_outputs[3045]);
    assign outputs[1669] = ~(layer6_outputs[232]);
    assign outputs[1670] = layer6_outputs[1763];
    assign outputs[1671] = layer6_outputs[5072];
    assign outputs[1672] = layer6_outputs[2771];
    assign outputs[1673] = ~((layer6_outputs[1575]) ^ (layer6_outputs[386]));
    assign outputs[1674] = ~(layer6_outputs[2391]) | (layer6_outputs[2023]);
    assign outputs[1675] = ~(layer6_outputs[787]);
    assign outputs[1676] = layer6_outputs[3421];
    assign outputs[1677] = ~(layer6_outputs[978]);
    assign outputs[1678] = (layer6_outputs[549]) & ~(layer6_outputs[4734]);
    assign outputs[1679] = ~((layer6_outputs[1707]) ^ (layer6_outputs[4845]));
    assign outputs[1680] = ~((layer6_outputs[4139]) ^ (layer6_outputs[4475]));
    assign outputs[1681] = ~((layer6_outputs[2143]) & (layer6_outputs[2384]));
    assign outputs[1682] = (layer6_outputs[730]) ^ (layer6_outputs[624]);
    assign outputs[1683] = layer6_outputs[68];
    assign outputs[1684] = ~((layer6_outputs[2281]) & (layer6_outputs[4261]));
    assign outputs[1685] = layer6_outputs[4077];
    assign outputs[1686] = ~(layer6_outputs[4754]);
    assign outputs[1687] = layer6_outputs[3397];
    assign outputs[1688] = ~(layer6_outputs[3711]);
    assign outputs[1689] = ~(layer6_outputs[2275]);
    assign outputs[1690] = layer6_outputs[1874];
    assign outputs[1691] = ~(layer6_outputs[4430]);
    assign outputs[1692] = (layer6_outputs[3750]) ^ (layer6_outputs[2660]);
    assign outputs[1693] = (layer6_outputs[3790]) ^ (layer6_outputs[1211]);
    assign outputs[1694] = ~((layer6_outputs[3444]) ^ (layer6_outputs[1007]));
    assign outputs[1695] = (layer6_outputs[2973]) ^ (layer6_outputs[4815]);
    assign outputs[1696] = ~(layer6_outputs[2279]);
    assign outputs[1697] = ~((layer6_outputs[1897]) | (layer6_outputs[2514]));
    assign outputs[1698] = ~((layer6_outputs[4321]) & (layer6_outputs[75]));
    assign outputs[1699] = (layer6_outputs[1564]) & ~(layer6_outputs[132]);
    assign outputs[1700] = (layer6_outputs[2413]) & (layer6_outputs[243]);
    assign outputs[1701] = ~(layer6_outputs[4762]);
    assign outputs[1702] = ~(layer6_outputs[3217]);
    assign outputs[1703] = ~(layer6_outputs[3319]);
    assign outputs[1704] = ~(layer6_outputs[5098]);
    assign outputs[1705] = (layer6_outputs[1605]) ^ (layer6_outputs[4116]);
    assign outputs[1706] = ~((layer6_outputs[1573]) ^ (layer6_outputs[3114]));
    assign outputs[1707] = ~((layer6_outputs[3152]) ^ (layer6_outputs[3583]));
    assign outputs[1708] = ~(layer6_outputs[3285]);
    assign outputs[1709] = ~((layer6_outputs[2779]) ^ (layer6_outputs[4922]));
    assign outputs[1710] = ~(layer6_outputs[2859]);
    assign outputs[1711] = ~(layer6_outputs[4842]);
    assign outputs[1712] = layer6_outputs[3685];
    assign outputs[1713] = (layer6_outputs[4669]) ^ (layer6_outputs[1396]);
    assign outputs[1714] = (layer6_outputs[1401]) ^ (layer6_outputs[2339]);
    assign outputs[1715] = ~(layer6_outputs[1617]);
    assign outputs[1716] = ~((layer6_outputs[966]) | (layer6_outputs[3609]));
    assign outputs[1717] = layer6_outputs[31];
    assign outputs[1718] = ~(layer6_outputs[2119]) | (layer6_outputs[817]);
    assign outputs[1719] = ~((layer6_outputs[932]) ^ (layer6_outputs[5013]));
    assign outputs[1720] = layer6_outputs[995];
    assign outputs[1721] = ~(layer6_outputs[3496]);
    assign outputs[1722] = (layer6_outputs[4449]) | (layer6_outputs[3154]);
    assign outputs[1723] = layer6_outputs[3203];
    assign outputs[1724] = layer6_outputs[2082];
    assign outputs[1725] = layer6_outputs[2451];
    assign outputs[1726] = (layer6_outputs[1815]) ^ (layer6_outputs[440]);
    assign outputs[1727] = layer6_outputs[4822];
    assign outputs[1728] = layer6_outputs[4413];
    assign outputs[1729] = ~(layer6_outputs[4799]);
    assign outputs[1730] = (layer6_outputs[505]) & ~(layer6_outputs[3041]);
    assign outputs[1731] = ~(layer6_outputs[3274]);
    assign outputs[1732] = ~((layer6_outputs[237]) ^ (layer6_outputs[3387]));
    assign outputs[1733] = layer6_outputs[381];
    assign outputs[1734] = ~(layer6_outputs[104]);
    assign outputs[1735] = layer6_outputs[2986];
    assign outputs[1736] = layer6_outputs[5110];
    assign outputs[1737] = ~(layer6_outputs[2342]);
    assign outputs[1738] = layer6_outputs[4766];
    assign outputs[1739] = ~(layer6_outputs[1355]);
    assign outputs[1740] = ~(layer6_outputs[187]);
    assign outputs[1741] = ~((layer6_outputs[2037]) ^ (layer6_outputs[1509]));
    assign outputs[1742] = (layer6_outputs[4242]) ^ (layer6_outputs[1758]);
    assign outputs[1743] = ~(layer6_outputs[2698]);
    assign outputs[1744] = layer6_outputs[1392];
    assign outputs[1745] = (layer6_outputs[1647]) & ~(layer6_outputs[2838]);
    assign outputs[1746] = ~(layer6_outputs[4497]);
    assign outputs[1747] = ~(layer6_outputs[1856]);
    assign outputs[1748] = ~(layer6_outputs[2352]);
    assign outputs[1749] = layer6_outputs[4334];
    assign outputs[1750] = (layer6_outputs[4772]) ^ (layer6_outputs[1323]);
    assign outputs[1751] = layer6_outputs[2155];
    assign outputs[1752] = layer6_outputs[4316];
    assign outputs[1753] = ~((layer6_outputs[2141]) ^ (layer6_outputs[1676]));
    assign outputs[1754] = ~(layer6_outputs[5053]);
    assign outputs[1755] = ~(layer6_outputs[1581]);
    assign outputs[1756] = ~(layer6_outputs[4081]);
    assign outputs[1757] = ~((layer6_outputs[4003]) ^ (layer6_outputs[4520]));
    assign outputs[1758] = layer6_outputs[3928];
    assign outputs[1759] = ~(layer6_outputs[423]);
    assign outputs[1760] = layer6_outputs[2834];
    assign outputs[1761] = ~((layer6_outputs[4480]) ^ (layer6_outputs[2786]));
    assign outputs[1762] = layer6_outputs[1737];
    assign outputs[1763] = layer6_outputs[1335];
    assign outputs[1764] = ~((layer6_outputs[2482]) | (layer6_outputs[507]));
    assign outputs[1765] = ~(layer6_outputs[800]);
    assign outputs[1766] = ~(layer6_outputs[2143]) | (layer6_outputs[1783]);
    assign outputs[1767] = layer6_outputs[1591];
    assign outputs[1768] = layer6_outputs[4629];
    assign outputs[1769] = layer6_outputs[2709];
    assign outputs[1770] = ~(layer6_outputs[1075]);
    assign outputs[1771] = ~(layer6_outputs[85]);
    assign outputs[1772] = layer6_outputs[3808];
    assign outputs[1773] = layer6_outputs[4085];
    assign outputs[1774] = ~(layer6_outputs[3765]) | (layer6_outputs[3194]);
    assign outputs[1775] = ~((layer6_outputs[1656]) ^ (layer6_outputs[1217]));
    assign outputs[1776] = ~(layer6_outputs[853]);
    assign outputs[1777] = ~((layer6_outputs[647]) | (layer6_outputs[3707]));
    assign outputs[1778] = ~(layer6_outputs[3793]);
    assign outputs[1779] = layer6_outputs[1658];
    assign outputs[1780] = ~(layer6_outputs[244]);
    assign outputs[1781] = layer6_outputs[4744];
    assign outputs[1782] = ~(layer6_outputs[1729]);
    assign outputs[1783] = ~(layer6_outputs[3898]);
    assign outputs[1784] = (layer6_outputs[2443]) ^ (layer6_outputs[5058]);
    assign outputs[1785] = layer6_outputs[2076];
    assign outputs[1786] = ~(layer6_outputs[2957]);
    assign outputs[1787] = ~(layer6_outputs[799]);
    assign outputs[1788] = ~((layer6_outputs[2728]) ^ (layer6_outputs[4230]));
    assign outputs[1789] = ~(layer6_outputs[1839]) | (layer6_outputs[4193]);
    assign outputs[1790] = (layer6_outputs[985]) & ~(layer6_outputs[2458]);
    assign outputs[1791] = ~(layer6_outputs[3601]) | (layer6_outputs[4943]);
    assign outputs[1792] = ~((layer6_outputs[5090]) ^ (layer6_outputs[3996]));
    assign outputs[1793] = ~(layer6_outputs[1484]);
    assign outputs[1794] = layer6_outputs[1620];
    assign outputs[1795] = ~(layer6_outputs[2394]);
    assign outputs[1796] = ~((layer6_outputs[4595]) | (layer6_outputs[2053]));
    assign outputs[1797] = ~(layer6_outputs[4644]);
    assign outputs[1798] = ~(layer6_outputs[1345]);
    assign outputs[1799] = layer6_outputs[3690];
    assign outputs[1800] = layer6_outputs[446];
    assign outputs[1801] = ~(layer6_outputs[171]);
    assign outputs[1802] = (layer6_outputs[3375]) ^ (layer6_outputs[2408]);
    assign outputs[1803] = layer6_outputs[1077];
    assign outputs[1804] = ~(layer6_outputs[3161]);
    assign outputs[1805] = layer6_outputs[1667];
    assign outputs[1806] = ~((layer6_outputs[3719]) ^ (layer6_outputs[2033]));
    assign outputs[1807] = layer6_outputs[3119];
    assign outputs[1808] = ~(layer6_outputs[4614]);
    assign outputs[1809] = ~(layer6_outputs[4641]);
    assign outputs[1810] = ~(layer6_outputs[465]);
    assign outputs[1811] = ~(layer6_outputs[1547]);
    assign outputs[1812] = layer6_outputs[2460];
    assign outputs[1813] = ~((layer6_outputs[2437]) ^ (layer6_outputs[1774]));
    assign outputs[1814] = ~(layer6_outputs[3953]);
    assign outputs[1815] = (layer6_outputs[3573]) ^ (layer6_outputs[360]);
    assign outputs[1816] = (layer6_outputs[53]) & ~(layer6_outputs[2001]);
    assign outputs[1817] = ~(layer6_outputs[4954]);
    assign outputs[1818] = layer6_outputs[2741];
    assign outputs[1819] = layer6_outputs[1492];
    assign outputs[1820] = layer6_outputs[444];
    assign outputs[1821] = ~(layer6_outputs[3019]);
    assign outputs[1822] = layer6_outputs[4400];
    assign outputs[1823] = layer6_outputs[4704];
    assign outputs[1824] = layer6_outputs[4745];
    assign outputs[1825] = (layer6_outputs[3762]) & ~(layer6_outputs[2671]);
    assign outputs[1826] = ~(layer6_outputs[825]) | (layer6_outputs[2502]);
    assign outputs[1827] = (layer6_outputs[1582]) ^ (layer6_outputs[965]);
    assign outputs[1828] = ~(layer6_outputs[2186]);
    assign outputs[1829] = (layer6_outputs[4827]) ^ (layer6_outputs[4041]);
    assign outputs[1830] = ~(layer6_outputs[3107]);
    assign outputs[1831] = layer6_outputs[4040];
    assign outputs[1832] = layer6_outputs[2810];
    assign outputs[1833] = (layer6_outputs[3518]) & (layer6_outputs[4667]);
    assign outputs[1834] = (layer6_outputs[250]) ^ (layer6_outputs[332]);
    assign outputs[1835] = ~(layer6_outputs[3943]);
    assign outputs[1836] = ~(layer6_outputs[5031]);
    assign outputs[1837] = ~((layer6_outputs[4060]) | (layer6_outputs[3696]));
    assign outputs[1838] = ~(layer6_outputs[3502]);
    assign outputs[1839] = ~((layer6_outputs[1399]) | (layer6_outputs[4275]));
    assign outputs[1840] = layer6_outputs[2291];
    assign outputs[1841] = (layer6_outputs[1422]) ^ (layer6_outputs[3665]);
    assign outputs[1842] = ~(layer6_outputs[1862]);
    assign outputs[1843] = ~(layer6_outputs[2072]);
    assign outputs[1844] = ~((layer6_outputs[3864]) ^ (layer6_outputs[3748]));
    assign outputs[1845] = layer6_outputs[1015];
    assign outputs[1846] = ~(layer6_outputs[1778]);
    assign outputs[1847] = (layer6_outputs[2753]) ^ (layer6_outputs[4187]);
    assign outputs[1848] = (layer6_outputs[331]) & ~(layer6_outputs[958]);
    assign outputs[1849] = ~(layer6_outputs[715]);
    assign outputs[1850] = layer6_outputs[4596];
    assign outputs[1851] = layer6_outputs[4237];
    assign outputs[1852] = layer6_outputs[2692];
    assign outputs[1853] = ~(layer6_outputs[2431]);
    assign outputs[1854] = layer6_outputs[3747];
    assign outputs[1855] = layer6_outputs[555];
    assign outputs[1856] = ~((layer6_outputs[4046]) ^ (layer6_outputs[3063]));
    assign outputs[1857] = ~(layer6_outputs[4507]);
    assign outputs[1858] = (layer6_outputs[2573]) ^ (layer6_outputs[4572]);
    assign outputs[1859] = layer6_outputs[1182];
    assign outputs[1860] = layer6_outputs[4981];
    assign outputs[1861] = ~(layer6_outputs[760]);
    assign outputs[1862] = ~(layer6_outputs[3252]);
    assign outputs[1863] = layer6_outputs[1833];
    assign outputs[1864] = layer6_outputs[3866];
    assign outputs[1865] = layer6_outputs[4055];
    assign outputs[1866] = ~(layer6_outputs[3966]);
    assign outputs[1867] = (layer6_outputs[780]) ^ (layer6_outputs[4451]);
    assign outputs[1868] = ~(layer6_outputs[3479]);
    assign outputs[1869] = (layer6_outputs[2432]) & ~(layer6_outputs[3562]);
    assign outputs[1870] = layer6_outputs[2474];
    assign outputs[1871] = ~((layer6_outputs[4893]) ^ (layer6_outputs[3975]));
    assign outputs[1872] = layer6_outputs[537];
    assign outputs[1873] = ~(layer6_outputs[3787]);
    assign outputs[1874] = ~(layer6_outputs[1382]);
    assign outputs[1875] = ~(layer6_outputs[2874]);
    assign outputs[1876] = layer6_outputs[2918];
    assign outputs[1877] = layer6_outputs[3977];
    assign outputs[1878] = layer6_outputs[212];
    assign outputs[1879] = layer6_outputs[1677];
    assign outputs[1880] = ~(layer6_outputs[633]);
    assign outputs[1881] = layer6_outputs[3342];
    assign outputs[1882] = layer6_outputs[1973];
    assign outputs[1883] = ~((layer6_outputs[2706]) ^ (layer6_outputs[2097]));
    assign outputs[1884] = ~((layer6_outputs[4721]) ^ (layer6_outputs[4297]));
    assign outputs[1885] = ~(layer6_outputs[792]) | (layer6_outputs[2376]);
    assign outputs[1886] = ~(layer6_outputs[5022]);
    assign outputs[1887] = ~((layer6_outputs[1311]) | (layer6_outputs[4752]));
    assign outputs[1888] = ~((layer6_outputs[1357]) ^ (layer6_outputs[765]));
    assign outputs[1889] = ~(layer6_outputs[33]);
    assign outputs[1890] = layer6_outputs[4647];
    assign outputs[1891] = layer6_outputs[3994];
    assign outputs[1892] = (layer6_outputs[1989]) ^ (layer6_outputs[4111]);
    assign outputs[1893] = layer6_outputs[5004];
    assign outputs[1894] = ~((layer6_outputs[4516]) | (layer6_outputs[4830]));
    assign outputs[1895] = (layer6_outputs[96]) ^ (layer6_outputs[3482]);
    assign outputs[1896] = layer6_outputs[4137];
    assign outputs[1897] = ~(layer6_outputs[4923]);
    assign outputs[1898] = layer6_outputs[3949];
    assign outputs[1899] = layer6_outputs[1557];
    assign outputs[1900] = layer6_outputs[4167];
    assign outputs[1901] = layer6_outputs[1141];
    assign outputs[1902] = layer6_outputs[1936];
    assign outputs[1903] = ~(layer6_outputs[2126]);
    assign outputs[1904] = ~((layer6_outputs[4032]) ^ (layer6_outputs[4602]));
    assign outputs[1905] = layer6_outputs[3355];
    assign outputs[1906] = layer6_outputs[1166];
    assign outputs[1907] = ~(layer6_outputs[4175]);
    assign outputs[1908] = ~(layer6_outputs[1117]);
    assign outputs[1909] = ~(layer6_outputs[3948]);
    assign outputs[1910] = layer6_outputs[4730];
    assign outputs[1911] = layer6_outputs[1307];
    assign outputs[1912] = layer6_outputs[4591];
    assign outputs[1913] = ~(layer6_outputs[3091]);
    assign outputs[1914] = layer6_outputs[4209];
    assign outputs[1915] = ~(layer6_outputs[2411]);
    assign outputs[1916] = (layer6_outputs[1492]) & (layer6_outputs[790]);
    assign outputs[1917] = layer6_outputs[2965];
    assign outputs[1918] = ~(layer6_outputs[4834]);
    assign outputs[1919] = ~(layer6_outputs[4639]);
    assign outputs[1920] = ~((layer6_outputs[5093]) | (layer6_outputs[3229]));
    assign outputs[1921] = layer6_outputs[3186];
    assign outputs[1922] = layer6_outputs[3050];
    assign outputs[1923] = ~(layer6_outputs[3704]);
    assign outputs[1924] = layer6_outputs[4122];
    assign outputs[1925] = layer6_outputs[2511];
    assign outputs[1926] = layer6_outputs[2237];
    assign outputs[1927] = layer6_outputs[3173];
    assign outputs[1928] = ~(layer6_outputs[3486]);
    assign outputs[1929] = layer6_outputs[4636];
    assign outputs[1930] = ~((layer6_outputs[2650]) ^ (layer6_outputs[2449]));
    assign outputs[1931] = layer6_outputs[930];
    assign outputs[1932] = ~(layer6_outputs[1972]);
    assign outputs[1933] = ~((layer6_outputs[2051]) & (layer6_outputs[661]));
    assign outputs[1934] = ~(layer6_outputs[2165]) | (layer6_outputs[214]);
    assign outputs[1935] = layer6_outputs[539];
    assign outputs[1936] = ~((layer6_outputs[677]) ^ (layer6_outputs[2131]));
    assign outputs[1937] = ~(layer6_outputs[1253]);
    assign outputs[1938] = ~(layer6_outputs[4829]);
    assign outputs[1939] = ~((layer6_outputs[2182]) ^ (layer6_outputs[2326]));
    assign outputs[1940] = ~(layer6_outputs[2966]);
    assign outputs[1941] = ~(layer6_outputs[2421]);
    assign outputs[1942] = ~(layer6_outputs[560]) | (layer6_outputs[4303]);
    assign outputs[1943] = ~((layer6_outputs[1054]) ^ (layer6_outputs[3560]));
    assign outputs[1944] = layer6_outputs[1303];
    assign outputs[1945] = ~((layer6_outputs[319]) | (layer6_outputs[3315]));
    assign outputs[1946] = layer6_outputs[844];
    assign outputs[1947] = layer6_outputs[3602];
    assign outputs[1948] = ~((layer6_outputs[1760]) ^ (layer6_outputs[2025]));
    assign outputs[1949] = layer6_outputs[199];
    assign outputs[1950] = ~((layer6_outputs[1871]) | (layer6_outputs[1712]));
    assign outputs[1951] = ~(layer6_outputs[323]);
    assign outputs[1952] = layer6_outputs[4705];
    assign outputs[1953] = ~(layer6_outputs[4807]);
    assign outputs[1954] = layer6_outputs[2700];
    assign outputs[1955] = ~(layer6_outputs[132]);
    assign outputs[1956] = layer6_outputs[2772];
    assign outputs[1957] = (layer6_outputs[3792]) & (layer6_outputs[1633]);
    assign outputs[1958] = ~(layer6_outputs[4779]);
    assign outputs[1959] = layer6_outputs[318];
    assign outputs[1960] = ~(layer6_outputs[1822]);
    assign outputs[1961] = layer6_outputs[1663];
    assign outputs[1962] = ~((layer6_outputs[3529]) | (layer6_outputs[538]));
    assign outputs[1963] = (layer6_outputs[2933]) ^ (layer6_outputs[252]);
    assign outputs[1964] = ~((layer6_outputs[5040]) ^ (layer6_outputs[306]));
    assign outputs[1965] = ~(layer6_outputs[3237]);
    assign outputs[1966] = ~(layer6_outputs[2684]);
    assign outputs[1967] = ~((layer6_outputs[1145]) ^ (layer6_outputs[666]));
    assign outputs[1968] = layer6_outputs[2878];
    assign outputs[1969] = ~(layer6_outputs[4851]);
    assign outputs[1970] = layer6_outputs[290];
    assign outputs[1971] = ~(layer6_outputs[339]);
    assign outputs[1972] = ~(layer6_outputs[4862]);
    assign outputs[1973] = layer6_outputs[1974];
    assign outputs[1974] = ~(layer6_outputs[2028]);
    assign outputs[1975] = ~(layer6_outputs[761]);
    assign outputs[1976] = (layer6_outputs[693]) ^ (layer6_outputs[1076]);
    assign outputs[1977] = ~((layer6_outputs[3260]) | (layer6_outputs[4481]));
    assign outputs[1978] = layer6_outputs[5051];
    assign outputs[1979] = layer6_outputs[967];
    assign outputs[1980] = (layer6_outputs[2732]) & (layer6_outputs[4174]);
    assign outputs[1981] = layer6_outputs[2822];
    assign outputs[1982] = layer6_outputs[2210];
    assign outputs[1983] = layer6_outputs[5081];
    assign outputs[1984] = layer6_outputs[13];
    assign outputs[1985] = ~((layer6_outputs[1540]) ^ (layer6_outputs[1366]));
    assign outputs[1986] = ~(layer6_outputs[2161]);
    assign outputs[1987] = ~(layer6_outputs[4087]);
    assign outputs[1988] = layer6_outputs[3289];
    assign outputs[1989] = ~(layer6_outputs[4157]);
    assign outputs[1990] = layer6_outputs[200];
    assign outputs[1991] = layer6_outputs[3320];
    assign outputs[1992] = (layer6_outputs[3220]) ^ (layer6_outputs[3265]);
    assign outputs[1993] = layer6_outputs[4449];
    assign outputs[1994] = layer6_outputs[904];
    assign outputs[1995] = ~(layer6_outputs[3770]);
    assign outputs[1996] = layer6_outputs[3119];
    assign outputs[1997] = (layer6_outputs[3273]) & ~(layer6_outputs[3668]);
    assign outputs[1998] = layer6_outputs[3377];
    assign outputs[1999] = layer6_outputs[1990];
    assign outputs[2000] = ~(layer6_outputs[2970]);
    assign outputs[2001] = layer6_outputs[5003];
    assign outputs[2002] = ~(layer6_outputs[4685]);
    assign outputs[2003] = layer6_outputs[1443];
    assign outputs[2004] = ~((layer6_outputs[2420]) ^ (layer6_outputs[3910]));
    assign outputs[2005] = layer6_outputs[1330];
    assign outputs[2006] = ~((layer6_outputs[1343]) ^ (layer6_outputs[3215]));
    assign outputs[2007] = ~((layer6_outputs[1267]) & (layer6_outputs[2258]));
    assign outputs[2008] = ~(layer6_outputs[1085]);
    assign outputs[2009] = ~(layer6_outputs[3540]);
    assign outputs[2010] = ~(layer6_outputs[4641]);
    assign outputs[2011] = layer6_outputs[3148];
    assign outputs[2012] = ~((layer6_outputs[4456]) ^ (layer6_outputs[4199]));
    assign outputs[2013] = ~((layer6_outputs[1162]) ^ (layer6_outputs[1246]));
    assign outputs[2014] = ~(layer6_outputs[3262]);
    assign outputs[2015] = ~((layer6_outputs[2130]) ^ (layer6_outputs[2974]));
    assign outputs[2016] = layer6_outputs[2866];
    assign outputs[2017] = ~((layer6_outputs[356]) ^ (layer6_outputs[3176]));
    assign outputs[2018] = (layer6_outputs[4037]) & ~(layer6_outputs[1192]);
    assign outputs[2019] = layer6_outputs[2569];
    assign outputs[2020] = (layer6_outputs[3832]) & ~(layer6_outputs[3316]);
    assign outputs[2021] = ~((layer6_outputs[2390]) ^ (layer6_outputs[2992]));
    assign outputs[2022] = ~((layer6_outputs[51]) ^ (layer6_outputs[832]));
    assign outputs[2023] = ~(layer6_outputs[4358]);
    assign outputs[2024] = ~(layer6_outputs[585]);
    assign outputs[2025] = ~(layer6_outputs[2465]);
    assign outputs[2026] = ~(layer6_outputs[3381]);
    assign outputs[2027] = (layer6_outputs[4620]) ^ (layer6_outputs[3978]);
    assign outputs[2028] = ~(layer6_outputs[4145]);
    assign outputs[2029] = ~(layer6_outputs[4333]);
    assign outputs[2030] = layer6_outputs[312];
    assign outputs[2031] = layer6_outputs[2963];
    assign outputs[2032] = layer6_outputs[1817];
    assign outputs[2033] = ~(layer6_outputs[3663]);
    assign outputs[2034] = ~(layer6_outputs[1151]);
    assign outputs[2035] = (layer6_outputs[4500]) | (layer6_outputs[3645]);
    assign outputs[2036] = layer6_outputs[4582];
    assign outputs[2037] = ~((layer6_outputs[4184]) | (layer6_outputs[711]));
    assign outputs[2038] = (layer6_outputs[74]) ^ (layer6_outputs[113]);
    assign outputs[2039] = layer6_outputs[3520];
    assign outputs[2040] = ~((layer6_outputs[441]) ^ (layer6_outputs[2067]));
    assign outputs[2041] = ~(layer6_outputs[3892]);
    assign outputs[2042] = (layer6_outputs[1951]) & ~(layer6_outputs[3559]);
    assign outputs[2043] = ~(layer6_outputs[28]) | (layer6_outputs[4056]);
    assign outputs[2044] = ~(layer6_outputs[813]);
    assign outputs[2045] = ~(layer6_outputs[4394]);
    assign outputs[2046] = ~(layer6_outputs[774]) | (layer6_outputs[2804]);
    assign outputs[2047] = (layer6_outputs[2787]) ^ (layer6_outputs[4223]);
    assign outputs[2048] = (layer6_outputs[1591]) & (layer6_outputs[1946]);
    assign outputs[2049] = (layer6_outputs[2661]) & ~(layer6_outputs[190]);
    assign outputs[2050] = layer6_outputs[1265];
    assign outputs[2051] = ~(layer6_outputs[3383]);
    assign outputs[2052] = layer6_outputs[2956];
    assign outputs[2053] = ~(layer6_outputs[283]);
    assign outputs[2054] = ~(layer6_outputs[3841]);
    assign outputs[2055] = ~((layer6_outputs[4136]) | (layer6_outputs[2073]));
    assign outputs[2056] = ~(layer6_outputs[2351]);
    assign outputs[2057] = layer6_outputs[701];
    assign outputs[2058] = (layer6_outputs[1994]) ^ (layer6_outputs[2270]);
    assign outputs[2059] = (layer6_outputs[316]) & (layer6_outputs[2299]);
    assign outputs[2060] = (layer6_outputs[816]) & ~(layer6_outputs[3688]);
    assign outputs[2061] = ~(layer6_outputs[2235]) | (layer6_outputs[2659]);
    assign outputs[2062] = ~((layer6_outputs[2592]) | (layer6_outputs[101]));
    assign outputs[2063] = layer6_outputs[770];
    assign outputs[2064] = ~(layer6_outputs[4630]);
    assign outputs[2065] = layer6_outputs[866];
    assign outputs[2066] = ~(layer6_outputs[3582]) | (layer6_outputs[1052]);
    assign outputs[2067] = ~(layer6_outputs[1917]);
    assign outputs[2068] = layer6_outputs[2240];
    assign outputs[2069] = layer6_outputs[1496];
    assign outputs[2070] = layer6_outputs[1978];
    assign outputs[2071] = ~(layer6_outputs[85]);
    assign outputs[2072] = (layer6_outputs[4710]) ^ (layer6_outputs[755]);
    assign outputs[2073] = ~(layer6_outputs[3983]);
    assign outputs[2074] = layer6_outputs[82];
    assign outputs[2075] = ~(layer6_outputs[4599]);
    assign outputs[2076] = layer6_outputs[1412];
    assign outputs[2077] = (layer6_outputs[1827]) ^ (layer6_outputs[2820]);
    assign outputs[2078] = (layer6_outputs[1034]) & ~(layer6_outputs[3992]);
    assign outputs[2079] = (layer6_outputs[2200]) & (layer6_outputs[4520]);
    assign outputs[2080] = ~(layer6_outputs[5033]);
    assign outputs[2081] = layer6_outputs[1155];
    assign outputs[2082] = layer6_outputs[2027];
    assign outputs[2083] = ~(layer6_outputs[3013]);
    assign outputs[2084] = layer6_outputs[4115];
    assign outputs[2085] = layer6_outputs[2983];
    assign outputs[2086] = ~((layer6_outputs[3582]) ^ (layer6_outputs[2826]));
    assign outputs[2087] = (layer6_outputs[5073]) & ~(layer6_outputs[803]);
    assign outputs[2088] = layer6_outputs[4462];
    assign outputs[2089] = ~(layer6_outputs[3588]);
    assign outputs[2090] = (layer6_outputs[4404]) ^ (layer6_outputs[3457]);
    assign outputs[2091] = layer6_outputs[1488];
    assign outputs[2092] = (layer6_outputs[2036]) & (layer6_outputs[1537]);
    assign outputs[2093] = layer6_outputs[3700];
    assign outputs[2094] = layer6_outputs[4155];
    assign outputs[2095] = layer6_outputs[1726];
    assign outputs[2096] = (layer6_outputs[1852]) | (layer6_outputs[4952]);
    assign outputs[2097] = ~(layer6_outputs[2904]);
    assign outputs[2098] = ~((layer6_outputs[4404]) ^ (layer6_outputs[2347]));
    assign outputs[2099] = (layer6_outputs[2653]) & ~(layer6_outputs[1609]);
    assign outputs[2100] = (layer6_outputs[1036]) ^ (layer6_outputs[712]);
    assign outputs[2101] = layer6_outputs[4793];
    assign outputs[2102] = ~((layer6_outputs[1141]) ^ (layer6_outputs[327]));
    assign outputs[2103] = ~(layer6_outputs[1227]) | (layer6_outputs[1183]);
    assign outputs[2104] = ~(layer6_outputs[4341]);
    assign outputs[2105] = (layer6_outputs[1901]) ^ (layer6_outputs[4952]);
    assign outputs[2106] = layer6_outputs[4288];
    assign outputs[2107] = layer6_outputs[43];
    assign outputs[2108] = layer6_outputs[4959];
    assign outputs[2109] = ~(layer6_outputs[1350]);
    assign outputs[2110] = layer6_outputs[5094];
    assign outputs[2111] = layer6_outputs[1454];
    assign outputs[2112] = ~((layer6_outputs[1114]) | (layer6_outputs[2239]));
    assign outputs[2113] = ~(layer6_outputs[1690]);
    assign outputs[2114] = layer6_outputs[2035];
    assign outputs[2115] = layer6_outputs[4183];
    assign outputs[2116] = ~(layer6_outputs[4794]);
    assign outputs[2117] = ~(layer6_outputs[3779]) | (layer6_outputs[2972]);
    assign outputs[2118] = ~(layer6_outputs[4826]);
    assign outputs[2119] = ~(layer6_outputs[1486]) | (layer6_outputs[1660]);
    assign outputs[2120] = ~((layer6_outputs[2303]) ^ (layer6_outputs[2101]));
    assign outputs[2121] = layer6_outputs[2777];
    assign outputs[2122] = ~(layer6_outputs[340]);
    assign outputs[2123] = layer6_outputs[1624];
    assign outputs[2124] = ~(layer6_outputs[3901]) | (layer6_outputs[3339]);
    assign outputs[2125] = layer6_outputs[2013];
    assign outputs[2126] = layer6_outputs[3465];
    assign outputs[2127] = ~(layer6_outputs[980]);
    assign outputs[2128] = ~(layer6_outputs[526]);
    assign outputs[2129] = ~((layer6_outputs[4649]) ^ (layer6_outputs[4208]));
    assign outputs[2130] = layer6_outputs[1968];
    assign outputs[2131] = layer6_outputs[2669];
    assign outputs[2132] = ~(layer6_outputs[1153]);
    assign outputs[2133] = ~(layer6_outputs[4438]) | (layer6_outputs[2091]);
    assign outputs[2134] = (layer6_outputs[1673]) & ~(layer6_outputs[251]);
    assign outputs[2135] = (layer6_outputs[380]) ^ (layer6_outputs[3708]);
    assign outputs[2136] = layer6_outputs[1210];
    assign outputs[2137] = ~((layer6_outputs[2242]) ^ (layer6_outputs[1383]));
    assign outputs[2138] = ~(layer6_outputs[3323]);
    assign outputs[2139] = ~(layer6_outputs[3049]);
    assign outputs[2140] = ~(layer6_outputs[2857]);
    assign outputs[2141] = layer6_outputs[478];
    assign outputs[2142] = (layer6_outputs[1195]) & ~(layer6_outputs[5069]);
    assign outputs[2143] = ~(layer6_outputs[1274]);
    assign outputs[2144] = ~((layer6_outputs[2115]) ^ (layer6_outputs[3278]));
    assign outputs[2145] = (layer6_outputs[2020]) & ~(layer6_outputs[4004]);
    assign outputs[2146] = ~(layer6_outputs[4134]);
    assign outputs[2147] = (layer6_outputs[262]) & ~(layer6_outputs[2762]);
    assign outputs[2148] = layer6_outputs[4216];
    assign outputs[2149] = ~(layer6_outputs[1847]) | (layer6_outputs[4076]);
    assign outputs[2150] = ~((layer6_outputs[1245]) ^ (layer6_outputs[1066]));
    assign outputs[2151] = ~(layer6_outputs[2490]);
    assign outputs[2152] = (layer6_outputs[3828]) & ~(layer6_outputs[4110]);
    assign outputs[2153] = layer6_outputs[4053];
    assign outputs[2154] = (layer6_outputs[5014]) & ~(layer6_outputs[1424]);
    assign outputs[2155] = ~((layer6_outputs[2172]) ^ (layer6_outputs[2587]));
    assign outputs[2156] = layer6_outputs[4267];
    assign outputs[2157] = ~(layer6_outputs[2535]);
    assign outputs[2158] = ~((layer6_outputs[2964]) ^ (layer6_outputs[4602]));
    assign outputs[2159] = layer6_outputs[1357];
    assign outputs[2160] = ~(layer6_outputs[4395]) | (layer6_outputs[156]);
    assign outputs[2161] = layer6_outputs[221];
    assign outputs[2162] = (layer6_outputs[2025]) ^ (layer6_outputs[298]);
    assign outputs[2163] = (layer6_outputs[4100]) & ~(layer6_outputs[5103]);
    assign outputs[2164] = ~(layer6_outputs[195]);
    assign outputs[2165] = ~(layer6_outputs[842]);
    assign outputs[2166] = ~((layer6_outputs[3111]) ^ (layer6_outputs[2592]));
    assign outputs[2167] = (layer6_outputs[4092]) ^ (layer6_outputs[3423]);
    assign outputs[2168] = ~((layer6_outputs[4836]) ^ (layer6_outputs[3576]));
    assign outputs[2169] = ~(layer6_outputs[1794]);
    assign outputs[2170] = ~(layer6_outputs[1067]);
    assign outputs[2171] = ~(layer6_outputs[322]);
    assign outputs[2172] = ~(layer6_outputs[426]);
    assign outputs[2173] = layer6_outputs[188];
    assign outputs[2174] = ~(layer6_outputs[3592]);
    assign outputs[2175] = (layer6_outputs[2924]) ^ (layer6_outputs[3904]);
    assign outputs[2176] = layer6_outputs[3729];
    assign outputs[2177] = ~((layer6_outputs[3605]) | (layer6_outputs[4724]));
    assign outputs[2178] = layer6_outputs[883];
    assign outputs[2179] = (layer6_outputs[772]) ^ (layer6_outputs[3439]);
    assign outputs[2180] = ~(layer6_outputs[3782]);
    assign outputs[2181] = layer6_outputs[2548];
    assign outputs[2182] = ~(layer6_outputs[79]);
    assign outputs[2183] = layer6_outputs[3993];
    assign outputs[2184] = ~(layer6_outputs[1090]);
    assign outputs[2185] = (layer6_outputs[4392]) ^ (layer6_outputs[4014]);
    assign outputs[2186] = ~((layer6_outputs[4756]) | (layer6_outputs[3211]));
    assign outputs[2187] = layer6_outputs[3364];
    assign outputs[2188] = (layer6_outputs[3036]) & ~(layer6_outputs[4469]);
    assign outputs[2189] = layer6_outputs[2459];
    assign outputs[2190] = ~(layer6_outputs[38]);
    assign outputs[2191] = ~((layer6_outputs[3178]) ^ (layer6_outputs[721]));
    assign outputs[2192] = ~(layer6_outputs[2267]);
    assign outputs[2193] = ~(layer6_outputs[4167]);
    assign outputs[2194] = (layer6_outputs[4248]) & ~(layer6_outputs[2769]);
    assign outputs[2195] = ~(layer6_outputs[4510]);
    assign outputs[2196] = ~(layer6_outputs[4143]);
    assign outputs[2197] = layer6_outputs[3222];
    assign outputs[2198] = layer6_outputs[2464];
    assign outputs[2199] = ~(layer6_outputs[968]);
    assign outputs[2200] = ~(layer6_outputs[3221]);
    assign outputs[2201] = (layer6_outputs[4179]) & ~(layer6_outputs[3277]);
    assign outputs[2202] = (layer6_outputs[2755]) ^ (layer6_outputs[4906]);
    assign outputs[2203] = (layer6_outputs[4399]) ^ (layer6_outputs[2238]);
    assign outputs[2204] = layer6_outputs[4633];
    assign outputs[2205] = layer6_outputs[5023];
    assign outputs[2206] = (layer6_outputs[2223]) & (layer6_outputs[856]);
    assign outputs[2207] = ~(layer6_outputs[3005]);
    assign outputs[2208] = layer6_outputs[3963];
    assign outputs[2209] = ~(layer6_outputs[3234]);
    assign outputs[2210] = ~(layer6_outputs[4101]);
    assign outputs[2211] = layer6_outputs[2700];
    assign outputs[2212] = layer6_outputs[4014];
    assign outputs[2213] = ~(layer6_outputs[4126]);
    assign outputs[2214] = ~(layer6_outputs[364]);
    assign outputs[2215] = ~((layer6_outputs[2192]) ^ (layer6_outputs[1709]));
    assign outputs[2216] = layer6_outputs[3851];
    assign outputs[2217] = layer6_outputs[763];
    assign outputs[2218] = ~(layer6_outputs[2007]);
    assign outputs[2219] = layer6_outputs[3831];
    assign outputs[2220] = ~(layer6_outputs[9]);
    assign outputs[2221] = ~(layer6_outputs[2480]);
    assign outputs[2222] = (layer6_outputs[740]) ^ (layer6_outputs[828]);
    assign outputs[2223] = ~((layer6_outputs[54]) & (layer6_outputs[1824]));
    assign outputs[2224] = ~(layer6_outputs[1131]);
    assign outputs[2225] = ~(layer6_outputs[1261]);
    assign outputs[2226] = layer6_outputs[1374];
    assign outputs[2227] = (layer6_outputs[4557]) & ~(layer6_outputs[1782]);
    assign outputs[2228] = ~(layer6_outputs[4965]);
    assign outputs[2229] = ~(layer6_outputs[4677]);
    assign outputs[2230] = ~(layer6_outputs[575]);
    assign outputs[2231] = (layer6_outputs[1975]) ^ (layer6_outputs[545]);
    assign outputs[2232] = ~(layer6_outputs[3633]);
    assign outputs[2233] = ~(layer6_outputs[2082]);
    assign outputs[2234] = ~(layer6_outputs[4984]);
    assign outputs[2235] = ~(layer6_outputs[4093]);
    assign outputs[2236] = layer6_outputs[1176];
    assign outputs[2237] = layer6_outputs[3529];
    assign outputs[2238] = layer6_outputs[4182];
    assign outputs[2239] = ~(layer6_outputs[1844]);
    assign outputs[2240] = layer6_outputs[1483];
    assign outputs[2241] = layer6_outputs[5051];
    assign outputs[2242] = ~((layer6_outputs[2182]) ^ (layer6_outputs[4208]));
    assign outputs[2243] = layer6_outputs[873];
    assign outputs[2244] = ~(layer6_outputs[3160]);
    assign outputs[2245] = layer6_outputs[4691];
    assign outputs[2246] = layer6_outputs[46];
    assign outputs[2247] = ~(layer6_outputs[226]);
    assign outputs[2248] = ~(layer6_outputs[2256]);
    assign outputs[2249] = layer6_outputs[3228];
    assign outputs[2250] = layer6_outputs[3269];
    assign outputs[2251] = layer6_outputs[846];
    assign outputs[2252] = ~(layer6_outputs[3130]);
    assign outputs[2253] = ~(layer6_outputs[2843]);
    assign outputs[2254] = layer6_outputs[4396];
    assign outputs[2255] = (layer6_outputs[3028]) & ~(layer6_outputs[1771]);
    assign outputs[2256] = layer6_outputs[521];
    assign outputs[2257] = (layer6_outputs[4945]) & ~(layer6_outputs[4697]);
    assign outputs[2258] = layer6_outputs[1125];
    assign outputs[2259] = layer6_outputs[813];
    assign outputs[2260] = layer6_outputs[770];
    assign outputs[2261] = ~(layer6_outputs[3783]);
    assign outputs[2262] = ~((layer6_outputs[3715]) ^ (layer6_outputs[169]));
    assign outputs[2263] = ~(layer6_outputs[2827]);
    assign outputs[2264] = (layer6_outputs[2203]) & (layer6_outputs[3868]);
    assign outputs[2265] = layer6_outputs[1586];
    assign outputs[2266] = layer6_outputs[1340];
    assign outputs[2267] = ~(layer6_outputs[3964]);
    assign outputs[2268] = ~((layer6_outputs[4399]) ^ (layer6_outputs[943]));
    assign outputs[2269] = ~(layer6_outputs[1333]);
    assign outputs[2270] = (layer6_outputs[4242]) & ~(layer6_outputs[315]);
    assign outputs[2271] = layer6_outputs[4854];
    assign outputs[2272] = (layer6_outputs[1849]) ^ (layer6_outputs[1873]);
    assign outputs[2273] = (layer6_outputs[2670]) ^ (layer6_outputs[3296]);
    assign outputs[2274] = layer6_outputs[3037];
    assign outputs[2275] = ~(layer6_outputs[2333]) | (layer6_outputs[3067]);
    assign outputs[2276] = layer6_outputs[215];
    assign outputs[2277] = layer6_outputs[220];
    assign outputs[2278] = ~(layer6_outputs[1489]);
    assign outputs[2279] = ~(layer6_outputs[1566]) | (layer6_outputs[466]);
    assign outputs[2280] = (layer6_outputs[4759]) & ~(layer6_outputs[3740]);
    assign outputs[2281] = layer6_outputs[2754];
    assign outputs[2282] = ~(layer6_outputs[7]);
    assign outputs[2283] = layer6_outputs[4171];
    assign outputs[2284] = (layer6_outputs[1045]) ^ (layer6_outputs[4385]);
    assign outputs[2285] = (layer6_outputs[1887]) & (layer6_outputs[2011]);
    assign outputs[2286] = (layer6_outputs[1371]) ^ (layer6_outputs[1575]);
    assign outputs[2287] = ~(layer6_outputs[437]);
    assign outputs[2288] = (layer6_outputs[3335]) ^ (layer6_outputs[4820]);
    assign outputs[2289] = (layer6_outputs[4956]) & ~(layer6_outputs[2858]);
    assign outputs[2290] = layer6_outputs[2171];
    assign outputs[2291] = ~(layer6_outputs[2904]);
    assign outputs[2292] = ~(layer6_outputs[2878]);
    assign outputs[2293] = (layer6_outputs[430]) & ~(layer6_outputs[4461]);
    assign outputs[2294] = layer6_outputs[1464];
    assign outputs[2295] = layer6_outputs[3981];
    assign outputs[2296] = layer6_outputs[71];
    assign outputs[2297] = layer6_outputs[2397];
    assign outputs[2298] = layer6_outputs[4536];
    assign outputs[2299] = ~(layer6_outputs[2328]);
    assign outputs[2300] = (layer6_outputs[321]) ^ (layer6_outputs[795]);
    assign outputs[2301] = (layer6_outputs[3013]) ^ (layer6_outputs[461]);
    assign outputs[2302] = (layer6_outputs[755]) & ~(layer6_outputs[1646]);
    assign outputs[2303] = layer6_outputs[791];
    assign outputs[2304] = ~(layer6_outputs[2893]);
    assign outputs[2305] = ~(layer6_outputs[4461]);
    assign outputs[2306] = ~(layer6_outputs[1314]);
    assign outputs[2307] = ~((layer6_outputs[4492]) ^ (layer6_outputs[2208]));
    assign outputs[2308] = (layer6_outputs[1219]) & ~(layer6_outputs[1296]);
    assign outputs[2309] = (layer6_outputs[757]) ^ (layer6_outputs[4005]);
    assign outputs[2310] = layer6_outputs[469];
    assign outputs[2311] = ~(layer6_outputs[4319]);
    assign outputs[2312] = ~(layer6_outputs[3116]);
    assign outputs[2313] = (layer6_outputs[4201]) & (layer6_outputs[4177]);
    assign outputs[2314] = layer6_outputs[4064];
    assign outputs[2315] = layer6_outputs[3789];
    assign outputs[2316] = layer6_outputs[3392];
    assign outputs[2317] = ~(layer6_outputs[942]);
    assign outputs[2318] = layer6_outputs[4430];
    assign outputs[2319] = layer6_outputs[1991];
    assign outputs[2320] = layer6_outputs[731];
    assign outputs[2321] = layer6_outputs[3207];
    assign outputs[2322] = ~(layer6_outputs[4408]);
    assign outputs[2323] = ~(layer6_outputs[4722]);
    assign outputs[2324] = (layer6_outputs[2172]) ^ (layer6_outputs[491]);
    assign outputs[2325] = layer6_outputs[584];
    assign outputs[2326] = (layer6_outputs[1853]) & ~(layer6_outputs[3921]);
    assign outputs[2327] = layer6_outputs[3412];
    assign outputs[2328] = layer6_outputs[2388];
    assign outputs[2329] = layer6_outputs[3197];
    assign outputs[2330] = layer6_outputs[1841];
    assign outputs[2331] = ~(layer6_outputs[3583]);
    assign outputs[2332] = layer6_outputs[2625];
    assign outputs[2333] = (layer6_outputs[631]) ^ (layer6_outputs[468]);
    assign outputs[2334] = 1'b0;
    assign outputs[2335] = ~(layer6_outputs[2959]);
    assign outputs[2336] = ~(layer6_outputs[2654]);
    assign outputs[2337] = layer6_outputs[2269];
    assign outputs[2338] = (layer6_outputs[2104]) ^ (layer6_outputs[4905]);
    assign outputs[2339] = layer6_outputs[4703];
    assign outputs[2340] = layer6_outputs[242];
    assign outputs[2341] = ~(layer6_outputs[4457]);
    assign outputs[2342] = ~(layer6_outputs[5057]);
    assign outputs[2343] = layer6_outputs[1353];
    assign outputs[2344] = ~(layer6_outputs[499]);
    assign outputs[2345] = layer6_outputs[871];
    assign outputs[2346] = layer6_outputs[4248];
    assign outputs[2347] = (layer6_outputs[2288]) & ~(layer6_outputs[5005]);
    assign outputs[2348] = layer6_outputs[3016];
    assign outputs[2349] = ~(layer6_outputs[3755]);
    assign outputs[2350] = (layer6_outputs[1878]) & (layer6_outputs[4518]);
    assign outputs[2351] = layer6_outputs[3945];
    assign outputs[2352] = ~((layer6_outputs[1053]) & (layer6_outputs[2867]));
    assign outputs[2353] = layer6_outputs[1316];
    assign outputs[2354] = ~(layer6_outputs[3343]);
    assign outputs[2355] = layer6_outputs[567];
    assign outputs[2356] = layer6_outputs[4765];
    assign outputs[2357] = (layer6_outputs[1696]) ^ (layer6_outputs[3677]);
    assign outputs[2358] = layer6_outputs[3972];
    assign outputs[2359] = layer6_outputs[2338];
    assign outputs[2360] = ~(layer6_outputs[5019]);
    assign outputs[2361] = layer6_outputs[3840];
    assign outputs[2362] = ~(layer6_outputs[2840]);
    assign outputs[2363] = layer6_outputs[3907];
    assign outputs[2364] = (layer6_outputs[4986]) & ~(layer6_outputs[1901]);
    assign outputs[2365] = layer6_outputs[3349];
    assign outputs[2366] = layer6_outputs[533];
    assign outputs[2367] = ~(layer6_outputs[3348]);
    assign outputs[2368] = layer6_outputs[560];
    assign outputs[2369] = ~(layer6_outputs[5043]) | (layer6_outputs[1202]);
    assign outputs[2370] = layer6_outputs[2726];
    assign outputs[2371] = (layer6_outputs[3653]) & (layer6_outputs[3429]);
    assign outputs[2372] = layer6_outputs[571];
    assign outputs[2373] = layer6_outputs[3953];
    assign outputs[2374] = ~(layer6_outputs[2845]);
    assign outputs[2375] = ~(layer6_outputs[1455]);
    assign outputs[2376] = ~(layer6_outputs[3125]);
    assign outputs[2377] = layer6_outputs[2464];
    assign outputs[2378] = layer6_outputs[3356];
    assign outputs[2379] = ~(layer6_outputs[556]);
    assign outputs[2380] = ~((layer6_outputs[1240]) ^ (layer6_outputs[3913]));
    assign outputs[2381] = ~(layer6_outputs[622]);
    assign outputs[2382] = (layer6_outputs[74]) & ~(layer6_outputs[3444]);
    assign outputs[2383] = layer6_outputs[856];
    assign outputs[2384] = layer6_outputs[1683];
    assign outputs[2385] = layer6_outputs[1155];
    assign outputs[2386] = ~((layer6_outputs[1466]) ^ (layer6_outputs[4715]));
    assign outputs[2387] = ~(layer6_outputs[4764]);
    assign outputs[2388] = (layer6_outputs[2542]) & ~(layer6_outputs[3266]);
    assign outputs[2389] = layer6_outputs[1885];
    assign outputs[2390] = ~((layer6_outputs[1574]) ^ (layer6_outputs[376]));
    assign outputs[2391] = (layer6_outputs[2708]) & ~(layer6_outputs[2243]);
    assign outputs[2392] = (layer6_outputs[2562]) & ~(layer6_outputs[2294]);
    assign outputs[2393] = ~(layer6_outputs[732]) | (layer6_outputs[700]);
    assign outputs[2394] = ~(layer6_outputs[4178]);
    assign outputs[2395] = layer6_outputs[121];
    assign outputs[2396] = ~(layer6_outputs[4138]);
    assign outputs[2397] = layer6_outputs[2958];
    assign outputs[2398] = ~(layer6_outputs[3939]);
    assign outputs[2399] = layer6_outputs[2984];
    assign outputs[2400] = layer6_outputs[5116];
    assign outputs[2401] = (layer6_outputs[3403]) & (layer6_outputs[4907]);
    assign outputs[2402] = ~(layer6_outputs[2289]);
    assign outputs[2403] = (layer6_outputs[2349]) & ~(layer6_outputs[4027]);
    assign outputs[2404] = layer6_outputs[3736];
    assign outputs[2405] = layer6_outputs[859];
    assign outputs[2406] = ~(layer6_outputs[4112]);
    assign outputs[2407] = (layer6_outputs[2707]) ^ (layer6_outputs[415]);
    assign outputs[2408] = ~(layer6_outputs[5087]);
    assign outputs[2409] = ~((layer6_outputs[1639]) ^ (layer6_outputs[296]));
    assign outputs[2410] = ~(layer6_outputs[4645]);
    assign outputs[2411] = ~((layer6_outputs[3802]) ^ (layer6_outputs[4705]));
    assign outputs[2412] = ~((layer6_outputs[2046]) ^ (layer6_outputs[1838]));
    assign outputs[2413] = ~(layer6_outputs[628]);
    assign outputs[2414] = (layer6_outputs[2137]) & ~(layer6_outputs[3986]);
    assign outputs[2415] = ~(layer6_outputs[314]);
    assign outputs[2416] = ~(layer6_outputs[2951]);
    assign outputs[2417] = ~((layer6_outputs[857]) ^ (layer6_outputs[2545]));
    assign outputs[2418] = ~(layer6_outputs[2267]);
    assign outputs[2419] = ~((layer6_outputs[1949]) ^ (layer6_outputs[2460]));
    assign outputs[2420] = ~(layer6_outputs[4599]);
    assign outputs[2421] = (layer6_outputs[4472]) ^ (layer6_outputs[3059]);
    assign outputs[2422] = ~(layer6_outputs[164]);
    assign outputs[2423] = (layer6_outputs[1708]) ^ (layer6_outputs[500]);
    assign outputs[2424] = layer6_outputs[4216];
    assign outputs[2425] = ~(layer6_outputs[841]);
    assign outputs[2426] = layer6_outputs[4941];
    assign outputs[2427] = ~(layer6_outputs[1504]);
    assign outputs[2428] = ~(layer6_outputs[2604]);
    assign outputs[2429] = (layer6_outputs[4584]) & (layer6_outputs[414]);
    assign outputs[2430] = (layer6_outputs[2219]) ^ (layer6_outputs[1928]);
    assign outputs[2431] = (layer6_outputs[906]) ^ (layer6_outputs[893]);
    assign outputs[2432] = ~(layer6_outputs[2860]);
    assign outputs[2433] = ~(layer6_outputs[1453]) | (layer6_outputs[1578]);
    assign outputs[2434] = ~(layer6_outputs[1765]);
    assign outputs[2435] = ~((layer6_outputs[2838]) ^ (layer6_outputs[725]));
    assign outputs[2436] = ~((layer6_outputs[3644]) ^ (layer6_outputs[4895]));
    assign outputs[2437] = ~(layer6_outputs[42]);
    assign outputs[2438] = layer6_outputs[3331];
    assign outputs[2439] = ~((layer6_outputs[3635]) ^ (layer6_outputs[796]));
    assign outputs[2440] = layer6_outputs[3464];
    assign outputs[2441] = ~(layer6_outputs[1808]);
    assign outputs[2442] = layer6_outputs[3820];
    assign outputs[2443] = layer6_outputs[4155];
    assign outputs[2444] = (layer6_outputs[2212]) ^ (layer6_outputs[3392]);
    assign outputs[2445] = layer6_outputs[1024];
    assign outputs[2446] = (layer6_outputs[2621]) ^ (layer6_outputs[1983]);
    assign outputs[2447] = (layer6_outputs[2181]) & (layer6_outputs[3141]);
    assign outputs[2448] = layer6_outputs[1494];
    assign outputs[2449] = layer6_outputs[5063];
    assign outputs[2450] = (layer6_outputs[2454]) | (layer6_outputs[2677]);
    assign outputs[2451] = ~(layer6_outputs[5109]);
    assign outputs[2452] = (layer6_outputs[1911]) & ~(layer6_outputs[4896]);
    assign outputs[2453] = (layer6_outputs[3256]) ^ (layer6_outputs[2531]);
    assign outputs[2454] = layer6_outputs[4678];
    assign outputs[2455] = (layer6_outputs[1861]) & (layer6_outputs[3311]);
    assign outputs[2456] = (layer6_outputs[4362]) & ~(layer6_outputs[4583]);
    assign outputs[2457] = ~(layer6_outputs[3383]);
    assign outputs[2458] = layer6_outputs[2186];
    assign outputs[2459] = ~(layer6_outputs[4193]);
    assign outputs[2460] = ~(layer6_outputs[2237]);
    assign outputs[2461] = (layer6_outputs[2585]) & ~(layer6_outputs[60]);
    assign outputs[2462] = ~(layer6_outputs[3226]);
    assign outputs[2463] = ~(layer6_outputs[380]);
    assign outputs[2464] = ~((layer6_outputs[547]) ^ (layer6_outputs[4794]));
    assign outputs[2465] = (layer6_outputs[4402]) & (layer6_outputs[521]);
    assign outputs[2466] = ~(layer6_outputs[3693]);
    assign outputs[2467] = (layer6_outputs[3749]) ^ (layer6_outputs[1590]);
    assign outputs[2468] = (layer6_outputs[3535]) & ~(layer6_outputs[840]);
    assign outputs[2469] = 1'b0;
    assign outputs[2470] = ~((layer6_outputs[911]) ^ (layer6_outputs[1397]));
    assign outputs[2471] = layer6_outputs[1187];
    assign outputs[2472] = (layer6_outputs[665]) ^ (layer6_outputs[3181]);
    assign outputs[2473] = ~((layer6_outputs[4464]) | (layer6_outputs[4519]));
    assign outputs[2474] = (layer6_outputs[2416]) & ~(layer6_outputs[4450]);
    assign outputs[2475] = layer6_outputs[2813];
    assign outputs[2476] = ~((layer6_outputs[5062]) | (layer6_outputs[138]));
    assign outputs[2477] = layer6_outputs[2142];
    assign outputs[2478] = (layer6_outputs[3889]) & ~(layer6_outputs[4173]);
    assign outputs[2479] = layer6_outputs[4537];
    assign outputs[2480] = (layer6_outputs[1447]) & ~(layer6_outputs[4089]);
    assign outputs[2481] = ~(layer6_outputs[1536]);
    assign outputs[2482] = layer6_outputs[2910];
    assign outputs[2483] = layer6_outputs[2510];
    assign outputs[2484] = layer6_outputs[4943];
    assign outputs[2485] = layer6_outputs[1648];
    assign outputs[2486] = ~((layer6_outputs[2675]) ^ (layer6_outputs[2727]));
    assign outputs[2487] = ~(layer6_outputs[4580]) | (layer6_outputs[5038]);
    assign outputs[2488] = layer6_outputs[1691];
    assign outputs[2489] = ~(layer6_outputs[4962]);
    assign outputs[2490] = layer6_outputs[923];
    assign outputs[2491] = (layer6_outputs[1520]) ^ (layer6_outputs[698]);
    assign outputs[2492] = (layer6_outputs[4099]) ^ (layer6_outputs[284]);
    assign outputs[2493] = ~(layer6_outputs[2148]);
    assign outputs[2494] = ~(layer6_outputs[3372]);
    assign outputs[2495] = (layer6_outputs[2040]) & ~(layer6_outputs[907]);
    assign outputs[2496] = layer6_outputs[5035];
    assign outputs[2497] = (layer6_outputs[1370]) & ~(layer6_outputs[964]);
    assign outputs[2498] = ~(layer6_outputs[4628]);
    assign outputs[2499] = ~((layer6_outputs[1545]) | (layer6_outputs[649]));
    assign outputs[2500] = layer6_outputs[2283];
    assign outputs[2501] = ~(layer6_outputs[95]);
    assign outputs[2502] = ~(layer6_outputs[4344]);
    assign outputs[2503] = ~((layer6_outputs[4295]) ^ (layer6_outputs[4717]));
    assign outputs[2504] = ~(layer6_outputs[4896]);
    assign outputs[2505] = layer6_outputs[4026];
    assign outputs[2506] = ~(layer6_outputs[4195]);
    assign outputs[2507] = layer6_outputs[193];
    assign outputs[2508] = layer6_outputs[2639];
    assign outputs[2509] = layer6_outputs[4684];
    assign outputs[2510] = layer6_outputs[3248];
    assign outputs[2511] = layer6_outputs[1814];
    assign outputs[2512] = ~(layer6_outputs[592]);
    assign outputs[2513] = layer6_outputs[3410];
    assign outputs[2514] = ~((layer6_outputs[1656]) | (layer6_outputs[2746]));
    assign outputs[2515] = (layer6_outputs[1865]) & ~(layer6_outputs[1604]);
    assign outputs[2516] = layer6_outputs[4611];
    assign outputs[2517] = ~(layer6_outputs[963]);
    assign outputs[2518] = ~(layer6_outputs[1082]);
    assign outputs[2519] = layer6_outputs[44];
    assign outputs[2520] = (layer6_outputs[146]) & ~(layer6_outputs[3591]);
    assign outputs[2521] = layer6_outputs[733];
    assign outputs[2522] = ~(layer6_outputs[4063]);
    assign outputs[2523] = (layer6_outputs[442]) & ~(layer6_outputs[1360]);
    assign outputs[2524] = layer6_outputs[1958];
    assign outputs[2525] = layer6_outputs[1684];
    assign outputs[2526] = (layer6_outputs[683]) ^ (layer6_outputs[4611]);
    assign outputs[2527] = ~((layer6_outputs[1697]) | (layer6_outputs[4679]));
    assign outputs[2528] = ~(layer6_outputs[3757]);
    assign outputs[2529] = ~((layer6_outputs[3908]) ^ (layer6_outputs[4114]));
    assign outputs[2530] = (layer6_outputs[2131]) & (layer6_outputs[1452]);
    assign outputs[2531] = layer6_outputs[1206];
    assign outputs[2532] = ~(layer6_outputs[1636]);
    assign outputs[2533] = ~(layer6_outputs[2734]);
    assign outputs[2534] = layer6_outputs[4692];
    assign outputs[2535] = ~(layer6_outputs[4636]);
    assign outputs[2536] = layer6_outputs[4200];
    assign outputs[2537] = ~(layer6_outputs[4012]);
    assign outputs[2538] = (layer6_outputs[3351]) ^ (layer6_outputs[3458]);
    assign outputs[2539] = ~(layer6_outputs[115]);
    assign outputs[2540] = (layer6_outputs[1315]) & ~(layer6_outputs[3528]);
    assign outputs[2541] = layer6_outputs[4411];
    assign outputs[2542] = (layer6_outputs[2696]) | (layer6_outputs[3846]);
    assign outputs[2543] = (layer6_outputs[819]) ^ (layer6_outputs[4362]);
    assign outputs[2544] = layer6_outputs[3648];
    assign outputs[2545] = layer6_outputs[3703];
    assign outputs[2546] = layer6_outputs[2058];
    assign outputs[2547] = (layer6_outputs[651]) ^ (layer6_outputs[2739]);
    assign outputs[2548] = ~(layer6_outputs[3298]);
    assign outputs[2549] = ~((layer6_outputs[3373]) | (layer6_outputs[3447]));
    assign outputs[2550] = ~(layer6_outputs[507]);
    assign outputs[2551] = (layer6_outputs[312]) ^ (layer6_outputs[4387]);
    assign outputs[2552] = (layer6_outputs[2214]) ^ (layer6_outputs[2485]);
    assign outputs[2553] = ~(layer6_outputs[308]);
    assign outputs[2554] = layer6_outputs[3691];
    assign outputs[2555] = ~(layer6_outputs[452]);
    assign outputs[2556] = layer6_outputs[2990];
    assign outputs[2557] = layer6_outputs[3187];
    assign outputs[2558] = ~(layer6_outputs[1417]);
    assign outputs[2559] = ~((layer6_outputs[1843]) ^ (layer6_outputs[366]));
    assign outputs[2560] = layer6_outputs[280];
    assign outputs[2561] = layer6_outputs[4469];
    assign outputs[2562] = layer6_outputs[2881];
    assign outputs[2563] = ~((layer6_outputs[3656]) ^ (layer6_outputs[2380]));
    assign outputs[2564] = (layer6_outputs[4529]) | (layer6_outputs[270]);
    assign outputs[2565] = layer6_outputs[3167];
    assign outputs[2566] = layer6_outputs[2316];
    assign outputs[2567] = ~(layer6_outputs[268]);
    assign outputs[2568] = (layer6_outputs[2516]) ^ (layer6_outputs[664]);
    assign outputs[2569] = ~(layer6_outputs[3440]);
    assign outputs[2570] = ~((layer6_outputs[4767]) & (layer6_outputs[4849]));
    assign outputs[2571] = ~(layer6_outputs[4230]);
    assign outputs[2572] = layer6_outputs[3951];
    assign outputs[2573] = ~(layer6_outputs[4448]);
    assign outputs[2574] = layer6_outputs[2309];
    assign outputs[2575] = ~(layer6_outputs[4812]);
    assign outputs[2576] = layer6_outputs[4675];
    assign outputs[2577] = ~(layer6_outputs[4400]);
    assign outputs[2578] = ~(layer6_outputs[144]) | (layer6_outputs[3154]);
    assign outputs[2579] = ~((layer6_outputs[843]) ^ (layer6_outputs[285]));
    assign outputs[2580] = (layer6_outputs[4024]) ^ (layer6_outputs[1027]);
    assign outputs[2581] = ~((layer6_outputs[672]) ^ (layer6_outputs[1770]));
    assign outputs[2582] = (layer6_outputs[4412]) & (layer6_outputs[1079]);
    assign outputs[2583] = layer6_outputs[1693];
    assign outputs[2584] = layer6_outputs[4360];
    assign outputs[2585] = layer6_outputs[4690];
    assign outputs[2586] = (layer6_outputs[1303]) ^ (layer6_outputs[3262]);
    assign outputs[2587] = layer6_outputs[4990];
    assign outputs[2588] = (layer6_outputs[3752]) ^ (layer6_outputs[3101]);
    assign outputs[2589] = ~(layer6_outputs[4203]);
    assign outputs[2590] = ~(layer6_outputs[1922]);
    assign outputs[2591] = layer6_outputs[3185];
    assign outputs[2592] = ~((layer6_outputs[3045]) & (layer6_outputs[4303]));
    assign outputs[2593] = ~(layer6_outputs[1937]) | (layer6_outputs[2412]);
    assign outputs[2594] = ~((layer6_outputs[589]) ^ (layer6_outputs[1791]));
    assign outputs[2595] = ~(layer6_outputs[2386]);
    assign outputs[2596] = layer6_outputs[478];
    assign outputs[2597] = layer6_outputs[1];
    assign outputs[2598] = (layer6_outputs[1924]) ^ (layer6_outputs[4681]);
    assign outputs[2599] = ~((layer6_outputs[4899]) ^ (layer6_outputs[2998]));
    assign outputs[2600] = layer6_outputs[4700];
    assign outputs[2601] = ~((layer6_outputs[1402]) ^ (layer6_outputs[3524]));
    assign outputs[2602] = (layer6_outputs[277]) ^ (layer6_outputs[1960]);
    assign outputs[2603] = layer6_outputs[2706];
    assign outputs[2604] = (layer6_outputs[4727]) & (layer6_outputs[909]);
    assign outputs[2605] = (layer6_outputs[1129]) ^ (layer6_outputs[3112]);
    assign outputs[2606] = ~((layer6_outputs[3829]) ^ (layer6_outputs[2488]));
    assign outputs[2607] = ~((layer6_outputs[4223]) ^ (layer6_outputs[3566]));
    assign outputs[2608] = (layer6_outputs[2688]) ^ (layer6_outputs[450]);
    assign outputs[2609] = (layer6_outputs[1490]) ^ (layer6_outputs[4724]);
    assign outputs[2610] = ~(layer6_outputs[3858]) | (layer6_outputs[903]);
    assign outputs[2611] = ~((layer6_outputs[4694]) ^ (layer6_outputs[108]));
    assign outputs[2612] = (layer6_outputs[4057]) & ~(layer6_outputs[3927]);
    assign outputs[2613] = ~(layer6_outputs[301]);
    assign outputs[2614] = ~(layer6_outputs[2611]);
    assign outputs[2615] = ~(layer6_outputs[3100]);
    assign outputs[2616] = layer6_outputs[2645];
    assign outputs[2617] = (layer6_outputs[1948]) | (layer6_outputs[435]);
    assign outputs[2618] = (layer6_outputs[4300]) ^ (layer6_outputs[4575]);
    assign outputs[2619] = (layer6_outputs[4900]) ^ (layer6_outputs[2489]);
    assign outputs[2620] = (layer6_outputs[404]) ^ (layer6_outputs[4483]);
    assign outputs[2621] = ~((layer6_outputs[2374]) ^ (layer6_outputs[3670]));
    assign outputs[2622] = layer6_outputs[808];
    assign outputs[2623] = ~(layer6_outputs[3846]);
    assign outputs[2624] = ~(layer6_outputs[1704]);
    assign outputs[2625] = (layer6_outputs[2048]) ^ (layer6_outputs[2788]);
    assign outputs[2626] = ~((layer6_outputs[997]) ^ (layer6_outputs[887]));
    assign outputs[2627] = layer6_outputs[3224];
    assign outputs[2628] = ~((layer6_outputs[288]) & (layer6_outputs[212]));
    assign outputs[2629] = layer6_outputs[3877];
    assign outputs[2630] = (layer6_outputs[632]) ^ (layer6_outputs[4607]);
    assign outputs[2631] = ~((layer6_outputs[1931]) ^ (layer6_outputs[1639]));
    assign outputs[2632] = (layer6_outputs[848]) ^ (layer6_outputs[4222]);
    assign outputs[2633] = layer6_outputs[4359];
    assign outputs[2634] = layer6_outputs[2652];
    assign outputs[2635] = ~((layer6_outputs[1053]) ^ (layer6_outputs[657]));
    assign outputs[2636] = ~(layer6_outputs[2150]);
    assign outputs[2637] = ~(layer6_outputs[4506]);
    assign outputs[2638] = ~(layer6_outputs[1102]);
    assign outputs[2639] = (layer6_outputs[2233]) ^ (layer6_outputs[600]);
    assign outputs[2640] = layer6_outputs[359];
    assign outputs[2641] = (layer6_outputs[2193]) ^ (layer6_outputs[1723]);
    assign outputs[2642] = ~(layer6_outputs[2155]);
    assign outputs[2643] = (layer6_outputs[1318]) ^ (layer6_outputs[3506]);
    assign outputs[2644] = ~((layer6_outputs[1448]) ^ (layer6_outputs[4229]));
    assign outputs[2645] = ~(layer6_outputs[1617]) | (layer6_outputs[4994]);
    assign outputs[2646] = ~(layer6_outputs[2877]);
    assign outputs[2647] = ~(layer6_outputs[4457]);
    assign outputs[2648] = ~(layer6_outputs[3320]) | (layer6_outputs[637]);
    assign outputs[2649] = ~((layer6_outputs[208]) | (layer6_outputs[381]));
    assign outputs[2650] = ~(layer6_outputs[1668]);
    assign outputs[2651] = (layer6_outputs[1932]) & (layer6_outputs[1316]);
    assign outputs[2652] = ~((layer6_outputs[1129]) ^ (layer6_outputs[4281]));
    assign outputs[2653] = ~(layer6_outputs[69]);
    assign outputs[2654] = layer6_outputs[3345];
    assign outputs[2655] = ~(layer6_outputs[3512]);
    assign outputs[2656] = (layer6_outputs[3984]) ^ (layer6_outputs[2224]);
    assign outputs[2657] = layer6_outputs[217];
    assign outputs[2658] = ~(layer6_outputs[2099]);
    assign outputs[2659] = ~((layer6_outputs[2747]) ^ (layer6_outputs[3276]));
    assign outputs[2660] = ~(layer6_outputs[2164]);
    assign outputs[2661] = layer6_outputs[3301];
    assign outputs[2662] = (layer6_outputs[2748]) ^ (layer6_outputs[4598]);
    assign outputs[2663] = (layer6_outputs[1706]) ^ (layer6_outputs[4985]);
    assign outputs[2664] = layer6_outputs[3048];
    assign outputs[2665] = (layer6_outputs[4039]) & ~(layer6_outputs[1991]);
    assign outputs[2666] = layer6_outputs[4239];
    assign outputs[2667] = ~(layer6_outputs[3959]);
    assign outputs[2668] = layer6_outputs[715];
    assign outputs[2669] = layer6_outputs[19];
    assign outputs[2670] = (layer6_outputs[1022]) ^ (layer6_outputs[4110]);
    assign outputs[2671] = (layer6_outputs[1558]) ^ (layer6_outputs[1587]);
    assign outputs[2672] = (layer6_outputs[1796]) ^ (layer6_outputs[3099]);
    assign outputs[2673] = ~(layer6_outputs[5045]);
    assign outputs[2674] = ~(layer6_outputs[5071]);
    assign outputs[2675] = (layer6_outputs[2413]) & (layer6_outputs[342]);
    assign outputs[2676] = ~(layer6_outputs[1277]);
    assign outputs[2677] = ~(layer6_outputs[3280]);
    assign outputs[2678] = ~(layer6_outputs[2829]);
    assign outputs[2679] = ~((layer6_outputs[941]) ^ (layer6_outputs[2999]));
    assign outputs[2680] = layer6_outputs[1814];
    assign outputs[2681] = ~(layer6_outputs[4862]);
    assign outputs[2682] = ~(layer6_outputs[5098]);
    assign outputs[2683] = ~((layer6_outputs[948]) | (layer6_outputs[3098]));
    assign outputs[2684] = layer6_outputs[2191];
    assign outputs[2685] = layer6_outputs[3831];
    assign outputs[2686] = ~(layer6_outputs[1369]);
    assign outputs[2687] = ~(layer6_outputs[3824]);
    assign outputs[2688] = ~(layer6_outputs[687]);
    assign outputs[2689] = ~((layer6_outputs[3500]) ^ (layer6_outputs[416]));
    assign outputs[2690] = ~(layer6_outputs[3308]);
    assign outputs[2691] = layer6_outputs[4975];
    assign outputs[2692] = ~(layer6_outputs[2358]);
    assign outputs[2693] = ~(layer6_outputs[1203]);
    assign outputs[2694] = (layer6_outputs[107]) ^ (layer6_outputs[986]);
    assign outputs[2695] = ~(layer6_outputs[4016]);
    assign outputs[2696] = layer6_outputs[2014];
    assign outputs[2697] = layer6_outputs[2508];
    assign outputs[2698] = ~((layer6_outputs[884]) ^ (layer6_outputs[5054]));
    assign outputs[2699] = ~(layer6_outputs[4921]);
    assign outputs[2700] = ~(layer6_outputs[1899]);
    assign outputs[2701] = ~((layer6_outputs[2083]) & (layer6_outputs[3206]));
    assign outputs[2702] = ~((layer6_outputs[142]) ^ (layer6_outputs[3189]));
    assign outputs[2703] = layer6_outputs[2332];
    assign outputs[2704] = layer6_outputs[2409];
    assign outputs[2705] = ~((layer6_outputs[2483]) ^ (layer6_outputs[4733]));
    assign outputs[2706] = layer6_outputs[4827];
    assign outputs[2707] = (layer6_outputs[1260]) ^ (layer6_outputs[2206]);
    assign outputs[2708] = (layer6_outputs[1728]) ^ (layer6_outputs[661]);
    assign outputs[2709] = ~(layer6_outputs[3530]);
    assign outputs[2710] = (layer6_outputs[4238]) ^ (layer6_outputs[2596]);
    assign outputs[2711] = layer6_outputs[2447];
    assign outputs[2712] = (layer6_outputs[4911]) ^ (layer6_outputs[583]);
    assign outputs[2713] = layer6_outputs[4841];
    assign outputs[2714] = layer6_outputs[2710];
    assign outputs[2715] = ~(layer6_outputs[1462]);
    assign outputs[2716] = ~(layer6_outputs[336]);
    assign outputs[2717] = layer6_outputs[3109];
    assign outputs[2718] = (layer6_outputs[834]) ^ (layer6_outputs[4021]);
    assign outputs[2719] = (layer6_outputs[1058]) ^ (layer6_outputs[2949]);
    assign outputs[2720] = (layer6_outputs[4702]) ^ (layer6_outputs[287]);
    assign outputs[2721] = layer6_outputs[273];
    assign outputs[2722] = (layer6_outputs[4873]) ^ (layer6_outputs[2499]);
    assign outputs[2723] = ~((layer6_outputs[727]) ^ (layer6_outputs[4905]));
    assign outputs[2724] = (layer6_outputs[2060]) ^ (layer6_outputs[151]);
    assign outputs[2725] = ~(layer6_outputs[494]);
    assign outputs[2726] = ~((layer6_outputs[4895]) & (layer6_outputs[4337]));
    assign outputs[2727] = ~(layer6_outputs[4670]);
    assign outputs[2728] = ~((layer6_outputs[3884]) ^ (layer6_outputs[456]));
    assign outputs[2729] = layer6_outputs[1747];
    assign outputs[2730] = ~((layer6_outputs[277]) ^ (layer6_outputs[2362]));
    assign outputs[2731] = layer6_outputs[3745];
    assign outputs[2732] = ~(layer6_outputs[3952]);
    assign outputs[2733] = ~(layer6_outputs[2389]);
    assign outputs[2734] = ~(layer6_outputs[3713]);
    assign outputs[2735] = (layer6_outputs[4857]) ^ (layer6_outputs[20]);
    assign outputs[2736] = ~(layer6_outputs[3485]);
    assign outputs[2737] = layer6_outputs[4940];
    assign outputs[2738] = layer6_outputs[4922];
    assign outputs[2739] = ~((layer6_outputs[3035]) ^ (layer6_outputs[3821]));
    assign outputs[2740] = ~(layer6_outputs[3353]);
    assign outputs[2741] = layer6_outputs[1101];
    assign outputs[2742] = ~(layer6_outputs[2595]);
    assign outputs[2743] = ~(layer6_outputs[4190]);
    assign outputs[2744] = (layer6_outputs[3909]) ^ (layer6_outputs[4428]);
    assign outputs[2745] = (layer6_outputs[881]) & (layer6_outputs[1246]);
    assign outputs[2746] = layer6_outputs[923];
    assign outputs[2747] = layer6_outputs[1002];
    assign outputs[2748] = layer6_outputs[5058];
    assign outputs[2749] = ~(layer6_outputs[2547]);
    assign outputs[2750] = layer6_outputs[2276];
    assign outputs[2751] = (layer6_outputs[2896]) ^ (layer6_outputs[4127]);
    assign outputs[2752] = layer6_outputs[3037];
    assign outputs[2753] = layer6_outputs[4533];
    assign outputs[2754] = layer6_outputs[4554];
    assign outputs[2755] = ~((layer6_outputs[4407]) ^ (layer6_outputs[183]));
    assign outputs[2756] = ~(layer6_outputs[2547]);
    assign outputs[2757] = (layer6_outputs[348]) ^ (layer6_outputs[2503]);
    assign outputs[2758] = (layer6_outputs[3786]) & ~(layer6_outputs[746]);
    assign outputs[2759] = ~(layer6_outputs[4507]) | (layer6_outputs[3115]);
    assign outputs[2760] = ~(layer6_outputs[3402]);
    assign outputs[2761] = layer6_outputs[4568];
    assign outputs[2762] = ~((layer6_outputs[5007]) ^ (layer6_outputs[1571]));
    assign outputs[2763] = ~(layer6_outputs[1350]);
    assign outputs[2764] = ~(layer6_outputs[2325]);
    assign outputs[2765] = ~(layer6_outputs[3441]) | (layer6_outputs[2344]);
    assign outputs[2766] = ~((layer6_outputs[2018]) & (layer6_outputs[5018]));
    assign outputs[2767] = ~((layer6_outputs[830]) ^ (layer6_outputs[3714]));
    assign outputs[2768] = layer6_outputs[2790];
    assign outputs[2769] = (layer6_outputs[1378]) ^ (layer6_outputs[1881]);
    assign outputs[2770] = layer6_outputs[4743];
    assign outputs[2771] = ~(layer6_outputs[471]);
    assign outputs[2772] = ~(layer6_outputs[610]);
    assign outputs[2773] = layer6_outputs[1164];
    assign outputs[2774] = layer6_outputs[2658];
    assign outputs[2775] = ~((layer6_outputs[1089]) ^ (layer6_outputs[2598]));
    assign outputs[2776] = ~(layer6_outputs[2386]);
    assign outputs[2777] = layer6_outputs[3940];
    assign outputs[2778] = ~(layer6_outputs[2808]);
    assign outputs[2779] = ~(layer6_outputs[3995]);
    assign outputs[2780] = ~(layer6_outputs[331]) | (layer6_outputs[1935]);
    assign outputs[2781] = ~((layer6_outputs[4213]) & (layer6_outputs[3359]));
    assign outputs[2782] = ~(layer6_outputs[1625]);
    assign outputs[2783] = layer6_outputs[432];
    assign outputs[2784] = ~(layer6_outputs[3737]);
    assign outputs[2785] = ~((layer6_outputs[3986]) ^ (layer6_outputs[557]));
    assign outputs[2786] = ~((layer6_outputs[2079]) ^ (layer6_outputs[4370]));
    assign outputs[2787] = ~(layer6_outputs[3771]);
    assign outputs[2788] = layer6_outputs[3564];
    assign outputs[2789] = layer6_outputs[4210];
    assign outputs[2790] = ~((layer6_outputs[2714]) ^ (layer6_outputs[1603]));
    assign outputs[2791] = layer6_outputs[1522];
    assign outputs[2792] = ~((layer6_outputs[860]) ^ (layer6_outputs[3020]));
    assign outputs[2793] = ~(layer6_outputs[3836]);
    assign outputs[2794] = ~(layer6_outputs[2559]);
    assign outputs[2795] = (layer6_outputs[3183]) ^ (layer6_outputs[3702]);
    assign outputs[2796] = layer6_outputs[2015];
    assign outputs[2797] = ~(layer6_outputs[5066]);
    assign outputs[2798] = ~(layer6_outputs[5012]);
    assign outputs[2799] = layer6_outputs[4441];
    assign outputs[2800] = ~((layer6_outputs[4645]) ^ (layer6_outputs[1607]));
    assign outputs[2801] = layer6_outputs[1235];
    assign outputs[2802] = layer6_outputs[4910];
    assign outputs[2803] = layer6_outputs[3717];
    assign outputs[2804] = (layer6_outputs[4809]) & ~(layer6_outputs[3087]);
    assign outputs[2805] = (layer6_outputs[13]) & ~(layer6_outputs[1269]);
    assign outputs[2806] = ~(layer6_outputs[3742]);
    assign outputs[2807] = layer6_outputs[5101];
    assign outputs[2808] = layer6_outputs[705];
    assign outputs[2809] = layer6_outputs[603];
    assign outputs[2810] = layer6_outputs[2117];
    assign outputs[2811] = ~(layer6_outputs[485]);
    assign outputs[2812] = ~(layer6_outputs[605]) | (layer6_outputs[4916]);
    assign outputs[2813] = ~(layer6_outputs[1531]);
    assign outputs[2814] = ~(layer6_outputs[4010]);
    assign outputs[2815] = layer6_outputs[3106];
    assign outputs[2816] = ~((layer6_outputs[3714]) ^ (layer6_outputs[56]));
    assign outputs[2817] = layer6_outputs[1072];
    assign outputs[2818] = ~(layer6_outputs[389]);
    assign outputs[2819] = ~(layer6_outputs[4080]);
    assign outputs[2820] = layer6_outputs[2697];
    assign outputs[2821] = ~((layer6_outputs[1670]) ^ (layer6_outputs[3504]));
    assign outputs[2822] = ~((layer6_outputs[2222]) ^ (layer6_outputs[146]));
    assign outputs[2823] = layer6_outputs[1378];
    assign outputs[2824] = ~(layer6_outputs[2525]) | (layer6_outputs[2010]);
    assign outputs[2825] = layer6_outputs[1554];
    assign outputs[2826] = ~(layer6_outputs[1485]);
    assign outputs[2827] = layer6_outputs[2268];
    assign outputs[2828] = layer6_outputs[651];
    assign outputs[2829] = (layer6_outputs[1654]) ^ (layer6_outputs[1471]);
    assign outputs[2830] = layer6_outputs[4017];
    assign outputs[2831] = ~(layer6_outputs[1236]);
    assign outputs[2832] = ~((layer6_outputs[4870]) ^ (layer6_outputs[4116]));
    assign outputs[2833] = (layer6_outputs[2912]) ^ (layer6_outputs[1748]);
    assign outputs[2834] = (layer6_outputs[2751]) & (layer6_outputs[4255]);
    assign outputs[2835] = (layer6_outputs[4198]) & ~(layer6_outputs[3675]);
    assign outputs[2836] = (layer6_outputs[1066]) ^ (layer6_outputs[3280]);
    assign outputs[2837] = ~((layer6_outputs[2950]) ^ (layer6_outputs[2314]));
    assign outputs[2838] = layer6_outputs[2601];
    assign outputs[2839] = layer6_outputs[4708];
    assign outputs[2840] = ~(layer6_outputs[1458]) | (layer6_outputs[3666]);
    assign outputs[2841] = ~(layer6_outputs[1229]);
    assign outputs[2842] = layer6_outputs[3679];
    assign outputs[2843] = ~((layer6_outputs[16]) ^ (layer6_outputs[4569]));
    assign outputs[2844] = ~(layer6_outputs[4479]);
    assign outputs[2845] = (layer6_outputs[2158]) ^ (layer6_outputs[3948]);
    assign outputs[2846] = layer6_outputs[3985];
    assign outputs[2847] = ~((layer6_outputs[4342]) ^ (layer6_outputs[4025]));
    assign outputs[2848] = (layer6_outputs[1692]) & (layer6_outputs[267]);
    assign outputs[2849] = ~(layer6_outputs[2089]);
    assign outputs[2850] = layer6_outputs[4815];
    assign outputs[2851] = layer6_outputs[2822];
    assign outputs[2852] = (layer6_outputs[4339]) | (layer6_outputs[1967]);
    assign outputs[2853] = layer6_outputs[1247];
    assign outputs[2854] = ~(layer6_outputs[4545]);
    assign outputs[2855] = ~(layer6_outputs[3315]);
    assign outputs[2856] = layer6_outputs[858];
    assign outputs[2857] = ~(layer6_outputs[4881]);
    assign outputs[2858] = (layer6_outputs[750]) ^ (layer6_outputs[1840]);
    assign outputs[2859] = (layer6_outputs[3734]) & (layer6_outputs[830]);
    assign outputs[2860] = ~(layer6_outputs[1566]);
    assign outputs[2861] = layer6_outputs[2550];
    assign outputs[2862] = (layer6_outputs[1059]) | (layer6_outputs[2969]);
    assign outputs[2863] = ~((layer6_outputs[4426]) ^ (layer6_outputs[62]));
    assign outputs[2864] = ~((layer6_outputs[10]) ^ (layer6_outputs[3661]));
    assign outputs[2865] = layer6_outputs[3823];
    assign outputs[2866] = ~((layer6_outputs[4612]) ^ (layer6_outputs[3430]));
    assign outputs[2867] = layer6_outputs[1450];
    assign outputs[2868] = ~(layer6_outputs[4848]) | (layer6_outputs[2837]);
    assign outputs[2869] = layer6_outputs[1985];
    assign outputs[2870] = (layer6_outputs[1665]) ^ (layer6_outputs[2452]);
    assign outputs[2871] = ~(layer6_outputs[2541]);
    assign outputs[2872] = layer6_outputs[3381];
    assign outputs[2873] = ~(layer6_outputs[10]) | (layer6_outputs[2406]);
    assign outputs[2874] = ~((layer6_outputs[470]) ^ (layer6_outputs[1993]));
    assign outputs[2875] = ~(layer6_outputs[2802]);
    assign outputs[2876] = layer6_outputs[927];
    assign outputs[2877] = ~(layer6_outputs[2190]) | (layer6_outputs[1686]);
    assign outputs[2878] = ~(layer6_outputs[2836]);
    assign outputs[2879] = ~((layer6_outputs[1109]) ^ (layer6_outputs[1301]));
    assign outputs[2880] = (layer6_outputs[2504]) & ~(layer6_outputs[2818]);
    assign outputs[2881] = ~(layer6_outputs[4616]);
    assign outputs[2882] = ~(layer6_outputs[4098]);
    assign outputs[2883] = (layer6_outputs[4704]) & ~(layer6_outputs[2024]);
    assign outputs[2884] = layer6_outputs[3106];
    assign outputs[2885] = ~(layer6_outputs[5061]);
    assign outputs[2886] = ~(layer6_outputs[4411]);
    assign outputs[2887] = ~((layer6_outputs[3415]) ^ (layer6_outputs[1392]));
    assign outputs[2888] = ~((layer6_outputs[2094]) ^ (layer6_outputs[902]));
    assign outputs[2889] = layer6_outputs[1907];
    assign outputs[2890] = ~((layer6_outputs[3907]) ^ (layer6_outputs[4433]));
    assign outputs[2891] = ~(layer6_outputs[4375]);
    assign outputs[2892] = ~(layer6_outputs[4444]);
    assign outputs[2893] = layer6_outputs[4228];
    assign outputs[2894] = (layer6_outputs[4861]) ^ (layer6_outputs[4646]);
    assign outputs[2895] = layer6_outputs[1907];
    assign outputs[2896] = layer6_outputs[3574];
    assign outputs[2897] = ~(layer6_outputs[2517]);
    assign outputs[2898] = (layer6_outputs[3919]) ^ (layer6_outputs[2614]);
    assign outputs[2899] = ~(layer6_outputs[800]);
    assign outputs[2900] = ~((layer6_outputs[437]) ^ (layer6_outputs[2622]));
    assign outputs[2901] = (layer6_outputs[92]) ^ (layer6_outputs[4199]);
    assign outputs[2902] = ~(layer6_outputs[522]);
    assign outputs[2903] = (layer6_outputs[718]) ^ (layer6_outputs[1103]);
    assign outputs[2904] = layer6_outputs[3411];
    assign outputs[2905] = ~((layer6_outputs[5104]) ^ (layer6_outputs[3926]));
    assign outputs[2906] = (layer6_outputs[3368]) ^ (layer6_outputs[1171]);
    assign outputs[2907] = ~((layer6_outputs[1488]) ^ (layer6_outputs[480]));
    assign outputs[2908] = ~((layer6_outputs[4201]) ^ (layer6_outputs[1416]));
    assign outputs[2909] = (layer6_outputs[175]) ^ (layer6_outputs[4914]);
    assign outputs[2910] = layer6_outputs[3245];
    assign outputs[2911] = ~(layer6_outputs[2990]);
    assign outputs[2912] = ~((layer6_outputs[2494]) ^ (layer6_outputs[1482]));
    assign outputs[2913] = (layer6_outputs[229]) ^ (layer6_outputs[544]);
    assign outputs[2914] = ~(layer6_outputs[3588]);
    assign outputs[2915] = ~(layer6_outputs[3271]);
    assign outputs[2916] = ~(layer6_outputs[4233]) | (layer6_outputs[1371]);
    assign outputs[2917] = layer6_outputs[1318];
    assign outputs[2918] = layer6_outputs[3942];
    assign outputs[2919] = ~((layer6_outputs[4840]) ^ (layer6_outputs[4043]));
    assign outputs[2920] = layer6_outputs[2495];
    assign outputs[2921] = ~(layer6_outputs[1196]);
    assign outputs[2922] = ~(layer6_outputs[2664]);
    assign outputs[2923] = layer6_outputs[3465];
    assign outputs[2924] = (layer6_outputs[1231]) | (layer6_outputs[4256]);
    assign outputs[2925] = ~(layer6_outputs[4440]);
    assign outputs[2926] = ~(layer6_outputs[4806]);
    assign outputs[2927] = ~(layer6_outputs[890]);
    assign outputs[2928] = ~(layer6_outputs[1292]);
    assign outputs[2929] = (layer6_outputs[4832]) ^ (layer6_outputs[4778]);
    assign outputs[2930] = ~(layer6_outputs[3924]);
    assign outputs[2931] = layer6_outputs[2729];
    assign outputs[2932] = ~((layer6_outputs[4268]) & (layer6_outputs[1084]));
    assign outputs[2933] = ~(layer6_outputs[1132]);
    assign outputs[2934] = (layer6_outputs[3695]) | (layer6_outputs[548]);
    assign outputs[2935] = (layer6_outputs[2282]) ^ (layer6_outputs[4865]);
    assign outputs[2936] = ~(layer6_outputs[3401]);
    assign outputs[2937] = ~(layer6_outputs[3656]);
    assign outputs[2938] = ~((layer6_outputs[4958]) ^ (layer6_outputs[4044]));
    assign outputs[2939] = (layer6_outputs[493]) ^ (layer6_outputs[1244]);
    assign outputs[2940] = ~(layer6_outputs[4437]);
    assign outputs[2941] = ~(layer6_outputs[1957]);
    assign outputs[2942] = ~(layer6_outputs[4]);
    assign outputs[2943] = ~((layer6_outputs[3466]) & (layer6_outputs[70]));
    assign outputs[2944] = ~(layer6_outputs[4329]);
    assign outputs[2945] = ~(layer6_outputs[356]);
    assign outputs[2946] = (layer6_outputs[5015]) ^ (layer6_outputs[614]);
    assign outputs[2947] = layer6_outputs[1802];
    assign outputs[2948] = ~(layer6_outputs[1191]);
    assign outputs[2949] = ~((layer6_outputs[3630]) ^ (layer6_outputs[1435]));
    assign outputs[2950] = ~(layer6_outputs[2824]);
    assign outputs[2951] = ~(layer6_outputs[2539]);
    assign outputs[2952] = layer6_outputs[2393];
    assign outputs[2953] = layer6_outputs[4717];
    assign outputs[2954] = ~((layer6_outputs[1584]) ^ (layer6_outputs[4468]));
    assign outputs[2955] = ~(layer6_outputs[2715]);
    assign outputs[2956] = (layer6_outputs[2466]) ^ (layer6_outputs[4103]);
    assign outputs[2957] = ~(layer6_outputs[1851]);
    assign outputs[2958] = layer6_outputs[935];
    assign outputs[2959] = layer6_outputs[4235];
    assign outputs[2960] = ~((layer6_outputs[4429]) ^ (layer6_outputs[3785]));
    assign outputs[2961] = ~(layer6_outputs[3064]);
    assign outputs[2962] = layer6_outputs[290];
    assign outputs[2963] = ~(layer6_outputs[3052]);
    assign outputs[2964] = layer6_outputs[4315];
    assign outputs[2965] = (layer6_outputs[2000]) & ~(layer6_outputs[3701]);
    assign outputs[2966] = layer6_outputs[2528];
    assign outputs[2967] = (layer6_outputs[751]) ^ (layer6_outputs[3105]);
    assign outputs[2968] = (layer6_outputs[4175]) & ~(layer6_outputs[1004]);
    assign outputs[2969] = ~(layer6_outputs[4318]);
    assign outputs[2970] = layer6_outputs[4819];
    assign outputs[2971] = ~(layer6_outputs[3126]);
    assign outputs[2972] = ~(layer6_outputs[1179]);
    assign outputs[2973] = ~(layer6_outputs[459]);
    assign outputs[2974] = layer6_outputs[835];
    assign outputs[2975] = ~(layer6_outputs[4857]) | (layer6_outputs[3306]);
    assign outputs[2976] = ~(layer6_outputs[4266]);
    assign outputs[2977] = ~(layer6_outputs[648]);
    assign outputs[2978] = (layer6_outputs[3657]) & ~(layer6_outputs[2733]);
    assign outputs[2979] = layer6_outputs[2304];
    assign outputs[2980] = layer6_outputs[3092];
    assign outputs[2981] = (layer6_outputs[1964]) | (layer6_outputs[4892]);
    assign outputs[2982] = layer6_outputs[787];
    assign outputs[2983] = ~((layer6_outputs[1210]) ^ (layer6_outputs[2830]));
    assign outputs[2984] = ~(layer6_outputs[3682]);
    assign outputs[2985] = ~((layer6_outputs[3406]) ^ (layer6_outputs[322]));
    assign outputs[2986] = ~(layer6_outputs[4490]);
    assign outputs[2987] = ~((layer6_outputs[4967]) ^ (layer6_outputs[2272]));
    assign outputs[2988] = (layer6_outputs[1855]) & ~(layer6_outputs[5036]);
    assign outputs[2989] = (layer6_outputs[444]) | (layer6_outputs[4357]);
    assign outputs[2990] = ~((layer6_outputs[922]) ^ (layer6_outputs[3316]));
    assign outputs[2991] = layer6_outputs[647];
    assign outputs[2992] = layer6_outputs[4567];
    assign outputs[2993] = ~(layer6_outputs[4744]);
    assign outputs[2994] = ~(layer6_outputs[3508]);
    assign outputs[2995] = (layer6_outputs[2832]) ^ (layer6_outputs[1085]);
    assign outputs[2996] = ~(layer6_outputs[1547]);
    assign outputs[2997] = ~(layer6_outputs[902]);
    assign outputs[2998] = layer6_outputs[992];
    assign outputs[2999] = (layer6_outputs[3916]) ^ (layer6_outputs[4798]);
    assign outputs[3000] = ~(layer6_outputs[4764]);
    assign outputs[3001] = (layer6_outputs[4125]) ^ (layer6_outputs[2071]);
    assign outputs[3002] = ~((layer6_outputs[3606]) ^ (layer6_outputs[850]));
    assign outputs[3003] = ~(layer6_outputs[403]) | (layer6_outputs[3553]);
    assign outputs[3004] = ~((layer6_outputs[2533]) ^ (layer6_outputs[4487]));
    assign outputs[3005] = ~(layer6_outputs[1130]);
    assign outputs[3006] = ~(layer6_outputs[1632]);
    assign outputs[3007] = ~(layer6_outputs[2925]);
    assign outputs[3008] = ~(layer6_outputs[914]);
    assign outputs[3009] = layer6_outputs[4569];
    assign outputs[3010] = layer6_outputs[1398];
    assign outputs[3011] = layer6_outputs[4674];
    assign outputs[3012] = (layer6_outputs[2396]) & (layer6_outputs[4445]);
    assign outputs[3013] = ~(layer6_outputs[2043]) | (layer6_outputs[2590]);
    assign outputs[3014] = (layer6_outputs[4776]) ^ (layer6_outputs[3590]);
    assign outputs[3015] = layer6_outputs[191];
    assign outputs[3016] = (layer6_outputs[3599]) ^ (layer6_outputs[1060]);
    assign outputs[3017] = ~(layer6_outputs[382]);
    assign outputs[3018] = ~(layer6_outputs[3974]);
    assign outputs[3019] = ~(layer6_outputs[2313]);
    assign outputs[3020] = ~(layer6_outputs[4782]);
    assign outputs[3021] = ~(layer6_outputs[387]);
    assign outputs[3022] = (layer6_outputs[1779]) ^ (layer6_outputs[3548]);
    assign outputs[3023] = layer6_outputs[523];
    assign outputs[3024] = ~((layer6_outputs[1395]) ^ (layer6_outputs[2163]));
    assign outputs[3025] = ~(layer6_outputs[793]);
    assign outputs[3026] = layer6_outputs[1336];
    assign outputs[3027] = (layer6_outputs[4254]) & (layer6_outputs[231]);
    assign outputs[3028] = ~((layer6_outputs[58]) ^ (layer6_outputs[2461]));
    assign outputs[3029] = ~(layer6_outputs[3641]);
    assign outputs[3030] = (layer6_outputs[2188]) ^ (layer6_outputs[2139]);
    assign outputs[3031] = layer6_outputs[98];
    assign outputs[3032] = ~((layer6_outputs[983]) ^ (layer6_outputs[4072]));
    assign outputs[3033] = ~((layer6_outputs[702]) ^ (layer6_outputs[3416]));
    assign outputs[3034] = ~(layer6_outputs[1621]);
    assign outputs[3035] = ~((layer6_outputs[3363]) ^ (layer6_outputs[4691]));
    assign outputs[3036] = (layer6_outputs[4456]) ^ (layer6_outputs[351]);
    assign outputs[3037] = layer6_outputs[3124];
    assign outputs[3038] = layer6_outputs[4975];
    assign outputs[3039] = ~((layer6_outputs[2996]) ^ (layer6_outputs[2021]));
    assign outputs[3040] = ~(layer6_outputs[282]);
    assign outputs[3041] = ~((layer6_outputs[484]) ^ (layer6_outputs[2667]));
    assign outputs[3042] = (layer6_outputs[2244]) & ~(layer6_outputs[3367]);
    assign outputs[3043] = (layer6_outputs[1980]) & ~(layer6_outputs[2372]);
    assign outputs[3044] = ~(layer6_outputs[4267]) | (layer6_outputs[4563]);
    assign outputs[3045] = (layer6_outputs[396]) ^ (layer6_outputs[2491]);
    assign outputs[3046] = layer6_outputs[4836];
    assign outputs[3047] = layer6_outputs[2890];
    assign outputs[3048] = layer6_outputs[4100];
    assign outputs[3049] = ~((layer6_outputs[767]) ^ (layer6_outputs[2348]));
    assign outputs[3050] = ~(layer6_outputs[1531]);
    assign outputs[3051] = ~((layer6_outputs[3324]) & (layer6_outputs[3427]));
    assign outputs[3052] = ~(layer6_outputs[2640]) | (layer6_outputs[4119]);
    assign outputs[3053] = ~((layer6_outputs[5062]) ^ (layer6_outputs[526]));
    assign outputs[3054] = layer6_outputs[747];
    assign outputs[3055] = ~(layer6_outputs[1095]);
    assign outputs[3056] = ~(layer6_outputs[1610]);
    assign outputs[3057] = ~((layer6_outputs[3169]) ^ (layer6_outputs[2501]));
    assign outputs[3058] = ~(layer6_outputs[3485]);
    assign outputs[3059] = layer6_outputs[325];
    assign outputs[3060] = ~((layer6_outputs[5106]) ^ (layer6_outputs[1226]));
    assign outputs[3061] = ~(layer6_outputs[3809]);
    assign outputs[3062] = (layer6_outputs[1393]) ^ (layer6_outputs[559]);
    assign outputs[3063] = ~(layer6_outputs[59]) | (layer6_outputs[2221]);
    assign outputs[3064] = ~(layer6_outputs[2029]);
    assign outputs[3065] = layer6_outputs[4048];
    assign outputs[3066] = ~((layer6_outputs[304]) ^ (layer6_outputs[1853]));
    assign outputs[3067] = ~(layer6_outputs[3278]);
    assign outputs[3068] = ~((layer6_outputs[259]) ^ (layer6_outputs[3445]));
    assign outputs[3069] = ~(layer6_outputs[2552]);
    assign outputs[3070] = ~((layer6_outputs[3940]) ^ (layer6_outputs[676]));
    assign outputs[3071] = ~(layer6_outputs[353]);
    assign outputs[3072] = layer6_outputs[339];
    assign outputs[3073] = (layer6_outputs[1007]) ^ (layer6_outputs[1033]);
    assign outputs[3074] = layer6_outputs[2862];
    assign outputs[3075] = ~(layer6_outputs[241]);
    assign outputs[3076] = layer6_outputs[95];
    assign outputs[3077] = ~(layer6_outputs[2768]);
    assign outputs[3078] = ~((layer6_outputs[4291]) | (layer6_outputs[1088]));
    assign outputs[3079] = (layer6_outputs[3941]) | (layer6_outputs[137]);
    assign outputs[3080] = ~((layer6_outputs[4712]) ^ (layer6_outputs[3773]));
    assign outputs[3081] = ~(layer6_outputs[3068]);
    assign outputs[3082] = layer6_outputs[2403];
    assign outputs[3083] = (layer6_outputs[1933]) ^ (layer6_outputs[125]);
    assign outputs[3084] = ~(layer6_outputs[3090]);
    assign outputs[3085] = layer6_outputs[2858];
    assign outputs[3086] = ~(layer6_outputs[2816]);
    assign outputs[3087] = layer6_outputs[1796];
    assign outputs[3088] = layer6_outputs[2342];
    assign outputs[3089] = ~(layer6_outputs[4973]);
    assign outputs[3090] = ~(layer6_outputs[1569]);
    assign outputs[3091] = ~(layer6_outputs[603]);
    assign outputs[3092] = (layer6_outputs[2534]) & ~(layer6_outputs[2745]);
    assign outputs[3093] = ~(layer6_outputs[1524]);
    assign outputs[3094] = ~((layer6_outputs[3594]) ^ (layer6_outputs[4917]));
    assign outputs[3095] = (layer6_outputs[2743]) & ~(layer6_outputs[2694]);
    assign outputs[3096] = layer6_outputs[4785];
    assign outputs[3097] = layer6_outputs[4995];
    assign outputs[3098] = layer6_outputs[3830];
    assign outputs[3099] = ~(layer6_outputs[2810]);
    assign outputs[3100] = layer6_outputs[4499];
    assign outputs[3101] = ~(layer6_outputs[2935]);
    assign outputs[3102] = ~((layer6_outputs[596]) ^ (layer6_outputs[3300]));
    assign outputs[3103] = (layer6_outputs[2035]) ^ (layer6_outputs[4960]);
    assign outputs[3104] = layer6_outputs[2000];
    assign outputs[3105] = ~(layer6_outputs[4119]);
    assign outputs[3106] = layer6_outputs[565];
    assign outputs[3107] = layer6_outputs[65];
    assign outputs[3108] = (layer6_outputs[2445]) & ~(layer6_outputs[5020]);
    assign outputs[3109] = ~(layer6_outputs[1057]);
    assign outputs[3110] = (layer6_outputs[4945]) | (layer6_outputs[2974]);
    assign outputs[3111] = layer6_outputs[3775];
    assign outputs[3112] = layer6_outputs[1380];
    assign outputs[3113] = ~(layer6_outputs[3001]);
    assign outputs[3114] = (layer6_outputs[908]) & ~(layer6_outputs[4937]);
    assign outputs[3115] = layer6_outputs[3131];
    assign outputs[3116] = (layer6_outputs[1365]) ^ (layer6_outputs[1074]);
    assign outputs[3117] = ~(layer6_outputs[5082]);
    assign outputs[3118] = (layer6_outputs[1895]) ^ (layer6_outputs[582]);
    assign outputs[3119] = ~(layer6_outputs[2125]);
    assign outputs[3120] = ~(layer6_outputs[1753]);
    assign outputs[3121] = ~((layer6_outputs[3886]) ^ (layer6_outputs[971]));
    assign outputs[3122] = layer6_outputs[0];
    assign outputs[3123] = layer6_outputs[2453];
    assign outputs[3124] = layer6_outputs[2742];
    assign outputs[3125] = layer6_outputs[2948];
    assign outputs[3126] = ~((layer6_outputs[2278]) & (layer6_outputs[1700]));
    assign outputs[3127] = ~(layer6_outputs[663]);
    assign outputs[3128] = layer6_outputs[622];
    assign outputs[3129] = ~(layer6_outputs[4923]);
    assign outputs[3130] = (layer6_outputs[5113]) ^ (layer6_outputs[4373]);
    assign outputs[3131] = ~(layer6_outputs[727]);
    assign outputs[3132] = ~((layer6_outputs[4207]) ^ (layer6_outputs[4951]));
    assign outputs[3133] = (layer6_outputs[3696]) ^ (layer6_outputs[1]);
    assign outputs[3134] = layer6_outputs[1175];
    assign outputs[3135] = layer6_outputs[530];
    assign outputs[3136] = ~((layer6_outputs[1287]) & (layer6_outputs[4538]));
    assign outputs[3137] = layer6_outputs[1736];
    assign outputs[3138] = layer6_outputs[681];
    assign outputs[3139] = ~(layer6_outputs[2655]);
    assign outputs[3140] = layer6_outputs[2159];
    assign outputs[3141] = layer6_outputs[411];
    assign outputs[3142] = layer6_outputs[1134];
    assign outputs[3143] = (layer6_outputs[848]) ^ (layer6_outputs[1279]);
    assign outputs[3144] = layer6_outputs[3428];
    assign outputs[3145] = (layer6_outputs[3860]) | (layer6_outputs[3854]);
    assign outputs[3146] = (layer6_outputs[953]) ^ (layer6_outputs[1619]);
    assign outputs[3147] = ~(layer6_outputs[4313]);
    assign outputs[3148] = layer6_outputs[2767];
    assign outputs[3149] = layer6_outputs[895];
    assign outputs[3150] = layer6_outputs[1504];
    assign outputs[3151] = layer6_outputs[1965];
    assign outputs[3152] = layer6_outputs[1301];
    assign outputs[3153] = ~(layer6_outputs[3945]);
    assign outputs[3154] = layer6_outputs[3282];
    assign outputs[3155] = ~(layer6_outputs[5068]);
    assign outputs[3156] = (layer6_outputs[4805]) | (layer6_outputs[582]);
    assign outputs[3157] = ~(layer6_outputs[2873]);
    assign outputs[3158] = ~(layer6_outputs[3171]);
    assign outputs[3159] = layer6_outputs[1339];
    assign outputs[3160] = ~(layer6_outputs[591]) | (layer6_outputs[1030]);
    assign outputs[3161] = ~(layer6_outputs[3081]);
    assign outputs[3162] = ~((layer6_outputs[2953]) ^ (layer6_outputs[2859]));
    assign outputs[3163] = layer6_outputs[3056];
    assign outputs[3164] = layer6_outputs[5069];
    assign outputs[3165] = layer6_outputs[458];
    assign outputs[3166] = ~(layer6_outputs[484]) | (layer6_outputs[3481]);
    assign outputs[3167] = layer6_outputs[4776];
    assign outputs[3168] = ~((layer6_outputs[4522]) ^ (layer6_outputs[4058]));
    assign outputs[3169] = layer6_outputs[2639];
    assign outputs[3170] = layer6_outputs[2813];
    assign outputs[3171] = ~(layer6_outputs[3904]);
    assign outputs[3172] = ~((layer6_outputs[4008]) ^ (layer6_outputs[783]));
    assign outputs[3173] = (layer6_outputs[3895]) & ~(layer6_outputs[1214]);
    assign outputs[3174] = ~((layer6_outputs[1866]) ^ (layer6_outputs[759]));
    assign outputs[3175] = layer6_outputs[862];
    assign outputs[3176] = layer6_outputs[369];
    assign outputs[3177] = (layer6_outputs[3581]) & (layer6_outputs[5039]);
    assign outputs[3178] = layer6_outputs[2300];
    assign outputs[3179] = (layer6_outputs[2466]) & ~(layer6_outputs[4001]);
    assign outputs[3180] = (layer6_outputs[341]) & (layer6_outputs[4761]);
    assign outputs[3181] = layer6_outputs[5063];
    assign outputs[3182] = (layer6_outputs[580]) ^ (layer6_outputs[3267]);
    assign outputs[3183] = layer6_outputs[3411];
    assign outputs[3184] = (layer6_outputs[569]) & ~(layer6_outputs[3577]);
    assign outputs[3185] = ~(layer6_outputs[812]);
    assign outputs[3186] = ~(layer6_outputs[730]);
    assign outputs[3187] = ~(layer6_outputs[425]);
    assign outputs[3188] = ~(layer6_outputs[240]);
    assign outputs[3189] = layer6_outputs[805];
    assign outputs[3190] = (layer6_outputs[4709]) ^ (layer6_outputs[4022]);
    assign outputs[3191] = layer6_outputs[1888];
    assign outputs[3192] = (layer6_outputs[4860]) ^ (layer6_outputs[1238]);
    assign outputs[3193] = layer6_outputs[2151];
    assign outputs[3194] = layer6_outputs[4335];
    assign outputs[3195] = ~((layer6_outputs[36]) | (layer6_outputs[1342]));
    assign outputs[3196] = (layer6_outputs[3777]) ^ (layer6_outputs[3990]);
    assign outputs[3197] = layer6_outputs[3476];
    assign outputs[3198] = ~(layer6_outputs[2929]);
    assign outputs[3199] = layer6_outputs[1431];
    assign outputs[3200] = layer6_outputs[1448];
    assign outputs[3201] = ~((layer6_outputs[36]) ^ (layer6_outputs[3250]));
    assign outputs[3202] = layer6_outputs[4398];
    assign outputs[3203] = ~(layer6_outputs[640]);
    assign outputs[3204] = (layer6_outputs[2949]) ^ (layer6_outputs[2752]);
    assign outputs[3205] = (layer6_outputs[4913]) ^ (layer6_outputs[1753]);
    assign outputs[3206] = ~(layer6_outputs[3944]);
    assign outputs[3207] = (layer6_outputs[1111]) | (layer6_outputs[3357]);
    assign outputs[3208] = (layer6_outputs[3463]) ^ (layer6_outputs[4687]);
    assign outputs[3209] = ~(layer6_outputs[2328]);
    assign outputs[3210] = ~(layer6_outputs[1508]);
    assign outputs[3211] = layer6_outputs[4401];
    assign outputs[3212] = layer6_outputs[3139];
    assign outputs[3213] = layer6_outputs[3991];
    assign outputs[3214] = ~(layer6_outputs[4203]);
    assign outputs[3215] = ~(layer6_outputs[1689]);
    assign outputs[3216] = layer6_outputs[1471];
    assign outputs[3217] = ~(layer6_outputs[4663]);
    assign outputs[3218] = (layer6_outputs[2576]) ^ (layer6_outputs[4732]);
    assign outputs[3219] = ~(layer6_outputs[838]);
    assign outputs[3220] = layer6_outputs[5112];
    assign outputs[3221] = (layer6_outputs[1589]) ^ (layer6_outputs[3010]);
    assign outputs[3222] = (layer6_outputs[4009]) & ~(layer6_outputs[4637]);
    assign outputs[3223] = (layer6_outputs[2565]) & ~(layer6_outputs[3249]);
    assign outputs[3224] = ~(layer6_outputs[3265]);
    assign outputs[3225] = (layer6_outputs[4468]) & (layer6_outputs[2854]);
    assign outputs[3226] = layer6_outputs[4535];
    assign outputs[3227] = layer6_outputs[3934];
    assign outputs[3228] = ~(layer6_outputs[3442]);
    assign outputs[3229] = ~((layer6_outputs[1522]) ^ (layer6_outputs[1043]));
    assign outputs[3230] = layer6_outputs[1622];
    assign outputs[3231] = (layer6_outputs[3853]) & (layer6_outputs[5088]);
    assign outputs[3232] = ~(layer6_outputs[3558]);
    assign outputs[3233] = ~(layer6_outputs[3643]);
    assign outputs[3234] = ~(layer6_outputs[4936]) | (layer6_outputs[4150]);
    assign outputs[3235] = layer6_outputs[4999];
    assign outputs[3236] = ~(layer6_outputs[738]);
    assign outputs[3237] = ~(layer6_outputs[3347]);
    assign outputs[3238] = ~((layer6_outputs[1546]) ^ (layer6_outputs[278]));
    assign outputs[3239] = ~(layer6_outputs[1443]);
    assign outputs[3240] = (layer6_outputs[4597]) & ~(layer6_outputs[1103]);
    assign outputs[3241] = ~(layer6_outputs[3075]);
    assign outputs[3242] = ~(layer6_outputs[4067]);
    assign outputs[3243] = layer6_outputs[3522];
    assign outputs[3244] = layer6_outputs[1717];
    assign outputs[3245] = ~(layer6_outputs[1979]);
    assign outputs[3246] = ~(layer6_outputs[4626]);
    assign outputs[3247] = layer6_outputs[1759];
    assign outputs[3248] = ~(layer6_outputs[4909]);
    assign outputs[3249] = ~(layer6_outputs[4210]);
    assign outputs[3250] = ~(layer6_outputs[2348]);
    assign outputs[3251] = layer6_outputs[2586];
    assign outputs[3252] = layer6_outputs[1349];
    assign outputs[3253] = ~(layer6_outputs[3936]);
    assign outputs[3254] = layer6_outputs[4588];
    assign outputs[3255] = layer6_outputs[120];
    assign outputs[3256] = layer6_outputs[3862];
    assign outputs[3257] = layer6_outputs[4021];
    assign outputs[3258] = layer6_outputs[226];
    assign outputs[3259] = ~(layer6_outputs[2197]);
    assign outputs[3260] = ~(layer6_outputs[3419]);
    assign outputs[3261] = ~((layer6_outputs[3770]) ^ (layer6_outputs[644]));
    assign outputs[3262] = ~(layer6_outputs[5020]);
    assign outputs[3263] = ~((layer6_outputs[3743]) ^ (layer6_outputs[4262]));
    assign outputs[3264] = layer6_outputs[4068];
    assign outputs[3265] = ~(layer6_outputs[1237]);
    assign outputs[3266] = (layer6_outputs[2122]) & (layer6_outputs[4120]);
    assign outputs[3267] = ~((layer6_outputs[553]) ^ (layer6_outputs[344]));
    assign outputs[3268] = ~(layer6_outputs[2711]) | (layer6_outputs[1784]);
    assign outputs[3269] = ~(layer6_outputs[3001]);
    assign outputs[3270] = layer6_outputs[1928];
    assign outputs[3271] = ~((layer6_outputs[1976]) ^ (layer6_outputs[4255]));
    assign outputs[3272] = layer6_outputs[3324];
    assign outputs[3273] = layer6_outputs[1172];
    assign outputs[3274] = ~(layer6_outputs[3171]);
    assign outputs[3275] = layer6_outputs[3456];
    assign outputs[3276] = ~((layer6_outputs[5093]) ^ (layer6_outputs[2762]));
    assign outputs[3277] = layer6_outputs[333];
    assign outputs[3278] = ~(layer6_outputs[128]);
    assign outputs[3279] = ~(layer6_outputs[2524]);
    assign outputs[3280] = layer6_outputs[1071];
    assign outputs[3281] = ~(layer6_outputs[1095]);
    assign outputs[3282] = ~(layer6_outputs[3318]);
    assign outputs[3283] = (layer6_outputs[3896]) & (layer6_outputs[1596]);
    assign outputs[3284] = layer6_outputs[3021];
    assign outputs[3285] = layer6_outputs[816];
    assign outputs[3286] = ~(layer6_outputs[4086]);
    assign outputs[3287] = ~(layer6_outputs[2590]);
    assign outputs[3288] = ~((layer6_outputs[1759]) ^ (layer6_outputs[4427]));
    assign outputs[3289] = layer6_outputs[2738];
    assign outputs[3290] = ~(layer6_outputs[2034]);
    assign outputs[3291] = (layer6_outputs[1481]) & ~(layer6_outputs[1854]);
    assign outputs[3292] = (layer6_outputs[1078]) & (layer6_outputs[4057]);
    assign outputs[3293] = ~(layer6_outputs[179]);
    assign outputs[3294] = ~((layer6_outputs[3237]) & (layer6_outputs[265]));
    assign outputs[3295] = (layer6_outputs[3541]) ^ (layer6_outputs[1986]);
    assign outputs[3296] = ~((layer6_outputs[2682]) ^ (layer6_outputs[2775]));
    assign outputs[3297] = layer6_outputs[2171];
    assign outputs[3298] = layer6_outputs[5017];
    assign outputs[3299] = layer6_outputs[4028];
    assign outputs[3300] = (layer6_outputs[138]) ^ (layer6_outputs[1961]);
    assign outputs[3301] = ~(layer6_outputs[179]);
    assign outputs[3302] = layer6_outputs[3530];
    assign outputs[3303] = ~((layer6_outputs[2060]) ^ (layer6_outputs[1948]));
    assign outputs[3304] = layer6_outputs[650];
    assign outputs[3305] = layer6_outputs[1515];
    assign outputs[3306] = ~(layer6_outputs[3962]);
    assign outputs[3307] = ~(layer6_outputs[2781]);
    assign outputs[3308] = (layer6_outputs[162]) & ~(layer6_outputs[2290]);
    assign outputs[3309] = ~((layer6_outputs[3199]) & (layer6_outputs[433]));
    assign outputs[3310] = layer6_outputs[2263];
    assign outputs[3311] = (layer6_outputs[3780]) & ~(layer6_outputs[453]);
    assign outputs[3312] = ~(layer6_outputs[448]);
    assign outputs[3313] = layer6_outputs[1588];
    assign outputs[3314] = ~(layer6_outputs[4405]);
    assign outputs[3315] = layer6_outputs[4015];
    assign outputs[3316] = layer6_outputs[2946];
    assign outputs[3317] = (layer6_outputs[291]) & ~(layer6_outputs[2975]);
    assign outputs[3318] = ~(layer6_outputs[1600]);
    assign outputs[3319] = ~(layer6_outputs[2783]);
    assign outputs[3320] = ~(layer6_outputs[3466]);
    assign outputs[3321] = layer6_outputs[1186];
    assign outputs[3322] = ~(layer6_outputs[3655]) | (layer6_outputs[2605]);
    assign outputs[3323] = layer6_outputs[3560];
    assign outputs[3324] = ~(layer6_outputs[947]);
    assign outputs[3325] = layer6_outputs[3161];
    assign outputs[3326] = layer6_outputs[4634];
    assign outputs[3327] = ~(layer6_outputs[155]);
    assign outputs[3328] = ~(layer6_outputs[4227]);
    assign outputs[3329] = ~(layer6_outputs[2389]);
    assign outputs[3330] = (layer6_outputs[2770]) ^ (layer6_outputs[4988]);
    assign outputs[3331] = layer6_outputs[2382];
    assign outputs[3332] = layer6_outputs[652];
    assign outputs[3333] = ~((layer6_outputs[206]) ^ (layer6_outputs[2434]));
    assign outputs[3334] = ~(layer6_outputs[3709]);
    assign outputs[3335] = ~((layer6_outputs[1145]) & (layer6_outputs[4299]));
    assign outputs[3336] = ~(layer6_outputs[2283]) | (layer6_outputs[4841]);
    assign outputs[3337] = ~(layer6_outputs[4403]);
    assign outputs[3338] = layer6_outputs[3979];
    assign outputs[3339] = ~(layer6_outputs[3400]);
    assign outputs[3340] = ~(layer6_outputs[186]);
    assign outputs[3341] = layer6_outputs[1280];
    assign outputs[3342] = ~((layer6_outputs[2533]) & (layer6_outputs[3819]));
    assign outputs[3343] = ~(layer6_outputs[4844]);
    assign outputs[3344] = ~(layer6_outputs[969]);
    assign outputs[3345] = (layer6_outputs[3187]) ^ (layer6_outputs[3141]);
    assign outputs[3346] = ~((layer6_outputs[3303]) | (layer6_outputs[1970]));
    assign outputs[3347] = layer6_outputs[2379];
    assign outputs[3348] = layer6_outputs[1846];
    assign outputs[3349] = layer6_outputs[2967];
    assign outputs[3350] = layer6_outputs[544];
    assign outputs[3351] = ~(layer6_outputs[515]) | (layer6_outputs[1269]);
    assign outputs[3352] = ~(layer6_outputs[293]);
    assign outputs[3353] = ~(layer6_outputs[1131]);
    assign outputs[3354] = ~(layer6_outputs[2750]);
    assign outputs[3355] = ~(layer6_outputs[2581]);
    assign outputs[3356] = layer6_outputs[4327];
    assign outputs[3357] = (layer6_outputs[997]) ^ (layer6_outputs[639]);
    assign outputs[3358] = ~((layer6_outputs[2242]) | (layer6_outputs[753]));
    assign outputs[3359] = ~((layer6_outputs[3586]) & (layer6_outputs[1716]));
    assign outputs[3360] = ~(layer6_outputs[4948]);
    assign outputs[3361] = layer6_outputs[1049];
    assign outputs[3362] = layer6_outputs[5040];
    assign outputs[3363] = ~(layer6_outputs[2247]);
    assign outputs[3364] = ~(layer6_outputs[4295]);
    assign outputs[3365] = ~((layer6_outputs[4309]) ^ (layer6_outputs[921]));
    assign outputs[3366] = (layer6_outputs[2431]) & ~(layer6_outputs[2808]);
    assign outputs[3367] = layer6_outputs[1742];
    assign outputs[3368] = ~(layer6_outputs[3367]);
    assign outputs[3369] = ~((layer6_outputs[3403]) | (layer6_outputs[4096]));
    assign outputs[3370] = ~(layer6_outputs[4631]);
    assign outputs[3371] = ~(layer6_outputs[1754]);
    assign outputs[3372] = layer6_outputs[1823];
    assign outputs[3373] = ~((layer6_outputs[1411]) | (layer6_outputs[3190]));
    assign outputs[3374] = ~(layer6_outputs[1287]);
    assign outputs[3375] = ~(layer6_outputs[2287]);
    assign outputs[3376] = ~((layer6_outputs[1011]) & (layer6_outputs[1564]));
    assign outputs[3377] = (layer6_outputs[2939]) ^ (layer6_outputs[4860]);
    assign outputs[3378] = layer6_outputs[1846];
    assign outputs[3379] = ~(layer6_outputs[2486]);
    assign outputs[3380] = ~(layer6_outputs[469]);
    assign outputs[3381] = ~((layer6_outputs[3928]) ^ (layer6_outputs[3667]));
    assign outputs[3382] = (layer6_outputs[2371]) & ~(layer6_outputs[1335]);
    assign outputs[3383] = ~(layer6_outputs[3925]);
    assign outputs[3384] = (layer6_outputs[2353]) ^ (layer6_outputs[2483]);
    assign outputs[3385] = ~(layer6_outputs[2160]) | (layer6_outputs[4553]);
    assign outputs[3386] = ~(layer6_outputs[839]);
    assign outputs[3387] = (layer6_outputs[76]) | (layer6_outputs[4858]);
    assign outputs[3388] = (layer6_outputs[1259]) & (layer6_outputs[2317]);
    assign outputs[3389] = ~(layer6_outputs[4746]);
    assign outputs[3390] = ~(layer6_outputs[4485]);
    assign outputs[3391] = ~(layer6_outputs[4020]);
    assign outputs[3392] = layer6_outputs[3098];
    assign outputs[3393] = ~(layer6_outputs[1390]);
    assign outputs[3394] = ~(layer6_outputs[4367]);
    assign outputs[3395] = layer6_outputs[2634];
    assign outputs[3396] = ~((layer6_outputs[307]) ^ (layer6_outputs[4919]));
    assign outputs[3397] = layer6_outputs[1317];
    assign outputs[3398] = ~((layer6_outputs[4530]) ^ (layer6_outputs[4105]));
    assign outputs[3399] = layer6_outputs[2885];
    assign outputs[3400] = (layer6_outputs[4658]) & (layer6_outputs[698]);
    assign outputs[3401] = (layer6_outputs[4389]) ^ (layer6_outputs[806]);
    assign outputs[3402] = ~(layer6_outputs[5106]);
    assign outputs[3403] = (layer6_outputs[1367]) | (layer6_outputs[3857]);
    assign outputs[3404] = ~((layer6_outputs[795]) ^ (layer6_outputs[1801]));
    assign outputs[3405] = ~(layer6_outputs[2497]);
    assign outputs[3406] = (layer6_outputs[3314]) & ~(layer6_outputs[1337]);
    assign outputs[3407] = layer6_outputs[1469];
    assign outputs[3408] = ~(layer6_outputs[4819]);
    assign outputs[3409] = (layer6_outputs[3446]) | (layer6_outputs[1374]);
    assign outputs[3410] = (layer6_outputs[2793]) & (layer6_outputs[4123]);
    assign outputs[3411] = layer6_outputs[1927];
    assign outputs[3412] = layer6_outputs[4742];
    assign outputs[3413] = ~(layer6_outputs[1766]);
    assign outputs[3414] = (layer6_outputs[287]) & ~(layer6_outputs[3552]);
    assign outputs[3415] = ~(layer6_outputs[229]);
    assign outputs[3416] = layer6_outputs[4353];
    assign outputs[3417] = ~(layer6_outputs[3617]);
    assign outputs[3418] = ~(layer6_outputs[1672]);
    assign outputs[3419] = layer6_outputs[2807];
    assign outputs[3420] = ~(layer6_outputs[2064]);
    assign outputs[3421] = ~(layer6_outputs[4737]);
    assign outputs[3422] = layer6_outputs[1008];
    assign outputs[3423] = ~(layer6_outputs[2750]);
    assign outputs[3424] = ~(layer6_outputs[634]);
    assign outputs[3425] = ~(layer6_outputs[4302]) | (layer6_outputs[948]);
    assign outputs[3426] = layer6_outputs[4244];
    assign outputs[3427] = ~(layer6_outputs[1495]);
    assign outputs[3428] = layer6_outputs[2946];
    assign outputs[3429] = layer6_outputs[1546];
    assign outputs[3430] = ~(layer6_outputs[2719]);
    assign outputs[3431] = ~(layer6_outputs[186]);
    assign outputs[3432] = ~((layer6_outputs[4651]) ^ (layer6_outputs[2774]));
    assign outputs[3433] = layer6_outputs[4912];
    assign outputs[3434] = layer6_outputs[1555];
    assign outputs[3435] = layer6_outputs[140];
    assign outputs[3436] = layer6_outputs[1911];
    assign outputs[3437] = ~(layer6_outputs[4319]);
    assign outputs[3438] = (layer6_outputs[4842]) & (layer6_outputs[1100]);
    assign outputs[3439] = ~(layer6_outputs[4727]);
    assign outputs[3440] = layer6_outputs[328];
    assign outputs[3441] = (layer6_outputs[1348]) & ~(layer6_outputs[1415]);
    assign outputs[3442] = ~((layer6_outputs[2879]) ^ (layer6_outputs[1724]));
    assign outputs[3443] = layer6_outputs[3241];
    assign outputs[3444] = layer6_outputs[1715];
    assign outputs[3445] = layer6_outputs[48];
    assign outputs[3446] = ~(layer6_outputs[4647]) | (layer6_outputs[2292]);
    assign outputs[3447] = ~(layer6_outputs[4802]);
    assign outputs[3448] = layer6_outputs[3328];
    assign outputs[3449] = layer6_outputs[4459];
    assign outputs[3450] = ~(layer6_outputs[3452]);
    assign outputs[3451] = (layer6_outputs[3448]) | (layer6_outputs[4211]);
    assign outputs[3452] = ~(layer6_outputs[3899]);
    assign outputs[3453] = ~(layer6_outputs[5097]);
    assign outputs[3454] = layer6_outputs[1785];
    assign outputs[3455] = layer6_outputs[1074];
    assign outputs[3456] = layer6_outputs[2647];
    assign outputs[3457] = layer6_outputs[4800];
    assign outputs[3458] = (layer6_outputs[836]) & ~(layer6_outputs[3998]);
    assign outputs[3459] = ~(layer6_outputs[3983]);
    assign outputs[3460] = layer6_outputs[3720];
    assign outputs[3461] = layer6_outputs[328];
    assign outputs[3462] = ~(layer6_outputs[3721]);
    assign outputs[3463] = layer6_outputs[4004];
    assign outputs[3464] = layer6_outputs[3938];
    assign outputs[3465] = ~(layer6_outputs[2929]);
    assign outputs[3466] = ~((layer6_outputs[1768]) ^ (layer6_outputs[1219]));
    assign outputs[3467] = (layer6_outputs[4608]) & ~(layer6_outputs[3832]);
    assign outputs[3468] = layer6_outputs[3627];
    assign outputs[3469] = layer6_outputs[223];
    assign outputs[3470] = layer6_outputs[4185];
    assign outputs[3471] = layer6_outputs[350];
    assign outputs[3472] = ~(layer6_outputs[127]);
    assign outputs[3473] = ~(layer6_outputs[4293]);
    assign outputs[3474] = ~(layer6_outputs[4477]);
    assign outputs[3475] = ~(layer6_outputs[5029]);
    assign outputs[3476] = ~((layer6_outputs[4161]) ^ (layer6_outputs[3389]));
    assign outputs[3477] = layer6_outputs[1704];
    assign outputs[3478] = layer6_outputs[2048];
    assign outputs[3479] = ~(layer6_outputs[952]);
    assign outputs[3480] = layer6_outputs[2566];
    assign outputs[3481] = layer6_outputs[2434];
    assign outputs[3482] = layer6_outputs[1115];
    assign outputs[3483] = ~(layer6_outputs[2412]) | (layer6_outputs[2067]);
    assign outputs[3484] = layer6_outputs[4185];
    assign outputs[3485] = (layer6_outputs[124]) | (layer6_outputs[5091]);
    assign outputs[3486] = (layer6_outputs[2332]) & ~(layer6_outputs[1215]);
    assign outputs[3487] = ~(layer6_outputs[198]) | (layer6_outputs[2919]);
    assign outputs[3488] = ~(layer6_outputs[106]) | (layer6_outputs[3746]);
    assign outputs[3489] = layer6_outputs[4283];
    assign outputs[3490] = ~(layer6_outputs[3800]);
    assign outputs[3491] = ~((layer6_outputs[523]) ^ (layer6_outputs[3359]));
    assign outputs[3492] = ~(layer6_outputs[4984]);
    assign outputs[3493] = ~(layer6_outputs[2385]);
    assign outputs[3494] = layer6_outputs[337];
    assign outputs[3495] = ~(layer6_outputs[1040]);
    assign outputs[3496] = ~(layer6_outputs[946]);
    assign outputs[3497] = ~((layer6_outputs[3350]) ^ (layer6_outputs[1696]));
    assign outputs[3498] = layer6_outputs[1181];
    assign outputs[3499] = layer6_outputs[1925];
    assign outputs[3500] = ~(layer6_outputs[466]);
    assign outputs[3501] = ~((layer6_outputs[2839]) ^ (layer6_outputs[2101]));
    assign outputs[3502] = layer6_outputs[2587];
    assign outputs[3503] = (layer6_outputs[209]) & ~(layer6_outputs[1905]);
    assign outputs[3504] = ~(layer6_outputs[3882]);
    assign outputs[3505] = ~(layer6_outputs[915]);
    assign outputs[3506] = ~(layer6_outputs[3142]);
    assign outputs[3507] = layer6_outputs[4928];
    assign outputs[3508] = ~(layer6_outputs[3919]);
    assign outputs[3509] = ~(layer6_outputs[3336]);
    assign outputs[3510] = layer6_outputs[2888];
    assign outputs[3511] = (layer6_outputs[4042]) ^ (layer6_outputs[3758]);
    assign outputs[3512] = ~(layer6_outputs[3294]);
    assign outputs[3513] = ~((layer6_outputs[3071]) ^ (layer6_outputs[2033]));
    assign outputs[3514] = (layer6_outputs[1752]) ^ (layer6_outputs[1181]);
    assign outputs[3515] = ~(layer6_outputs[4876]);
    assign outputs[3516] = ~((layer6_outputs[2358]) ^ (layer6_outputs[4664]));
    assign outputs[3517] = (layer6_outputs[3463]) ^ (layer6_outputs[1984]);
    assign outputs[3518] = (layer6_outputs[3732]) | (layer6_outputs[2520]);
    assign outputs[3519] = ~(layer6_outputs[3386]);
    assign outputs[3520] = (layer6_outputs[2433]) ^ (layer6_outputs[1003]);
    assign outputs[3521] = layer6_outputs[4662];
    assign outputs[3522] = (layer6_outputs[3883]) & (layer6_outputs[1012]);
    assign outputs[3523] = (layer6_outputs[2673]) & ~(layer6_outputs[2228]);
    assign outputs[3524] = ~(layer6_outputs[2931]);
    assign outputs[3525] = layer6_outputs[3652];
    assign outputs[3526] = layer6_outputs[3285];
    assign outputs[3527] = ~(layer6_outputs[5080]);
    assign outputs[3528] = ~(layer6_outputs[169]);
    assign outputs[3529] = ~(layer6_outputs[2054]);
    assign outputs[3530] = layer6_outputs[725];
    assign outputs[3531] = ~(layer6_outputs[3321]);
    assign outputs[3532] = layer6_outputs[2853];
    assign outputs[3533] = ~(layer6_outputs[20]);
    assign outputs[3534] = ~(layer6_outputs[3097]);
    assign outputs[3535] = ~(layer6_outputs[2077]);
    assign outputs[3536] = ~((layer6_outputs[1914]) & (layer6_outputs[3713]));
    assign outputs[3537] = (layer6_outputs[4740]) & (layer6_outputs[3550]);
    assign outputs[3538] = ~(layer6_outputs[2541]);
    assign outputs[3539] = layer6_outputs[4589];
    assign outputs[3540] = (layer6_outputs[357]) ^ (layer6_outputs[3148]);
    assign outputs[3541] = layer6_outputs[1762];
    assign outputs[3542] = layer6_outputs[1627];
    assign outputs[3543] = layer6_outputs[61];
    assign outputs[3544] = (layer6_outputs[4832]) & ~(layer6_outputs[2335]);
    assign outputs[3545] = ~((layer6_outputs[2850]) & (layer6_outputs[2207]));
    assign outputs[3546] = ~(layer6_outputs[4773]);
    assign outputs[3547] = layer6_outputs[3366];
    assign outputs[3548] = ~(layer6_outputs[2365]);
    assign outputs[3549] = layer6_outputs[1884];
    assign outputs[3550] = layer6_outputs[3368];
    assign outputs[3551] = layer6_outputs[2307];
    assign outputs[3552] = layer6_outputs[4068];
    assign outputs[3553] = (layer6_outputs[1908]) & ~(layer6_outputs[1125]);
    assign outputs[3554] = ~(layer6_outputs[4948]);
    assign outputs[3555] = ~(layer6_outputs[2481]);
    assign outputs[3556] = (layer6_outputs[2306]) ^ (layer6_outputs[1971]);
    assign outputs[3557] = (layer6_outputs[3253]) ^ (layer6_outputs[4426]);
    assign outputs[3558] = ~((layer6_outputs[3000]) ^ (layer6_outputs[3661]));
    assign outputs[3559] = layer6_outputs[4882];
    assign outputs[3560] = layer6_outputs[872];
    assign outputs[3561] = layer6_outputs[2523];
    assign outputs[3562] = ~(layer6_outputs[358]);
    assign outputs[3563] = layer6_outputs[262];
    assign outputs[3564] = layer6_outputs[517];
    assign outputs[3565] = ~(layer6_outputs[4177]);
    assign outputs[3566] = layer6_outputs[4990];
    assign outputs[3567] = ~(layer6_outputs[4909]);
    assign outputs[3568] = layer6_outputs[4274];
    assign outputs[3569] = layer6_outputs[2716];
    assign outputs[3570] = ~((layer6_outputs[1049]) ^ (layer6_outputs[1215]));
    assign outputs[3571] = (layer6_outputs[251]) ^ (layer6_outputs[2960]);
    assign outputs[3572] = ~(layer6_outputs[1229]);
    assign outputs[3573] = ~((layer6_outputs[286]) ^ (layer6_outputs[3034]));
    assign outputs[3574] = (layer6_outputs[4951]) | (layer6_outputs[2211]);
    assign outputs[3575] = ~(layer6_outputs[4474]);
    assign outputs[3576] = (layer6_outputs[5032]) ^ (layer6_outputs[29]);
    assign outputs[3577] = ~(layer6_outputs[1094]);
    assign outputs[3578] = ~(layer6_outputs[4181]);
    assign outputs[3579] = layer6_outputs[3858];
    assign outputs[3580] = (layer6_outputs[1321]) & ~(layer6_outputs[1776]);
    assign outputs[3581] = ~((layer6_outputs[241]) | (layer6_outputs[1387]));
    assign outputs[3582] = ~(layer6_outputs[4166]);
    assign outputs[3583] = layer6_outputs[3517];
    assign outputs[3584] = layer6_outputs[4837];
    assign outputs[3585] = layer6_outputs[1426];
    assign outputs[3586] = layer6_outputs[2449];
    assign outputs[3587] = ~(layer6_outputs[4536]);
    assign outputs[3588] = layer6_outputs[1359];
    assign outputs[3589] = ~((layer6_outputs[2106]) | (layer6_outputs[12]));
    assign outputs[3590] = layer6_outputs[4356];
    assign outputs[3591] = layer6_outputs[959];
    assign outputs[3592] = layer6_outputs[1950];
    assign outputs[3593] = layer6_outputs[3090];
    assign outputs[3594] = ~((layer6_outputs[3137]) ^ (layer6_outputs[1784]));
    assign outputs[3595] = layer6_outputs[1754];
    assign outputs[3596] = ~(layer6_outputs[1679]);
    assign outputs[3597] = layer6_outputs[4690];
    assign outputs[3598] = ~(layer6_outputs[2179]);
    assign outputs[3599] = ~(layer6_outputs[562]);
    assign outputs[3600] = ~(layer6_outputs[3888]);
    assign outputs[3601] = ~(layer6_outputs[2717]);
    assign outputs[3602] = ~((layer6_outputs[2041]) | (layer6_outputs[1772]));
    assign outputs[3603] = layer6_outputs[1794];
    assign outputs[3604] = (layer6_outputs[497]) & ~(layer6_outputs[159]);
    assign outputs[3605] = (layer6_outputs[994]) & ~(layer6_outputs[773]);
    assign outputs[3606] = layer6_outputs[4331];
    assign outputs[3607] = (layer6_outputs[4892]) ^ (layer6_outputs[4525]);
    assign outputs[3608] = ~((layer6_outputs[1332]) | (layer6_outputs[390]));
    assign outputs[3609] = ~(layer6_outputs[514]);
    assign outputs[3610] = ~((layer6_outputs[2220]) ^ (layer6_outputs[4736]));
    assign outputs[3611] = layer6_outputs[3777];
    assign outputs[3612] = (layer6_outputs[4866]) ^ (layer6_outputs[785]);
    assign outputs[3613] = ~(layer6_outputs[1977]);
    assign outputs[3614] = layer6_outputs[2844];
    assign outputs[3615] = layer6_outputs[1480];
    assign outputs[3616] = (layer6_outputs[1850]) & ~(layer6_outputs[3414]);
    assign outputs[3617] = ~((layer6_outputs[4883]) ^ (layer6_outputs[4918]));
    assign outputs[3618] = ~(layer6_outputs[2299]);
    assign outputs[3619] = ~((layer6_outputs[2088]) ^ (layer6_outputs[3805]));
    assign outputs[3620] = ~(layer6_outputs[5118]);
    assign outputs[3621] = ~(layer6_outputs[419]);
    assign outputs[3622] = (layer6_outputs[433]) ^ (layer6_outputs[1525]);
    assign outputs[3623] = ~(layer6_outputs[2318]);
    assign outputs[3624] = ~(layer6_outputs[143]);
    assign outputs[3625] = layer6_outputs[462];
    assign outputs[3626] = layer6_outputs[3692];
    assign outputs[3627] = layer6_outputs[3219];
    assign outputs[3628] = layer6_outputs[236];
    assign outputs[3629] = ~(layer6_outputs[2258]);
    assign outputs[3630] = (layer6_outputs[3881]) & ~(layer6_outputs[2404]);
    assign outputs[3631] = ~(layer6_outputs[4768]);
    assign outputs[3632] = layer6_outputs[1113];
    assign outputs[3633] = layer6_outputs[3134];
    assign outputs[3634] = layer6_outputs[3809];
    assign outputs[3635] = ~(layer6_outputs[4676]);
    assign outputs[3636] = ~(layer6_outputs[2066]);
    assign outputs[3637] = ~(layer6_outputs[187]);
    assign outputs[3638] = layer6_outputs[4782];
    assign outputs[3639] = (layer6_outputs[1746]) | (layer6_outputs[2578]);
    assign outputs[3640] = layer6_outputs[3835];
    assign outputs[3641] = layer6_outputs[1737];
    assign outputs[3642] = layer6_outputs[4683];
    assign outputs[3643] = ~(layer6_outputs[4270]) | (layer6_outputs[1542]);
    assign outputs[3644] = ~(layer6_outputs[3614]);
    assign outputs[3645] = ~(layer6_outputs[168]);
    assign outputs[3646] = ~(layer6_outputs[2049]);
    assign outputs[3647] = ~(layer6_outputs[4780]);
    assign outputs[3648] = ~(layer6_outputs[1529]);
    assign outputs[3649] = ~(layer6_outputs[3443]);
    assign outputs[3650] = (layer6_outputs[695]) & ~(layer6_outputs[21]);
    assign outputs[3651] = ~(layer6_outputs[3310]) | (layer6_outputs[4899]);
    assign outputs[3652] = layer6_outputs[2138];
    assign outputs[3653] = (layer6_outputs[2970]) & ~(layer6_outputs[1813]);
    assign outputs[3654] = ~(layer6_outputs[130]);
    assign outputs[3655] = ~(layer6_outputs[4651]);
    assign outputs[3656] = layer6_outputs[942];
    assign outputs[3657] = ~(layer6_outputs[2100]);
    assign outputs[3658] = ~(layer6_outputs[2010]);
    assign outputs[3659] = layer6_outputs[3967];
    assign outputs[3660] = layer6_outputs[1133];
    assign outputs[3661] = layer6_outputs[2150];
    assign outputs[3662] = layer6_outputs[2759];
    assign outputs[3663] = ~(layer6_outputs[2200]);
    assign outputs[3664] = ~(layer6_outputs[4287]);
    assign outputs[3665] = layer6_outputs[660];
    assign outputs[3666] = ~(layer6_outputs[3568]);
    assign outputs[3667] = (layer6_outputs[1208]) & ~(layer6_outputs[4686]);
    assign outputs[3668] = ~((layer6_outputs[1161]) ^ (layer6_outputs[1993]));
    assign outputs[3669] = ~(layer6_outputs[868]);
    assign outputs[3670] = ~(layer6_outputs[1308]);
    assign outputs[3671] = (layer6_outputs[2806]) ^ (layer6_outputs[4045]);
    assign outputs[3672] = ~(layer6_outputs[2179]);
    assign outputs[3673] = ~(layer6_outputs[1482]);
    assign outputs[3674] = (layer6_outputs[1187]) & ~(layer6_outputs[1497]);
    assign outputs[3675] = ~((layer6_outputs[3172]) ^ (layer6_outputs[5100]));
    assign outputs[3676] = layer6_outputs[3338];
    assign outputs[3677] = ~(layer6_outputs[3108]);
    assign outputs[3678] = layer6_outputs[4711];
    assign outputs[3679] = layer6_outputs[4190];
    assign outputs[3680] = ~(layer6_outputs[2226]);
    assign outputs[3681] = ~(layer6_outputs[4932]);
    assign outputs[3682] = layer6_outputs[3993];
    assign outputs[3683] = layer6_outputs[3306];
    assign outputs[3684] = layer6_outputs[177];
    assign outputs[3685] = ~((layer6_outputs[1104]) | (layer6_outputs[1512]));
    assign outputs[3686] = ~(layer6_outputs[3826]);
    assign outputs[3687] = ~(layer6_outputs[1607]);
    assign outputs[3688] = ~(layer6_outputs[1225]);
    assign outputs[3689] = ~((layer6_outputs[2095]) ^ (layer6_outputs[3843]));
    assign outputs[3690] = ~((layer6_outputs[2134]) | (layer6_outputs[562]));
    assign outputs[3691] = ~(layer6_outputs[892]);
    assign outputs[3692] = ~(layer6_outputs[3620]);
    assign outputs[3693] = layer6_outputs[234];
    assign outputs[3694] = ~((layer6_outputs[2983]) & (layer6_outputs[2714]));
    assign outputs[3695] = ~((layer6_outputs[1002]) & (layer6_outputs[1254]));
    assign outputs[3696] = (layer6_outputs[4929]) & ~(layer6_outputs[4007]);
    assign outputs[3697] = layer6_outputs[3957];
    assign outputs[3698] = layer6_outputs[2261];
    assign outputs[3699] = (layer6_outputs[4356]) & ~(layer6_outputs[4095]);
    assign outputs[3700] = layer6_outputs[4872];
    assign outputs[3701] = ~(layer6_outputs[3117]);
    assign outputs[3702] = ~(layer6_outputs[1805]);
    assign outputs[3703] = layer6_outputs[4723];
    assign outputs[3704] = ~((layer6_outputs[3972]) | (layer6_outputs[204]));
    assign outputs[3705] = ~(layer6_outputs[3476]);
    assign outputs[3706] = ~(layer6_outputs[2643]);
    assign outputs[3707] = ~((layer6_outputs[2245]) ^ (layer6_outputs[1671]));
    assign outputs[3708] = layer6_outputs[4147];
    assign outputs[3709] = layer6_outputs[4981];
    assign outputs[3710] = ~(layer6_outputs[3162]);
    assign outputs[3711] = ~(layer6_outputs[3845]);
    assign outputs[3712] = ~(layer6_outputs[1903]);
    assign outputs[3713] = layer6_outputs[1811];
    assign outputs[3714] = layer6_outputs[3721];
    assign outputs[3715] = ~((layer6_outputs[1915]) | (layer6_outputs[4312]));
    assign outputs[3716] = (layer6_outputs[977]) ^ (layer6_outputs[4760]);
    assign outputs[3717] = layer6_outputs[2006];
    assign outputs[3718] = (layer6_outputs[424]) & ~(layer6_outputs[662]);
    assign outputs[3719] = ~(layer6_outputs[2210]);
    assign outputs[3720] = layer6_outputs[1645];
    assign outputs[3721] = ~(layer6_outputs[2720]);
    assign outputs[3722] = ~(layer6_outputs[1184]);
    assign outputs[3723] = ~((layer6_outputs[2430]) | (layer6_outputs[736]));
    assign outputs[3724] = layer6_outputs[782];
    assign outputs[3725] = layer6_outputs[1121];
    assign outputs[3726] = (layer6_outputs[1369]) & ~(layer6_outputs[3030]);
    assign outputs[3727] = layer6_outputs[3897];
    assign outputs[3728] = layer6_outputs[3039];
    assign outputs[3729] = layer6_outputs[807];
    assign outputs[3730] = (layer6_outputs[3437]) & ~(layer6_outputs[1515]);
    assign outputs[3731] = ~(layer6_outputs[1884]);
    assign outputs[3732] = ~((layer6_outputs[3034]) | (layer6_outputs[1222]));
    assign outputs[3733] = ~(layer6_outputs[4548]);
    assign outputs[3734] = ~(layer6_outputs[3323]);
    assign outputs[3735] = (layer6_outputs[4423]) ^ (layer6_outputs[719]);
    assign outputs[3736] = layer6_outputs[2886];
    assign outputs[3737] = (layer6_outputs[833]) & (layer6_outputs[2255]);
    assign outputs[3738] = ~(layer6_outputs[4673]);
    assign outputs[3739] = ~(layer6_outputs[2223]);
    assign outputs[3740] = ~(layer6_outputs[4650]);
    assign outputs[3741] = layer6_outputs[382];
    assign outputs[3742] = layer6_outputs[648];
    assign outputs[3743] = ~(layer6_outputs[2066]);
    assign outputs[3744] = layer6_outputs[4573];
    assign outputs[3745] = (layer6_outputs[1168]) & ~(layer6_outputs[3123]);
    assign outputs[3746] = ~(layer6_outputs[2290]);
    assign outputs[3747] = ~((layer6_outputs[3734]) & (layer6_outputs[680]));
    assign outputs[3748] = ~(layer6_outputs[1995]);
    assign outputs[3749] = layer6_outputs[2668];
    assign outputs[3750] = layer6_outputs[3833];
    assign outputs[3751] = ~(layer6_outputs[1832]);
    assign outputs[3752] = layer6_outputs[3872];
    assign outputs[3753] = layer6_outputs[4311];
    assign outputs[3754] = (layer6_outputs[3827]) & (layer6_outputs[2157]);
    assign outputs[3755] = layer6_outputs[4238];
    assign outputs[3756] = ~(layer6_outputs[3951]);
    assign outputs[3757] = (layer6_outputs[3670]) ^ (layer6_outputs[1192]);
    assign outputs[3758] = (layer6_outputs[4561]) & ~(layer6_outputs[4392]);
    assign outputs[3759] = ~(layer6_outputs[2145]);
    assign outputs[3760] = layer6_outputs[4670];
    assign outputs[3761] = layer6_outputs[4341];
    assign outputs[3762] = (layer6_outputs[2913]) & ~(layer6_outputs[2322]);
    assign outputs[3763] = (layer6_outputs[3123]) ^ (layer6_outputs[4786]);
    assign outputs[3764] = ~(layer6_outputs[0]);
    assign outputs[3765] = (layer6_outputs[3550]) & ~(layer6_outputs[4968]);
    assign outputs[3766] = ~(layer6_outputs[988]);
    assign outputs[3767] = (layer6_outputs[2408]) & ~(layer6_outputs[2098]);
    assign outputs[3768] = (layer6_outputs[4078]) & ~(layer6_outputs[2410]);
    assign outputs[3769] = (layer6_outputs[2916]) ^ (layer6_outputs[3026]);
    assign outputs[3770] = layer6_outputs[702];
    assign outputs[3771] = ~(layer6_outputs[1745]);
    assign outputs[3772] = ~(layer6_outputs[367]);
    assign outputs[3773] = ~((layer6_outputs[2112]) | (layer6_outputs[426]));
    assign outputs[3774] = ~(layer6_outputs[2478]);
    assign outputs[3775] = (layer6_outputs[4054]) ^ (layer6_outputs[5088]);
    assign outputs[3776] = (layer6_outputs[1970]) & ~(layer6_outputs[2861]);
    assign outputs[3777] = layer6_outputs[4902];
    assign outputs[3778] = layer6_outputs[416];
    assign outputs[3779] = ~((layer6_outputs[50]) & (layer6_outputs[3310]));
    assign outputs[3780] = ~(layer6_outputs[2803]);
    assign outputs[3781] = layer6_outputs[991];
    assign outputs[3782] = ~(layer6_outputs[3108]);
    assign outputs[3783] = ~(layer6_outputs[3511]);
    assign outputs[3784] = (layer6_outputs[4614]) & (layer6_outputs[5059]);
    assign outputs[3785] = ~(layer6_outputs[2729]);
    assign outputs[3786] = ~((layer6_outputs[939]) & (layer6_outputs[3036]));
    assign outputs[3787] = layer6_outputs[905];
    assign outputs[3788] = layer6_outputs[4374];
    assign outputs[3789] = ~(layer6_outputs[4787]);
    assign outputs[3790] = (layer6_outputs[2875]) & (layer6_outputs[1081]);
    assign outputs[3791] = ~(layer6_outputs[2982]);
    assign outputs[3792] = ~(layer6_outputs[2558]) | (layer6_outputs[3111]);
    assign outputs[3793] = ~(layer6_outputs[4332]);
    assign outputs[3794] = ~(layer6_outputs[1439]);
    assign outputs[3795] = (layer6_outputs[1611]) & ~(layer6_outputs[4926]);
    assign outputs[3796] = ~((layer6_outputs[2792]) ^ (layer6_outputs[4582]));
    assign outputs[3797] = layer6_outputs[4955];
    assign outputs[3798] = (layer6_outputs[630]) ^ (layer6_outputs[1175]);
    assign outputs[3799] = layer6_outputs[3536];
    assign outputs[3800] = ~(layer6_outputs[1969]);
    assign outputs[3801] = ~((layer6_outputs[482]) ^ (layer6_outputs[2004]));
    assign outputs[3802] = (layer6_outputs[1706]) & ~(layer6_outputs[4791]);
    assign outputs[3803] = ~(layer6_outputs[1324]);
    assign outputs[3804] = (layer6_outputs[1826]) & ~(layer6_outputs[4971]);
    assign outputs[3805] = ~(layer6_outputs[2321]);
    assign outputs[3806] = ~(layer6_outputs[3230]);
    assign outputs[3807] = layer6_outputs[494];
    assign outputs[3808] = (layer6_outputs[2588]) | (layer6_outputs[827]);
    assign outputs[3809] = ~(layer6_outputs[3791]);
    assign outputs[3810] = layer6_outputs[879];
    assign outputs[3811] = ~((layer6_outputs[528]) ^ (layer6_outputs[541]));
    assign outputs[3812] = ~(layer6_outputs[4056]);
    assign outputs[3813] = ~(layer6_outputs[4823]);
    assign outputs[3814] = layer6_outputs[2144];
    assign outputs[3815] = layer6_outputs[694];
    assign outputs[3816] = ~(layer6_outputs[3168]) | (layer6_outputs[3254]);
    assign outputs[3817] = ~(layer6_outputs[3853]) | (layer6_outputs[4264]);
    assign outputs[3818] = ~((layer6_outputs[3622]) ^ (layer6_outputs[5054]));
    assign outputs[3819] = ~((layer6_outputs[1890]) ^ (layer6_outputs[929]));
    assign outputs[3820] = (layer6_outputs[3793]) ^ (layer6_outputs[4422]);
    assign outputs[3821] = layer6_outputs[1777];
    assign outputs[3822] = layer6_outputs[975];
    assign outputs[3823] = layer6_outputs[2971];
    assign outputs[3824] = layer6_outputs[2152];
    assign outputs[3825] = (layer6_outputs[4442]) & ~(layer6_outputs[3068]);
    assign outputs[3826] = (layer6_outputs[205]) & (layer6_outputs[4653]);
    assign outputs[3827] = ~(layer6_outputs[4290]);
    assign outputs[3828] = layer6_outputs[301];
    assign outputs[3829] = ~(layer6_outputs[184]);
    assign outputs[3830] = (layer6_outputs[2846]) & ~(layer6_outputs[3135]);
    assign outputs[3831] = layer6_outputs[3142];
    assign outputs[3832] = ~(layer6_outputs[2569]);
    assign outputs[3833] = layer6_outputs[3088];
    assign outputs[3834] = (layer6_outputs[1945]) ^ (layer6_outputs[2749]);
    assign outputs[3835] = ~((layer6_outputs[3740]) & (layer6_outputs[1904]));
    assign outputs[3836] = ~(layer6_outputs[939]);
    assign outputs[3837] = layer6_outputs[4861];
    assign outputs[3838] = layer6_outputs[2170];
    assign outputs[3839] = (layer6_outputs[4256]) & (layer6_outputs[3432]);
    assign outputs[3840] = ~((layer6_outputs[2168]) ^ (layer6_outputs[4672]));
    assign outputs[3841] = ~(layer6_outputs[4091]);
    assign outputs[3842] = ~(layer6_outputs[1694]);
    assign outputs[3843] = layer6_outputs[2921];
    assign outputs[3844] = layer6_outputs[3548];
    assign outputs[3845] = ~(layer6_outputs[3785]);
    assign outputs[3846] = ~(layer6_outputs[182]);
    assign outputs[3847] = (layer6_outputs[1347]) ^ (layer6_outputs[2993]);
    assign outputs[3848] = ~((layer6_outputs[1655]) ^ (layer6_outputs[4124]));
    assign outputs[3849] = layer6_outputs[4617];
    assign outputs[3850] = ~(layer6_outputs[1112]);
    assign outputs[3851] = ~(layer6_outputs[3206]);
    assign outputs[3852] = ~(layer6_outputs[1035]);
    assign outputs[3853] = layer6_outputs[1886];
    assign outputs[3854] = ~(layer6_outputs[1252]);
    assign outputs[3855] = layer6_outputs[1484];
    assign outputs[3856] = ~(layer6_outputs[3906]);
    assign outputs[3857] = ~((layer6_outputs[4688]) & (layer6_outputs[5076]));
    assign outputs[3858] = layer6_outputs[113];
    assign outputs[3859] = layer6_outputs[886];
    assign outputs[3860] = layer6_outputs[1336];
    assign outputs[3861] = (layer6_outputs[4735]) ^ (layer6_outputs[1006]);
    assign outputs[3862] = ~(layer6_outputs[1036]);
    assign outputs[3863] = ~(layer6_outputs[624]);
    assign outputs[3864] = ~(layer6_outputs[2370]);
    assign outputs[3865] = layer6_outputs[2192];
    assign outputs[3866] = ~(layer6_outputs[86]);
    assign outputs[3867] = ~(layer6_outputs[1226]) | (layer6_outputs[660]);
    assign outputs[3868] = ~(layer6_outputs[4517]) | (layer6_outputs[3414]);
    assign outputs[3869] = ~(layer6_outputs[3941]);
    assign outputs[3870] = layer6_outputs[3327];
    assign outputs[3871] = ~(layer6_outputs[3963]);
    assign outputs[3872] = ~(layer6_outputs[3158]);
    assign outputs[3873] = (layer6_outputs[1429]) | (layer6_outputs[2900]);
    assign outputs[3874] = layer6_outputs[1779];
    assign outputs[3875] = ~((layer6_outputs[2085]) ^ (layer6_outputs[2805]));
    assign outputs[3876] = ~((layer6_outputs[516]) & (layer6_outputs[2363]));
    assign outputs[3877] = layer6_outputs[3484];
    assign outputs[3878] = ~((layer6_outputs[3567]) ^ (layer6_outputs[3279]));
    assign outputs[3879] = layer6_outputs[194];
    assign outputs[3880] = layer6_outputs[970];
    assign outputs[3881] = ~(layer6_outputs[1792]);
    assign outputs[3882] = layer6_outputs[4380];
    assign outputs[3883] = layer6_outputs[3924];
    assign outputs[3884] = layer6_outputs[2405];
    assign outputs[3885] = ~(layer6_outputs[2814]);
    assign outputs[3886] = (layer6_outputs[1431]) ^ (layer6_outputs[3259]);
    assign outputs[3887] = (layer6_outputs[677]) | (layer6_outputs[343]);
    assign outputs[3888] = layer6_outputs[3488];
    assign outputs[3889] = layer6_outputs[1579];
    assign outputs[3890] = layer6_outputs[2718];
    assign outputs[3891] = layer6_outputs[3477];
    assign outputs[3892] = (layer6_outputs[5095]) ^ (layer6_outputs[3533]);
    assign outputs[3893] = ~(layer6_outputs[2704]);
    assign outputs[3894] = layer6_outputs[64];
    assign outputs[3895] = ~(layer6_outputs[1164]);
    assign outputs[3896] = (layer6_outputs[4099]) ^ (layer6_outputs[1498]);
    assign outputs[3897] = (layer6_outputs[4112]) & (layer6_outputs[1142]);
    assign outputs[3898] = layer6_outputs[650];
    assign outputs[3899] = layer6_outputs[1135];
    assign outputs[3900] = ~(layer6_outputs[4334]);
    assign outputs[3901] = ~(layer6_outputs[4893]);
    assign outputs[3902] = layer6_outputs[4439];
    assign outputs[3903] = ~(layer6_outputs[4677]);
    assign outputs[3904] = layer6_outputs[3596];
    assign outputs[3905] = ~(layer6_outputs[4296]);
    assign outputs[3906] = ~(layer6_outputs[216]);
    assign outputs[3907] = layer6_outputs[5061];
    assign outputs[3908] = layer6_outputs[2504];
    assign outputs[3909] = layer6_outputs[636];
    assign outputs[3910] = layer6_outputs[3501];
    assign outputs[3911] = layer6_outputs[3937];
    assign outputs[3912] = ~(layer6_outputs[3954]);
    assign outputs[3913] = layer6_outputs[2611];
    assign outputs[3914] = layer6_outputs[3057];
    assign outputs[3915] = ~(layer6_outputs[3140]);
    assign outputs[3916] = ~(layer6_outputs[3342]);
    assign outputs[3917] = ~(layer6_outputs[1385]);
    assign outputs[3918] = ~(layer6_outputs[3599]);
    assign outputs[3919] = ~(layer6_outputs[788]);
    assign outputs[3920] = (layer6_outputs[2421]) | (layer6_outputs[2105]);
    assign outputs[3921] = layer6_outputs[3514];
    assign outputs[3922] = layer6_outputs[5105];
    assign outputs[3923] = ~(layer6_outputs[4576]);
    assign outputs[3924] = (layer6_outputs[3258]) | (layer6_outputs[4482]);
    assign outputs[3925] = ~(layer6_outputs[3425]);
    assign outputs[3926] = layer6_outputs[2666];
    assign outputs[3927] = ~(layer6_outputs[4626]);
    assign outputs[3928] = layer6_outputs[2766];
    assign outputs[3929] = (layer6_outputs[505]) ^ (layer6_outputs[78]);
    assign outputs[3930] = (layer6_outputs[3578]) | (layer6_outputs[2847]);
    assign outputs[3931] = ~(layer6_outputs[397]);
    assign outputs[3932] = layer6_outputs[2926];
    assign outputs[3933] = (layer6_outputs[3369]) ^ (layer6_outputs[2891]);
    assign outputs[3934] = (layer6_outputs[3027]) & ~(layer6_outputs[4932]);
    assign outputs[3935] = ~(layer6_outputs[3380]);
    assign outputs[3936] = ~((layer6_outputs[5119]) ^ (layer6_outputs[1415]));
    assign outputs[3937] = layer6_outputs[2502];
    assign outputs[3938] = layer6_outputs[1714];
    assign outputs[3939] = layer6_outputs[2703];
    assign outputs[3940] = ~((layer6_outputs[1185]) ^ (layer6_outputs[1290]));
    assign outputs[3941] = layer6_outputs[3287];
    assign outputs[3942] = layer6_outputs[353];
    assign outputs[3943] = ~(layer6_outputs[823]);
    assign outputs[3944] = ~((layer6_outputs[496]) ^ (layer6_outputs[2444]));
    assign outputs[3945] = ~(layer6_outputs[495]);
    assign outputs[3946] = ~(layer6_outputs[3232]);
    assign outputs[3947] = ~(layer6_outputs[2942]);
    assign outputs[3948] = ~(layer6_outputs[4225]);
    assign outputs[3949] = (layer6_outputs[3654]) & ~(layer6_outputs[4501]);
    assign outputs[3950] = (layer6_outputs[61]) ^ (layer6_outputs[2927]);
    assign outputs[3951] = ~(layer6_outputs[3231]) | (layer6_outputs[1545]);
    assign outputs[3952] = layer6_outputs[3914];
    assign outputs[3953] = layer6_outputs[4224];
    assign outputs[3954] = ~(layer6_outputs[4898]);
    assign outputs[3955] = ~(layer6_outputs[2907]);
    assign outputs[3956] = ~(layer6_outputs[4900]);
    assign outputs[3957] = ~(layer6_outputs[490]);
    assign outputs[3958] = layer6_outputs[4292];
    assign outputs[3959] = (layer6_outputs[5028]) ^ (layer6_outputs[1509]);
    assign outputs[3960] = ~(layer6_outputs[4775]) | (layer6_outputs[791]);
    assign outputs[3961] = ~((layer6_outputs[993]) ^ (layer6_outputs[1365]));
    assign outputs[3962] = layer6_outputs[3578];
    assign outputs[3963] = ~((layer6_outputs[673]) ^ (layer6_outputs[369]));
    assign outputs[3964] = ~(layer6_outputs[1061]);
    assign outputs[3965] = ~(layer6_outputs[4868]);
    assign outputs[3966] = ~(layer6_outputs[4164]);
    assign outputs[3967] = layer6_outputs[655];
    assign outputs[3968] = ~(layer6_outputs[1451]) | (layer6_outputs[185]);
    assign outputs[3969] = layer6_outputs[4284];
    assign outputs[3970] = (layer6_outputs[4567]) & (layer6_outputs[4748]);
    assign outputs[3971] = ~(layer6_outputs[3151]);
    assign outputs[3972] = layer6_outputs[1408];
    assign outputs[3973] = ~((layer6_outputs[1174]) ^ (layer6_outputs[1864]));
    assign outputs[3974] = (layer6_outputs[3971]) ^ (layer6_outputs[2280]);
    assign outputs[3975] = ~(layer6_outputs[4735]);
    assign outputs[3976] = ~(layer6_outputs[1203]);
    assign outputs[3977] = ~(layer6_outputs[2019]);
    assign outputs[3978] = ~(layer6_outputs[3974]);
    assign outputs[3979] = ~(layer6_outputs[2007]);
    assign outputs[3980] = ~(layer6_outputs[1563]);
    assign outputs[3981] = (layer6_outputs[4566]) & (layer6_outputs[1232]);
    assign outputs[3982] = ~(layer6_outputs[334]);
    assign outputs[3983] = ~((layer6_outputs[2723]) | (layer6_outputs[4104]));
    assign outputs[3984] = ~(layer6_outputs[784]);
    assign outputs[3985] = layer6_outputs[2898];
    assign outputs[3986] = ~(layer6_outputs[3635]);
    assign outputs[3987] = layer6_outputs[4098];
    assign outputs[3988] = ~(layer6_outputs[3631]);
    assign outputs[3989] = ~(layer6_outputs[1615]);
    assign outputs[3990] = ~((layer6_outputs[4251]) | (layer6_outputs[1673]));
    assign outputs[3991] = ~(layer6_outputs[3203]);
    assign outputs[3992] = (layer6_outputs[519]) & ~(layer6_outputs[4153]);
    assign outputs[3993] = layer6_outputs[810];
    assign outputs[3994] = layer6_outputs[999];
    assign outputs[3995] = layer6_outputs[126];
    assign outputs[3996] = (layer6_outputs[746]) & (layer6_outputs[1442]);
    assign outputs[3997] = layer6_outputs[4908];
    assign outputs[3998] = ~((layer6_outputs[2084]) ^ (layer6_outputs[3640]));
    assign outputs[3999] = layer6_outputs[4881];
    assign outputs[4000] = (layer6_outputs[4132]) & (layer6_outputs[957]);
    assign outputs[4001] = layer6_outputs[3408];
    assign outputs[4002] = ~(layer6_outputs[4714]);
    assign outputs[4003] = layer6_outputs[1821];
    assign outputs[4004] = layer6_outputs[4770];
    assign outputs[4005] = ~((layer6_outputs[2442]) ^ (layer6_outputs[2839]));
    assign outputs[4006] = ~((layer6_outputs[182]) | (layer6_outputs[5086]));
    assign outputs[4007] = (layer6_outputs[2893]) ^ (layer6_outputs[4354]);
    assign outputs[4008] = ~(layer6_outputs[3818]);
    assign outputs[4009] = layer6_outputs[258];
    assign outputs[4010] = layer6_outputs[4890];
    assign outputs[4011] = ~((layer6_outputs[2398]) | (layer6_outputs[4452]));
    assign outputs[4012] = ~(layer6_outputs[4051]);
    assign outputs[4013] = ~(layer6_outputs[4279]);
    assign outputs[4014] = layer6_outputs[4746];
    assign outputs[4015] = ~(layer6_outputs[3049]);
    assign outputs[4016] = ~(layer6_outputs[1058]);
    assign outputs[4017] = layer6_outputs[2988];
    assign outputs[4018] = ~((layer6_outputs[1463]) ^ (layer6_outputs[2758]));
    assign outputs[4019] = layer6_outputs[1212];
    assign outputs[4020] = ~(layer6_outputs[2052]);
    assign outputs[4021] = (layer6_outputs[2403]) & ~(layer6_outputs[4342]);
    assign outputs[4022] = (layer6_outputs[2087]) ^ (layer6_outputs[3047]);
    assign outputs[4023] = ~((layer6_outputs[941]) ^ (layer6_outputs[4871]));
    assign outputs[4024] = ~((layer6_outputs[1764]) & (layer6_outputs[5070]));
    assign outputs[4025] = layer6_outputs[2248];
    assign outputs[4026] = ~(layer6_outputs[1285]);
    assign outputs[4027] = (layer6_outputs[889]) ^ (layer6_outputs[177]);
    assign outputs[4028] = (layer6_outputs[4001]) & ~(layer6_outputs[1353]);
    assign outputs[4029] = ~((layer6_outputs[2296]) | (layer6_outputs[4323]));
    assign outputs[4030] = ~((layer6_outputs[1518]) ^ (layer6_outputs[1858]));
    assign outputs[4031] = (layer6_outputs[32]) & (layer6_outputs[1685]);
    assign outputs[4032] = ~((layer6_outputs[154]) | (layer6_outputs[4431]));
    assign outputs[4033] = ~((layer6_outputs[3880]) ^ (layer6_outputs[2363]));
    assign outputs[4034] = layer6_outputs[2351];
    assign outputs[4035] = ~(layer6_outputs[1552]);
    assign outputs[4036] = ~(layer6_outputs[3923]);
    assign outputs[4037] = ~(layer6_outputs[392]);
    assign outputs[4038] = layer6_outputs[3937];
    assign outputs[4039] = layer6_outputs[2661];
    assign outputs[4040] = (layer6_outputs[2512]) & (layer6_outputs[4503]);
    assign outputs[4041] = ~(layer6_outputs[4818]);
    assign outputs[4042] = ~(layer6_outputs[1242]);
    assign outputs[4043] = ~(layer6_outputs[2746]);
    assign outputs[4044] = ~(layer6_outputs[4970]);
    assign outputs[4045] = (layer6_outputs[4555]) ^ (layer6_outputs[561]);
    assign outputs[4046] = ~(layer6_outputs[613]);
    assign outputs[4047] = (layer6_outputs[981]) & ~(layer6_outputs[2229]);
    assign outputs[4048] = ~(layer6_outputs[2169]);
    assign outputs[4049] = layer6_outputs[1128];
    assign outputs[4050] = layer6_outputs[2377];
    assign outputs[4051] = ~(layer6_outputs[2416]);
    assign outputs[4052] = layer6_outputs[2613];
    assign outputs[4053] = (layer6_outputs[2833]) | (layer6_outputs[4618]);
    assign outputs[4054] = (layer6_outputs[370]) ^ (layer6_outputs[37]);
    assign outputs[4055] = (layer6_outputs[3343]) & (layer6_outputs[2608]);
    assign outputs[4056] = ~((layer6_outputs[4745]) | (layer6_outputs[993]));
    assign outputs[4057] = layer6_outputs[5023];
    assign outputs[4058] = ~(layer6_outputs[4131]) | (layer6_outputs[1714]);
    assign outputs[4059] = ~(layer6_outputs[2288]);
    assign outputs[4060] = ~(layer6_outputs[3177]);
    assign outputs[4061] = ~(layer6_outputs[4790]);
    assign outputs[4062] = ~(layer6_outputs[390]);
    assign outputs[4063] = (layer6_outputs[2054]) & (layer6_outputs[2921]);
    assign outputs[4064] = layer6_outputs[3538];
    assign outputs[4065] = ~(layer6_outputs[1093]);
    assign outputs[4066] = layer6_outputs[3681];
    assign outputs[4067] = ~(layer6_outputs[1556]);
    assign outputs[4068] = layer6_outputs[757];
    assign outputs[4069] = ~(layer6_outputs[410]);
    assign outputs[4070] = (layer6_outputs[1270]) & ~(layer6_outputs[362]);
    assign outputs[4071] = ~(layer6_outputs[3689]);
    assign outputs[4072] = layer6_outputs[2298];
    assign outputs[4073] = ~(layer6_outputs[1253]);
    assign outputs[4074] = layer6_outputs[2110];
    assign outputs[4075] = layer6_outputs[638];
    assign outputs[4076] = (layer6_outputs[3884]) & ~(layer6_outputs[1507]);
    assign outputs[4077] = ~((layer6_outputs[1176]) ^ (layer6_outputs[3673]));
    assign outputs[4078] = layer6_outputs[2036];
    assign outputs[4079] = ~(layer6_outputs[3534]);
    assign outputs[4080] = ~((layer6_outputs[3547]) ^ (layer6_outputs[1923]));
    assign outputs[4081] = layer6_outputs[4901];
    assign outputs[4082] = (layer6_outputs[1420]) & (layer6_outputs[2369]);
    assign outputs[4083] = layer6_outputs[4394];
    assign outputs[4084] = layer6_outputs[4623];
    assign outputs[4085] = ~(layer6_outputs[2347]);
    assign outputs[4086] = layer6_outputs[1543];
    assign outputs[4087] = layer6_outputs[125];
    assign outputs[4088] = ~(layer6_outputs[4376]);
    assign outputs[4089] = layer6_outputs[2325];
    assign outputs[4090] = layer6_outputs[4024];
    assign outputs[4091] = (layer6_outputs[2691]) & ~(layer6_outputs[2969]);
    assign outputs[4092] = layer6_outputs[1900];
    assign outputs[4093] = layer6_outputs[3293];
    assign outputs[4094] = (layer6_outputs[1198]) ^ (layer6_outputs[1258]);
    assign outputs[4095] = ~(layer6_outputs[888]);
    assign outputs[4096] = ~(layer6_outputs[4187]);
    assign outputs[4097] = layer6_outputs[1526];
    assign outputs[4098] = ~(layer6_outputs[2619]);
    assign outputs[4099] = layer6_outputs[4953];
    assign outputs[4100] = ~((layer6_outputs[992]) & (layer6_outputs[3432]));
    assign outputs[4101] = (layer6_outputs[2627]) ^ (layer6_outputs[3586]);
    assign outputs[4102] = ~(layer6_outputs[5]);
    assign outputs[4103] = (layer6_outputs[439]) ^ (layer6_outputs[1132]);
    assign outputs[4104] = layer6_outputs[3103];
    assign outputs[4105] = ~(layer6_outputs[4240]) | (layer6_outputs[1987]);
    assign outputs[4106] = ~(layer6_outputs[3137]);
    assign outputs[4107] = ~(layer6_outputs[3655]) | (layer6_outputs[4215]);
    assign outputs[4108] = ~((layer6_outputs[100]) ^ (layer6_outputs[4847]));
    assign outputs[4109] = ~(layer6_outputs[4587]) | (layer6_outputs[1845]);
    assign outputs[4110] = layer6_outputs[1614];
    assign outputs[4111] = ~(layer6_outputs[1932]);
    assign outputs[4112] = ~(layer6_outputs[1068]);
    assign outputs[4113] = ~(layer6_outputs[1957]);
    assign outputs[4114] = ~(layer6_outputs[4150]);
    assign outputs[4115] = ~(layer6_outputs[4084]);
    assign outputs[4116] = (layer6_outputs[586]) ^ (layer6_outputs[3422]);
    assign outputs[4117] = layer6_outputs[1868];
    assign outputs[4118] = ~(layer6_outputs[4245]);
    assign outputs[4119] = ~((layer6_outputs[5019]) ^ (layer6_outputs[3950]));
    assign outputs[4120] = (layer6_outputs[620]) & (layer6_outputs[2648]);
    assign outputs[4121] = layer6_outputs[2572];
    assign outputs[4122] = layer6_outputs[971];
    assign outputs[4123] = layer6_outputs[5075];
    assign outputs[4124] = layer6_outputs[3915];
    assign outputs[4125] = layer6_outputs[3683];
    assign outputs[4126] = layer6_outputs[1565];
    assign outputs[4127] = layer6_outputs[2295];
    assign outputs[4128] = ~(layer6_outputs[2370]);
    assign outputs[4129] = (layer6_outputs[2536]) & ~(layer6_outputs[233]);
    assign outputs[4130] = 1'b1;
    assign outputs[4131] = ~(layer6_outputs[305]);
    assign outputs[4132] = layer6_outputs[3820];
    assign outputs[4133] = layer6_outputs[1615];
    assign outputs[4134] = (layer6_outputs[4370]) ^ (layer6_outputs[481]);
    assign outputs[4135] = layer6_outputs[3760];
    assign outputs[4136] = layer6_outputs[2821];
    assign outputs[4137] = ~(layer6_outputs[3522]);
    assign outputs[4138] = layer6_outputs[1693];
    assign outputs[4139] = layer6_outputs[566];
    assign outputs[4140] = layer6_outputs[82];
    assign outputs[4141] = ~(layer6_outputs[1453]);
    assign outputs[4142] = ~(layer6_outputs[2966]);
    assign outputs[4143] = ~((layer6_outputs[3920]) ^ (layer6_outputs[3859]));
    assign outputs[4144] = ~((layer6_outputs[3460]) ^ (layer6_outputs[3191]));
    assign outputs[4145] = (layer6_outputs[3415]) ^ (layer6_outputs[4508]);
    assign outputs[4146] = ~((layer6_outputs[3665]) ^ (layer6_outputs[337]));
    assign outputs[4147] = layer6_outputs[3625];
    assign outputs[4148] = ~(layer6_outputs[3650]);
    assign outputs[4149] = ~(layer6_outputs[1849]);
    assign outputs[4150] = ~(layer6_outputs[2954]);
    assign outputs[4151] = ~(layer6_outputs[3122]);
    assign outputs[4152] = ~(layer6_outputs[4566]) | (layer6_outputs[3843]);
    assign outputs[4153] = (layer6_outputs[1389]) & ~(layer6_outputs[1889]);
    assign outputs[4154] = ~((layer6_outputs[3614]) ^ (layer6_outputs[909]));
    assign outputs[4155] = ~(layer6_outputs[829]);
    assign outputs[4156] = ~((layer6_outputs[789]) ^ (layer6_outputs[1571]));
    assign outputs[4157] = layer6_outputs[5057];
    assign outputs[4158] = layer6_outputs[3893];
    assign outputs[4159] = ~(layer6_outputs[5079]);
    assign outputs[4160] = layer6_outputs[1620];
    assign outputs[4161] = (layer6_outputs[1472]) | (layer6_outputs[5077]);
    assign outputs[4162] = ~((layer6_outputs[142]) ^ (layer6_outputs[3518]));
    assign outputs[4163] = ~(layer6_outputs[5102]);
    assign outputs[4164] = layer6_outputs[824];
    assign outputs[4165] = ~(layer6_outputs[2539]);
    assign outputs[4166] = (layer6_outputs[2662]) ^ (layer6_outputs[2540]);
    assign outputs[4167] = ~(layer6_outputs[1285]) | (layer6_outputs[2735]);
    assign outputs[4168] = ~(layer6_outputs[5111]);
    assign outputs[4169] = (layer6_outputs[2135]) ^ (layer6_outputs[374]);
    assign outputs[4170] = ~(layer6_outputs[1376]);
    assign outputs[4171] = layer6_outputs[3829];
    assign outputs[4172] = layer6_outputs[4668];
    assign outputs[4173] = ~(layer6_outputs[5010]);
    assign outputs[4174] = ~(layer6_outputs[4192]);
    assign outputs[4175] = layer6_outputs[2281];
    assign outputs[4176] = layer6_outputs[2417];
    assign outputs[4177] = layer6_outputs[4653];
    assign outputs[4178] = layer6_outputs[2494];
    assign outputs[4179] = ~(layer6_outputs[4882]);
    assign outputs[4180] = ~(layer6_outputs[4117]);
    assign outputs[4181] = layer6_outputs[1749];
    assign outputs[4182] = ~(layer6_outputs[642]);
    assign outputs[4183] = ~((layer6_outputs[692]) ^ (layer6_outputs[2976]));
    assign outputs[4184] = ~(layer6_outputs[1908]) | (layer6_outputs[378]);
    assign outputs[4185] = ~((layer6_outputs[272]) & (layer6_outputs[3393]));
    assign outputs[4186] = layer6_outputs[3800];
    assign outputs[4187] = (layer6_outputs[275]) | (layer6_outputs[3730]);
    assign outputs[4188] = (layer6_outputs[3671]) ^ (layer6_outputs[2612]);
    assign outputs[4189] = layer6_outputs[4023];
    assign outputs[4190] = layer6_outputs[2572];
    assign outputs[4191] = layer6_outputs[4863];
    assign outputs[4192] = ~((layer6_outputs[3395]) ^ (layer6_outputs[1976]));
    assign outputs[4193] = (layer6_outputs[2889]) ^ (layer6_outputs[4830]);
    assign outputs[4194] = layer6_outputs[1848];
    assign outputs[4195] = 1'b0;
    assign outputs[4196] = layer6_outputs[2870];
    assign outputs[4197] = (layer6_outputs[1516]) ^ (layer6_outputs[1892]);
    assign outputs[4198] = layer6_outputs[1632];
    assign outputs[4199] = ~((layer6_outputs[4398]) ^ (layer6_outputs[2792]));
    assign outputs[4200] = ~(layer6_outputs[2378]);
    assign outputs[4201] = ~((layer6_outputs[4284]) ^ (layer6_outputs[843]));
    assign outputs[4202] = layer6_outputs[1997];
    assign outputs[4203] = layer6_outputs[210];
    assign outputs[4204] = ~(layer6_outputs[2305]);
    assign outputs[4205] = ~((layer6_outputs[3482]) & (layer6_outputs[2233]));
    assign outputs[4206] = (layer6_outputs[3481]) ^ (layer6_outputs[1499]);
    assign outputs[4207] = ~(layer6_outputs[1014]);
    assign outputs[4208] = ~(layer6_outputs[2188]) | (layer6_outputs[2574]);
    assign outputs[4209] = ~(layer6_outputs[3240]);
    assign outputs[4210] = ~((layer6_outputs[223]) | (layer6_outputs[5107]));
    assign outputs[4211] = layer6_outputs[4162];
    assign outputs[4212] = ~(layer6_outputs[2885]);
    assign outputs[4213] = ~(layer6_outputs[1177]);
    assign outputs[4214] = ~(layer6_outputs[1880]);
    assign outputs[4215] = ~(layer6_outputs[2259]) | (layer6_outputs[2452]);
    assign outputs[4216] = layer6_outputs[4371];
    assign outputs[4217] = ~(layer6_outputs[522]);
    assign outputs[4218] = (layer6_outputs[3927]) | (layer6_outputs[551]);
    assign outputs[4219] = (layer6_outputs[1051]) & (layer6_outputs[3741]);
    assign outputs[4220] = layer6_outputs[94];
    assign outputs[4221] = layer6_outputs[4781];
    assign outputs[4222] = ~(layer6_outputs[4817]);
    assign outputs[4223] = ~(layer6_outputs[1183]);
    assign outputs[4224] = ~(layer6_outputs[2360]) | (layer6_outputs[2842]);
    assign outputs[4225] = ~(layer6_outputs[443]);
    assign outputs[4226] = layer6_outputs[1275];
    assign outputs[4227] = ~((layer6_outputs[1235]) ^ (layer6_outputs[2807]));
    assign outputs[4228] = ~(layer6_outputs[1300]);
    assign outputs[4229] = ~((layer6_outputs[1500]) ^ (layer6_outputs[248]));
    assign outputs[4230] = layer6_outputs[3286];
    assign outputs[4231] = layer6_outputs[3608];
    assign outputs[4232] = layer6_outputs[1209];
    assign outputs[4233] = layer6_outputs[1875];
    assign outputs[4234] = ~((layer6_outputs[2818]) ^ (layer6_outputs[2208]));
    assign outputs[4235] = (layer6_outputs[1295]) ^ (layer6_outputs[579]);
    assign outputs[4236] = ~((layer6_outputs[1250]) ^ (layer6_outputs[785]));
    assign outputs[4237] = layer6_outputs[1767];
    assign outputs[4238] = ~(layer6_outputs[3121]);
    assign outputs[4239] = layer6_outputs[3887];
    assign outputs[4240] = ~(layer6_outputs[2626]);
    assign outputs[4241] = ~(layer6_outputs[3921]);
    assign outputs[4242] = ~(layer6_outputs[2228]);
    assign outputs[4243] = ~((layer6_outputs[2988]) ^ (layer6_outputs[1249]));
    assign outputs[4244] = (layer6_outputs[3574]) & ~(layer6_outputs[1341]);
    assign outputs[4245] = ~((layer6_outputs[3238]) ^ (layer6_outputs[569]));
    assign outputs[4246] = ~(layer6_outputs[3240]);
    assign outputs[4247] = layer6_outputs[3399];
    assign outputs[4248] = ~((layer6_outputs[3067]) ^ (layer6_outputs[1633]));
    assign outputs[4249] = (layer6_outputs[1475]) & ~(layer6_outputs[2868]);
    assign outputs[4250] = ~(layer6_outputs[879]);
    assign outputs[4251] = ~(layer6_outputs[1570]);
    assign outputs[4252] = (layer6_outputs[1205]) ^ (layer6_outputs[644]);
    assign outputs[4253] = layer6_outputs[4125];
    assign outputs[4254] = layer6_outputs[2651];
    assign outputs[4255] = layer6_outputs[3917];
    assign outputs[4256] = ~(layer6_outputs[1834]);
    assign outputs[4257] = (layer6_outputs[2991]) ^ (layer6_outputs[781]);
    assign outputs[4258] = (layer6_outputs[889]) ^ (layer6_outputs[2942]);
    assign outputs[4259] = ~((layer6_outputs[4419]) ^ (layer6_outputs[4496]));
    assign outputs[4260] = ~((layer6_outputs[3224]) & (layer6_outputs[1559]));
    assign outputs[4261] = (layer6_outputs[2545]) ^ (layer6_outputs[893]);
    assign outputs[4262] = layer6_outputs[4206];
    assign outputs[4263] = layer6_outputs[3163];
    assign outputs[4264] = layer6_outputs[4535];
    assign outputs[4265] = layer6_outputs[606];
    assign outputs[4266] = ~(layer6_outputs[3360]);
    assign outputs[4267] = ~(layer6_outputs[4890]);
    assign outputs[4268] = layer6_outputs[3736];
    assign outputs[4269] = (layer6_outputs[3062]) ^ (layer6_outputs[1781]);
    assign outputs[4270] = ~((layer6_outputs[1349]) | (layer6_outputs[4888]));
    assign outputs[4271] = layer6_outputs[931];
    assign outputs[4272] = (layer6_outputs[2648]) & (layer6_outputs[626]);
    assign outputs[4273] = ~((layer6_outputs[1751]) & (layer6_outputs[2549]));
    assign outputs[4274] = ~(layer6_outputs[2300]);
    assign outputs[4275] = ~(layer6_outputs[4706]);
    assign outputs[4276] = layer6_outputs[1676];
    assign outputs[4277] = layer6_outputs[3719];
    assign outputs[4278] = (layer6_outputs[2560]) ^ (layer6_outputs[4880]);
    assign outputs[4279] = layer6_outputs[156];
    assign outputs[4280] = (layer6_outputs[2320]) ^ (layer6_outputs[1110]);
    assign outputs[4281] = (layer6_outputs[4324]) & ~(layer6_outputs[2118]);
    assign outputs[4282] = ~(layer6_outputs[3209]);
    assign outputs[4283] = ~((layer6_outputs[4161]) & (layer6_outputs[2984]));
    assign outputs[4284] = layer6_outputs[3105];
    assign outputs[4285] = layer6_outputs[1681];
    assign outputs[4286] = ~(layer6_outputs[3646]);
    assign outputs[4287] = layer6_outputs[63];
    assign outputs[4288] = layer6_outputs[3133];
    assign outputs[4289] = ~(layer6_outputs[3128]) | (layer6_outputs[474]);
    assign outputs[4290] = ~((layer6_outputs[1933]) ^ (layer6_outputs[1722]));
    assign outputs[4291] = layer6_outputs[3903];
    assign outputs[4292] = ~(layer6_outputs[2864]);
    assign outputs[4293] = ~((layer6_outputs[2630]) ^ (layer6_outputs[4209]));
    assign outputs[4294] = layer6_outputs[3330];
    assign outputs[4295] = (layer6_outputs[4178]) ^ (layer6_outputs[1587]);
    assign outputs[4296] = layer6_outputs[4685];
    assign outputs[4297] = layer6_outputs[607];
    assign outputs[4298] = (layer6_outputs[4700]) ^ (layer6_outputs[2799]);
    assign outputs[4299] = ~(layer6_outputs[2229]);
    assign outputs[4300] = ~(layer6_outputs[4348]);
    assign outputs[4301] = ~(layer6_outputs[4731]);
    assign outputs[4302] = ~((layer6_outputs[256]) & (layer6_outputs[4889]));
    assign outputs[4303] = ~(layer6_outputs[2159]);
    assign outputs[4304] = ~(layer6_outputs[4474]);
    assign outputs[4305] = layer6_outputs[3070];
    assign outputs[4306] = ~(layer6_outputs[1120]);
    assign outputs[4307] = layer6_outputs[1086];
    assign outputs[4308] = ~(layer6_outputs[2189]);
    assign outputs[4309] = (layer6_outputs[160]) ^ (layer6_outputs[3180]);
    assign outputs[4310] = ~(layer6_outputs[2652]);
    assign outputs[4311] = layer6_outputs[1806];
    assign outputs[4312] = ~(layer6_outputs[4937]);
    assign outputs[4313] = layer6_outputs[3436];
    assign outputs[4314] = ~((layer6_outputs[3702]) & (layer6_outputs[1535]));
    assign outputs[4315] = layer6_outputs[3766];
    assign outputs[4316] = ~((layer6_outputs[4788]) ^ (layer6_outputs[2162]));
    assign outputs[4317] = ~((layer6_outputs[77]) ^ (layer6_outputs[1585]));
    assign outputs[4318] = ~((layer6_outputs[3870]) & (layer6_outputs[4551]));
    assign outputs[4319] = ~((layer6_outputs[4176]) ^ (layer6_outputs[2377]));
    assign outputs[4320] = layer6_outputs[1879];
    assign outputs[4321] = ~((layer6_outputs[2031]) ^ (layer6_outputs[1406]));
    assign outputs[4322] = layer6_outputs[3244];
    assign outputs[4323] = ~(layer6_outputs[1337]);
    assign outputs[4324] = (layer6_outputs[4246]) | (layer6_outputs[4008]);
    assign outputs[4325] = ~(layer6_outputs[114]) | (layer6_outputs[1758]);
    assign outputs[4326] = ~(layer6_outputs[1071]);
    assign outputs[4327] = ~(layer6_outputs[1622]);
    assign outputs[4328] = layer6_outputs[3636];
    assign outputs[4329] = (layer6_outputs[1836]) | (layer6_outputs[98]);
    assign outputs[4330] = ~((layer6_outputs[120]) ^ (layer6_outputs[1837]));
    assign outputs[4331] = ~(layer6_outputs[499]);
    assign outputs[4332] = layer6_outputs[4417];
    assign outputs[4333] = ~(layer6_outputs[2378]);
    assign outputs[4334] = ~(layer6_outputs[2800]);
    assign outputs[4335] = ~(layer6_outputs[2613]);
    assign outputs[4336] = (layer6_outputs[1551]) ^ (layer6_outputs[2279]);
    assign outputs[4337] = (layer6_outputs[1228]) & ~(layer6_outputs[741]);
    assign outputs[4338] = layer6_outputs[3475];
    assign outputs[4339] = ~(layer6_outputs[4767]);
    assign outputs[4340] = layer6_outputs[119];
    assign outputs[4341] = (layer6_outputs[4355]) ^ (layer6_outputs[178]);
    assign outputs[4342] = (layer6_outputs[2728]) & ~(layer6_outputs[1496]);
    assign outputs[4343] = layer6_outputs[2687];
    assign outputs[4344] = layer6_outputs[4289];
    assign outputs[4345] = layer6_outputs[2981];
    assign outputs[4346] = ~(layer6_outputs[982]);
    assign outputs[4347] = (layer6_outputs[222]) ^ (layer6_outputs[397]);
    assign outputs[4348] = ~(layer6_outputs[2835]);
    assign outputs[4349] = (layer6_outputs[646]) ^ (layer6_outputs[4715]);
    assign outputs[4350] = layer6_outputs[3231];
    assign outputs[4351] = ~(layer6_outputs[1718]);
    assign outputs[4352] = ~(layer6_outputs[766]);
    assign outputs[4353] = (layer6_outputs[2021]) & ~(layer6_outputs[3011]);
    assign outputs[4354] = ~((layer6_outputs[4778]) ^ (layer6_outputs[2968]));
    assign outputs[4355] = layer6_outputs[4689];
    assign outputs[4356] = ~(layer6_outputs[914]);
    assign outputs[4357] = ~(layer6_outputs[97]);
    assign outputs[4358] = layer6_outputs[3625];
    assign outputs[4359] = ~((layer6_outputs[2617]) ^ (layer6_outputs[576]));
    assign outputs[4360] = ~(layer6_outputs[2163]);
    assign outputs[4361] = ~((layer6_outputs[1971]) ^ (layer6_outputs[4886]));
    assign outputs[4362] = ~((layer6_outputs[1651]) ^ (layer6_outputs[3555]));
    assign outputs[4363] = (layer6_outputs[4471]) | (layer6_outputs[4859]);
    assign outputs[4364] = layer6_outputs[5045];
    assign outputs[4365] = ~(layer6_outputs[1168]) | (layer6_outputs[3247]);
    assign outputs[4366] = ~(layer6_outputs[4143]);
    assign outputs[4367] = ~(layer6_outputs[2800]);
    assign outputs[4368] = ~(layer6_outputs[2619]);
    assign outputs[4369] = (layer6_outputs[2994]) ^ (layer6_outputs[756]);
    assign outputs[4370] = layer6_outputs[2604];
    assign outputs[4371] = ~(layer6_outputs[3649]);
    assign outputs[4372] = ~(layer6_outputs[4997]);
    assign outputs[4373] = (layer6_outputs[1562]) | (layer6_outputs[1030]);
    assign outputs[4374] = ~((layer6_outputs[4924]) ^ (layer6_outputs[3313]));
    assign outputs[4375] = ~(layer6_outputs[1485]);
    assign outputs[4376] = ~((layer6_outputs[2216]) ^ (layer6_outputs[1574]));
    assign outputs[4377] = ~((layer6_outputs[1136]) ^ (layer6_outputs[407]));
    assign outputs[4378] = layer6_outputs[3293];
    assign outputs[4379] = ~((layer6_outputs[1743]) ^ (layer6_outputs[195]));
    assign outputs[4380] = layer6_outputs[3404];
    assign outputs[4381] = ~((layer6_outputs[1133]) & (layer6_outputs[2580]));
    assign outputs[4382] = ~(layer6_outputs[1510]);
    assign outputs[4383] = layer6_outputs[709];
    assign outputs[4384] = layer6_outputs[2078];
    assign outputs[4385] = ~((layer6_outputs[2432]) ^ (layer6_outputs[1563]));
    assign outputs[4386] = (layer6_outputs[1272]) ^ (layer6_outputs[4961]);
    assign outputs[4387] = ~(layer6_outputs[4797]) | (layer6_outputs[960]);
    assign outputs[4388] = ~(layer6_outputs[3637]);
    assign outputs[4389] = layer6_outputs[2926];
    assign outputs[4390] = ~(layer6_outputs[300]);
    assign outputs[4391] = layer6_outputs[1781];
    assign outputs[4392] = layer6_outputs[1056];
    assign outputs[4393] = ~((layer6_outputs[2789]) ^ (layer6_outputs[736]));
    assign outputs[4394] = layer6_outputs[579];
    assign outputs[4395] = (layer6_outputs[1157]) ^ (layer6_outputs[2071]);
    assign outputs[4396] = ~(layer6_outputs[3767]);
    assign outputs[4397] = layer6_outputs[151];
    assign outputs[4398] = ~(layer6_outputs[1098]);
    assign outputs[4399] = layer6_outputs[3056];
    assign outputs[4400] = ~((layer6_outputs[4702]) ^ (layer6_outputs[2244]));
    assign outputs[4401] = layer6_outputs[3302];
    assign outputs[4402] = ~(layer6_outputs[929]);
    assign outputs[4403] = ~(layer6_outputs[891]);
    assign outputs[4404] = ~((layer6_outputs[1553]) ^ (layer6_outputs[4642]));
    assign outputs[4405] = (layer6_outputs[2705]) | (layer6_outputs[1592]);
    assign outputs[4406] = layer6_outputs[6];
    assign outputs[4407] = (layer6_outputs[5043]) ^ (layer6_outputs[2015]);
    assign outputs[4408] = ~(layer6_outputs[4234]);
    assign outputs[4409] = ~(layer6_outputs[733]);
    assign outputs[4410] = layer6_outputs[1124];
    assign outputs[4411] = layer6_outputs[3870];
    assign outputs[4412] = layer6_outputs[3642];
    assign outputs[4413] = ~((layer6_outputs[3439]) | (layer6_outputs[4891]));
    assign outputs[4414] = ~(layer6_outputs[4084]);
    assign outputs[4415] = ~(layer6_outputs[5046]);
    assign outputs[4416] = (layer6_outputs[1000]) ^ (layer6_outputs[877]);
    assign outputs[4417] = layer6_outputs[2761];
    assign outputs[4418] = ~((layer6_outputs[1384]) ^ (layer6_outputs[2438]));
    assign outputs[4419] = ~((layer6_outputs[862]) ^ (layer6_outputs[1099]));
    assign outputs[4420] = (layer6_outputs[1572]) & ~(layer6_outputs[2312]);
    assign outputs[4421] = layer6_outputs[794];
    assign outputs[4422] = layer6_outputs[1465];
    assign outputs[4423] = ~((layer6_outputs[4780]) ^ (layer6_outputs[2086]));
    assign outputs[4424] = layer6_outputs[1191];
    assign outputs[4425] = ~((layer6_outputs[4019]) ^ (layer6_outputs[4252]));
    assign outputs[4426] = layer6_outputs[3595];
    assign outputs[4427] = (layer6_outputs[4166]) & ~(layer6_outputs[2089]);
    assign outputs[4428] = ~((layer6_outputs[2012]) ^ (layer6_outputs[2754]));
    assign outputs[4429] = 1'b1;
    assign outputs[4430] = (layer6_outputs[4552]) ^ (layer6_outputs[3075]);
    assign outputs[4431] = ~(layer6_outputs[4499]);
    assign outputs[4432] = ~(layer6_outputs[3462]);
    assign outputs[4433] = ~(layer6_outputs[2373]);
    assign outputs[4434] = ~(layer6_outputs[347]);
    assign outputs[4435] = ~(layer6_outputs[2874]);
    assign outputs[4436] = ~((layer6_outputs[2886]) ^ (layer6_outputs[3761]));
    assign outputs[4437] = ~(layer6_outputs[1134]);
    assign outputs[4438] = ~((layer6_outputs[2641]) ^ (layer6_outputs[2287]));
    assign outputs[4439] = ~(layer6_outputs[4578]);
    assign outputs[4440] = ~(layer6_outputs[4453]);
    assign outputs[4441] = ~(layer6_outputs[3212]) | (layer6_outputs[4306]);
    assign outputs[4442] = layer6_outputs[3718];
    assign outputs[4443] = ~(layer6_outputs[2459]);
    assign outputs[4444] = ~(layer6_outputs[4027]);
    assign outputs[4445] = layer6_outputs[876];
    assign outputs[4446] = ~(layer6_outputs[4386]);
    assign outputs[4447] = ~((layer6_outputs[3100]) & (layer6_outputs[557]));
    assign outputs[4448] = (layer6_outputs[33]) ^ (layer6_outputs[3572]);
    assign outputs[4449] = ~((layer6_outputs[3792]) ^ (layer6_outputs[5]));
    assign outputs[4450] = ~((layer6_outputs[4542]) | (layer6_outputs[2566]));
    assign outputs[4451] = layer6_outputs[4435];
    assign outputs[4452] = ~((layer6_outputs[3409]) ^ (layer6_outputs[672]));
    assign outputs[4453] = ~((layer6_outputs[683]) | (layer6_outputs[1419]));
    assign outputs[4454] = (layer6_outputs[340]) | (layer6_outputs[2561]);
    assign outputs[4455] = ~((layer6_outputs[3549]) & (layer6_outputs[4560]));
    assign outputs[4456] = ~(layer6_outputs[1766]);
    assign outputs[4457] = (layer6_outputs[784]) ^ (layer6_outputs[2003]);
    assign outputs[4458] = ~(layer6_outputs[3042]);
    assign outputs[4459] = (layer6_outputs[3259]) ^ (layer6_outputs[4665]);
    assign outputs[4460] = layer6_outputs[1195];
    assign outputs[4461] = layer6_outputs[3930];
    assign outputs[4462] = layer6_outputs[2842];
    assign outputs[4463] = layer6_outputs[3028];
    assign outputs[4464] = ~((layer6_outputs[1381]) ^ (layer6_outputs[2529]));
    assign outputs[4465] = ~((layer6_outputs[3118]) ^ (layer6_outputs[934]));
    assign outputs[4466] = ~(layer6_outputs[4792]);
    assign outputs[4467] = ~(layer6_outputs[3093]);
    assign outputs[4468] = ~(layer6_outputs[3365]);
    assign outputs[4469] = layer6_outputs[1166];
    assign outputs[4470] = layer6_outputs[1818];
    assign outputs[4471] = (layer6_outputs[510]) ^ (layer6_outputs[1800]);
    assign outputs[4472] = layer6_outputs[926];
    assign outputs[4473] = (layer6_outputs[4508]) | (layer6_outputs[4069]);
    assign outputs[4474] = ~(layer6_outputs[3966]);
    assign outputs[4475] = ~(layer6_outputs[546]);
    assign outputs[4476] = layer6_outputs[302];
    assign outputs[4477] = (layer6_outputs[2176]) ^ (layer6_outputs[4157]);
    assign outputs[4478] = layer6_outputs[3058];
    assign outputs[4479] = (layer6_outputs[1070]) ^ (layer6_outputs[2083]);
    assign outputs[4480] = (layer6_outputs[4045]) | (layer6_outputs[552]);
    assign outputs[4481] = layer6_outputs[4243];
    assign outputs[4482] = ~((layer6_outputs[5038]) & (layer6_outputs[4470]));
    assign outputs[4483] = ~(layer6_outputs[1505]);
    assign outputs[4484] = (layer6_outputs[1703]) ^ (layer6_outputs[2928]);
    assign outputs[4485] = ~((layer6_outputs[1608]) ^ (layer6_outputs[4692]));
    assign outputs[4486] = layer6_outputs[4090];
    assign outputs[4487] = ~(layer6_outputs[945]) | (layer6_outputs[4918]);
    assign outputs[4488] = layer6_outputs[2947];
    assign outputs[4489] = ~(layer6_outputs[2068]);
    assign outputs[4490] = ~(layer6_outputs[2871]);
    assign outputs[4491] = layer6_outputs[1893];
    assign outputs[4492] = ~(layer6_outputs[3925]);
    assign outputs[4493] = ~((layer6_outputs[3018]) ^ (layer6_outputs[3453]));
    assign outputs[4494] = ~((layer6_outputs[1491]) ^ (layer6_outputs[5116]));
    assign outputs[4495] = ~(layer6_outputs[3764]);
    assign outputs[4496] = ~(layer6_outputs[818]);
    assign outputs[4497] = layer6_outputs[2745];
    assign outputs[4498] = layer6_outputs[3085];
    assign outputs[4499] = ~(layer6_outputs[1869]);
    assign outputs[4500] = (layer6_outputs[2979]) & ~(layer6_outputs[202]);
    assign outputs[4501] = ~(layer6_outputs[4549]) | (layer6_outputs[2968]);
    assign outputs[4502] = (layer6_outputs[2471]) & (layer6_outputs[4822]);
    assign outputs[4503] = layer6_outputs[2558];
    assign outputs[4504] = ~(layer6_outputs[3722]);
    assign outputs[4505] = (layer6_outputs[4174]) & ~(layer6_outputs[1750]);
    assign outputs[4506] = layer6_outputs[587];
    assign outputs[4507] = (layer6_outputs[3192]) ^ (layer6_outputs[3341]);
    assign outputs[4508] = ~(layer6_outputs[537]) | (layer6_outputs[1987]);
    assign outputs[4509] = ~(layer6_outputs[2153]) | (layer6_outputs[1249]);
    assign outputs[4510] = ~(layer6_outputs[1498]);
    assign outputs[4511] = layer6_outputs[3932];
    assign outputs[4512] = ~(layer6_outputs[1126]);
    assign outputs[4513] = ~(layer6_outputs[4486]) | (layer6_outputs[710]);
    assign outputs[4514] = layer6_outputs[4526];
    assign outputs[4515] = layer6_outputs[2612];
    assign outputs[4516] = 1'b1;
    assign outputs[4517] = layer6_outputs[2107];
    assign outputs[4518] = ~(layer6_outputs[329]);
    assign outputs[4519] = (layer6_outputs[536]) ^ (layer6_outputs[3480]);
    assign outputs[4520] = ~(layer6_outputs[3129]) | (layer6_outputs[358]);
    assign outputs[4521] = (layer6_outputs[2232]) ^ (layer6_outputs[2388]);
    assign outputs[4522] = ~(layer6_outputs[5004]);
    assign outputs[4523] = layer6_outputs[2636];
    assign outputs[4524] = layer6_outputs[2527];
    assign outputs[4525] = layer6_outputs[4241];
    assign outputs[4526] = ~((layer6_outputs[1713]) ^ (layer6_outputs[2812]));
    assign outputs[4527] = layer6_outputs[520];
    assign outputs[4528] = ~(layer6_outputs[764]);
    assign outputs[4529] = layer6_outputs[4160];
    assign outputs[4530] = layer6_outputs[3478];
    assign outputs[4531] = ~(layer6_outputs[2293]);
    assign outputs[4532] = ~(layer6_outputs[2110]);
    assign outputs[4533] = (layer6_outputs[2809]) ^ (layer6_outputs[395]);
    assign outputs[4534] = ~((layer6_outputs[555]) & (layer6_outputs[3677]));
    assign outputs[4535] = ~(layer6_outputs[2405]) | (layer6_outputs[276]);
    assign outputs[4536] = ~(layer6_outputs[1122]);
    assign outputs[4537] = layer6_outputs[1044];
    assign outputs[4538] = layer6_outputs[1404];
    assign outputs[4539] = 1'b1;
    assign outputs[4540] = layer6_outputs[3456];
    assign outputs[4541] = layer6_outputs[4495];
    assign outputs[4542] = ~(layer6_outputs[3460]);
    assign outputs[4543] = ~(layer6_outputs[298]) | (layer6_outputs[3484]);
    assign outputs[4544] = ~(layer6_outputs[384]);
    assign outputs[4545] = layer6_outputs[2193];
    assign outputs[4546] = ~(layer6_outputs[1410]);
    assign outputs[4547] = ~((layer6_outputs[1885]) & (layer6_outputs[3041]));
    assign outputs[4548] = layer6_outputs[1257];
    assign outputs[4549] = layer6_outputs[265];
    assign outputs[4550] = layer6_outputs[4459];
    assign outputs[4551] = ~(layer6_outputs[839]);
    assign outputs[4552] = ~(layer6_outputs[1618]);
    assign outputs[4553] = ~((layer6_outputs[1744]) & (layer6_outputs[4579]));
    assign outputs[4554] = ~(layer6_outputs[4375]);
    assign outputs[4555] = layer6_outputs[4369];
    assign outputs[4556] = layer6_outputs[4512];
    assign outputs[4557] = layer6_outputs[2316];
    assign outputs[4558] = layer6_outputs[1291];
    assign outputs[4559] = layer6_outputs[1739];
    assign outputs[4560] = ~((layer6_outputs[4107]) ^ (layer6_outputs[1407]));
    assign outputs[4561] = ~((layer6_outputs[3139]) ^ (layer6_outputs[349]));
    assign outputs[4562] = (layer6_outputs[4788]) ^ (layer6_outputs[2375]);
    assign outputs[4563] = ~(layer6_outputs[3576]);
    assign outputs[4564] = layer6_outputs[4790];
    assign outputs[4565] = layer6_outputs[3327];
    assign outputs[4566] = ~(layer6_outputs[405]);
    assign outputs[4567] = ~(layer6_outputs[3609]) | (layer6_outputs[391]);
    assign outputs[4568] = ~(layer6_outputs[329]);
    assign outputs[4569] = ~(layer6_outputs[3202]);
    assign outputs[4570] = layer6_outputs[2480];
    assign outputs[4571] = layer6_outputs[270];
    assign outputs[4572] = layer6_outputs[2819];
    assign outputs[4573] = ~(layer6_outputs[2944]) | (layer6_outputs[3434]);
    assign outputs[4574] = layer6_outputs[2236];
    assign outputs[4575] = ~((layer6_outputs[1479]) | (layer6_outputs[3235]));
    assign outputs[4576] = ~(layer6_outputs[1268]);
    assign outputs[4577] = (layer6_outputs[5036]) & ~(layer6_outputs[4113]);
    assign outputs[4578] = (layer6_outputs[692]) ^ (layer6_outputs[3336]);
    assign outputs[4579] = ~(layer6_outputs[1017]);
    assign outputs[4580] = (layer6_outputs[706]) ^ (layer6_outputs[5083]);
    assign outputs[4581] = layer6_outputs[7];
    assign outputs[4582] = ~((layer6_outputs[3406]) ^ (layer6_outputs[2215]));
    assign outputs[4583] = ~(layer6_outputs[3685]);
    assign outputs[4584] = layer6_outputs[520];
    assign outputs[4585] = layer6_outputs[4239];
    assign outputs[4586] = ~((layer6_outputs[3759]) ^ (layer6_outputs[1466]));
    assign outputs[4587] = layer6_outputs[3508];
    assign outputs[4588] = layer6_outputs[1291];
    assign outputs[4589] = ~(layer6_outputs[2682]) | (layer6_outputs[2633]);
    assign outputs[4590] = (layer6_outputs[203]) ^ (layer6_outputs[5079]);
    assign outputs[4591] = (layer6_outputs[1919]) ^ (layer6_outputs[4455]);
    assign outputs[4592] = (layer6_outputs[1638]) & ~(layer6_outputs[1815]);
    assign outputs[4593] = (layer6_outputs[2637]) ^ (layer6_outputs[488]);
    assign outputs[4594] = ~(layer6_outputs[1833]);
    assign outputs[4595] = (layer6_outputs[2385]) ^ (layer6_outputs[1543]);
    assign outputs[4596] = (layer6_outputs[1362]) & ~(layer6_outputs[1399]);
    assign outputs[4597] = (layer6_outputs[836]) | (layer6_outputs[3066]);
    assign outputs[4598] = ~(layer6_outputs[3776]);
    assign outputs[4599] = ~(layer6_outputs[2475]);
    assign outputs[4600] = ~(layer6_outputs[3337]);
    assign outputs[4601] = (layer6_outputs[3751]) ^ (layer6_outputs[777]);
    assign outputs[4602] = layer6_outputs[3570];
    assign outputs[4603] = ~(layer6_outputs[4328]);
    assign outputs[4604] = ~(layer6_outputs[1996]);
    assign outputs[4605] = ~(layer6_outputs[3978]);
    assign outputs[4606] = ~((layer6_outputs[4610]) ^ (layer6_outputs[3563]));
    assign outputs[4607] = (layer6_outputs[4515]) ^ (layer6_outputs[4522]);
    assign outputs[4608] = layer6_outputs[244];
    assign outputs[4609] = (layer6_outputs[4680]) ^ (layer6_outputs[1157]);
    assign outputs[4610] = layer6_outputs[2473];
    assign outputs[4611] = ~((layer6_outputs[65]) ^ (layer6_outputs[1835]));
    assign outputs[4612] = layer6_outputs[1628];
    assign outputs[4613] = ~(layer6_outputs[2493]);
    assign outputs[4614] = ~(layer6_outputs[4974]);
    assign outputs[4615] = layer6_outputs[112];
    assign outputs[4616] = layer6_outputs[1358];
    assign outputs[4617] = layer6_outputs[1324];
    assign outputs[4618] = ~(layer6_outputs[230]);
    assign outputs[4619] = (layer6_outputs[2814]) ^ (layer6_outputs[4786]);
    assign outputs[4620] = ~((layer6_outputs[3669]) | (layer6_outputs[1565]));
    assign outputs[4621] = ~((layer6_outputs[586]) ^ (layer6_outputs[1816]));
    assign outputs[4622] = layer6_outputs[2934];
    assign outputs[4623] = ~(layer6_outputs[3247]);
    assign outputs[4624] = (layer6_outputs[2989]) ^ (layer6_outputs[4880]);
    assign outputs[4625] = layer6_outputs[4031];
    assign outputs[4626] = layer6_outputs[1162];
    assign outputs[4627] = (layer6_outputs[201]) & ~(layer6_outputs[5015]);
    assign outputs[4628] = layer6_outputs[2923];
    assign outputs[4629] = ~(layer6_outputs[1013]) | (layer6_outputs[5066]);
    assign outputs[4630] = ~(layer6_outputs[2537]);
    assign outputs[4631] = ~(layer6_outputs[824]);
    assign outputs[4632] = layer6_outputs[3557];
    assign outputs[4633] = layer6_outputs[3061];
    assign outputs[4634] = layer6_outputs[1728];
    assign outputs[4635] = ~(layer6_outputs[3094]) | (layer6_outputs[2621]);
    assign outputs[4636] = layer6_outputs[3840];
    assign outputs[4637] = ~(layer6_outputs[3496]);
    assign outputs[4638] = (layer6_outputs[4379]) & ~(layer6_outputs[1694]);
    assign outputs[4639] = ~(layer6_outputs[2574]);
    assign outputs[4640] = layer6_outputs[1422];
    assign outputs[4641] = layer6_outputs[1551];
    assign outputs[4642] = (layer6_outputs[389]) | (layer6_outputs[3371]);
    assign outputs[4643] = layer6_outputs[3922];
    assign outputs[4644] = ~(layer6_outputs[3895]);
    assign outputs[4645] = ~(layer6_outputs[985]);
    assign outputs[4646] = layer6_outputs[3078];
    assign outputs[4647] = layer6_outputs[3658];
    assign outputs[4648] = ~((layer6_outputs[737]) ^ (layer6_outputs[4581]));
    assign outputs[4649] = layer6_outputs[2248];
    assign outputs[4650] = ~(layer6_outputs[3127]);
    assign outputs[4651] = ~(layer6_outputs[1342]);
    assign outputs[4652] = ~(layer6_outputs[2550]);
    assign outputs[4653] = layer6_outputs[3258];
    assign outputs[4654] = layer6_outputs[1364];
    assign outputs[4655] = ~(layer6_outputs[4228]);
    assign outputs[4656] = layer6_outputs[2104];
    assign outputs[4657] = layer6_outputs[2738];
    assign outputs[4658] = layer6_outputs[2];
    assign outputs[4659] = ~(layer6_outputs[1680]);
    assign outputs[4660] = ~(layer6_outputs[2294]);
    assign outputs[4661] = ~(layer6_outputs[4072]) | (layer6_outputs[3543]);
    assign outputs[4662] = layer6_outputs[4964];
    assign outputs[4663] = layer6_outputs[64];
    assign outputs[4664] = layer6_outputs[4086];
    assign outputs[4665] = ~(layer6_outputs[4236]);
    assign outputs[4666] = layer6_outputs[1200];
    assign outputs[4667] = ~(layer6_outputs[348]);
    assign outputs[4668] = (layer6_outputs[1154]) ^ (layer6_outputs[2722]);
    assign outputs[4669] = ~(layer6_outputs[3816]);
    assign outputs[4670] = (layer6_outputs[5039]) & ~(layer6_outputs[4389]);
    assign outputs[4671] = ~((layer6_outputs[4043]) & (layer6_outputs[221]));
    assign outputs[4672] = (layer6_outputs[568]) ^ (layer6_outputs[27]);
    assign outputs[4673] = layer6_outputs[1641];
    assign outputs[4674] = (layer6_outputs[3429]) | (layer6_outputs[3645]);
    assign outputs[4675] = layer6_outputs[3082];
    assign outputs[4676] = ~(layer6_outputs[1344]);
    assign outputs[4677] = layer6_outputs[4972];
    assign outputs[4678] = ~(layer6_outputs[2394]);
    assign outputs[4679] = ~(layer6_outputs[901]);
    assign outputs[4680] = layer6_outputs[3492];
    assign outputs[4681] = ~(layer6_outputs[1820]);
    assign outputs[4682] = layer6_outputs[1403];
    assign outputs[4683] = ~(layer6_outputs[4390]);
    assign outputs[4684] = (layer6_outputs[2917]) & ~(layer6_outputs[1138]);
    assign outputs[4685] = ~(layer6_outputs[55]);
    assign outputs[4686] = ~((layer6_outputs[2759]) ^ (layer6_outputs[2165]));
    assign outputs[4687] = ~((layer6_outputs[2653]) ^ (layer6_outputs[3074]));
    assign outputs[4688] = ~((layer6_outputs[4791]) | (layer6_outputs[700]));
    assign outputs[4689] = ~(layer6_outputs[3787]);
    assign outputs[4690] = ~(layer6_outputs[1653]);
    assign outputs[4691] = ~(layer6_outputs[4138]);
    assign outputs[4692] = ~((layer6_outputs[511]) ^ (layer6_outputs[1189]));
    assign outputs[4693] = ~((layer6_outputs[3308]) | (layer6_outputs[4397]));
    assign outputs[4694] = ~((layer6_outputs[1207]) ^ (layer6_outputs[1478]));
    assign outputs[4695] = (layer6_outputs[3089]) ^ (layer6_outputs[955]);
    assign outputs[4696] = layer6_outputs[4444];
    assign outputs[4697] = layer6_outputs[3122];
    assign outputs[4698] = (layer6_outputs[1931]) ^ (layer6_outputs[760]);
    assign outputs[4699] = layer6_outputs[3052];
    assign outputs[4700] = (layer6_outputs[3179]) & (layer6_outputs[1274]);
    assign outputs[4701] = (layer6_outputs[4560]) & ~(layer6_outputs[2933]);
    assign outputs[4702] = layer6_outputs[1081];
    assign outputs[4703] = layer6_outputs[129];
    assign outputs[4704] = ~((layer6_outputs[4577]) ^ (layer6_outputs[980]));
    assign outputs[4705] = (layer6_outputs[4875]) ^ (layer6_outputs[3750]);
    assign outputs[4706] = ~((layer6_outputs[2340]) | (layer6_outputs[613]));
    assign outputs[4707] = (layer6_outputs[2985]) & ~(layer6_outputs[1867]);
    assign outputs[4708] = (layer6_outputs[1041]) ^ (layer6_outputs[516]);
    assign outputs[4709] = ~(layer6_outputs[1028]);
    assign outputs[4710] = ~(layer6_outputs[3479]);
    assign outputs[4711] = layer6_outputs[57];
    assign outputs[4712] = layer6_outputs[890];
    assign outputs[4713] = ~((layer6_outputs[3062]) | (layer6_outputs[797]));
    assign outputs[4714] = ~(layer6_outputs[4829]);
    assign outputs[4715] = layer6_outputs[764];
    assign outputs[4716] = (layer6_outputs[479]) ^ (layer6_outputs[1462]);
    assign outputs[4717] = layer6_outputs[573];
    assign outputs[4718] = (layer6_outputs[1705]) & (layer6_outputs[2749]);
    assign outputs[4719] = layer6_outputs[3791];
    assign outputs[4720] = layer6_outputs[2943];
    assign outputs[4721] = ~((layer6_outputs[3632]) ^ (layer6_outputs[384]));
    assign outputs[4722] = ~(layer6_outputs[3226]);
    assign outputs[4723] = layer6_outputs[1512];
    assign outputs[4724] = layer6_outputs[3070];
    assign outputs[4725] = (layer6_outputs[189]) | (layer6_outputs[2901]);
    assign outputs[4726] = (layer6_outputs[5046]) | (layer6_outputs[2241]);
    assign outputs[4727] = ~(layer6_outputs[42]);
    assign outputs[4728] = ~(layer6_outputs[3628]);
    assign outputs[4729] = ~(layer6_outputs[45]);
    assign outputs[4730] = (layer6_outputs[3113]) ^ (layer6_outputs[1010]);
    assign outputs[4731] = layer6_outputs[2231];
    assign outputs[4732] = ~((layer6_outputs[3807]) ^ (layer6_outputs[2476]));
    assign outputs[4733] = ~(layer6_outputs[2093]);
    assign outputs[4734] = layer6_outputs[2472];
    assign outputs[4735] = (layer6_outputs[2747]) ^ (layer6_outputs[1809]);
    assign outputs[4736] = ~((layer6_outputs[1782]) ^ (layer6_outputs[451]));
    assign outputs[4737] = (layer6_outputs[4369]) ^ (layer6_outputs[3402]);
    assign outputs[4738] = ~(layer6_outputs[1308]);
    assign outputs[4739] = ~(layer6_outputs[2195]);
    assign outputs[4740] = ~(layer6_outputs[1917]);
    assign outputs[4741] = layer6_outputs[4686];
    assign outputs[4742] = ~((layer6_outputs[172]) ^ (layer6_outputs[3942]));
    assign outputs[4743] = layer6_outputs[3546];
    assign outputs[4744] = ~(layer6_outputs[2151]);
    assign outputs[4745] = ~(layer6_outputs[704]) | (layer6_outputs[2987]);
    assign outputs[4746] = ~(layer6_outputs[3145]);
    assign outputs[4747] = (layer6_outputs[3393]) & ~(layer6_outputs[3024]);
    assign outputs[4748] = ~(layer6_outputs[2869]);
    assign outputs[4749] = ~((layer6_outputs[3944]) ^ (layer6_outputs[4154]));
    assign outputs[4750] = ~(layer6_outputs[4091]);
    assign outputs[4751] = (layer6_outputs[3513]) & ~(layer6_outputs[3521]);
    assign outputs[4752] = ~(layer6_outputs[946]) | (layer6_outputs[3602]);
    assign outputs[4753] = ~(layer6_outputs[3405]);
    assign outputs[4754] = layer6_outputs[2663];
    assign outputs[4755] = ~(layer6_outputs[3066]);
    assign outputs[4756] = ~(layer6_outputs[3102]);
    assign outputs[4757] = ~(layer6_outputs[4509]);
    assign outputs[4758] = ~(layer6_outputs[4946]);
    assign outputs[4759] = layer6_outputs[1742];
    assign outputs[4760] = layer6_outputs[3639];
    assign outputs[4761] = ~((layer6_outputs[850]) ^ (layer6_outputs[3017]));
    assign outputs[4762] = ~((layer6_outputs[1083]) | (layer6_outputs[1143]));
    assign outputs[4763] = layer6_outputs[2059];
    assign outputs[4764] = ~((layer6_outputs[1491]) ^ (layer6_outputs[2256]));
    assign outputs[4765] = layer6_outputs[1581];
    assign outputs[4766] = (layer6_outputs[3281]) | (layer6_outputs[385]);
    assign outputs[4767] = (layer6_outputs[2472]) ^ (layer6_outputs[1643]);
    assign outputs[4768] = (layer6_outputs[4849]) ^ (layer6_outputs[2400]);
    assign outputs[4769] = ~(layer6_outputs[4755]);
    assign outputs[4770] = layer6_outputs[3624];
    assign outputs[4771] = ~(layer6_outputs[530]);
    assign outputs[4772] = (layer6_outputs[1657]) ^ (layer6_outputs[2511]);
    assign outputs[4773] = ~(layer6_outputs[4360]);
    assign outputs[4774] = layer6_outputs[1237];
    assign outputs[4775] = ~(layer6_outputs[3664]);
    assign outputs[4776] = ~((layer6_outputs[577]) ^ (layer6_outputs[447]));
    assign outputs[4777] = ~(layer6_outputs[2198]) | (layer6_outputs[1207]);
    assign outputs[4778] = layer6_outputs[2631];
    assign outputs[4779] = (layer6_outputs[2938]) ^ (layer6_outputs[4130]);
    assign outputs[4780] = (layer6_outputs[1382]) ^ (layer6_outputs[4763]);
    assign outputs[4781] = layer6_outputs[3492];
    assign outputs[4782] = (layer6_outputs[386]) ^ (layer6_outputs[1313]);
    assign outputs[4783] = ~(layer6_outputs[1804]);
    assign outputs[4784] = ~((layer6_outputs[2406]) ^ (layer6_outputs[4590]));
    assign outputs[4785] = layer6_outputs[3255];
    assign outputs[4786] = ~(layer6_outputs[772]);
    assign outputs[4787] = ~(layer6_outputs[1609]);
    assign outputs[4788] = (layer6_outputs[801]) & ~(layer6_outputs[415]);
    assign outputs[4789] = 1'b0;
    assign outputs[4790] = (layer6_outputs[2717]) ^ (layer6_outputs[4562]);
    assign outputs[4791] = layer6_outputs[2735];
    assign outputs[4792] = ~(layer6_outputs[1834]);
    assign outputs[4793] = ~(layer6_outputs[4141]);
    assign outputs[4794] = layer6_outputs[5000];
    assign outputs[4795] = layer6_outputs[5049];
    assign outputs[4796] = layer6_outputs[664];
    assign outputs[4797] = ~(layer6_outputs[2938]);
    assign outputs[4798] = ~(layer6_outputs[3896]);
    assign outputs[4799] = layer6_outputs[1403];
    assign outputs[4800] = (layer6_outputs[907]) ^ (layer6_outputs[1691]);
    assign outputs[4801] = layer6_outputs[3147];
    assign outputs[4802] = ~(layer6_outputs[492]);
    assign outputs[4803] = ~(layer6_outputs[2538]);
    assign outputs[4804] = ~((layer6_outputs[4527]) ^ (layer6_outputs[4808]));
    assign outputs[4805] = layer6_outputs[2586];
    assign outputs[4806] = layer6_outputs[2514];
    assign outputs[4807] = layer6_outputs[5085];
    assign outputs[4808] = (layer6_outputs[3050]) & (layer6_outputs[309]);
    assign outputs[4809] = layer6_outputs[663];
    assign outputs[4810] = layer6_outputs[2384];
    assign outputs[4811] = layer6_outputs[3572];
    assign outputs[4812] = ~(layer6_outputs[3856]);
    assign outputs[4813] = ~(layer6_outputs[4606]);
    assign outputs[4814] = ~((layer6_outputs[1047]) | (layer6_outputs[3767]));
    assign outputs[4815] = ~(layer6_outputs[919]);
    assign outputs[4816] = layer6_outputs[1630];
    assign outputs[4817] = ~(layer6_outputs[2669]);
    assign outputs[4818] = ~((layer6_outputs[2445]) & (layer6_outputs[878]));
    assign outputs[4819] = layer6_outputs[3018];
    assign outputs[4820] = ~(layer6_outputs[1857]);
    assign outputs[4821] = ~(layer6_outputs[2594]);
    assign outputs[4822] = layer6_outputs[546];
    assign outputs[4823] = ~(layer6_outputs[2873]);
    assign outputs[4824] = layer6_outputs[3165];
    assign outputs[4825] = (layer6_outputs[1334]) & (layer6_outputs[3120]);
    assign outputs[4826] = ~(layer6_outputs[1555]);
    assign outputs[4827] = layer6_outputs[527];
    assign outputs[4828] = ~((layer6_outputs[1558]) ^ (layer6_outputs[3083]));
    assign outputs[4829] = (layer6_outputs[2702]) ^ (layer6_outputs[2183]);
    assign outputs[4830] = layer6_outputs[2570];
    assign outputs[4831] = (layer6_outputs[2685]) | (layer6_outputs[805]);
    assign outputs[4832] = ~((layer6_outputs[3600]) | (layer6_outputs[5037]));
    assign outputs[4833] = (layer6_outputs[2034]) ^ (layer6_outputs[2606]);
    assign outputs[4834] = (layer6_outputs[4363]) & (layer6_outputs[5073]);
    assign outputs[4835] = ~((layer6_outputs[4925]) ^ (layer6_outputs[1243]));
    assign outputs[4836] = (layer6_outputs[707]) & ~(layer6_outputs[2018]);
    assign outputs[4837] = ~((layer6_outputs[2601]) ^ (layer6_outputs[3969]));
    assign outputs[4838] = (layer6_outputs[4638]) & ~(layer6_outputs[4903]);
    assign outputs[4839] = ~(layer6_outputs[471]);
    assign outputs[4840] = (layer6_outputs[1227]) ^ (layer6_outputs[425]);
    assign outputs[4841] = layer6_outputs[1299];
    assign outputs[4842] = layer6_outputs[3681];
    assign outputs[4843] = layer6_outputs[553];
    assign outputs[4844] = (layer6_outputs[1872]) ^ (layer6_outputs[3430]);
    assign outputs[4845] = layer6_outputs[2373];
    assign outputs[4846] = layer6_outputs[3629];
    assign outputs[4847] = layer6_outputs[4954];
    assign outputs[4848] = layer6_outputs[3503];
    assign outputs[4849] = ~((layer6_outputs[4247]) ^ (layer6_outputs[671]));
    assign outputs[4850] = ~((layer6_outputs[3981]) ^ (layer6_outputs[2506]));
    assign outputs[4851] = layer6_outputs[4926];
    assign outputs[4852] = layer6_outputs[872];
    assign outputs[4853] = ~((layer6_outputs[1044]) ^ (layer6_outputs[3053]));
    assign outputs[4854] = ~(layer6_outputs[4544]);
    assign outputs[4855] = layer6_outputs[24];
    assign outputs[4856] = layer6_outputs[4292];
    assign outputs[4857] = layer6_outputs[354];
    assign outputs[4858] = (layer6_outputs[1380]) ^ (layer6_outputs[1413]);
    assign outputs[4859] = ~((layer6_outputs[4797]) & (layer6_outputs[1182]));
    assign outputs[4860] = ~(layer6_outputs[860]);
    assign outputs[4861] = ~(layer6_outputs[2799]);
    assign outputs[4862] = ~(layer6_outputs[1955]);
    assign outputs[4863] = ~((layer6_outputs[608]) ^ (layer6_outputs[2542]));
    assign outputs[4864] = ~(layer6_outputs[1264]);
    assign outputs[4865] = layer6_outputs[3910];
    assign outputs[4866] = ~(layer6_outputs[3287]);
    assign outputs[4867] = ~(layer6_outputs[3607]) | (layer6_outputs[2154]);
    assign outputs[4868] = (layer6_outputs[2897]) ^ (layer6_outputs[4935]);
    assign outputs[4869] = (layer6_outputs[2178]) & ~(layer6_outputs[1083]);
    assign outputs[4870] = layer6_outputs[3140];
    assign outputs[4871] = ~(layer6_outputs[3248]);
    assign outputs[4872] = ~((layer6_outputs[493]) ^ (layer6_outputs[3086]));
    assign outputs[4873] = layer6_outputs[297];
    assign outputs[4874] = (layer6_outputs[3871]) & ~(layer6_outputs[3363]);
    assign outputs[4875] = ~(layer6_outputs[3307]);
    assign outputs[4876] = ~((layer6_outputs[96]) | (layer6_outputs[1426]));
    assign outputs[4877] = ~(layer6_outputs[4495]);
    assign outputs[4878] = ~(layer6_outputs[4034]);
    assign outputs[4879] = layer6_outputs[1238];
    assign outputs[4880] = ~(layer6_outputs[1583]);
    assign outputs[4881] = ~((layer6_outputs[3527]) ^ (layer6_outputs[4421]));
    assign outputs[4882] = layer6_outputs[3844];
    assign outputs[4883] = layer6_outputs[1042];
    assign outputs[4884] = ~((layer6_outputs[1338]) | (layer6_outputs[3024]));
    assign outputs[4885] = ~((layer6_outputs[3649]) ^ (layer6_outputs[2271]));
    assign outputs[4886] = (layer6_outputs[264]) & (layer6_outputs[3379]);
    assign outputs[4887] = ~(layer6_outputs[4225]);
    assign outputs[4888] = (layer6_outputs[1051]) & ~(layer6_outputs[542]);
    assign outputs[4889] = layer6_outputs[2435];
    assign outputs[4890] = ~((layer6_outputs[2791]) ^ (layer6_outputs[2961]));
    assign outputs[4891] = layer6_outputs[1224];
    assign outputs[4892] = (layer6_outputs[4040]) ^ (layer6_outputs[4473]);
    assign outputs[4893] = layer6_outputs[1592];
    assign outputs[4894] = ~(layer6_outputs[4047]);
    assign outputs[4895] = (layer6_outputs[4350]) ^ (layer6_outputs[249]);
    assign outputs[4896] = layer6_outputs[3865];
    assign outputs[4897] = ~(layer6_outputs[3144]);
    assign outputs[4898] = (layer6_outputs[2644]) & ~(layer6_outputs[227]);
    assign outputs[4899] = ~(layer6_outputs[1968]);
    assign outputs[4900] = layer6_outputs[1156];
    assign outputs[4901] = ~((layer6_outputs[903]) ^ (layer6_outputs[1039]));
    assign outputs[4902] = layer6_outputs[4345];
    assign outputs[4903] = (layer6_outputs[3334]) & ~(layer6_outputs[1062]);
    assign outputs[4904] = layer6_outputs[3256];
    assign outputs[4905] = ~(layer6_outputs[2692]);
    assign outputs[4906] = ~((layer6_outputs[4578]) | (layer6_outputs[611]));
    assign outputs[4907] = ~(layer6_outputs[4410]);
    assign outputs[4908] = layer6_outputs[3709];
    assign outputs[4909] = layer6_outputs[274];
    assign outputs[4910] = (layer6_outputs[2585]) & ~(layer6_outputs[3756]);
    assign outputs[4911] = layer6_outputs[129];
    assign outputs[4912] = layer6_outputs[3834];
    assign outputs[4913] = (layer6_outputs[2783]) & ~(layer6_outputs[2401]);
    assign outputs[4914] = layer6_outputs[859];
    assign outputs[4915] = layer6_outputs[1225];
    assign outputs[4916] = layer6_outputs[2030];
    assign outputs[4917] = layer6_outputs[3229];
    assign outputs[4918] = ~(layer6_outputs[3532]);
    assign outputs[4919] = ~(layer6_outputs[3138]);
    assign outputs[4920] = ~(layer6_outputs[4120]);
    assign outputs[4921] = layer6_outputs[3079];
    assign outputs[4922] = layer6_outputs[1441];
    assign outputs[4923] = ~(layer6_outputs[1028]);
    assign outputs[4924] = ~(layer6_outputs[63]);
    assign outputs[4925] = ~(layer6_outputs[1550]);
    assign outputs[4926] = (layer6_outputs[2836]) ^ (layer6_outputs[1652]);
    assign outputs[4927] = layer6_outputs[4136];
    assign outputs[4928] = ~(layer6_outputs[4728]);
    assign outputs[4929] = ~(layer6_outputs[2087]);
    assign outputs[4930] = layer6_outputs[3274];
    assign outputs[4931] = (layer6_outputs[73]) & (layer6_outputs[2560]);
    assign outputs[4932] = (layer6_outputs[4620]) & ~(layer6_outputs[2113]);
    assign outputs[4933] = ~((layer6_outputs[3135]) | (layer6_outputs[3358]));
    assign outputs[4934] = ~(layer6_outputs[362]);
    assign outputs[4935] = (layer6_outputs[2543]) & ~(layer6_outputs[2551]);
    assign outputs[4936] = (layer6_outputs[3443]) & (layer6_outputs[4571]);
    assign outputs[4937] = ~(layer6_outputs[1832]);
    assign outputs[4938] = ~(layer6_outputs[1810]);
    assign outputs[4939] = ~(layer6_outputs[1347]);
    assign outputs[4940] = ~(layer6_outputs[2253]);
    assign outputs[4941] = ~(layer6_outputs[4226]) | (layer6_outputs[1981]);
    assign outputs[4942] = ~(layer6_outputs[3425]) | (layer6_outputs[1663]);
    assign outputs[4943] = layer6_outputs[4260];
    assign outputs[4944] = ~(layer6_outputs[2679]);
    assign outputs[4945] = (layer6_outputs[1944]) ^ (layer6_outputs[1370]);
    assign outputs[4946] = ~((layer6_outputs[2364]) ^ (layer6_outputs[199]));
    assign outputs[4947] = (layer6_outputs[3622]) ^ (layer6_outputs[3738]);
    assign outputs[4948] = layer6_outputs[2853];
    assign outputs[4949] = ~(layer6_outputs[2903]);
    assign outputs[4950] = (layer6_outputs[5090]) ^ (layer6_outputs[3251]);
    assign outputs[4951] = ~(layer6_outputs[194]);
    assign outputs[4952] = layer6_outputs[4182];
    assign outputs[4953] = (layer6_outputs[3998]) & ~(layer6_outputs[4966]);
    assign outputs[4954] = ~(layer6_outputs[1087]);
    assign outputs[4955] = layer6_outputs[2703];
    assign outputs[4956] = ~(layer6_outputs[3376]);
    assign outputs[4957] = layer6_outputs[1628];
    assign outputs[4958] = ~((layer6_outputs[2211]) ^ (layer6_outputs[1956]));
    assign outputs[4959] = ~(layer6_outputs[924]);
    assign outputs[4960] = ~(layer6_outputs[2170]) | (layer6_outputs[2508]);
    assign outputs[4961] = (layer6_outputs[2823]) ^ (layer6_outputs[3902]);
    assign outputs[4962] = layer6_outputs[2900];
    assign outputs[4963] = layer6_outputs[2884];
    assign outputs[4964] = (layer6_outputs[974]) ^ (layer6_outputs[3181]);
    assign outputs[4965] = ~((layer6_outputs[4787]) ^ (layer6_outputs[126]));
    assign outputs[4966] = ~(layer6_outputs[114]);
    assign outputs[4967] = layer6_outputs[1669];
    assign outputs[4968] = ~((layer6_outputs[1955]) | (layer6_outputs[3620]));
    assign outputs[4969] = layer6_outputs[2181];
    assign outputs[4970] = ~(layer6_outputs[4249]);
    assign outputs[4971] = (layer6_outputs[1902]) ^ (layer6_outputs[104]);
    assign outputs[4972] = (layer6_outputs[4579]) ^ (layer6_outputs[3774]);
    assign outputs[4973] = ~(layer6_outputs[1528]);
    assign outputs[4974] = layer6_outputs[3804];
    assign outputs[4975] = layer6_outputs[2713];
    assign outputs[4976] = ~(layer6_outputs[1327]);
    assign outputs[4977] = ~(layer6_outputs[419]);
    assign outputs[4978] = ~(layer6_outputs[4006]);
    assign outputs[4979] = (layer6_outputs[5009]) ^ (layer6_outputs[509]);
    assign outputs[4980] = ~((layer6_outputs[1852]) ^ (layer6_outputs[1659]));
    assign outputs[4981] = layer6_outputs[3356];
    assign outputs[4982] = layer6_outputs[4345];
    assign outputs[4983] = layer6_outputs[4030];
    assign outputs[4984] = (layer6_outputs[3284]) ^ (layer6_outputs[2391]);
    assign outputs[4985] = layer6_outputs[4032];
    assign outputs[4986] = ~((layer6_outputs[3175]) | (layer6_outputs[3515]));
    assign outputs[4987] = layer6_outputs[2687];
    assign outputs[4988] = (layer6_outputs[1216]) & (layer6_outputs[3269]);
    assign outputs[4989] = ~((layer6_outputs[4232]) | (layer6_outputs[458]));
    assign outputs[4990] = (layer6_outputs[4011]) ^ (layer6_outputs[1685]);
    assign outputs[4991] = ~(layer6_outputs[2618]);
    assign outputs[4992] = layer6_outputs[3438];
    assign outputs[4993] = layer6_outputs[2176];
    assign outputs[4994] = layer6_outputs[4604];
    assign outputs[4995] = layer6_outputs[2568];
    assign outputs[4996] = ~((layer6_outputs[3389]) ^ (layer6_outputs[4159]));
    assign outputs[4997] = (layer6_outputs[524]) ^ (layer6_outputs[4048]);
    assign outputs[4998] = (layer6_outputs[1541]) & ~(layer6_outputs[831]);
    assign outputs[4999] = layer6_outputs[2831];
    assign outputs[5000] = layer6_outputs[1560];
    assign outputs[5001] = ~(layer6_outputs[1140]);
    assign outputs[5002] = (layer6_outputs[2487]) ^ (layer6_outputs[1115]);
    assign outputs[5003] = ~((layer6_outputs[2456]) ^ (layer6_outputs[4432]));
    assign outputs[5004] = layer6_outputs[2589];
    assign outputs[5005] = (layer6_outputs[1524]) & (layer6_outputs[2530]);
    assign outputs[5006] = (layer6_outputs[3686]) | (layer6_outputs[2580]);
    assign outputs[5007] = layer6_outputs[1231];
    assign outputs[5008] = layer6_outputs[3914];
    assign outputs[5009] = ~((layer6_outputs[2866]) | (layer6_outputs[379]));
    assign outputs[5010] = layer6_outputs[738];
    assign outputs[5011] = layer6_outputs[4992];
    assign outputs[5012] = ~((layer6_outputs[263]) ^ (layer6_outputs[2324]));
    assign outputs[5013] = ~(layer6_outputs[876]);
    assign outputs[5014] = layer6_outputs[3547];
    assign outputs[5015] = (layer6_outputs[2793]) & ~(layer6_outputs[1732]);
    assign outputs[5016] = layer6_outputs[2008];
    assign outputs[5017] = ~((layer6_outputs[2301]) | (layer6_outputs[5076]));
    assign outputs[5018] = layer6_outputs[2462];
    assign outputs[5019] = ~((layer6_outputs[5097]) & (layer6_outputs[4993]));
    assign outputs[5020] = ~(layer6_outputs[2368]);
    assign outputs[5021] = ~(layer6_outputs[1680]);
    assign outputs[5022] = (layer6_outputs[706]) & (layer6_outputs[4597]);
    assign outputs[5023] = layer6_outputs[3239];
    assign outputs[5024] = ~(layer6_outputs[4028]);
    assign outputs[5025] = ~(layer6_outputs[588]);
    assign outputs[5026] = (layer6_outputs[3077]) ^ (layer6_outputs[1822]);
    assign outputs[5027] = layer6_outputs[1429];
    assign outputs[5028] = 1'b0;
    assign outputs[5029] = layer6_outputs[2184];
    assign outputs[5030] = ~((layer6_outputs[3970]) ^ (layer6_outputs[1636]));
    assign outputs[5031] = layer6_outputs[2663];
    assign outputs[5032] = layer6_outputs[3575];
    assign outputs[5033] = ~(layer6_outputs[4296]) | (layer6_outputs[3705]);
    assign outputs[5034] = layer6_outputs[2530];
    assign outputs[5035] = layer6_outputs[154];
    assign outputs[5036] = ~((layer6_outputs[4837]) ^ (layer6_outputs[1688]));
    assign outputs[5037] = ~(layer6_outputs[2955]);
    assign outputs[5038] = ~((layer6_outputs[4619]) ^ (layer6_outputs[1768]));
    assign outputs[5039] = (layer6_outputs[1719]) & (layer6_outputs[327]);
    assign outputs[5040] = ~(layer6_outputs[937]);
    assign outputs[5041] = layer6_outputs[1886];
    assign outputs[5042] = ~((layer6_outputs[1650]) ^ (layer6_outputs[4541]));
    assign outputs[5043] = ~(layer6_outputs[4550]);
    assign outputs[5044] = layer6_outputs[3639];
    assign outputs[5045] = ~(layer6_outputs[3589]);
    assign outputs[5046] = ~((layer6_outputs[4049]) ^ (layer6_outputs[4682]));
    assign outputs[5047] = (layer6_outputs[2952]) ^ (layer6_outputs[3632]);
    assign outputs[5048] = layer6_outputs[609];
    assign outputs[5049] = layer6_outputs[3227];
    assign outputs[5050] = ~((layer6_outputs[1069]) ^ (layer6_outputs[1021]));
    assign outputs[5051] = ~((layer6_outputs[4164]) ^ (layer6_outputs[1070]));
    assign outputs[5052] = (layer6_outputs[2213]) ^ (layer6_outputs[2207]);
    assign outputs[5053] = ~(layer6_outputs[3745]);
    assign outputs[5054] = layer6_outputs[67];
    assign outputs[5055] = ~(layer6_outputs[3291]);
    assign outputs[5056] = layer6_outputs[4152];
    assign outputs[5057] = (layer6_outputs[2387]) ^ (layer6_outputs[3592]);
    assign outputs[5058] = ~(layer6_outputs[2537]);
    assign outputs[5059] = ~(layer6_outputs[2467]);
    assign outputs[5060] = layer6_outputs[636];
    assign outputs[5061] = ~((layer6_outputs[2860]) | (layer6_outputs[4869]));
    assign outputs[5062] = ~(layer6_outputs[2314]);
    assign outputs[5063] = ~((layer6_outputs[3382]) ^ (layer6_outputs[3346]));
    assign outputs[5064] = ~(layer6_outputs[4047]);
    assign outputs[5065] = ~(layer6_outputs[2202]);
    assign outputs[5066] = layer6_outputs[2631];
    assign outputs[5067] = layer6_outputs[3042];
    assign outputs[5068] = (layer6_outputs[407]) ^ (layer6_outputs[3657]);
    assign outputs[5069] = layer6_outputs[731];
    assign outputs[5070] = layer6_outputs[4071];
    assign outputs[5071] = ~(layer6_outputs[2257]);
    assign outputs[5072] = layer6_outputs[2234];
    assign outputs[5073] = ~((layer6_outputs[4843]) ^ (layer6_outputs[2438]));
    assign outputs[5074] = ~(layer6_outputs[3980]) | (layer6_outputs[213]);
    assign outputs[5075] = ~(layer6_outputs[4876]);
    assign outputs[5076] = ~((layer6_outputs[2365]) ^ (layer6_outputs[781]));
    assign outputs[5077] = ~(layer6_outputs[4997]);
    assign outputs[5078] = (layer6_outputs[2713]) & ~(layer6_outputs[3264]);
    assign outputs[5079] = ~(layer6_outputs[1562]);
    assign outputs[5080] = ~(layer6_outputs[2355]);
    assign outputs[5081] = (layer6_outputs[4504]) & (layer6_outputs[261]);
    assign outputs[5082] = (layer6_outputs[2577]) ^ (layer6_outputs[1912]);
    assign outputs[5083] = ~(layer6_outputs[4967]) | (layer6_outputs[3095]);
    assign outputs[5084] = layer6_outputs[1213];
    assign outputs[5085] = ~(layer6_outputs[3009]);
    assign outputs[5086] = ~(layer6_outputs[574]);
    assign outputs[5087] = layer6_outputs[1530];
    assign outputs[5088] = (layer6_outputs[931]) & ~(layer6_outputs[1570]);
    assign outputs[5089] = layer6_outputs[3682];
    assign outputs[5090] = layer6_outputs[5016];
    assign outputs[5091] = ~((layer6_outputs[1138]) | (layer6_outputs[4774]));
    assign outputs[5092] = ~(layer6_outputs[4243]);
    assign outputs[5093] = (layer6_outputs[1014]) ^ (layer6_outputs[4606]);
    assign outputs[5094] = ~(layer6_outputs[295]);
    assign outputs[5095] = (layer6_outputs[4993]) ^ (layer6_outputs[1819]);
    assign outputs[5096] = ~((layer6_outputs[2811]) | (layer6_outputs[1201]));
    assign outputs[5097] = ~(layer6_outputs[361]);
    assign outputs[5098] = ~(layer6_outputs[3254]);
    assign outputs[5099] = ~(layer6_outputs[1896]) | (layer6_outputs[193]);
    assign outputs[5100] = layer6_outputs[4172];
    assign outputs[5101] = layer6_outputs[1761];
    assign outputs[5102] = ~(layer6_outputs[1697]);
    assign outputs[5103] = layer6_outputs[2199];
    assign outputs[5104] = ~(layer6_outputs[4454]);
    assign outputs[5105] = ~(layer6_outputs[159]);
    assign outputs[5106] = (layer6_outputs[2953]) ^ (layer6_outputs[1630]);
    assign outputs[5107] = ~((layer6_outputs[5005]) & (layer6_outputs[3841]));
    assign outputs[5108] = ~(layer6_outputs[295]);
    assign outputs[5109] = (layer6_outputs[1598]) ^ (layer6_outputs[1356]);
    assign outputs[5110] = ~(layer6_outputs[3464]);
    assign outputs[5111] = (layer6_outputs[180]) ^ (layer6_outputs[2162]);
    assign outputs[5112] = ~(layer6_outputs[3331]);
    assign outputs[5113] = ~(layer6_outputs[2257]);
    assign outputs[5114] = ~(layer6_outputs[2977]);
    assign outputs[5115] = (layer6_outputs[491]) & (layer6_outputs[4218]);
    assign outputs[5116] = ~(layer6_outputs[3475]);
    assign outputs[5117] = ~(layer6_outputs[2618]);
    assign outputs[5118] = ~(layer6_outputs[4936]);
    assign outputs[5119] = ~((layer6_outputs[4266]) ^ (layer6_outputs[4406]));
endmodule
