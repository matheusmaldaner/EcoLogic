module logic_network(
	// Whatever i need for input SRAM
   // input wire [399:0] inputs,
    output reg [9:0] classification
);

	 wire [399:0] inputs;
    wire [2499:0] layer0_outputs;
	 wire [2499:0] outputs;

    assign layer0_outputs[0] = ~(inputs[303]) | (inputs[179]);
    assign layer0_outputs[1] = inputs[193];
    assign layer0_outputs[2] = (inputs[66]) & (inputs[72]);
    assign layer0_outputs[3] = ~(inputs[199]);
    assign layer0_outputs[4] = ~((inputs[361]) | (inputs[30]));
    assign layer0_outputs[5] = ~(inputs[244]);
    assign layer0_outputs[6] = (inputs[196]) ^ (inputs[8]);
    assign layer0_outputs[7] = ~(inputs[173]) | (inputs[378]);
    assign layer0_outputs[8] = (inputs[228]) & ~(inputs[356]);
    assign layer0_outputs[9] = ~(inputs[114]) | (inputs[332]);
    assign layer0_outputs[10] = (inputs[73]) | (inputs[284]);
    assign layer0_outputs[11] = ~(inputs[207]) | (inputs[24]);
    assign layer0_outputs[12] = (inputs[328]) & ~(inputs[398]);
    assign layer0_outputs[13] = (inputs[167]) | (inputs[106]);
    assign layer0_outputs[14] = (inputs[367]) ^ (inputs[161]);
    assign layer0_outputs[15] = inputs[116];
    assign layer0_outputs[16] = (inputs[1]) | (inputs[398]);
    assign layer0_outputs[17] = ~(inputs[156]);
    assign layer0_outputs[18] = (inputs[245]) & ~(inputs[292]);
    assign layer0_outputs[19] = (inputs[275]) ^ (inputs[153]);
    assign layer0_outputs[20] = (inputs[144]) | (inputs[247]);
    assign layer0_outputs[21] = ~(inputs[206]);
    assign layer0_outputs[22] = ~((inputs[29]) | (inputs[101]));
    assign layer0_outputs[23] = inputs[4];
    assign layer0_outputs[24] = ~((inputs[357]) & (inputs[83]));
    assign layer0_outputs[25] = inputs[177];
    assign layer0_outputs[26] = inputs[272];
    assign layer0_outputs[27] = ~(inputs[346]) | (inputs[57]);
    assign layer0_outputs[28] = inputs[115];
    assign layer0_outputs[29] = ~(inputs[133]);
    assign layer0_outputs[30] = inputs[363];
    assign layer0_outputs[31] = ~(inputs[137]);
    assign layer0_outputs[32] = (inputs[106]) | (inputs[178]);
    assign layer0_outputs[33] = ~(inputs[207]);
    assign layer0_outputs[34] = ~(inputs[388]) | (inputs[5]);
    assign layer0_outputs[35] = ~(inputs[345]);
    assign layer0_outputs[36] = (inputs[127]) & ~(inputs[238]);
    assign layer0_outputs[37] = (inputs[66]) | (inputs[119]);
    assign layer0_outputs[38] = (inputs[269]) & (inputs[172]);
    assign layer0_outputs[39] = (inputs[304]) | (inputs[341]);
    assign layer0_outputs[40] = ~(inputs[135]);
    assign layer0_outputs[41] = ~((inputs[8]) | (inputs[191]));
    assign layer0_outputs[42] = ~((inputs[389]) | (inputs[239]));
    assign layer0_outputs[43] = ~(inputs[108]) | (inputs[378]);
    assign layer0_outputs[44] = inputs[210];
    assign layer0_outputs[45] = (inputs[333]) | (inputs[354]);
    assign layer0_outputs[46] = inputs[175];
    assign layer0_outputs[47] = inputs[163];
    assign layer0_outputs[48] = inputs[366];
    assign layer0_outputs[49] = inputs[245];
    assign layer0_outputs[50] = ~(inputs[64]);
    assign layer0_outputs[51] = (inputs[76]) ^ (inputs[177]);
    assign layer0_outputs[52] = (inputs[210]) & ~(inputs[63]);
    assign layer0_outputs[53] = ~(inputs[288]);
    assign layer0_outputs[54] = (inputs[192]) | (inputs[327]);
    assign layer0_outputs[55] = (inputs[85]) | (inputs[143]);
    assign layer0_outputs[56] = ~((inputs[184]) | (inputs[301]));
    assign layer0_outputs[57] = ~((inputs[161]) | (inputs[395]));
    assign layer0_outputs[58] = 1'b0;
    assign layer0_outputs[59] = ~((inputs[158]) | (inputs[67]));
    assign layer0_outputs[60] = (inputs[119]) ^ (inputs[30]);
    assign layer0_outputs[61] = ~((inputs[287]) ^ (inputs[44]));
    assign layer0_outputs[62] = ~(inputs[134]);
    assign layer0_outputs[63] = (inputs[60]) ^ (inputs[117]);
    assign layer0_outputs[64] = ~((inputs[302]) | (inputs[87]));
    assign layer0_outputs[65] = (inputs[398]) | (inputs[73]);
    assign layer0_outputs[66] = ~(inputs[150]);
    assign layer0_outputs[67] = (inputs[287]) & ~(inputs[77]);
    assign layer0_outputs[68] = inputs[375];
    assign layer0_outputs[69] = ~(inputs[47]) | (inputs[241]);
    assign layer0_outputs[70] = inputs[222];
    assign layer0_outputs[71] = inputs[393];
    assign layer0_outputs[72] = (inputs[223]) | (inputs[201]);
    assign layer0_outputs[73] = (inputs[274]) | (inputs[363]);
    assign layer0_outputs[74] = ~((inputs[344]) | (inputs[197]));
    assign layer0_outputs[75] = ~((inputs[279]) ^ (inputs[386]));
    assign layer0_outputs[76] = (inputs[119]) | (inputs[384]);
    assign layer0_outputs[77] = ~(inputs[136]);
    assign layer0_outputs[78] = ~(inputs[308]) | (inputs[199]);
    assign layer0_outputs[79] = ~(inputs[323]);
    assign layer0_outputs[80] = (inputs[199]) | (inputs[330]);
    assign layer0_outputs[81] = ~((inputs[61]) & (inputs[381]));
    assign layer0_outputs[82] = ~(inputs[186]) | (inputs[281]);
    assign layer0_outputs[83] = (inputs[263]) | (inputs[157]);
    assign layer0_outputs[84] = (inputs[174]) | (inputs[157]);
    assign layer0_outputs[85] = (inputs[167]) | (inputs[144]);
    assign layer0_outputs[86] = inputs[267];
    assign layer0_outputs[87] = (inputs[358]) & ~(inputs[136]);
    assign layer0_outputs[88] = ~((inputs[84]) | (inputs[287]));
    assign layer0_outputs[89] = (inputs[206]) & (inputs[93]);
    assign layer0_outputs[90] = 1'b0;
    assign layer0_outputs[91] = (inputs[225]) & ~(inputs[239]);
    assign layer0_outputs[92] = inputs[273];
    assign layer0_outputs[93] = inputs[205];
    assign layer0_outputs[94] = ~(inputs[50]) | (inputs[26]);
    assign layer0_outputs[95] = inputs[177];
    assign layer0_outputs[96] = (inputs[258]) ^ (inputs[49]);
    assign layer0_outputs[97] = ~((inputs[373]) ^ (inputs[303]));
    assign layer0_outputs[98] = (inputs[218]) & ~(inputs[2]);
    assign layer0_outputs[99] = (inputs[284]) ^ (inputs[293]);
    assign layer0_outputs[100] = ~(inputs[325]);
    assign layer0_outputs[101] = ~(inputs[287]) | (inputs[232]);
    assign layer0_outputs[102] = 1'b1;
    assign layer0_outputs[103] = ~(inputs[171]);
    assign layer0_outputs[104] = ~(inputs[169]);
    assign layer0_outputs[105] = (inputs[185]) ^ (inputs[130]);
    assign layer0_outputs[106] = (inputs[195]) & ~(inputs[358]);
    assign layer0_outputs[107] = inputs[313];
    assign layer0_outputs[108] = ~(inputs[326]) | (inputs[220]);
    assign layer0_outputs[109] = ~((inputs[45]) | (inputs[111]));
    assign layer0_outputs[110] = ~(inputs[312]);
    assign layer0_outputs[111] = ~(inputs[267]);
    assign layer0_outputs[112] = ~((inputs[77]) ^ (inputs[162]));
    assign layer0_outputs[113] = inputs[189];
    assign layer0_outputs[114] = (inputs[68]) & (inputs[15]);
    assign layer0_outputs[115] = ~((inputs[197]) | (inputs[76]));
    assign layer0_outputs[116] = (inputs[57]) | (inputs[23]);
    assign layer0_outputs[117] = (inputs[350]) ^ (inputs[390]);
    assign layer0_outputs[118] = (inputs[385]) | (inputs[263]);
    assign layer0_outputs[119] = (inputs[205]) | (inputs[88]);
    assign layer0_outputs[120] = (inputs[239]) & ~(inputs[71]);
    assign layer0_outputs[121] = (inputs[65]) & ~(inputs[58]);
    assign layer0_outputs[122] = (inputs[115]) | (inputs[398]);
    assign layer0_outputs[123] = (inputs[70]) & ~(inputs[388]);
    assign layer0_outputs[124] = (inputs[279]) | (inputs[356]);
    assign layer0_outputs[125] = inputs[136];
    assign layer0_outputs[126] = inputs[284];
    assign layer0_outputs[127] = ~((inputs[45]) | (inputs[33]));
    assign layer0_outputs[128] = inputs[245];
    assign layer0_outputs[129] = inputs[164];
    assign layer0_outputs[130] = (inputs[210]) & ~(inputs[213]);
    assign layer0_outputs[131] = ~(inputs[371]);
    assign layer0_outputs[132] = (inputs[175]) & ~(inputs[257]);
    assign layer0_outputs[133] = (inputs[50]) & ~(inputs[396]);
    assign layer0_outputs[134] = ~((inputs[121]) | (inputs[208]));
    assign layer0_outputs[135] = inputs[145];
    assign layer0_outputs[136] = ~(inputs[350]) | (inputs[47]);
    assign layer0_outputs[137] = ~(inputs[170]);
    assign layer0_outputs[138] = (inputs[284]) & ~(inputs[22]);
    assign layer0_outputs[139] = (inputs[391]) | (inputs[266]);
    assign layer0_outputs[140] = ~((inputs[210]) ^ (inputs[224]));
    assign layer0_outputs[141] = (inputs[258]) & ~(inputs[149]);
    assign layer0_outputs[142] = ~(inputs[168]) | (inputs[343]);
    assign layer0_outputs[143] = inputs[186];
    assign layer0_outputs[144] = (inputs[150]) ^ (inputs[80]);
    assign layer0_outputs[145] = ~((inputs[218]) | (inputs[14]));
    assign layer0_outputs[146] = ~((inputs[347]) | (inputs[281]));
    assign layer0_outputs[147] = inputs[38];
    assign layer0_outputs[148] = (inputs[316]) | (inputs[27]);
    assign layer0_outputs[149] = ~((inputs[267]) ^ (inputs[96]));
    assign layer0_outputs[150] = ~(inputs[390]);
    assign layer0_outputs[151] = inputs[202];
    assign layer0_outputs[152] = (inputs[114]) | (inputs[290]);
    assign layer0_outputs[153] = ~((inputs[47]) ^ (inputs[256]));
    assign layer0_outputs[154] = (inputs[200]) | (inputs[205]);
    assign layer0_outputs[155] = (inputs[96]) | (inputs[237]);
    assign layer0_outputs[156] = (inputs[328]) & ~(inputs[75]);
    assign layer0_outputs[157] = ~(inputs[360]);
    assign layer0_outputs[158] = (inputs[293]) & ~(inputs[201]);
    assign layer0_outputs[159] = ~(inputs[9]);
    assign layer0_outputs[160] = (inputs[314]) ^ (inputs[79]);
    assign layer0_outputs[161] = ~(inputs[113]) | (inputs[223]);
    assign layer0_outputs[162] = ~((inputs[24]) | (inputs[304]));
    assign layer0_outputs[163] = ~(inputs[203]);
    assign layer0_outputs[164] = ~((inputs[67]) ^ (inputs[63]));
    assign layer0_outputs[165] = (inputs[311]) | (inputs[161]);
    assign layer0_outputs[166] = ~((inputs[42]) ^ (inputs[83]));
    assign layer0_outputs[167] = ~((inputs[266]) | (inputs[19]));
    assign layer0_outputs[168] = (inputs[366]) ^ (inputs[347]);
    assign layer0_outputs[169] = inputs[361];
    assign layer0_outputs[170] = ~(inputs[186]) | (inputs[281]);
    assign layer0_outputs[171] = (inputs[44]) & ~(inputs[161]);
    assign layer0_outputs[172] = (inputs[371]) ^ (inputs[361]);
    assign layer0_outputs[173] = (inputs[321]) | (inputs[42]);
    assign layer0_outputs[174] = ~(inputs[231]);
    assign layer0_outputs[175] = ~(inputs[50]);
    assign layer0_outputs[176] = (inputs[364]) | (inputs[209]);
    assign layer0_outputs[177] = inputs[274];
    assign layer0_outputs[178] = (inputs[377]) & (inputs[385]);
    assign layer0_outputs[179] = (inputs[169]) & (inputs[371]);
    assign layer0_outputs[180] = ~(inputs[142]);
    assign layer0_outputs[181] = inputs[44];
    assign layer0_outputs[182] = inputs[66];
    assign layer0_outputs[183] = inputs[37];
    assign layer0_outputs[184] = inputs[36];
    assign layer0_outputs[185] = ~(inputs[307]);
    assign layer0_outputs[186] = ~(inputs[372]);
    assign layer0_outputs[187] = 1'b1;
    assign layer0_outputs[188] = ~(inputs[30]);
    assign layer0_outputs[189] = ~(inputs[318]);
    assign layer0_outputs[190] = inputs[157];
    assign layer0_outputs[191] = inputs[257];
    assign layer0_outputs[192] = ~(inputs[89]) | (inputs[5]);
    assign layer0_outputs[193] = ~(inputs[284]);
    assign layer0_outputs[194] = inputs[31];
    assign layer0_outputs[195] = ~(inputs[106]);
    assign layer0_outputs[196] = (inputs[205]) & ~(inputs[299]);
    assign layer0_outputs[197] = ~((inputs[385]) | (inputs[326]));
    assign layer0_outputs[198] = ~((inputs[12]) ^ (inputs[311]));
    assign layer0_outputs[199] = ~((inputs[320]) | (inputs[260]));
    assign layer0_outputs[200] = ~(inputs[350]);
    assign layer0_outputs[201] = ~((inputs[5]) ^ (inputs[33]));
    assign layer0_outputs[202] = ~(inputs[264]) | (inputs[92]);
    assign layer0_outputs[203] = ~((inputs[236]) ^ (inputs[177]));
    assign layer0_outputs[204] = (inputs[51]) & ~(inputs[220]);
    assign layer0_outputs[205] = ~(inputs[26]) | (inputs[75]);
    assign layer0_outputs[206] = inputs[269];
    assign layer0_outputs[207] = ~((inputs[77]) ^ (inputs[34]));
    assign layer0_outputs[208] = (inputs[138]) | (inputs[312]);
    assign layer0_outputs[209] = inputs[39];
    assign layer0_outputs[210] = inputs[210];
    assign layer0_outputs[211] = ~(inputs[105]) | (inputs[394]);
    assign layer0_outputs[212] = ~((inputs[79]) | (inputs[323]));
    assign layer0_outputs[213] = ~((inputs[167]) | (inputs[19]));
    assign layer0_outputs[214] = ~((inputs[397]) | (inputs[104]));
    assign layer0_outputs[215] = ~(inputs[384]);
    assign layer0_outputs[216] = (inputs[375]) ^ (inputs[366]);
    assign layer0_outputs[217] = (inputs[399]) ^ (inputs[150]);
    assign layer0_outputs[218] = (inputs[74]) & ~(inputs[147]);
    assign layer0_outputs[219] = ~((inputs[61]) | (inputs[259]));
    assign layer0_outputs[220] = (inputs[36]) | (inputs[287]);
    assign layer0_outputs[221] = (inputs[286]) & ~(inputs[79]);
    assign layer0_outputs[222] = (inputs[364]) & ~(inputs[83]);
    assign layer0_outputs[223] = (inputs[389]) ^ (inputs[197]);
    assign layer0_outputs[224] = (inputs[6]) | (inputs[133]);
    assign layer0_outputs[225] = (inputs[376]) ^ (inputs[106]);
    assign layer0_outputs[226] = ~((inputs[180]) | (inputs[206]));
    assign layer0_outputs[227] = ~(inputs[220]) | (inputs[339]);
    assign layer0_outputs[228] = ~(inputs[165]);
    assign layer0_outputs[229] = ~(inputs[289]);
    assign layer0_outputs[230] = ~(inputs[345]) | (inputs[70]);
    assign layer0_outputs[231] = inputs[68];
    assign layer0_outputs[232] = inputs[86];
    assign layer0_outputs[233] = 1'b1;
    assign layer0_outputs[234] = ~((inputs[78]) ^ (inputs[58]));
    assign layer0_outputs[235] = (inputs[192]) & ~(inputs[348]);
    assign layer0_outputs[236] = ~(inputs[138]);
    assign layer0_outputs[237] = ~((inputs[158]) | (inputs[20]));
    assign layer0_outputs[238] = (inputs[250]) ^ (inputs[35]);
    assign layer0_outputs[239] = ~((inputs[221]) | (inputs[144]));
    assign layer0_outputs[240] = (inputs[345]) ^ (inputs[102]);
    assign layer0_outputs[241] = (inputs[295]) ^ (inputs[324]);
    assign layer0_outputs[242] = ~((inputs[198]) | (inputs[255]));
    assign layer0_outputs[243] = inputs[51];
    assign layer0_outputs[244] = ~(inputs[134]) | (inputs[351]);
    assign layer0_outputs[245] = (inputs[253]) ^ (inputs[354]);
    assign layer0_outputs[246] = ~((inputs[4]) | (inputs[126]));
    assign layer0_outputs[247] = inputs[58];
    assign layer0_outputs[248] = ~((inputs[1]) ^ (inputs[328]));
    assign layer0_outputs[249] = ~((inputs[63]) | (inputs[255]));
    assign layer0_outputs[250] = inputs[23];
    assign layer0_outputs[251] = inputs[155];
    assign layer0_outputs[252] = (inputs[131]) & ~(inputs[375]);
    assign layer0_outputs[253] = inputs[253];
    assign layer0_outputs[254] = (inputs[197]) | (inputs[28]);
    assign layer0_outputs[255] = (inputs[2]) | (inputs[9]);
    assign layer0_outputs[256] = (inputs[54]) & ~(inputs[311]);
    assign layer0_outputs[257] = ~(inputs[18]);
    assign layer0_outputs[258] = ~(inputs[33]);
    assign layer0_outputs[259] = ~(inputs[304]);
    assign layer0_outputs[260] = (inputs[382]) | (inputs[332]);
    assign layer0_outputs[261] = ~((inputs[349]) & (inputs[29]));
    assign layer0_outputs[262] = (inputs[338]) & ~(inputs[16]);
    assign layer0_outputs[263] = ~(inputs[87]) | (inputs[373]);
    assign layer0_outputs[264] = (inputs[146]) & ~(inputs[215]);
    assign layer0_outputs[265] = (inputs[107]) | (inputs[11]);
    assign layer0_outputs[266] = ~((inputs[214]) | (inputs[88]));
    assign layer0_outputs[267] = ~(inputs[262]);
    assign layer0_outputs[268] = ~(inputs[317]);
    assign layer0_outputs[269] = (inputs[189]) & ~(inputs[383]);
    assign layer0_outputs[270] = ~(inputs[143]);
    assign layer0_outputs[271] = inputs[167];
    assign layer0_outputs[272] = (inputs[208]) ^ (inputs[244]);
    assign layer0_outputs[273] = inputs[287];
    assign layer0_outputs[274] = (inputs[185]) & ~(inputs[339]);
    assign layer0_outputs[275] = (inputs[364]) ^ (inputs[13]);
    assign layer0_outputs[276] = ~(inputs[190]);
    assign layer0_outputs[277] = (inputs[241]) ^ (inputs[283]);
    assign layer0_outputs[278] = ~(inputs[52]) | (inputs[206]);
    assign layer0_outputs[279] = ~(inputs[231]);
    assign layer0_outputs[280] = ~(inputs[136]) | (inputs[338]);
    assign layer0_outputs[281] = inputs[243];
    assign layer0_outputs[282] = inputs[159];
    assign layer0_outputs[283] = inputs[23];
    assign layer0_outputs[284] = ~(inputs[17]) | (inputs[242]);
    assign layer0_outputs[285] = ~((inputs[338]) ^ (inputs[201]));
    assign layer0_outputs[286] = (inputs[70]) ^ (inputs[69]);
    assign layer0_outputs[287] = ~(inputs[86]) | (inputs[277]);
    assign layer0_outputs[288] = ~(inputs[228]) | (inputs[377]);
    assign layer0_outputs[289] = (inputs[240]) | (inputs[82]);
    assign layer0_outputs[290] = (inputs[222]) | (inputs[297]);
    assign layer0_outputs[291] = inputs[111];
    assign layer0_outputs[292] = inputs[329];
    assign layer0_outputs[293] = ~(inputs[255]);
    assign layer0_outputs[294] = inputs[231];
    assign layer0_outputs[295] = inputs[325];
    assign layer0_outputs[296] = ~((inputs[313]) | (inputs[301]));
    assign layer0_outputs[297] = ~(inputs[267]) | (inputs[43]);
    assign layer0_outputs[298] = inputs[193];
    assign layer0_outputs[299] = (inputs[101]) & (inputs[79]);
    assign layer0_outputs[300] = ~(inputs[352]) | (inputs[157]);
    assign layer0_outputs[301] = ~(inputs[249]);
    assign layer0_outputs[302] = inputs[155];
    assign layer0_outputs[303] = (inputs[243]) & ~(inputs[129]);
    assign layer0_outputs[304] = ~((inputs[254]) | (inputs[186]));
    assign layer0_outputs[305] = ~((inputs[301]) ^ (inputs[354]));
    assign layer0_outputs[306] = (inputs[98]) | (inputs[293]);
    assign layer0_outputs[307] = (inputs[246]) | (inputs[297]);
    assign layer0_outputs[308] = inputs[53];
    assign layer0_outputs[309] = 1'b1;
    assign layer0_outputs[310] = (inputs[85]) & ~(inputs[229]);
    assign layer0_outputs[311] = ~(inputs[31]);
    assign layer0_outputs[312] = (inputs[100]) | (inputs[81]);
    assign layer0_outputs[313] = ~(inputs[285]) | (inputs[156]);
    assign layer0_outputs[314] = inputs[232];
    assign layer0_outputs[315] = ~(inputs[49]);
    assign layer0_outputs[316] = ~(inputs[352]);
    assign layer0_outputs[317] = inputs[138];
    assign layer0_outputs[318] = (inputs[101]) | (inputs[22]);
    assign layer0_outputs[319] = ~(inputs[144]);
    assign layer0_outputs[320] = (inputs[83]) & ~(inputs[181]);
    assign layer0_outputs[321] = ~(inputs[325]) | (inputs[294]);
    assign layer0_outputs[322] = (inputs[310]) | (inputs[397]);
    assign layer0_outputs[323] = ~(inputs[139]);
    assign layer0_outputs[324] = ~(inputs[286]) | (inputs[153]);
    assign layer0_outputs[325] = ~(inputs[27]);
    assign layer0_outputs[326] = inputs[265];
    assign layer0_outputs[327] = (inputs[345]) & ~(inputs[198]);
    assign layer0_outputs[328] = (inputs[104]) & ~(inputs[248]);
    assign layer0_outputs[329] = (inputs[296]) | (inputs[77]);
    assign layer0_outputs[330] = inputs[203];
    assign layer0_outputs[331] = ~(inputs[192]) | (inputs[206]);
    assign layer0_outputs[332] = ~((inputs[294]) | (inputs[157]));
    assign layer0_outputs[333] = ~(inputs[289]) | (inputs[74]);
    assign layer0_outputs[334] = ~(inputs[134]);
    assign layer0_outputs[335] = (inputs[242]) | (inputs[122]);
    assign layer0_outputs[336] = ~((inputs[53]) & (inputs[87]));
    assign layer0_outputs[337] = inputs[361];
    assign layer0_outputs[338] = (inputs[371]) & ~(inputs[118]);
    assign layer0_outputs[339] = ~((inputs[357]) ^ (inputs[223]));
    assign layer0_outputs[340] = ~((inputs[292]) ^ (inputs[61]));
    assign layer0_outputs[341] = (inputs[38]) | (inputs[394]);
    assign layer0_outputs[342] = (inputs[204]) & ~(inputs[383]);
    assign layer0_outputs[343] = (inputs[61]) | (inputs[290]);
    assign layer0_outputs[344] = ~(inputs[254]) | (inputs[362]);
    assign layer0_outputs[345] = ~(inputs[155]);
    assign layer0_outputs[346] = ~(inputs[297]);
    assign layer0_outputs[347] = ~(inputs[140]) | (inputs[118]);
    assign layer0_outputs[348] = inputs[11];
    assign layer0_outputs[349] = (inputs[340]) | (inputs[135]);
    assign layer0_outputs[350] = ~((inputs[110]) | (inputs[92]));
    assign layer0_outputs[351] = (inputs[232]) | (inputs[94]);
    assign layer0_outputs[352] = (inputs[256]) | (inputs[305]);
    assign layer0_outputs[353] = inputs[162];
    assign layer0_outputs[354] = (inputs[375]) | (inputs[368]);
    assign layer0_outputs[355] = ~((inputs[307]) ^ (inputs[350]));
    assign layer0_outputs[356] = ~(inputs[106]);
    assign layer0_outputs[357] = inputs[74];
    assign layer0_outputs[358] = ~(inputs[344]);
    assign layer0_outputs[359] = (inputs[291]) & (inputs[296]);
    assign layer0_outputs[360] = (inputs[52]) & ~(inputs[132]);
    assign layer0_outputs[361] = ~(inputs[308]) | (inputs[299]);
    assign layer0_outputs[362] = (inputs[349]) & (inputs[116]);
    assign layer0_outputs[363] = ~(inputs[175]) | (inputs[63]);
    assign layer0_outputs[364] = inputs[188];
    assign layer0_outputs[365] = (inputs[324]) & ~(inputs[399]);
    assign layer0_outputs[366] = ~((inputs[110]) | (inputs[315]));
    assign layer0_outputs[367] = (inputs[318]) | (inputs[362]);
    assign layer0_outputs[368] = (inputs[74]) ^ (inputs[21]);
    assign layer0_outputs[369] = (inputs[109]) & ~(inputs[46]);
    assign layer0_outputs[370] = (inputs[237]) | (inputs[333]);
    assign layer0_outputs[371] = inputs[135];
    assign layer0_outputs[372] = ~(inputs[46]);
    assign layer0_outputs[373] = inputs[191];
    assign layer0_outputs[374] = ~((inputs[180]) ^ (inputs[234]));
    assign layer0_outputs[375] = (inputs[230]) | (inputs[269]);
    assign layer0_outputs[376] = inputs[397];
    assign layer0_outputs[377] = ~((inputs[20]) ^ (inputs[390]));
    assign layer0_outputs[378] = ~(inputs[109]);
    assign layer0_outputs[379] = ~(inputs[229]);
    assign layer0_outputs[380] = (inputs[274]) | (inputs[255]);
    assign layer0_outputs[381] = ~(inputs[186]);
    assign layer0_outputs[382] = ~(inputs[391]);
    assign layer0_outputs[383] = inputs[94];
    assign layer0_outputs[384] = ~((inputs[96]) & (inputs[49]));
    assign layer0_outputs[385] = (inputs[328]) & (inputs[363]);
    assign layer0_outputs[386] = inputs[43];
    assign layer0_outputs[387] = inputs[310];
    assign layer0_outputs[388] = (inputs[91]) & (inputs[279]);
    assign layer0_outputs[389] = ~(inputs[169]);
    assign layer0_outputs[390] = (inputs[394]) ^ (inputs[289]);
    assign layer0_outputs[391] = inputs[13];
    assign layer0_outputs[392] = (inputs[214]) | (inputs[218]);
    assign layer0_outputs[393] = (inputs[163]) ^ (inputs[131]);
    assign layer0_outputs[394] = inputs[208];
    assign layer0_outputs[395] = (inputs[137]) | (inputs[38]);
    assign layer0_outputs[396] = (inputs[158]) & ~(inputs[42]);
    assign layer0_outputs[397] = ~(inputs[390]) | (inputs[119]);
    assign layer0_outputs[398] = ~(inputs[315]) | (inputs[124]);
    assign layer0_outputs[399] = ~(inputs[148]) | (inputs[110]);
    assign layer0_outputs[400] = ~((inputs[53]) ^ (inputs[90]));
    assign layer0_outputs[401] = ~(inputs[335]);
    assign layer0_outputs[402] = (inputs[131]) & ~(inputs[373]);
    assign layer0_outputs[403] = ~(inputs[219]) | (inputs[266]);
    assign layer0_outputs[404] = ~(inputs[6]) | (inputs[179]);
    assign layer0_outputs[405] = (inputs[369]) & ~(inputs[398]);
    assign layer0_outputs[406] = ~(inputs[350]);
    assign layer0_outputs[407] = ~(inputs[134]);
    assign layer0_outputs[408] = ~((inputs[2]) ^ (inputs[67]));
    assign layer0_outputs[409] = (inputs[89]) ^ (inputs[50]);
    assign layer0_outputs[410] = inputs[84];
    assign layer0_outputs[411] = ~(inputs[47]);
    assign layer0_outputs[412] = ~(inputs[144]) | (inputs[363]);
    assign layer0_outputs[413] = ~(inputs[37]);
    assign layer0_outputs[414] = inputs[326];
    assign layer0_outputs[415] = ~((inputs[352]) ^ (inputs[87]));
    assign layer0_outputs[416] = ~((inputs[293]) ^ (inputs[300]));
    assign layer0_outputs[417] = inputs[211];
    assign layer0_outputs[418] = ~((inputs[304]) | (inputs[286]));
    assign layer0_outputs[419] = (inputs[271]) | (inputs[78]);
    assign layer0_outputs[420] = ~(inputs[134]);
    assign layer0_outputs[421] = (inputs[41]) | (inputs[357]);
    assign layer0_outputs[422] = ~(inputs[143]);
    assign layer0_outputs[423] = (inputs[343]) & ~(inputs[37]);
    assign layer0_outputs[424] = (inputs[109]) & ~(inputs[256]);
    assign layer0_outputs[425] = (inputs[220]) & ~(inputs[311]);
    assign layer0_outputs[426] = (inputs[32]) & ~(inputs[263]);
    assign layer0_outputs[427] = ~(inputs[378]) | (inputs[104]);
    assign layer0_outputs[428] = ~(inputs[373]);
    assign layer0_outputs[429] = ~((inputs[1]) | (inputs[257]));
    assign layer0_outputs[430] = (inputs[299]) & ~(inputs[262]);
    assign layer0_outputs[431] = ~((inputs[117]) | (inputs[203]));
    assign layer0_outputs[432] = ~(inputs[391]);
    assign layer0_outputs[433] = ~(inputs[55]);
    assign layer0_outputs[434] = ~(inputs[150]);
    assign layer0_outputs[435] = ~(inputs[351]);
    assign layer0_outputs[436] = (inputs[213]) & ~(inputs[259]);
    assign layer0_outputs[437] = (inputs[186]) ^ (inputs[141]);
    assign layer0_outputs[438] = ~(inputs[84]);
    assign layer0_outputs[439] = (inputs[49]) & ~(inputs[43]);
    assign layer0_outputs[440] = ~((inputs[312]) | (inputs[74]));
    assign layer0_outputs[441] = ~(inputs[104]);
    assign layer0_outputs[442] = 1'b0;
    assign layer0_outputs[443] = (inputs[42]) | (inputs[255]);
    assign layer0_outputs[444] = (inputs[59]) & ~(inputs[116]);
    assign layer0_outputs[445] = ~(inputs[90]);
    assign layer0_outputs[446] = inputs[56];
    assign layer0_outputs[447] = ~(inputs[140]);
    assign layer0_outputs[448] = (inputs[327]) & ~(inputs[397]);
    assign layer0_outputs[449] = ~(inputs[190]) | (inputs[100]);
    assign layer0_outputs[450] = ~(inputs[347]) | (inputs[218]);
    assign layer0_outputs[451] = ~(inputs[324]) | (inputs[1]);
    assign layer0_outputs[452] = (inputs[255]) ^ (inputs[372]);
    assign layer0_outputs[453] = ~(inputs[244]);
    assign layer0_outputs[454] = ~(inputs[305]) | (inputs[0]);
    assign layer0_outputs[455] = ~(inputs[342]);
    assign layer0_outputs[456] = inputs[170];
    assign layer0_outputs[457] = inputs[374];
    assign layer0_outputs[458] = inputs[356];
    assign layer0_outputs[459] = (inputs[108]) | (inputs[254]);
    assign layer0_outputs[460] = (inputs[179]) ^ (inputs[50]);
    assign layer0_outputs[461] = inputs[243];
    assign layer0_outputs[462] = ~(inputs[268]) | (inputs[199]);
    assign layer0_outputs[463] = ~((inputs[337]) | (inputs[224]));
    assign layer0_outputs[464] = ~(inputs[344]) | (inputs[30]);
    assign layer0_outputs[465] = ~(inputs[129]);
    assign layer0_outputs[466] = inputs[235];
    assign layer0_outputs[467] = inputs[112];
    assign layer0_outputs[468] = (inputs[147]) ^ (inputs[161]);
    assign layer0_outputs[469] = (inputs[124]) & ~(inputs[100]);
    assign layer0_outputs[470] = ~((inputs[353]) | (inputs[157]));
    assign layer0_outputs[471] = ~(inputs[182]);
    assign layer0_outputs[472] = inputs[2];
    assign layer0_outputs[473] = ~(inputs[340]);
    assign layer0_outputs[474] = ~(inputs[250]) | (inputs[361]);
    assign layer0_outputs[475] = (inputs[380]) & (inputs[118]);
    assign layer0_outputs[476] = (inputs[283]) & (inputs[124]);
    assign layer0_outputs[477] = (inputs[60]) & (inputs[64]);
    assign layer0_outputs[478] = (inputs[23]) | (inputs[353]);
    assign layer0_outputs[479] = (inputs[293]) ^ (inputs[353]);
    assign layer0_outputs[480] = ~((inputs[39]) | (inputs[174]));
    assign layer0_outputs[481] = ~(inputs[75]);
    assign layer0_outputs[482] = ~(inputs[243]) | (inputs[177]);
    assign layer0_outputs[483] = inputs[284];
    assign layer0_outputs[484] = ~(inputs[197]) | (inputs[271]);
    assign layer0_outputs[485] = ~(inputs[166]);
    assign layer0_outputs[486] = ~(inputs[279]) | (inputs[183]);
    assign layer0_outputs[487] = inputs[97];
    assign layer0_outputs[488] = (inputs[390]) | (inputs[299]);
    assign layer0_outputs[489] = inputs[240];
    assign layer0_outputs[490] = ~((inputs[217]) | (inputs[168]));
    assign layer0_outputs[491] = inputs[9];
    assign layer0_outputs[492] = (inputs[398]) | (inputs[208]);
    assign layer0_outputs[493] = ~(inputs[201]);
    assign layer0_outputs[494] = (inputs[15]) | (inputs[113]);
    assign layer0_outputs[495] = ~(inputs[189]);
    assign layer0_outputs[496] = (inputs[147]) & ~(inputs[297]);
    assign layer0_outputs[497] = inputs[314];
    assign layer0_outputs[498] = inputs[185];
    assign layer0_outputs[499] = (inputs[62]) | (inputs[51]);
    assign layer0_outputs[500] = (inputs[151]) & ~(inputs[60]);
    assign layer0_outputs[501] = ~((inputs[152]) & (inputs[366]));
    assign layer0_outputs[502] = (inputs[10]) & ~(inputs[156]);
    assign layer0_outputs[503] = ~((inputs[306]) | (inputs[292]));
    assign layer0_outputs[504] = ~(inputs[31]);
    assign layer0_outputs[505] = inputs[335];
    assign layer0_outputs[506] = ~(inputs[302]) | (inputs[363]);
    assign layer0_outputs[507] = (inputs[42]) ^ (inputs[190]);
    assign layer0_outputs[508] = ~((inputs[233]) | (inputs[149]));
    assign layer0_outputs[509] = ~(inputs[313]) | (inputs[176]);
    assign layer0_outputs[510] = ~(inputs[172]) | (inputs[246]);
    assign layer0_outputs[511] = inputs[183];
    assign layer0_outputs[512] = ~(inputs[399]) | (inputs[373]);
    assign layer0_outputs[513] = ~(inputs[108]);
    assign layer0_outputs[514] = ~((inputs[147]) ^ (inputs[241]));
    assign layer0_outputs[515] = ~(inputs[324]) | (inputs[160]);
    assign layer0_outputs[516] = inputs[116];
    assign layer0_outputs[517] = ~((inputs[108]) | (inputs[122]));
    assign layer0_outputs[518] = ~((inputs[212]) | (inputs[105]));
    assign layer0_outputs[519] = ~(inputs[306]);
    assign layer0_outputs[520] = (inputs[236]) & ~(inputs[208]);
    assign layer0_outputs[521] = ~(inputs[50]) | (inputs[126]);
    assign layer0_outputs[522] = (inputs[399]) | (inputs[290]);
    assign layer0_outputs[523] = (inputs[146]) & ~(inputs[259]);
    assign layer0_outputs[524] = ~(inputs[13]) | (inputs[61]);
    assign layer0_outputs[525] = inputs[302];
    assign layer0_outputs[526] = ~(inputs[212]) | (inputs[294]);
    assign layer0_outputs[527] = inputs[182];
    assign layer0_outputs[528] = (inputs[349]) & ~(inputs[224]);
    assign layer0_outputs[529] = ~(inputs[52]);
    assign layer0_outputs[530] = ~(inputs[353]) | (inputs[84]);
    assign layer0_outputs[531] = inputs[192];
    assign layer0_outputs[532] = inputs[314];
    assign layer0_outputs[533] = (inputs[164]) & ~(inputs[6]);
    assign layer0_outputs[534] = (inputs[359]) ^ (inputs[84]);
    assign layer0_outputs[535] = ~((inputs[11]) | (inputs[63]));
    assign layer0_outputs[536] = (inputs[43]) ^ (inputs[127]);
    assign layer0_outputs[537] = (inputs[46]) & (inputs[326]);
    assign layer0_outputs[538] = ~(inputs[35]) | (inputs[342]);
    assign layer0_outputs[539] = (inputs[144]) & ~(inputs[399]);
    assign layer0_outputs[540] = (inputs[89]) & (inputs[329]);
    assign layer0_outputs[541] = ~(inputs[231]) | (inputs[398]);
    assign layer0_outputs[542] = (inputs[361]) | (inputs[399]);
    assign layer0_outputs[543] = ~((inputs[300]) | (inputs[292]));
    assign layer0_outputs[544] = ~((inputs[85]) | (inputs[242]));
    assign layer0_outputs[545] = inputs[250];
    assign layer0_outputs[546] = ~(inputs[32]);
    assign layer0_outputs[547] = ~(inputs[148]) | (inputs[64]);
    assign layer0_outputs[548] = ~((inputs[302]) ^ (inputs[240]));
    assign layer0_outputs[549] = inputs[194];
    assign layer0_outputs[550] = ~(inputs[176]) | (inputs[357]);
    assign layer0_outputs[551] = ~((inputs[345]) | (inputs[315]));
    assign layer0_outputs[552] = ~(inputs[376]);
    assign layer0_outputs[553] = ~((inputs[341]) ^ (inputs[168]));
    assign layer0_outputs[554] = (inputs[209]) | (inputs[80]);
    assign layer0_outputs[555] = ~((inputs[123]) ^ (inputs[314]));
    assign layer0_outputs[556] = ~(inputs[146]) | (inputs[277]);
    assign layer0_outputs[557] = (inputs[320]) | (inputs[273]);
    assign layer0_outputs[558] = ~((inputs[58]) | (inputs[24]));
    assign layer0_outputs[559] = ~(inputs[127]);
    assign layer0_outputs[560] = ~(inputs[389]);
    assign layer0_outputs[561] = ~((inputs[284]) ^ (inputs[380]));
    assign layer0_outputs[562] = ~((inputs[134]) | (inputs[249]));
    assign layer0_outputs[563] = (inputs[392]) & ~(inputs[365]);
    assign layer0_outputs[564] = ~((inputs[367]) & (inputs[86]));
    assign layer0_outputs[565] = (inputs[28]) & ~(inputs[257]);
    assign layer0_outputs[566] = (inputs[100]) ^ (inputs[351]);
    assign layer0_outputs[567] = ~(inputs[17]) | (inputs[118]);
    assign layer0_outputs[568] = ~((inputs[208]) | (inputs[116]));
    assign layer0_outputs[569] = ~(inputs[274]) | (inputs[380]);
    assign layer0_outputs[570] = ~((inputs[31]) | (inputs[23]));
    assign layer0_outputs[571] = (inputs[332]) ^ (inputs[181]);
    assign layer0_outputs[572] = ~((inputs[197]) | (inputs[199]));
    assign layer0_outputs[573] = ~(inputs[202]);
    assign layer0_outputs[574] = ~(inputs[307]) | (inputs[109]);
    assign layer0_outputs[575] = (inputs[349]) & ~(inputs[194]);
    assign layer0_outputs[576] = (inputs[170]) & ~(inputs[44]);
    assign layer0_outputs[577] = (inputs[268]) ^ (inputs[337]);
    assign layer0_outputs[578] = ~((inputs[387]) | (inputs[383]));
    assign layer0_outputs[579] = (inputs[149]) & ~(inputs[23]);
    assign layer0_outputs[580] = (inputs[17]) & ~(inputs[15]);
    assign layer0_outputs[581] = (inputs[307]) & (inputs[330]);
    assign layer0_outputs[582] = inputs[257];
    assign layer0_outputs[583] = inputs[385];
    assign layer0_outputs[584] = inputs[184];
    assign layer0_outputs[585] = (inputs[94]) & ~(inputs[19]);
    assign layer0_outputs[586] = ~(inputs[174]) | (inputs[261]);
    assign layer0_outputs[587] = (inputs[251]) & ~(inputs[388]);
    assign layer0_outputs[588] = ~((inputs[327]) | (inputs[323]));
    assign layer0_outputs[589] = ~(inputs[195]) | (inputs[323]);
    assign layer0_outputs[590] = ~(inputs[241]);
    assign layer0_outputs[591] = ~(inputs[14]);
    assign layer0_outputs[592] = ~((inputs[32]) | (inputs[157]));
    assign layer0_outputs[593] = inputs[226];
    assign layer0_outputs[594] = (inputs[55]) ^ (inputs[274]);
    assign layer0_outputs[595] = ~((inputs[196]) ^ (inputs[295]));
    assign layer0_outputs[596] = inputs[134];
    assign layer0_outputs[597] = ~(inputs[356]) | (inputs[70]);
    assign layer0_outputs[598] = (inputs[234]) | (inputs[26]);
    assign layer0_outputs[599] = (inputs[254]) | (inputs[180]);
    assign layer0_outputs[600] = ~(inputs[372]);
    assign layer0_outputs[601] = ~(inputs[321]);
    assign layer0_outputs[602] = (inputs[371]) & ~(inputs[21]);
    assign layer0_outputs[603] = ~(inputs[240]);
    assign layer0_outputs[604] = ~(inputs[200]) | (inputs[139]);
    assign layer0_outputs[605] = (inputs[275]) | (inputs[202]);
    assign layer0_outputs[606] = ~(inputs[95]) | (inputs[183]);
    assign layer0_outputs[607] = ~((inputs[192]) ^ (inputs[196]));
    assign layer0_outputs[608] = ~((inputs[258]) ^ (inputs[291]));
    assign layer0_outputs[609] = ~(inputs[198]);
    assign layer0_outputs[610] = ~(inputs[247]) | (inputs[392]);
    assign layer0_outputs[611] = (inputs[368]) ^ (inputs[99]);
    assign layer0_outputs[612] = (inputs[381]) | (inputs[260]);
    assign layer0_outputs[613] = ~(inputs[48]);
    assign layer0_outputs[614] = inputs[391];
    assign layer0_outputs[615] = (inputs[376]) | (inputs[378]);
    assign layer0_outputs[616] = inputs[107];
    assign layer0_outputs[617] = (inputs[135]) ^ (inputs[41]);
    assign layer0_outputs[618] = 1'b1;
    assign layer0_outputs[619] = ~(inputs[291]);
    assign layer0_outputs[620] = ~((inputs[248]) & (inputs[305]));
    assign layer0_outputs[621] = ~((inputs[185]) | (inputs[343]));
    assign layer0_outputs[622] = ~(inputs[47]) | (inputs[278]);
    assign layer0_outputs[623] = (inputs[40]) | (inputs[391]);
    assign layer0_outputs[624] = ~((inputs[16]) ^ (inputs[71]));
    assign layer0_outputs[625] = ~(inputs[268]);
    assign layer0_outputs[626] = inputs[147];
    assign layer0_outputs[627] = ~((inputs[252]) | (inputs[117]));
    assign layer0_outputs[628] = ~(inputs[12]);
    assign layer0_outputs[629] = (inputs[336]) | (inputs[211]);
    assign layer0_outputs[630] = (inputs[117]) ^ (inputs[315]);
    assign layer0_outputs[631] = ~(inputs[49]) | (inputs[145]);
    assign layer0_outputs[632] = ~(inputs[12]) | (inputs[123]);
    assign layer0_outputs[633] = ~(inputs[190]);
    assign layer0_outputs[634] = (inputs[98]) & ~(inputs[80]);
    assign layer0_outputs[635] = ~((inputs[222]) | (inputs[284]));
    assign layer0_outputs[636] = (inputs[132]) & ~(inputs[314]);
    assign layer0_outputs[637] = ~(inputs[72]);
    assign layer0_outputs[638] = ~((inputs[357]) ^ (inputs[298]));
    assign layer0_outputs[639] = (inputs[80]) ^ (inputs[41]);
    assign layer0_outputs[640] = inputs[284];
    assign layer0_outputs[641] = ~(inputs[131]) | (inputs[105]);
    assign layer0_outputs[642] = ~((inputs[229]) | (inputs[121]));
    assign layer0_outputs[643] = inputs[225];
    assign layer0_outputs[644] = inputs[210];
    assign layer0_outputs[645] = ~(inputs[165]);
    assign layer0_outputs[646] = ~(inputs[156]);
    assign layer0_outputs[647] = inputs[274];
    assign layer0_outputs[648] = ~((inputs[319]) | (inputs[384]));
    assign layer0_outputs[649] = ~((inputs[359]) | (inputs[46]));
    assign layer0_outputs[650] = inputs[366];
    assign layer0_outputs[651] = (inputs[279]) | (inputs[335]);
    assign layer0_outputs[652] = ~((inputs[65]) | (inputs[51]));
    assign layer0_outputs[653] = (inputs[127]) ^ (inputs[103]);
    assign layer0_outputs[654] = inputs[162];
    assign layer0_outputs[655] = ~(inputs[370]);
    assign layer0_outputs[656] = ~((inputs[297]) | (inputs[391]));
    assign layer0_outputs[657] = inputs[124];
    assign layer0_outputs[658] = ~(inputs[118]);
    assign layer0_outputs[659] = inputs[354];
    assign layer0_outputs[660] = ~(inputs[172]);
    assign layer0_outputs[661] = ~((inputs[145]) & (inputs[55]));
    assign layer0_outputs[662] = ~(inputs[302]);
    assign layer0_outputs[663] = ~(inputs[83]);
    assign layer0_outputs[664] = (inputs[356]) | (inputs[365]);
    assign layer0_outputs[665] = ~((inputs[81]) | (inputs[113]));
    assign layer0_outputs[666] = ~(inputs[140]);
    assign layer0_outputs[667] = ~(inputs[327]) | (inputs[249]);
    assign layer0_outputs[668] = (inputs[349]) & ~(inputs[62]);
    assign layer0_outputs[669] = (inputs[336]) | (inputs[337]);
    assign layer0_outputs[670] = ~((inputs[135]) & (inputs[99]));
    assign layer0_outputs[671] = (inputs[283]) | (inputs[235]);
    assign layer0_outputs[672] = ~((inputs[358]) | (inputs[380]));
    assign layer0_outputs[673] = (inputs[83]) | (inputs[355]);
    assign layer0_outputs[674] = (inputs[289]) & ~(inputs[163]);
    assign layer0_outputs[675] = (inputs[107]) | (inputs[67]);
    assign layer0_outputs[676] = (inputs[3]) | (inputs[347]);
    assign layer0_outputs[677] = (inputs[262]) & ~(inputs[378]);
    assign layer0_outputs[678] = 1'b1;
    assign layer0_outputs[679] = (inputs[279]) | (inputs[132]);
    assign layer0_outputs[680] = ~(inputs[202]) | (inputs[262]);
    assign layer0_outputs[681] = (inputs[325]) | (inputs[281]);
    assign layer0_outputs[682] = (inputs[145]) & ~(inputs[219]);
    assign layer0_outputs[683] = ~(inputs[154]);
    assign layer0_outputs[684] = ~((inputs[143]) | (inputs[28]));
    assign layer0_outputs[685] = ~((inputs[174]) & (inputs[117]));
    assign layer0_outputs[686] = (inputs[97]) | (inputs[138]);
    assign layer0_outputs[687] = ~((inputs[4]) ^ (inputs[40]));
    assign layer0_outputs[688] = inputs[383];
    assign layer0_outputs[689] = ~(inputs[318]) | (inputs[82]);
    assign layer0_outputs[690] = inputs[325];
    assign layer0_outputs[691] = (inputs[215]) & ~(inputs[367]);
    assign layer0_outputs[692] = (inputs[313]) & (inputs[362]);
    assign layer0_outputs[693] = ~(inputs[244]);
    assign layer0_outputs[694] = ~(inputs[6]);
    assign layer0_outputs[695] = ~(inputs[337]) | (inputs[27]);
    assign layer0_outputs[696] = ~((inputs[355]) | (inputs[338]));
    assign layer0_outputs[697] = ~((inputs[149]) | (inputs[169]));
    assign layer0_outputs[698] = (inputs[58]) | (inputs[160]);
    assign layer0_outputs[699] = (inputs[322]) | (inputs[316]);
    assign layer0_outputs[700] = (inputs[387]) & ~(inputs[296]);
    assign layer0_outputs[701] = ~((inputs[296]) | (inputs[62]));
    assign layer0_outputs[702] = (inputs[378]) | (inputs[174]);
    assign layer0_outputs[703] = ~(inputs[315]);
    assign layer0_outputs[704] = ~((inputs[5]) | (inputs[25]));
    assign layer0_outputs[705] = (inputs[332]) | (inputs[352]);
    assign layer0_outputs[706] = inputs[171];
    assign layer0_outputs[707] = (inputs[295]) | (inputs[326]);
    assign layer0_outputs[708] = (inputs[138]) | (inputs[20]);
    assign layer0_outputs[709] = ~(inputs[245]);
    assign layer0_outputs[710] = ~(inputs[41]);
    assign layer0_outputs[711] = (inputs[215]) & ~(inputs[67]);
    assign layer0_outputs[712] = ~((inputs[398]) ^ (inputs[151]));
    assign layer0_outputs[713] = (inputs[314]) & (inputs[350]);
    assign layer0_outputs[714] = ~(inputs[166]);
    assign layer0_outputs[715] = inputs[42];
    assign layer0_outputs[716] = (inputs[69]) ^ (inputs[144]);
    assign layer0_outputs[717] = (inputs[332]) & ~(inputs[203]);
    assign layer0_outputs[718] = inputs[351];
    assign layer0_outputs[719] = (inputs[97]) | (inputs[27]);
    assign layer0_outputs[720] = ~((inputs[241]) ^ (inputs[264]));
    assign layer0_outputs[721] = ~(inputs[9]) | (inputs[72]);
    assign layer0_outputs[722] = inputs[243];
    assign layer0_outputs[723] = (inputs[308]) & ~(inputs[273]);
    assign layer0_outputs[724] = inputs[133];
    assign layer0_outputs[725] = ~((inputs[158]) | (inputs[378]));
    assign layer0_outputs[726] = (inputs[10]) & ~(inputs[3]);
    assign layer0_outputs[727] = (inputs[174]) & ~(inputs[51]);
    assign layer0_outputs[728] = ~((inputs[151]) ^ (inputs[111]));
    assign layer0_outputs[729] = ~(inputs[132]) | (inputs[217]);
    assign layer0_outputs[730] = inputs[35];
    assign layer0_outputs[731] = ~((inputs[288]) | (inputs[227]));
    assign layer0_outputs[732] = ~(inputs[248]) | (inputs[184]);
    assign layer0_outputs[733] = (inputs[55]) ^ (inputs[153]);
    assign layer0_outputs[734] = (inputs[168]) | (inputs[370]);
    assign layer0_outputs[735] = inputs[333];
    assign layer0_outputs[736] = ~(inputs[387]);
    assign layer0_outputs[737] = ~(inputs[265]) | (inputs[86]);
    assign layer0_outputs[738] = (inputs[107]) | (inputs[222]);
    assign layer0_outputs[739] = ~(inputs[264]);
    assign layer0_outputs[740] = (inputs[212]) & ~(inputs[364]);
    assign layer0_outputs[741] = (inputs[95]) & ~(inputs[396]);
    assign layer0_outputs[742] = ~(inputs[358]);
    assign layer0_outputs[743] = inputs[103];
    assign layer0_outputs[744] = ~(inputs[366]);
    assign layer0_outputs[745] = ~((inputs[140]) | (inputs[221]));
    assign layer0_outputs[746] = (inputs[86]) ^ (inputs[66]);
    assign layer0_outputs[747] = (inputs[306]) & ~(inputs[118]);
    assign layer0_outputs[748] = ~(inputs[137]);
    assign layer0_outputs[749] = ~(inputs[151]) | (inputs[217]);
    assign layer0_outputs[750] = ~(inputs[115]);
    assign layer0_outputs[751] = ~(inputs[13]);
    assign layer0_outputs[752] = inputs[211];
    assign layer0_outputs[753] = (inputs[324]) & ~(inputs[357]);
    assign layer0_outputs[754] = (inputs[199]) | (inputs[18]);
    assign layer0_outputs[755] = ~(inputs[288]);
    assign layer0_outputs[756] = inputs[91];
    assign layer0_outputs[757] = ~((inputs[209]) | (inputs[157]));
    assign layer0_outputs[758] = ~((inputs[230]) | (inputs[4]));
    assign layer0_outputs[759] = (inputs[131]) & ~(inputs[219]);
    assign layer0_outputs[760] = ~((inputs[256]) ^ (inputs[364]));
    assign layer0_outputs[761] = ~((inputs[280]) | (inputs[10]));
    assign layer0_outputs[762] = 1'b1;
    assign layer0_outputs[763] = ~(inputs[368]);
    assign layer0_outputs[764] = ~((inputs[198]) | (inputs[0]));
    assign layer0_outputs[765] = (inputs[307]) & ~(inputs[170]);
    assign layer0_outputs[766] = (inputs[98]) | (inputs[74]);
    assign layer0_outputs[767] = (inputs[146]) | (inputs[216]);
    assign layer0_outputs[768] = inputs[126];
    assign layer0_outputs[769] = inputs[116];
    assign layer0_outputs[770] = (inputs[201]) | (inputs[115]);
    assign layer0_outputs[771] = (inputs[268]) & ~(inputs[298]);
    assign layer0_outputs[772] = inputs[106];
    assign layer0_outputs[773] = inputs[217];
    assign layer0_outputs[774] = ~((inputs[127]) | (inputs[167]));
    assign layer0_outputs[775] = (inputs[384]) | (inputs[209]);
    assign layer0_outputs[776] = (inputs[21]) ^ (inputs[316]);
    assign layer0_outputs[777] = ~((inputs[112]) & (inputs[188]));
    assign layer0_outputs[778] = ~((inputs[359]) | (inputs[40]));
    assign layer0_outputs[779] = inputs[250];
    assign layer0_outputs[780] = ~(inputs[301]);
    assign layer0_outputs[781] = (inputs[53]) & (inputs[333]);
    assign layer0_outputs[782] = (inputs[4]) | (inputs[338]);
    assign layer0_outputs[783] = (inputs[240]) | (inputs[115]);
    assign layer0_outputs[784] = ~((inputs[171]) | (inputs[45]));
    assign layer0_outputs[785] = inputs[182];
    assign layer0_outputs[786] = ~(inputs[223]);
    assign layer0_outputs[787] = (inputs[319]) & ~(inputs[161]);
    assign layer0_outputs[788] = ~(inputs[312]);
    assign layer0_outputs[789] = (inputs[380]) ^ (inputs[341]);
    assign layer0_outputs[790] = inputs[144];
    assign layer0_outputs[791] = ~(inputs[389]);
    assign layer0_outputs[792] = inputs[282];
    assign layer0_outputs[793] = ~(inputs[247]);
    assign layer0_outputs[794] = ~((inputs[343]) | (inputs[225]));
    assign layer0_outputs[795] = (inputs[14]) & ~(inputs[382]);
    assign layer0_outputs[796] = inputs[93];
    assign layer0_outputs[797] = ~(inputs[105]);
    assign layer0_outputs[798] = ~((inputs[395]) | (inputs[310]));
    assign layer0_outputs[799] = (inputs[25]) & ~(inputs[172]);
    assign layer0_outputs[800] = ~((inputs[43]) ^ (inputs[100]));
    assign layer0_outputs[801] = ~((inputs[19]) | (inputs[336]));
    assign layer0_outputs[802] = inputs[305];
    assign layer0_outputs[803] = ~(inputs[213]);
    assign layer0_outputs[804] = ~(inputs[122]);
    assign layer0_outputs[805] = inputs[26];
    assign layer0_outputs[806] = (inputs[99]) | (inputs[241]);
    assign layer0_outputs[807] = (inputs[324]) | (inputs[280]);
    assign layer0_outputs[808] = ~(inputs[111]) | (inputs[294]);
    assign layer0_outputs[809] = inputs[72];
    assign layer0_outputs[810] = (inputs[292]) ^ (inputs[187]);
    assign layer0_outputs[811] = inputs[111];
    assign layer0_outputs[812] = (inputs[103]) | (inputs[327]);
    assign layer0_outputs[813] = ~(inputs[174]) | (inputs[349]);
    assign layer0_outputs[814] = ~((inputs[174]) & (inputs[95]));
    assign layer0_outputs[815] = (inputs[395]) | (inputs[21]);
    assign layer0_outputs[816] = ~(inputs[172]);
    assign layer0_outputs[817] = (inputs[195]) | (inputs[323]);
    assign layer0_outputs[818] = ~(inputs[306]);
    assign layer0_outputs[819] = (inputs[39]) | (inputs[195]);
    assign layer0_outputs[820] = inputs[181];
    assign layer0_outputs[821] = inputs[1];
    assign layer0_outputs[822] = (inputs[75]) & (inputs[373]);
    assign layer0_outputs[823] = ~(inputs[300]);
    assign layer0_outputs[824] = (inputs[165]) | (inputs[117]);
    assign layer0_outputs[825] = inputs[168];
    assign layer0_outputs[826] = (inputs[250]) | (inputs[42]);
    assign layer0_outputs[827] = inputs[167];
    assign layer0_outputs[828] = ~((inputs[252]) | (inputs[215]));
    assign layer0_outputs[829] = (inputs[168]) | (inputs[373]);
    assign layer0_outputs[830] = inputs[251];
    assign layer0_outputs[831] = ~(inputs[196]);
    assign layer0_outputs[832] = ~((inputs[365]) & (inputs[283]));
    assign layer0_outputs[833] = ~((inputs[15]) ^ (inputs[158]));
    assign layer0_outputs[834] = ~((inputs[97]) | (inputs[314]));
    assign layer0_outputs[835] = 1'b0;
    assign layer0_outputs[836] = inputs[55];
    assign layer0_outputs[837] = ~(inputs[5]) | (inputs[376]);
    assign layer0_outputs[838] = (inputs[40]) | (inputs[88]);
    assign layer0_outputs[839] = ~((inputs[312]) | (inputs[293]));
    assign layer0_outputs[840] = ~(inputs[283]);
    assign layer0_outputs[841] = 1'b1;
    assign layer0_outputs[842] = ~((inputs[220]) | (inputs[126]));
    assign layer0_outputs[843] = (inputs[187]) & ~(inputs[337]);
    assign layer0_outputs[844] = ~((inputs[145]) | (inputs[253]));
    assign layer0_outputs[845] = (inputs[119]) & ~(inputs[178]);
    assign layer0_outputs[846] = inputs[102];
    assign layer0_outputs[847] = ~(inputs[202]) | (inputs[240]);
    assign layer0_outputs[848] = ~(inputs[390]) | (inputs[175]);
    assign layer0_outputs[849] = (inputs[281]) | (inputs[34]);
    assign layer0_outputs[850] = (inputs[28]) & ~(inputs[17]);
    assign layer0_outputs[851] = inputs[168];
    assign layer0_outputs[852] = (inputs[285]) & ~(inputs[139]);
    assign layer0_outputs[853] = (inputs[16]) ^ (inputs[26]);
    assign layer0_outputs[854] = (inputs[276]) & ~(inputs[398]);
    assign layer0_outputs[855] = inputs[370];
    assign layer0_outputs[856] = inputs[267];
    assign layer0_outputs[857] = (inputs[371]) | (inputs[284]);
    assign layer0_outputs[858] = (inputs[304]) & ~(inputs[112]);
    assign layer0_outputs[859] = ~((inputs[110]) & (inputs[288]));
    assign layer0_outputs[860] = (inputs[375]) & ~(inputs[27]);
    assign layer0_outputs[861] = inputs[164];
    assign layer0_outputs[862] = (inputs[184]) | (inputs[242]);
    assign layer0_outputs[863] = inputs[114];
    assign layer0_outputs[864] = inputs[204];
    assign layer0_outputs[865] = ~((inputs[99]) ^ (inputs[22]));
    assign layer0_outputs[866] = inputs[176];
    assign layer0_outputs[867] = ~((inputs[140]) ^ (inputs[356]));
    assign layer0_outputs[868] = inputs[260];
    assign layer0_outputs[869] = ~(inputs[73]) | (inputs[274]);
    assign layer0_outputs[870] = (inputs[243]) & (inputs[389]);
    assign layer0_outputs[871] = ~((inputs[27]) ^ (inputs[365]));
    assign layer0_outputs[872] = ~(inputs[10]);
    assign layer0_outputs[873] = inputs[29];
    assign layer0_outputs[874] = ~(inputs[87]);
    assign layer0_outputs[875] = ~((inputs[294]) & (inputs[270]));
    assign layer0_outputs[876] = inputs[296];
    assign layer0_outputs[877] = ~(inputs[367]);
    assign layer0_outputs[878] = (inputs[204]) & ~(inputs[101]);
    assign layer0_outputs[879] = ~(inputs[204]);
    assign layer0_outputs[880] = ~(inputs[34]);
    assign layer0_outputs[881] = (inputs[258]) | (inputs[254]);
    assign layer0_outputs[882] = inputs[22];
    assign layer0_outputs[883] = (inputs[386]) & (inputs[207]);
    assign layer0_outputs[884] = ~((inputs[306]) | (inputs[257]));
    assign layer0_outputs[885] = (inputs[237]) & ~(inputs[246]);
    assign layer0_outputs[886] = ~((inputs[73]) ^ (inputs[75]));
    assign layer0_outputs[887] = (inputs[52]) & (inputs[75]);
    assign layer0_outputs[888] = inputs[348];
    assign layer0_outputs[889] = inputs[395];
    assign layer0_outputs[890] = inputs[303];
    assign layer0_outputs[891] = ~((inputs[307]) | (inputs[122]));
    assign layer0_outputs[892] = inputs[72];
    assign layer0_outputs[893] = ~(inputs[334]);
    assign layer0_outputs[894] = inputs[388];
    assign layer0_outputs[895] = ~((inputs[13]) | (inputs[186]));
    assign layer0_outputs[896] = ~(inputs[92]);
    assign layer0_outputs[897] = (inputs[27]) | (inputs[377]);
    assign layer0_outputs[898] = ~(inputs[59]);
    assign layer0_outputs[899] = inputs[131];
    assign layer0_outputs[900] = (inputs[40]) & ~(inputs[95]);
    assign layer0_outputs[901] = (inputs[103]) & (inputs[328]);
    assign layer0_outputs[902] = ~((inputs[362]) ^ (inputs[95]));
    assign layer0_outputs[903] = inputs[248];
    assign layer0_outputs[904] = ~((inputs[148]) ^ (inputs[158]));
    assign layer0_outputs[905] = inputs[366];
    assign layer0_outputs[906] = ~(inputs[25]) | (inputs[217]);
    assign layer0_outputs[907] = ~(inputs[229]) | (inputs[60]);
    assign layer0_outputs[908] = (inputs[339]) ^ (inputs[165]);
    assign layer0_outputs[909] = inputs[137];
    assign layer0_outputs[910] = inputs[368];
    assign layer0_outputs[911] = ~(inputs[13]);
    assign layer0_outputs[912] = (inputs[31]) | (inputs[380]);
    assign layer0_outputs[913] = inputs[156];
    assign layer0_outputs[914] = ~((inputs[250]) & (inputs[322]));
    assign layer0_outputs[915] = (inputs[384]) | (inputs[243]);
    assign layer0_outputs[916] = ~(inputs[321]);
    assign layer0_outputs[917] = inputs[349];
    assign layer0_outputs[918] = 1'b0;
    assign layer0_outputs[919] = ~((inputs[282]) ^ (inputs[16]));
    assign layer0_outputs[920] = ~(inputs[17]);
    assign layer0_outputs[921] = (inputs[151]) | (inputs[67]);
    assign layer0_outputs[922] = ~((inputs[397]) | (inputs[396]));
    assign layer0_outputs[923] = ~((inputs[393]) | (inputs[395]));
    assign layer0_outputs[924] = ~(inputs[358]);
    assign layer0_outputs[925] = (inputs[221]) ^ (inputs[211]);
    assign layer0_outputs[926] = (inputs[54]) | (inputs[260]);
    assign layer0_outputs[927] = inputs[169];
    assign layer0_outputs[928] = ~(inputs[229]);
    assign layer0_outputs[929] = inputs[291];
    assign layer0_outputs[930] = inputs[183];
    assign layer0_outputs[931] = ~(inputs[41]) | (inputs[180]);
    assign layer0_outputs[932] = ~((inputs[213]) ^ (inputs[211]));
    assign layer0_outputs[933] = ~((inputs[244]) ^ (inputs[344]));
    assign layer0_outputs[934] = ~(inputs[375]);
    assign layer0_outputs[935] = inputs[281];
    assign layer0_outputs[936] = inputs[114];
    assign layer0_outputs[937] = inputs[234];
    assign layer0_outputs[938] = inputs[128];
    assign layer0_outputs[939] = ~(inputs[266]) | (inputs[320]);
    assign layer0_outputs[940] = ~(inputs[335]) | (inputs[85]);
    assign layer0_outputs[941] = (inputs[27]) & ~(inputs[15]);
    assign layer0_outputs[942] = ~(inputs[230]);
    assign layer0_outputs[943] = (inputs[3]) | (inputs[280]);
    assign layer0_outputs[944] = inputs[293];
    assign layer0_outputs[945] = ~(inputs[128]);
    assign layer0_outputs[946] = ~((inputs[66]) | (inputs[44]));
    assign layer0_outputs[947] = (inputs[193]) ^ (inputs[256]);
    assign layer0_outputs[948] = ~(inputs[85]);
    assign layer0_outputs[949] = ~((inputs[369]) | (inputs[140]));
    assign layer0_outputs[950] = inputs[319];
    assign layer0_outputs[951] = (inputs[133]) & ~(inputs[334]);
    assign layer0_outputs[952] = inputs[113];
    assign layer0_outputs[953] = ~((inputs[82]) & (inputs[91]));
    assign layer0_outputs[954] = ~((inputs[149]) ^ (inputs[106]));
    assign layer0_outputs[955] = (inputs[71]) | (inputs[190]);
    assign layer0_outputs[956] = ~((inputs[395]) ^ (inputs[295]));
    assign layer0_outputs[957] = ~(inputs[186]) | (inputs[158]);
    assign layer0_outputs[958] = (inputs[83]) & ~(inputs[198]);
    assign layer0_outputs[959] = (inputs[276]) & ~(inputs[152]);
    assign layer0_outputs[960] = ~((inputs[151]) ^ (inputs[201]));
    assign layer0_outputs[961] = inputs[192];
    assign layer0_outputs[962] = (inputs[149]) ^ (inputs[283]);
    assign layer0_outputs[963] = ~(inputs[22]);
    assign layer0_outputs[964] = inputs[143];
    assign layer0_outputs[965] = inputs[264];
    assign layer0_outputs[966] = ~(inputs[267]) | (inputs[79]);
    assign layer0_outputs[967] = ~(inputs[162]);
    assign layer0_outputs[968] = (inputs[349]) ^ (inputs[373]);
    assign layer0_outputs[969] = ~(inputs[68]) | (inputs[159]);
    assign layer0_outputs[970] = ~((inputs[194]) | (inputs[201]));
    assign layer0_outputs[971] = ~(inputs[70]);
    assign layer0_outputs[972] = (inputs[114]) | (inputs[99]);
    assign layer0_outputs[973] = inputs[374];
    assign layer0_outputs[974] = ~(inputs[85]);
    assign layer0_outputs[975] = ~(inputs[334]) | (inputs[350]);
    assign layer0_outputs[976] = inputs[157];
    assign layer0_outputs[977] = inputs[184];
    assign layer0_outputs[978] = ~(inputs[34]);
    assign layer0_outputs[979] = inputs[359];
    assign layer0_outputs[980] = (inputs[348]) & ~(inputs[173]);
    assign layer0_outputs[981] = ~(inputs[262]);
    assign layer0_outputs[982] = inputs[154];
    assign layer0_outputs[983] = (inputs[133]) & ~(inputs[304]);
    assign layer0_outputs[984] = inputs[12];
    assign layer0_outputs[985] = inputs[207];
    assign layer0_outputs[986] = ~((inputs[264]) | (inputs[237]));
    assign layer0_outputs[987] = ~((inputs[37]) | (inputs[15]));
    assign layer0_outputs[988] = ~((inputs[295]) | (inputs[242]));
    assign layer0_outputs[989] = (inputs[32]) & (inputs[57]);
    assign layer0_outputs[990] = ~(inputs[120]) | (inputs[295]);
    assign layer0_outputs[991] = inputs[227];
    assign layer0_outputs[992] = ~(inputs[11]) | (inputs[381]);
    assign layer0_outputs[993] = ~((inputs[25]) ^ (inputs[216]));
    assign layer0_outputs[994] = ~(inputs[389]) | (inputs[89]);
    assign layer0_outputs[995] = (inputs[298]) | (inputs[316]);
    assign layer0_outputs[996] = (inputs[71]) & (inputs[167]);
    assign layer0_outputs[997] = ~(inputs[17]) | (inputs[300]);
    assign layer0_outputs[998] = (inputs[356]) ^ (inputs[217]);
    assign layer0_outputs[999] = ~(inputs[245]) | (inputs[100]);
    assign layer0_outputs[1000] = 1'b1;
    assign layer0_outputs[1001] = ~((inputs[121]) ^ (inputs[28]));
    assign layer0_outputs[1002] = ~(inputs[142]);
    assign layer0_outputs[1003] = ~((inputs[101]) | (inputs[387]));
    assign layer0_outputs[1004] = (inputs[136]) | (inputs[235]);
    assign layer0_outputs[1005] = ~(inputs[139]);
    assign layer0_outputs[1006] = (inputs[234]) & ~(inputs[92]);
    assign layer0_outputs[1007] = (inputs[141]) & (inputs[258]);
    assign layer0_outputs[1008] = ~((inputs[34]) | (inputs[132]));
    assign layer0_outputs[1009] = ~(inputs[251]);
    assign layer0_outputs[1010] = ~((inputs[394]) | (inputs[305]));
    assign layer0_outputs[1011] = ~((inputs[259]) ^ (inputs[277]));
    assign layer0_outputs[1012] = inputs[322];
    assign layer0_outputs[1013] = inputs[150];
    assign layer0_outputs[1014] = (inputs[249]) ^ (inputs[210]);
    assign layer0_outputs[1015] = ~(inputs[285]);
    assign layer0_outputs[1016] = ~(inputs[321]) | (inputs[141]);
    assign layer0_outputs[1017] = (inputs[336]) | (inputs[336]);
    assign layer0_outputs[1018] = ~(inputs[219]);
    assign layer0_outputs[1019] = (inputs[363]) | (inputs[341]);
    assign layer0_outputs[1020] = ~(inputs[173]);
    assign layer0_outputs[1021] = ~(inputs[354]) | (inputs[20]);
    assign layer0_outputs[1022] = (inputs[310]) ^ (inputs[356]);
    assign layer0_outputs[1023] = inputs[149];
    assign layer0_outputs[1024] = ~((inputs[345]) | (inputs[279]));
    assign layer0_outputs[1025] = ~(inputs[84]);
    assign layer0_outputs[1026] = inputs[367];
    assign layer0_outputs[1027] = (inputs[37]) | (inputs[317]);
    assign layer0_outputs[1028] = (inputs[141]) | (inputs[392]);
    assign layer0_outputs[1029] = inputs[117];
    assign layer0_outputs[1030] = (inputs[388]) & ~(inputs[54]);
    assign layer0_outputs[1031] = (inputs[266]) | (inputs[361]);
    assign layer0_outputs[1032] = inputs[153];
    assign layer0_outputs[1033] = (inputs[82]) | (inputs[80]);
    assign layer0_outputs[1034] = ~(inputs[331]);
    assign layer0_outputs[1035] = (inputs[93]) & ~(inputs[316]);
    assign layer0_outputs[1036] = (inputs[339]) ^ (inputs[216]);
    assign layer0_outputs[1037] = (inputs[89]) ^ (inputs[360]);
    assign layer0_outputs[1038] = ~((inputs[141]) | (inputs[190]));
    assign layer0_outputs[1039] = inputs[326];
    assign layer0_outputs[1040] = ~((inputs[159]) ^ (inputs[136]));
    assign layer0_outputs[1041] = ~(inputs[269]);
    assign layer0_outputs[1042] = ~(inputs[166]) | (inputs[249]);
    assign layer0_outputs[1043] = (inputs[331]) ^ (inputs[312]);
    assign layer0_outputs[1044] = (inputs[285]) & ~(inputs[359]);
    assign layer0_outputs[1045] = ~(inputs[47]);
    assign layer0_outputs[1046] = ~(inputs[197]) | (inputs[101]);
    assign layer0_outputs[1047] = ~(inputs[68]);
    assign layer0_outputs[1048] = ~((inputs[396]) | (inputs[276]));
    assign layer0_outputs[1049] = inputs[309];
    assign layer0_outputs[1050] = ~(inputs[360]);
    assign layer0_outputs[1051] = ~(inputs[377]) | (inputs[340]);
    assign layer0_outputs[1052] = inputs[264];
    assign layer0_outputs[1053] = ~(inputs[162]);
    assign layer0_outputs[1054] = ~(inputs[91]) | (inputs[22]);
    assign layer0_outputs[1055] = ~(inputs[345]);
    assign layer0_outputs[1056] = inputs[209];
    assign layer0_outputs[1057] = ~(inputs[338]);
    assign layer0_outputs[1058] = ~((inputs[155]) ^ (inputs[2]));
    assign layer0_outputs[1059] = ~(inputs[95]) | (inputs[142]);
    assign layer0_outputs[1060] = ~(inputs[371]) | (inputs[238]);
    assign layer0_outputs[1061] = ~((inputs[96]) | (inputs[126]));
    assign layer0_outputs[1062] = (inputs[204]) ^ (inputs[294]);
    assign layer0_outputs[1063] = ~((inputs[346]) | (inputs[392]));
    assign layer0_outputs[1064] = (inputs[6]) ^ (inputs[84]);
    assign layer0_outputs[1065] = ~(inputs[272]) | (inputs[119]);
    assign layer0_outputs[1066] = ~(inputs[286]);
    assign layer0_outputs[1067] = ~((inputs[182]) | (inputs[59]));
    assign layer0_outputs[1068] = (inputs[11]) ^ (inputs[301]);
    assign layer0_outputs[1069] = ~(inputs[30]) | (inputs[264]);
    assign layer0_outputs[1070] = inputs[220];
    assign layer0_outputs[1071] = inputs[276];
    assign layer0_outputs[1072] = (inputs[156]) ^ (inputs[130]);
    assign layer0_outputs[1073] = ~(inputs[170]);
    assign layer0_outputs[1074] = (inputs[143]) & ~(inputs[344]);
    assign layer0_outputs[1075] = (inputs[245]) & ~(inputs[64]);
    assign layer0_outputs[1076] = ~(inputs[151]);
    assign layer0_outputs[1077] = (inputs[86]) & ~(inputs[298]);
    assign layer0_outputs[1078] = (inputs[70]) & ~(inputs[337]);
    assign layer0_outputs[1079] = inputs[48];
    assign layer0_outputs[1080] = ~(inputs[283]) | (inputs[116]);
    assign layer0_outputs[1081] = ~(inputs[353]) | (inputs[396]);
    assign layer0_outputs[1082] = ~(inputs[249]) | (inputs[226]);
    assign layer0_outputs[1083] = ~((inputs[136]) | (inputs[389]));
    assign layer0_outputs[1084] = (inputs[34]) & ~(inputs[180]);
    assign layer0_outputs[1085] = (inputs[142]) & ~(inputs[139]);
    assign layer0_outputs[1086] = inputs[128];
    assign layer0_outputs[1087] = ~(inputs[10]);
    assign layer0_outputs[1088] = ~((inputs[52]) | (inputs[318]));
    assign layer0_outputs[1089] = inputs[297];
    assign layer0_outputs[1090] = (inputs[301]) | (inputs[317]);
    assign layer0_outputs[1091] = inputs[184];
    assign layer0_outputs[1092] = ~(inputs[261]);
    assign layer0_outputs[1093] = ~(inputs[193]);
    assign layer0_outputs[1094] = (inputs[308]) & ~(inputs[191]);
    assign layer0_outputs[1095] = inputs[207];
    assign layer0_outputs[1096] = ~(inputs[191]);
    assign layer0_outputs[1097] = ~(inputs[145]);
    assign layer0_outputs[1098] = (inputs[32]) ^ (inputs[121]);
    assign layer0_outputs[1099] = ~(inputs[146]) | (inputs[179]);
    assign layer0_outputs[1100] = ~((inputs[33]) ^ (inputs[52]));
    assign layer0_outputs[1101] = (inputs[252]) & ~(inputs[130]);
    assign layer0_outputs[1102] = inputs[153];
    assign layer0_outputs[1103] = (inputs[381]) | (inputs[24]);
    assign layer0_outputs[1104] = ~(inputs[10]) | (inputs[303]);
    assign layer0_outputs[1105] = inputs[165];
    assign layer0_outputs[1106] = ~((inputs[195]) | (inputs[198]));
    assign layer0_outputs[1107] = inputs[365];
    assign layer0_outputs[1108] = ~(inputs[18]);
    assign layer0_outputs[1109] = (inputs[130]) & ~(inputs[317]);
    assign layer0_outputs[1110] = (inputs[161]) | (inputs[297]);
    assign layer0_outputs[1111] = 1'b0;
    assign layer0_outputs[1112] = (inputs[154]) & (inputs[210]);
    assign layer0_outputs[1113] = ~((inputs[99]) | (inputs[200]));
    assign layer0_outputs[1114] = ~(inputs[351]);
    assign layer0_outputs[1115] = inputs[11];
    assign layer0_outputs[1116] = ~(inputs[280]);
    assign layer0_outputs[1117] = ~(inputs[376]);
    assign layer0_outputs[1118] = (inputs[213]) & ~(inputs[160]);
    assign layer0_outputs[1119] = (inputs[89]) | (inputs[348]);
    assign layer0_outputs[1120] = ~((inputs[294]) ^ (inputs[332]));
    assign layer0_outputs[1121] = ~((inputs[337]) | (inputs[296]));
    assign layer0_outputs[1122] = (inputs[269]) ^ (inputs[22]);
    assign layer0_outputs[1123] = ~((inputs[26]) | (inputs[3]));
    assign layer0_outputs[1124] = inputs[0];
    assign layer0_outputs[1125] = ~(inputs[39]);
    assign layer0_outputs[1126] = (inputs[306]) & ~(inputs[132]);
    assign layer0_outputs[1127] = inputs[106];
    assign layer0_outputs[1128] = 1'b1;
    assign layer0_outputs[1129] = (inputs[171]) ^ (inputs[289]);
    assign layer0_outputs[1130] = ~((inputs[270]) ^ (inputs[289]));
    assign layer0_outputs[1131] = (inputs[159]) ^ (inputs[131]);
    assign layer0_outputs[1132] = inputs[114];
    assign layer0_outputs[1133] = ~(inputs[130]) | (inputs[101]);
    assign layer0_outputs[1134] = ~(inputs[130]) | (inputs[142]);
    assign layer0_outputs[1135] = inputs[193];
    assign layer0_outputs[1136] = ~(inputs[307]);
    assign layer0_outputs[1137] = (inputs[265]) & ~(inputs[380]);
    assign layer0_outputs[1138] = inputs[245];
    assign layer0_outputs[1139] = ~(inputs[373]);
    assign layer0_outputs[1140] = ~((inputs[333]) | (inputs[261]));
    assign layer0_outputs[1141] = ~((inputs[270]) ^ (inputs[99]));
    assign layer0_outputs[1142] = inputs[54];
    assign layer0_outputs[1143] = ~(inputs[81]);
    assign layer0_outputs[1144] = (inputs[217]) ^ (inputs[331]);
    assign layer0_outputs[1145] = ~(inputs[27]);
    assign layer0_outputs[1146] = inputs[129];
    assign layer0_outputs[1147] = ~((inputs[331]) ^ (inputs[287]));
    assign layer0_outputs[1148] = inputs[278];
    assign layer0_outputs[1149] = inputs[247];
    assign layer0_outputs[1150] = (inputs[295]) | (inputs[363]);
    assign layer0_outputs[1151] = ~(inputs[325]) | (inputs[226]);
    assign layer0_outputs[1152] = ~(inputs[358]);
    assign layer0_outputs[1153] = ~((inputs[21]) | (inputs[78]));
    assign layer0_outputs[1154] = ~((inputs[281]) | (inputs[290]));
    assign layer0_outputs[1155] = ~(inputs[121]);
    assign layer0_outputs[1156] = ~((inputs[174]) ^ (inputs[285]));
    assign layer0_outputs[1157] = ~(inputs[216]);
    assign layer0_outputs[1158] = ~((inputs[275]) ^ (inputs[45]));
    assign layer0_outputs[1159] = (inputs[244]) & ~(inputs[137]);
    assign layer0_outputs[1160] = inputs[369];
    assign layer0_outputs[1161] = ~((inputs[181]) | (inputs[278]));
    assign layer0_outputs[1162] = inputs[197];
    assign layer0_outputs[1163] = ~((inputs[320]) | (inputs[15]));
    assign layer0_outputs[1164] = inputs[92];
    assign layer0_outputs[1165] = (inputs[289]) & ~(inputs[298]);
    assign layer0_outputs[1166] = ~(inputs[10]);
    assign layer0_outputs[1167] = (inputs[79]) & ~(inputs[105]);
    assign layer0_outputs[1168] = (inputs[178]) ^ (inputs[121]);
    assign layer0_outputs[1169] = ~(inputs[340]);
    assign layer0_outputs[1170] = (inputs[346]) & ~(inputs[118]);
    assign layer0_outputs[1171] = ~(inputs[92]) | (inputs[123]);
    assign layer0_outputs[1172] = inputs[267];
    assign layer0_outputs[1173] = (inputs[326]) & ~(inputs[178]);
    assign layer0_outputs[1174] = ~(inputs[29]);
    assign layer0_outputs[1175] = (inputs[190]) | (inputs[130]);
    assign layer0_outputs[1176] = 1'b0;
    assign layer0_outputs[1177] = ~(inputs[88]) | (inputs[234]);
    assign layer0_outputs[1178] = (inputs[262]) | (inputs[280]);
    assign layer0_outputs[1179] = ~(inputs[94]);
    assign layer0_outputs[1180] = (inputs[214]) | (inputs[101]);
    assign layer0_outputs[1181] = inputs[42];
    assign layer0_outputs[1182] = (inputs[188]) ^ (inputs[195]);
    assign layer0_outputs[1183] = inputs[89];
    assign layer0_outputs[1184] = inputs[211];
    assign layer0_outputs[1185] = ~(inputs[364]) | (inputs[283]);
    assign layer0_outputs[1186] = ~((inputs[40]) ^ (inputs[68]));
    assign layer0_outputs[1187] = ~((inputs[258]) | (inputs[329]));
    assign layer0_outputs[1188] = ~(inputs[73]);
    assign layer0_outputs[1189] = inputs[134];
    assign layer0_outputs[1190] = ~(inputs[268]);
    assign layer0_outputs[1191] = (inputs[26]) & ~(inputs[127]);
    assign layer0_outputs[1192] = (inputs[150]) | (inputs[59]);
    assign layer0_outputs[1193] = inputs[153];
    assign layer0_outputs[1194] = ~(inputs[355]);
    assign layer0_outputs[1195] = (inputs[249]) & ~(inputs[202]);
    assign layer0_outputs[1196] = ~((inputs[222]) ^ (inputs[246]));
    assign layer0_outputs[1197] = inputs[242];
    assign layer0_outputs[1198] = (inputs[102]) ^ (inputs[297]);
    assign layer0_outputs[1199] = ~(inputs[73]);
    assign layer0_outputs[1200] = ~(inputs[114]);
    assign layer0_outputs[1201] = ~(inputs[178]);
    assign layer0_outputs[1202] = ~((inputs[179]) | (inputs[135]));
    assign layer0_outputs[1203] = inputs[275];
    assign layer0_outputs[1204] = (inputs[213]) & ~(inputs[11]);
    assign layer0_outputs[1205] = ~(inputs[217]);
    assign layer0_outputs[1206] = (inputs[390]) & ~(inputs[200]);
    assign layer0_outputs[1207] = (inputs[91]) ^ (inputs[66]);
    assign layer0_outputs[1208] = ~((inputs[292]) | (inputs[7]));
    assign layer0_outputs[1209] = ~((inputs[307]) | (inputs[396]));
    assign layer0_outputs[1210] = (inputs[272]) & ~(inputs[145]);
    assign layer0_outputs[1211] = ~(inputs[327]) | (inputs[153]);
    assign layer0_outputs[1212] = (inputs[396]) ^ (inputs[111]);
    assign layer0_outputs[1213] = (inputs[226]) ^ (inputs[325]);
    assign layer0_outputs[1214] = (inputs[310]) & ~(inputs[216]);
    assign layer0_outputs[1215] = ~(inputs[152]);
    assign layer0_outputs[1216] = (inputs[252]) & ~(inputs[123]);
    assign layer0_outputs[1217] = ~((inputs[60]) | (inputs[217]));
    assign layer0_outputs[1218] = ~(inputs[117]);
    assign layer0_outputs[1219] = ~((inputs[178]) | (inputs[136]));
    assign layer0_outputs[1220] = (inputs[194]) ^ (inputs[275]);
    assign layer0_outputs[1221] = ~(inputs[303]);
    assign layer0_outputs[1222] = inputs[285];
    assign layer0_outputs[1223] = ~(inputs[90]);
    assign layer0_outputs[1224] = inputs[51];
    assign layer0_outputs[1225] = (inputs[30]) & ~(inputs[220]);
    assign layer0_outputs[1226] = 1'b0;
    assign layer0_outputs[1227] = ~((inputs[97]) | (inputs[285]));
    assign layer0_outputs[1228] = ~(inputs[90]) | (inputs[62]);
    assign layer0_outputs[1229] = (inputs[64]) ^ (inputs[14]);
    assign layer0_outputs[1230] = inputs[90];
    assign layer0_outputs[1231] = inputs[347];
    assign layer0_outputs[1232] = (inputs[323]) & ~(inputs[162]);
    assign layer0_outputs[1233] = ~(inputs[130]);
    assign layer0_outputs[1234] = ~((inputs[24]) | (inputs[293]));
    assign layer0_outputs[1235] = (inputs[309]) & ~(inputs[182]);
    assign layer0_outputs[1236] = (inputs[187]) & ~(inputs[365]);
    assign layer0_outputs[1237] = inputs[305];
    assign layer0_outputs[1238] = ~(inputs[29]);
    assign layer0_outputs[1239] = inputs[119];
    assign layer0_outputs[1240] = ~(inputs[353]);
    assign layer0_outputs[1241] = (inputs[122]) | (inputs[396]);
    assign layer0_outputs[1242] = ~(inputs[223]) | (inputs[140]);
    assign layer0_outputs[1243] = (inputs[333]) & ~(inputs[217]);
    assign layer0_outputs[1244] = ~(inputs[47]);
    assign layer0_outputs[1245] = ~((inputs[45]) | (inputs[35]));
    assign layer0_outputs[1246] = ~((inputs[145]) & (inputs[374]));
    assign layer0_outputs[1247] = inputs[264];
    assign layer0_outputs[1248] = ~(inputs[36]) | (inputs[365]);
    assign layer0_outputs[1249] = inputs[4];
    assign layer0_outputs[1250] = inputs[94];
    assign layer0_outputs[1251] = ~(inputs[40]) | (inputs[180]);
    assign layer0_outputs[1252] = ~(inputs[285]);
    assign layer0_outputs[1253] = inputs[109];
    assign layer0_outputs[1254] = ~(inputs[237]);
    assign layer0_outputs[1255] = (inputs[218]) | (inputs[314]);
    assign layer0_outputs[1256] = (inputs[270]) | (inputs[17]);
    assign layer0_outputs[1257] = (inputs[369]) | (inputs[218]);
    assign layer0_outputs[1258] = ~((inputs[340]) | (inputs[255]));
    assign layer0_outputs[1259] = ~(inputs[169]) | (inputs[257]);
    assign layer0_outputs[1260] = ~((inputs[339]) | (inputs[209]));
    assign layer0_outputs[1261] = inputs[226];
    assign layer0_outputs[1262] = (inputs[281]) ^ (inputs[196]);
    assign layer0_outputs[1263] = (inputs[163]) | (inputs[376]);
    assign layer0_outputs[1264] = (inputs[390]) | (inputs[160]);
    assign layer0_outputs[1265] = ~(inputs[317]);
    assign layer0_outputs[1266] = ~(inputs[200]) | (inputs[331]);
    assign layer0_outputs[1267] = (inputs[104]) | (inputs[259]);
    assign layer0_outputs[1268] = inputs[225];
    assign layer0_outputs[1269] = (inputs[254]) & ~(inputs[8]);
    assign layer0_outputs[1270] = (inputs[61]) ^ (inputs[392]);
    assign layer0_outputs[1271] = 1'b1;
    assign layer0_outputs[1272] = (inputs[192]) & ~(inputs[314]);
    assign layer0_outputs[1273] = ~(inputs[304]);
    assign layer0_outputs[1274] = (inputs[243]) ^ (inputs[348]);
    assign layer0_outputs[1275] = ~(inputs[73]) | (inputs[160]);
    assign layer0_outputs[1276] = ~(inputs[12]) | (inputs[357]);
    assign layer0_outputs[1277] = inputs[30];
    assign layer0_outputs[1278] = ~(inputs[265]);
    assign layer0_outputs[1279] = inputs[34];
    assign layer0_outputs[1280] = ~((inputs[167]) ^ (inputs[227]));
    assign layer0_outputs[1281] = inputs[65];
    assign layer0_outputs[1282] = (inputs[266]) & (inputs[266]);
    assign layer0_outputs[1283] = ~((inputs[213]) | (inputs[59]));
    assign layer0_outputs[1284] = ~((inputs[176]) | (inputs[261]));
    assign layer0_outputs[1285] = ~((inputs[215]) ^ (inputs[177]));
    assign layer0_outputs[1286] = ~(inputs[189]);
    assign layer0_outputs[1287] = ~(inputs[224]);
    assign layer0_outputs[1288] = (inputs[175]) | (inputs[25]);
    assign layer0_outputs[1289] = ~((inputs[69]) & (inputs[47]));
    assign layer0_outputs[1290] = (inputs[297]) ^ (inputs[323]);
    assign layer0_outputs[1291] = (inputs[179]) ^ (inputs[355]);
    assign layer0_outputs[1292] = ~(inputs[92]) | (inputs[280]);
    assign layer0_outputs[1293] = inputs[368];
    assign layer0_outputs[1294] = (inputs[341]) | (inputs[140]);
    assign layer0_outputs[1295] = ~(inputs[93]) | (inputs[298]);
    assign layer0_outputs[1296] = ~(inputs[265]) | (inputs[102]);
    assign layer0_outputs[1297] = ~(inputs[246]);
    assign layer0_outputs[1298] = ~(inputs[269]);
    assign layer0_outputs[1299] = ~((inputs[173]) | (inputs[156]));
    assign layer0_outputs[1300] = ~(inputs[56]);
    assign layer0_outputs[1301] = ~(inputs[193]);
    assign layer0_outputs[1302] = (inputs[206]) & (inputs[98]);
    assign layer0_outputs[1303] = inputs[226];
    assign layer0_outputs[1304] = ~((inputs[183]) | (inputs[244]));
    assign layer0_outputs[1305] = ~((inputs[206]) | (inputs[115]));
    assign layer0_outputs[1306] = ~(inputs[125]);
    assign layer0_outputs[1307] = inputs[251];
    assign layer0_outputs[1308] = ~((inputs[329]) | (inputs[324]));
    assign layer0_outputs[1309] = ~(inputs[156]);
    assign layer0_outputs[1310] = (inputs[121]) | (inputs[184]);
    assign layer0_outputs[1311] = ~(inputs[48]);
    assign layer0_outputs[1312] = ~(inputs[315]);
    assign layer0_outputs[1313] = ~(inputs[98]);
    assign layer0_outputs[1314] = ~(inputs[26]);
    assign layer0_outputs[1315] = (inputs[154]) ^ (inputs[74]);
    assign layer0_outputs[1316] = inputs[71];
    assign layer0_outputs[1317] = ~(inputs[32]) | (inputs[152]);
    assign layer0_outputs[1318] = inputs[240];
    assign layer0_outputs[1319] = ~((inputs[308]) | (inputs[328]));
    assign layer0_outputs[1320] = inputs[69];
    assign layer0_outputs[1321] = ~(inputs[34]) | (inputs[259]);
    assign layer0_outputs[1322] = inputs[366];
    assign layer0_outputs[1323] = ~(inputs[272]) | (inputs[389]);
    assign layer0_outputs[1324] = ~((inputs[360]) | (inputs[352]));
    assign layer0_outputs[1325] = ~(inputs[51]);
    assign layer0_outputs[1326] = (inputs[175]) | (inputs[367]);
    assign layer0_outputs[1327] = inputs[386];
    assign layer0_outputs[1328] = ~(inputs[224]);
    assign layer0_outputs[1329] = (inputs[149]) & ~(inputs[224]);
    assign layer0_outputs[1330] = (inputs[9]) & ~(inputs[39]);
    assign layer0_outputs[1331] = (inputs[154]) | (inputs[18]);
    assign layer0_outputs[1332] = ~((inputs[305]) & (inputs[268]));
    assign layer0_outputs[1333] = ~(inputs[205]);
    assign layer0_outputs[1334] = inputs[356];
    assign layer0_outputs[1335] = ~((inputs[332]) & (inputs[265]));
    assign layer0_outputs[1336] = ~((inputs[318]) | (inputs[28]));
    assign layer0_outputs[1337] = ~((inputs[30]) | (inputs[253]));
    assign layer0_outputs[1338] = ~(inputs[284]);
    assign layer0_outputs[1339] = (inputs[387]) & ~(inputs[77]);
    assign layer0_outputs[1340] = inputs[149];
    assign layer0_outputs[1341] = (inputs[345]) & ~(inputs[61]);
    assign layer0_outputs[1342] = ~(inputs[124]) | (inputs[338]);
    assign layer0_outputs[1343] = inputs[142];
    assign layer0_outputs[1344] = ~((inputs[259]) ^ (inputs[155]));
    assign layer0_outputs[1345] = (inputs[257]) | (inputs[278]);
    assign layer0_outputs[1346] = inputs[315];
    assign layer0_outputs[1347] = ~((inputs[299]) | (inputs[150]));
    assign layer0_outputs[1348] = ~((inputs[352]) ^ (inputs[381]));
    assign layer0_outputs[1349] = ~(inputs[322]);
    assign layer0_outputs[1350] = (inputs[93]) | (inputs[320]);
    assign layer0_outputs[1351] = inputs[323];
    assign layer0_outputs[1352] = ~((inputs[100]) ^ (inputs[138]));
    assign layer0_outputs[1353] = (inputs[336]) ^ (inputs[395]);
    assign layer0_outputs[1354] = ~(inputs[188]);
    assign layer0_outputs[1355] = ~((inputs[65]) | (inputs[136]));
    assign layer0_outputs[1356] = (inputs[118]) | (inputs[228]);
    assign layer0_outputs[1357] = inputs[205];
    assign layer0_outputs[1358] = inputs[239];
    assign layer0_outputs[1359] = ~(inputs[346]);
    assign layer0_outputs[1360] = (inputs[107]) | (inputs[125]);
    assign layer0_outputs[1361] = ~(inputs[177]);
    assign layer0_outputs[1362] = ~((inputs[337]) ^ (inputs[349]));
    assign layer0_outputs[1363] = (inputs[394]) & ~(inputs[242]);
    assign layer0_outputs[1364] = ~(inputs[281]);
    assign layer0_outputs[1365] = (inputs[277]) ^ (inputs[315]);
    assign layer0_outputs[1366] = ~(inputs[56]) | (inputs[399]);
    assign layer0_outputs[1367] = ~((inputs[240]) | (inputs[219]));
    assign layer0_outputs[1368] = inputs[8];
    assign layer0_outputs[1369] = inputs[146];
    assign layer0_outputs[1370] = ~((inputs[221]) | (inputs[398]));
    assign layer0_outputs[1371] = ~(inputs[266]) | (inputs[94]);
    assign layer0_outputs[1372] = ~(inputs[59]);
    assign layer0_outputs[1373] = ~(inputs[50]);
    assign layer0_outputs[1374] = ~(inputs[201]) | (inputs[176]);
    assign layer0_outputs[1375] = inputs[202];
    assign layer0_outputs[1376] = ~((inputs[297]) | (inputs[221]));
    assign layer0_outputs[1377] = ~((inputs[257]) & (inputs[109]));
    assign layer0_outputs[1378] = inputs[114];
    assign layer0_outputs[1379] = (inputs[87]) & (inputs[146]);
    assign layer0_outputs[1380] = (inputs[183]) | (inputs[185]);
    assign layer0_outputs[1381] = inputs[163];
    assign layer0_outputs[1382] = ~(inputs[228]);
    assign layer0_outputs[1383] = (inputs[98]) & ~(inputs[374]);
    assign layer0_outputs[1384] = (inputs[345]) & ~(inputs[63]);
    assign layer0_outputs[1385] = inputs[9];
    assign layer0_outputs[1386] = ~(inputs[163]);
    assign layer0_outputs[1387] = (inputs[63]) | (inputs[37]);
    assign layer0_outputs[1388] = (inputs[203]) & ~(inputs[61]);
    assign layer0_outputs[1389] = (inputs[167]) & ~(inputs[286]);
    assign layer0_outputs[1390] = (inputs[105]) ^ (inputs[100]);
    assign layer0_outputs[1391] = ~(inputs[133]);
    assign layer0_outputs[1392] = ~(inputs[115]) | (inputs[187]);
    assign layer0_outputs[1393] = ~((inputs[59]) | (inputs[192]));
    assign layer0_outputs[1394] = ~((inputs[38]) | (inputs[17]));
    assign layer0_outputs[1395] = (inputs[173]) & ~(inputs[20]);
    assign layer0_outputs[1396] = ~(inputs[161]);
    assign layer0_outputs[1397] = ~((inputs[112]) & (inputs[292]));
    assign layer0_outputs[1398] = (inputs[36]) & ~(inputs[379]);
    assign layer0_outputs[1399] = ~(inputs[238]);
    assign layer0_outputs[1400] = ~(inputs[190]);
    assign layer0_outputs[1401] = inputs[196];
    assign layer0_outputs[1402] = (inputs[359]) | (inputs[338]);
    assign layer0_outputs[1403] = ~(inputs[192]) | (inputs[390]);
    assign layer0_outputs[1404] = ~(inputs[267]);
    assign layer0_outputs[1405] = (inputs[253]) | (inputs[17]);
    assign layer0_outputs[1406] = (inputs[122]) ^ (inputs[323]);
    assign layer0_outputs[1407] = inputs[158];
    assign layer0_outputs[1408] = ~(inputs[395]) | (inputs[44]);
    assign layer0_outputs[1409] = (inputs[316]) & ~(inputs[272]);
    assign layer0_outputs[1410] = ~(inputs[77]);
    assign layer0_outputs[1411] = (inputs[185]) ^ (inputs[160]);
    assign layer0_outputs[1412] = (inputs[146]) ^ (inputs[82]);
    assign layer0_outputs[1413] = ~(inputs[126]);
    assign layer0_outputs[1414] = ~((inputs[152]) | (inputs[101]));
    assign layer0_outputs[1415] = ~((inputs[295]) ^ (inputs[136]));
    assign layer0_outputs[1416] = ~(inputs[32]);
    assign layer0_outputs[1417] = ~((inputs[46]) ^ (inputs[60]));
    assign layer0_outputs[1418] = ~((inputs[220]) | (inputs[267]));
    assign layer0_outputs[1419] = (inputs[207]) ^ (inputs[331]);
    assign layer0_outputs[1420] = ~((inputs[309]) | (inputs[265]));
    assign layer0_outputs[1421] = ~(inputs[195]);
    assign layer0_outputs[1422] = ~(inputs[205]) | (inputs[110]);
    assign layer0_outputs[1423] = (inputs[180]) ^ (inputs[295]);
    assign layer0_outputs[1424] = inputs[227];
    assign layer0_outputs[1425] = (inputs[62]) | (inputs[286]);
    assign layer0_outputs[1426] = ~(inputs[96]) | (inputs[208]);
    assign layer0_outputs[1427] = (inputs[37]) & ~(inputs[265]);
    assign layer0_outputs[1428] = ~(inputs[347]);
    assign layer0_outputs[1429] = ~(inputs[290]) | (inputs[346]);
    assign layer0_outputs[1430] = inputs[334];
    assign layer0_outputs[1431] = (inputs[14]) | (inputs[302]);
    assign layer0_outputs[1432] = 1'b1;
    assign layer0_outputs[1433] = inputs[189];
    assign layer0_outputs[1434] = ~(inputs[137]);
    assign layer0_outputs[1435] = ~(inputs[33]);
    assign layer0_outputs[1436] = ~(inputs[131]);
    assign layer0_outputs[1437] = (inputs[399]) | (inputs[231]);
    assign layer0_outputs[1438] = ~(inputs[319]);
    assign layer0_outputs[1439] = ~((inputs[191]) ^ (inputs[313]));
    assign layer0_outputs[1440] = ~(inputs[265]);
    assign layer0_outputs[1441] = inputs[46];
    assign layer0_outputs[1442] = (inputs[310]) ^ (inputs[241]);
    assign layer0_outputs[1443] = (inputs[308]) & (inputs[291]);
    assign layer0_outputs[1444] = inputs[369];
    assign layer0_outputs[1445] = (inputs[209]) & ~(inputs[166]);
    assign layer0_outputs[1446] = ~(inputs[254]);
    assign layer0_outputs[1447] = (inputs[284]) ^ (inputs[91]);
    assign layer0_outputs[1448] = ~(inputs[382]) | (inputs[66]);
    assign layer0_outputs[1449] = ~((inputs[299]) ^ (inputs[198]));
    assign layer0_outputs[1450] = ~(inputs[163]);
    assign layer0_outputs[1451] = ~(inputs[387]);
    assign layer0_outputs[1452] = ~(inputs[190]) | (inputs[120]);
    assign layer0_outputs[1453] = inputs[60];
    assign layer0_outputs[1454] = (inputs[273]) ^ (inputs[350]);
    assign layer0_outputs[1455] = inputs[133];
    assign layer0_outputs[1456] = (inputs[158]) | (inputs[24]);
    assign layer0_outputs[1457] = (inputs[228]) | (inputs[22]);
    assign layer0_outputs[1458] = inputs[39];
    assign layer0_outputs[1459] = inputs[142];
    assign layer0_outputs[1460] = ~(inputs[231]) | (inputs[151]);
    assign layer0_outputs[1461] = ~((inputs[321]) ^ (inputs[123]));
    assign layer0_outputs[1462] = (inputs[372]) | (inputs[386]);
    assign layer0_outputs[1463] = ~((inputs[6]) ^ (inputs[336]));
    assign layer0_outputs[1464] = inputs[261];
    assign layer0_outputs[1465] = ~((inputs[225]) ^ (inputs[65]));
    assign layer0_outputs[1466] = ~((inputs[212]) | (inputs[155]));
    assign layer0_outputs[1467] = ~((inputs[209]) ^ (inputs[207]));
    assign layer0_outputs[1468] = (inputs[194]) & ~(inputs[19]);
    assign layer0_outputs[1469] = ~((inputs[94]) & (inputs[167]));
    assign layer0_outputs[1470] = inputs[31];
    assign layer0_outputs[1471] = 1'b1;
    assign layer0_outputs[1472] = ~((inputs[131]) | (inputs[92]));
    assign layer0_outputs[1473] = inputs[134];
    assign layer0_outputs[1474] = ~((inputs[265]) | (inputs[374]));
    assign layer0_outputs[1475] = ~(inputs[147]) | (inputs[38]);
    assign layer0_outputs[1476] = ~((inputs[322]) | (inputs[227]));
    assign layer0_outputs[1477] = ~((inputs[110]) | (inputs[259]));
    assign layer0_outputs[1478] = (inputs[260]) ^ (inputs[300]);
    assign layer0_outputs[1479] = ~(inputs[354]);
    assign layer0_outputs[1480] = ~(inputs[144]);
    assign layer0_outputs[1481] = (inputs[141]) | (inputs[103]);
    assign layer0_outputs[1482] = (inputs[106]) & ~(inputs[91]);
    assign layer0_outputs[1483] = ~(inputs[218]);
    assign layer0_outputs[1484] = ~((inputs[189]) | (inputs[383]));
    assign layer0_outputs[1485] = inputs[230];
    assign layer0_outputs[1486] = inputs[204];
    assign layer0_outputs[1487] = inputs[375];
    assign layer0_outputs[1488] = (inputs[165]) & ~(inputs[178]);
    assign layer0_outputs[1489] = ~(inputs[256]);
    assign layer0_outputs[1490] = (inputs[296]) ^ (inputs[50]);
    assign layer0_outputs[1491] = (inputs[46]) & ~(inputs[184]);
    assign layer0_outputs[1492] = ~((inputs[132]) | (inputs[224]));
    assign layer0_outputs[1493] = ~(inputs[276]);
    assign layer0_outputs[1494] = ~(inputs[317]) | (inputs[220]);
    assign layer0_outputs[1495] = (inputs[231]) & ~(inputs[287]);
    assign layer0_outputs[1496] = (inputs[341]) | (inputs[41]);
    assign layer0_outputs[1497] = ~((inputs[232]) ^ (inputs[210]));
    assign layer0_outputs[1498] = ~(inputs[148]) | (inputs[2]);
    assign layer0_outputs[1499] = ~((inputs[269]) & (inputs[171]));
    assign layer0_outputs[1500] = (inputs[64]) & ~(inputs[342]);
    assign layer0_outputs[1501] = (inputs[124]) | (inputs[180]);
    assign layer0_outputs[1502] = (inputs[229]) ^ (inputs[251]);
    assign layer0_outputs[1503] = ~(inputs[6]);
    assign layer0_outputs[1504] = inputs[83];
    assign layer0_outputs[1505] = ~((inputs[303]) | (inputs[325]));
    assign layer0_outputs[1506] = (inputs[324]) | (inputs[282]);
    assign layer0_outputs[1507] = (inputs[7]) | (inputs[189]);
    assign layer0_outputs[1508] = (inputs[360]) & (inputs[93]);
    assign layer0_outputs[1509] = inputs[227];
    assign layer0_outputs[1510] = (inputs[67]) | (inputs[57]);
    assign layer0_outputs[1511] = ~(inputs[298]);
    assign layer0_outputs[1512] = ~((inputs[305]) | (inputs[305]));
    assign layer0_outputs[1513] = ~((inputs[38]) & (inputs[365]));
    assign layer0_outputs[1514] = (inputs[277]) & ~(inputs[119]);
    assign layer0_outputs[1515] = ~(inputs[94]) | (inputs[376]);
    assign layer0_outputs[1516] = ~(inputs[129]);
    assign layer0_outputs[1517] = ~(inputs[166]);
    assign layer0_outputs[1518] = ~(inputs[280]);
    assign layer0_outputs[1519] = ~(inputs[29]) | (inputs[198]);
    assign layer0_outputs[1520] = (inputs[70]) | (inputs[388]);
    assign layer0_outputs[1521] = ~(inputs[33]);
    assign layer0_outputs[1522] = ~(inputs[226]) | (inputs[398]);
    assign layer0_outputs[1523] = ~(inputs[298]) | (inputs[137]);
    assign layer0_outputs[1524] = inputs[329];
    assign layer0_outputs[1525] = ~(inputs[367]);
    assign layer0_outputs[1526] = inputs[58];
    assign layer0_outputs[1527] = ~(inputs[388]) | (inputs[270]);
    assign layer0_outputs[1528] = (inputs[367]) & ~(inputs[160]);
    assign layer0_outputs[1529] = ~(inputs[173]);
    assign layer0_outputs[1530] = (inputs[179]) | (inputs[127]);
    assign layer0_outputs[1531] = ~(inputs[74]);
    assign layer0_outputs[1532] = ~((inputs[116]) & (inputs[355]));
    assign layer0_outputs[1533] = ~(inputs[118]);
    assign layer0_outputs[1534] = (inputs[32]) & ~(inputs[321]);
    assign layer0_outputs[1535] = ~((inputs[165]) ^ (inputs[95]));
    assign layer0_outputs[1536] = inputs[233];
    assign layer0_outputs[1537] = inputs[249];
    assign layer0_outputs[1538] = inputs[2];
    assign layer0_outputs[1539] = 1'b1;
    assign layer0_outputs[1540] = ~((inputs[80]) | (inputs[49]));
    assign layer0_outputs[1541] = inputs[344];
    assign layer0_outputs[1542] = ~((inputs[356]) ^ (inputs[306]));
    assign layer0_outputs[1543] = (inputs[7]) & ~(inputs[25]);
    assign layer0_outputs[1544] = ~(inputs[306]);
    assign layer0_outputs[1545] = (inputs[229]) & ~(inputs[4]);
    assign layer0_outputs[1546] = ~((inputs[281]) ^ (inputs[254]));
    assign layer0_outputs[1547] = 1'b0;
    assign layer0_outputs[1548] = (inputs[148]) & ~(inputs[258]);
    assign layer0_outputs[1549] = 1'b0;
    assign layer0_outputs[1550] = (inputs[181]) & (inputs[238]);
    assign layer0_outputs[1551] = ~(inputs[95]);
    assign layer0_outputs[1552] = ~((inputs[113]) ^ (inputs[97]));
    assign layer0_outputs[1553] = (inputs[43]) & (inputs[26]);
    assign layer0_outputs[1554] = 1'b1;
    assign layer0_outputs[1555] = ~(inputs[267]);
    assign layer0_outputs[1556] = ~(inputs[388]) | (inputs[380]);
    assign layer0_outputs[1557] = inputs[378];
    assign layer0_outputs[1558] = inputs[143];
    assign layer0_outputs[1559] = ~((inputs[213]) | (inputs[241]));
    assign layer0_outputs[1560] = (inputs[122]) & ~(inputs[369]);
    assign layer0_outputs[1561] = ~(inputs[233]);
    assign layer0_outputs[1562] = (inputs[135]) & ~(inputs[220]);
    assign layer0_outputs[1563] = (inputs[96]) & ~(inputs[202]);
    assign layer0_outputs[1564] = ~(inputs[347]);
    assign layer0_outputs[1565] = (inputs[6]) | (inputs[254]);
    assign layer0_outputs[1566] = ~(inputs[200]);
    assign layer0_outputs[1567] = ~((inputs[192]) | (inputs[105]));
    assign layer0_outputs[1568] = inputs[183];
    assign layer0_outputs[1569] = ~(inputs[245]) | (inputs[329]);
    assign layer0_outputs[1570] = inputs[46];
    assign layer0_outputs[1571] = (inputs[21]) | (inputs[173]);
    assign layer0_outputs[1572] = (inputs[208]) | (inputs[162]);
    assign layer0_outputs[1573] = ~(inputs[371]);
    assign layer0_outputs[1574] = (inputs[239]) | (inputs[386]);
    assign layer0_outputs[1575] = (inputs[262]) | (inputs[185]);
    assign layer0_outputs[1576] = ~(inputs[225]);
    assign layer0_outputs[1577] = (inputs[258]) | (inputs[363]);
    assign layer0_outputs[1578] = inputs[93];
    assign layer0_outputs[1579] = ~((inputs[348]) & (inputs[147]));
    assign layer0_outputs[1580] = ~(inputs[153]);
    assign layer0_outputs[1581] = (inputs[205]) | (inputs[78]);
    assign layer0_outputs[1582] = inputs[189];
    assign layer0_outputs[1583] = (inputs[77]) & (inputs[110]);
    assign layer0_outputs[1584] = (inputs[288]) & ~(inputs[116]);
    assign layer0_outputs[1585] = 1'b1;
    assign layer0_outputs[1586] = (inputs[394]) | (inputs[381]);
    assign layer0_outputs[1587] = ~(inputs[156]);
    assign layer0_outputs[1588] = (inputs[256]) | (inputs[379]);
    assign layer0_outputs[1589] = ~((inputs[116]) | (inputs[179]));
    assign layer0_outputs[1590] = ~((inputs[178]) | (inputs[213]));
    assign layer0_outputs[1591] = ~((inputs[214]) | (inputs[184]));
    assign layer0_outputs[1592] = (inputs[367]) & ~(inputs[135]);
    assign layer0_outputs[1593] = ~(inputs[11]) | (inputs[276]);
    assign layer0_outputs[1594] = (inputs[203]) | (inputs[166]);
    assign layer0_outputs[1595] = (inputs[263]) & ~(inputs[160]);
    assign layer0_outputs[1596] = inputs[138];
    assign layer0_outputs[1597] = ~((inputs[393]) ^ (inputs[294]));
    assign layer0_outputs[1598] = ~((inputs[8]) ^ (inputs[283]));
    assign layer0_outputs[1599] = inputs[69];
    assign layer0_outputs[1600] = (inputs[309]) | (inputs[227]);
    assign layer0_outputs[1601] = ~((inputs[75]) | (inputs[59]));
    assign layer0_outputs[1602] = (inputs[291]) ^ (inputs[228]);
    assign layer0_outputs[1603] = ~((inputs[392]) & (inputs[330]));
    assign layer0_outputs[1604] = (inputs[391]) ^ (inputs[56]);
    assign layer0_outputs[1605] = ~((inputs[181]) | (inputs[91]));
    assign layer0_outputs[1606] = ~(inputs[313]);
    assign layer0_outputs[1607] = inputs[37];
    assign layer0_outputs[1608] = (inputs[154]) | (inputs[242]);
    assign layer0_outputs[1609] = ~((inputs[52]) & (inputs[150]));
    assign layer0_outputs[1610] = (inputs[368]) | (inputs[52]);
    assign layer0_outputs[1611] = ~(inputs[222]);
    assign layer0_outputs[1612] = (inputs[41]) ^ (inputs[22]);
    assign layer0_outputs[1613] = (inputs[375]) | (inputs[343]);
    assign layer0_outputs[1614] = ~((inputs[367]) ^ (inputs[49]));
    assign layer0_outputs[1615] = ~(inputs[228]);
    assign layer0_outputs[1616] = inputs[269];
    assign layer0_outputs[1617] = inputs[194];
    assign layer0_outputs[1618] = (inputs[204]) & ~(inputs[342]);
    assign layer0_outputs[1619] = inputs[286];
    assign layer0_outputs[1620] = ~((inputs[362]) ^ (inputs[309]));
    assign layer0_outputs[1621] = ~((inputs[53]) | (inputs[292]));
    assign layer0_outputs[1622] = ~(inputs[346]);
    assign layer0_outputs[1623] = 1'b0;
    assign layer0_outputs[1624] = (inputs[87]) & ~(inputs[243]);
    assign layer0_outputs[1625] = (inputs[321]) | (inputs[188]);
    assign layer0_outputs[1626] = inputs[229];
    assign layer0_outputs[1627] = (inputs[113]) ^ (inputs[52]);
    assign layer0_outputs[1628] = (inputs[242]) ^ (inputs[210]);
    assign layer0_outputs[1629] = (inputs[213]) & (inputs[369]);
    assign layer0_outputs[1630] = ~(inputs[364]);
    assign layer0_outputs[1631] = inputs[230];
    assign layer0_outputs[1632] = ~(inputs[171]);
    assign layer0_outputs[1633] = (inputs[94]) ^ (inputs[150]);
    assign layer0_outputs[1634] = inputs[230];
    assign layer0_outputs[1635] = ~(inputs[211]);
    assign layer0_outputs[1636] = ~((inputs[338]) | (inputs[137]));
    assign layer0_outputs[1637] = inputs[251];
    assign layer0_outputs[1638] = ~(inputs[353]) | (inputs[191]);
    assign layer0_outputs[1639] = inputs[217];
    assign layer0_outputs[1640] = ~((inputs[210]) & (inputs[308]));
    assign layer0_outputs[1641] = inputs[163];
    assign layer0_outputs[1642] = ~((inputs[32]) | (inputs[76]));
    assign layer0_outputs[1643] = inputs[228];
    assign layer0_outputs[1644] = (inputs[97]) | (inputs[3]);
    assign layer0_outputs[1645] = ~((inputs[191]) ^ (inputs[235]));
    assign layer0_outputs[1646] = (inputs[33]) | (inputs[120]);
    assign layer0_outputs[1647] = inputs[29];
    assign layer0_outputs[1648] = ~((inputs[353]) | (inputs[343]));
    assign layer0_outputs[1649] = ~((inputs[345]) | (inputs[288]));
    assign layer0_outputs[1650] = ~((inputs[264]) ^ (inputs[128]));
    assign layer0_outputs[1651] = (inputs[65]) & ~(inputs[139]);
    assign layer0_outputs[1652] = ~((inputs[221]) & (inputs[372]));
    assign layer0_outputs[1653] = ~((inputs[219]) | (inputs[270]));
    assign layer0_outputs[1654] = ~(inputs[308]) | (inputs[54]);
    assign layer0_outputs[1655] = inputs[322];
    assign layer0_outputs[1656] = ~((inputs[167]) | (inputs[237]));
    assign layer0_outputs[1657] = ~(inputs[311]);
    assign layer0_outputs[1658] = ~(inputs[107]) | (inputs[62]);
    assign layer0_outputs[1659] = (inputs[183]) | (inputs[278]);
    assign layer0_outputs[1660] = inputs[164];
    assign layer0_outputs[1661] = inputs[89];
    assign layer0_outputs[1662] = ~((inputs[154]) ^ (inputs[166]));
    assign layer0_outputs[1663] = (inputs[214]) & ~(inputs[45]);
    assign layer0_outputs[1664] = inputs[375];
    assign layer0_outputs[1665] = ~((inputs[124]) | (inputs[139]));
    assign layer0_outputs[1666] = inputs[148];
    assign layer0_outputs[1667] = ~(inputs[75]) | (inputs[29]);
    assign layer0_outputs[1668] = ~(inputs[387]);
    assign layer0_outputs[1669] = (inputs[390]) & ~(inputs[16]);
    assign layer0_outputs[1670] = (inputs[119]) | (inputs[237]);
    assign layer0_outputs[1671] = (inputs[148]) & ~(inputs[120]);
    assign layer0_outputs[1672] = inputs[163];
    assign layer0_outputs[1673] = (inputs[253]) & ~(inputs[86]);
    assign layer0_outputs[1674] = (inputs[16]) ^ (inputs[48]);
    assign layer0_outputs[1675] = ~(inputs[168]);
    assign layer0_outputs[1676] = ~(inputs[65]);
    assign layer0_outputs[1677] = ~((inputs[385]) | (inputs[391]));
    assign layer0_outputs[1678] = ~((inputs[387]) ^ (inputs[200]));
    assign layer0_outputs[1679] = ~((inputs[318]) | (inputs[85]));
    assign layer0_outputs[1680] = ~(inputs[66]);
    assign layer0_outputs[1681] = ~((inputs[187]) & (inputs[185]));
    assign layer0_outputs[1682] = (inputs[28]) | (inputs[339]);
    assign layer0_outputs[1683] = (inputs[381]) | (inputs[351]);
    assign layer0_outputs[1684] = (inputs[309]) ^ (inputs[302]);
    assign layer0_outputs[1685] = ~(inputs[249]) | (inputs[146]);
    assign layer0_outputs[1686] = ~((inputs[273]) | (inputs[281]));
    assign layer0_outputs[1687] = ~(inputs[223]) | (inputs[120]);
    assign layer0_outputs[1688] = inputs[331];
    assign layer0_outputs[1689] = ~((inputs[266]) | (inputs[229]));
    assign layer0_outputs[1690] = ~(inputs[31]);
    assign layer0_outputs[1691] = ~((inputs[306]) | (inputs[198]));
    assign layer0_outputs[1692] = ~((inputs[293]) ^ (inputs[392]));
    assign layer0_outputs[1693] = inputs[89];
    assign layer0_outputs[1694] = 1'b0;
    assign layer0_outputs[1695] = (inputs[106]) | (inputs[146]);
    assign layer0_outputs[1696] = inputs[255];
    assign layer0_outputs[1697] = ~((inputs[322]) & (inputs[128]));
    assign layer0_outputs[1698] = ~(inputs[121]);
    assign layer0_outputs[1699] = ~(inputs[104]);
    assign layer0_outputs[1700] = ~(inputs[96]) | (inputs[370]);
    assign layer0_outputs[1701] = inputs[20];
    assign layer0_outputs[1702] = inputs[166];
    assign layer0_outputs[1703] = (inputs[115]) ^ (inputs[78]);
    assign layer0_outputs[1704] = (inputs[172]) & ~(inputs[82]);
    assign layer0_outputs[1705] = (inputs[258]) | (inputs[282]);
    assign layer0_outputs[1706] = inputs[351];
    assign layer0_outputs[1707] = ~(inputs[188]) | (inputs[200]);
    assign layer0_outputs[1708] = ~(inputs[224]) | (inputs[80]);
    assign layer0_outputs[1709] = (inputs[24]) ^ (inputs[363]);
    assign layer0_outputs[1710] = ~(inputs[349]) | (inputs[79]);
    assign layer0_outputs[1711] = ~((inputs[141]) ^ (inputs[388]));
    assign layer0_outputs[1712] = ~(inputs[161]);
    assign layer0_outputs[1713] = ~((inputs[248]) & (inputs[278]));
    assign layer0_outputs[1714] = ~(inputs[213]) | (inputs[84]);
    assign layer0_outputs[1715] = ~((inputs[259]) ^ (inputs[5]));
    assign layer0_outputs[1716] = (inputs[396]) | (inputs[106]);
    assign layer0_outputs[1717] = ~((inputs[194]) | (inputs[242]));
    assign layer0_outputs[1718] = (inputs[241]) ^ (inputs[68]);
    assign layer0_outputs[1719] = ~(inputs[253]) | (inputs[348]);
    assign layer0_outputs[1720] = ~(inputs[222]) | (inputs[20]);
    assign layer0_outputs[1721] = ~(inputs[61]);
    assign layer0_outputs[1722] = ~(inputs[95]);
    assign layer0_outputs[1723] = (inputs[215]) ^ (inputs[162]);
    assign layer0_outputs[1724] = (inputs[226]) ^ (inputs[254]);
    assign layer0_outputs[1725] = (inputs[221]) | (inputs[379]);
    assign layer0_outputs[1726] = ~((inputs[175]) ^ (inputs[138]));
    assign layer0_outputs[1727] = (inputs[318]) ^ (inputs[214]);
    assign layer0_outputs[1728] = ~((inputs[185]) ^ (inputs[222]));
    assign layer0_outputs[1729] = ~(inputs[207]) | (inputs[297]);
    assign layer0_outputs[1730] = ~(inputs[355]) | (inputs[161]);
    assign layer0_outputs[1731] = inputs[327];
    assign layer0_outputs[1732] = ~(inputs[260]) | (inputs[372]);
    assign layer0_outputs[1733] = ~((inputs[194]) | (inputs[161]));
    assign layer0_outputs[1734] = inputs[88];
    assign layer0_outputs[1735] = inputs[43];
    assign layer0_outputs[1736] = (inputs[130]) | (inputs[303]);
    assign layer0_outputs[1737] = ~((inputs[117]) | (inputs[370]));
    assign layer0_outputs[1738] = (inputs[10]) & ~(inputs[18]);
    assign layer0_outputs[1739] = (inputs[145]) & ~(inputs[237]);
    assign layer0_outputs[1740] = (inputs[203]) & ~(inputs[233]);
    assign layer0_outputs[1741] = ~(inputs[236]);
    assign layer0_outputs[1742] = ~((inputs[143]) | (inputs[170]));
    assign layer0_outputs[1743] = (inputs[124]) | (inputs[341]);
    assign layer0_outputs[1744] = (inputs[379]) | (inputs[172]);
    assign layer0_outputs[1745] = ~(inputs[244]);
    assign layer0_outputs[1746] = (inputs[123]) ^ (inputs[88]);
    assign layer0_outputs[1747] = ~(inputs[388]) | (inputs[288]);
    assign layer0_outputs[1748] = inputs[301];
    assign layer0_outputs[1749] = inputs[291];
    assign layer0_outputs[1750] = inputs[182];
    assign layer0_outputs[1751] = ~((inputs[81]) | (inputs[272]));
    assign layer0_outputs[1752] = ~((inputs[226]) | (inputs[369]));
    assign layer0_outputs[1753] = (inputs[205]) | (inputs[246]);
    assign layer0_outputs[1754] = (inputs[119]) | (inputs[103]);
    assign layer0_outputs[1755] = inputs[90];
    assign layer0_outputs[1756] = (inputs[317]) | (inputs[335]);
    assign layer0_outputs[1757] = ~(inputs[47]);
    assign layer0_outputs[1758] = (inputs[197]) & ~(inputs[80]);
    assign layer0_outputs[1759] = ~((inputs[212]) | (inputs[270]));
    assign layer0_outputs[1760] = (inputs[188]) | (inputs[379]);
    assign layer0_outputs[1761] = ~((inputs[3]) | (inputs[386]));
    assign layer0_outputs[1762] = inputs[258];
    assign layer0_outputs[1763] = (inputs[124]) & ~(inputs[341]);
    assign layer0_outputs[1764] = inputs[185];
    assign layer0_outputs[1765] = ~(inputs[75]);
    assign layer0_outputs[1766] = inputs[122];
    assign layer0_outputs[1767] = (inputs[7]) | (inputs[235]);
    assign layer0_outputs[1768] = ~(inputs[176]) | (inputs[362]);
    assign layer0_outputs[1769] = ~(inputs[302]);
    assign layer0_outputs[1770] = ~(inputs[268]);
    assign layer0_outputs[1771] = ~(inputs[96]);
    assign layer0_outputs[1772] = inputs[144];
    assign layer0_outputs[1773] = ~(inputs[9]) | (inputs[246]);
    assign layer0_outputs[1774] = ~((inputs[344]) & (inputs[260]));
    assign layer0_outputs[1775] = inputs[48];
    assign layer0_outputs[1776] = inputs[13];
    assign layer0_outputs[1777] = ~((inputs[118]) | (inputs[266]));
    assign layer0_outputs[1778] = (inputs[153]) & ~(inputs[98]);
    assign layer0_outputs[1779] = (inputs[366]) & ~(inputs[134]);
    assign layer0_outputs[1780] = ~((inputs[202]) | (inputs[368]));
    assign layer0_outputs[1781] = (inputs[366]) | (inputs[275]);
    assign layer0_outputs[1782] = inputs[89];
    assign layer0_outputs[1783] = ~(inputs[57]) | (inputs[396]);
    assign layer0_outputs[1784] = (inputs[151]) & ~(inputs[164]);
    assign layer0_outputs[1785] = inputs[351];
    assign layer0_outputs[1786] = ~((inputs[328]) | (inputs[260]));
    assign layer0_outputs[1787] = ~(inputs[262]);
    assign layer0_outputs[1788] = ~(inputs[212]) | (inputs[359]);
    assign layer0_outputs[1789] = (inputs[97]) & ~(inputs[4]);
    assign layer0_outputs[1790] = (inputs[390]) & ~(inputs[137]);
    assign layer0_outputs[1791] = ~((inputs[120]) | (inputs[321]));
    assign layer0_outputs[1792] = inputs[370];
    assign layer0_outputs[1793] = inputs[46];
    assign layer0_outputs[1794] = ~(inputs[13]) | (inputs[162]);
    assign layer0_outputs[1795] = (inputs[293]) & ~(inputs[177]);
    assign layer0_outputs[1796] = (inputs[282]) ^ (inputs[395]);
    assign layer0_outputs[1797] = ~(inputs[313]) | (inputs[352]);
    assign layer0_outputs[1798] = (inputs[32]) & ~(inputs[350]);
    assign layer0_outputs[1799] = ~((inputs[381]) | (inputs[181]));
    assign layer0_outputs[1800] = (inputs[323]) ^ (inputs[55]);
    assign layer0_outputs[1801] = (inputs[113]) | (inputs[23]);
    assign layer0_outputs[1802] = (inputs[153]) & ~(inputs[398]);
    assign layer0_outputs[1803] = ~((inputs[88]) ^ (inputs[24]));
    assign layer0_outputs[1804] = (inputs[276]) & ~(inputs[82]);
    assign layer0_outputs[1805] = ~(inputs[191]) | (inputs[222]);
    assign layer0_outputs[1806] = (inputs[233]) | (inputs[18]);
    assign layer0_outputs[1807] = ~(inputs[127]) | (inputs[214]);
    assign layer0_outputs[1808] = ~(inputs[60]);
    assign layer0_outputs[1809] = (inputs[113]) & ~(inputs[42]);
    assign layer0_outputs[1810] = (inputs[235]) & ~(inputs[0]);
    assign layer0_outputs[1811] = ~(inputs[159]);
    assign layer0_outputs[1812] = (inputs[329]) & ~(inputs[78]);
    assign layer0_outputs[1813] = ~((inputs[140]) ^ (inputs[286]));
    assign layer0_outputs[1814] = (inputs[104]) | (inputs[271]);
    assign layer0_outputs[1815] = (inputs[358]) | (inputs[211]);
    assign layer0_outputs[1816] = inputs[136];
    assign layer0_outputs[1817] = ~((inputs[251]) ^ (inputs[232]));
    assign layer0_outputs[1818] = ~(inputs[247]);
    assign layer0_outputs[1819] = ~((inputs[140]) ^ (inputs[187]));
    assign layer0_outputs[1820] = inputs[218];
    assign layer0_outputs[1821] = ~((inputs[214]) ^ (inputs[178]));
    assign layer0_outputs[1822] = inputs[335];
    assign layer0_outputs[1823] = ~(inputs[203]) | (inputs[62]);
    assign layer0_outputs[1824] = ~(inputs[184]);
    assign layer0_outputs[1825] = inputs[252];
    assign layer0_outputs[1826] = (inputs[243]) & ~(inputs[397]);
    assign layer0_outputs[1827] = ~(inputs[382]);
    assign layer0_outputs[1828] = ~((inputs[272]) ^ (inputs[262]));
    assign layer0_outputs[1829] = ~((inputs[39]) | (inputs[22]));
    assign layer0_outputs[1830] = ~(inputs[317]);
    assign layer0_outputs[1831] = (inputs[207]) ^ (inputs[247]);
    assign layer0_outputs[1832] = inputs[193];
    assign layer0_outputs[1833] = inputs[105];
    assign layer0_outputs[1834] = (inputs[168]) ^ (inputs[108]);
    assign layer0_outputs[1835] = ~(inputs[14]);
    assign layer0_outputs[1836] = ~((inputs[66]) ^ (inputs[68]));
    assign layer0_outputs[1837] = ~((inputs[377]) | (inputs[195]));
    assign layer0_outputs[1838] = (inputs[303]) | (inputs[286]);
    assign layer0_outputs[1839] = (inputs[352]) & ~(inputs[66]);
    assign layer0_outputs[1840] = ~((inputs[204]) | (inputs[233]));
    assign layer0_outputs[1841] = ~((inputs[366]) ^ (inputs[260]));
    assign layer0_outputs[1842] = ~((inputs[21]) | (inputs[36]));
    assign layer0_outputs[1843] = (inputs[24]) & ~(inputs[242]);
    assign layer0_outputs[1844] = ~(inputs[125]) | (inputs[361]);
    assign layer0_outputs[1845] = ~(inputs[66]) | (inputs[370]);
    assign layer0_outputs[1846] = ~((inputs[48]) | (inputs[204]));
    assign layer0_outputs[1847] = ~((inputs[175]) ^ (inputs[279]));
    assign layer0_outputs[1848] = (inputs[240]) ^ (inputs[206]);
    assign layer0_outputs[1849] = ~((inputs[165]) ^ (inputs[129]));
    assign layer0_outputs[1850] = ~((inputs[332]) | (inputs[123]));
    assign layer0_outputs[1851] = (inputs[20]) | (inputs[113]);
    assign layer0_outputs[1852] = 1'b1;
    assign layer0_outputs[1853] = ~(inputs[94]);
    assign layer0_outputs[1854] = ~(inputs[157]);
    assign layer0_outputs[1855] = ~(inputs[41]) | (inputs[326]);
    assign layer0_outputs[1856] = inputs[172];
    assign layer0_outputs[1857] = (inputs[48]) ^ (inputs[120]);
    assign layer0_outputs[1858] = (inputs[303]) & ~(inputs[36]);
    assign layer0_outputs[1859] = ~(inputs[343]);
    assign layer0_outputs[1860] = ~((inputs[300]) | (inputs[0]));
    assign layer0_outputs[1861] = inputs[19];
    assign layer0_outputs[1862] = ~((inputs[359]) | (inputs[83]));
    assign layer0_outputs[1863] = (inputs[73]) | (inputs[3]);
    assign layer0_outputs[1864] = inputs[9];
    assign layer0_outputs[1865] = ~(inputs[369]);
    assign layer0_outputs[1866] = ~((inputs[31]) | (inputs[305]));
    assign layer0_outputs[1867] = inputs[13];
    assign layer0_outputs[1868] = ~(inputs[45]);
    assign layer0_outputs[1869] = inputs[148];
    assign layer0_outputs[1870] = inputs[152];
    assign layer0_outputs[1871] = ~(inputs[257]) | (inputs[188]);
    assign layer0_outputs[1872] = ~(inputs[370]) | (inputs[15]);
    assign layer0_outputs[1873] = ~(inputs[77]);
    assign layer0_outputs[1874] = ~((inputs[246]) | (inputs[341]));
    assign layer0_outputs[1875] = (inputs[86]) ^ (inputs[28]);
    assign layer0_outputs[1876] = inputs[310];
    assign layer0_outputs[1877] = ~((inputs[88]) ^ (inputs[83]));
    assign layer0_outputs[1878] = inputs[86];
    assign layer0_outputs[1879] = (inputs[388]) & ~(inputs[0]);
    assign layer0_outputs[1880] = inputs[344];
    assign layer0_outputs[1881] = ~((inputs[399]) | (inputs[202]));
    assign layer0_outputs[1882] = ~(inputs[116]);
    assign layer0_outputs[1883] = inputs[239];
    assign layer0_outputs[1884] = ~(inputs[188]) | (inputs[60]);
    assign layer0_outputs[1885] = ~(inputs[109]);
    assign layer0_outputs[1886] = ~(inputs[368]) | (inputs[136]);
    assign layer0_outputs[1887] = (inputs[97]) | (inputs[320]);
    assign layer0_outputs[1888] = ~(inputs[278]) | (inputs[178]);
    assign layer0_outputs[1889] = inputs[335];
    assign layer0_outputs[1890] = ~(inputs[320]);
    assign layer0_outputs[1891] = (inputs[251]) | (inputs[212]);
    assign layer0_outputs[1892] = ~(inputs[270]);
    assign layer0_outputs[1893] = inputs[96];
    assign layer0_outputs[1894] = ~((inputs[291]) | (inputs[379]));
    assign layer0_outputs[1895] = ~(inputs[186]) | (inputs[262]);
    assign layer0_outputs[1896] = (inputs[370]) & ~(inputs[40]);
    assign layer0_outputs[1897] = ~(inputs[184]) | (inputs[136]);
    assign layer0_outputs[1898] = (inputs[59]) | (inputs[261]);
    assign layer0_outputs[1899] = inputs[319];
    assign layer0_outputs[1900] = (inputs[16]) ^ (inputs[227]);
    assign layer0_outputs[1901] = inputs[123];
    assign layer0_outputs[1902] = (inputs[279]) & ~(inputs[325]);
    assign layer0_outputs[1903] = inputs[23];
    assign layer0_outputs[1904] = ~((inputs[195]) | (inputs[39]));
    assign layer0_outputs[1905] = ~((inputs[357]) | (inputs[126]));
    assign layer0_outputs[1906] = ~(inputs[74]);
    assign layer0_outputs[1907] = ~((inputs[240]) | (inputs[232]));
    assign layer0_outputs[1908] = ~(inputs[120]);
    assign layer0_outputs[1909] = (inputs[272]) & ~(inputs[69]);
    assign layer0_outputs[1910] = (inputs[121]) | (inputs[367]);
    assign layer0_outputs[1911] = ~(inputs[76]);
    assign layer0_outputs[1912] = inputs[52];
    assign layer0_outputs[1913] = ~((inputs[205]) | (inputs[376]));
    assign layer0_outputs[1914] = ~(inputs[386]) | (inputs[124]);
    assign layer0_outputs[1915] = ~(inputs[329]);
    assign layer0_outputs[1916] = ~((inputs[316]) | (inputs[3]));
    assign layer0_outputs[1917] = ~(inputs[102]);
    assign layer0_outputs[1918] = ~(inputs[29]);
    assign layer0_outputs[1919] = ~(inputs[125]) | (inputs[40]);
    assign layer0_outputs[1920] = ~((inputs[78]) | (inputs[237]));
    assign layer0_outputs[1921] = ~((inputs[353]) | (inputs[340]));
    assign layer0_outputs[1922] = ~((inputs[45]) | (inputs[98]));
    assign layer0_outputs[1923] = inputs[301];
    assign layer0_outputs[1924] = ~((inputs[231]) | (inputs[215]));
    assign layer0_outputs[1925] = (inputs[64]) | (inputs[41]);
    assign layer0_outputs[1926] = 1'b0;
    assign layer0_outputs[1927] = inputs[351];
    assign layer0_outputs[1928] = ~(inputs[348]) | (inputs[2]);
    assign layer0_outputs[1929] = ~(inputs[45]);
    assign layer0_outputs[1930] = ~((inputs[14]) ^ (inputs[243]));
    assign layer0_outputs[1931] = (inputs[3]) | (inputs[79]);
    assign layer0_outputs[1932] = (inputs[69]) | (inputs[390]);
    assign layer0_outputs[1933] = (inputs[196]) | (inputs[159]);
    assign layer0_outputs[1934] = ~(inputs[48]) | (inputs[162]);
    assign layer0_outputs[1935] = inputs[320];
    assign layer0_outputs[1936] = ~((inputs[343]) ^ (inputs[351]));
    assign layer0_outputs[1937] = (inputs[179]) | (inputs[294]);
    assign layer0_outputs[1938] = (inputs[383]) & (inputs[299]);
    assign layer0_outputs[1939] = ~(inputs[268]);
    assign layer0_outputs[1940] = (inputs[43]) & ~(inputs[275]);
    assign layer0_outputs[1941] = inputs[24];
    assign layer0_outputs[1942] = ~((inputs[397]) ^ (inputs[287]));
    assign layer0_outputs[1943] = ~((inputs[393]) ^ (inputs[341]));
    assign layer0_outputs[1944] = (inputs[253]) ^ (inputs[131]);
    assign layer0_outputs[1945] = ~(inputs[332]);
    assign layer0_outputs[1946] = ~(inputs[290]);
    assign layer0_outputs[1947] = inputs[71];
    assign layer0_outputs[1948] = ~(inputs[368]);
    assign layer0_outputs[1949] = ~((inputs[399]) | (inputs[329]));
    assign layer0_outputs[1950] = (inputs[248]) | (inputs[339]);
    assign layer0_outputs[1951] = (inputs[264]) | (inputs[181]);
    assign layer0_outputs[1952] = inputs[125];
    assign layer0_outputs[1953] = ~(inputs[130]) | (inputs[159]);
    assign layer0_outputs[1954] = ~(inputs[261]);
    assign layer0_outputs[1955] = ~(inputs[294]) | (inputs[101]);
    assign layer0_outputs[1956] = ~(inputs[84]);
    assign layer0_outputs[1957] = inputs[285];
    assign layer0_outputs[1958] = 1'b0;
    assign layer0_outputs[1959] = 1'b1;
    assign layer0_outputs[1960] = ~(inputs[104]) | (inputs[69]);
    assign layer0_outputs[1961] = (inputs[293]) & ~(inputs[126]);
    assign layer0_outputs[1962] = ~(inputs[163]);
    assign layer0_outputs[1963] = ~((inputs[187]) | (inputs[372]));
    assign layer0_outputs[1964] = (inputs[361]) | (inputs[98]);
    assign layer0_outputs[1965] = ~((inputs[331]) | (inputs[18]));
    assign layer0_outputs[1966] = (inputs[169]) ^ (inputs[103]);
    assign layer0_outputs[1967] = ~(inputs[114]) | (inputs[199]);
    assign layer0_outputs[1968] = inputs[246];
    assign layer0_outputs[1969] = ~((inputs[117]) | (inputs[384]));
    assign layer0_outputs[1970] = 1'b0;
    assign layer0_outputs[1971] = ~((inputs[150]) ^ (inputs[216]));
    assign layer0_outputs[1972] = ~((inputs[273]) | (inputs[33]));
    assign layer0_outputs[1973] = ~((inputs[45]) ^ (inputs[274]));
    assign layer0_outputs[1974] = ~((inputs[263]) ^ (inputs[184]));
    assign layer0_outputs[1975] = ~(inputs[225]) | (inputs[37]);
    assign layer0_outputs[1976] = ~(inputs[234]) | (inputs[12]);
    assign layer0_outputs[1977] = (inputs[344]) & ~(inputs[31]);
    assign layer0_outputs[1978] = ~(inputs[190]) | (inputs[277]);
    assign layer0_outputs[1979] = 1'b1;
    assign layer0_outputs[1980] = ~(inputs[263]);
    assign layer0_outputs[1981] = (inputs[187]) & ~(inputs[145]);
    assign layer0_outputs[1982] = inputs[346];
    assign layer0_outputs[1983] = ~((inputs[372]) & (inputs[372]));
    assign layer0_outputs[1984] = ~(inputs[133]);
    assign layer0_outputs[1985] = (inputs[384]) | (inputs[102]);
    assign layer0_outputs[1986] = inputs[9];
    assign layer0_outputs[1987] = (inputs[112]) & ~(inputs[313]);
    assign layer0_outputs[1988] = ~((inputs[319]) ^ (inputs[44]));
    assign layer0_outputs[1989] = inputs[162];
    assign layer0_outputs[1990] = ~(inputs[168]);
    assign layer0_outputs[1991] = 1'b1;
    assign layer0_outputs[1992] = inputs[208];
    assign layer0_outputs[1993] = (inputs[105]) & ~(inputs[175]);
    assign layer0_outputs[1994] = 1'b0;
    assign layer0_outputs[1995] = ~(inputs[80]) | (inputs[161]);
    assign layer0_outputs[1996] = ~((inputs[334]) | (inputs[393]));
    assign layer0_outputs[1997] = ~((inputs[262]) | (inputs[387]));
    assign layer0_outputs[1998] = ~(inputs[160]) | (inputs[289]);
    assign layer0_outputs[1999] = inputs[286];
    assign layer0_outputs[2000] = ~(inputs[45]);
    assign layer0_outputs[2001] = (inputs[33]) ^ (inputs[258]);
    assign layer0_outputs[2002] = ~(inputs[392]);
    assign layer0_outputs[2003] = ~((inputs[372]) | (inputs[342]));
    assign layer0_outputs[2004] = (inputs[2]) | (inputs[121]);
    assign layer0_outputs[2005] = ~(inputs[48]) | (inputs[200]);
    assign layer0_outputs[2006] = ~(inputs[147]);
    assign layer0_outputs[2007] = (inputs[168]) | (inputs[228]);
    assign layer0_outputs[2008] = (inputs[1]) | (inputs[23]);
    assign layer0_outputs[2009] = ~(inputs[347]);
    assign layer0_outputs[2010] = (inputs[29]) & ~(inputs[145]);
    assign layer0_outputs[2011] = (inputs[148]) ^ (inputs[129]);
    assign layer0_outputs[2012] = ~((inputs[324]) | (inputs[304]));
    assign layer0_outputs[2013] = (inputs[143]) | (inputs[396]);
    assign layer0_outputs[2014] = inputs[348];
    assign layer0_outputs[2015] = ~(inputs[120]);
    assign layer0_outputs[2016] = ~(inputs[49]);
    assign layer0_outputs[2017] = ~(inputs[43]);
    assign layer0_outputs[2018] = ~(inputs[170]);
    assign layer0_outputs[2019] = inputs[282];
    assign layer0_outputs[2020] = ~(inputs[199]);
    assign layer0_outputs[2021] = (inputs[13]) ^ (inputs[9]);
    assign layer0_outputs[2022] = ~((inputs[90]) & (inputs[342]));
    assign layer0_outputs[2023] = inputs[316];
    assign layer0_outputs[2024] = (inputs[172]) & ~(inputs[8]);
    assign layer0_outputs[2025] = (inputs[325]) & ~(inputs[378]);
    assign layer0_outputs[2026] = ~(inputs[89]);
    assign layer0_outputs[2027] = inputs[234];
    assign layer0_outputs[2028] = inputs[127];
    assign layer0_outputs[2029] = (inputs[330]) & ~(inputs[247]);
    assign layer0_outputs[2030] = ~(inputs[166]);
    assign layer0_outputs[2031] = ~(inputs[128]) | (inputs[43]);
    assign layer0_outputs[2032] = ~((inputs[201]) ^ (inputs[204]));
    assign layer0_outputs[2033] = ~((inputs[309]) ^ (inputs[382]));
    assign layer0_outputs[2034] = inputs[5];
    assign layer0_outputs[2035] = (inputs[63]) | (inputs[90]);
    assign layer0_outputs[2036] = ~((inputs[108]) | (inputs[159]));
    assign layer0_outputs[2037] = ~(inputs[4]) | (inputs[271]);
    assign layer0_outputs[2038] = ~(inputs[302]);
    assign layer0_outputs[2039] = ~((inputs[236]) | (inputs[200]));
    assign layer0_outputs[2040] = ~((inputs[171]) | (inputs[232]));
    assign layer0_outputs[2041] = inputs[170];
    assign layer0_outputs[2042] = ~(inputs[6]) | (inputs[296]);
    assign layer0_outputs[2043] = ~(inputs[335]) | (inputs[177]);
    assign layer0_outputs[2044] = (inputs[296]) | (inputs[333]);
    assign layer0_outputs[2045] = inputs[326];
    assign layer0_outputs[2046] = (inputs[275]) & ~(inputs[105]);
    assign layer0_outputs[2047] = (inputs[220]) ^ (inputs[7]);
    assign layer0_outputs[2048] = (inputs[369]) & ~(inputs[379]);
    assign layer0_outputs[2049] = (inputs[263]) | (inputs[386]);
    assign layer0_outputs[2050] = ~(inputs[118]) | (inputs[393]);
    assign layer0_outputs[2051] = inputs[92];
    assign layer0_outputs[2052] = (inputs[153]) | (inputs[111]);
    assign layer0_outputs[2053] = 1'b0;
    assign layer0_outputs[2054] = ~(inputs[227]) | (inputs[8]);
    assign layer0_outputs[2055] = (inputs[333]) & ~(inputs[56]);
    assign layer0_outputs[2056] = ~(inputs[288]) | (inputs[38]);
    assign layer0_outputs[2057] = inputs[223];
    assign layer0_outputs[2058] = ~((inputs[71]) | (inputs[23]));
    assign layer0_outputs[2059] = ~((inputs[63]) ^ (inputs[28]));
    assign layer0_outputs[2060] = ~((inputs[155]) | (inputs[143]));
    assign layer0_outputs[2061] = inputs[307];
    assign layer0_outputs[2062] = 1'b0;
    assign layer0_outputs[2063] = (inputs[219]) & ~(inputs[98]);
    assign layer0_outputs[2064] = inputs[27];
    assign layer0_outputs[2065] = (inputs[81]) | (inputs[116]);
    assign layer0_outputs[2066] = inputs[190];
    assign layer0_outputs[2067] = (inputs[371]) & ~(inputs[382]);
    assign layer0_outputs[2068] = (inputs[171]) & ~(inputs[87]);
    assign layer0_outputs[2069] = inputs[269];
    assign layer0_outputs[2070] = (inputs[64]) ^ (inputs[362]);
    assign layer0_outputs[2071] = ~(inputs[203]) | (inputs[34]);
    assign layer0_outputs[2072] = ~(inputs[27]);
    assign layer0_outputs[2073] = inputs[25];
    assign layer0_outputs[2074] = inputs[112];
    assign layer0_outputs[2075] = inputs[364];
    assign layer0_outputs[2076] = inputs[280];
    assign layer0_outputs[2077] = ~((inputs[220]) | (inputs[252]));
    assign layer0_outputs[2078] = ~((inputs[346]) ^ (inputs[103]));
    assign layer0_outputs[2079] = ~(inputs[87]) | (inputs[382]);
    assign layer0_outputs[2080] = (inputs[125]) | (inputs[168]);
    assign layer0_outputs[2081] = (inputs[114]) | (inputs[42]);
    assign layer0_outputs[2082] = inputs[269];
    assign layer0_outputs[2083] = inputs[125];
    assign layer0_outputs[2084] = ~((inputs[166]) | (inputs[391]));
    assign layer0_outputs[2085] = (inputs[325]) & ~(inputs[75]);
    assign layer0_outputs[2086] = ~(inputs[163]);
    assign layer0_outputs[2087] = (inputs[79]) ^ (inputs[82]);
    assign layer0_outputs[2088] = ~(inputs[21]);
    assign layer0_outputs[2089] = ~((inputs[160]) ^ (inputs[108]));
    assign layer0_outputs[2090] = (inputs[385]) ^ (inputs[310]);
    assign layer0_outputs[2091] = ~(inputs[391]) | (inputs[319]);
    assign layer0_outputs[2092] = ~(inputs[34]);
    assign layer0_outputs[2093] = inputs[56];
    assign layer0_outputs[2094] = (inputs[238]) | (inputs[274]);
    assign layer0_outputs[2095] = ~(inputs[166]);
    assign layer0_outputs[2096] = ~((inputs[203]) & (inputs[223]));
    assign layer0_outputs[2097] = inputs[154];
    assign layer0_outputs[2098] = (inputs[100]) & ~(inputs[141]);
    assign layer0_outputs[2099] = (inputs[392]) ^ (inputs[99]);
    assign layer0_outputs[2100] = (inputs[317]) & ~(inputs[121]);
    assign layer0_outputs[2101] = ~((inputs[303]) ^ (inputs[48]));
    assign layer0_outputs[2102] = ~(inputs[273]);
    assign layer0_outputs[2103] = (inputs[273]) & ~(inputs[358]);
    assign layer0_outputs[2104] = inputs[111];
    assign layer0_outputs[2105] = inputs[229];
    assign layer0_outputs[2106] = ~(inputs[101]);
    assign layer0_outputs[2107] = ~((inputs[245]) ^ (inputs[241]));
    assign layer0_outputs[2108] = ~((inputs[205]) ^ (inputs[102]));
    assign layer0_outputs[2109] = inputs[36];
    assign layer0_outputs[2110] = inputs[182];
    assign layer0_outputs[2111] = inputs[133];
    assign layer0_outputs[2112] = (inputs[368]) & ~(inputs[177]);
    assign layer0_outputs[2113] = (inputs[248]) | (inputs[44]);
    assign layer0_outputs[2114] = ~((inputs[367]) ^ (inputs[216]));
    assign layer0_outputs[2115] = (inputs[375]) & ~(inputs[238]);
    assign layer0_outputs[2116] = (inputs[265]) ^ (inputs[304]);
    assign layer0_outputs[2117] = (inputs[261]) ^ (inputs[65]);
    assign layer0_outputs[2118] = ~(inputs[80]) | (inputs[1]);
    assign layer0_outputs[2119] = ~((inputs[51]) ^ (inputs[86]));
    assign layer0_outputs[2120] = ~(inputs[244]);
    assign layer0_outputs[2121] = ~((inputs[56]) | (inputs[290]));
    assign layer0_outputs[2122] = ~(inputs[393]) | (inputs[236]);
    assign layer0_outputs[2123] = ~(inputs[115]);
    assign layer0_outputs[2124] = (inputs[129]) | (inputs[286]);
    assign layer0_outputs[2125] = (inputs[198]) ^ (inputs[274]);
    assign layer0_outputs[2126] = ~(inputs[145]);
    assign layer0_outputs[2127] = (inputs[46]) & ~(inputs[241]);
    assign layer0_outputs[2128] = ~(inputs[191]);
    assign layer0_outputs[2129] = (inputs[66]) | (inputs[38]);
    assign layer0_outputs[2130] = inputs[196];
    assign layer0_outputs[2131] = (inputs[117]) | (inputs[372]);
    assign layer0_outputs[2132] = ~(inputs[191]) | (inputs[245]);
    assign layer0_outputs[2133] = (inputs[64]) | (inputs[76]);
    assign layer0_outputs[2134] = (inputs[298]) & ~(inputs[56]);
    assign layer0_outputs[2135] = 1'b0;
    assign layer0_outputs[2136] = (inputs[250]) ^ (inputs[385]);
    assign layer0_outputs[2137] = ~(inputs[274]);
    assign layer0_outputs[2138] = ~((inputs[26]) & (inputs[5]));
    assign layer0_outputs[2139] = ~(inputs[117]);
    assign layer0_outputs[2140] = (inputs[222]) ^ (inputs[5]);
    assign layer0_outputs[2141] = ~((inputs[12]) | (inputs[31]));
    assign layer0_outputs[2142] = ~(inputs[196]) | (inputs[189]);
    assign layer0_outputs[2143] = ~(inputs[387]) | (inputs[228]);
    assign layer0_outputs[2144] = ~((inputs[264]) | (inputs[110]));
    assign layer0_outputs[2145] = ~((inputs[25]) & (inputs[188]));
    assign layer0_outputs[2146] = ~((inputs[107]) | (inputs[165]));
    assign layer0_outputs[2147] = ~(inputs[396]) | (inputs[312]);
    assign layer0_outputs[2148] = inputs[362];
    assign layer0_outputs[2149] = ~((inputs[135]) | (inputs[115]));
    assign layer0_outputs[2150] = inputs[316];
    assign layer0_outputs[2151] = ~(inputs[245]);
    assign layer0_outputs[2152] = (inputs[46]) | (inputs[139]);
    assign layer0_outputs[2153] = ~(inputs[331]) | (inputs[381]);
    assign layer0_outputs[2154] = (inputs[331]) | (inputs[100]);
    assign layer0_outputs[2155] = (inputs[256]) & ~(inputs[270]);
    assign layer0_outputs[2156] = (inputs[129]) & ~(inputs[198]);
    assign layer0_outputs[2157] = ~(inputs[49]);
    assign layer0_outputs[2158] = ~(inputs[12]) | (inputs[235]);
    assign layer0_outputs[2159] = 1'b0;
    assign layer0_outputs[2160] = inputs[224];
    assign layer0_outputs[2161] = ~(inputs[70]) | (inputs[76]);
    assign layer0_outputs[2162] = (inputs[224]) ^ (inputs[282]);
    assign layer0_outputs[2163] = (inputs[90]) | (inputs[308]);
    assign layer0_outputs[2164] = ~(inputs[175]) | (inputs[239]);
    assign layer0_outputs[2165] = (inputs[327]) | (inputs[309]);
    assign layer0_outputs[2166] = ~(inputs[90]);
    assign layer0_outputs[2167] = ~(inputs[26]) | (inputs[379]);
    assign layer0_outputs[2168] = ~((inputs[30]) ^ (inputs[160]));
    assign layer0_outputs[2169] = ~((inputs[382]) ^ (inputs[189]));
    assign layer0_outputs[2170] = ~(inputs[371]);
    assign layer0_outputs[2171] = ~(inputs[339]);
    assign layer0_outputs[2172] = ~(inputs[335]);
    assign layer0_outputs[2173] = inputs[37];
    assign layer0_outputs[2174] = ~(inputs[98]) | (inputs[154]);
    assign layer0_outputs[2175] = ~((inputs[171]) ^ (inputs[169]));
    assign layer0_outputs[2176] = (inputs[242]) ^ (inputs[350]);
    assign layer0_outputs[2177] = ~((inputs[269]) | (inputs[376]));
    assign layer0_outputs[2178] = ~(inputs[30]) | (inputs[358]);
    assign layer0_outputs[2179] = (inputs[385]) | (inputs[203]);
    assign layer0_outputs[2180] = (inputs[334]) & ~(inputs[118]);
    assign layer0_outputs[2181] = ~((inputs[229]) ^ (inputs[261]));
    assign layer0_outputs[2182] = ~((inputs[349]) & (inputs[52]));
    assign layer0_outputs[2183] = inputs[60];
    assign layer0_outputs[2184] = ~((inputs[69]) | (inputs[26]));
    assign layer0_outputs[2185] = inputs[395];
    assign layer0_outputs[2186] = inputs[9];
    assign layer0_outputs[2187] = ~(inputs[169]);
    assign layer0_outputs[2188] = inputs[25];
    assign layer0_outputs[2189] = ~(inputs[53]);
    assign layer0_outputs[2190] = inputs[131];
    assign layer0_outputs[2191] = ~((inputs[59]) | (inputs[10]));
    assign layer0_outputs[2192] = (inputs[97]) & ~(inputs[289]);
    assign layer0_outputs[2193] = (inputs[348]) ^ (inputs[288]);
    assign layer0_outputs[2194] = ~((inputs[241]) ^ (inputs[107]));
    assign layer0_outputs[2195] = (inputs[271]) ^ (inputs[108]);
    assign layer0_outputs[2196] = (inputs[218]) & ~(inputs[247]);
    assign layer0_outputs[2197] = inputs[108];
    assign layer0_outputs[2198] = (inputs[371]) & ~(inputs[159]);
    assign layer0_outputs[2199] = (inputs[187]) | (inputs[151]);
    assign layer0_outputs[2200] = (inputs[105]) ^ (inputs[19]);
    assign layer0_outputs[2201] = inputs[67];
    assign layer0_outputs[2202] = (inputs[21]) | (inputs[7]);
    assign layer0_outputs[2203] = ~(inputs[244]);
    assign layer0_outputs[2204] = ~(inputs[282]) | (inputs[389]);
    assign layer0_outputs[2205] = (inputs[141]) & (inputs[340]);
    assign layer0_outputs[2206] = ~(inputs[168]);
    assign layer0_outputs[2207] = ~(inputs[275]);
    assign layer0_outputs[2208] = ~(inputs[186]);
    assign layer0_outputs[2209] = ~(inputs[171]) | (inputs[375]);
    assign layer0_outputs[2210] = ~(inputs[15]) | (inputs[393]);
    assign layer0_outputs[2211] = inputs[35];
    assign layer0_outputs[2212] = (inputs[48]) ^ (inputs[54]);
    assign layer0_outputs[2213] = inputs[7];
    assign layer0_outputs[2214] = inputs[8];
    assign layer0_outputs[2215] = inputs[126];
    assign layer0_outputs[2216] = ~(inputs[342]) | (inputs[263]);
    assign layer0_outputs[2217] = ~((inputs[268]) & (inputs[328]));
    assign layer0_outputs[2218] = ~((inputs[299]) | (inputs[297]));
    assign layer0_outputs[2219] = ~(inputs[310]);
    assign layer0_outputs[2220] = ~(inputs[322]);
    assign layer0_outputs[2221] = inputs[235];
    assign layer0_outputs[2222] = (inputs[125]) & ~(inputs[51]);
    assign layer0_outputs[2223] = ~((inputs[35]) ^ (inputs[261]));
    assign layer0_outputs[2224] = inputs[157];
    assign layer0_outputs[2225] = (inputs[281]) & ~(inputs[198]);
    assign layer0_outputs[2226] = ~(inputs[305]);
    assign layer0_outputs[2227] = ~((inputs[40]) ^ (inputs[134]));
    assign layer0_outputs[2228] = ~((inputs[162]) | (inputs[54]));
    assign layer0_outputs[2229] = ~((inputs[147]) | (inputs[298]));
    assign layer0_outputs[2230] = inputs[165];
    assign layer0_outputs[2231] = (inputs[171]) & ~(inputs[139]);
    assign layer0_outputs[2232] = inputs[350];
    assign layer0_outputs[2233] = inputs[363];
    assign layer0_outputs[2234] = inputs[49];
    assign layer0_outputs[2235] = ~((inputs[77]) ^ (inputs[135]));
    assign layer0_outputs[2236] = ~((inputs[55]) | (inputs[300]));
    assign layer0_outputs[2237] = inputs[31];
    assign layer0_outputs[2238] = ~((inputs[215]) | (inputs[393]));
    assign layer0_outputs[2239] = (inputs[25]) ^ (inputs[54]);
    assign layer0_outputs[2240] = ~((inputs[318]) | (inputs[10]));
    assign layer0_outputs[2241] = inputs[364];
    assign layer0_outputs[2242] = ~((inputs[73]) | (inputs[3]));
    assign layer0_outputs[2243] = inputs[211];
    assign layer0_outputs[2244] = ~((inputs[336]) | (inputs[341]));
    assign layer0_outputs[2245] = inputs[389];
    assign layer0_outputs[2246] = (inputs[59]) | (inputs[189]);
    assign layer0_outputs[2247] = 1'b0;
    assign layer0_outputs[2248] = ~((inputs[231]) | (inputs[21]));
    assign layer0_outputs[2249] = (inputs[5]) | (inputs[340]);
    assign layer0_outputs[2250] = (inputs[91]) & (inputs[172]);
    assign layer0_outputs[2251] = ~((inputs[333]) ^ (inputs[118]));
    assign layer0_outputs[2252] = (inputs[158]) & ~(inputs[74]);
    assign layer0_outputs[2253] = inputs[249];
    assign layer0_outputs[2254] = (inputs[282]) | (inputs[321]);
    assign layer0_outputs[2255] = (inputs[119]) ^ (inputs[259]);
    assign layer0_outputs[2256] = (inputs[21]) & ~(inputs[123]);
    assign layer0_outputs[2257] = (inputs[115]) & ~(inputs[302]);
    assign layer0_outputs[2258] = (inputs[13]) & ~(inputs[128]);
    assign layer0_outputs[2259] = (inputs[322]) | (inputs[70]);
    assign layer0_outputs[2260] = inputs[164];
    assign layer0_outputs[2261] = ~((inputs[327]) | (inputs[63]));
    assign layer0_outputs[2262] = inputs[357];
    assign layer0_outputs[2263] = ~((inputs[335]) | (inputs[179]));
    assign layer0_outputs[2264] = ~((inputs[164]) ^ (inputs[270]));
    assign layer0_outputs[2265] = inputs[265];
    assign layer0_outputs[2266] = ~((inputs[43]) ^ (inputs[355]));
    assign layer0_outputs[2267] = (inputs[144]) ^ (inputs[263]);
    assign layer0_outputs[2268] = inputs[155];
    assign layer0_outputs[2269] = (inputs[239]) | (inputs[183]);
    assign layer0_outputs[2270] = ~((inputs[242]) & (inputs[338]));
    assign layer0_outputs[2271] = ~((inputs[271]) | (inputs[236]));
    assign layer0_outputs[2272] = (inputs[252]) & ~(inputs[102]);
    assign layer0_outputs[2273] = inputs[288];
    assign layer0_outputs[2274] = ~((inputs[354]) | (inputs[232]));
    assign layer0_outputs[2275] = (inputs[194]) & ~(inputs[306]);
    assign layer0_outputs[2276] = ~(inputs[102]);
    assign layer0_outputs[2277] = ~(inputs[220]);
    assign layer0_outputs[2278] = ~(inputs[112]);
    assign layer0_outputs[2279] = ~(inputs[18]) | (inputs[225]);
    assign layer0_outputs[2280] = inputs[267];
    assign layer0_outputs[2281] = (inputs[147]) | (inputs[264]);
    assign layer0_outputs[2282] = (inputs[125]) | (inputs[53]);
    assign layer0_outputs[2283] = ~((inputs[311]) | (inputs[13]));
    assign layer0_outputs[2284] = ~(inputs[390]) | (inputs[268]);
    assign layer0_outputs[2285] = ~(inputs[270]);
    assign layer0_outputs[2286] = ~((inputs[146]) ^ (inputs[130]));
    assign layer0_outputs[2287] = inputs[267];
    assign layer0_outputs[2288] = ~((inputs[285]) | (inputs[280]));
    assign layer0_outputs[2289] = (inputs[364]) & (inputs[244]);
    assign layer0_outputs[2290] = (inputs[35]) ^ (inputs[311]);
    assign layer0_outputs[2291] = ~(inputs[333]);
    assign layer0_outputs[2292] = ~(inputs[75]);
    assign layer0_outputs[2293] = (inputs[368]) | (inputs[81]);
    assign layer0_outputs[2294] = ~((inputs[185]) | (inputs[182]));
    assign layer0_outputs[2295] = ~(inputs[156]);
    assign layer0_outputs[2296] = ~(inputs[343]);
    assign layer0_outputs[2297] = (inputs[263]) & ~(inputs[155]);
    assign layer0_outputs[2298] = inputs[39];
    assign layer0_outputs[2299] = ~(inputs[317]);
    assign layer0_outputs[2300] = ~(inputs[182]);
    assign layer0_outputs[2301] = (inputs[276]) ^ (inputs[214]);
    assign layer0_outputs[2302] = ~(inputs[29]) | (inputs[188]);
    assign layer0_outputs[2303] = ~(inputs[321]);
    assign layer0_outputs[2304] = inputs[271];
    assign layer0_outputs[2305] = ~(inputs[319]);
    assign layer0_outputs[2306] = ~((inputs[126]) ^ (inputs[47]));
    assign layer0_outputs[2307] = ~(inputs[167]);
    assign layer0_outputs[2308] = (inputs[245]) ^ (inputs[160]);
    assign layer0_outputs[2309] = (inputs[57]) & (inputs[173]);
    assign layer0_outputs[2310] = ~(inputs[186]) | (inputs[0]);
    assign layer0_outputs[2311] = ~(inputs[152]) | (inputs[187]);
    assign layer0_outputs[2312] = inputs[366];
    assign layer0_outputs[2313] = ~((inputs[4]) | (inputs[320]));
    assign layer0_outputs[2314] = ~(inputs[150]) | (inputs[360]);
    assign layer0_outputs[2315] = (inputs[65]) & ~(inputs[143]);
    assign layer0_outputs[2316] = inputs[359];
    assign layer0_outputs[2317] = ~((inputs[70]) ^ (inputs[330]));
    assign layer0_outputs[2318] = ~(inputs[243]);
    assign layer0_outputs[2319] = ~(inputs[368]);
    assign layer0_outputs[2320] = (inputs[111]) & ~(inputs[331]);
    assign layer0_outputs[2321] = (inputs[3]) & ~(inputs[374]);
    assign layer0_outputs[2322] = ~((inputs[255]) ^ (inputs[12]));
    assign layer0_outputs[2323] = ~((inputs[57]) | (inputs[189]));
    assign layer0_outputs[2324] = ~(inputs[142]);
    assign layer0_outputs[2325] = inputs[267];
    assign layer0_outputs[2326] = inputs[76];
    assign layer0_outputs[2327] = (inputs[394]) & ~(inputs[121]);
    assign layer0_outputs[2328] = (inputs[293]) & ~(inputs[211]);
    assign layer0_outputs[2329] = inputs[314];
    assign layer0_outputs[2330] = (inputs[82]) & ~(inputs[324]);
    assign layer0_outputs[2331] = (inputs[285]) & (inputs[233]);
    assign layer0_outputs[2332] = inputs[192];
    assign layer0_outputs[2333] = ~((inputs[115]) | (inputs[60]));
    assign layer0_outputs[2334] = (inputs[248]) & (inputs[247]);
    assign layer0_outputs[2335] = ~(inputs[98]);
    assign layer0_outputs[2336] = 1'b0;
    assign layer0_outputs[2337] = ~((inputs[10]) | (inputs[77]));
    assign layer0_outputs[2338] = ~(inputs[112]) | (inputs[149]);
    assign layer0_outputs[2339] = (inputs[273]) | (inputs[336]);
    assign layer0_outputs[2340] = inputs[102];
    assign layer0_outputs[2341] = (inputs[35]) ^ (inputs[77]);
    assign layer0_outputs[2342] = ~(inputs[282]);
    assign layer0_outputs[2343] = ~(inputs[311]) | (inputs[139]);
    assign layer0_outputs[2344] = ~(inputs[95]);
    assign layer0_outputs[2345] = ~(inputs[253]) | (inputs[18]);
    assign layer0_outputs[2346] = ~(inputs[55]) | (inputs[178]);
    assign layer0_outputs[2347] = (inputs[201]) & ~(inputs[81]);
    assign layer0_outputs[2348] = inputs[278];
    assign layer0_outputs[2349] = ~(inputs[323]);
    assign layer0_outputs[2350] = (inputs[266]) | (inputs[0]);
    assign layer0_outputs[2351] = ~((inputs[362]) ^ (inputs[304]));
    assign layer0_outputs[2352] = 1'b0;
    assign layer0_outputs[2353] = ~(inputs[291]);
    assign layer0_outputs[2354] = (inputs[335]) | (inputs[378]);
    assign layer0_outputs[2355] = ~((inputs[236]) | (inputs[58]));
    assign layer0_outputs[2356] = ~(inputs[291]);
    assign layer0_outputs[2357] = (inputs[237]) ^ (inputs[59]);
    assign layer0_outputs[2358] = (inputs[397]) | (inputs[247]);
    assign layer0_outputs[2359] = ~((inputs[35]) ^ (inputs[113]));
    assign layer0_outputs[2360] = ~(inputs[377]);
    assign layer0_outputs[2361] = ~(inputs[276]);
    assign layer0_outputs[2362] = ~(inputs[230]);
    assign layer0_outputs[2363] = inputs[128];
    assign layer0_outputs[2364] = ~(inputs[138]);
    assign layer0_outputs[2365] = (inputs[184]) | (inputs[397]);
    assign layer0_outputs[2366] = ~(inputs[322]) | (inputs[177]);
    assign layer0_outputs[2367] = (inputs[50]) & ~(inputs[303]);
    assign layer0_outputs[2368] = ~(inputs[339]) | (inputs[76]);
    assign layer0_outputs[2369] = ~((inputs[371]) & (inputs[224]));
    assign layer0_outputs[2370] = ~((inputs[318]) ^ (inputs[30]));
    assign layer0_outputs[2371] = inputs[230];
    assign layer0_outputs[2372] = ~(inputs[301]);
    assign layer0_outputs[2373] = ~((inputs[377]) ^ (inputs[19]));
    assign layer0_outputs[2374] = inputs[356];
    assign layer0_outputs[2375] = (inputs[322]) & (inputs[134]);
    assign layer0_outputs[2376] = ~(inputs[182]);
    assign layer0_outputs[2377] = ~(inputs[143]);
    assign layer0_outputs[2378] = ~(inputs[342]);
    assign layer0_outputs[2379] = (inputs[132]) & (inputs[385]);
    assign layer0_outputs[2380] = (inputs[53]) & (inputs[68]);
    assign layer0_outputs[2381] = inputs[377];
    assign layer0_outputs[2382] = (inputs[20]) ^ (inputs[36]);
    assign layer0_outputs[2383] = (inputs[218]) & ~(inputs[11]);
    assign layer0_outputs[2384] = ~(inputs[58]);
    assign layer0_outputs[2385] = inputs[57];
    assign layer0_outputs[2386] = ~((inputs[394]) & (inputs[354]));
    assign layer0_outputs[2387] = (inputs[358]) | (inputs[154]);
    assign layer0_outputs[2388] = (inputs[4]) | (inputs[341]);
    assign layer0_outputs[2389] = ~((inputs[387]) | (inputs[263]));
    assign layer0_outputs[2390] = inputs[324];
    assign layer0_outputs[2391] = ~((inputs[156]) | (inputs[67]));
    assign layer0_outputs[2392] = inputs[287];
    assign layer0_outputs[2393] = ~((inputs[272]) | (inputs[221]));
    assign layer0_outputs[2394] = ~((inputs[334]) | (inputs[195]));
    assign layer0_outputs[2395] = (inputs[16]) | (inputs[300]);
    assign layer0_outputs[2396] = ~(inputs[394]) | (inputs[60]);
    assign layer0_outputs[2397] = ~(inputs[71]);
    assign layer0_outputs[2398] = ~((inputs[172]) ^ (inputs[338]));
    assign layer0_outputs[2399] = ~((inputs[182]) | (inputs[169]));
    assign layer0_outputs[2400] = ~(inputs[202]);
    assign layer0_outputs[2401] = ~(inputs[112]) | (inputs[334]);
    assign layer0_outputs[2402] = ~((inputs[304]) | (inputs[290]));
    assign layer0_outputs[2403] = ~(inputs[230]);
    assign layer0_outputs[2404] = ~(inputs[229]);
    assign layer0_outputs[2405] = (inputs[397]) | (inputs[111]);
    assign layer0_outputs[2406] = ~((inputs[162]) | (inputs[294]));
    assign layer0_outputs[2407] = inputs[224];
    assign layer0_outputs[2408] = ~(inputs[8]) | (inputs[251]);
    assign layer0_outputs[2409] = inputs[40];
    assign layer0_outputs[2410] = ~(inputs[273]) | (inputs[1]);
    assign layer0_outputs[2411] = ~(inputs[333]);
    assign layer0_outputs[2412] = (inputs[284]) ^ (inputs[170]);
    assign layer0_outputs[2413] = ~((inputs[1]) & (inputs[190]));
    assign layer0_outputs[2414] = inputs[103];
    assign layer0_outputs[2415] = ~(inputs[57]) | (inputs[206]);
    assign layer0_outputs[2416] = ~(inputs[150]) | (inputs[313]);
    assign layer0_outputs[2417] = (inputs[239]) | (inputs[44]);
    assign layer0_outputs[2418] = ~(inputs[45]) | (inputs[301]);
    assign layer0_outputs[2419] = inputs[201];
    assign layer0_outputs[2420] = ~(inputs[291]) | (inputs[364]);
    assign layer0_outputs[2421] = (inputs[78]) | (inputs[1]);
    assign layer0_outputs[2422] = inputs[103];
    assign layer0_outputs[2423] = ~(inputs[38]);
    assign layer0_outputs[2424] = (inputs[17]) & ~(inputs[102]);
    assign layer0_outputs[2425] = ~((inputs[50]) | (inputs[159]));
    assign layer0_outputs[2426] = (inputs[393]) | (inputs[311]);
    assign layer0_outputs[2427] = ~(inputs[176]);
    assign layer0_outputs[2428] = inputs[310];
    assign layer0_outputs[2429] = ~(inputs[106]);
    assign layer0_outputs[2430] = (inputs[282]) ^ (inputs[377]);
    assign layer0_outputs[2431] = ~(inputs[241]);
    assign layer0_outputs[2432] = (inputs[110]) & ~(inputs[238]);
    assign layer0_outputs[2433] = inputs[206];
    assign layer0_outputs[2434] = inputs[374];
    assign layer0_outputs[2435] = inputs[31];
    assign layer0_outputs[2436] = (inputs[214]) | (inputs[109]);
    assign layer0_outputs[2437] = inputs[131];
    assign layer0_outputs[2438] = (inputs[132]) & ~(inputs[239]);
    assign layer0_outputs[2439] = inputs[351];
    assign layer0_outputs[2440] = ~((inputs[138]) & (inputs[342]));
    assign layer0_outputs[2441] = ~((inputs[185]) | (inputs[178]));
    assign layer0_outputs[2442] = (inputs[299]) | (inputs[389]);
    assign layer0_outputs[2443] = ~(inputs[193]) | (inputs[199]);
    assign layer0_outputs[2444] = ~((inputs[343]) | (inputs[296]));
    assign layer0_outputs[2445] = (inputs[352]) & ~(inputs[34]);
    assign layer0_outputs[2446] = ~((inputs[347]) | (inputs[355]));
    assign layer0_outputs[2447] = (inputs[99]) | (inputs[365]);
    assign layer0_outputs[2448] = (inputs[81]) | (inputs[173]);
    assign layer0_outputs[2449] = (inputs[240]) | (inputs[187]);
    assign layer0_outputs[2450] = inputs[90];
    assign layer0_outputs[2451] = (inputs[263]) | (inputs[39]);
    assign layer0_outputs[2452] = ~((inputs[12]) ^ (inputs[89]));
    assign layer0_outputs[2453] = ~(inputs[347]);
    assign layer0_outputs[2454] = ~(inputs[54]) | (inputs[301]);
    assign layer0_outputs[2455] = ~(inputs[216]) | (inputs[379]);
    assign layer0_outputs[2456] = (inputs[137]) ^ (inputs[282]);
    assign layer0_outputs[2457] = ~((inputs[192]) ^ (inputs[327]));
    assign layer0_outputs[2458] = inputs[179];
    assign layer0_outputs[2459] = 1'b0;
    assign layer0_outputs[2460] = (inputs[48]) ^ (inputs[351]);
    assign layer0_outputs[2461] = ~((inputs[261]) ^ (inputs[288]));
    assign layer0_outputs[2462] = ~(inputs[53]);
    assign layer0_outputs[2463] = (inputs[93]) & ~(inputs[342]);
    assign layer0_outputs[2464] = (inputs[330]) & ~(inputs[127]);
    assign layer0_outputs[2465] = (inputs[2]) ^ (inputs[176]);
    assign layer0_outputs[2466] = ~((inputs[57]) | (inputs[252]));
    assign layer0_outputs[2467] = (inputs[170]) & ~(inputs[299]);
    assign layer0_outputs[2468] = ~(inputs[128]);
    assign layer0_outputs[2469] = (inputs[326]) ^ (inputs[384]);
    assign layer0_outputs[2470] = inputs[209];
    assign layer0_outputs[2471] = ~(inputs[383]);
    assign layer0_outputs[2472] = (inputs[169]) | (inputs[169]);
    assign layer0_outputs[2473] = ~((inputs[395]) & (inputs[377]));
    assign layer0_outputs[2474] = (inputs[141]) | (inputs[187]);
    assign layer0_outputs[2475] = ~(inputs[256]);
    assign layer0_outputs[2476] = ~(inputs[149]);
    assign layer0_outputs[2477] = inputs[384];
    assign layer0_outputs[2478] = ~(inputs[33]);
    assign layer0_outputs[2479] = ~(inputs[49]);
    assign layer0_outputs[2480] = inputs[123];
    assign layer0_outputs[2481] = (inputs[246]) | (inputs[247]);
    assign layer0_outputs[2482] = ~(inputs[250]);
    assign layer0_outputs[2483] = ~((inputs[259]) ^ (inputs[98]));
    assign layer0_outputs[2484] = inputs[337];
    assign layer0_outputs[2485] = ~(inputs[51]) | (inputs[316]);
    assign layer0_outputs[2486] = (inputs[315]) & ~(inputs[181]);
    assign layer0_outputs[2487] = ~(inputs[28]);
    assign layer0_outputs[2488] = (inputs[249]) ^ (inputs[360]);
    assign layer0_outputs[2489] = inputs[183];
    assign layer0_outputs[2490] = ~(inputs[11]);
    assign layer0_outputs[2491] = ~(inputs[270]);
    assign layer0_outputs[2492] = ~((inputs[7]) | (inputs[146]));
    assign layer0_outputs[2493] = ~((inputs[231]) ^ (inputs[359]));
    assign layer0_outputs[2494] = ~((inputs[195]) | (inputs[68]));
    assign layer0_outputs[2495] = ~(inputs[109]) | (inputs[235]);
    assign layer0_outputs[2496] = (inputs[94]) | (inputs[68]);
    assign layer0_outputs[2497] = (inputs[90]) & ~(inputs[159]);
    assign layer0_outputs[2498] = (inputs[196]) | (inputs[140]);
    assign layer0_outputs[2499] = ~(inputs[358]);
    assign outputs[0] = (layer0_outputs[1719]) & ~(layer0_outputs[1616]);
    assign outputs[1] = ~(layer0_outputs[1891]);
    assign outputs[2] = ~(layer0_outputs[1352]);
    assign outputs[3] = ~((layer0_outputs[2137]) & (layer0_outputs[2011]));
    assign outputs[4] = layer0_outputs[1378];
    assign outputs[5] = (layer0_outputs[104]) | (layer0_outputs[1167]);
    assign outputs[6] = (layer0_outputs[1372]) & ~(layer0_outputs[192]);
    assign outputs[7] = (layer0_outputs[2463]) & ~(layer0_outputs[2211]);
    assign outputs[8] = layer0_outputs[2128];
    assign outputs[9] = (layer0_outputs[2025]) | (layer0_outputs[281]);
    assign outputs[10] = (layer0_outputs[1942]) & (layer0_outputs[349]);
    assign outputs[11] = ~(layer0_outputs[1944]) | (layer0_outputs[1324]);
    assign outputs[12] = ~(layer0_outputs[456]);
    assign outputs[13] = ~(layer0_outputs[1882]);
    assign outputs[14] = ~(layer0_outputs[2249]) | (layer0_outputs[935]);
    assign outputs[15] = (layer0_outputs[308]) & (layer0_outputs[157]);
    assign outputs[16] = ~((layer0_outputs[2087]) | (layer0_outputs[1252]));
    assign outputs[17] = (layer0_outputs[1201]) ^ (layer0_outputs[2295]);
    assign outputs[18] = layer0_outputs[2145];
    assign outputs[19] = (layer0_outputs[2196]) ^ (layer0_outputs[302]);
    assign outputs[20] = ~(layer0_outputs[1457]);
    assign outputs[21] = layer0_outputs[1318];
    assign outputs[22] = ~(layer0_outputs[723]);
    assign outputs[23] = ~((layer0_outputs[1399]) | (layer0_outputs[825]));
    assign outputs[24] = ~(layer0_outputs[1478]);
    assign outputs[25] = ~((layer0_outputs[1807]) ^ (layer0_outputs[2111]));
    assign outputs[26] = ~(layer0_outputs[986]);
    assign outputs[27] = ~((layer0_outputs[180]) & (layer0_outputs[1515]));
    assign outputs[28] = layer0_outputs[70];
    assign outputs[29] = (layer0_outputs[1529]) & ~(layer0_outputs[505]);
    assign outputs[30] = layer0_outputs[783];
    assign outputs[31] = ~((layer0_outputs[2459]) ^ (layer0_outputs[2107]));
    assign outputs[32] = (layer0_outputs[137]) & ~(layer0_outputs[2143]);
    assign outputs[33] = layer0_outputs[1400];
    assign outputs[34] = ~(layer0_outputs[31]) | (layer0_outputs[2383]);
    assign outputs[35] = ~((layer0_outputs[614]) ^ (layer0_outputs[1221]));
    assign outputs[36] = (layer0_outputs[2088]) & (layer0_outputs[2323]);
    assign outputs[37] = (layer0_outputs[2197]) & (layer0_outputs[278]);
    assign outputs[38] = layer0_outputs[2104];
    assign outputs[39] = (layer0_outputs[803]) & (layer0_outputs[1827]);
    assign outputs[40] = (layer0_outputs[365]) | (layer0_outputs[996]);
    assign outputs[41] = (layer0_outputs[2312]) & (layer0_outputs[1956]);
    assign outputs[42] = ~(layer0_outputs[1389]);
    assign outputs[43] = (layer0_outputs[1143]) & ~(layer0_outputs[871]);
    assign outputs[44] = layer0_outputs[354];
    assign outputs[45] = ~((layer0_outputs[1357]) ^ (layer0_outputs[1742]));
    assign outputs[46] = ~((layer0_outputs[318]) | (layer0_outputs[75]));
    assign outputs[47] = ~(layer0_outputs[453]) | (layer0_outputs[1994]);
    assign outputs[48] = layer0_outputs[2496];
    assign outputs[49] = (layer0_outputs[2169]) & ~(layer0_outputs[1903]);
    assign outputs[50] = ~(layer0_outputs[2039]);
    assign outputs[51] = (layer0_outputs[1401]) & (layer0_outputs[2080]);
    assign outputs[52] = ~((layer0_outputs[2189]) | (layer0_outputs[598]));
    assign outputs[53] = ~((layer0_outputs[2110]) ^ (layer0_outputs[666]));
    assign outputs[54] = ~((layer0_outputs[2456]) | (layer0_outputs[2470]));
    assign outputs[55] = layer0_outputs[928];
    assign outputs[56] = ~(layer0_outputs[1180]) | (layer0_outputs[1411]);
    assign outputs[57] = ~((layer0_outputs[458]) | (layer0_outputs[674]));
    assign outputs[58] = ~(layer0_outputs[1505]);
    assign outputs[59] = ~(layer0_outputs[1140]) | (layer0_outputs[836]);
    assign outputs[60] = ~((layer0_outputs[544]) ^ (layer0_outputs[1261]));
    assign outputs[61] = layer0_outputs[207];
    assign outputs[62] = (layer0_outputs[977]) & ~(layer0_outputs[1697]);
    assign outputs[63] = ~((layer0_outputs[1825]) | (layer0_outputs[958]));
    assign outputs[64] = ~((layer0_outputs[1002]) ^ (layer0_outputs[1916]));
    assign outputs[65] = (layer0_outputs[1464]) | (layer0_outputs[668]);
    assign outputs[66] = (layer0_outputs[1463]) & ~(layer0_outputs[1192]);
    assign outputs[67] = layer0_outputs[154];
    assign outputs[68] = ~(layer0_outputs[737]) | (layer0_outputs[66]);
    assign outputs[69] = layer0_outputs[1758];
    assign outputs[70] = ~(layer0_outputs[629]);
    assign outputs[71] = (layer0_outputs[1411]) & ~(layer0_outputs[1184]);
    assign outputs[72] = ~(layer0_outputs[776]) | (layer0_outputs[504]);
    assign outputs[73] = ~(layer0_outputs[2358]) | (layer0_outputs[1455]);
    assign outputs[74] = ~(layer0_outputs[2069]);
    assign outputs[75] = (layer0_outputs[676]) & ~(layer0_outputs[884]);
    assign outputs[76] = (layer0_outputs[20]) | (layer0_outputs[524]);
    assign outputs[77] = ~(layer0_outputs[400]);
    assign outputs[78] = (layer0_outputs[2049]) | (layer0_outputs[653]);
    assign outputs[79] = ~((layer0_outputs[2460]) ^ (layer0_outputs[984]));
    assign outputs[80] = ~(layer0_outputs[1200]);
    assign outputs[81] = (layer0_outputs[1583]) | (layer0_outputs[1659]);
    assign outputs[82] = (layer0_outputs[1615]) & ~(layer0_outputs[2199]);
    assign outputs[83] = ~(layer0_outputs[2303]) | (layer0_outputs[798]);
    assign outputs[84] = ~((layer0_outputs[370]) ^ (layer0_outputs[2102]));
    assign outputs[85] = ~(layer0_outputs[1774]) | (layer0_outputs[277]);
    assign outputs[86] = layer0_outputs[165];
    assign outputs[87] = layer0_outputs[2362];
    assign outputs[88] = layer0_outputs[2362];
    assign outputs[89] = ~((layer0_outputs[1364]) & (layer0_outputs[1273]));
    assign outputs[90] = ~((layer0_outputs[2105]) | (layer0_outputs[1363]));
    assign outputs[91] = (layer0_outputs[1575]) & (layer0_outputs[670]);
    assign outputs[92] = (layer0_outputs[1414]) & (layer0_outputs[1293]);
    assign outputs[93] = layer0_outputs[1164];
    assign outputs[94] = layer0_outputs[2404];
    assign outputs[95] = ~((layer0_outputs[419]) & (layer0_outputs[1774]));
    assign outputs[96] = layer0_outputs[1444];
    assign outputs[97] = ~(layer0_outputs[706]);
    assign outputs[98] = layer0_outputs[1879];
    assign outputs[99] = layer0_outputs[229];
    assign outputs[100] = (layer0_outputs[1818]) & (layer0_outputs[2269]);
    assign outputs[101] = (layer0_outputs[956]) ^ (layer0_outputs[1794]);
    assign outputs[102] = ~((layer0_outputs[203]) & (layer0_outputs[1074]));
    assign outputs[103] = ~((layer0_outputs[1531]) ^ (layer0_outputs[2]));
    assign outputs[104] = layer0_outputs[1026];
    assign outputs[105] = layer0_outputs[461];
    assign outputs[106] = ~(layer0_outputs[1228]);
    assign outputs[107] = ~(layer0_outputs[1419]);
    assign outputs[108] = ~((layer0_outputs[1894]) ^ (layer0_outputs[1345]));
    assign outputs[109] = ~(layer0_outputs[242]);
    assign outputs[110] = ~(layer0_outputs[2182]);
    assign outputs[111] = (layer0_outputs[1669]) & ~(layer0_outputs[644]);
    assign outputs[112] = (layer0_outputs[1646]) ^ (layer0_outputs[198]);
    assign outputs[113] = ~(layer0_outputs[280]) | (layer0_outputs[731]);
    assign outputs[114] = layer0_outputs[2419];
    assign outputs[115] = (layer0_outputs[2396]) & ~(layer0_outputs[550]);
    assign outputs[116] = layer0_outputs[1251];
    assign outputs[117] = layer0_outputs[2458];
    assign outputs[118] = ~((layer0_outputs[1235]) ^ (layer0_outputs[1210]));
    assign outputs[119] = ~(layer0_outputs[2243]);
    assign outputs[120] = (layer0_outputs[1114]) ^ (layer0_outputs[2261]);
    assign outputs[121] = ~((layer0_outputs[1997]) & (layer0_outputs[261]));
    assign outputs[122] = layer0_outputs[369];
    assign outputs[123] = ~(layer0_outputs[750]);
    assign outputs[124] = (layer0_outputs[701]) | (layer0_outputs[1740]);
    assign outputs[125] = layer0_outputs[2493];
    assign outputs[126] = (layer0_outputs[1120]) & (layer0_outputs[1117]);
    assign outputs[127] = (layer0_outputs[942]) & (layer0_outputs[2266]);
    assign outputs[128] = ~((layer0_outputs[1666]) & (layer0_outputs[2238]));
    assign outputs[129] = ~((layer0_outputs[1043]) | (layer0_outputs[1458]));
    assign outputs[130] = ~(layer0_outputs[752]);
    assign outputs[131] = layer0_outputs[894];
    assign outputs[132] = ~(layer0_outputs[1745]);
    assign outputs[133] = ~(layer0_outputs[1256]);
    assign outputs[134] = (layer0_outputs[439]) & ~(layer0_outputs[2185]);
    assign outputs[135] = ~((layer0_outputs[334]) | (layer0_outputs[376]));
    assign outputs[136] = (layer0_outputs[1949]) | (layer0_outputs[2191]);
    assign outputs[137] = (layer0_outputs[2140]) & ~(layer0_outputs[2022]);
    assign outputs[138] = layer0_outputs[733];
    assign outputs[139] = ~(layer0_outputs[1518]) | (layer0_outputs[2236]);
    assign outputs[140] = (layer0_outputs[965]) | (layer0_outputs[1883]);
    assign outputs[141] = (layer0_outputs[279]) & ~(layer0_outputs[312]);
    assign outputs[142] = (layer0_outputs[479]) & ~(layer0_outputs[1195]);
    assign outputs[143] = ~((layer0_outputs[1854]) & (layer0_outputs[403]));
    assign outputs[144] = layer0_outputs[785];
    assign outputs[145] = ~(layer0_outputs[2332]);
    assign outputs[146] = ~(layer0_outputs[2020]) | (layer0_outputs[190]);
    assign outputs[147] = (layer0_outputs[867]) & ~(layer0_outputs[1856]);
    assign outputs[148] = ~((layer0_outputs[1534]) & (layer0_outputs[1385]));
    assign outputs[149] = ~((layer0_outputs[2308]) ^ (layer0_outputs[661]));
    assign outputs[150] = ~((layer0_outputs[2108]) | (layer0_outputs[1631]));
    assign outputs[151] = ~((layer0_outputs[918]) | (layer0_outputs[961]));
    assign outputs[152] = (layer0_outputs[770]) & (layer0_outputs[640]);
    assign outputs[153] = ~(layer0_outputs[752]);
    assign outputs[154] = (layer0_outputs[2130]) | (layer0_outputs[2282]);
    assign outputs[155] = (layer0_outputs[69]) & ~(layer0_outputs[27]);
    assign outputs[156] = (layer0_outputs[301]) & ~(layer0_outputs[1458]);
    assign outputs[157] = ~((layer0_outputs[1414]) ^ (layer0_outputs[923]));
    assign outputs[158] = (layer0_outputs[2210]) ^ (layer0_outputs[59]);
    assign outputs[159] = ~((layer0_outputs[723]) | (layer0_outputs[1427]));
    assign outputs[160] = ~(layer0_outputs[1359]);
    assign outputs[161] = (layer0_outputs[910]) & ~(layer0_outputs[1056]);
    assign outputs[162] = ~(layer0_outputs[1334]);
    assign outputs[163] = ~((layer0_outputs[323]) & (layer0_outputs[332]));
    assign outputs[164] = (layer0_outputs[997]) & (layer0_outputs[1286]);
    assign outputs[165] = ~(layer0_outputs[1720]) | (layer0_outputs[1123]);
    assign outputs[166] = ~(layer0_outputs[210]);
    assign outputs[167] = (layer0_outputs[104]) & ~(layer0_outputs[2173]);
    assign outputs[168] = layer0_outputs[1550];
    assign outputs[169] = (layer0_outputs[2365]) & ~(layer0_outputs[363]);
    assign outputs[170] = layer0_outputs[510];
    assign outputs[171] = (layer0_outputs[1932]) & (layer0_outputs[234]);
    assign outputs[172] = ~(layer0_outputs[1182]);
    assign outputs[173] = layer0_outputs[379];
    assign outputs[174] = layer0_outputs[1316];
    assign outputs[175] = layer0_outputs[98];
    assign outputs[176] = ~(layer0_outputs[1566]);
    assign outputs[177] = ~((layer0_outputs[1088]) ^ (layer0_outputs[217]));
    assign outputs[178] = ~((layer0_outputs[1434]) & (layer0_outputs[1060]));
    assign outputs[179] = layer0_outputs[1096];
    assign outputs[180] = (layer0_outputs[2030]) ^ (layer0_outputs[1480]);
    assign outputs[181] = ~(layer0_outputs[1397]) | (layer0_outputs[792]);
    assign outputs[182] = ~((layer0_outputs[1101]) | (layer0_outputs[635]));
    assign outputs[183] = (layer0_outputs[78]) & (layer0_outputs[583]);
    assign outputs[184] = layer0_outputs[1896];
    assign outputs[185] = layer0_outputs[1826];
    assign outputs[186] = ~((layer0_outputs[2436]) ^ (layer0_outputs[1983]));
    assign outputs[187] = ~(layer0_outputs[2441]) | (layer0_outputs[2121]);
    assign outputs[188] = ~(layer0_outputs[2475]) | (layer0_outputs[1379]);
    assign outputs[189] = (layer0_outputs[618]) ^ (layer0_outputs[35]);
    assign outputs[190] = (layer0_outputs[2247]) ^ (layer0_outputs[1164]);
    assign outputs[191] = (layer0_outputs[1671]) ^ (layer0_outputs[788]);
    assign outputs[192] = (layer0_outputs[697]) & (layer0_outputs[2015]);
    assign outputs[193] = layer0_outputs[753];
    assign outputs[194] = (layer0_outputs[1109]) & ~(layer0_outputs[897]);
    assign outputs[195] = layer0_outputs[1156];
    assign outputs[196] = layer0_outputs[758];
    assign outputs[197] = (layer0_outputs[1685]) & (layer0_outputs[2482]);
    assign outputs[198] = layer0_outputs[95];
    assign outputs[199] = layer0_outputs[1609];
    assign outputs[200] = ~((layer0_outputs[1284]) | (layer0_outputs[588]));
    assign outputs[201] = (layer0_outputs[553]) & (layer0_outputs[934]);
    assign outputs[202] = ~(layer0_outputs[1046]);
    assign outputs[203] = ~(layer0_outputs[830]);
    assign outputs[204] = ~((layer0_outputs[985]) ^ (layer0_outputs[786]));
    assign outputs[205] = ~(layer0_outputs[810]);
    assign outputs[206] = ~(layer0_outputs[1033]);
    assign outputs[207] = (layer0_outputs[1357]) & ~(layer0_outputs[1059]);
    assign outputs[208] = ~(layer0_outputs[1717]);
    assign outputs[209] = ~((layer0_outputs[876]) ^ (layer0_outputs[1337]));
    assign outputs[210] = ~(layer0_outputs[564]) | (layer0_outputs[48]);
    assign outputs[211] = ~(layer0_outputs[1692]);
    assign outputs[212] = ~(layer0_outputs[1304]) | (layer0_outputs[1222]);
    assign outputs[213] = ~((layer0_outputs[2020]) & (layer0_outputs[1544]));
    assign outputs[214] = layer0_outputs[2248];
    assign outputs[215] = ~(layer0_outputs[2344]);
    assign outputs[216] = (layer0_outputs[1662]) & ~(layer0_outputs[273]);
    assign outputs[217] = ~(layer0_outputs[1975]);
    assign outputs[218] = layer0_outputs[816];
    assign outputs[219] = layer0_outputs[1298];
    assign outputs[220] = ~(layer0_outputs[1993]);
    assign outputs[221] = ~((layer0_outputs[1307]) | (layer0_outputs[210]));
    assign outputs[222] = ~(layer0_outputs[1199]) | (layer0_outputs[1743]);
    assign outputs[223] = ~(layer0_outputs[573]);
    assign outputs[224] = layer0_outputs[2122];
    assign outputs[225] = ~((layer0_outputs[2183]) | (layer0_outputs[1399]));
    assign outputs[226] = ~(layer0_outputs[573]);
    assign outputs[227] = ~(layer0_outputs[1367]);
    assign outputs[228] = (layer0_outputs[215]) ^ (layer0_outputs[1087]);
    assign outputs[229] = ~(layer0_outputs[1485]);
    assign outputs[230] = layer0_outputs[2074];
    assign outputs[231] = (layer0_outputs[801]) & ~(layer0_outputs[1522]);
    assign outputs[232] = (layer0_outputs[111]) ^ (layer0_outputs[566]);
    assign outputs[233] = (layer0_outputs[1051]) & (layer0_outputs[930]);
    assign outputs[234] = (layer0_outputs[2017]) & ~(layer0_outputs[417]);
    assign outputs[235] = ~((layer0_outputs[1354]) ^ (layer0_outputs[1310]));
    assign outputs[236] = ~((layer0_outputs[2075]) ^ (layer0_outputs[1431]));
    assign outputs[237] = ~((layer0_outputs[293]) ^ (layer0_outputs[1806]));
    assign outputs[238] = (layer0_outputs[2384]) & (layer0_outputs[996]);
    assign outputs[239] = layer0_outputs[396];
    assign outputs[240] = ~(layer0_outputs[1579]) | (layer0_outputs[1550]);
    assign outputs[241] = ~(layer0_outputs[2066]);
    assign outputs[242] = (layer0_outputs[1601]) ^ (layer0_outputs[1779]);
    assign outputs[243] = ~((layer0_outputs[1537]) | (layer0_outputs[373]));
    assign outputs[244] = (layer0_outputs[1260]) & ~(layer0_outputs[1941]);
    assign outputs[245] = ~(layer0_outputs[1198]);
    assign outputs[246] = ~((layer0_outputs[1850]) ^ (layer0_outputs[1526]));
    assign outputs[247] = ~(layer0_outputs[236]);
    assign outputs[248] = layer0_outputs[2065];
    assign outputs[249] = (layer0_outputs[448]) & (layer0_outputs[963]);
    assign outputs[250] = (layer0_outputs[176]) & ~(layer0_outputs[1141]);
    assign outputs[251] = layer0_outputs[2306];
    assign outputs[252] = (layer0_outputs[1305]) & (layer0_outputs[1078]);
    assign outputs[253] = (layer0_outputs[399]) ^ (layer0_outputs[641]);
    assign outputs[254] = (layer0_outputs[874]) & ~(layer0_outputs[1931]);
    assign outputs[255] = (layer0_outputs[2271]) & ~(layer0_outputs[255]);
    assign outputs[256] = ~(layer0_outputs[1603]);
    assign outputs[257] = ~(layer0_outputs[1326]);
    assign outputs[258] = (layer0_outputs[130]) & ~(layer0_outputs[243]);
    assign outputs[259] = (layer0_outputs[219]) & ~(layer0_outputs[585]);
    assign outputs[260] = (layer0_outputs[2163]) & ~(layer0_outputs[1501]);
    assign outputs[261] = (layer0_outputs[2369]) & (layer0_outputs[602]);
    assign outputs[262] = (layer0_outputs[2208]) & ~(layer0_outputs[1620]);
    assign outputs[263] = (layer0_outputs[2434]) & ~(layer0_outputs[596]);
    assign outputs[264] = (layer0_outputs[1987]) & (layer0_outputs[1966]);
    assign outputs[265] = ~((layer0_outputs[2016]) ^ (layer0_outputs[1885]));
    assign outputs[266] = (layer0_outputs[2431]) & ~(layer0_outputs[1617]);
    assign outputs[267] = ~((layer0_outputs[1041]) | (layer0_outputs[253]));
    assign outputs[268] = (layer0_outputs[684]) & ~(layer0_outputs[950]);
    assign outputs[269] = (layer0_outputs[2472]) & ~(layer0_outputs[1004]);
    assign outputs[270] = 1'b0;
    assign outputs[271] = (layer0_outputs[1066]) & ~(layer0_outputs[54]);
    assign outputs[272] = (layer0_outputs[844]) ^ (layer0_outputs[1617]);
    assign outputs[273] = (layer0_outputs[2290]) & (layer0_outputs[228]);
    assign outputs[274] = ~((layer0_outputs[317]) | (layer0_outputs[391]));
    assign outputs[275] = (layer0_outputs[1564]) & (layer0_outputs[803]);
    assign outputs[276] = (layer0_outputs[801]) ^ (layer0_outputs[101]);
    assign outputs[277] = ~((layer0_outputs[951]) ^ (layer0_outputs[1282]));
    assign outputs[278] = (layer0_outputs[1589]) & ~(layer0_outputs[2417]);
    assign outputs[279] = ~((layer0_outputs[789]) ^ (layer0_outputs[2315]));
    assign outputs[280] = ~(layer0_outputs[1286]);
    assign outputs[281] = ~(layer0_outputs[2001]) | (layer0_outputs[2494]);
    assign outputs[282] = (layer0_outputs[1543]) & (layer0_outputs[962]);
    assign outputs[283] = (layer0_outputs[1635]) ^ (layer0_outputs[1802]);
    assign outputs[284] = (layer0_outputs[2370]) & (layer0_outputs[1721]);
    assign outputs[285] = (layer0_outputs[1551]) & ~(layer0_outputs[995]);
    assign outputs[286] = ~((layer0_outputs[2116]) | (layer0_outputs[2458]));
    assign outputs[287] = (layer0_outputs[756]) & ~(layer0_outputs[2399]);
    assign outputs[288] = (layer0_outputs[1502]) & ~(layer0_outputs[1315]);
    assign outputs[289] = (layer0_outputs[122]) & (layer0_outputs[629]);
    assign outputs[290] = ~(layer0_outputs[1133]);
    assign outputs[291] = (layer0_outputs[839]) & (layer0_outputs[249]);
    assign outputs[292] = ~(layer0_outputs[290]);
    assign outputs[293] = (layer0_outputs[1866]) & (layer0_outputs[710]);
    assign outputs[294] = ~(layer0_outputs[599]) | (layer0_outputs[1334]);
    assign outputs[295] = ~(layer0_outputs[1288]);
    assign outputs[296] = layer0_outputs[1445];
    assign outputs[297] = ~((layer0_outputs[479]) | (layer0_outputs[1986]));
    assign outputs[298] = (layer0_outputs[2434]) | (layer0_outputs[170]);
    assign outputs[299] = (layer0_outputs[709]) & ~(layer0_outputs[2421]);
    assign outputs[300] = ~(layer0_outputs[2166]);
    assign outputs[301] = (layer0_outputs[1584]) & (layer0_outputs[863]);
    assign outputs[302] = (layer0_outputs[1127]) ^ (layer0_outputs[514]);
    assign outputs[303] = ~((layer0_outputs[939]) ^ (layer0_outputs[101]));
    assign outputs[304] = (layer0_outputs[238]) & ~(layer0_outputs[1510]);
    assign outputs[305] = (layer0_outputs[1521]) & ~(layer0_outputs[959]);
    assign outputs[306] = (layer0_outputs[589]) & (layer0_outputs[2148]);
    assign outputs[307] = ~((layer0_outputs[1134]) | (layer0_outputs[858]));
    assign outputs[308] = ~(layer0_outputs[2416]);
    assign outputs[309] = layer0_outputs[1465];
    assign outputs[310] = (layer0_outputs[416]) & ~(layer0_outputs[1427]);
    assign outputs[311] = (layer0_outputs[2425]) & (layer0_outputs[564]);
    assign outputs[312] = (layer0_outputs[2243]) & ~(layer0_outputs[562]);
    assign outputs[313] = (layer0_outputs[2024]) ^ (layer0_outputs[1078]);
    assign outputs[314] = layer0_outputs[2337];
    assign outputs[315] = ~((layer0_outputs[329]) | (layer0_outputs[140]));
    assign outputs[316] = (layer0_outputs[1955]) & (layer0_outputs[2477]);
    assign outputs[317] = (layer0_outputs[2029]) & ~(layer0_outputs[1627]);
    assign outputs[318] = (layer0_outputs[2376]) & (layer0_outputs[162]);
    assign outputs[319] = (layer0_outputs[2437]) & ~(layer0_outputs[1004]);
    assign outputs[320] = (layer0_outputs[506]) & ~(layer0_outputs[1610]);
    assign outputs[321] = ~((layer0_outputs[1467]) | (layer0_outputs[599]));
    assign outputs[322] = (layer0_outputs[1711]) & ~(layer0_outputs[1979]);
    assign outputs[323] = (layer0_outputs[902]) & ~(layer0_outputs[1029]);
    assign outputs[324] = layer0_outputs[145];
    assign outputs[325] = (layer0_outputs[1083]) & ~(layer0_outputs[1673]);
    assign outputs[326] = ~((layer0_outputs[390]) ^ (layer0_outputs[1349]));
    assign outputs[327] = ~(layer0_outputs[593]) | (layer0_outputs[139]);
    assign outputs[328] = (layer0_outputs[1024]) & (layer0_outputs[1493]);
    assign outputs[329] = ~((layer0_outputs[1836]) ^ (layer0_outputs[530]));
    assign outputs[330] = (layer0_outputs[1410]) & ~(layer0_outputs[1800]);
    assign outputs[331] = (layer0_outputs[1023]) | (layer0_outputs[1549]);
    assign outputs[332] = (layer0_outputs[463]) & ~(layer0_outputs[1936]);
    assign outputs[333] = ~(layer0_outputs[598]);
    assign outputs[334] = (layer0_outputs[205]) & ~(layer0_outputs[168]);
    assign outputs[335] = (layer0_outputs[1986]) ^ (layer0_outputs[2157]);
    assign outputs[336] = ~((layer0_outputs[1565]) | (layer0_outputs[1560]));
    assign outputs[337] = ~((layer0_outputs[686]) | (layer0_outputs[901]));
    assign outputs[338] = (layer0_outputs[1426]) & ~(layer0_outputs[1310]);
    assign outputs[339] = (layer0_outputs[1975]) & (layer0_outputs[1956]);
    assign outputs[340] = ~((layer0_outputs[66]) | (layer0_outputs[2357]));
    assign outputs[341] = ~((layer0_outputs[2394]) ^ (layer0_outputs[8]));
    assign outputs[342] = (layer0_outputs[975]) & (layer0_outputs[1602]);
    assign outputs[343] = (layer0_outputs[771]) & ~(layer0_outputs[965]);
    assign outputs[344] = layer0_outputs[2149];
    assign outputs[345] = (layer0_outputs[59]) & ~(layer0_outputs[1685]);
    assign outputs[346] = (layer0_outputs[2424]) ^ (layer0_outputs[1037]);
    assign outputs[347] = (layer0_outputs[468]) ^ (layer0_outputs[149]);
    assign outputs[348] = (layer0_outputs[577]) & ~(layer0_outputs[1659]);
    assign outputs[349] = (layer0_outputs[1342]) & (layer0_outputs[2342]);
    assign outputs[350] = (layer0_outputs[1227]) & ~(layer0_outputs[785]);
    assign outputs[351] = (layer0_outputs[2189]) & (layer0_outputs[1433]);
    assign outputs[352] = (layer0_outputs[10]) ^ (layer0_outputs[512]);
    assign outputs[353] = ~((layer0_outputs[967]) ^ (layer0_outputs[1751]));
    assign outputs[354] = ~((layer0_outputs[1910]) | (layer0_outputs[2044]));
    assign outputs[355] = (layer0_outputs[2262]) & (layer0_outputs[1829]);
    assign outputs[356] = ~((layer0_outputs[225]) | (layer0_outputs[1110]));
    assign outputs[357] = ~((layer0_outputs[1504]) | (layer0_outputs[173]));
    assign outputs[358] = (layer0_outputs[415]) & (layer0_outputs[714]);
    assign outputs[359] = (layer0_outputs[1806]) ^ (layer0_outputs[2443]);
    assign outputs[360] = layer0_outputs[2406];
    assign outputs[361] = (layer0_outputs[1539]) ^ (layer0_outputs[1021]);
    assign outputs[362] = (layer0_outputs[1916]) & (layer0_outputs[1756]);
    assign outputs[363] = (layer0_outputs[1165]) & ~(layer0_outputs[1764]);
    assign outputs[364] = (layer0_outputs[834]) & ~(layer0_outputs[1026]);
    assign outputs[365] = (layer0_outputs[1212]) & ~(layer0_outputs[1887]);
    assign outputs[366] = (layer0_outputs[258]) & ~(layer0_outputs[1180]);
    assign outputs[367] = ~((layer0_outputs[1834]) | (layer0_outputs[671]));
    assign outputs[368] = ~((layer0_outputs[2094]) | (layer0_outputs[1189]));
    assign outputs[369] = (layer0_outputs[2306]) & ~(layer0_outputs[123]);
    assign outputs[370] = (layer0_outputs[2408]) & ~(layer0_outputs[2329]);
    assign outputs[371] = 1'b0;
    assign outputs[372] = ~((layer0_outputs[1792]) ^ (layer0_outputs[2028]));
    assign outputs[373] = ~((layer0_outputs[729]) ^ (layer0_outputs[941]));
    assign outputs[374] = (layer0_outputs[2406]) & ~(layer0_outputs[13]);
    assign outputs[375] = ~((layer0_outputs[2451]) | (layer0_outputs[849]));
    assign outputs[376] = (layer0_outputs[1730]) ^ (layer0_outputs[182]);
    assign outputs[377] = (layer0_outputs[2184]) & (layer0_outputs[2174]);
    assign outputs[378] = (layer0_outputs[1906]) & (layer0_outputs[115]);
    assign outputs[379] = ~((layer0_outputs[2442]) | (layer0_outputs[1754]));
    assign outputs[380] = ~((layer0_outputs[1060]) | (layer0_outputs[1962]));
    assign outputs[381] = (layer0_outputs[902]) & ~(layer0_outputs[1709]);
    assign outputs[382] = (layer0_outputs[1679]) & ~(layer0_outputs[289]);
    assign outputs[383] = ~((layer0_outputs[1329]) ^ (layer0_outputs[1515]));
    assign outputs[384] = (layer0_outputs[339]) & ~(layer0_outputs[1082]);
    assign outputs[385] = ~((layer0_outputs[57]) | (layer0_outputs[2253]));
    assign outputs[386] = ~((layer0_outputs[2047]) | (layer0_outputs[605]));
    assign outputs[387] = (layer0_outputs[311]) & (layer0_outputs[1920]);
    assign outputs[388] = (layer0_outputs[627]) & (layer0_outputs[1868]);
    assign outputs[389] = 1'b0;
    assign outputs[390] = ~((layer0_outputs[2281]) | (layer0_outputs[1406]));
    assign outputs[391] = ~((layer0_outputs[2093]) ^ (layer0_outputs[1350]));
    assign outputs[392] = (layer0_outputs[1580]) & ~(layer0_outputs[1965]);
    assign outputs[393] = ~((layer0_outputs[817]) | (layer0_outputs[23]));
    assign outputs[394] = (layer0_outputs[2429]) & (layer0_outputs[1808]);
    assign outputs[395] = ~((layer0_outputs[98]) | (layer0_outputs[681]));
    assign outputs[396] = ~((layer0_outputs[1615]) | (layer0_outputs[1640]));
    assign outputs[397] = layer0_outputs[727];
    assign outputs[398] = ~((layer0_outputs[1735]) | (layer0_outputs[1268]));
    assign outputs[399] = (layer0_outputs[2068]) & (layer0_outputs[339]);
    assign outputs[400] = ~((layer0_outputs[1641]) | (layer0_outputs[932]));
    assign outputs[401] = ~((layer0_outputs[2261]) ^ (layer0_outputs[1927]));
    assign outputs[402] = ~((layer0_outputs[1833]) | (layer0_outputs[910]));
    assign outputs[403] = layer0_outputs[761];
    assign outputs[404] = (layer0_outputs[795]) & (layer0_outputs[1294]);
    assign outputs[405] = ~(layer0_outputs[194]);
    assign outputs[406] = (layer0_outputs[951]) & (layer0_outputs[759]);
    assign outputs[407] = (layer0_outputs[2457]) & (layer0_outputs[720]);
    assign outputs[408] = ~((layer0_outputs[675]) ^ (layer0_outputs[1241]));
    assign outputs[409] = ~((layer0_outputs[2394]) ^ (layer0_outputs[543]));
    assign outputs[410] = (layer0_outputs[703]) & (layer0_outputs[1106]);
    assign outputs[411] = (layer0_outputs[1143]) & (layer0_outputs[1417]);
    assign outputs[412] = layer0_outputs[1280];
    assign outputs[413] = (layer0_outputs[1974]) & ~(layer0_outputs[405]);
    assign outputs[414] = (layer0_outputs[1545]) & (layer0_outputs[1416]);
    assign outputs[415] = 1'b0;
    assign outputs[416] = layer0_outputs[1895];
    assign outputs[417] = ~((layer0_outputs[1001]) ^ (layer0_outputs[2356]));
    assign outputs[418] = ~((layer0_outputs[1079]) | (layer0_outputs[1062]));
    assign outputs[419] = ~((layer0_outputs[766]) ^ (layer0_outputs[1977]));
    assign outputs[420] = ~(layer0_outputs[2396]);
    assign outputs[421] = layer0_outputs[1960];
    assign outputs[422] = (layer0_outputs[961]) ^ (layer0_outputs[1551]);
    assign outputs[423] = (layer0_outputs[2345]) & ~(layer0_outputs[2484]);
    assign outputs[424] = (layer0_outputs[2371]) & (layer0_outputs[2146]);
    assign outputs[425] = (layer0_outputs[895]) & (layer0_outputs[2317]);
    assign outputs[426] = (layer0_outputs[684]) ^ (layer0_outputs[2180]);
    assign outputs[427] = ~(layer0_outputs[1147]);
    assign outputs[428] = (layer0_outputs[1336]) & (layer0_outputs[1791]);
    assign outputs[429] = (layer0_outputs[103]) ^ (layer0_outputs[1244]);
    assign outputs[430] = (layer0_outputs[2204]) & ~(layer0_outputs[2297]);
    assign outputs[431] = ~((layer0_outputs[1232]) | (layer0_outputs[1082]));
    assign outputs[432] = ~((layer0_outputs[1983]) | (layer0_outputs[192]));
    assign outputs[433] = ~((layer0_outputs[2328]) | (layer0_outputs[342]));
    assign outputs[434] = ~(layer0_outputs[1651]);
    assign outputs[435] = ~((layer0_outputs[372]) ^ (layer0_outputs[304]));
    assign outputs[436] = layer0_outputs[1097];
    assign outputs[437] = ~((layer0_outputs[6]) | (layer0_outputs[1899]));
    assign outputs[438] = (layer0_outputs[493]) & ~(layer0_outputs[2]);
    assign outputs[439] = (layer0_outputs[2115]) & ~(layer0_outputs[394]);
    assign outputs[440] = (layer0_outputs[1145]) & ~(layer0_outputs[1110]);
    assign outputs[441] = ~((layer0_outputs[2340]) | (layer0_outputs[567]));
    assign outputs[442] = (layer0_outputs[1654]) & ~(layer0_outputs[716]);
    assign outputs[443] = ~((layer0_outputs[501]) & (layer0_outputs[2499]));
    assign outputs[444] = ~((layer0_outputs[265]) ^ (layer0_outputs[2099]));
    assign outputs[445] = (layer0_outputs[2273]) & ~(layer0_outputs[1793]);
    assign outputs[446] = (layer0_outputs[701]) & ~(layer0_outputs[2116]);
    assign outputs[447] = (layer0_outputs[745]) & (layer0_outputs[1684]);
    assign outputs[448] = (layer0_outputs[777]) & ~(layer0_outputs[498]);
    assign outputs[449] = (layer0_outputs[1355]) & ~(layer0_outputs[533]);
    assign outputs[450] = (layer0_outputs[2060]) & ~(layer0_outputs[2081]);
    assign outputs[451] = ~((layer0_outputs[138]) | (layer0_outputs[208]));
    assign outputs[452] = (layer0_outputs[1054]) ^ (layer0_outputs[1125]);
    assign outputs[453] = (layer0_outputs[2317]) & (layer0_outputs[2345]);
    assign outputs[454] = (layer0_outputs[2371]) & ~(layer0_outputs[1388]);
    assign outputs[455] = (layer0_outputs[40]) & ~(layer0_outputs[539]);
    assign outputs[456] = (layer0_outputs[172]) & ~(layer0_outputs[2085]);
    assign outputs[457] = (layer0_outputs[748]) & ~(layer0_outputs[1900]);
    assign outputs[458] = (layer0_outputs[2334]) & (layer0_outputs[2410]);
    assign outputs[459] = (layer0_outputs[848]) & ~(layer0_outputs[1781]);
    assign outputs[460] = 1'b0;
    assign outputs[461] = (layer0_outputs[838]) ^ (layer0_outputs[945]);
    assign outputs[462] = (layer0_outputs[1415]) & ~(layer0_outputs[1267]);
    assign outputs[463] = (layer0_outputs[829]) ^ (layer0_outputs[1122]);
    assign outputs[464] = (layer0_outputs[1837]) & (layer0_outputs[1797]);
    assign outputs[465] = (layer0_outputs[421]) & ~(layer0_outputs[1055]);
    assign outputs[466] = (layer0_outputs[497]) ^ (layer0_outputs[2006]);
    assign outputs[467] = ~(layer0_outputs[1923]);
    assign outputs[468] = (layer0_outputs[440]) ^ (layer0_outputs[1704]);
    assign outputs[469] = (layer0_outputs[2274]) & ~(layer0_outputs[2034]);
    assign outputs[470] = layer0_outputs[1726];
    assign outputs[471] = ~((layer0_outputs[2217]) & (layer0_outputs[186]));
    assign outputs[472] = layer0_outputs[246];
    assign outputs[473] = layer0_outputs[1686];
    assign outputs[474] = (layer0_outputs[1665]) & ~(layer0_outputs[410]);
    assign outputs[475] = ~(layer0_outputs[60]);
    assign outputs[476] = (layer0_outputs[56]) & ~(layer0_outputs[605]);
    assign outputs[477] = ~((layer0_outputs[870]) | (layer0_outputs[1279]));
    assign outputs[478] = ~((layer0_outputs[2293]) ^ (layer0_outputs[448]));
    assign outputs[479] = (layer0_outputs[2136]) & ~(layer0_outputs[730]);
    assign outputs[480] = (layer0_outputs[1902]) ^ (layer0_outputs[628]);
    assign outputs[481] = (layer0_outputs[1460]) & ~(layer0_outputs[767]);
    assign outputs[482] = ~((layer0_outputs[255]) | (layer0_outputs[715]));
    assign outputs[483] = (layer0_outputs[1015]) ^ (layer0_outputs[1039]);
    assign outputs[484] = (layer0_outputs[2408]) & (layer0_outputs[946]);
    assign outputs[485] = (layer0_outputs[1922]) & ~(layer0_outputs[979]);
    assign outputs[486] = (layer0_outputs[992]) & ~(layer0_outputs[1610]);
    assign outputs[487] = (layer0_outputs[842]) & ~(layer0_outputs[2398]);
    assign outputs[488] = (layer0_outputs[2236]) & (layer0_outputs[2355]);
    assign outputs[489] = (layer0_outputs[2156]) & (layer0_outputs[590]);
    assign outputs[490] = ~((layer0_outputs[1301]) ^ (layer0_outputs[1984]));
    assign outputs[491] = ~((layer0_outputs[1439]) ^ (layer0_outputs[2271]));
    assign outputs[492] = (layer0_outputs[1561]) & (layer0_outputs[1306]);
    assign outputs[493] = layer0_outputs[2168];
    assign outputs[494] = ~((layer0_outputs[90]) ^ (layer0_outputs[355]));
    assign outputs[495] = ~((layer0_outputs[733]) | (layer0_outputs[2004]));
    assign outputs[496] = (layer0_outputs[429]) & ~(layer0_outputs[808]);
    assign outputs[497] = (layer0_outputs[2372]) & (layer0_outputs[2233]);
    assign outputs[498] = ~((layer0_outputs[2215]) ^ (layer0_outputs[938]));
    assign outputs[499] = (layer0_outputs[345]) & ~(layer0_outputs[1400]);
    assign outputs[500] = (layer0_outputs[1445]) | (layer0_outputs[1724]);
    assign outputs[501] = ~((layer0_outputs[183]) | (layer0_outputs[1762]));
    assign outputs[502] = ~((layer0_outputs[1142]) & (layer0_outputs[8]));
    assign outputs[503] = (layer0_outputs[1284]) ^ (layer0_outputs[1261]);
    assign outputs[504] = layer0_outputs[145];
    assign outputs[505] = ~(layer0_outputs[1323]);
    assign outputs[506] = (layer0_outputs[483]) | (layer0_outputs[2115]);
    assign outputs[507] = layer0_outputs[967];
    assign outputs[508] = (layer0_outputs[697]) & ~(layer0_outputs[2363]);
    assign outputs[509] = ~(layer0_outputs[620]) | (layer0_outputs[1073]);
    assign outputs[510] = (layer0_outputs[96]) | (layer0_outputs[2183]);
    assign outputs[511] = (layer0_outputs[1179]) & ~(layer0_outputs[819]);
    assign outputs[512] = (layer0_outputs[1656]) & (layer0_outputs[1667]);
    assign outputs[513] = layer0_outputs[514];
    assign outputs[514] = ~(layer0_outputs[1440]);
    assign outputs[515] = (layer0_outputs[1496]) & (layer0_outputs[480]);
    assign outputs[516] = ~((layer0_outputs[1337]) & (layer0_outputs[1102]));
    assign outputs[517] = layer0_outputs[242];
    assign outputs[518] = ~(layer0_outputs[521]);
    assign outputs[519] = ~((layer0_outputs[330]) | (layer0_outputs[2318]));
    assign outputs[520] = ~(layer0_outputs[1404]);
    assign outputs[521] = layer0_outputs[1214];
    assign outputs[522] = ~((layer0_outputs[110]) & (layer0_outputs[1116]));
    assign outputs[523] = ~(layer0_outputs[2246]) | (layer0_outputs[376]);
    assign outputs[524] = ~(layer0_outputs[1194]) | (layer0_outputs[2254]);
    assign outputs[525] = layer0_outputs[1113];
    assign outputs[526] = (layer0_outputs[2443]) & ~(layer0_outputs[1777]);
    assign outputs[527] = layer0_outputs[1454];
    assign outputs[528] = (layer0_outputs[943]) & ~(layer0_outputs[348]);
    assign outputs[529] = ~(layer0_outputs[357]);
    assign outputs[530] = (layer0_outputs[1900]) & (layer0_outputs[1858]);
    assign outputs[531] = ~((layer0_outputs[470]) ^ (layer0_outputs[1481]));
    assign outputs[532] = ~((layer0_outputs[1409]) | (layer0_outputs[1666]));
    assign outputs[533] = ~(layer0_outputs[1158]) | (layer0_outputs[262]);
    assign outputs[534] = ~((layer0_outputs[184]) ^ (layer0_outputs[806]));
    assign outputs[535] = ~(layer0_outputs[1209]) | (layer0_outputs[1509]);
    assign outputs[536] = ~((layer0_outputs[614]) | (layer0_outputs[1582]));
    assign outputs[537] = layer0_outputs[1365];
    assign outputs[538] = ~((layer0_outputs[1208]) | (layer0_outputs[350]));
    assign outputs[539] = ~(layer0_outputs[2244]);
    assign outputs[540] = ~(layer0_outputs[53]) | (layer0_outputs[980]);
    assign outputs[541] = (layer0_outputs[973]) | (layer0_outputs[1188]);
    assign outputs[542] = (layer0_outputs[457]) ^ (layer0_outputs[532]);
    assign outputs[543] = ~((layer0_outputs[1870]) & (layer0_outputs[1428]));
    assign outputs[544] = ~((layer0_outputs[2175]) ^ (layer0_outputs[1876]));
    assign outputs[545] = layer0_outputs[1274];
    assign outputs[546] = (layer0_outputs[483]) & ~(layer0_outputs[795]);
    assign outputs[547] = ~(layer0_outputs[1649]);
    assign outputs[548] = ~((layer0_outputs[864]) | (layer0_outputs[197]));
    assign outputs[549] = ~(layer0_outputs[1209]);
    assign outputs[550] = (layer0_outputs[80]) & ~(layer0_outputs[2309]);
    assign outputs[551] = ~(layer0_outputs[2389]) | (layer0_outputs[2178]);
    assign outputs[552] = ~((layer0_outputs[758]) & (layer0_outputs[1131]));
    assign outputs[553] = (layer0_outputs[2092]) & (layer0_outputs[2466]);
    assign outputs[554] = ~((layer0_outputs[408]) ^ (layer0_outputs[1915]));
    assign outputs[555] = layer0_outputs[2400];
    assign outputs[556] = ~(layer0_outputs[2230]);
    assign outputs[557] = ~((layer0_outputs[347]) ^ (layer0_outputs[2019]));
    assign outputs[558] = layer0_outputs[1664];
    assign outputs[559] = layer0_outputs[1600];
    assign outputs[560] = (layer0_outputs[641]) & (layer0_outputs[991]);
    assign outputs[561] = ~((layer0_outputs[52]) ^ (layer0_outputs[744]));
    assign outputs[562] = ~(layer0_outputs[400]);
    assign outputs[563] = ~((layer0_outputs[547]) ^ (layer0_outputs[1386]));
    assign outputs[564] = ~(layer0_outputs[725]) | (layer0_outputs[1122]);
    assign outputs[565] = layer0_outputs[807];
    assign outputs[566] = ~(layer0_outputs[1408]) | (layer0_outputs[1557]);
    assign outputs[567] = ~(layer0_outputs[755]);
    assign outputs[568] = ~((layer0_outputs[2204]) | (layer0_outputs[885]));
    assign outputs[569] = (layer0_outputs[81]) & ~(layer0_outputs[2260]);
    assign outputs[570] = ~(layer0_outputs[1798]) | (layer0_outputs[1346]);
    assign outputs[571] = (layer0_outputs[207]) & ~(layer0_outputs[503]);
    assign outputs[572] = ~((layer0_outputs[274]) | (layer0_outputs[1861]));
    assign outputs[573] = ~(layer0_outputs[364]) | (layer0_outputs[421]);
    assign outputs[574] = ~(layer0_outputs[788]);
    assign outputs[575] = (layer0_outputs[2128]) & (layer0_outputs[1108]);
    assign outputs[576] = layer0_outputs[1858];
    assign outputs[577] = ~(layer0_outputs[1874]);
    assign outputs[578] = layer0_outputs[538];
    assign outputs[579] = ~(layer0_outputs[2012]) | (layer0_outputs[699]);
    assign outputs[580] = ~(layer0_outputs[742]) | (layer0_outputs[856]);
    assign outputs[581] = (layer0_outputs[401]) ^ (layer0_outputs[268]);
    assign outputs[582] = layer0_outputs[1353];
    assign outputs[583] = ~(layer0_outputs[129]);
    assign outputs[584] = layer0_outputs[352];
    assign outputs[585] = ~(layer0_outputs[1660]);
    assign outputs[586] = layer0_outputs[1517];
    assign outputs[587] = ~(layer0_outputs[2491]) | (layer0_outputs[569]);
    assign outputs[588] = (layer0_outputs[1133]) | (layer0_outputs[799]);
    assign outputs[589] = ~((layer0_outputs[189]) & (layer0_outputs[2333]));
    assign outputs[590] = ~(layer0_outputs[2182]) | (layer0_outputs[382]);
    assign outputs[591] = layer0_outputs[746];
    assign outputs[592] = (layer0_outputs[743]) ^ (layer0_outputs[2152]);
    assign outputs[593] = (layer0_outputs[239]) & (layer0_outputs[485]);
    assign outputs[594] = ~(layer0_outputs[2385]);
    assign outputs[595] = layer0_outputs[148];
    assign outputs[596] = ~(layer0_outputs[2366]) | (layer0_outputs[130]);
    assign outputs[597] = (layer0_outputs[1633]) & ~(layer0_outputs[1066]);
    assign outputs[598] = (layer0_outputs[244]) & ~(layer0_outputs[1989]);
    assign outputs[599] = layer0_outputs[423];
    assign outputs[600] = ~(layer0_outputs[1265]) | (layer0_outputs[449]);
    assign outputs[601] = layer0_outputs[1126];
    assign outputs[602] = (layer0_outputs[337]) | (layer0_outputs[1191]);
    assign outputs[603] = ~(layer0_outputs[1109]) | (layer0_outputs[16]);
    assign outputs[604] = ~(layer0_outputs[1344]) | (layer0_outputs[2486]);
    assign outputs[605] = (layer0_outputs[2277]) & ~(layer0_outputs[1240]);
    assign outputs[606] = (layer0_outputs[670]) & (layer0_outputs[2413]);
    assign outputs[607] = (layer0_outputs[2006]) ^ (layer0_outputs[1672]);
    assign outputs[608] = layer0_outputs[2241];
    assign outputs[609] = ~(layer0_outputs[619]) | (layer0_outputs[1197]);
    assign outputs[610] = ~(layer0_outputs[51]);
    assign outputs[611] = ~((layer0_outputs[846]) ^ (layer0_outputs[1202]));
    assign outputs[612] = ~((layer0_outputs[654]) | (layer0_outputs[1629]));
    assign outputs[613] = (layer0_outputs[1537]) | (layer0_outputs[181]);
    assign outputs[614] = ~((layer0_outputs[496]) ^ (layer0_outputs[2063]));
    assign outputs[615] = ~(layer0_outputs[778]) | (layer0_outputs[1783]);
    assign outputs[616] = layer0_outputs[1950];
    assign outputs[617] = ~(layer0_outputs[1139]) | (layer0_outputs[1467]);
    assign outputs[618] = ~(layer0_outputs[316]) | (layer0_outputs[232]);
    assign outputs[619] = ~(layer0_outputs[653]);
    assign outputs[620] = (layer0_outputs[403]) & ~(layer0_outputs[2359]);
    assign outputs[621] = layer0_outputs[432];
    assign outputs[622] = ~(layer0_outputs[2220]) | (layer0_outputs[822]);
    assign outputs[623] = ~(layer0_outputs[1518]) | (layer0_outputs[979]);
    assign outputs[624] = layer0_outputs[68];
    assign outputs[625] = layer0_outputs[1591];
    assign outputs[626] = (layer0_outputs[1844]) ^ (layer0_outputs[2336]);
    assign outputs[627] = (layer0_outputs[191]) ^ (layer0_outputs[148]);
    assign outputs[628] = ~(layer0_outputs[1015]) | (layer0_outputs[273]);
    assign outputs[629] = layer0_outputs[2148];
    assign outputs[630] = layer0_outputs[452];
    assign outputs[631] = ~(layer0_outputs[1221]) | (layer0_outputs[1880]);
    assign outputs[632] = layer0_outputs[954];
    assign outputs[633] = (layer0_outputs[1824]) & ~(layer0_outputs[503]);
    assign outputs[634] = (layer0_outputs[240]) & ~(layer0_outputs[563]);
    assign outputs[635] = layer0_outputs[2089];
    assign outputs[636] = (layer0_outputs[1300]) ^ (layer0_outputs[1789]);
    assign outputs[637] = ~(layer0_outputs[1440]) | (layer0_outputs[2316]);
    assign outputs[638] = ~((layer0_outputs[1946]) | (layer0_outputs[1572]));
    assign outputs[639] = layer0_outputs[1990];
    assign outputs[640] = ~(layer0_outputs[1628]) | (layer0_outputs[781]);
    assign outputs[641] = ~(layer0_outputs[2460]) | (layer0_outputs[388]);
    assign outputs[642] = (layer0_outputs[1908]) ^ (layer0_outputs[1338]);
    assign outputs[643] = layer0_outputs[409];
    assign outputs[644] = ~(layer0_outputs[864]);
    assign outputs[645] = (layer0_outputs[1652]) & ~(layer0_outputs[1568]);
    assign outputs[646] = ~((layer0_outputs[2285]) ^ (layer0_outputs[80]));
    assign outputs[647] = layer0_outputs[245];
    assign outputs[648] = layer0_outputs[1215];
    assign outputs[649] = ~(layer0_outputs[576]) | (layer0_outputs[943]);
    assign outputs[650] = ~(layer0_outputs[625]);
    assign outputs[651] = layer0_outputs[2082];
    assign outputs[652] = layer0_outputs[1038];
    assign outputs[653] = ~((layer0_outputs[1658]) ^ (layer0_outputs[611]));
    assign outputs[654] = (layer0_outputs[775]) & ~(layer0_outputs[316]);
    assign outputs[655] = ~(layer0_outputs[271]) | (layer0_outputs[669]);
    assign outputs[656] = ~(layer0_outputs[840]) | (layer0_outputs[1822]);
    assign outputs[657] = (layer0_outputs[2324]) ^ (layer0_outputs[2083]);
    assign outputs[658] = ~((layer0_outputs[404]) | (layer0_outputs[450]));
    assign outputs[659] = (layer0_outputs[30]) & ~(layer0_outputs[2298]);
    assign outputs[660] = ~(layer0_outputs[1135]);
    assign outputs[661] = ~((layer0_outputs[778]) & (layer0_outputs[2360]));
    assign outputs[662] = (layer0_outputs[685]) & (layer0_outputs[852]);
    assign outputs[663] = layer0_outputs[2464];
    assign outputs[664] = ~(layer0_outputs[500]);
    assign outputs[665] = layer0_outputs[1450];
    assign outputs[666] = (layer0_outputs[912]) | (layer0_outputs[1421]);
    assign outputs[667] = layer0_outputs[2176];
    assign outputs[668] = (layer0_outputs[213]) & (layer0_outputs[1871]);
    assign outputs[669] = (layer0_outputs[203]) & ~(layer0_outputs[1302]);
    assign outputs[670] = layer0_outputs[1748];
    assign outputs[671] = ~(layer0_outputs[398]) | (layer0_outputs[900]);
    assign outputs[672] = ~(layer0_outputs[469]);
    assign outputs[673] = layer0_outputs[1838];
    assign outputs[674] = (layer0_outputs[1067]) & ~(layer0_outputs[74]);
    assign outputs[675] = ~(layer0_outputs[437]);
    assign outputs[676] = ~((layer0_outputs[579]) ^ (layer0_outputs[790]));
    assign outputs[677] = ~(layer0_outputs[1988]) | (layer0_outputs[2114]);
    assign outputs[678] = ~(layer0_outputs[2444]);
    assign outputs[679] = (layer0_outputs[9]) & ~(layer0_outputs[531]);
    assign outputs[680] = (layer0_outputs[1935]) & ~(layer0_outputs[2389]);
    assign outputs[681] = layer0_outputs[1354];
    assign outputs[682] = ~(layer0_outputs[1966]);
    assign outputs[683] = (layer0_outputs[1429]) & ~(layer0_outputs[1459]);
    assign outputs[684] = (layer0_outputs[1466]) | (layer0_outputs[587]);
    assign outputs[685] = ~(layer0_outputs[1057]) | (layer0_outputs[1179]);
    assign outputs[686] = ~(layer0_outputs[2219]);
    assign outputs[687] = ~(layer0_outputs[548]);
    assign outputs[688] = (layer0_outputs[1173]) ^ (layer0_outputs[1162]);
    assign outputs[689] = layer0_outputs[833];
    assign outputs[690] = (layer0_outputs[1972]) | (layer0_outputs[1781]);
    assign outputs[691] = (layer0_outputs[152]) & ~(layer0_outputs[1618]);
    assign outputs[692] = (layer0_outputs[1687]) & ~(layer0_outputs[1946]);
    assign outputs[693] = ~(layer0_outputs[324]) | (layer0_outputs[747]);
    assign outputs[694] = ~(layer0_outputs[1023]);
    assign outputs[695] = ~(layer0_outputs[1091]);
    assign outputs[696] = (layer0_outputs[915]) & (layer0_outputs[1632]);
    assign outputs[697] = ~((layer0_outputs[2177]) | (layer0_outputs[1764]));
    assign outputs[698] = ~((layer0_outputs[1038]) ^ (layer0_outputs[1687]));
    assign outputs[699] = ~(layer0_outputs[1945]);
    assign outputs[700] = (layer0_outputs[2084]) & ~(layer0_outputs[2053]);
    assign outputs[701] = ~(layer0_outputs[2499]);
    assign outputs[702] = layer0_outputs[11];
    assign outputs[703] = ~(layer0_outputs[2372]) | (layer0_outputs[1039]);
    assign outputs[704] = layer0_outputs[1831];
    assign outputs[705] = ~((layer0_outputs[516]) ^ (layer0_outputs[1072]));
    assign outputs[706] = (layer0_outputs[2423]) & ~(layer0_outputs[89]);
    assign outputs[707] = ~(layer0_outputs[2275]) | (layer0_outputs[1437]);
    assign outputs[708] = ~(layer0_outputs[51]);
    assign outputs[709] = (layer0_outputs[2284]) & (layer0_outputs[413]);
    assign outputs[710] = (layer0_outputs[2023]) ^ (layer0_outputs[876]);
    assign outputs[711] = (layer0_outputs[1684]) | (layer0_outputs[1402]);
    assign outputs[712] = layer0_outputs[1205];
    assign outputs[713] = (layer0_outputs[1378]) ^ (layer0_outputs[188]);
    assign outputs[714] = (layer0_outputs[1205]) & ~(layer0_outputs[22]);
    assign outputs[715] = layer0_outputs[287];
    assign outputs[716] = layer0_outputs[2228];
    assign outputs[717] = layer0_outputs[547];
    assign outputs[718] = ~(layer0_outputs[549]) | (layer0_outputs[2319]);
    assign outputs[719] = ~((layer0_outputs[427]) & (layer0_outputs[1627]));
    assign outputs[720] = ~(layer0_outputs[1332]) | (layer0_outputs[2098]);
    assign outputs[721] = layer0_outputs[2030];
    assign outputs[722] = ~((layer0_outputs[2452]) | (layer0_outputs[983]));
    assign outputs[723] = layer0_outputs[1728];
    assign outputs[724] = ~(layer0_outputs[166]) | (layer0_outputs[1812]);
    assign outputs[725] = ~(layer0_outputs[1702]);
    assign outputs[726] = (layer0_outputs[777]) & (layer0_outputs[244]);
    assign outputs[727] = layer0_outputs[226];
    assign outputs[728] = ~(layer0_outputs[657]);
    assign outputs[729] = (layer0_outputs[1553]) | (layer0_outputs[1595]);
    assign outputs[730] = layer0_outputs[1579];
    assign outputs[731] = layer0_outputs[158];
    assign outputs[732] = ~((layer0_outputs[1680]) ^ (layer0_outputs[1570]));
    assign outputs[733] = ~(layer0_outputs[2353]);
    assign outputs[734] = ~(layer0_outputs[462]) | (layer0_outputs[1825]);
    assign outputs[735] = (layer0_outputs[610]) ^ (layer0_outputs[108]);
    assign outputs[736] = ~(layer0_outputs[1154]);
    assign outputs[737] = layer0_outputs[1243];
    assign outputs[738] = ~((layer0_outputs[584]) & (layer0_outputs[1797]));
    assign outputs[739] = layer0_outputs[1011];
    assign outputs[740] = ~(layer0_outputs[247]);
    assign outputs[741] = (layer0_outputs[1168]) ^ (layer0_outputs[815]);
    assign outputs[742] = layer0_outputs[2086];
    assign outputs[743] = (layer0_outputs[2262]) & ~(layer0_outputs[881]);
    assign outputs[744] = ~(layer0_outputs[875]);
    assign outputs[745] = (layer0_outputs[1422]) & (layer0_outputs[833]);
    assign outputs[746] = ~((layer0_outputs[648]) & (layer0_outputs[436]));
    assign outputs[747] = (layer0_outputs[1742]) & (layer0_outputs[170]);
    assign outputs[748] = ~(layer0_outputs[913]) | (layer0_outputs[1320]);
    assign outputs[749] = ~(layer0_outputs[1569]) | (layer0_outputs[367]);
    assign outputs[750] = ~(layer0_outputs[1721]) | (layer0_outputs[2225]);
    assign outputs[751] = (layer0_outputs[1688]) & ~(layer0_outputs[436]);
    assign outputs[752] = ~(layer0_outputs[1957]);
    assign outputs[753] = (layer0_outputs[2054]) & ~(layer0_outputs[1390]);
    assign outputs[754] = ~((layer0_outputs[1172]) | (layer0_outputs[1814]));
    assign outputs[755] = ~((layer0_outputs[1168]) | (layer0_outputs[1234]));
    assign outputs[756] = ~((layer0_outputs[2260]) | (layer0_outputs[1672]));
    assign outputs[757] = (layer0_outputs[1802]) & ~(layer0_outputs[2057]);
    assign outputs[758] = (layer0_outputs[2079]) & (layer0_outputs[193]);
    assign outputs[759] = ~((layer0_outputs[1412]) | (layer0_outputs[1508]));
    assign outputs[760] = ~(layer0_outputs[2361]);
    assign outputs[761] = (layer0_outputs[739]) & ~(layer0_outputs[1660]);
    assign outputs[762] = layer0_outputs[208];
    assign outputs[763] = (layer0_outputs[1555]) & ~(layer0_outputs[1725]);
    assign outputs[764] = ~((layer0_outputs[18]) & (layer0_outputs[323]));
    assign outputs[765] = (layer0_outputs[1232]) & (layer0_outputs[2067]);
    assign outputs[766] = (layer0_outputs[321]) & ~(layer0_outputs[1530]);
    assign outputs[767] = (layer0_outputs[680]) & (layer0_outputs[1696]);
    assign outputs[768] = (layer0_outputs[499]) & (layer0_outputs[804]);
    assign outputs[769] = (layer0_outputs[1341]) | (layer0_outputs[367]);
    assign outputs[770] = (layer0_outputs[713]) & ~(layer0_outputs[1263]);
    assign outputs[771] = layer0_outputs[229];
    assign outputs[772] = (layer0_outputs[1611]) & ~(layer0_outputs[1369]);
    assign outputs[773] = (layer0_outputs[693]) & ~(layer0_outputs[2240]);
    assign outputs[774] = (layer0_outputs[1569]) & ~(layer0_outputs[232]);
    assign outputs[775] = ~(layer0_outputs[1138]);
    assign outputs[776] = ~(layer0_outputs[806]) | (layer0_outputs[594]);
    assign outputs[777] = (layer0_outputs[37]) ^ (layer0_outputs[1904]);
    assign outputs[778] = layer0_outputs[1287];
    assign outputs[779] = (layer0_outputs[2449]) & (layer0_outputs[181]);
    assign outputs[780] = (layer0_outputs[1832]) & ~(layer0_outputs[47]);
    assign outputs[781] = ~(layer0_outputs[760]);
    assign outputs[782] = (layer0_outputs[2379]) | (layer0_outputs[639]);
    assign outputs[783] = (layer0_outputs[696]) ^ (layer0_outputs[1163]);
    assign outputs[784] = ~(layer0_outputs[1805]);
    assign outputs[785] = (layer0_outputs[1394]) & ~(layer0_outputs[1362]);
    assign outputs[786] = ~(layer0_outputs[1817]) | (layer0_outputs[362]);
    assign outputs[787] = layer0_outputs[1350];
    assign outputs[788] = ~(layer0_outputs[667]);
    assign outputs[789] = layer0_outputs[1002];
    assign outputs[790] = (layer0_outputs[721]) & (layer0_outputs[2448]);
    assign outputs[791] = layer0_outputs[117];
    assign outputs[792] = ~((layer0_outputs[964]) | (layer0_outputs[1075]));
    assign outputs[793] = (layer0_outputs[1947]) & (layer0_outputs[590]);
    assign outputs[794] = ~((layer0_outputs[1558]) | (layer0_outputs[1969]));
    assign outputs[795] = (layer0_outputs[526]) ^ (layer0_outputs[1215]);
    assign outputs[796] = layer0_outputs[2151];
    assign outputs[797] = (layer0_outputs[891]) & ~(layer0_outputs[738]);
    assign outputs[798] = layer0_outputs[609];
    assign outputs[799] = (layer0_outputs[809]) & ~(layer0_outputs[1773]);
    assign outputs[800] = ~(layer0_outputs[1081]) | (layer0_outputs[1596]);
    assign outputs[801] = (layer0_outputs[333]) & ~(layer0_outputs[1668]);
    assign outputs[802] = layer0_outputs[679];
    assign outputs[803] = layer0_outputs[1203];
    assign outputs[804] = ~((layer0_outputs[2321]) ^ (layer0_outputs[1746]));
    assign outputs[805] = (layer0_outputs[1265]) ^ (layer0_outputs[618]);
    assign outputs[806] = ~((layer0_outputs[282]) | (layer0_outputs[633]));
    assign outputs[807] = ~((layer0_outputs[1483]) & (layer0_outputs[1165]));
    assign outputs[808] = (layer0_outputs[1981]) | (layer0_outputs[1789]);
    assign outputs[809] = ~((layer0_outputs[1253]) ^ (layer0_outputs[862]));
    assign outputs[810] = ~(layer0_outputs[595]);
    assign outputs[811] = ~(layer0_outputs[560]);
    assign outputs[812] = (layer0_outputs[2100]) & ~(layer0_outputs[1749]);
    assign outputs[813] = ~((layer0_outputs[1918]) ^ (layer0_outputs[2476]));
    assign outputs[814] = (layer0_outputs[881]) | (layer0_outputs[106]);
    assign outputs[815] = ~(layer0_outputs[1076]) | (layer0_outputs[1628]);
    assign outputs[816] = ~(layer0_outputs[1901]);
    assign outputs[817] = ~(layer0_outputs[1171]);
    assign outputs[818] = (layer0_outputs[1186]) & ~(layer0_outputs[1431]);
    assign outputs[819] = layer0_outputs[1430];
    assign outputs[820] = ~(layer0_outputs[1725]);
    assign outputs[821] = ~(layer0_outputs[930]);
    assign outputs[822] = ~((layer0_outputs[1025]) ^ (layer0_outputs[969]));
    assign outputs[823] = layer0_outputs[1072];
    assign outputs[824] = (layer0_outputs[2386]) & ~(layer0_outputs[86]);
    assign outputs[825] = (layer0_outputs[118]) & ~(layer0_outputs[93]);
    assign outputs[826] = ~(layer0_outputs[142]);
    assign outputs[827] = ~((layer0_outputs[1016]) & (layer0_outputs[1535]));
    assign outputs[828] = layer0_outputs[1930];
    assign outputs[829] = (layer0_outputs[955]) & ~(layer0_outputs[802]);
    assign outputs[830] = layer0_outputs[224];
    assign outputs[831] = ~((layer0_outputs[631]) ^ (layer0_outputs[1940]));
    assign outputs[832] = (layer0_outputs[1555]) & ~(layer0_outputs[1525]);
    assign outputs[833] = (layer0_outputs[1982]) & ~(layer0_outputs[408]);
    assign outputs[834] = (layer0_outputs[974]) & ~(layer0_outputs[1800]);
    assign outputs[835] = (layer0_outputs[1404]) & ~(layer0_outputs[964]);
    assign outputs[836] = layer0_outputs[2151];
    assign outputs[837] = ~((layer0_outputs[827]) ^ (layer0_outputs[977]));
    assign outputs[838] = (layer0_outputs[689]) ^ (layer0_outputs[2216]);
    assign outputs[839] = ~(layer0_outputs[536]);
    assign outputs[840] = layer0_outputs[739];
    assign outputs[841] = ~(layer0_outputs[812]);
    assign outputs[842] = ~((layer0_outputs[534]) | (layer0_outputs[206]));
    assign outputs[843] = ~(layer0_outputs[161]);
    assign outputs[844] = (layer0_outputs[1248]) & ~(layer0_outputs[256]);
    assign outputs[845] = layer0_outputs[1562];
    assign outputs[846] = (layer0_outputs[604]) & ~(layer0_outputs[2273]);
    assign outputs[847] = (layer0_outputs[1574]) & ~(layer0_outputs[1393]);
    assign outputs[848] = ~(layer0_outputs[142]) | (layer0_outputs[1022]);
    assign outputs[849] = layer0_outputs[1939];
    assign outputs[850] = ~((layer0_outputs[2278]) & (layer0_outputs[606]));
    assign outputs[851] = ~((layer0_outputs[341]) ^ (layer0_outputs[1446]));
    assign outputs[852] = (layer0_outputs[2033]) & (layer0_outputs[1156]);
    assign outputs[853] = (layer0_outputs[1394]) & ~(layer0_outputs[1436]);
    assign outputs[854] = ~(layer0_outputs[1722]);
    assign outputs[855] = ~(layer0_outputs[1632]);
    assign outputs[856] = (layer0_outputs[1361]) & ~(layer0_outputs[1675]);
    assign outputs[857] = (layer0_outputs[2348]) | (layer0_outputs[2375]);
    assign outputs[858] = (layer0_outputs[2373]) & ~(layer0_outputs[1185]);
    assign outputs[859] = (layer0_outputs[2239]) & ~(layer0_outputs[2451]);
    assign outputs[860] = ~(layer0_outputs[2487]) | (layer0_outputs[1118]);
    assign outputs[861] = ~(layer0_outputs[1753]);
    assign outputs[862] = ~(layer0_outputs[682]) | (layer0_outputs[2409]);
    assign outputs[863] = (layer0_outputs[2402]) & ~(layer0_outputs[691]);
    assign outputs[864] = ~(layer0_outputs[1888]);
    assign outputs[865] = ~(layer0_outputs[2422]);
    assign outputs[866] = (layer0_outputs[1770]) & ~(layer0_outputs[67]);
    assign outputs[867] = layer0_outputs[15];
    assign outputs[868] = (layer0_outputs[976]) ^ (layer0_outputs[1570]);
    assign outputs[869] = ~(layer0_outputs[523]);
    assign outputs[870] = layer0_outputs[854];
    assign outputs[871] = ~(layer0_outputs[1794]) | (layer0_outputs[171]);
    assign outputs[872] = layer0_outputs[453];
    assign outputs[873] = ~((layer0_outputs[1178]) ^ (layer0_outputs[708]));
    assign outputs[874] = ~((layer0_outputs[1104]) & (layer0_outputs[1494]));
    assign outputs[875] = ~(layer0_outputs[1091]) | (layer0_outputs[1958]);
    assign outputs[876] = layer0_outputs[239];
    assign outputs[877] = (layer0_outputs[574]) & ~(layer0_outputs[1424]);
    assign outputs[878] = ~(layer0_outputs[2187]);
    assign outputs[879] = layer0_outputs[2300];
    assign outputs[880] = ~((layer0_outputs[2395]) ^ (layer0_outputs[2061]));
    assign outputs[881] = (layer0_outputs[2190]) & ~(layer0_outputs[957]);
    assign outputs[882] = ~((layer0_outputs[259]) ^ (layer0_outputs[117]));
    assign outputs[883] = (layer0_outputs[1282]) ^ (layer0_outputs[981]);
    assign outputs[884] = (layer0_outputs[661]) & ~(layer0_outputs[2110]);
    assign outputs[885] = ~((layer0_outputs[2444]) | (layer0_outputs[1838]));
    assign outputs[886] = layer0_outputs[301];
    assign outputs[887] = layer0_outputs[64];
    assign outputs[888] = layer0_outputs[2264];
    assign outputs[889] = ~((layer0_outputs[1872]) & (layer0_outputs[1702]));
    assign outputs[890] = ~(layer0_outputs[1489]);
    assign outputs[891] = ~(layer0_outputs[2050]) | (layer0_outputs[1669]);
    assign outputs[892] = ~(layer0_outputs[276]);
    assign outputs[893] = ~((layer0_outputs[722]) | (layer0_outputs[20]));
    assign outputs[894] = ~((layer0_outputs[2164]) | (layer0_outputs[861]));
    assign outputs[895] = (layer0_outputs[2246]) ^ (layer0_outputs[1701]);
    assign outputs[896] = ~(layer0_outputs[1952]);
    assign outputs[897] = (layer0_outputs[2130]) ^ (layer0_outputs[1010]);
    assign outputs[898] = ~(layer0_outputs[119]);
    assign outputs[899] = layer0_outputs[945];
    assign outputs[900] = ~(layer0_outputs[1619]);
    assign outputs[901] = layer0_outputs[164];
    assign outputs[902] = (layer0_outputs[1020]) ^ (layer0_outputs[371]);
    assign outputs[903] = (layer0_outputs[1571]) & (layer0_outputs[1582]);
    assign outputs[904] = ~(layer0_outputs[340]);
    assign outputs[905] = ~((layer0_outputs[1629]) ^ (layer0_outputs[157]));
    assign outputs[906] = ~((layer0_outputs[1379]) ^ (layer0_outputs[2008]));
    assign outputs[907] = layer0_outputs[1960];
    assign outputs[908] = ~((layer0_outputs[1587]) ^ (layer0_outputs[454]));
    assign outputs[909] = (layer0_outputs[133]) & ~(layer0_outputs[501]);
    assign outputs[910] = (layer0_outputs[2376]) & ~(layer0_outputs[1757]);
    assign outputs[911] = (layer0_outputs[2270]) & ~(layer0_outputs[1747]);
    assign outputs[912] = ~((layer0_outputs[147]) ^ (layer0_outputs[508]));
    assign outputs[913] = ~(layer0_outputs[2355]);
    assign outputs[914] = layer0_outputs[2286];
    assign outputs[915] = ~(layer0_outputs[1360]);
    assign outputs[916] = ~(layer0_outputs[1236]) | (layer0_outputs[477]);
    assign outputs[917] = layer0_outputs[6];
    assign outputs[918] = ~(layer0_outputs[736]);
    assign outputs[919] = ~((layer0_outputs[2045]) ^ (layer0_outputs[1608]));
    assign outputs[920] = ~(layer0_outputs[62]) | (layer0_outputs[2033]);
    assign outputs[921] = (layer0_outputs[2091]) & ~(layer0_outputs[1348]);
    assign outputs[922] = (layer0_outputs[1497]) | (layer0_outputs[487]);
    assign outputs[923] = ~(layer0_outputs[377]) | (layer0_outputs[871]);
    assign outputs[924] = (layer0_outputs[2495]) & ~(layer0_outputs[2252]);
    assign outputs[925] = (layer0_outputs[1670]) & (layer0_outputs[1908]);
    assign outputs[926] = ~((layer0_outputs[810]) ^ (layer0_outputs[12]));
    assign outputs[927] = (layer0_outputs[2359]) & ~(layer0_outputs[282]);
    assign outputs[928] = layer0_outputs[1190];
    assign outputs[929] = (layer0_outputs[2177]) & ~(layer0_outputs[221]);
    assign outputs[930] = (layer0_outputs[2393]) & ~(layer0_outputs[2325]);
    assign outputs[931] = layer0_outputs[1257];
    assign outputs[932] = ~((layer0_outputs[1101]) | (layer0_outputs[1677]));
    assign outputs[933] = ~((layer0_outputs[1169]) ^ (layer0_outputs[1755]));
    assign outputs[934] = layer0_outputs[422];
    assign outputs[935] = ~((layer0_outputs[1606]) ^ (layer0_outputs[1536]));
    assign outputs[936] = (layer0_outputs[1317]) & ~(layer0_outputs[1618]);
    assign outputs[937] = layer0_outputs[699];
    assign outputs[938] = (layer0_outputs[1328]) & ~(layer0_outputs[1134]);
    assign outputs[939] = (layer0_outputs[2092]) & (layer0_outputs[1346]);
    assign outputs[940] = ~(layer0_outputs[1086]) | (layer0_outputs[2255]);
    assign outputs[941] = ~(layer0_outputs[2453]) | (layer0_outputs[393]);
    assign outputs[942] = ~((layer0_outputs[2480]) | (layer0_outputs[858]));
    assign outputs[943] = ~((layer0_outputs[2407]) | (layer0_outputs[178]));
    assign outputs[944] = layer0_outputs[155];
    assign outputs[945] = layer0_outputs[1041];
    assign outputs[946] = layer0_outputs[1189];
    assign outputs[947] = ~((layer0_outputs[2476]) ^ (layer0_outputs[1626]));
    assign outputs[948] = ~(layer0_outputs[1482]);
    assign outputs[949] = ~(layer0_outputs[1968]);
    assign outputs[950] = ~(layer0_outputs[1814]);
    assign outputs[951] = (layer0_outputs[561]) & ~(layer0_outputs[522]);
    assign outputs[952] = layer0_outputs[1875];
    assign outputs[953] = ~(layer0_outputs[933]) | (layer0_outputs[1345]);
    assign outputs[954] = ~((layer0_outputs[1739]) | (layer0_outputs[335]));
    assign outputs[955] = layer0_outputs[1818];
    assign outputs[956] = ~((layer0_outputs[1312]) ^ (layer0_outputs[1963]));
    assign outputs[957] = ~(layer0_outputs[206]);
    assign outputs[958] = ~(layer0_outputs[201]);
    assign outputs[959] = (layer0_outputs[936]) | (layer0_outputs[824]);
    assign outputs[960] = layer0_outputs[554];
    assign outputs[961] = (layer0_outputs[989]) | (layer0_outputs[443]);
    assign outputs[962] = layer0_outputs[1013];
    assign outputs[963] = (layer0_outputs[1099]) & (layer0_outputs[111]);
    assign outputs[964] = ~((layer0_outputs[332]) & (layer0_outputs[603]));
    assign outputs[965] = (layer0_outputs[374]) ^ (layer0_outputs[2432]);
    assign outputs[966] = (layer0_outputs[582]) | (layer0_outputs[1150]);
    assign outputs[967] = layer0_outputs[1614];
    assign outputs[968] = (layer0_outputs[2125]) & (layer0_outputs[502]);
    assign outputs[969] = ~(layer0_outputs[828]);
    assign outputs[970] = ~((layer0_outputs[161]) | (layer0_outputs[1772]));
    assign outputs[971] = (layer0_outputs[922]) & (layer0_outputs[430]);
    assign outputs[972] = ~((layer0_outputs[1044]) | (layer0_outputs[2340]));
    assign outputs[973] = (layer0_outputs[147]) ^ (layer0_outputs[2439]);
    assign outputs[974] = (layer0_outputs[842]) & ~(layer0_outputs[281]);
    assign outputs[975] = (layer0_outputs[1144]) ^ (layer0_outputs[124]);
    assign outputs[976] = ~((layer0_outputs[511]) | (layer0_outputs[1519]));
    assign outputs[977] = ~(layer0_outputs[1953]);
    assign outputs[978] = (layer0_outputs[1933]) ^ (layer0_outputs[1709]);
    assign outputs[979] = (layer0_outputs[1839]) & (layer0_outputs[428]);
    assign outputs[980] = ~((layer0_outputs[496]) | (layer0_outputs[310]));
    assign outputs[981] = (layer0_outputs[172]) & (layer0_outputs[645]);
    assign outputs[982] = ~(layer0_outputs[2430]) | (layer0_outputs[114]);
    assign outputs[983] = (layer0_outputs[663]) ^ (layer0_outputs[1083]);
    assign outputs[984] = (layer0_outputs[1647]) & (layer0_outputs[1962]);
    assign outputs[985] = layer0_outputs[2048];
    assign outputs[986] = ~((layer0_outputs[873]) ^ (layer0_outputs[734]));
    assign outputs[987] = layer0_outputs[1653];
    assign outputs[988] = (layer0_outputs[2147]) & ~(layer0_outputs[1001]);
    assign outputs[989] = ~((layer0_outputs[387]) ^ (layer0_outputs[843]));
    assign outputs[990] = (layer0_outputs[1201]) & ~(layer0_outputs[2475]);
    assign outputs[991] = ~(layer0_outputs[1662]);
    assign outputs[992] = (layer0_outputs[1704]) & (layer0_outputs[2081]);
    assign outputs[993] = ~((layer0_outputs[1074]) | (layer0_outputs[722]));
    assign outputs[994] = (layer0_outputs[1939]) ^ (layer0_outputs[128]);
    assign outputs[995] = ~((layer0_outputs[2335]) | (layer0_outputs[1302]));
    assign outputs[996] = ~(layer0_outputs[486]);
    assign outputs[997] = (layer0_outputs[2026]) ^ (layer0_outputs[1674]);
    assign outputs[998] = ~(layer0_outputs[2114]) | (layer0_outputs[1883]);
    assign outputs[999] = layer0_outputs[441];
    assign outputs[1000] = ~(layer0_outputs[2176]) | (layer0_outputs[1256]);
    assign outputs[1001] = ~((layer0_outputs[2447]) | (layer0_outputs[1409]));
    assign outputs[1002] = ~(layer0_outputs[1406]);
    assign outputs[1003] = ~(layer0_outputs[611]);
    assign outputs[1004] = ~(layer0_outputs[1720]);
    assign outputs[1005] = (layer0_outputs[1505]) & ~(layer0_outputs[275]);
    assign outputs[1006] = ~((layer0_outputs[2205]) ^ (layer0_outputs[2259]));
    assign outputs[1007] = layer0_outputs[728];
    assign outputs[1008] = ~((layer0_outputs[228]) | (layer0_outputs[360]));
    assign outputs[1009] = ~(layer0_outputs[1115]);
    assign outputs[1010] = ~(layer0_outputs[1322]);
    assign outputs[1011] = ~((layer0_outputs[1511]) ^ (layer0_outputs[507]));
    assign outputs[1012] = (layer0_outputs[1778]) & ~(layer0_outputs[250]);
    assign outputs[1013] = layer0_outputs[1866];
    assign outputs[1014] = layer0_outputs[272];
    assign outputs[1015] = ~(layer0_outputs[556]);
    assign outputs[1016] = (layer0_outputs[2160]) & ~(layer0_outputs[283]);
    assign outputs[1017] = (layer0_outputs[1236]) & ~(layer0_outputs[1425]);
    assign outputs[1018] = (layer0_outputs[2365]) & ~(layer0_outputs[537]);
    assign outputs[1019] = (layer0_outputs[1951]) | (layer0_outputs[613]);
    assign outputs[1020] = ~(layer0_outputs[1093]) | (layer0_outputs[294]);
    assign outputs[1021] = ~(layer0_outputs[1927]);
    assign outputs[1022] = (layer0_outputs[2184]) & (layer0_outputs[841]);
    assign outputs[1023] = ~((layer0_outputs[2420]) | (layer0_outputs[368]));
    assign outputs[1024] = (layer0_outputs[1876]) ^ (layer0_outputs[34]);
    assign outputs[1025] = layer0_outputs[2267];
    assign outputs[1026] = layer0_outputs[504];
    assign outputs[1027] = (layer0_outputs[2397]) & ~(layer0_outputs[1840]);
    assign outputs[1028] = (layer0_outputs[272]) & ~(layer0_outputs[857]);
    assign outputs[1029] = (layer0_outputs[2024]) & ~(layer0_outputs[612]);
    assign outputs[1030] = (layer0_outputs[872]) & (layer0_outputs[1886]);
    assign outputs[1031] = (layer0_outputs[2212]) & ~(layer0_outputs[1932]);
    assign outputs[1032] = (layer0_outputs[1319]) & ~(layer0_outputs[477]);
    assign outputs[1033] = ~(layer0_outputs[389]) | (layer0_outputs[1623]);
    assign outputs[1034] = ~((layer0_outputs[1631]) ^ (layer0_outputs[975]));
    assign outputs[1035] = layer0_outputs[637];
    assign outputs[1036] = layer0_outputs[2050];
    assign outputs[1037] = ~(layer0_outputs[2493]);
    assign outputs[1038] = ~((layer0_outputs[1745]) | (layer0_outputs[1064]));
    assign outputs[1039] = ~(layer0_outputs[348]);
    assign outputs[1040] = ~((layer0_outputs[1290]) & (layer0_outputs[814]));
    assign outputs[1041] = ~((layer0_outputs[1324]) ^ (layer0_outputs[1860]));
    assign outputs[1042] = ~(layer0_outputs[1661]);
    assign outputs[1043] = ~(layer0_outputs[499]);
    assign outputs[1044] = ~((layer0_outputs[592]) ^ (layer0_outputs[1862]));
    assign outputs[1045] = (layer0_outputs[823]) & (layer0_outputs[450]);
    assign outputs[1046] = (layer0_outputs[1760]) & (layer0_outputs[61]);
    assign outputs[1047] = ~(layer0_outputs[493]);
    assign outputs[1048] = ~((layer0_outputs[1020]) | (layer0_outputs[1443]));
    assign outputs[1049] = (layer0_outputs[2069]) & ~(layer0_outputs[167]);
    assign outputs[1050] = ~((layer0_outputs[1455]) ^ (layer0_outputs[1250]));
    assign outputs[1051] = (layer0_outputs[2453]) & ~(layer0_outputs[87]);
    assign outputs[1052] = ~((layer0_outputs[2229]) | (layer0_outputs[1466]));
    assign outputs[1053] = (layer0_outputs[205]) & (layer0_outputs[143]);
    assign outputs[1054] = layer0_outputs[1336];
    assign outputs[1055] = ~((layer0_outputs[762]) ^ (layer0_outputs[667]));
    assign outputs[1056] = (layer0_outputs[2263]) ^ (layer0_outputs[2447]);
    assign outputs[1057] = ~((layer0_outputs[467]) ^ (layer0_outputs[490]));
    assign outputs[1058] = ~(layer0_outputs[449]);
    assign outputs[1059] = ~(layer0_outputs[1973]);
    assign outputs[1060] = layer0_outputs[1389];
    assign outputs[1061] = (layer0_outputs[212]) & ~(layer0_outputs[2087]);
    assign outputs[1062] = (layer0_outputs[1366]) & ~(layer0_outputs[1318]);
    assign outputs[1063] = layer0_outputs[498];
    assign outputs[1064] = (layer0_outputs[1461]) ^ (layer0_outputs[1208]);
    assign outputs[1065] = ~((layer0_outputs[1183]) | (layer0_outputs[1924]));
    assign outputs[1066] = (layer0_outputs[1732]) & (layer0_outputs[2478]);
    assign outputs[1067] = (layer0_outputs[773]) | (layer0_outputs[251]);
    assign outputs[1068] = (layer0_outputs[1377]) & ~(layer0_outputs[29]);
    assign outputs[1069] = (layer0_outputs[22]) & ~(layer0_outputs[12]);
    assign outputs[1070] = ~(layer0_outputs[96]);
    assign outputs[1071] = layer0_outputs[1006];
    assign outputs[1072] = layer0_outputs[1671];
    assign outputs[1073] = (layer0_outputs[1325]) & ~(layer0_outputs[1796]);
    assign outputs[1074] = layer0_outputs[1438];
    assign outputs[1075] = (layer0_outputs[197]) & ~(layer0_outputs[639]);
    assign outputs[1076] = ~(layer0_outputs[2071]) | (layer0_outputs[843]);
    assign outputs[1077] = layer0_outputs[527];
    assign outputs[1078] = ~((layer0_outputs[916]) ^ (layer0_outputs[1251]));
    assign outputs[1079] = layer0_outputs[4];
    assign outputs[1080] = layer0_outputs[2304];
    assign outputs[1081] = ~(layer0_outputs[886]);
    assign outputs[1082] = layer0_outputs[1412];
    assign outputs[1083] = layer0_outputs[2118];
    assign outputs[1084] = (layer0_outputs[2027]) ^ (layer0_outputs[2336]);
    assign outputs[1085] = (layer0_outputs[515]) & ~(layer0_outputs[2466]);
    assign outputs[1086] = ~((layer0_outputs[1592]) | (layer0_outputs[926]));
    assign outputs[1087] = layer0_outputs[527];
    assign outputs[1088] = ~(layer0_outputs[1524]);
    assign outputs[1089] = ~(layer0_outputs[1635]) | (layer0_outputs[1027]);
    assign outputs[1090] = ~(layer0_outputs[879]);
    assign outputs[1091] = layer0_outputs[1105];
    assign outputs[1092] = (layer0_outputs[2335]) & ~(layer0_outputs[1759]);
    assign outputs[1093] = ~((layer0_outputs[1341]) | (layer0_outputs[789]));
    assign outputs[1094] = ~((layer0_outputs[1877]) | (layer0_outputs[853]));
    assign outputs[1095] = ~(layer0_outputs[1042]) | (layer0_outputs[600]);
    assign outputs[1096] = ~((layer0_outputs[2101]) ^ (layer0_outputs[473]));
    assign outputs[1097] = (layer0_outputs[2407]) & (layer0_outputs[64]);
    assign outputs[1098] = (layer0_outputs[829]) ^ (layer0_outputs[1203]);
    assign outputs[1099] = ~(layer0_outputs[45]) | (layer0_outputs[1608]);
    assign outputs[1100] = (layer0_outputs[1697]) & (layer0_outputs[2222]);
    assign outputs[1101] = (layer0_outputs[914]) & ~(layer0_outputs[845]);
    assign outputs[1102] = layer0_outputs[2003];
    assign outputs[1103] = ~((layer0_outputs[911]) ^ (layer0_outputs[1113]));
    assign outputs[1104] = (layer0_outputs[189]) & ~(layer0_outputs[1577]);
    assign outputs[1105] = (layer0_outputs[2313]) & ~(layer0_outputs[1553]);
    assign outputs[1106] = (layer0_outputs[1557]) | (layer0_outputs[657]);
    assign outputs[1107] = ~(layer0_outputs[21]) | (layer0_outputs[968]);
    assign outputs[1108] = ~(layer0_outputs[1591]);
    assign outputs[1109] = ~((layer0_outputs[634]) ^ (layer0_outputs[917]));
    assign outputs[1110] = ~((layer0_outputs[2018]) & (layer0_outputs[892]));
    assign outputs[1111] = ~(layer0_outputs[719]);
    assign outputs[1112] = (layer0_outputs[695]) ^ (layer0_outputs[907]);
    assign outputs[1113] = ~(layer0_outputs[1693]);
    assign outputs[1114] = ~(layer0_outputs[984]);
    assign outputs[1115] = ~(layer0_outputs[2399]);
    assign outputs[1116] = ~(layer0_outputs[589]);
    assign outputs[1117] = ~(layer0_outputs[1718]);
    assign outputs[1118] = (layer0_outputs[990]) & (layer0_outputs[445]);
    assign outputs[1119] = ~((layer0_outputs[755]) | (layer0_outputs[555]));
    assign outputs[1120] = (layer0_outputs[1851]) & ~(layer0_outputs[1650]);
    assign outputs[1121] = ~(layer0_outputs[1645]);
    assign outputs[1122] = (layer0_outputs[124]) ^ (layer0_outputs[1950]);
    assign outputs[1123] = ~(layer0_outputs[1291]);
    assign outputs[1124] = (layer0_outputs[1395]) | (layer0_outputs[2381]);
    assign outputs[1125] = layer0_outputs[150];
    assign outputs[1126] = ~(layer0_outputs[491]);
    assign outputs[1127] = ~(layer0_outputs[1973]);
    assign outputs[1128] = (layer0_outputs[38]) & (layer0_outputs[1914]);
    assign outputs[1129] = ~(layer0_outputs[211]) | (layer0_outputs[860]);
    assign outputs[1130] = (layer0_outputs[1634]) | (layer0_outputs[1761]);
    assign outputs[1131] = (layer0_outputs[465]) & ~(layer0_outputs[2255]);
    assign outputs[1132] = (layer0_outputs[455]) & ~(layer0_outputs[2256]);
    assign outputs[1133] = (layer0_outputs[1811]) & ~(layer0_outputs[10]);
    assign outputs[1134] = ~(layer0_outputs[886]);
    assign outputs[1135] = ~(layer0_outputs[2430]);
    assign outputs[1136] = layer0_outputs[626];
    assign outputs[1137] = ~(layer0_outputs[1541]);
    assign outputs[1138] = (layer0_outputs[587]) | (layer0_outputs[132]);
    assign outputs[1139] = layer0_outputs[1600];
    assign outputs[1140] = layer0_outputs[325];
    assign outputs[1141] = layer0_outputs[1174];
    assign outputs[1142] = (layer0_outputs[375]) & ~(layer0_outputs[2075]);
    assign outputs[1143] = ~(layer0_outputs[1552]);
    assign outputs[1144] = (layer0_outputs[79]) & ~(layer0_outputs[540]);
    assign outputs[1145] = ~(layer0_outputs[2293]);
    assign outputs[1146] = layer0_outputs[305];
    assign outputs[1147] = ~((layer0_outputs[518]) | (layer0_outputs[873]));
    assign outputs[1148] = (layer0_outputs[2251]) & ~(layer0_outputs[2193]);
    assign outputs[1149] = layer0_outputs[2009];
    assign outputs[1150] = ~(layer0_outputs[1098]);
    assign outputs[1151] = ~((layer0_outputs[202]) ^ (layer0_outputs[2041]));
    assign outputs[1152] = ~(layer0_outputs[1190]) | (layer0_outputs[1869]);
    assign outputs[1153] = (layer0_outputs[1943]) & ~(layer0_outputs[2377]);
    assign outputs[1154] = ~(layer0_outputs[1429]);
    assign outputs[1155] = ~((layer0_outputs[2323]) | (layer0_outputs[17]));
    assign outputs[1156] = ~(layer0_outputs[2196]);
    assign outputs[1157] = layer0_outputs[1573];
    assign outputs[1158] = ~(layer0_outputs[847]) | (layer0_outputs[1841]);
    assign outputs[1159] = layer0_outputs[1204];
    assign outputs[1160] = (layer0_outputs[551]) & ~(layer0_outputs[581]);
    assign outputs[1161] = (layer0_outputs[2231]) & ~(layer0_outputs[292]);
    assign outputs[1162] = layer0_outputs[626];
    assign outputs[1163] = ~((layer0_outputs[1870]) ^ (layer0_outputs[40]));
    assign outputs[1164] = (layer0_outputs[166]) | (layer0_outputs[2013]);
    assign outputs[1165] = (layer0_outputs[1218]) ^ (layer0_outputs[1756]);
    assign outputs[1166] = ~(layer0_outputs[1084]);
    assign outputs[1167] = (layer0_outputs[1827]) ^ (layer0_outputs[489]);
    assign outputs[1168] = (layer0_outputs[1415]) & ~(layer0_outputs[717]);
    assign outputs[1169] = ~(layer0_outputs[460]);
    assign outputs[1170] = (layer0_outputs[315]) & ~(layer0_outputs[1320]);
    assign outputs[1171] = (layer0_outputs[1648]) & ~(layer0_outputs[845]);
    assign outputs[1172] = (layer0_outputs[880]) & (layer0_outputs[662]);
    assign outputs[1173] = ~(layer0_outputs[1788]) | (layer0_outputs[2309]);
    assign outputs[1174] = ~(layer0_outputs[1913]);
    assign outputs[1175] = (layer0_outputs[560]) & ~(layer0_outputs[171]);
    assign outputs[1176] = (layer0_outputs[196]) & ~(layer0_outputs[707]);
    assign outputs[1177] = (layer0_outputs[1622]) & (layer0_outputs[658]);
    assign outputs[1178] = ~((layer0_outputs[1898]) & (layer0_outputs[1578]));
    assign outputs[1179] = layer0_outputs[1943];
    assign outputs[1180] = ~((layer0_outputs[1824]) & (layer0_outputs[556]));
    assign outputs[1181] = (layer0_outputs[2173]) | (layer0_outputs[515]);
    assign outputs[1182] = (layer0_outputs[638]) & ~(layer0_outputs[2194]);
    assign outputs[1183] = (layer0_outputs[153]) ^ (layer0_outputs[893]);
    assign outputs[1184] = layer0_outputs[1690];
    assign outputs[1185] = ~((layer0_outputs[1148]) ^ (layer0_outputs[1383]));
    assign outputs[1186] = layer0_outputs[1069];
    assign outputs[1187] = (layer0_outputs[2168]) & ~(layer0_outputs[900]);
    assign outputs[1188] = ~((layer0_outputs[325]) ^ (layer0_outputs[1418]));
    assign outputs[1189] = ~(layer0_outputs[1119]) | (layer0_outputs[1159]);
    assign outputs[1190] = ~(layer0_outputs[2423]) | (layer0_outputs[406]);
    assign outputs[1191] = (layer0_outputs[85]) & ~(layer0_outputs[2442]);
    assign outputs[1192] = layer0_outputs[971];
    assign outputs[1193] = layer0_outputs[251];
    assign outputs[1194] = ~(layer0_outputs[993]);
    assign outputs[1195] = (layer0_outputs[1869]) & ~(layer0_outputs[813]);
    assign outputs[1196] = ~(layer0_outputs[82]);
    assign outputs[1197] = layer0_outputs[1087];
    assign outputs[1198] = ~((layer0_outputs[1263]) ^ (layer0_outputs[1471]));
    assign outputs[1199] = layer0_outputs[1641];
    assign outputs[1200] = layer0_outputs[358];
    assign outputs[1201] = ~((layer0_outputs[857]) | (layer0_outputs[2053]));
    assign outputs[1202] = ~(layer0_outputs[1717]);
    assign outputs[1203] = (layer0_outputs[1269]) & ~(layer0_outputs[528]);
    assign outputs[1204] = ~(layer0_outputs[713]);
    assign outputs[1205] = layer0_outputs[628];
    assign outputs[1206] = (layer0_outputs[1848]) & (layer0_outputs[1598]);
    assign outputs[1207] = layer0_outputs[1238];
    assign outputs[1208] = ~(layer0_outputs[2237]);
    assign outputs[1209] = (layer0_outputs[36]) & (layer0_outputs[1003]);
    assign outputs[1210] = (layer0_outputs[314]) & ~(layer0_outputs[1173]);
    assign outputs[1211] = ~(layer0_outputs[850]);
    assign outputs[1212] = (layer0_outputs[2203]) ^ (layer0_outputs[1919]);
    assign outputs[1213] = (layer0_outputs[1732]) & ~(layer0_outputs[528]);
    assign outputs[1214] = (layer0_outputs[1438]) & ~(layer0_outputs[2095]);
    assign outputs[1215] = ~(layer0_outputs[645]);
    assign outputs[1216] = (layer0_outputs[1027]) ^ (layer0_outputs[1136]);
    assign outputs[1217] = layer0_outputs[767];
    assign outputs[1218] = (layer0_outputs[1831]) & ~(layer0_outputs[262]);
    assign outputs[1219] = (layer0_outputs[2218]) & (layer0_outputs[2299]);
    assign outputs[1220] = ~((layer0_outputs[2099]) | (layer0_outputs[2126]));
    assign outputs[1221] = layer0_outputs[727];
    assign outputs[1222] = layer0_outputs[1088];
    assign outputs[1223] = (layer0_outputs[1813]) & (layer0_outputs[1437]);
    assign outputs[1224] = ~(layer0_outputs[1964]) | (layer0_outputs[465]);
    assign outputs[1225] = layer0_outputs[2157];
    assign outputs[1226] = (layer0_outputs[127]) & ~(layer0_outputs[1176]);
    assign outputs[1227] = (layer0_outputs[2440]) & (layer0_outputs[469]);
    assign outputs[1228] = layer0_outputs[1272];
    assign outputs[1229] = layer0_outputs[1885];
    assign outputs[1230] = ~((layer0_outputs[257]) & (layer0_outputs[1879]));
    assign outputs[1231] = ~((layer0_outputs[2007]) ^ (layer0_outputs[1364]));
    assign outputs[1232] = ~((layer0_outputs[270]) & (layer0_outputs[920]));
    assign outputs[1233] = (layer0_outputs[2013]) | (layer0_outputs[1482]);
    assign outputs[1234] = (layer0_outputs[305]) & ~(layer0_outputs[2155]);
    assign outputs[1235] = layer0_outputs[856];
    assign outputs[1236] = ~(layer0_outputs[2126]);
    assign outputs[1237] = ~((layer0_outputs[1007]) | (layer0_outputs[2213]));
    assign outputs[1238] = (layer0_outputs[35]) & ~(layer0_outputs[320]);
    assign outputs[1239] = ~(layer0_outputs[163]) | (layer0_outputs[889]);
    assign outputs[1240] = layer0_outputs[151];
    assign outputs[1241] = (layer0_outputs[2078]) & (layer0_outputs[2483]);
    assign outputs[1242] = ~(layer0_outputs[2112]);
    assign outputs[1243] = (layer0_outputs[1692]) & (layer0_outputs[971]);
    assign outputs[1244] = ~((layer0_outputs[1835]) ^ (layer0_outputs[184]));
    assign outputs[1245] = ~(layer0_outputs[1452]);
    assign outputs[1246] = ~((layer0_outputs[776]) | (layer0_outputs[1297]));
    assign outputs[1247] = (layer0_outputs[2138]) & ~(layer0_outputs[1068]);
    assign outputs[1248] = (layer0_outputs[1311]) & (layer0_outputs[1678]);
    assign outputs[1249] = ~((layer0_outputs[311]) ^ (layer0_outputs[1080]));
    assign outputs[1250] = ~((layer0_outputs[2171]) ^ (layer0_outputs[1449]));
    assign outputs[1251] = ~(layer0_outputs[2022]);
    assign outputs[1252] = (layer0_outputs[1490]) ^ (layer0_outputs[153]);
    assign outputs[1253] = ~(layer0_outputs[1863]) | (layer0_outputs[1766]);
    assign outputs[1254] = layer0_outputs[1080];
    assign outputs[1255] = (layer0_outputs[1264]) & ~(layer0_outputs[1780]);
    assign outputs[1256] = layer0_outputs[474];
    assign outputs[1257] = layer0_outputs[1014];
    assign outputs[1258] = layer0_outputs[1572];
    assign outputs[1259] = ~(layer0_outputs[546]) | (layer0_outputs[159]);
    assign outputs[1260] = (layer0_outputs[574]) & ~(layer0_outputs[925]);
    assign outputs[1261] = ~((layer0_outputs[1747]) | (layer0_outputs[1803]));
    assign outputs[1262] = layer0_outputs[149];
    assign outputs[1263] = layer0_outputs[1381];
    assign outputs[1264] = (layer0_outputs[1003]) ^ (layer0_outputs[267]);
    assign outputs[1265] = (layer0_outputs[1770]) & (layer0_outputs[2282]);
    assign outputs[1266] = (layer0_outputs[732]) & ~(layer0_outputs[1832]);
    assign outputs[1267] = layer0_outputs[1207];
    assign outputs[1268] = ~((layer0_outputs[1835]) ^ (layer0_outputs[911]));
    assign outputs[1269] = layer0_outputs[5];
    assign outputs[1270] = (layer0_outputs[1260]) | (layer0_outputs[2247]);
    assign outputs[1271] = ~((layer0_outputs[1643]) | (layer0_outputs[253]));
    assign outputs[1272] = (layer0_outputs[1258]) ^ (layer0_outputs[2303]);
    assign outputs[1273] = (layer0_outputs[1488]) | (layer0_outputs[1970]);
    assign outputs[1274] = ~((layer0_outputs[1359]) & (layer0_outputs[1053]));
    assign outputs[1275] = ~((layer0_outputs[1707]) ^ (layer0_outputs[1493]));
    assign outputs[1276] = ~(layer0_outputs[1112]);
    assign outputs[1277] = ~((layer0_outputs[1673]) | (layer0_outputs[952]));
    assign outputs[1278] = ~(layer0_outputs[1396]) | (layer0_outputs[114]);
    assign outputs[1279] = ~((layer0_outputs[1196]) ^ (layer0_outputs[233]));
    assign outputs[1280] = (layer0_outputs[1371]) & (layer0_outputs[1854]);
    assign outputs[1281] = layer0_outputs[2461];
    assign outputs[1282] = ~((layer0_outputs[860]) | (layer0_outputs[277]));
    assign outputs[1283] = (layer0_outputs[1434]) & ~(layer0_outputs[1435]);
    assign outputs[1284] = ~(layer0_outputs[2257]);
    assign outputs[1285] = (layer0_outputs[1390]) & (layer0_outputs[1107]);
    assign outputs[1286] = ~((layer0_outputs[703]) ^ (layer0_outputs[41]));
    assign outputs[1287] = ~(layer0_outputs[347]) | (layer0_outputs[209]);
    assign outputs[1288] = (layer0_outputs[338]) ^ (layer0_outputs[2391]);
    assign outputs[1289] = (layer0_outputs[1594]) | (layer0_outputs[732]);
    assign outputs[1290] = layer0_outputs[685];
    assign outputs[1291] = (layer0_outputs[2385]) ^ (layer0_outputs[1596]);
    assign outputs[1292] = layer0_outputs[1971];
    assign outputs[1293] = layer0_outputs[2028];
    assign outputs[1294] = layer0_outputs[2119];
    assign outputs[1295] = layer0_outputs[1391];
    assign outputs[1296] = ~(layer0_outputs[1372]);
    assign outputs[1297] = ~(layer0_outputs[726]);
    assign outputs[1298] = (layer0_outputs[1830]) & ~(layer0_outputs[736]);
    assign outputs[1299] = layer0_outputs[1552];
    assign outputs[1300] = ~((layer0_outputs[651]) | (layer0_outputs[1681]));
    assign outputs[1301] = ~(layer0_outputs[740]);
    assign outputs[1302] = (layer0_outputs[2295]) & (layer0_outputs[1991]);
    assign outputs[1303] = (layer0_outputs[1715]) & ~(layer0_outputs[520]);
    assign outputs[1304] = ~((layer0_outputs[651]) ^ (layer0_outputs[659]));
    assign outputs[1305] = (layer0_outputs[1937]) ^ (layer0_outputs[63]);
    assign outputs[1306] = ~(layer0_outputs[234]);
    assign outputs[1307] = (layer0_outputs[5]) & ~(layer0_outputs[983]);
    assign outputs[1308] = (layer0_outputs[632]) & ~(layer0_outputs[2132]);
    assign outputs[1309] = ~((layer0_outputs[1996]) ^ (layer0_outputs[346]));
    assign outputs[1310] = layer0_outputs[2474];
    assign outputs[1311] = (layer0_outputs[136]) ^ (layer0_outputs[1961]);
    assign outputs[1312] = ~((layer0_outputs[913]) ^ (layer0_outputs[2062]));
    assign outputs[1313] = ~(layer0_outputs[2350]);
    assign outputs[1314] = (layer0_outputs[163]) ^ (layer0_outputs[1999]);
    assign outputs[1315] = ~(layer0_outputs[1195]);
    assign outputs[1316] = ~((layer0_outputs[1217]) ^ (layer0_outputs[201]));
    assign outputs[1317] = (layer0_outputs[2162]) | (layer0_outputs[1779]);
    assign outputs[1318] = layer0_outputs[2341];
    assign outputs[1319] = ~(layer0_outputs[125]);
    assign outputs[1320] = layer0_outputs[536];
    assign outputs[1321] = (layer0_outputs[1237]) ^ (layer0_outputs[905]);
    assign outputs[1322] = ~((layer0_outputs[156]) | (layer0_outputs[2438]));
    assign outputs[1323] = ~((layer0_outputs[791]) ^ (layer0_outputs[1442]));
    assign outputs[1324] = ~(layer0_outputs[218]);
    assign outputs[1325] = (layer0_outputs[1614]) & ~(layer0_outputs[2307]);
    assign outputs[1326] = (layer0_outputs[631]) & ~(layer0_outputs[1776]);
    assign outputs[1327] = ~(layer0_outputs[2429]);
    assign outputs[1328] = layer0_outputs[328];
    assign outputs[1329] = (layer0_outputs[1787]) & ~(layer0_outputs[2010]);
    assign outputs[1330] = ~(layer0_outputs[555]);
    assign outputs[1331] = ~((layer0_outputs[1009]) ^ (layer0_outputs[245]));
    assign outputs[1332] = ~((layer0_outputs[1142]) ^ (layer0_outputs[243]));
    assign outputs[1333] = ~((layer0_outputs[940]) ^ (layer0_outputs[1366]));
    assign outputs[1334] = layer0_outputs[630];
    assign outputs[1335] = ~((layer0_outputs[433]) & (layer0_outputs[102]));
    assign outputs[1336] = (layer0_outputs[694]) & ~(layer0_outputs[54]);
    assign outputs[1337] = ~((layer0_outputs[2321]) | (layer0_outputs[1043]));
    assign outputs[1338] = (layer0_outputs[2490]) & ~(layer0_outputs[702]);
    assign outputs[1339] = ~((layer0_outputs[601]) ^ (layer0_outputs[868]));
    assign outputs[1340] = (layer0_outputs[1229]) ^ (layer0_outputs[721]);
    assign outputs[1341] = layer0_outputs[1392];
    assign outputs[1342] = (layer0_outputs[877]) ^ (layer0_outputs[1367]);
    assign outputs[1343] = ~((layer0_outputs[2403]) ^ (layer0_outputs[33]));
    assign outputs[1344] = (layer0_outputs[2294]) ^ (layer0_outputs[1590]);
    assign outputs[1345] = ~((layer0_outputs[826]) | (layer0_outputs[746]));
    assign outputs[1346] = ~(layer0_outputs[1061]) | (layer0_outputs[1360]);
    assign outputs[1347] = layer0_outputs[1589];
    assign outputs[1348] = (layer0_outputs[1439]) | (layer0_outputs[444]);
    assign outputs[1349] = layer0_outputs[698];
    assign outputs[1350] = (layer0_outputs[2322]) & (layer0_outputs[1278]);
    assign outputs[1351] = (layer0_outputs[921]) ^ (layer0_outputs[2283]);
    assign outputs[1352] = (layer0_outputs[73]) & ~(layer0_outputs[1417]);
    assign outputs[1353] = ~((layer0_outputs[456]) ^ (layer0_outputs[702]));
    assign outputs[1354] = layer0_outputs[327];
    assign outputs[1355] = ~((layer0_outputs[898]) & (layer0_outputs[994]));
    assign outputs[1356] = (layer0_outputs[1688]) & ~(layer0_outputs[2419]);
    assign outputs[1357] = ~(layer0_outputs[38]);
    assign outputs[1358] = ~((layer0_outputs[998]) | (layer0_outputs[1272]));
    assign outputs[1359] = (layer0_outputs[1271]) & ~(layer0_outputs[1151]);
    assign outputs[1360] = ~((layer0_outputs[299]) ^ (layer0_outputs[2280]));
    assign outputs[1361] = ~((layer0_outputs[1542]) | (layer0_outputs[79]));
    assign outputs[1362] = ~(layer0_outputs[1578]);
    assign outputs[1363] = ~((layer0_outputs[1178]) ^ (layer0_outputs[1163]));
    assign outputs[1364] = layer0_outputs[2175];
    assign outputs[1365] = (layer0_outputs[907]) & (layer0_outputs[710]);
    assign outputs[1366] = ~((layer0_outputs[2296]) | (layer0_outputs[1758]));
    assign outputs[1367] = ~((layer0_outputs[623]) ^ (layer0_outputs[1470]));
    assign outputs[1368] = layer0_outputs[1499];
    assign outputs[1369] = ~(layer0_outputs[797]) | (layer0_outputs[2076]);
    assign outputs[1370] = layer0_outputs[2109];
    assign outputs[1371] = (layer0_outputs[230]) & ~(layer0_outputs[2301]);
    assign outputs[1372] = ~((layer0_outputs[1928]) | (layer0_outputs[43]));
    assign outputs[1373] = ~((layer0_outputs[990]) & (layer0_outputs[1266]));
    assign outputs[1374] = ~(layer0_outputs[1447]);
    assign outputs[1375] = (layer0_outputs[1418]) & (layer0_outputs[1980]);
    assign outputs[1376] = layer0_outputs[562];
    assign outputs[1377] = (layer0_outputs[1380]) & (layer0_outputs[1934]);
    assign outputs[1378] = (layer0_outputs[1911]) ^ (layer0_outputs[529]);
    assign outputs[1379] = (layer0_outputs[1532]) & (layer0_outputs[2209]);
    assign outputs[1380] = ~((layer0_outputs[2364]) ^ (layer0_outputs[333]));
    assign outputs[1381] = layer0_outputs[2117];
    assign outputs[1382] = layer0_outputs[1278];
    assign outputs[1383] = ~(layer0_outputs[84]);
    assign outputs[1384] = (layer0_outputs[1576]) & ~(layer0_outputs[1968]);
    assign outputs[1385] = ~((layer0_outputs[2498]) & (layer0_outputs[987]));
    assign outputs[1386] = layer0_outputs[999];
    assign outputs[1387] = ~((layer0_outputs[81]) & (layer0_outputs[46]));
    assign outputs[1388] = layer0_outputs[851];
    assign outputs[1389] = (layer0_outputs[2078]) & ~(layer0_outputs[1368]);
    assign outputs[1390] = (layer0_outputs[852]) ^ (layer0_outputs[1370]);
    assign outputs[1391] = (layer0_outputs[924]) & (layer0_outputs[2032]);
    assign outputs[1392] = ~(layer0_outputs[1513]);
    assign outputs[1393] = ~(layer0_outputs[257]) | (layer0_outputs[1766]);
    assign outputs[1394] = ~((layer0_outputs[2450]) ^ (layer0_outputs[559]));
    assign outputs[1395] = ~(layer0_outputs[1456]) | (layer0_outputs[1651]);
    assign outputs[1396] = (layer0_outputs[1149]) ^ (layer0_outputs[1175]);
    assign outputs[1397] = layer0_outputs[1580];
    assign outputs[1398] = ~(layer0_outputs[774]);
    assign outputs[1399] = ~((layer0_outputs[2224]) | (layer0_outputs[1358]));
    assign outputs[1400] = ~(layer0_outputs[1502]);
    assign outputs[1401] = (layer0_outputs[2346]) ^ (layer0_outputs[1255]);
    assign outputs[1402] = (layer0_outputs[1247]) ^ (layer0_outputs[154]);
    assign outputs[1403] = ~(layer0_outputs[141]);
    assign outputs[1404] = ~(layer0_outputs[585]) | (layer0_outputs[103]);
    assign outputs[1405] = layer0_outputs[1202];
    assign outputs[1406] = ~(layer0_outputs[1137]);
    assign outputs[1407] = (layer0_outputs[1123]) | (layer0_outputs[135]);
    assign outputs[1408] = (layer0_outputs[1748]) & ~(layer0_outputs[805]);
    assign outputs[1409] = ~(layer0_outputs[373]) | (layer0_outputs[2390]);
    assign outputs[1410] = (layer0_outputs[1387]) & ~(layer0_outputs[70]);
    assign outputs[1411] = layer0_outputs[2193];
    assign outputs[1412] = ~(layer0_outputs[1368]) | (layer0_outputs[1861]);
    assign outputs[1413] = ~((layer0_outputs[578]) ^ (layer0_outputs[1581]));
    assign outputs[1414] = ~(layer0_outputs[2481]);
    assign outputs[1415] = (layer0_outputs[1433]) ^ (layer0_outputs[743]);
    assign outputs[1416] = layer0_outputs[2040];
    assign outputs[1417] = (layer0_outputs[520]) ^ (layer0_outputs[616]);
    assign outputs[1418] = layer0_outputs[1436];
    assign outputs[1419] = (layer0_outputs[1462]) ^ (layer0_outputs[1479]);
    assign outputs[1420] = ~((layer0_outputs[1875]) | (layer0_outputs[83]));
    assign outputs[1421] = ~(layer0_outputs[997]);
    assign outputs[1422] = ~((layer0_outputs[2265]) | (layer0_outputs[1468]));
    assign outputs[1423] = (layer0_outputs[2305]) ^ (layer0_outputs[1815]);
    assign outputs[1424] = ~(layer0_outputs[947]);
    assign outputs[1425] = (layer0_outputs[1016]) ^ (layer0_outputs[383]);
    assign outputs[1426] = layer0_outputs[1085];
    assign outputs[1427] = layer0_outputs[1309];
    assign outputs[1428] = layer0_outputs[1568];
    assign outputs[1429] = ~((layer0_outputs[2051]) & (layer0_outputs[2213]));
    assign outputs[1430] = (layer0_outputs[1760]) | (layer0_outputs[1398]);
    assign outputs[1431] = (layer0_outputs[664]) & ~(layer0_outputs[546]);
    assign outputs[1432] = ~(layer0_outputs[2465]);
    assign outputs[1433] = ~((layer0_outputs[1845]) ^ (layer0_outputs[2471]));
    assign outputs[1434] = layer0_outputs[2083];
    assign outputs[1435] = (layer0_outputs[1730]) & (layer0_outputs[2398]);
    assign outputs[1436] = ~((layer0_outputs[660]) ^ (layer0_outputs[986]));
    assign outputs[1437] = (layer0_outputs[1750]) & ~(layer0_outputs[1036]);
    assign outputs[1438] = ~((layer0_outputs[586]) ^ (layer0_outputs[346]));
    assign outputs[1439] = ~(layer0_outputs[302]);
    assign outputs[1440] = ~((layer0_outputs[872]) ^ (layer0_outputs[2072]));
    assign outputs[1441] = (layer0_outputs[2129]) & ~(layer0_outputs[25]);
    assign outputs[1442] = (layer0_outputs[634]) ^ (layer0_outputs[1577]);
    assign outputs[1443] = ~(layer0_outputs[596]);
    assign outputs[1444] = (layer0_outputs[1019]) ^ (layer0_outputs[671]);
    assign outputs[1445] = ~((layer0_outputs[359]) ^ (layer0_outputs[1407]));
    assign outputs[1446] = ~(layer0_outputs[955]) | (layer0_outputs[568]);
    assign outputs[1447] = (layer0_outputs[1329]) & ~(layer0_outputs[2010]);
    assign outputs[1448] = ~(layer0_outputs[2015]) | (layer0_outputs[2333]);
    assign outputs[1449] = ~((layer0_outputs[859]) & (layer0_outputs[1461]));
    assign outputs[1450] = (layer0_outputs[1509]) ^ (layer0_outputs[1225]);
    assign outputs[1451] = (layer0_outputs[2190]) ^ (layer0_outputs[407]);
    assign outputs[1452] = (layer0_outputs[539]) & (layer0_outputs[1529]);
    assign outputs[1453] = (layer0_outputs[291]) ^ (layer0_outputs[921]);
    assign outputs[1454] = layer0_outputs[1478];
    assign outputs[1455] = ~((layer0_outputs[647]) ^ (layer0_outputs[392]));
    assign outputs[1456] = ~((layer0_outputs[2435]) ^ (layer0_outputs[2484]));
    assign outputs[1457] = (layer0_outputs[953]) & ~(layer0_outputs[317]);
    assign outputs[1458] = (layer0_outputs[122]) ^ (layer0_outputs[378]);
    assign outputs[1459] = ~((layer0_outputs[779]) & (layer0_outputs[358]));
    assign outputs[1460] = (layer0_outputs[1275]) & ~(layer0_outputs[1280]);
    assign outputs[1461] = ~((layer0_outputs[2046]) ^ (layer0_outputs[381]));
    assign outputs[1462] = (layer0_outputs[993]) & (layer0_outputs[1652]);
    assign outputs[1463] = (layer0_outputs[2472]) & ~(layer0_outputs[1737]);
    assign outputs[1464] = ~(layer0_outputs[97]) | (layer0_outputs[683]);
    assign outputs[1465] = layer0_outputs[966];
    assign outputs[1466] = (layer0_outputs[1734]) | (layer0_outputs[1323]);
    assign outputs[1467] = ~((layer0_outputs[2464]) | (layer0_outputs[131]));
    assign outputs[1468] = layer0_outputs[2080];
    assign outputs[1469] = layer0_outputs[831];
    assign outputs[1470] = (layer0_outputs[1842]) ^ (layer0_outputs[1771]);
    assign outputs[1471] = ~(layer0_outputs[1247]);
    assign outputs[1472] = layer0_outputs[1590];
    assign outputs[1473] = (layer0_outputs[460]) ^ (layer0_outputs[2207]);
    assign outputs[1474] = ~((layer0_outputs[212]) ^ (layer0_outputs[141]));
    assign outputs[1475] = ~((layer0_outputs[1233]) ^ (layer0_outputs[1040]));
    assign outputs[1476] = (layer0_outputs[1477]) ^ (layer0_outputs[811]);
    assign outputs[1477] = (layer0_outputs[28]) ^ (layer0_outputs[2439]);
    assign outputs[1478] = ~((layer0_outputs[248]) ^ (layer0_outputs[2048]));
    assign outputs[1479] = (layer0_outputs[1448]) & ~(layer0_outputs[2090]);
    assign outputs[1480] = (layer0_outputs[707]) ^ (layer0_outputs[1393]);
    assign outputs[1481] = (layer0_outputs[2290]) ^ (layer0_outputs[2446]);
    assign outputs[1482] = ~((layer0_outputs[351]) & (layer0_outputs[1036]));
    assign outputs[1483] = ~(layer0_outputs[1099]);
    assign outputs[1484] = (layer0_outputs[328]) ^ (layer0_outputs[487]);
    assign outputs[1485] = ~(layer0_outputs[1895]);
    assign outputs[1486] = (layer0_outputs[1239]) & (layer0_outputs[592]);
    assign outputs[1487] = (layer0_outputs[2137]) & ~(layer0_outputs[2448]);
    assign outputs[1488] = (layer0_outputs[42]) ^ (layer0_outputs[1520]);
    assign outputs[1489] = ~((layer0_outputs[1057]) ^ (layer0_outputs[1583]));
    assign outputs[1490] = ~((layer0_outputs[19]) | (layer0_outputs[2379]));
    assign outputs[1491] = ~((layer0_outputs[1373]) ^ (layer0_outputs[1132]));
    assign outputs[1492] = ~((layer0_outputs[1865]) | (layer0_outputs[1545]));
    assign outputs[1493] = ~(layer0_outputs[50]);
    assign outputs[1494] = ~(layer0_outputs[2223]);
    assign outputs[1495] = layer0_outputs[725];
    assign outputs[1496] = ~((layer0_outputs[513]) | (layer0_outputs[1358]));
    assign outputs[1497] = ~((layer0_outputs[2279]) & (layer0_outputs[261]));
    assign outputs[1498] = (layer0_outputs[1492]) & ~(layer0_outputs[2327]);
    assign outputs[1499] = (layer0_outputs[620]) & ~(layer0_outputs[485]);
    assign outputs[1500] = layer0_outputs[1388];
    assign outputs[1501] = layer0_outputs[1327];
    assign outputs[1502] = (layer0_outputs[1974]) & ~(layer0_outputs[595]);
    assign outputs[1503] = ~((layer0_outputs[357]) | (layer0_outputs[1964]));
    assign outputs[1504] = ~(layer0_outputs[230]);
    assign outputs[1505] = ~(layer0_outputs[1084]);
    assign outputs[1506] = ~((layer0_outputs[3]) ^ (layer0_outputs[2297]));
    assign outputs[1507] = ~(layer0_outputs[2402]);
    assign outputs[1508] = ~((layer0_outputs[11]) ^ (layer0_outputs[2348]));
    assign outputs[1509] = ~(layer0_outputs[708]);
    assign outputs[1510] = ~((layer0_outputs[297]) & (layer0_outputs[2056]));
    assign outputs[1511] = ~((layer0_outputs[1813]) & (layer0_outputs[914]));
    assign outputs[1512] = ~(layer0_outputs[2455]) | (layer0_outputs[1216]);
    assign outputs[1513] = layer0_outputs[1410];
    assign outputs[1514] = (layer0_outputs[1219]) & (layer0_outputs[680]);
    assign outputs[1515] = ~(layer0_outputs[1497]) | (layer0_outputs[550]);
    assign outputs[1516] = ~((layer0_outputs[1246]) & (layer0_outputs[2410]));
    assign outputs[1517] = ~((layer0_outputs[1018]) ^ (layer0_outputs[1834]));
    assign outputs[1518] = (layer0_outputs[214]) & ~(layer0_outputs[787]);
    assign outputs[1519] = (layer0_outputs[660]) & ~(layer0_outputs[1296]);
    assign outputs[1520] = ~((layer0_outputs[530]) | (layer0_outputs[1181]));
    assign outputs[1521] = (layer0_outputs[2112]) & (layer0_outputs[622]);
    assign outputs[1522] = ~(layer0_outputs[1865]);
    assign outputs[1523] = ~(layer0_outputs[1624]);
    assign outputs[1524] = ~((layer0_outputs[1301]) ^ (layer0_outputs[572]));
    assign outputs[1525] = (layer0_outputs[1259]) ^ (layer0_outputs[1643]);
    assign outputs[1526] = layer0_outputs[1313];
    assign outputs[1527] = layer0_outputs[2452];
    assign outputs[1528] = (layer0_outputs[2415]) & ~(layer0_outputs[2343]);
    assign outputs[1529] = (layer0_outputs[823]) & ~(layer0_outputs[2320]);
    assign outputs[1530] = (layer0_outputs[413]) & ~(layer0_outputs[2268]);
    assign outputs[1531] = (layer0_outputs[1126]) | (layer0_outputs[870]);
    assign outputs[1532] = ~(layer0_outputs[324]);
    assign outputs[1533] = (layer0_outputs[233]) & (layer0_outputs[2227]);
    assign outputs[1534] = layer0_outputs[1049];
    assign outputs[1535] = ~((layer0_outputs[1710]) ^ (layer0_outputs[1938]));
    assign outputs[1536] = ~(layer0_outputs[617]);
    assign outputs[1537] = layer0_outputs[2280];
    assign outputs[1538] = ~((layer0_outputs[1803]) ^ (layer0_outputs[579]));
    assign outputs[1539] = layer0_outputs[2292];
    assign outputs[1540] = layer0_outputs[2055];
    assign outputs[1541] = (layer0_outputs[502]) ^ (layer0_outputs[94]);
    assign outputs[1542] = layer0_outputs[2016];
    assign outputs[1543] = ~((layer0_outputs[1850]) & (layer0_outputs[2356]));
    assign outputs[1544] = ~(layer0_outputs[796]);
    assign outputs[1545] = ~((layer0_outputs[335]) ^ (layer0_outputs[1297]));
    assign outputs[1546] = layer0_outputs[602];
    assign outputs[1547] = (layer0_outputs[774]) & ~(layer0_outputs[1118]);
    assign outputs[1548] = ~(layer0_outputs[464]);
    assign outputs[1549] = (layer0_outputs[31]) & ~(layer0_outputs[1224]);
    assign outputs[1550] = ~(layer0_outputs[509]);
    assign outputs[1551] = (layer0_outputs[1210]) ^ (layer0_outputs[461]);
    assign outputs[1552] = layer0_outputs[2085];
    assign outputs[1553] = (layer0_outputs[704]) & ~(layer0_outputs[1744]);
    assign outputs[1554] = ~((layer0_outputs[420]) ^ (layer0_outputs[1005]));
    assign outputs[1555] = ~(layer0_outputs[1708]) | (layer0_outputs[476]);
    assign outputs[1556] = layer0_outputs[2426];
    assign outputs[1557] = (layer0_outputs[1145]) & ~(layer0_outputs[1135]);
    assign outputs[1558] = layer0_outputs[1929];
    assign outputs[1559] = layer0_outputs[420];
    assign outputs[1560] = ~(layer0_outputs[42]);
    assign outputs[1561] = (layer0_outputs[1995]) & ~(layer0_outputs[1754]);
    assign outputs[1562] = ~(layer0_outputs[426]) | (layer0_outputs[2061]);
    assign outputs[1563] = ~(layer0_outputs[2380]) | (layer0_outputs[1464]);
    assign outputs[1564] = (layer0_outputs[1762]) & ~(layer0_outputs[1530]);
    assign outputs[1565] = (layer0_outputs[2019]) | (layer0_outputs[1519]);
    assign outputs[1566] = layer0_outputs[1853];
    assign outputs[1567] = (layer0_outputs[331]) & (layer0_outputs[1846]);
    assign outputs[1568] = (layer0_outputs[1473]) ^ (layer0_outputs[865]);
    assign outputs[1569] = (layer0_outputs[1071]) & ~(layer0_outputs[882]);
    assign outputs[1570] = ~(layer0_outputs[1032]);
    assign outputs[1571] = ~(layer0_outputs[1296]);
    assign outputs[1572] = layer0_outputs[1058];
    assign outputs[1573] = (layer0_outputs[658]) & (layer0_outputs[343]);
    assign outputs[1574] = ~(layer0_outputs[1225]);
    assign outputs[1575] = layer0_outputs[2392];
    assign outputs[1576] = ~(layer0_outputs[1512]);
    assign outputs[1577] = layer0_outputs[2164];
    assign outputs[1578] = ~(layer0_outputs[1823]);
    assign outputs[1579] = layer0_outputs[334];
    assign outputs[1580] = (layer0_outputs[1188]) & (layer0_outputs[2067]);
    assign outputs[1581] = ~(layer0_outputs[200]);
    assign outputs[1582] = ~((layer0_outputs[1594]) ^ (layer0_outputs[109]));
    assign outputs[1583] = layer0_outputs[263];
    assign outputs[1584] = (layer0_outputs[1300]) & ~(layer0_outputs[756]);
    assign outputs[1585] = layer0_outputs[2165];
    assign outputs[1586] = ~(layer0_outputs[34]) | (layer0_outputs[2014]);
    assign outputs[1587] = ~(layer0_outputs[2012]);
    assign outputs[1588] = (layer0_outputs[352]) & ~(layer0_outputs[65]);
    assign outputs[1589] = (layer0_outputs[1790]) & (layer0_outputs[159]);
    assign outputs[1590] = ~(layer0_outputs[1316]);
    assign outputs[1591] = ~(layer0_outputs[2422]);
    assign outputs[1592] = (layer0_outputs[1637]) & ~(layer0_outputs[2316]);
    assign outputs[1593] = ~(layer0_outputs[1712]);
    assign outputs[1594] = layer0_outputs[607];
    assign outputs[1595] = ~(layer0_outputs[1338]);
    assign outputs[1596] = (layer0_outputs[2118]) & ~(layer0_outputs[1053]);
    assign outputs[1597] = layer0_outputs[757];
    assign outputs[1598] = (layer0_outputs[1380]) & ~(layer0_outputs[794]);
    assign outputs[1599] = ~(layer0_outputs[769]);
    assign outputs[1600] = layer0_outputs[350];
    assign outputs[1601] = layer0_outputs[905];
    assign outputs[1602] = ~((layer0_outputs[1356]) ^ (layer0_outputs[1507]));
    assign outputs[1603] = ~((layer0_outputs[1868]) ^ (layer0_outputs[1219]));
    assign outputs[1604] = ~(layer0_outputs[939]) | (layer0_outputs[2141]);
    assign outputs[1605] = ~(layer0_outputs[1864]);
    assign outputs[1606] = ~(layer0_outputs[848]);
    assign outputs[1607] = ~((layer0_outputs[846]) | (layer0_outputs[2369]));
    assign outputs[1608] = (layer0_outputs[2018]) & ~(layer0_outputs[1878]);
    assign outputs[1609] = (layer0_outputs[414]) & (layer0_outputs[2276]);
    assign outputs[1610] = ~(layer0_outputs[772]) | (layer0_outputs[624]);
    assign outputs[1611] = ~((layer0_outputs[937]) ^ (layer0_outputs[416]));
    assign outputs[1612] = layer0_outputs[2242];
    assign outputs[1613] = layer0_outputs[1880];
    assign outputs[1614] = ~((layer0_outputs[1886]) | (layer0_outputs[1470]));
    assign outputs[1615] = layer0_outputs[2125];
    assign outputs[1616] = layer0_outputs[1472];
    assign outputs[1617] = ~(layer0_outputs[1638]) | (layer0_outputs[1588]);
    assign outputs[1618] = (layer0_outputs[580]) | (layer0_outputs[784]);
    assign outputs[1619] = (layer0_outputs[1873]) & ~(layer0_outputs[2127]);
    assign outputs[1620] = (layer0_outputs[1061]) | (layer0_outputs[91]);
    assign outputs[1621] = (layer0_outputs[1765]) & ~(layer0_outputs[2056]);
    assign outputs[1622] = ~((layer0_outputs[877]) | (layer0_outputs[1623]));
    assign outputs[1623] = ~((layer0_outputs[2438]) | (layer0_outputs[1801]));
    assign outputs[1624] = ~((layer0_outputs[604]) & (layer0_outputs[1914]));
    assign outputs[1625] = ~((layer0_outputs[1843]) | (layer0_outputs[2129]));
    assign outputs[1626] = ~(layer0_outputs[313]);
    assign outputs[1627] = (layer0_outputs[816]) ^ (layer0_outputs[106]);
    assign outputs[1628] = ~((layer0_outputs[246]) ^ (layer0_outputs[1714]));
    assign outputs[1629] = (layer0_outputs[865]) & (layer0_outputs[2445]);
    assign outputs[1630] = (layer0_outputs[2142]) & ~(layer0_outputs[2291]);
    assign outputs[1631] = (layer0_outputs[2308]) & ~(layer0_outputs[1262]);
    assign outputs[1632] = (layer0_outputs[1185]) & ~(layer0_outputs[131]);
    assign outputs[1633] = ~(layer0_outputs[2153]);
    assign outputs[1634] = (layer0_outputs[1559]) ^ (layer0_outputs[1561]);
    assign outputs[1635] = layer0_outputs[1207];
    assign outputs[1636] = layer0_outputs[2469];
    assign outputs[1637] = (layer0_outputs[2037]) ^ (layer0_outputs[500]);
    assign outputs[1638] = (layer0_outputs[1177]) | (layer0_outputs[1971]);
    assign outputs[1639] = ~((layer0_outputs[320]) | (layer0_outputs[377]));
    assign outputs[1640] = ~((layer0_outputs[379]) | (layer0_outputs[296]));
    assign outputs[1641] = ~(layer0_outputs[1546]);
    assign outputs[1642] = ~(layer0_outputs[1948]);
    assign outputs[1643] = ~((layer0_outputs[2206]) ^ (layer0_outputs[612]));
    assign outputs[1644] = ~((layer0_outputs[2395]) | (layer0_outputs[1625]));
    assign outputs[1645] = (layer0_outputs[1050]) & ~(layer0_outputs[418]);
    assign outputs[1646] = ~((layer0_outputs[1734]) | (layer0_outputs[1786]));
    assign outputs[1647] = ~(layer0_outputs[1211]) | (layer0_outputs[792]);
    assign outputs[1648] = layer0_outputs[518];
    assign outputs[1649] = ~((layer0_outputs[1419]) | (layer0_outputs[1451]));
    assign outputs[1650] = ~((layer0_outputs[1703]) | (layer0_outputs[2192]));
    assign outputs[1651] = (layer0_outputs[1375]) ^ (layer0_outputs[946]);
    assign outputs[1652] = layer0_outputs[1040];
    assign outputs[1653] = layer0_outputs[1384];
    assign outputs[1654] = ~(layer0_outputs[1250]);
    assign outputs[1655] = (layer0_outputs[466]) & ~(layer0_outputs[2382]);
    assign outputs[1656] = ~((layer0_outputs[570]) ^ (layer0_outputs[2420]));
    assign outputs[1657] = ~(layer0_outputs[2380]);
    assign outputs[1658] = (layer0_outputs[1052]) | (layer0_outputs[1162]);
    assign outputs[1659] = (layer0_outputs[1842]) & ~(layer0_outputs[1034]);
    assign outputs[1660] = layer0_outputs[529];
    assign outputs[1661] = ~((layer0_outputs[383]) | (layer0_outputs[252]));
    assign outputs[1662] = ~(layer0_outputs[1874]) | (layer0_outputs[1353]);
    assign outputs[1663] = (layer0_outputs[1517]) ^ (layer0_outputs[1712]);
    assign outputs[1664] = ~((layer0_outputs[1175]) & (layer0_outputs[1606]));
    assign outputs[1665] = ~(layer0_outputs[899]);
    assign outputs[1666] = ~((layer0_outputs[2276]) ^ (layer0_outputs[831]));
    assign outputs[1667] = (layer0_outputs[1616]) & (layer0_outputs[1982]);
    assign outputs[1668] = layer0_outputs[2232];
    assign outputs[1669] = ~(layer0_outputs[1032]);
    assign outputs[1670] = ~(layer0_outputs[972]);
    assign outputs[1671] = (layer0_outputs[2312]) & ~(layer0_outputs[312]);
    assign outputs[1672] = layer0_outputs[69];
    assign outputs[1673] = ~(layer0_outputs[2367]);
    assign outputs[1674] = (layer0_outputs[632]) & (layer0_outputs[275]);
    assign outputs[1675] = (layer0_outputs[1222]) & (layer0_outputs[1268]);
    assign outputs[1676] = layer0_outputs[2245];
    assign outputs[1677] = (layer0_outputs[2191]) & (layer0_outputs[2139]);
    assign outputs[1678] = layer0_outputs[1829];
    assign outputs[1679] = ~(layer0_outputs[805]);
    assign outputs[1680] = ~(layer0_outputs[2326]);
    assign outputs[1681] = ~((layer0_outputs[2405]) & (layer0_outputs[2117]));
    assign outputs[1682] = ~((layer0_outputs[110]) | (layer0_outputs[2250]));
    assign outputs[1683] = ~((layer0_outputs[780]) ^ (layer0_outputs[1044]));
    assign outputs[1684] = (layer0_outputs[2278]) ^ (layer0_outputs[836]);
    assign outputs[1685] = ~(layer0_outputs[1193]);
    assign outputs[1686] = ~((layer0_outputs[47]) ^ (layer0_outputs[1819]));
    assign outputs[1687] = ~((layer0_outputs[738]) & (layer0_outputs[1192]));
    assign outputs[1688] = ~(layer0_outputs[2249]);
    assign outputs[1689] = ~((layer0_outputs[394]) ^ (layer0_outputs[962]));
    assign outputs[1690] = layer0_outputs[1484];
    assign outputs[1691] = ~(layer0_outputs[27]);
    assign outputs[1692] = ~((layer0_outputs[1611]) & (layer0_outputs[288]));
    assign outputs[1693] = ~(layer0_outputs[988]);
    assign outputs[1694] = ~(layer0_outputs[1599]);
    assign outputs[1695] = (layer0_outputs[1174]) & ~(layer0_outputs[2170]);
    assign outputs[1696] = layer0_outputs[646];
    assign outputs[1697] = ~(layer0_outputs[397]);
    assign outputs[1698] = (layer0_outputs[882]) ^ (layer0_outputs[1059]);
    assign outputs[1699] = layer0_outputs[1531];
    assign outputs[1700] = ~(layer0_outputs[655]);
    assign outputs[1701] = ~(layer0_outputs[2071]);
    assign outputs[1702] = ~(layer0_outputs[897]);
    assign outputs[1703] = ~(layer0_outputs[1633]);
    assign outputs[1704] = layer0_outputs[1757];
    assign outputs[1705] = (layer0_outputs[1094]) | (layer0_outputs[1373]);
    assign outputs[1706] = layer0_outputs[1873];
    assign outputs[1707] = ~(layer0_outputs[1782]);
    assign outputs[1708] = (layer0_outputs[1576]) ^ (layer0_outputs[1386]);
    assign outputs[1709] = (layer0_outputs[223]) & (layer0_outputs[1821]);
    assign outputs[1710] = (layer0_outputs[1153]) & ~(layer0_outputs[1476]);
    assign outputs[1711] = ~((layer0_outputs[621]) | (layer0_outputs[1859]));
    assign outputs[1712] = layer0_outputs[1339];
    assign outputs[1713] = (layer0_outputs[1093]) & ~(layer0_outputs[1940]);
    assign outputs[1714] = ~(layer0_outputs[1332]);
    assign outputs[1715] = ~(layer0_outputs[1571]);
    assign outputs[1716] = layer0_outputs[2180];
    assign outputs[1717] = (layer0_outputs[1771]) & ~(layer0_outputs[116]);
    assign outputs[1718] = (layer0_outputs[287]) & ~(layer0_outputs[1775]);
    assign outputs[1719] = layer0_outputs[705];
    assign outputs[1720] = (layer0_outputs[1472]) & ~(layer0_outputs[2202]);
    assign outputs[1721] = (layer0_outputs[1276]) & ~(layer0_outputs[2102]);
    assign outputs[1722] = ~(layer0_outputs[2143]) | (layer0_outputs[1516]);
    assign outputs[1723] = ~((layer0_outputs[673]) & (layer0_outputs[267]));
    assign outputs[1724] = ~((layer0_outputs[720]) | (layer0_outputs[763]));
    assign outputs[1725] = (layer0_outputs[2289]) | (layer0_outputs[1514]);
    assign outputs[1726] = ~(layer0_outputs[1285]) | (layer0_outputs[883]);
    assign outputs[1727] = (layer0_outputs[438]) & (layer0_outputs[1006]);
    assign outputs[1728] = ~((layer0_outputs[1131]) | (layer0_outputs[1491]));
    assign outputs[1729] = (layer0_outputs[199]) & ~(layer0_outputs[1456]);
    assign outputs[1730] = (layer0_outputs[1811]) & (layer0_outputs[575]);
    assign outputs[1731] = layer0_outputs[2370];
    assign outputs[1732] = ~((layer0_outputs[2098]) | (layer0_outputs[1254]));
    assign outputs[1733] = layer0_outputs[156];
    assign outputs[1734] = ~(layer0_outputs[1328]);
    assign outputs[1735] = layer0_outputs[1967];
    assign outputs[1736] = ~(layer0_outputs[1566]) | (layer0_outputs[1255]);
    assign outputs[1737] = ~(layer0_outputs[2152]);
    assign outputs[1738] = ~(layer0_outputs[818]);
    assign outputs[1739] = ~(layer0_outputs[2320]);
    assign outputs[1740] = ~(layer0_outputs[2274]);
    assign outputs[1741] = (layer0_outputs[510]) & ~(layer0_outputs[1136]);
    assign outputs[1742] = ~((layer0_outputs[892]) & (layer0_outputs[2491]));
    assign outputs[1743] = layer0_outputs[1030];
    assign outputs[1744] = layer0_outputs[649];
    assign outputs[1745] = layer0_outputs[2240];
    assign outputs[1746] = layer0_outputs[338];
    assign outputs[1747] = ~(layer0_outputs[361]) | (layer0_outputs[72]);
    assign outputs[1748] = (layer0_outputs[2366]) ^ (layer0_outputs[1371]);
    assign outputs[1749] = (layer0_outputs[1307]) & ~(layer0_outputs[2097]);
    assign outputs[1750] = ~((layer0_outputs[484]) & (layer0_outputs[1223]));
    assign outputs[1751] = ~((layer0_outputs[39]) | (layer0_outputs[890]));
    assign outputs[1752] = (layer0_outputs[1468]) & ~(layer0_outputs[380]);
    assign outputs[1753] = layer0_outputs[2084];
    assign outputs[1754] = (layer0_outputs[1024]) & (layer0_outputs[2495]);
    assign outputs[1755] = (layer0_outputs[427]) & ~(layer0_outputs[1292]);
    assign outputs[1756] = (layer0_outputs[2043]) & ~(layer0_outputs[2156]);
    assign outputs[1757] = (layer0_outputs[28]) & ~(layer0_outputs[425]);
    assign outputs[1758] = layer0_outputs[2127];
    assign outputs[1759] = ~(layer0_outputs[1934]);
    assign outputs[1760] = ~(layer0_outputs[158]) | (layer0_outputs[2065]);
    assign outputs[1761] = ~(layer0_outputs[734]);
    assign outputs[1762] = (layer0_outputs[2463]) & ~(layer0_outputs[2135]);
    assign outputs[1763] = (layer0_outputs[696]) & ~(layer0_outputs[1961]);
    assign outputs[1764] = ~((layer0_outputs[999]) ^ (layer0_outputs[276]));
    assign outputs[1765] = (layer0_outputs[1872]) & ~(layer0_outputs[2100]);
    assign outputs[1766] = ~(layer0_outputs[2302]);
    assign outputs[1767] = ~((layer0_outputs[1508]) ^ (layer0_outputs[593]));
    assign outputs[1768] = ~(layer0_outputs[664]);
    assign outputs[1769] = ~((layer0_outputs[2241]) | (layer0_outputs[1548]));
    assign outputs[1770] = (layer0_outputs[1602]) & ~(layer0_outputs[1089]);
    assign outputs[1771] = (layer0_outputs[2258]) & ~(layer0_outputs[1487]);
    assign outputs[1772] = (layer0_outputs[1376]) & ~(layer0_outputs[557]);
    assign outputs[1773] = (layer0_outputs[155]) & (layer0_outputs[642]);
    assign outputs[1774] = (layer0_outputs[2479]) ^ (layer0_outputs[804]);
    assign outputs[1775] = ~(layer0_outputs[1147]) | (layer0_outputs[289]);
    assign outputs[1776] = (layer0_outputs[1859]) & ~(layer0_outputs[43]);
    assign outputs[1777] = (layer0_outputs[2095]) ^ (layer0_outputs[424]);
    assign outputs[1778] = layer0_outputs[1064];
    assign outputs[1779] = (layer0_outputs[1630]) & (layer0_outputs[1494]);
    assign outputs[1780] = layer0_outputs[1564];
    assign outputs[1781] = ~((layer0_outputs[705]) | (layer0_outputs[1753]));
    assign outputs[1782] = (layer0_outputs[1767]) & ~(layer0_outputs[2150]);
    assign outputs[1783] = (layer0_outputs[459]) ^ (layer0_outputs[2483]);
    assign outputs[1784] = layer0_outputs[318];
    assign outputs[1785] = ~((layer0_outputs[1137]) | (layer0_outputs[583]));
    assign outputs[1786] = layer0_outputs[463];
    assign outputs[1787] = (layer0_outputs[1308]) & ~(layer0_outputs[2215]);
    assign outputs[1788] = ~((layer0_outputs[2418]) & (layer0_outputs[1217]));
    assign outputs[1789] = (layer0_outputs[893]) & (layer0_outputs[2341]);
    assign outputs[1790] = ~(layer0_outputs[1558]);
    assign outputs[1791] = ~(layer0_outputs[687]) | (layer0_outputs[472]);
    assign outputs[1792] = ~((layer0_outputs[60]) ^ (layer0_outputs[2393]));
    assign outputs[1793] = (layer0_outputs[904]) & ~(layer0_outputs[1989]);
    assign outputs[1794] = (layer0_outputs[435]) ^ (layer0_outputs[1749]);
    assign outputs[1795] = ~((layer0_outputs[586]) & (layer0_outputs[9]));
    assign outputs[1796] = (layer0_outputs[1152]) & ~(layer0_outputs[668]);
    assign outputs[1797] = ~(layer0_outputs[372]);
    assign outputs[1798] = (layer0_outputs[689]) & ~(layer0_outputs[571]);
    assign outputs[1799] = layer0_outputs[621];
    assign outputs[1800] = layer0_outputs[226];
    assign outputs[1801] = (layer0_outputs[1374]) & (layer0_outputs[2378]);
    assign outputs[1802] = (layer0_outputs[1949]) & ~(layer0_outputs[995]);
    assign outputs[1803] = ~((layer0_outputs[126]) | (layer0_outputs[359]));
    assign outputs[1804] = (layer0_outputs[794]) & (layer0_outputs[1140]);
    assign outputs[1805] = ~(layer0_outputs[45]);
    assign outputs[1806] = (layer0_outputs[1063]) & (layer0_outputs[875]);
    assign outputs[1807] = ~((layer0_outputs[1462]) | (layer0_outputs[1560]));
    assign outputs[1808] = ~(layer0_outputs[2046]);
    assign outputs[1809] = layer0_outputs[887];
    assign outputs[1810] = ~((layer0_outputs[1642]) | (layer0_outputs[385]));
    assign outputs[1811] = ~(layer0_outputs[694]);
    assign outputs[1812] = ~(layer0_outputs[800]);
    assign outputs[1813] = ~((layer0_outputs[2044]) | (layer0_outputs[643]));
    assign outputs[1814] = layer0_outputs[2064];
    assign outputs[1815] = ~(layer0_outputs[1700]) | (layer0_outputs[949]);
    assign outputs[1816] = ~((layer0_outputs[1114]) ^ (layer0_outputs[304]));
    assign outputs[1817] = (layer0_outputs[146]) & ~(layer0_outputs[269]);
    assign outputs[1818] = layer0_outputs[719];
    assign outputs[1819] = ~((layer0_outputs[2338]) & (layer0_outputs[2199]));
    assign outputs[1820] = (layer0_outputs[1538]) | (layer0_outputs[866]);
    assign outputs[1821] = (layer0_outputs[1013]) ^ (layer0_outputs[561]);
    assign outputs[1822] = ~(layer0_outputs[814]) | (layer0_outputs[2298]);
    assign outputs[1823] = (layer0_outputs[1912]) & ~(layer0_outputs[1514]);
    assign outputs[1824] = (layer0_outputs[786]) & (layer0_outputs[924]);
    assign outputs[1825] = (layer0_outputs[742]) & ~(layer0_outputs[1795]);
    assign outputs[1826] = (layer0_outputs[186]) & ~(layer0_outputs[1935]);
    assign outputs[1827] = (layer0_outputs[231]) & (layer0_outputs[123]);
    assign outputs[1828] = ~((layer0_outputs[1213]) | (layer0_outputs[266]));
    assign outputs[1829] = layer0_outputs[200];
    assign outputs[1830] = ~(layer0_outputs[1289]);
    assign outputs[1831] = (layer0_outputs[300]) & ~(layer0_outputs[862]);
    assign outputs[1832] = ~((layer0_outputs[1788]) ^ (layer0_outputs[2200]));
    assign outputs[1833] = layer0_outputs[218];
    assign outputs[1834] = layer0_outputs[1718];
    assign outputs[1835] = (layer0_outputs[1312]) & ~(layer0_outputs[14]);
    assign outputs[1836] = ~(layer0_outputs[354]) | (layer0_outputs[2008]);
    assign outputs[1837] = (layer0_outputs[1335]) & ~(layer0_outputs[2391]);
    assign outputs[1838] = layer0_outputs[401];
    assign outputs[1839] = (layer0_outputs[2272]) ^ (layer0_outputs[688]);
    assign outputs[1840] = (layer0_outputs[1146]) ^ (layer0_outputs[447]);
    assign outputs[1841] = (layer0_outputs[2052]) & ~(layer0_outputs[445]);
    assign outputs[1842] = (layer0_outputs[866]) & ~(layer0_outputs[1167]);
    assign outputs[1843] = layer0_outputs[2172];
    assign outputs[1844] = ~((layer0_outputs[474]) ^ (layer0_outputs[99]));
    assign outputs[1845] = (layer0_outputs[395]) & ~(layer0_outputs[1197]);
    assign outputs[1846] = layer0_outputs[1752];
    assign outputs[1847] = ~(layer0_outputs[2131]) | (layer0_outputs[960]);
    assign outputs[1848] = (layer0_outputs[1077]) & (layer0_outputs[957]);
    assign outputs[1849] = ~((layer0_outputs[1183]) ^ (layer0_outputs[55]));
    assign outputs[1850] = ~((layer0_outputs[2390]) | (layer0_outputs[2058]));
    assign outputs[1851] = ~(layer0_outputs[2021]);
    assign outputs[1852] = ~((layer0_outputs[700]) | (layer0_outputs[109]));
    assign outputs[1853] = (layer0_outputs[840]) & ~(layer0_outputs[71]);
    assign outputs[1854] = (layer0_outputs[2093]) & ~(layer0_outputs[2412]);
    assign outputs[1855] = (layer0_outputs[1620]) ^ (layer0_outputs[2253]);
    assign outputs[1856] = (layer0_outputs[1304]) ^ (layer0_outputs[424]);
    assign outputs[1857] = (layer0_outputs[1830]) & ~(layer0_outputs[49]);
    assign outputs[1858] = (layer0_outputs[296]) & (layer0_outputs[1807]);
    assign outputs[1859] = layer0_outputs[730];
    assign outputs[1860] = (layer0_outputs[1048]) & ~(layer0_outputs[1290]);
    assign outputs[1861] = (layer0_outputs[2133]) & ~(layer0_outputs[1488]);
    assign outputs[1862] = layer0_outputs[1498];
    assign outputs[1863] = (layer0_outputs[2349]) & ~(layer0_outputs[1613]);
    assign outputs[1864] = layer0_outputs[1921];
    assign outputs[1865] = ~(layer0_outputs[812]);
    assign outputs[1866] = ~(layer0_outputs[2042]) | (layer0_outputs[1644]);
    assign outputs[1867] = layer0_outputs[1905];
    assign outputs[1868] = layer0_outputs[32];
    assign outputs[1869] = ~((layer0_outputs[890]) | (layer0_outputs[1715]));
    assign outputs[1870] = (layer0_outputs[2343]) | (layer0_outputs[1298]);
    assign outputs[1871] = ~(layer0_outputs[1483]) | (layer0_outputs[656]);
    assign outputs[1872] = (layer0_outputs[2319]) & ~(layer0_outputs[1303]);
    assign outputs[1873] = ~(layer0_outputs[2397]);
    assign outputs[1874] = ~(layer0_outputs[1588]) | (layer0_outputs[2383]);
    assign outputs[1875] = layer0_outputs[1333];
    assign outputs[1876] = (layer0_outputs[2488]) ^ (layer0_outputs[1816]);
    assign outputs[1877] = ~((layer0_outputs[113]) ^ (layer0_outputs[1031]));
    assign outputs[1878] = layer0_outputs[1851];
    assign outputs[1879] = (layer0_outputs[2315]) | (layer0_outputs[1035]);
    assign outputs[1880] = ~((layer0_outputs[1625]) & (layer0_outputs[1808]));
    assign outputs[1881] = (layer0_outputs[1723]) & (layer0_outputs[1823]);
    assign outputs[1882] = (layer0_outputs[2144]) | (layer0_outputs[2250]);
    assign outputs[1883] = ~(layer0_outputs[264]);
    assign outputs[1884] = ~(layer0_outputs[295]) | (layer0_outputs[1907]);
    assign outputs[1885] = layer0_outputs[2035];
    assign outputs[1886] = ~(layer0_outputs[1292]) | (layer0_outputs[741]);
    assign outputs[1887] = ~((layer0_outputs[266]) | (layer0_outputs[2166]));
    assign outputs[1888] = (layer0_outputs[1728]) | (layer0_outputs[2047]);
    assign outputs[1889] = (layer0_outputs[2096]) & ~(layer0_outputs[1985]);
    assign outputs[1890] = ~(layer0_outputs[1726]);
    assign outputs[1891] = ~(layer0_outputs[837]);
    assign outputs[1892] = ~(layer0_outputs[1683]) | (layer0_outputs[1931]);
    assign outputs[1893] = ~((layer0_outputs[2462]) ^ (layer0_outputs[582]));
    assign outputs[1894] = (layer0_outputs[1374]) & (layer0_outputs[2192]);
    assign outputs[1895] = layer0_outputs[2109];
    assign outputs[1896] = layer0_outputs[2361];
    assign outputs[1897] = ~(layer0_outputs[1344]);
    assign outputs[1898] = (layer0_outputs[1769]) & ~(layer0_outputs[584]);
    assign outputs[1899] = layer0_outputs[1793];
    assign outputs[1900] = (layer0_outputs[1011]) & ~(layer0_outputs[2485]);
    assign outputs[1901] = ~((layer0_outputs[105]) | (layer0_outputs[1655]));
    assign outputs[1902] = ~(layer0_outputs[1443]);
    assign outputs[1903] = ~(layer0_outputs[1645]);
    assign outputs[1904] = (layer0_outputs[1130]) & ~(layer0_outputs[677]);
    assign outputs[1905] = (layer0_outputs[608]) & ~(layer0_outputs[2363]);
    assign outputs[1906] = (layer0_outputs[1193]) & ~(layer0_outputs[307]);
    assign outputs[1907] = ~((layer0_outputs[1833]) ^ (layer0_outputs[1729]));
    assign outputs[1908] = ~((layer0_outputs[2331]) | (layer0_outputs[869]));
    assign outputs[1909] = (layer0_outputs[247]) & ~(layer0_outputs[688]);
    assign outputs[1910] = ~((layer0_outputs[1277]) ^ (layer0_outputs[2468]));
    assign outputs[1911] = ~(layer0_outputs[896]);
    assign outputs[1912] = (layer0_outputs[1782]) & (layer0_outputs[2038]);
    assign outputs[1913] = ~((layer0_outputs[1540]) | (layer0_outputs[1340]));
    assign outputs[1914] = ~((layer0_outputs[1621]) | (layer0_outputs[927]));
    assign outputs[1915] = layer0_outputs[2140];
    assign outputs[1916] = (layer0_outputs[1095]) ^ (layer0_outputs[960]);
    assign outputs[1917] = ~(layer0_outputs[615]);
    assign outputs[1918] = layer0_outputs[2188];
    assign outputs[1919] = (layer0_outputs[1849]) & (layer0_outputs[1857]);
    assign outputs[1920] = ~(layer0_outputs[274]) | (layer0_outputs[616]);
    assign outputs[1921] = layer0_outputs[1849];
    assign outputs[1922] = layer0_outputs[1686];
    assign outputs[1923] = (layer0_outputs[1954]) & ~(layer0_outputs[525]);
    assign outputs[1924] = layer0_outputs[2229];
    assign outputs[1925] = (layer0_outputs[2002]) & ~(layer0_outputs[682]);
    assign outputs[1926] = (layer0_outputs[1791]) & (layer0_outputs[1921]);
    assign outputs[1927] = ~((layer0_outputs[1657]) ^ (layer0_outputs[1573]));
    assign outputs[1928] = ~(layer0_outputs[931]);
    assign outputs[1929] = ~(layer0_outputs[1426]);
    assign outputs[1930] = layer0_outputs[2373];
    assign outputs[1931] = (layer0_outputs[204]) & ~(layer0_outputs[2179]);
    assign outputs[1932] = ~((layer0_outputs[2310]) ^ (layer0_outputs[1287]));
    assign outputs[1933] = layer0_outputs[1525];
    assign outputs[1934] = ~(layer0_outputs[2162]);
    assign outputs[1935] = ~((layer0_outputs[1826]) | (layer0_outputs[1213]));
    assign outputs[1936] = ~((layer0_outputs[681]) | (layer0_outputs[901]));
    assign outputs[1937] = (layer0_outputs[1562]) | (layer0_outputs[2330]);
    assign outputs[1938] = (layer0_outputs[1526]) | (layer0_outputs[386]);
    assign outputs[1939] = (layer0_outputs[1784]) ^ (layer0_outputs[419]);
    assign outputs[1940] = (layer0_outputs[1500]) & (layer0_outputs[1919]);
    assign outputs[1941] = ~(layer0_outputs[1768]);
    assign outputs[1942] = (layer0_outputs[879]) & ~(layer0_outputs[1845]);
    assign outputs[1943] = ~((layer0_outputs[1796]) | (layer0_outputs[1951]));
    assign outputs[1944] = ~((layer0_outputs[1768]) & (layer0_outputs[1295]));
    assign outputs[1945] = ~((layer0_outputs[322]) | (layer0_outputs[2344]));
    assign outputs[1946] = (layer0_outputs[1492]) & ~(layer0_outputs[542]);
    assign outputs[1947] = ~((layer0_outputs[581]) | (layer0_outputs[1848]));
    assign outputs[1948] = (layer0_outputs[1996]) & (layer0_outputs[952]);
    assign outputs[1949] = (layer0_outputs[1161]) & (layer0_outputs[285]);
    assign outputs[1950] = ~(layer0_outputs[704]);
    assign outputs[1951] = ~((layer0_outputs[2427]) & (layer0_outputs[278]));
    assign outputs[1952] = (layer0_outputs[2275]) ^ (layer0_outputs[1763]);
    assign outputs[1953] = layer0_outputs[446];
    assign outputs[1954] = (layer0_outputs[1928]) & ~(layer0_outputs[1245]);
    assign outputs[1955] = (layer0_outputs[75]) & ~(layer0_outputs[615]);
    assign outputs[1956] = (layer0_outputs[78]) & ~(layer0_outputs[489]);
    assign outputs[1957] = ~((layer0_outputs[237]) | (layer0_outputs[2347]));
    assign outputs[1958] = (layer0_outputs[1220]) & ~(layer0_outputs[303]);
    assign outputs[1959] = (layer0_outputs[2468]) & (layer0_outputs[1527]);
    assign outputs[1960] = (layer0_outputs[793]) ^ (layer0_outputs[2007]);
    assign outputs[1961] = (layer0_outputs[1335]) & ~(layer0_outputs[2245]);
    assign outputs[1962] = (layer0_outputs[1780]) & (layer0_outputs[399]);
    assign outputs[1963] = ~((layer0_outputs[1548]) ^ (layer0_outputs[353]));
    assign outputs[1964] = (layer0_outputs[2197]) ^ (layer0_outputs[2237]);
    assign outputs[1965] = ~((layer0_outputs[2433]) | (layer0_outputs[1264]));
    assign outputs[1966] = ~(layer0_outputs[1089]);
    assign outputs[1967] = (layer0_outputs[2234]) & ~(layer0_outputs[511]);
    assign outputs[1968] = ~(layer0_outputs[1340]);
    assign outputs[1969] = ~(layer0_outputs[521]) | (layer0_outputs[2498]);
    assign outputs[1970] = (layer0_outputs[1331]) & ~(layer0_outputs[222]);
    assign outputs[1971] = (layer0_outputs[2307]) & ~(layer0_outputs[2412]);
    assign outputs[1972] = ~(layer0_outputs[1129]);
    assign outputs[1973] = (layer0_outputs[1890]) & (layer0_outputs[1474]);
    assign outputs[1974] = (layer0_outputs[1347]) & ~(layer0_outputs[138]);
    assign outputs[1975] = ~(layer0_outputs[1107]);
    assign outputs[1976] = ~(layer0_outputs[609]);
    assign outputs[1977] = layer0_outputs[675];
    assign outputs[1978] = ~((layer0_outputs[1922]) ^ (layer0_outputs[1330]));
    assign outputs[1979] = (layer0_outputs[1624]) & (layer0_outputs[1713]);
    assign outputs[1980] = ~((layer0_outputs[107]) | (layer0_outputs[1705]));
    assign outputs[1981] = ~(layer0_outputs[143]);
    assign outputs[1982] = (layer0_outputs[1650]) & (layer0_outputs[1857]);
    assign outputs[1983] = (layer0_outputs[762]) & (layer0_outputs[1597]);
    assign outputs[1984] = (layer0_outputs[724]) ^ (layer0_outputs[2437]);
    assign outputs[1985] = ~(layer0_outputs[2425]);
    assign outputs[1986] = (layer0_outputs[1681]) & ~(layer0_outputs[2449]);
    assign outputs[1987] = ~((layer0_outputs[533]) | (layer0_outputs[1017]));
    assign outputs[1988] = (layer0_outputs[254]) & (layer0_outputs[2220]);
    assign outputs[1989] = (layer0_outputs[541]) ^ (layer0_outputs[779]);
    assign outputs[1990] = layer0_outputs[1420];
    assign outputs[1991] = (layer0_outputs[1913]) ^ (layer0_outputs[291]);
    assign outputs[1992] = (layer0_outputs[451]) & (layer0_outputs[343]);
    assign outputs[1993] = (layer0_outputs[1522]) & (layer0_outputs[731]);
    assign outputs[1994] = (layer0_outputs[432]) & (layer0_outputs[2351]);
    assign outputs[1995] = ~(layer0_outputs[1906]) | (layer0_outputs[2221]);
    assign outputs[1996] = ~(layer0_outputs[2000]) | (layer0_outputs[1884]);
    assign outputs[1997] = (layer0_outputs[1963]) | (layer0_outputs[472]);
    assign outputs[1998] = (layer0_outputs[565]) & (layer0_outputs[1527]);
    assign outputs[1999] = ~(layer0_outputs[1384]);
    assign outputs[2000] = ~(layer0_outputs[389]);
    assign outputs[2001] = layer0_outputs[264];
    assign outputs[2002] = ~((layer0_outputs[944]) & (layer0_outputs[1696]));
    assign outputs[2003] = (layer0_outputs[1266]) & ~(layer0_outputs[2357]);
    assign outputs[2004] = ~((layer0_outputs[88]) | (layer0_outputs[2489]));
    assign outputs[2005] = layer0_outputs[2287];
    assign outputs[2006] = (layer0_outputs[1361]) & ~(layer0_outputs[295]);
    assign outputs[2007] = (layer0_outputs[640]) & (layer0_outputs[531]);
    assign outputs[2008] = ~(layer0_outputs[2328]);
    assign outputs[2009] = ~((layer0_outputs[238]) & (layer0_outputs[2073]));
    assign outputs[2010] = ~(layer0_outputs[1882]) | (layer0_outputs[1798]);
    assign outputs[2011] = layer0_outputs[1033];
    assign outputs[2012] = layer0_outputs[293];
    assign outputs[2013] = ~((layer0_outputs[2329]) ^ (layer0_outputs[259]));
    assign outputs[2014] = (layer0_outputs[828]) ^ (layer0_outputs[505]);
    assign outputs[2015] = ~((layer0_outputs[437]) & (layer0_outputs[382]));
    assign outputs[2016] = (layer0_outputs[1187]) | (layer0_outputs[936]);
    assign outputs[2017] = layer0_outputs[558];
    assign outputs[2018] = (layer0_outputs[603]) & (layer0_outputs[48]);
    assign outputs[2019] = (layer0_outputs[476]) | (layer0_outputs[1856]);
    assign outputs[2020] = (layer0_outputs[144]) | (layer0_outputs[1559]);
    assign outputs[2021] = ~((layer0_outputs[2068]) ^ (layer0_outputs[434]));
    assign outputs[2022] = (layer0_outputs[2474]) ^ (layer0_outputs[1755]);
    assign outputs[2023] = (layer0_outputs[580]) | (layer0_outputs[152]);
    assign outputs[2024] = (layer0_outputs[1977]) ^ (layer0_outputs[1146]);
    assign outputs[2025] = ~(layer0_outputs[1100]);
    assign outputs[2026] = layer0_outputs[1724];
    assign outputs[2027] = (layer0_outputs[1069]) ^ (layer0_outputs[2005]);
    assign outputs[2028] = layer0_outputs[2311];
    assign outputs[2029] = ~((layer0_outputs[2259]) ^ (layer0_outputs[896]));
    assign outputs[2030] = ~((layer0_outputs[2031]) ^ (layer0_outputs[271]));
    assign outputs[2031] = (layer0_outputs[1904]) ^ (layer0_outputs[1058]);
    assign outputs[2032] = ~(layer0_outputs[1451]) | (layer0_outputs[1442]);
    assign outputs[2033] = ~(layer0_outputs[1936]);
    assign outputs[2034] = layer0_outputs[507];
    assign outputs[2035] = 1'b1;
    assign outputs[2036] = (layer0_outputs[2252]) | (layer0_outputs[1303]);
    assign outputs[2037] = layer0_outputs[903];
    assign outputs[2038] = ~((layer0_outputs[2120]) ^ (layer0_outputs[1216]));
    assign outputs[2039] = (layer0_outputs[1230]) | (layer0_outputs[1847]);
    assign outputs[2040] = (layer0_outputs[1138]) & (layer0_outputs[1821]);
    assign outputs[2041] = (layer0_outputs[2368]) & ~(layer0_outputs[1699]);
    assign outputs[2042] = ~((layer0_outputs[1096]) | (layer0_outputs[1196]));
    assign outputs[2043] = (layer0_outputs[2076]) ^ (layer0_outputs[2326]);
    assign outputs[2044] = layer0_outputs[1619];
    assign outputs[2045] = ~(layer0_outputs[1723]);
    assign outputs[2046] = ~((layer0_outputs[1809]) ^ (layer0_outputs[1984]));
    assign outputs[2047] = ~((layer0_outputs[1607]) | (layer0_outputs[1820]));
    assign outputs[2048] = ~(layer0_outputs[654]) | (layer0_outputs[1065]);
    assign outputs[2049] = (layer0_outputs[14]) | (layer0_outputs[855]);
    assign outputs[2050] = ~(layer0_outputs[904]);
    assign outputs[2051] = (layer0_outputs[2411]) ^ (layer0_outputs[679]);
    assign outputs[2052] = ~(layer0_outputs[1490]) | (layer0_outputs[1054]);
    assign outputs[2053] = ~((layer0_outputs[1473]) ^ (layer0_outputs[2454]));
    assign outputs[2054] = (layer0_outputs[1465]) & ~(layer0_outputs[895]);
    assign outputs[2055] = ~((layer0_outputs[160]) ^ (layer0_outputs[1121]));
    assign outputs[2056] = layer0_outputs[1563];
    assign outputs[2057] = ~(layer0_outputs[97]);
    assign outputs[2058] = ~(layer0_outputs[928]) | (layer0_outputs[1383]);
    assign outputs[2059] = ~(layer0_outputs[832]) | (layer0_outputs[362]);
    assign outputs[2060] = ~(layer0_outputs[1348]) | (layer0_outputs[2368]);
    assign outputs[2061] = ~((layer0_outputs[1998]) ^ (layer0_outputs[1299]));
    assign outputs[2062] = layer0_outputs[1743];
    assign outputs[2063] = (layer0_outputs[744]) ^ (layer0_outputs[2124]);
    assign outputs[2064] = ~(layer0_outputs[1351]) | (layer0_outputs[2299]);
    assign outputs[2065] = (layer0_outputs[2239]) & (layer0_outputs[2266]);
    assign outputs[2066] = ~(layer0_outputs[497]) | (layer0_outputs[1604]);
    assign outputs[2067] = ~(layer0_outputs[1]) | (layer0_outputs[1327]);
    assign outputs[2068] = ~((layer0_outputs[1352]) & (layer0_outputs[1238]));
    assign outputs[2069] = ~((layer0_outputs[1047]) ^ (layer0_outputs[1441]));
    assign outputs[2070] = ~(layer0_outputs[2206]);
    assign outputs[2071] = layer0_outputs[2147];
    assign outputs[2072] = ~(layer0_outputs[1227]);
    assign outputs[2073] = (layer0_outputs[1157]) & ~(layer0_outputs[1070]);
    assign outputs[2074] = ~(layer0_outputs[1693]);
    assign outputs[2075] = ~((layer0_outputs[71]) ^ (layer0_outputs[94]));
    assign outputs[2076] = ~(layer0_outputs[2436]) | (layer0_outputs[2219]);
    assign outputs[2077] = ~(layer0_outputs[1689]);
    assign outputs[2078] = (layer0_outputs[1691]) | (layer0_outputs[366]);
    assign outputs[2079] = (layer0_outputs[1421]) & ~(layer0_outputs[1381]);
    assign outputs[2080] = (layer0_outputs[1254]) & (layer0_outputs[1194]);
    assign outputs[2081] = ~((layer0_outputs[2094]) | (layer0_outputs[1362]));
    assign outputs[2082] = (layer0_outputs[958]) | (layer0_outputs[1993]);
    assign outputs[2083] = ~((layer0_outputs[782]) ^ (layer0_outputs[1269]));
    assign outputs[2084] = (layer0_outputs[1586]) ^ (layer0_outputs[1031]);
    assign outputs[2085] = ~((layer0_outputs[2235]) & (layer0_outputs[412]));
    assign outputs[2086] = (layer0_outputs[1897]) & (layer0_outputs[813]);
    assign outputs[2087] = ~((layer0_outputs[552]) ^ (layer0_outputs[365]));
    assign outputs[2088] = layer0_outputs[545];
    assign outputs[2089] = ~(layer0_outputs[1828]) | (layer0_outputs[1239]);
    assign outputs[2090] = ~(layer0_outputs[1836]) | (layer0_outputs[1923]);
    assign outputs[2091] = ~(layer0_outputs[2235]) | (layer0_outputs[286]);
    assign outputs[2092] = ~(layer0_outputs[1853]) | (layer0_outputs[1240]);
    assign outputs[2093] = layer0_outputs[1896];
    assign outputs[2094] = ~(layer0_outputs[1045]) | (layer0_outputs[2070]);
    assign outputs[2095] = ~((layer0_outputs[1170]) | (layer0_outputs[929]));
    assign outputs[2096] = ~(layer0_outputs[540]);
    assign outputs[2097] = ~((layer0_outputs[748]) | (layer0_outputs[1750]));
    assign outputs[2098] = (layer0_outputs[179]) & (layer0_outputs[2455]);
    assign outputs[2099] = ~(layer0_outputs[1130]);
    assign outputs[2100] = ~((layer0_outputs[1604]) ^ (layer0_outputs[2014]));
    assign outputs[2101] = ~(layer0_outputs[709]);
    assign outputs[2102] = ~((layer0_outputs[2123]) & (layer0_outputs[88]));
    assign outputs[2103] = (layer0_outputs[969]) & ~(layer0_outputs[2040]);
    assign outputs[2104] = (layer0_outputs[1920]) & (layer0_outputs[1160]);
    assign outputs[2105] = (layer0_outputs[1804]) ^ (layer0_outputs[1403]);
    assign outputs[2106] = ~(layer0_outputs[998]);
    assign outputs[2107] = ~((layer0_outputs[337]) ^ (layer0_outputs[2181]));
    assign outputs[2108] = layer0_outputs[185];
    assign outputs[2109] = ~((layer0_outputs[2106]) & (layer0_outputs[633]));
    assign outputs[2110] = (layer0_outputs[2351]) ^ (layer0_outputs[2238]);
    assign outputs[2111] = ~((layer0_outputs[495]) & (layer0_outputs[1729]));
    assign outputs[2112] = ~((layer0_outputs[1556]) & (layer0_outputs[397]));
    assign outputs[2113] = ~((layer0_outputs[2091]) ^ (layer0_outputs[698]));
    assign outputs[2114] = ~((layer0_outputs[1822]) ^ (layer0_outputs[861]));
    assign outputs[2115] = (layer0_outputs[196]) ^ (layer0_outputs[1184]);
    assign outputs[2116] = ~((layer0_outputs[548]) | (layer0_outputs[2256]));
    assign outputs[2117] = layer0_outputs[374];
    assign outputs[2118] = ~((layer0_outputs[2339]) & (layer0_outputs[535]));
    assign outputs[2119] = ~(layer0_outputs[544]);
    assign outputs[2120] = ~(layer0_outputs[1100]);
    assign outputs[2121] = layer0_outputs[1062];
    assign outputs[2122] = (layer0_outputs[1978]) ^ (layer0_outputs[1605]);
    assign outputs[2123] = ~(layer0_outputs[1567]) | (layer0_outputs[2375]);
    assign outputs[2124] = ~(layer0_outputs[2029]) | (layer0_outputs[1172]);
    assign outputs[2125] = ~(layer0_outputs[1942]) | (layer0_outputs[1540]);
    assign outputs[2126] = ~(layer0_outputs[1081]) | (layer0_outputs[519]);
    assign outputs[2127] = ~((layer0_outputs[457]) ^ (layer0_outputs[2342]));
    assign outputs[2128] = layer0_outputs[216];
    assign outputs[2129] = ~(layer0_outputs[676]) | (layer0_outputs[2287]);
    assign outputs[2130] = ~((layer0_outputs[522]) ^ (layer0_outputs[647]));
    assign outputs[2131] = layer0_outputs[837];
    assign outputs[2132] = (layer0_outputs[284]) & (layer0_outputs[2454]);
    assign outputs[2133] = (layer0_outputs[220]) ^ (layer0_outputs[1541]);
    assign outputs[2134] = layer0_outputs[417];
    assign outputs[2135] = ~(layer0_outputs[517]);
    assign outputs[2136] = (layer0_outputs[464]) ^ (layer0_outputs[2450]);
    assign outputs[2137] = (layer0_outputs[968]) & ~(layer0_outputs[1249]);
    assign outputs[2138] = ~(layer0_outputs[2139]);
    assign outputs[2139] = (layer0_outputs[2097]) | (layer0_outputs[451]);
    assign outputs[2140] = (layer0_outputs[1902]) ^ (layer0_outputs[768]);
    assign outputs[2141] = (layer0_outputs[0]) ^ (layer0_outputs[313]);
    assign outputs[2142] = (layer0_outputs[1248]) & (layer0_outputs[554]);
    assign outputs[2143] = ~(layer0_outputs[258]) | (layer0_outputs[1224]);
    assign outputs[2144] = (layer0_outputs[1881]) & ~(layer0_outputs[571]);
    assign outputs[2145] = 1'b1;
    assign outputs[2146] = (layer0_outputs[764]) & ~(layer0_outputs[878]);
    assign outputs[2147] = ~((layer0_outputs[711]) | (layer0_outputs[763]));
    assign outputs[2148] = (layer0_outputs[2131]) ^ (layer0_outputs[1237]);
    assign outputs[2149] = ~(layer0_outputs[854]);
    assign outputs[2150] = layer0_outputs[933];
    assign outputs[2151] = (layer0_outputs[85]) ^ (layer0_outputs[2103]);
    assign outputs[2152] = ~(layer0_outputs[134]);
    assign outputs[2153] = ~(layer0_outputs[1612]) | (layer0_outputs[1909]);
    assign outputs[2154] = (layer0_outputs[1051]) ^ (layer0_outputs[1944]);
    assign outputs[2155] = (layer0_outputs[1199]) ^ (layer0_outputs[481]);
    assign outputs[2156] = (layer0_outputs[1028]) | (layer0_outputs[2435]);
    assign outputs[2157] = (layer0_outputs[2132]) ^ (layer0_outputs[2339]);
    assign outputs[2158] = (layer0_outputs[3]) & ~(layer0_outputs[2036]);
    assign outputs[2159] = (layer0_outputs[1511]) & ~(layer0_outputs[140]);
    assign outputs[2160] = layer0_outputs[1792];
    assign outputs[2161] = ~((layer0_outputs[213]) | (layer0_outputs[1727]));
    assign outputs[2162] = (layer0_outputs[2226]) ^ (layer0_outputs[112]);
    assign outputs[2163] = layer0_outputs[1392];
    assign outputs[2164] = (layer0_outputs[1014]) ^ (layer0_outputs[532]);
    assign outputs[2165] = ~((layer0_outputs[270]) ^ (layer0_outputs[1501]));
    assign outputs[2166] = layer0_outputs[1910];
    assign outputs[2167] = (layer0_outputs[981]) ^ (layer0_outputs[1010]);
    assign outputs[2168] = layer0_outputs[1315];
    assign outputs[2169] = ~((layer0_outputs[1477]) ^ (layer0_outputs[2167]));
    assign outputs[2170] = ~(layer0_outputs[17]) | (layer0_outputs[13]);
    assign outputs[2171] = (layer0_outputs[72]) ^ (layer0_outputs[1634]);
    assign outputs[2172] = (layer0_outputs[1095]) | (layer0_outputs[405]);
    assign outputs[2173] = (layer0_outputs[2470]) & (layer0_outputs[1520]);
    assign outputs[2174] = layer0_outputs[1695];
    assign outputs[2175] = layer0_outputs[1106];
    assign outputs[2176] = ~(layer0_outputs[749]) | (layer0_outputs[1739]);
    assign outputs[2177] = (layer0_outputs[1738]) & ~(layer0_outputs[989]);
    assign outputs[2178] = (layer0_outputs[1370]) & (layer0_outputs[44]);
    assign outputs[2179] = ~((layer0_outputs[807]) & (layer0_outputs[92]));
    assign outputs[2180] = layer0_outputs[825];
    assign outputs[2181] = (layer0_outputs[2154]) ^ (layer0_outputs[808]);
    assign outputs[2182] = layer0_outputs[1119];
    assign outputs[2183] = layer0_outputs[2289];
    assign outputs[2184] = (layer0_outputs[2497]) ^ (layer0_outputs[431]);
    assign outputs[2185] = ~((layer0_outputs[2414]) ^ (layer0_outputs[211]));
    assign outputs[2186] = ~(layer0_outputs[1401]);
    assign outputs[2187] = ~((layer0_outputs[2194]) & (layer0_outputs[2473]));
    assign outputs[2188] = (layer0_outputs[2001]) ^ (layer0_outputs[435]);
    assign outputs[2189] = ~((layer0_outputs[2492]) & (layer0_outputs[7]));
    assign outputs[2190] = (layer0_outputs[1491]) ^ (layer0_outputs[844]);
    assign outputs[2191] = (layer0_outputs[1917]) ^ (layer0_outputs[524]);
    assign outputs[2192] = ~(layer0_outputs[780]) | (layer0_outputs[1086]);
    assign outputs[2193] = (layer0_outputs[970]) & ~(layer0_outputs[1212]);
    assign outputs[2194] = (layer0_outputs[466]) ^ (layer0_outputs[177]);
    assign outputs[2195] = layer0_outputs[18];
    assign outputs[2196] = (layer0_outputs[798]) ^ (layer0_outputs[594]);
    assign outputs[2197] = ~((layer0_outputs[665]) | (layer0_outputs[791]));
    assign outputs[2198] = ~(layer0_outputs[1486]);
    assign outputs[2199] = ~((layer0_outputs[1892]) ^ (layer0_outputs[2134]));
    assign outputs[2200] = 1'b1;
    assign outputs[2201] = (layer0_outputs[1664]) ^ (layer0_outputs[126]);
    assign outputs[2202] = ~((layer0_outputs[1382]) & (layer0_outputs[1532]));
    assign outputs[2203] = ~((layer0_outputs[1663]) ^ (layer0_outputs[2388]));
    assign outputs[2204] = (layer0_outputs[1504]) & ~(layer0_outputs[120]);
    assign outputs[2205] = layer0_outputs[2011];
    assign outputs[2206] = (layer0_outputs[2268]) | (layer0_outputs[1077]);
    assign outputs[2207] = ~((layer0_outputs[1339]) ^ (layer0_outputs[906]));
    assign outputs[2208] = ~(layer0_outputs[517]) | (layer0_outputs[1622]);
    assign outputs[2209] = (layer0_outputs[1204]) ^ (layer0_outputs[859]);
    assign outputs[2210] = (layer0_outputs[1407]) | (layer0_outputs[1897]);
    assign outputs[2211] = layer0_outputs[2195];
    assign outputs[2212] = ~((layer0_outputs[2440]) & (layer0_outputs[1862]));
    assign outputs[2213] = layer0_outputs[1799];
    assign outputs[2214] = (layer0_outputs[1214]) & ~(layer0_outputs[642]);
    assign outputs[2215] = (layer0_outputs[86]) ^ (layer0_outputs[326]);
    assign outputs[2216] = ~(layer0_outputs[402]);
    assign outputs[2217] = ~(layer0_outputs[728]);
    assign outputs[2218] = (layer0_outputs[2281]) & ~(layer0_outputs[16]);
    assign outputs[2219] = ~((layer0_outputs[151]) & (layer0_outputs[1890]));
    assign outputs[2220] = (layer0_outputs[2374]) ^ (layer0_outputs[1322]);
    assign outputs[2221] = layer0_outputs[768];
    assign outputs[2222] = ~((layer0_outputs[1073]) & (layer0_outputs[314]));
    assign outputs[2223] = ~(layer0_outputs[2310]) | (layer0_outputs[700]);
    assign outputs[2224] = layer0_outputs[991];
    assign outputs[2225] = (layer0_outputs[765]) | (layer0_outputs[1171]);
    assign outputs[2226] = layer0_outputs[198];
    assign outputs[2227] = ~(layer0_outputs[2327]) | (layer0_outputs[759]);
    assign outputs[2228] = (layer0_outputs[1408]) & ~(layer0_outputs[750]);
    assign outputs[2229] = ~((layer0_outputs[2186]) ^ (layer0_outputs[1271]));
    assign outputs[2230] = ~((layer0_outputs[772]) ^ (layer0_outputs[1306]));
    assign outputs[2231] = layer0_outputs[1992];
    assign outputs[2232] = (layer0_outputs[144]) ^ (layer0_outputs[1710]);
    assign outputs[2233] = layer0_outputs[1741];
    assign outputs[2234] = ~(layer0_outputs[1484]);
    assign outputs[2235] = ~((layer0_outputs[2392]) ^ (layer0_outputs[193]));
    assign outputs[2236] = ~(layer0_outputs[462]);
    assign outputs[2237] = layer0_outputs[179];
    assign outputs[2238] = (layer0_outputs[361]) | (layer0_outputs[2214]);
    assign outputs[2239] = (layer0_outputs[1815]) & ~(layer0_outputs[926]);
    assign outputs[2240] = ~(layer0_outputs[1777]);
    assign outputs[2241] = layer0_outputs[1356];
    assign outputs[2242] = (layer0_outputs[1270]) | (layer0_outputs[1646]);
    assign outputs[2243] = ~((layer0_outputs[327]) & (layer0_outputs[2264]));
    assign outputs[2244] = ~(layer0_outputs[1025]) | (layer0_outputs[741]);
    assign outputs[2245] = ~(layer0_outputs[1609]);
    assign outputs[2246] = ~(layer0_outputs[495]);
    assign outputs[2247] = ~(layer0_outputs[1503]) | (layer0_outputs[2467]);
    assign outputs[2248] = ~(layer0_outputs[1765]);
    assign outputs[2249] = (layer0_outputs[672]) & ~(layer0_outputs[1355]);
    assign outputs[2250] = ~(layer0_outputs[948]);
    assign outputs[2251] = (layer0_outputs[1769]) & (layer0_outputs[46]);
    assign outputs[2252] = (layer0_outputs[1092]) & (layer0_outputs[863]);
    assign outputs[2253] = (layer0_outputs[2350]) ^ (layer0_outputs[1955]);
    assign outputs[2254] = ~(layer0_outputs[888]);
    assign outputs[2255] = ~(layer0_outputs[1706]);
    assign outputs[2256] = ~((layer0_outputs[1783]) ^ (layer0_outputs[978]));
    assign outputs[2257] = (layer0_outputs[135]) & (layer0_outputs[1708]);
    assign outputs[2258] = layer0_outputs[1965];
    assign outputs[2259] = (layer0_outputs[2170]) & ~(layer0_outputs[2233]);
    assign outputs[2260] = ~((layer0_outputs[176]) & (layer0_outputs[1733]));
    assign outputs[2261] = layer0_outputs[1534];
    assign outputs[2262] = ~((layer0_outputs[1999]) | (layer0_outputs[370]));
    assign outputs[2263] = ~((layer0_outputs[241]) & (layer0_outputs[970]));
    assign outputs[2264] = (layer0_outputs[2203]) & (layer0_outputs[2432]);
    assign outputs[2265] = ~(layer0_outputs[29]);
    assign outputs[2266] = layer0_outputs[2059];
    assign outputs[2267] = layer0_outputs[2111];
    assign outputs[2268] = layer0_outputs[2043];
    assign outputs[2269] = (layer0_outputs[2144]) & ~(layer0_outputs[674]);
    assign outputs[2270] = layer0_outputs[1763];
    assign outputs[2271] = ~((layer0_outputs[62]) | (layer0_outputs[1805]));
    assign outputs[2272] = layer0_outputs[1674];
    assign outputs[2273] = layer0_outputs[588];
    assign outputs[2274] = ~((layer0_outputs[326]) | (layer0_outputs[2055]));
    assign outputs[2275] = (layer0_outputs[793]) | (layer0_outputs[1281]);
    assign outputs[2276] = layer0_outputs[608];
    assign outputs[2277] = ~(layer0_outputs[1698]);
    assign outputs[2278] = ~(layer0_outputs[712]);
    assign outputs[2279] = ~((layer0_outputs[24]) & (layer0_outputs[992]));
    assign outputs[2280] = (layer0_outputs[2231]) & ~(layer0_outputs[1453]);
    assign outputs[2281] = (layer0_outputs[2038]) & (layer0_outputs[919]);
    assign outputs[2282] = layer0_outputs[1420];
    assign outputs[2283] = (layer0_outputs[286]) | (layer0_outputs[909]);
    assign outputs[2284] = ~((layer0_outputs[1220]) | (layer0_outputs[76]));
    assign outputs[2285] = (layer0_outputs[1888]) & ~(layer0_outputs[1206]);
    assign outputs[2286] = (layer0_outputs[1387]) ^ (layer0_outputs[1267]);
    assign outputs[2287] = ~((layer0_outputs[751]) ^ (layer0_outputs[87]));
    assign outputs[2288] = ~(layer0_outputs[2158]);
    assign outputs[2289] = ~(layer0_outputs[1592]);
    assign outputs[2290] = ~(layer0_outputs[1170]);
    assign outputs[2291] = (layer0_outputs[1513]) & ~(layer0_outputs[356]);
    assign outputs[2292] = (layer0_outputs[61]) ^ (layer0_outputs[2354]);
    assign outputs[2293] = ~(layer0_outputs[26]) | (layer0_outputs[1141]);
    assign outputs[2294] = (layer0_outputs[600]) & ~(layer0_outputs[2388]);
    assign outputs[2295] = (layer0_outputs[2002]) & ~(layer0_outputs[677]);
    assign outputs[2296] = (layer0_outputs[1035]) | (layer0_outputs[636]);
    assign outputs[2297] = layer0_outputs[351];
    assign outputs[2298] = layer0_outputs[1682];
    assign outputs[2299] = ~(layer0_outputs[2136]);
    assign outputs[2300] = layer0_outputs[887];
    assign outputs[2301] = layer0_outputs[662];
    assign outputs[2302] = layer0_outputs[956];
    assign outputs[2303] = ~(layer0_outputs[1785]);
    assign outputs[2304] = (layer0_outputs[1867]) & (layer0_outputs[832]);
    assign outputs[2305] = ~((layer0_outputs[2330]) ^ (layer0_outputs[1640]));
    assign outputs[2306] = layer0_outputs[2167];
    assign outputs[2307] = ~(layer0_outputs[50]) | (layer0_outputs[636]);
    assign outputs[2308] = ~((layer0_outputs[576]) ^ (layer0_outputs[953]));
    assign outputs[2309] = (layer0_outputs[1997]) & ~(layer0_outputs[41]);
    assign outputs[2310] = (layer0_outputs[687]) & ~(layer0_outputs[319]);
    assign outputs[2311] = ~((layer0_outputs[2270]) & (layer0_outputs[1321]));
    assign outputs[2312] = ~((layer0_outputs[1097]) ^ (layer0_outputs[1639]));
    assign outputs[2313] = ~(layer0_outputs[2377]);
    assign outputs[2314] = ~(layer0_outputs[292]);
    assign outputs[2315] = ~(layer0_outputs[1231]);
    assign outputs[2316] = (layer0_outputs[1029]) | (layer0_outputs[2201]);
    assign outputs[2317] = (layer0_outputs[1252]) & ~(layer0_outputs[1181]);
    assign outputs[2318] = layer0_outputs[1055];
    assign outputs[2319] = ~(layer0_outputs[345]);
    assign outputs[2320] = (layer0_outputs[820]) ^ (layer0_outputs[235]);
    assign outputs[2321] = ~((layer0_outputs[2198]) | (layer0_outputs[690]));
    assign outputs[2322] = ~((layer0_outputs[1423]) ^ (layer0_outputs[1595]));
    assign outputs[2323] = ~(layer0_outputs[765]);
    assign outputs[2324] = (layer0_outputs[726]) & ~(layer0_outputs[183]);
    assign outputs[2325] = layer0_outputs[724];
    assign outputs[2326] = ~(layer0_outputs[188]);
    assign outputs[2327] = ~((layer0_outputs[36]) ^ (layer0_outputs[384]));
    assign outputs[2328] = (layer0_outputs[418]) & (layer0_outputs[1050]);
    assign outputs[2329] = layer0_outputs[1809];
    assign outputs[2330] = ~((layer0_outputs[2405]) ^ (layer0_outputs[1636]));
    assign outputs[2331] = (layer0_outputs[1273]) & ~(layer0_outputs[1012]);
    assign outputs[2332] = ~(layer0_outputs[650]);
    assign outputs[2333] = (layer0_outputs[443]) ^ (layer0_outputs[298]);
    assign outputs[2334] = ~(layer0_outputs[216]);
    assign outputs[2335] = ~(layer0_outputs[77]);
    assign outputs[2336] = (layer0_outputs[1187]) & ~(layer0_outputs[1528]);
    assign outputs[2337] = ~(layer0_outputs[2478]);
    assign outputs[2338] = (layer0_outputs[619]) | (layer0_outputs[908]);
    assign outputs[2339] = ~((layer0_outputs[319]) | (layer0_outputs[2421]));
    assign outputs[2340] = ~(layer0_outputs[1309]);
    assign outputs[2341] = ~(layer0_outputs[488]);
    assign outputs[2342] = (layer0_outputs[963]) & ~(layer0_outputs[2163]);
    assign outputs[2343] = (layer0_outputs[824]) & ~(layer0_outputs[591]);
    assign outputs[2344] = (layer0_outputs[2105]) ^ (layer0_outputs[2331]);
    assign outputs[2345] = (layer0_outputs[2251]) & ~(layer0_outputs[1970]);
    assign outputs[2346] = ~(layer0_outputs[1177]);
    assign outputs[2347] = ~((layer0_outputs[659]) | (layer0_outputs[1351]));
    assign outputs[2348] = (layer0_outputs[2212]) & (layer0_outputs[2384]);
    assign outputs[2349] = layer0_outputs[770];
    assign outputs[2350] = ~((layer0_outputs[753]) | (layer0_outputs[1699]));
    assign outputs[2351] = (layer0_outputs[1486]) & (layer0_outputs[1901]);
    assign outputs[2352] = (layer0_outputs[1893]) & ~(layer0_outputs[306]);
    assign outputs[2353] = ~((layer0_outputs[650]) | (layer0_outputs[1325]));
    assign outputs[2354] = layer0_outputs[2387];
    assign outputs[2355] = ~((layer0_outputs[57]) | (layer0_outputs[2032]));
    assign outputs[2356] = (layer0_outputs[1495]) & ~(layer0_outputs[1889]);
    assign outputs[2357] = (layer0_outputs[1864]) ^ (layer0_outputs[1070]);
    assign outputs[2358] = (layer0_outputs[695]) & ~(layer0_outputs[221]);
    assign outputs[2359] = (layer0_outputs[1772]) & (layer0_outputs[199]);
    assign outputs[2360] = ~((layer0_outputs[1094]) | (layer0_outputs[1475]));
    assign outputs[2361] = (layer0_outputs[2367]) & (layer0_outputs[2244]);
    assign outputs[2362] = layer0_outputs[1649];
    assign outputs[2363] = (layer0_outputs[1691]) & ~(layer0_outputs[2005]);
    assign outputs[2364] = ~((layer0_outputs[2150]) | (layer0_outputs[1104]));
    assign outputs[2365] = (layer0_outputs[1176]) | (layer0_outputs[1542]);
    assign outputs[2366] = ~((layer0_outputs[2027]) ^ (layer0_outputs[815]));
    assign outputs[2367] = (layer0_outputs[1817]) & ~(layer0_outputs[369]);
    assign outputs[2368] = ~((layer0_outputs[714]) | (layer0_outputs[1144]));
    assign outputs[2369] = ~(layer0_outputs[39]);
    assign outputs[2370] = ~((layer0_outputs[1705]) ^ (layer0_outputs[1124]));
    assign outputs[2371] = ~((layer0_outputs[1299]) | (layer0_outputs[388]));
    assign outputs[2372] = (layer0_outputs[1523]) & ~(layer0_outputs[1506]);
    assign outputs[2373] = layer0_outputs[982];
    assign outputs[2374] = (layer0_outputs[1363]) | (layer0_outputs[2414]);
    assign outputs[2375] = ~(layer0_outputs[1506]);
    assign outputs[2376] = ~(layer0_outputs[1444]);
    assign outputs[2377] = (layer0_outputs[1]) & (layer0_outputs[1108]);
    assign outputs[2378] = (layer0_outputs[100]) | (layer0_outputs[938]);
    assign outputs[2379] = (layer0_outputs[2052]) & (layer0_outputs[1277]);
    assign outputs[2380] = (layer0_outputs[1597]) | (layer0_outputs[686]);
    assign outputs[2381] = (layer0_outputs[2467]) & ~(layer0_outputs[1008]);
    assign outputs[2382] = ~(layer0_outputs[139]) | (layer0_outputs[1479]);
    assign outputs[2383] = (layer0_outputs[1474]) & ~(layer0_outputs[749]);
    assign outputs[2384] = (layer0_outputs[1127]) & ~(layer0_outputs[1259]);
    assign outputs[2385] = ~((layer0_outputs[1524]) & (layer0_outputs[2123]));
    assign outputs[2386] = (layer0_outputs[1395]) & ~(layer0_outputs[1839]);
    assign outputs[2387] = layer0_outputs[982];
    assign outputs[2388] = ~(layer0_outputs[2428]);
    assign outputs[2389] = ~((layer0_outputs[2433]) ^ (layer0_outputs[1512]));
    assign outputs[2390] = (layer0_outputs[2234]) & ~(layer0_outputs[2469]);
    assign outputs[2391] = (layer0_outputs[2313]) & (layer0_outputs[491]);
    assign outputs[2392] = ~(layer0_outputs[718]);
    assign outputs[2393] = (layer0_outputs[624]) | (layer0_outputs[2121]);
    assign outputs[2394] = ~(layer0_outputs[1148]);
    assign outputs[2395] = (layer0_outputs[1871]) & ~(layer0_outputs[2254]);
    assign outputs[2396] = ~(layer0_outputs[1844]);
    assign outputs[2397] = ~((layer0_outputs[1510]) ^ (layer0_outputs[2000]));
    assign outputs[2398] = (layer0_outputs[1761]) & ~(layer0_outputs[1245]);
    assign outputs[2399] = ~((layer0_outputs[1262]) | (layer0_outputs[91]));
    assign outputs[2400] = (layer0_outputs[551]) | (layer0_outputs[2221]);
    assign outputs[2401] = (layer0_outputs[393]) & (layer0_outputs[1860]);
    assign outputs[2402] = (layer0_outputs[428]) & (layer0_outputs[454]);
    assign outputs[2403] = ~(layer0_outputs[2165]);
    assign outputs[2404] = (layer0_outputs[2153]) & ~(layer0_outputs[1430]);
    assign outputs[2405] = (layer0_outputs[1079]) ^ (layer0_outputs[1385]);
    assign outputs[2406] = ~((layer0_outputs[297]) ^ (layer0_outputs[644]));
    assign outputs[2407] = (layer0_outputs[1158]) & ~(layer0_outputs[787]);
    assign outputs[2408] = layer0_outputs[769];
    assign outputs[2409] = layer0_outputs[783];
    assign outputs[2410] = ~(layer0_outputs[488]);
    assign outputs[2411] = ~(layer0_outputs[260]);
    assign outputs[2412] = ~((layer0_outputs[1253]) ^ (layer0_outputs[1498]));
    assign outputs[2413] = ~((layer0_outputs[669]) | (layer0_outputs[336]));
    assign outputs[2414] = ~((layer0_outputs[512]) & (layer0_outputs[1581]));
    assign outputs[2415] = ~(layer0_outputs[932]);
    assign outputs[2416] = ~(layer0_outputs[2277]) | (layer0_outputs[1063]);
    assign outputs[2417] = (layer0_outputs[519]) | (layer0_outputs[390]);
    assign outputs[2418] = ~((layer0_outputs[757]) ^ (layer0_outputs[1311]));
    assign outputs[2419] = layer0_outputs[439];
    assign outputs[2420] = ~((layer0_outputs[643]) ^ (layer0_outputs[434]));
    assign outputs[2421] = (layer0_outputs[884]) & ~(layer0_outputs[868]);
    assign outputs[2422] = (layer0_outputs[2088]) & ~(layer0_outputs[2417]);
    assign outputs[2423] = (layer0_outputs[558]) & ~(layer0_outputs[944]);
    assign outputs[2424] = ~((layer0_outputs[1533]) & (layer0_outputs[754]));
    assign outputs[2425] = ~(layer0_outputs[894]);
    assign outputs[2426] = ~((layer0_outputs[784]) ^ (layer0_outputs[1639]));
    assign outputs[2427] = (layer0_outputs[1258]) & (layer0_outputs[1463]);
    assign outputs[2428] = (layer0_outputs[2346]) | (layer0_outputs[1105]);
    assign outputs[2429] = (layer0_outputs[2181]) & ~(layer0_outputs[1103]);
    assign outputs[2430] = (layer0_outputs[2138]) & ~(layer0_outputs[1166]);
    assign outputs[2431] = (layer0_outputs[1308]) & ~(layer0_outputs[423]);
    assign outputs[2432] = layer0_outputs[468];
    assign outputs[2433] = ~((layer0_outputs[2003]) ^ (layer0_outputs[227]));
    assign outputs[2434] = (layer0_outputs[2039]) & (layer0_outputs[392]);
    assign outputs[2435] = (layer0_outputs[162]) & ~(layer0_outputs[168]);
    assign outputs[2436] = layer0_outputs[1677];
    assign outputs[2437] = (layer0_outputs[2185]) | (layer0_outputs[426]);
    assign outputs[2438] = ~(layer0_outputs[77]);
    assign outputs[2439] = (layer0_outputs[252]) ^ (layer0_outputs[937]);
    assign outputs[2440] = (layer0_outputs[482]) & ~(layer0_outputs[2294]);
    assign outputs[2441] = (layer0_outputs[1489]) | (layer0_outputs[1343]);
    assign outputs[2442] = ~(layer0_outputs[1293]);
    assign outputs[2443] = ~((layer0_outputs[922]) & (layer0_outputs[2416]));
    assign outputs[2444] = ~((layer0_outputs[1675]) ^ (layer0_outputs[2124]));
    assign outputs[2445] = layer0_outputs[1459];
    assign outputs[2446] = layer0_outputs[248];
    assign outputs[2447] = layer0_outputs[1987];
    assign outputs[2448] = (layer0_outputs[2217]) & ~(layer0_outputs[2023]);
    assign outputs[2449] = ~((layer0_outputs[1295]) & (layer0_outputs[1978]));
    assign outputs[2450] = (layer0_outputs[1405]) ^ (layer0_outputs[2161]);
    assign outputs[2451] = (layer0_outputs[1707]) ^ (layer0_outputs[2401]);
    assign outputs[2452] = (layer0_outputs[217]) & ~(layer0_outputs[26]);
    assign outputs[2453] = ~(layer0_outputs[1042]) | (layer0_outputs[925]);
    assign outputs[2454] = (layer0_outputs[2496]) & (layer0_outputs[1242]);
    assign outputs[2455] = ~((layer0_outputs[1957]) ^ (layer0_outputs[1607]));
    assign outputs[2456] = ~((layer0_outputs[1090]) ^ (layer0_outputs[2073]));
    assign outputs[2457] = (layer0_outputs[2354]) ^ (layer0_outputs[2041]);
    assign outputs[2458] = (layer0_outputs[2378]) & (layer0_outputs[2461]);
    assign outputs[2459] = ~((layer0_outputs[2113]) & (layer0_outputs[1155]));
    assign outputs[2460] = ~(layer0_outputs[1231]) | (layer0_outputs[909]);
    assign outputs[2461] = ~((layer0_outputs[1810]) ^ (layer0_outputs[195]));
    assign outputs[2462] = (layer0_outputs[1654]) & ~(layer0_outputs[299]);
    assign outputs[2463] = layer0_outputs[850];
    assign outputs[2464] = (layer0_outputs[908]) & ~(layer0_outputs[2486]);
    assign outputs[2465] = (layer0_outputs[2216]) & ~(layer0_outputs[441]);
    assign outputs[2466] = (layer0_outputs[898]) & ~(layer0_outputs[175]);
    assign outputs[2467] = ~((layer0_outputs[1516]) ^ (layer0_outputs[49]));
    assign outputs[2468] = ~(layer0_outputs[1103]) | (layer0_outputs[1893]);
    assign outputs[2469] = layer0_outputs[2288];
    assign outputs[2470] = ~((layer0_outputs[2120]) ^ (layer0_outputs[2228]));
    assign outputs[2471] = (layer0_outputs[711]) ^ (layer0_outputs[906]);
    assign outputs[2472] = layer0_outputs[1349];
    assign outputs[2473] = ~(layer0_outputs[1911]) | (layer0_outputs[565]);
    assign outputs[2474] = (layer0_outputs[2172]) & ~(layer0_outputs[82]);
    assign outputs[2475] = (layer0_outputs[285]) & (layer0_outputs[402]);
    assign outputs[2476] = ~(layer0_outputs[1567]);
    assign outputs[2477] = layer0_outputs[406];
    assign outputs[2478] = ~((layer0_outputs[797]) | (layer0_outputs[508]));
    assign outputs[2479] = ~((layer0_outputs[569]) ^ (layer0_outputs[1741]));
    assign outputs[2480] = ~(layer0_outputs[481]) | (layer0_outputs[167]);
    assign outputs[2481] = (layer0_outputs[597]) & ~(layer0_outputs[1469]);
    assign outputs[2482] = ~(layer0_outputs[652]);
    assign outputs[2483] = ~((layer0_outputs[2209]) | (layer0_outputs[2409]));
    assign outputs[2484] = ~((layer0_outputs[717]) | (layer0_outputs[1291]));
    assign outputs[2485] = layer0_outputs[976];
    assign outputs[2486] = layer0_outputs[1648];
    assign outputs[2487] = ~(layer0_outputs[1521]);
    assign outputs[2488] = layer0_outputs[578];
    assign outputs[2489] = layer0_outputs[15];
    assign outputs[2490] = ~(layer0_outputs[1593]);
    assign outputs[2491] = ~(layer0_outputs[356]);
    assign outputs[2492] = (layer0_outputs[1773]) ^ (layer0_outputs[471]);
    assign outputs[2493] = layer0_outputs[2230];
    assign outputs[2494] = (layer0_outputs[1653]) & ~(layer0_outputs[411]);
    assign outputs[2495] = (layer0_outputs[190]) | (layer0_outputs[2009]);
    assign outputs[2496] = (layer0_outputs[2415]) & ~(layer0_outputs[444]);
    assign outputs[2497] = ~((layer0_outputs[2089]) & (layer0_outputs[2049]));
    assign outputs[2498] = (layer0_outputs[1314]) & ~(layer0_outputs[537]);
    assign outputs[2499] = ~((layer0_outputs[535]) | (layer0_outputs[1655]));
	 
	 // Sum and argmax logic
	 reg [9:0] sums [0:9];                     // Array to store sums for each group of 250 bits
    reg [9:0] max_sum;                        // Variable for the maximum sum
    reg [3:0] max_index;                      // 4-bit output for index of maximum sum (0 to 9)
    integer i, j;
	 
    always @* begin
        // Initialize sums
        for (i = 0; i < 10; i = i + 1) begin
            sums[i] = 0; // Reset each sum to 0
        end

        // Sum each group of 250 bits in outputs
        for (i = 0; i < 10; i = i + 1) begin
            for (j = 0; j < 250; j = j + 1) begin
                sums[i] = sums[i] + outputs[i * 250 + j]; // Sum the elements in each group
            end
        end

        // Find argmax
        max_index = 0;
        max_sum = sums[0];
        for (i = 1; i < 10; i = i + 1) begin
            if (sums[i] > max_sum) begin
                max_sum = sums[i];
                max_index = i;
            end
        end
		  
		  // Generate one-hot encoding for classification
        classification = 10'b0; // Reset classification
        classification[max_index] = 1'b1; // Set the corresponding index to 1
    end
	 
endmodule
